module SPEEDY_Rounds6_0 ( Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  wire   \RI1[1][179] , \RI1[1][149] , \RI1[1][47] , \RI1[1][23] ,
         \RI1[1][11] , \RI1[2][191] , \RI1[2][185] , \RI1[2][149] ,
         \RI1[2][125] , \RI1[2][119] , \RI1[2][116] , \RI1[2][107] ,
         \RI1[2][101] , \RI1[2][59] , \RI1[2][17] , \RI1[2][9] , \RI1[2][5] ,
         \RI1[3][191] , \RI1[3][167] , \RI1[3][165] , \RI1[3][161] ,
         \RI1[3][107] , \RI1[3][101] , \RI1[3][17] , \RI1[3][5] ,
         \RI1[4][191] , \RI1[4][173] , \RI1[4][155] , \RI1[4][141] ,
         \RI1[4][140] , \RI1[4][131] , \RI1[4][119] , \RI1[4][105] ,
         \RI1[4][65] , \RI1[4][59] , \RI1[4][53] , \RI1[4][41] , \RI1[4][26] ,
         \RI1[4][17] , \RI1[4][5] , \RI1[5][185] , \RI1[5][179] ,
         \RI1[5][173] , \RI1[5][167] , \RI1[5][155] , \RI1[5][137] ,
         \RI1[5][119] , \RI1[5][113] , \RI1[5][107] , \RI1[5][89] ,
         \RI1[5][80] , \RI1[5][77] , \RI1[5][59] , \RI1[5][53] , \RI1[5][41] ,
         \RI1[5][35] , \RI1[5][17] , \RI1[5][11] , \RI3[0][190] ,
         \RI3[0][189] , \RI3[0][188] , \RI3[0][187] , \RI3[0][184] ,
         \RI3[0][183] , \RI3[0][182] , \RI3[0][179] , \RI3[0][178] ,
         \RI3[0][177] , \RI3[0][176] , \RI3[0][175] , \RI3[0][174] ,
         \RI3[0][173] , \RI3[0][172] , \RI3[0][171] , \RI3[0][170] ,
         \RI3[0][169] , \RI3[0][167] , \RI3[0][166] , \RI3[0][163] ,
         \RI3[0][158] , \RI3[0][155] , \RI3[0][154] , \RI3[0][153] ,
         \RI3[0][152] , \RI3[0][151] , \RI3[0][150] , \RI3[0][149] ,
         \RI3[0][148] , \RI3[0][147] , \RI3[0][144] , \RI3[0][143] ,
         \RI3[0][142] , \RI3[0][141] , \RI3[0][140] , \RI3[0][139] ,
         \RI3[0][136] , \RI3[0][133] , \RI3[0][131] , \RI3[0][129] ,
         \RI3[0][128] , \RI3[0][127] , \RI3[0][126] , \RI3[0][125] ,
         \RI3[0][123] , \RI3[0][122] , \RI3[0][121] , \RI3[0][120] ,
         \RI3[0][119] , \RI3[0][118] , \RI3[0][117] , \RI3[0][116] ,
         \RI3[0][115] , \RI3[0][114] , \RI3[0][113] , \RI3[0][112] ,
         \RI3[0][111] , \RI3[0][110] , \RI3[0][109] , \RI3[0][101] ,
         \RI3[0][100] , \RI3[0][99] , \RI3[0][97] , \RI3[0][96] , \RI3[0][95] ,
         \RI3[0][93] , \RI3[0][91] , \RI3[0][90] , \RI3[0][89] , \RI3[0][88] ,
         \RI3[0][87] , \RI3[0][86] , \RI3[0][83] , \RI3[0][82] , \RI3[0][81] ,
         \RI3[0][78] , \RI3[0][77] , \RI3[0][76] , \RI3[0][75] , \RI3[0][72] ,
         \RI3[0][71] , \RI3[0][70] , \RI3[0][68] , \RI3[0][67] , \RI3[0][65] ,
         \RI3[0][63] , \RI3[0][62] , \RI3[0][60] , \RI3[0][58] , \RI3[0][57] ,
         \RI3[0][56] , \RI3[0][55] , \RI3[0][53] , \RI3[0][52] , \RI3[0][50] ,
         \RI3[0][49] , \RI3[0][47] , \RI3[0][46] , \RI3[0][44] , \RI3[0][42] ,
         \RI3[0][41] , \RI3[0][39] , \RI3[0][38] , \RI3[0][35] , \RI3[0][33] ,
         \RI3[0][30] , \RI3[0][29] , \RI3[0][28] , \RI3[0][27] , \RI3[0][21] ,
         \RI3[0][19] , \RI3[0][18] , \RI3[0][15] , \RI3[0][10] , \RI3[0][9] ,
         \RI3[0][8] , \RI3[0][5] , \RI3[0][4] , \RI3[0][3] , \RI3[0][1] ,
         \RI3[0][0] , \RI3[1][152] , \RI3[1][111] , \RI3[1][26] ,
         \RI3[2][131] , \RI3[2][121] , \RI3[2][97] , \RI3[2][95] ,
         \RI3[2][88] , \RI3[3][70] , \RI3[3][64] , \RI3[3][58] , \RI3[4][188] ,
         \RI3[4][148] , \RI3[4][127] , \RI3[5][171] , \RI3[5][149] ,
         \RI3[5][128] , \RI3[5][73] , \RI5[0][191] , \RI5[0][190] ,
         \RI5[0][189] , \RI5[0][188] , \RI5[0][187] , \RI5[0][186] ,
         \RI5[0][185] , \RI5[0][184] , \RI5[0][183] , \RI5[0][182] ,
         \RI5[0][181] , \RI5[0][180] , \RI5[0][179] , \RI5[0][178] ,
         \RI5[0][177] , \RI5[0][176] , \RI5[0][175] , \RI5[0][174] ,
         \RI5[0][173] , \RI5[0][172] , \RI5[0][171] , \RI5[0][170] ,
         \RI5[0][169] , \RI5[0][168] , \RI5[0][167] , \RI5[0][166] ,
         \RI5[0][165] , \RI5[0][164] , \RI5[0][163] , \RI5[0][162] ,
         \RI5[0][161] , \RI5[0][160] , \RI5[0][159] , \RI5[0][158] ,
         \RI5[0][157] , \RI5[0][156] , \RI5[0][155] , \RI5[0][154] ,
         \RI5[0][153] , \RI5[0][152] , \RI5[0][151] , \RI5[0][150] ,
         \RI5[0][149] , \RI5[0][148] , \RI5[0][147] , \RI5[0][146] ,
         \RI5[0][145] , \RI5[0][144] , \RI5[0][143] , \RI5[0][142] ,
         \RI5[0][141] , \RI5[0][140] , \RI5[0][138] , \RI5[0][136] ,
         \RI5[0][135] , \RI5[0][134] , \RI5[0][133] , \RI5[0][132] ,
         \RI5[0][131] , \RI5[0][130] , \RI5[0][129] , \RI5[0][128] ,
         \RI5[0][127] , \RI5[0][126] , \RI5[0][125] , \RI5[0][124] ,
         \RI5[0][123] , \RI5[0][122] , \RI5[0][121] , \RI5[0][120] ,
         \RI5[0][119] , \RI5[0][118] , \RI5[0][117] , \RI5[0][116] ,
         \RI5[0][115] , \RI5[0][114] , \RI5[0][112] , \RI5[0][111] ,
         \RI5[0][110] , \RI5[0][109] , \RI5[0][107] , \RI5[0][106] ,
         \RI5[0][105] , \RI5[0][104] , \RI5[0][103] , \RI5[0][101] ,
         \RI5[0][100] , \RI5[0][99] , \RI5[0][98] , \RI5[0][96] , \RI5[0][95] ,
         \RI5[0][94] , \RI5[0][93] , \RI5[0][92] , \RI5[0][91] , \RI5[0][90] ,
         \RI5[0][89] , \RI5[0][88] , \RI5[0][87] , \RI5[0][86] , \RI5[0][85] ,
         \RI5[0][83] , \RI5[0][82] , \RI5[0][81] , \RI5[0][80] , \RI5[0][79] ,
         \RI5[0][78] , \RI5[0][76] , \RI5[0][74] , \RI5[0][73] , \RI5[0][72] ,
         \RI5[0][69] , \RI5[0][68] , \RI5[0][66] , \RI5[0][65] , \RI5[0][63] ,
         \RI5[0][62] , \RI5[0][61] , \RI5[0][60] , \RI5[0][59] , \RI5[0][58] ,
         \RI5[0][57] , \RI5[0][56] , \RI5[0][55] , \RI5[0][54] , \RI5[0][53] ,
         \RI5[0][52] , \RI5[0][51] , \RI5[0][50] , \RI5[0][49] , \RI5[0][48] ,
         \RI5[0][47] , \RI5[0][46] , \RI5[0][45] , \RI5[0][44] , \RI5[0][42] ,
         \RI5[0][40] , \RI5[0][39] , \RI5[0][38] , \RI5[0][37] , \RI5[0][36] ,
         \RI5[0][34] , \RI5[0][33] , \RI5[0][32] , \RI5[0][30] , \RI5[0][29] ,
         \RI5[0][28] , \RI5[0][27] , \RI5[0][26] , \RI5[0][25] , \RI5[0][24] ,
         \RI5[0][23] , \RI5[0][22] , \RI5[0][21] , \RI5[0][20] , \RI5[0][19] ,
         \RI5[0][18] , \RI5[0][17] , \RI5[0][16] , \RI5[0][15] , \RI5[0][14] ,
         \RI5[0][13] , \RI5[0][12] , \RI5[0][11] , \RI5[0][10] , \RI5[0][9] ,
         \RI5[0][8] , \RI5[0][7] , \RI5[0][6] , \RI5[0][5] , \RI5[0][4] ,
         \RI5[0][3] , \RI5[0][2] , \RI5[0][1] , \RI5[0][0] , \RI5[1][191] ,
         \RI5[1][190] , \RI5[1][186] , \RI5[1][185] , \RI5[1][184] ,
         \RI5[1][183] , \RI5[1][181] , \RI5[1][180] , \RI5[1][179] ,
         \RI5[1][176] , \RI5[1][175] , \RI5[1][174] , \RI5[1][173] ,
         \RI5[1][171] , \RI5[1][170] , \RI5[1][169] , \RI5[1][167] ,
         \RI5[1][166] , \RI5[1][165] , \RI5[1][161] , \RI5[1][160] ,
         \RI5[1][159] , \RI5[1][158] , \RI5[1][157] , \RI5[1][156] ,
         \RI5[1][155] , \RI5[1][154] , \RI5[1][153] , \RI5[1][149] ,
         \RI5[1][148] , \RI5[1][147] , \RI5[1][144] , \RI5[1][143] ,
         \RI5[1][142] , \RI5[1][140] , \RI5[1][139] , \RI5[1][138] ,
         \RI5[1][137] , \RI5[1][136] , \RI5[1][135] , \RI5[1][134] ,
         \RI5[1][133] , \RI5[1][132] , \RI5[1][131] , \RI5[1][130] ,
         \RI5[1][129] , \RI5[1][128] , \RI5[1][127] , \RI5[1][126] ,
         \RI5[1][123] , \RI5[1][121] , \RI5[1][120] , \RI5[1][119] ,
         \RI5[1][118] , \RI5[1][116] , \RI5[1][115] , \RI5[1][114] ,
         \RI5[1][113] , \RI5[1][112] , \RI5[1][111] , \RI5[1][109] ,
         \RI5[1][107] , \RI5[1][106] , \RI5[1][105] , \RI5[1][104] ,
         \RI5[1][102] , \RI5[1][101] , \RI5[1][100] , \RI5[1][99] ,
         \RI5[1][98] , \RI5[1][97] , \RI5[1][96] , \RI5[1][95] , \RI5[1][93] ,
         \RI5[1][92] , \RI5[1][91] , \RI5[1][90] , \RI5[1][89] , \RI5[1][88] ,
         \RI5[1][87] , \RI5[1][86] , \RI5[1][85] , \RI5[1][82] , \RI5[1][81] ,
         \RI5[1][80] , \RI5[1][79] , \RI5[1][78] , \RI5[1][77] , \RI5[1][75] ,
         \RI5[1][70] , \RI5[1][69] , \RI5[1][68] , \RI5[1][67] , \RI5[1][66] ,
         \RI5[1][65] , \RI5[1][64] , \RI5[1][63] , \RI5[1][61] , \RI5[1][60] ,
         \RI5[1][59] , \RI5[1][57] , \RI5[1][56] , \RI5[1][55] , \RI5[1][54] ,
         \RI5[1][53] , \RI5[1][52] , \RI5[1][51] , \RI5[1][49] , \RI5[1][47] ,
         \RI5[1][46] , \RI5[1][43] , \RI5[1][42] , \RI5[1][41] , \RI5[1][40] ,
         \RI5[1][39] , \RI5[1][35] , \RI5[1][33] , \RI5[1][31] , \RI5[1][30] ,
         \RI5[1][29] , \RI5[1][28] , \RI5[1][27] , \RI5[1][26] , \RI5[1][25] ,
         \RI5[1][24] , \RI5[1][23] , \RI5[1][20] , \RI5[1][19] , \RI5[1][18] ,
         \RI5[1][17] , \RI5[1][16] , \RI5[1][14] , \RI5[1][13] , \RI5[1][12] ,
         \RI5[1][11] , \RI5[1][10] , \RI5[1][9] , \RI5[1][8] , \RI5[1][6] ,
         \RI5[1][5] , \RI5[1][2] , \RI5[2][191] , \RI5[2][190] , \RI5[2][189] ,
         \RI5[2][188] , \RI5[2][187] , \RI5[2][186] , \RI5[2][185] ,
         \RI5[2][184] , \RI5[2][182] , \RI5[2][180] , \RI5[2][178] ,
         \RI5[2][177] , \RI5[2][176] , \RI5[2][175] , \RI5[2][174] ,
         \RI5[2][173] , \RI5[2][170] , \RI5[2][169] , \RI5[2][168] ,
         \RI5[2][167] , \RI5[2][166] , \RI5[2][165] , \RI5[2][163] ,
         \RI5[2][161] , \RI5[2][160] , \RI5[2][159] , \RI5[2][158] ,
         \RI5[2][157] , \RI5[2][156] , \RI5[2][155] , \RI5[2][154] ,
         \RI5[2][153] , \RI5[2][152] , \RI5[2][149] , \RI5[2][148] ,
         \RI5[2][145] , \RI5[2][144] , \RI5[2][142] , \RI5[2][140] ,
         \RI5[2][139] , \RI5[2][138] , \RI5[2][137] , \RI5[2][136] ,
         \RI5[2][135] , \RI5[2][134] , \RI5[2][132] , \RI5[2][130] ,
         \RI5[2][129] , \RI5[2][128] , \RI5[2][127] , \RI5[2][126] ,
         \RI5[2][125] , \RI5[2][123] , \RI5[2][119] , \RI5[2][118] ,
         \RI5[2][117] , \RI5[2][116] , \RI5[2][114] , \RI5[2][113] ,
         \RI5[2][111] , \RI5[2][109] , \RI5[2][108] , \RI5[2][107] ,
         \RI5[2][105] , \RI5[2][104] , \RI5[2][103] , \RI5[2][102] ,
         \RI5[2][101] , \RI5[2][97] , \RI5[2][96] , \RI5[2][95] , \RI5[2][94] ,
         \RI5[2][93] , \RI5[2][91] , \RI5[2][90] , \RI5[2][88] , \RI5[2][87] ,
         \RI5[2][86] , \RI5[2][85] , \RI5[2][83] , \RI5[2][82] , \RI5[2][81] ,
         \RI5[2][80] , \RI5[2][78] , \RI5[2][77] , \RI5[2][76] , \RI5[2][75] ,
         \RI5[2][73] , \RI5[2][72] , \RI5[2][71] , \RI5[2][69] , \RI5[2][67] ,
         \RI5[2][66] , \RI5[2][64] , \RI5[2][62] , \RI5[2][59] , \RI5[2][58] ,
         \RI5[2][57] , \RI5[2][54] , \RI5[2][53] , \RI5[2][51] , \RI5[2][50] ,
         \RI5[2][48] , \RI5[2][47] , \RI5[2][46] , \RI5[2][44] , \RI5[2][43] ,
         \RI5[2][42] , \RI5[2][39] , \RI5[2][38] , \RI5[2][37] , \RI5[2][36] ,
         \RI5[2][34] , \RI5[2][33] , \RI5[2][32] , \RI5[2][31] , \RI5[2][30] ,
         \RI5[2][27] , \RI5[2][26] , \RI5[2][21] , \RI5[2][20] , \RI5[2][19] ,
         \RI5[2][18] , \RI5[2][17] , \RI5[2][16] , \RI5[2][15] , \RI5[2][13] ,
         \RI5[2][12] , \RI5[2][11] , \RI5[2][9] , \RI5[2][8] , \RI5[2][6] ,
         \RI5[2][5] , \RI5[2][4] , \RI5[2][2] , \RI5[2][1] , \RI5[2][0] ,
         \RI5[3][191] , \RI5[3][190] , \RI5[3][189] , \RI5[3][186] ,
         \RI5[3][185] , \RI5[3][181] , \RI5[3][180] , \RI5[3][179] ,
         \RI5[3][175] , \RI5[3][174] , \RI5[3][173] , \RI5[3][172] ,
         \RI5[3][171] , \RI5[3][169] , \RI5[3][168] , \RI5[3][167] ,
         \RI5[3][166] , \RI5[3][165] , \RI5[3][163] , \RI5[3][162] ,
         \RI5[3][161] , \RI5[3][160] , \RI5[3][154] , \RI5[3][153] ,
         \RI5[3][152] , \RI5[3][150] , \RI5[3][149] , \RI5[3][148] ,
         \RI5[3][146] , \RI5[3][145] , \RI5[3][139] , \RI5[3][138] ,
         \RI5[3][137] , \RI5[3][136] , \RI5[3][135] , \RI5[3][134] ,
         \RI5[3][132] , \RI5[3][131] , \RI5[3][130] , \RI5[3][127] ,
         \RI5[3][126] , \RI5[3][125] , \RI5[3][124] , \RI5[3][123] ,
         \RI5[3][122] , \RI5[3][121] , \RI5[3][120] , \RI5[3][119] ,
         \RI5[3][117] , \RI5[3][114] , \RI5[3][113] , \RI5[3][112] ,
         \RI5[3][111] , \RI5[3][110] , \RI5[3][108] , \RI5[3][107] ,
         \RI5[3][106] , \RI5[3][104] , \RI5[3][103] , \RI5[3][101] ,
         \RI5[3][100] , \RI5[3][98] , \RI5[3][97] , \RI5[3][95] , \RI5[3][93] ,
         \RI5[3][92] , \RI5[3][91] , \RI5[3][90] , \RI5[3][89] , \RI5[3][88] ,
         \RI5[3][87] , \RI5[3][86] , \RI5[3][85] , \RI5[3][84] , \RI5[3][83] ,
         \RI5[3][82] , \RI5[3][81] , \RI5[3][79] , \RI5[3][78] , \RI5[3][77] ,
         \RI5[3][76] , \RI5[3][75] , \RI5[3][74] , \RI5[3][73] , \RI5[3][72] ,
         \RI5[3][70] , \RI5[3][68] , \RI5[3][67] , \RI5[3][66] , \RI5[3][65] ,
         \RI5[3][64] , \RI5[3][63] , \RI5[3][61] , \RI5[3][60] , \RI5[3][59] ,
         \RI5[3][58] , \RI5[3][57] , \RI5[3][56] , \RI5[3][55] , \RI5[3][54] ,
         \RI5[3][52] , \RI5[3][51] , \RI5[3][50] , \RI5[3][48] , \RI5[3][47] ,
         \RI5[3][45] , \RI5[3][44] , \RI5[3][42] , \RI5[3][41] , \RI5[3][40] ,
         \RI5[3][38] , \RI5[3][36] , \RI5[3][35] , \RI5[3][34] , \RI5[3][33] ,
         \RI5[3][31] , \RI5[3][30] , \RI5[3][28] , \RI5[3][27] , \RI5[3][26] ,
         \RI5[3][25] , \RI5[3][23] , \RI5[3][22] , \RI5[3][18] , \RI5[3][17] ,
         \RI5[3][16] , \RI5[3][14] , \RI5[3][13] , \RI5[3][12] , \RI5[3][11] ,
         \RI5[3][10] , \RI5[3][9] , \RI5[3][8] , \RI5[3][6] , \RI5[3][4] ,
         \RI5[3][3] , \RI5[3][2] , \RI5[4][191] , \RI5[4][190] , \RI5[4][189] ,
         \RI5[4][187] , \RI5[4][186] , \RI5[4][185] , \RI5[4][182] ,
         \RI5[4][181] , \RI5[4][180] , \RI5[4][179] , \RI5[4][178] ,
         \RI5[4][175] , \RI5[4][174] , \RI5[4][172] , \RI5[4][166] ,
         \RI5[4][164] , \RI5[4][163] , \RI5[4][162] , \RI5[4][161] ,
         \RI5[4][159] , \RI5[4][158] , \RI5[4][157] , \RI5[4][156] ,
         \RI5[4][155] , \RI5[4][153] , \RI5[4][152] , \RI5[4][151] ,
         \RI5[4][150] , \RI5[4][149] , \RI5[4][147] , \RI5[4][146] ,
         \RI5[4][145] , \RI5[4][144] , \RI5[4][143] , \RI5[4][142] ,
         \RI5[4][140] , \RI5[4][139] , \RI5[4][138] , \RI5[4][137] ,
         \RI5[4][136] , \RI5[4][134] , \RI5[4][133] , \RI5[4][131] ,
         \RI5[4][130] , \RI5[4][128] , \RI5[4][127] , \RI5[4][126] ,
         \RI5[4][125] , \RI5[4][124] , \RI5[4][123] , \RI5[4][122] ,
         \RI5[4][121] , \RI5[4][119] , \RI5[4][116] , \RI5[4][115] ,
         \RI5[4][114] , \RI5[4][113] , \RI5[4][112] , \RI5[4][111] ,
         \RI5[4][110] , \RI5[4][109] , \RI5[4][107] , \RI5[4][106] ,
         \RI5[4][105] , \RI5[4][104] , \RI5[4][103] , \RI5[4][102] ,
         \RI5[4][101] , \RI5[4][100] , \RI5[4][99] , \RI5[4][98] ,
         \RI5[4][96] , \RI5[4][95] , \RI5[4][92] , \RI5[4][91] , \RI5[4][90] ,
         \RI5[4][89] , \RI5[4][88] , \RI5[4][85] , \RI5[4][84] , \RI5[4][83] ,
         \RI5[4][82] , \RI5[4][81] , \RI5[4][80] , \RI5[4][79] , \RI5[4][78] ,
         \RI5[4][74] , \RI5[4][72] , \RI5[4][71] , \RI5[4][70] , \RI5[4][69] ,
         \RI5[4][68] , \RI5[4][67] , \RI5[4][66] , \RI5[4][65] , \RI5[4][62] ,
         \RI5[4][61] , \RI5[4][60] , \RI5[4][59] , \RI5[4][58] , \RI5[4][57] ,
         \RI5[4][56] , \RI5[4][52] , \RI5[4][51] , \RI5[4][50] , \RI5[4][49] ,
         \RI5[4][48] , \RI5[4][47] , \RI5[4][46] , \RI5[4][44] , \RI5[4][42] ,
         \RI5[4][41] , \RI5[4][40] , \RI5[4][38] , \RI5[4][37] , \RI5[4][36] ,
         \RI5[4][35] , \RI5[4][34] , \RI5[4][33] , \RI5[4][32] , \RI5[4][31] ,
         \RI5[4][30] , \RI5[4][29] , \RI5[4][28] , \RI5[4][26] , \RI5[4][25] ,
         \RI5[4][24] , \RI5[4][21] , \RI5[4][20] , \RI5[4][19] , \RI5[4][17] ,
         \RI5[4][16] , \RI5[4][14] , \RI5[4][13] , \RI5[4][11] , \RI5[4][10] ,
         \RI5[4][8] , \RI5[4][7] , \RI5[4][6] , \RI5[4][5] , \RI5[4][4] ,
         \RI5[4][1] , \RI5[4][0] , \MC_ARK_ARC_1_0/buf_output[191] ,
         \MC_ARK_ARC_1_0/buf_output[190] , \MC_ARK_ARC_1_0/buf_output[189] ,
         \MC_ARK_ARC_1_0/buf_output[188] , \MC_ARK_ARC_1_0/buf_output[187] ,
         \MC_ARK_ARC_1_0/buf_output[186] , \MC_ARK_ARC_1_0/buf_output[185] ,
         \MC_ARK_ARC_1_0/buf_output[184] , \MC_ARK_ARC_1_0/buf_output[183] ,
         \MC_ARK_ARC_1_0/buf_output[182] , \MC_ARK_ARC_1_0/buf_output[181] ,
         \MC_ARK_ARC_1_0/buf_output[180] , \MC_ARK_ARC_1_0/buf_output[178] ,
         \MC_ARK_ARC_1_0/buf_output[177] , \MC_ARK_ARC_1_0/buf_output[176] ,
         \MC_ARK_ARC_1_0/buf_output[175] , \MC_ARK_ARC_1_0/buf_output[174] ,
         \MC_ARK_ARC_1_0/buf_output[173] , \MC_ARK_ARC_1_0/buf_output[172] ,
         \MC_ARK_ARC_1_0/buf_output[171] , \MC_ARK_ARC_1_0/buf_output[170] ,
         \MC_ARK_ARC_1_0/buf_output[169] , \MC_ARK_ARC_1_0/buf_output[168] ,
         \MC_ARK_ARC_1_0/buf_output[167] , \MC_ARK_ARC_1_0/buf_output[166] ,
         \MC_ARK_ARC_1_0/buf_output[165] , \MC_ARK_ARC_1_0/buf_output[164] ,
         \MC_ARK_ARC_1_0/buf_output[163] , \MC_ARK_ARC_1_0/buf_output[162] ,
         \MC_ARK_ARC_1_0/buf_output[161] , \MC_ARK_ARC_1_0/buf_output[160] ,
         \MC_ARK_ARC_1_0/buf_output[159] , \MC_ARK_ARC_1_0/buf_output[158] ,
         \MC_ARK_ARC_1_0/buf_output[157] , \MC_ARK_ARC_1_0/buf_output[156] ,
         \MC_ARK_ARC_1_0/buf_output[155] , \MC_ARK_ARC_1_0/buf_output[154] ,
         \MC_ARK_ARC_1_0/buf_output[153] , \MC_ARK_ARC_1_0/buf_output[152] ,
         \MC_ARK_ARC_1_0/buf_output[151] , \MC_ARK_ARC_1_0/buf_output[150] ,
         \MC_ARK_ARC_1_0/buf_output[148] , \MC_ARK_ARC_1_0/buf_output[147] ,
         \MC_ARK_ARC_1_0/buf_output[146] , \MC_ARK_ARC_1_0/buf_output[145] ,
         \MC_ARK_ARC_1_0/buf_output[144] , \MC_ARK_ARC_1_0/buf_output[143] ,
         \MC_ARK_ARC_1_0/buf_output[142] , \MC_ARK_ARC_1_0/buf_output[141] ,
         \MC_ARK_ARC_1_0/buf_output[140] , \MC_ARK_ARC_1_0/buf_output[139] ,
         \MC_ARK_ARC_1_0/buf_output[138] , \MC_ARK_ARC_1_0/buf_output[137] ,
         \MC_ARK_ARC_1_0/buf_output[136] , \MC_ARK_ARC_1_0/buf_output[135] ,
         \MC_ARK_ARC_1_0/buf_output[134] , \MC_ARK_ARC_1_0/buf_output[133] ,
         \MC_ARK_ARC_1_0/buf_output[132] , \MC_ARK_ARC_1_0/buf_output[131] ,
         \MC_ARK_ARC_1_0/buf_output[130] , \MC_ARK_ARC_1_0/buf_output[129] ,
         \MC_ARK_ARC_1_0/buf_output[128] , \MC_ARK_ARC_1_0/buf_output[127] ,
         \MC_ARK_ARC_1_0/buf_output[126] , \MC_ARK_ARC_1_0/buf_output[125] ,
         \MC_ARK_ARC_1_0/buf_output[124] , \MC_ARK_ARC_1_0/buf_output[123] ,
         \MC_ARK_ARC_1_0/buf_output[122] , \MC_ARK_ARC_1_0/buf_output[121] ,
         \MC_ARK_ARC_1_0/buf_output[120] , \MC_ARK_ARC_1_0/buf_output[119] ,
         \MC_ARK_ARC_1_0/buf_output[118] , \MC_ARK_ARC_1_0/buf_output[117] ,
         \MC_ARK_ARC_1_0/buf_output[116] , \MC_ARK_ARC_1_0/buf_output[115] ,
         \MC_ARK_ARC_1_0/buf_output[114] , \MC_ARK_ARC_1_0/buf_output[113] ,
         \MC_ARK_ARC_1_0/buf_output[112] , \MC_ARK_ARC_1_0/buf_output[111] ,
         \MC_ARK_ARC_1_0/buf_output[110] , \MC_ARK_ARC_1_0/buf_output[109] ,
         \MC_ARK_ARC_1_0/buf_output[108] , \MC_ARK_ARC_1_0/buf_output[107] ,
         \MC_ARK_ARC_1_0/buf_output[106] , \MC_ARK_ARC_1_0/buf_output[105] ,
         \MC_ARK_ARC_1_0/buf_output[104] , \MC_ARK_ARC_1_0/buf_output[103] ,
         \MC_ARK_ARC_1_0/buf_output[102] , \MC_ARK_ARC_1_0/buf_output[101] ,
         \MC_ARK_ARC_1_0/buf_output[100] , \MC_ARK_ARC_1_0/buf_output[99] ,
         \MC_ARK_ARC_1_0/buf_output[98] , \MC_ARK_ARC_1_0/buf_output[97] ,
         \MC_ARK_ARC_1_0/buf_output[96] , \MC_ARK_ARC_1_0/buf_output[95] ,
         \MC_ARK_ARC_1_0/buf_output[94] , \MC_ARK_ARC_1_0/buf_output[93] ,
         \MC_ARK_ARC_1_0/buf_output[92] , \MC_ARK_ARC_1_0/buf_output[91] ,
         \MC_ARK_ARC_1_0/buf_output[90] , \MC_ARK_ARC_1_0/buf_output[89] ,
         \MC_ARK_ARC_1_0/buf_output[88] , \MC_ARK_ARC_1_0/buf_output[87] ,
         \MC_ARK_ARC_1_0/buf_output[86] , \MC_ARK_ARC_1_0/buf_output[85] ,
         \MC_ARK_ARC_1_0/buf_output[84] , \MC_ARK_ARC_1_0/buf_output[83] ,
         \MC_ARK_ARC_1_0/buf_output[82] , \MC_ARK_ARC_1_0/buf_output[81] ,
         \MC_ARK_ARC_1_0/buf_output[80] , \MC_ARK_ARC_1_0/buf_output[79] ,
         \MC_ARK_ARC_1_0/buf_output[78] , \MC_ARK_ARC_1_0/buf_output[77] ,
         \MC_ARK_ARC_1_0/buf_output[76] , \MC_ARK_ARC_1_0/buf_output[75] ,
         \MC_ARK_ARC_1_0/buf_output[74] , \MC_ARK_ARC_1_0/buf_output[73] ,
         \MC_ARK_ARC_1_0/buf_output[72] , \MC_ARK_ARC_1_0/buf_output[71] ,
         \MC_ARK_ARC_1_0/buf_output[70] , \MC_ARK_ARC_1_0/buf_output[69] ,
         \MC_ARK_ARC_1_0/buf_output[68] , \MC_ARK_ARC_1_0/buf_output[67] ,
         \MC_ARK_ARC_1_0/buf_output[66] , \MC_ARK_ARC_1_0/buf_output[65] ,
         \MC_ARK_ARC_1_0/buf_output[64] , \MC_ARK_ARC_1_0/buf_output[63] ,
         \MC_ARK_ARC_1_0/buf_output[62] , \MC_ARK_ARC_1_0/buf_output[61] ,
         \MC_ARK_ARC_1_0/buf_output[60] , \MC_ARK_ARC_1_0/buf_output[59] ,
         \MC_ARK_ARC_1_0/buf_output[58] , \MC_ARK_ARC_1_0/buf_output[57] ,
         \MC_ARK_ARC_1_0/buf_output[56] , \MC_ARK_ARC_1_0/buf_output[55] ,
         \MC_ARK_ARC_1_0/buf_output[54] , \MC_ARK_ARC_1_0/buf_output[53] ,
         \MC_ARK_ARC_1_0/buf_output[52] , \MC_ARK_ARC_1_0/buf_output[51] ,
         \MC_ARK_ARC_1_0/buf_output[50] , \MC_ARK_ARC_1_0/buf_output[49] ,
         \MC_ARK_ARC_1_0/buf_output[48] , \MC_ARK_ARC_1_0/buf_output[47] ,
         \MC_ARK_ARC_1_0/buf_output[46] , \MC_ARK_ARC_1_0/buf_output[45] ,
         \MC_ARK_ARC_1_0/buf_output[44] , \MC_ARK_ARC_1_0/buf_output[43] ,
         \MC_ARK_ARC_1_0/buf_output[42] , \MC_ARK_ARC_1_0/buf_output[41] ,
         \MC_ARK_ARC_1_0/buf_output[40] , \MC_ARK_ARC_1_0/buf_output[39] ,
         \MC_ARK_ARC_1_0/buf_output[38] , \MC_ARK_ARC_1_0/buf_output[37] ,
         \MC_ARK_ARC_1_0/buf_output[36] , \MC_ARK_ARC_1_0/buf_output[35] ,
         \MC_ARK_ARC_1_0/buf_output[34] , \MC_ARK_ARC_1_0/buf_output[33] ,
         \MC_ARK_ARC_1_0/buf_output[32] , \MC_ARK_ARC_1_0/buf_output[31] ,
         \MC_ARK_ARC_1_0/buf_output[30] , \MC_ARK_ARC_1_0/buf_output[29] ,
         \MC_ARK_ARC_1_0/buf_output[28] , \MC_ARK_ARC_1_0/buf_output[27] ,
         \MC_ARK_ARC_1_0/buf_output[26] , \MC_ARK_ARC_1_0/buf_output[25] ,
         \MC_ARK_ARC_1_0/buf_output[24] , \MC_ARK_ARC_1_0/buf_output[22] ,
         \MC_ARK_ARC_1_0/buf_output[21] , \MC_ARK_ARC_1_0/buf_output[20] ,
         \MC_ARK_ARC_1_0/buf_output[19] , \MC_ARK_ARC_1_0/buf_output[18] ,
         \MC_ARK_ARC_1_0/buf_output[17] , \MC_ARK_ARC_1_0/buf_output[16] ,
         \MC_ARK_ARC_1_0/buf_output[15] , \MC_ARK_ARC_1_0/buf_output[14] ,
         \MC_ARK_ARC_1_0/buf_output[13] , \MC_ARK_ARC_1_0/buf_output[12] ,
         \MC_ARK_ARC_1_0/buf_output[10] , \MC_ARK_ARC_1_0/buf_output[9] ,
         \MC_ARK_ARC_1_0/buf_output[8] , \MC_ARK_ARC_1_0/buf_output[7] ,
         \MC_ARK_ARC_1_0/buf_output[6] , \MC_ARK_ARC_1_0/buf_output[5] ,
         \MC_ARK_ARC_1_0/buf_output[4] , \MC_ARK_ARC_1_0/buf_output[3] ,
         \MC_ARK_ARC_1_0/buf_output[2] , \MC_ARK_ARC_1_0/buf_output[1] ,
         \MC_ARK_ARC_1_0/buf_output[0] , \MC_ARK_ARC_1_0/temp6[190] ,
         \MC_ARK_ARC_1_0/temp6[189] , \MC_ARK_ARC_1_0/temp6[187] ,
         \MC_ARK_ARC_1_0/temp6[186] , \MC_ARK_ARC_1_0/temp6[185] ,
         \MC_ARK_ARC_1_0/temp6[184] , \MC_ARK_ARC_1_0/temp6[183] ,
         \MC_ARK_ARC_1_0/temp6[182] , \MC_ARK_ARC_1_0/temp6[180] ,
         \MC_ARK_ARC_1_0/temp6[178] , \MC_ARK_ARC_1_0/temp6[177] ,
         \MC_ARK_ARC_1_0/temp6[175] , \MC_ARK_ARC_1_0/temp6[174] ,
         \MC_ARK_ARC_1_0/temp6[171] , \MC_ARK_ARC_1_0/temp6[169] ,
         \MC_ARK_ARC_1_0/temp6[163] , \MC_ARK_ARC_1_0/temp6[162] ,
         \MC_ARK_ARC_1_0/temp6[161] , \MC_ARK_ARC_1_0/temp6[160] ,
         \MC_ARK_ARC_1_0/temp6[157] , \MC_ARK_ARC_1_0/temp6[155] ,
         \MC_ARK_ARC_1_0/temp6[154] , \MC_ARK_ARC_1_0/temp6[151] ,
         \MC_ARK_ARC_1_0/temp6[150] , \MC_ARK_ARC_1_0/temp6[147] ,
         \MC_ARK_ARC_1_0/temp6[145] , \MC_ARK_ARC_1_0/temp6[144] ,
         \MC_ARK_ARC_1_0/temp6[143] , \MC_ARK_ARC_1_0/temp6[142] ,
         \MC_ARK_ARC_1_0/temp6[139] , \MC_ARK_ARC_1_0/temp6[137] ,
         \MC_ARK_ARC_1_0/temp6[135] , \MC_ARK_ARC_1_0/temp6[133] ,
         \MC_ARK_ARC_1_0/temp6[130] , \MC_ARK_ARC_1_0/temp6[129] ,
         \MC_ARK_ARC_1_0/temp6[127] , \MC_ARK_ARC_1_0/temp6[126] ,
         \MC_ARK_ARC_1_0/temp6[124] , \MC_ARK_ARC_1_0/temp6[121] ,
         \MC_ARK_ARC_1_0/temp6[120] , \MC_ARK_ARC_1_0/temp6[119] ,
         \MC_ARK_ARC_1_0/temp6[118] , \MC_ARK_ARC_1_0/temp6[115] ,
         \MC_ARK_ARC_1_0/temp6[114] , \MC_ARK_ARC_1_0/temp6[113] ,
         \MC_ARK_ARC_1_0/temp6[111] , \MC_ARK_ARC_1_0/temp6[108] ,
         \MC_ARK_ARC_1_0/temp6[106] , \MC_ARK_ARC_1_0/temp6[101] ,
         \MC_ARK_ARC_1_0/temp6[100] , \MC_ARK_ARC_1_0/temp6[98] ,
         \MC_ARK_ARC_1_0/temp6[97] , \MC_ARK_ARC_1_0/temp6[95] ,
         \MC_ARK_ARC_1_0/temp6[91] , \MC_ARK_ARC_1_0/temp6[87] ,
         \MC_ARK_ARC_1_0/temp6[85] , \MC_ARK_ARC_1_0/temp6[84] ,
         \MC_ARK_ARC_1_0/temp6[83] , \MC_ARK_ARC_1_0/temp6[82] ,
         \MC_ARK_ARC_1_0/temp6[78] , \MC_ARK_ARC_1_0/temp6[77] ,
         \MC_ARK_ARC_1_0/temp6[76] , \MC_ARK_ARC_1_0/temp6[72] ,
         \MC_ARK_ARC_1_0/temp6[70] , \MC_ARK_ARC_1_0/temp6[67] ,
         \MC_ARK_ARC_1_0/temp6[63] , \MC_ARK_ARC_1_0/temp6[62] ,
         \MC_ARK_ARC_1_0/temp6[61] , \MC_ARK_ARC_1_0/temp6[60] ,
         \MC_ARK_ARC_1_0/temp6[58] , \MC_ARK_ARC_1_0/temp6[56] ,
         \MC_ARK_ARC_1_0/temp6[54] , \MC_ARK_ARC_1_0/temp6[52] ,
         \MC_ARK_ARC_1_0/temp6[51] , \MC_ARK_ARC_1_0/temp6[49] ,
         \MC_ARK_ARC_1_0/temp6[48] , \MC_ARK_ARC_1_0/temp6[47] ,
         \MC_ARK_ARC_1_0/temp6[46] , \MC_ARK_ARC_1_0/temp6[45] ,
         \MC_ARK_ARC_1_0/temp6[43] , \MC_ARK_ARC_1_0/temp6[40] ,
         \MC_ARK_ARC_1_0/temp6[39] , \MC_ARK_ARC_1_0/temp6[37] ,
         \MC_ARK_ARC_1_0/temp6[36] , \MC_ARK_ARC_1_0/temp6[35] ,
         \MC_ARK_ARC_1_0/temp6[33] , \MC_ARK_ARC_1_0/temp6[32] ,
         \MC_ARK_ARC_1_0/temp6[26] , \MC_ARK_ARC_1_0/temp6[25] ,
         \MC_ARK_ARC_1_0/temp6[24] , \MC_ARK_ARC_1_0/temp6[21] ,
         \MC_ARK_ARC_1_0/temp6[19] , \MC_ARK_ARC_1_0/temp6[16] ,
         \MC_ARK_ARC_1_0/temp6[13] , \MC_ARK_ARC_1_0/temp6[12] ,
         \MC_ARK_ARC_1_0/temp6[8] , \MC_ARK_ARC_1_0/temp6[7] ,
         \MC_ARK_ARC_1_0/temp6[6] , \MC_ARK_ARC_1_0/temp6[5] ,
         \MC_ARK_ARC_1_0/temp6[3] , \MC_ARK_ARC_1_0/temp6[2] ,
         \MC_ARK_ARC_1_0/temp6[0] , \MC_ARK_ARC_1_0/temp5[190] ,
         \MC_ARK_ARC_1_0/temp5[187] , \MC_ARK_ARC_1_0/temp5[185] ,
         \MC_ARK_ARC_1_0/temp5[184] , \MC_ARK_ARC_1_0/temp5[182] ,
         \MC_ARK_ARC_1_0/temp5[181] , \MC_ARK_ARC_1_0/temp5[180] ,
         \MC_ARK_ARC_1_0/temp5[179] , \MC_ARK_ARC_1_0/temp5[178] ,
         \MC_ARK_ARC_1_0/temp5[176] , \MC_ARK_ARC_1_0/temp5[175] ,
         \MC_ARK_ARC_1_0/temp5[174] , \MC_ARK_ARC_1_0/temp5[169] ,
         \MC_ARK_ARC_1_0/temp5[168] , \MC_ARK_ARC_1_0/temp5[167] ,
         \MC_ARK_ARC_1_0/temp5[166] , \MC_ARK_ARC_1_0/temp5[162] ,
         \MC_ARK_ARC_1_0/temp5[161] , \MC_ARK_ARC_1_0/temp5[158] ,
         \MC_ARK_ARC_1_0/temp5[157] , \MC_ARK_ARC_1_0/temp5[156] ,
         \MC_ARK_ARC_1_0/temp5[154] , \MC_ARK_ARC_1_0/temp5[153] ,
         \MC_ARK_ARC_1_0/temp5[151] , \MC_ARK_ARC_1_0/temp5[150] ,
         \MC_ARK_ARC_1_0/temp5[149] , \MC_ARK_ARC_1_0/temp5[148] ,
         \MC_ARK_ARC_1_0/temp5[146] , \MC_ARK_ARC_1_0/temp5[145] ,
         \MC_ARK_ARC_1_0/temp5[144] , \MC_ARK_ARC_1_0/temp5[142] ,
         \MC_ARK_ARC_1_0/temp5[140] , \MC_ARK_ARC_1_0/temp5[133] ,
         \MC_ARK_ARC_1_0/temp5[130] , \MC_ARK_ARC_1_0/temp5[129] ,
         \MC_ARK_ARC_1_0/temp5[128] , \MC_ARK_ARC_1_0/temp5[124] ,
         \MC_ARK_ARC_1_0/temp5[122] , \MC_ARK_ARC_1_0/temp5[121] ,
         \MC_ARK_ARC_1_0/temp5[120] , \MC_ARK_ARC_1_0/temp5[119] ,
         \MC_ARK_ARC_1_0/temp5[118] , \MC_ARK_ARC_1_0/temp5[116] ,
         \MC_ARK_ARC_1_0/temp5[115] , \MC_ARK_ARC_1_0/temp5[114] ,
         \MC_ARK_ARC_1_0/temp5[112] , \MC_ARK_ARC_1_0/temp5[111] ,
         \MC_ARK_ARC_1_0/temp5[106] , \MC_ARK_ARC_1_0/temp5[105] ,
         \MC_ARK_ARC_1_0/temp5[104] , \MC_ARK_ARC_1_0/temp5[103] ,
         \MC_ARK_ARC_1_0/temp5[101] , \MC_ARK_ARC_1_0/temp5[97] ,
         \MC_ARK_ARC_1_0/temp5[96] , \MC_ARK_ARC_1_0/temp5[93] ,
         \MC_ARK_ARC_1_0/temp5[91] , \MC_ARK_ARC_1_0/temp5[88] ,
         \MC_ARK_ARC_1_0/temp5[85] , \MC_ARK_ARC_1_0/temp5[84] ,
         \MC_ARK_ARC_1_0/temp5[83] , \MC_ARK_ARC_1_0/temp5[77] ,
         \MC_ARK_ARC_1_0/temp5[76] , \MC_ARK_ARC_1_0/temp5[74] ,
         \MC_ARK_ARC_1_0/temp5[73] , \MC_ARK_ARC_1_0/temp5[72] ,
         \MC_ARK_ARC_1_0/temp5[71] , \MC_ARK_ARC_1_0/temp5[70] ,
         \MC_ARK_ARC_1_0/temp5[69] , \MC_ARK_ARC_1_0/temp5[65] ,
         \MC_ARK_ARC_1_0/temp5[64] , \MC_ARK_ARC_1_0/temp5[62] ,
         \MC_ARK_ARC_1_0/temp5[61] , \MC_ARK_ARC_1_0/temp5[59] ,
         \MC_ARK_ARC_1_0/temp5[58] , \MC_ARK_ARC_1_0/temp5[55] ,
         \MC_ARK_ARC_1_0/temp5[54] , \MC_ARK_ARC_1_0/temp5[53] ,
         \MC_ARK_ARC_1_0/temp5[48] , \MC_ARK_ARC_1_0/temp5[46] ,
         \MC_ARK_ARC_1_0/temp5[45] , \MC_ARK_ARC_1_0/temp5[43] ,
         \MC_ARK_ARC_1_0/temp5[40] , \MC_ARK_ARC_1_0/temp5[39] ,
         \MC_ARK_ARC_1_0/temp5[37] , \MC_ARK_ARC_1_0/temp5[33] ,
         \MC_ARK_ARC_1_0/temp5[30] , \MC_ARK_ARC_1_0/temp5[25] ,
         \MC_ARK_ARC_1_0/temp5[23] , \MC_ARK_ARC_1_0/temp5[19] ,
         \MC_ARK_ARC_1_0/temp5[18] , \MC_ARK_ARC_1_0/temp5[16] ,
         \MC_ARK_ARC_1_0/temp5[15] , \MC_ARK_ARC_1_0/temp5[13] ,
         \MC_ARK_ARC_1_0/temp5[12] , \MC_ARK_ARC_1_0/temp5[8] ,
         \MC_ARK_ARC_1_0/temp5[7] , \MC_ARK_ARC_1_0/temp5[2] ,
         \MC_ARK_ARC_1_0/temp5[0] , \MC_ARK_ARC_1_0/temp4[191] ,
         \MC_ARK_ARC_1_0/temp4[190] , \MC_ARK_ARC_1_0/temp4[189] ,
         \MC_ARK_ARC_1_0/temp4[188] , \MC_ARK_ARC_1_0/temp4[187] ,
         \MC_ARK_ARC_1_0/temp4[186] , \MC_ARK_ARC_1_0/temp4[185] ,
         \MC_ARK_ARC_1_0/temp4[184] , \MC_ARK_ARC_1_0/temp4[183] ,
         \MC_ARK_ARC_1_0/temp4[182] , \MC_ARK_ARC_1_0/temp4[181] ,
         \MC_ARK_ARC_1_0/temp4[180] , \MC_ARK_ARC_1_0/temp4[179] ,
         \MC_ARK_ARC_1_0/temp4[178] , \MC_ARK_ARC_1_0/temp4[177] ,
         \MC_ARK_ARC_1_0/temp4[175] , \MC_ARK_ARC_1_0/temp4[174] ,
         \MC_ARK_ARC_1_0/temp4[173] , \MC_ARK_ARC_1_0/temp4[172] ,
         \MC_ARK_ARC_1_0/temp4[171] , \MC_ARK_ARC_1_0/temp4[170] ,
         \MC_ARK_ARC_1_0/temp4[169] , \MC_ARK_ARC_1_0/temp4[168] ,
         \MC_ARK_ARC_1_0/temp4[167] , \MC_ARK_ARC_1_0/temp4[165] ,
         \MC_ARK_ARC_1_0/temp4[163] , \MC_ARK_ARC_1_0/temp4[162] ,
         \MC_ARK_ARC_1_0/temp4[161] , \MC_ARK_ARC_1_0/temp4[160] ,
         \MC_ARK_ARC_1_0/temp4[159] , \MC_ARK_ARC_1_0/temp4[158] ,
         \MC_ARK_ARC_1_0/temp4[157] , \MC_ARK_ARC_1_0/temp4[156] ,
         \MC_ARK_ARC_1_0/temp4[154] , \MC_ARK_ARC_1_0/temp4[153] ,
         \MC_ARK_ARC_1_0/temp4[152] , \MC_ARK_ARC_1_0/temp4[151] ,
         \MC_ARK_ARC_1_0/temp4[150] , \MC_ARK_ARC_1_0/temp4[148] ,
         \MC_ARK_ARC_1_0/temp4[147] , \MC_ARK_ARC_1_0/temp4[146] ,
         \MC_ARK_ARC_1_0/temp4[145] , \MC_ARK_ARC_1_0/temp4[144] ,
         \MC_ARK_ARC_1_0/temp4[143] , \MC_ARK_ARC_1_0/temp4[142] ,
         \MC_ARK_ARC_1_0/temp4[141] , \MC_ARK_ARC_1_0/temp4[140] ,
         \MC_ARK_ARC_1_0/temp4[139] , \MC_ARK_ARC_1_0/temp4[138] ,
         \MC_ARK_ARC_1_0/temp4[137] , \MC_ARK_ARC_1_0/temp4[136] ,
         \MC_ARK_ARC_1_0/temp4[135] , \MC_ARK_ARC_1_0/temp4[133] ,
         \MC_ARK_ARC_1_0/temp4[132] , \MC_ARK_ARC_1_0/temp4[131] ,
         \MC_ARK_ARC_1_0/temp4[130] , \MC_ARK_ARC_1_0/temp4[129] ,
         \MC_ARK_ARC_1_0/temp4[128] , \MC_ARK_ARC_1_0/temp4[127] ,
         \MC_ARK_ARC_1_0/temp4[126] , \MC_ARK_ARC_1_0/temp4[125] ,
         \MC_ARK_ARC_1_0/temp4[124] , \MC_ARK_ARC_1_0/temp4[123] ,
         \MC_ARK_ARC_1_0/temp4[122] , \MC_ARK_ARC_1_0/temp4[121] ,
         \MC_ARK_ARC_1_0/temp4[120] , \MC_ARK_ARC_1_0/temp4[119] ,
         \MC_ARK_ARC_1_0/temp4[118] , \MC_ARK_ARC_1_0/temp4[117] ,
         \MC_ARK_ARC_1_0/temp4[116] , \MC_ARK_ARC_1_0/temp4[115] ,
         \MC_ARK_ARC_1_0/temp4[114] , \MC_ARK_ARC_1_0/temp4[113] ,
         \MC_ARK_ARC_1_0/temp4[112] , \MC_ARK_ARC_1_0/temp4[111] ,
         \MC_ARK_ARC_1_0/temp4[110] , \MC_ARK_ARC_1_0/temp4[109] ,
         \MC_ARK_ARC_1_0/temp4[108] , \MC_ARK_ARC_1_0/temp4[107] ,
         \MC_ARK_ARC_1_0/temp4[106] , \MC_ARK_ARC_1_0/temp4[105] ,
         \MC_ARK_ARC_1_0/temp4[104] , \MC_ARK_ARC_1_0/temp4[103] ,
         \MC_ARK_ARC_1_0/temp4[102] , \MC_ARK_ARC_1_0/temp4[101] ,
         \MC_ARK_ARC_1_0/temp4[100] , \MC_ARK_ARC_1_0/temp4[99] ,
         \MC_ARK_ARC_1_0/temp4[98] , \MC_ARK_ARC_1_0/temp4[97] ,
         \MC_ARK_ARC_1_0/temp4[96] , \MC_ARK_ARC_1_0/temp4[95] ,
         \MC_ARK_ARC_1_0/temp4[94] , \MC_ARK_ARC_1_0/temp4[93] ,
         \MC_ARK_ARC_1_0/temp4[92] , \MC_ARK_ARC_1_0/temp4[91] ,
         \MC_ARK_ARC_1_0/temp4[90] , \MC_ARK_ARC_1_0/temp4[88] ,
         \MC_ARK_ARC_1_0/temp4[86] , \MC_ARK_ARC_1_0/temp4[85] ,
         \MC_ARK_ARC_1_0/temp4[84] , \MC_ARK_ARC_1_0/temp4[83] ,
         \MC_ARK_ARC_1_0/temp4[82] , \MC_ARK_ARC_1_0/temp4[81] ,
         \MC_ARK_ARC_1_0/temp4[80] , \MC_ARK_ARC_1_0/temp4[79] ,
         \MC_ARK_ARC_1_0/temp4[78] , \MC_ARK_ARC_1_0/temp4[77] ,
         \MC_ARK_ARC_1_0/temp4[76] , \MC_ARK_ARC_1_0/temp4[75] ,
         \MC_ARK_ARC_1_0/temp4[74] , \MC_ARK_ARC_1_0/temp4[73] ,
         \MC_ARK_ARC_1_0/temp4[72] , \MC_ARK_ARC_1_0/temp4[71] ,
         \MC_ARK_ARC_1_0/temp4[70] , \MC_ARK_ARC_1_0/temp4[69] ,
         \MC_ARK_ARC_1_0/temp4[68] , \MC_ARK_ARC_1_0/temp4[67] ,
         \MC_ARK_ARC_1_0/temp4[66] , \MC_ARK_ARC_1_0/temp4[64] ,
         \MC_ARK_ARC_1_0/temp4[63] , \MC_ARK_ARC_1_0/temp4[62] ,
         \MC_ARK_ARC_1_0/temp4[61] , \MC_ARK_ARC_1_0/temp4[60] ,
         \MC_ARK_ARC_1_0/temp4[58] , \MC_ARK_ARC_1_0/temp4[57] ,
         \MC_ARK_ARC_1_0/temp4[55] , \MC_ARK_ARC_1_0/temp4[54] ,
         \MC_ARK_ARC_1_0/temp4[53] , \MC_ARK_ARC_1_0/temp4[52] ,
         \MC_ARK_ARC_1_0/temp4[51] , \MC_ARK_ARC_1_0/temp4[50] ,
         \MC_ARK_ARC_1_0/temp4[49] , \MC_ARK_ARC_1_0/temp4[48] ,
         \MC_ARK_ARC_1_0/temp4[46] , \MC_ARK_ARC_1_0/temp4[45] ,
         \MC_ARK_ARC_1_0/temp4[44] , \MC_ARK_ARC_1_0/temp4[43] ,
         \MC_ARK_ARC_1_0/temp4[42] , \MC_ARK_ARC_1_0/temp4[41] ,
         \MC_ARK_ARC_1_0/temp4[40] , \MC_ARK_ARC_1_0/temp4[39] ,
         \MC_ARK_ARC_1_0/temp4[37] , \MC_ARK_ARC_1_0/temp4[36] ,
         \MC_ARK_ARC_1_0/temp4[35] , \MC_ARK_ARC_1_0/temp4[33] ,
         \MC_ARK_ARC_1_0/temp4[31] , \MC_ARK_ARC_1_0/temp4[28] ,
         \MC_ARK_ARC_1_0/temp4[27] , \MC_ARK_ARC_1_0/temp4[25] ,
         \MC_ARK_ARC_1_0/temp4[24] , \MC_ARK_ARC_1_0/temp4[23] ,
         \MC_ARK_ARC_1_0/temp4[22] , \MC_ARK_ARC_1_0/temp4[21] ,
         \MC_ARK_ARC_1_0/temp4[19] , \MC_ARK_ARC_1_0/temp4[18] ,
         \MC_ARK_ARC_1_0/temp4[16] , \MC_ARK_ARC_1_0/temp4[15] ,
         \MC_ARK_ARC_1_0/temp4[14] , \MC_ARK_ARC_1_0/temp4[13] ,
         \MC_ARK_ARC_1_0/temp4[12] , \MC_ARK_ARC_1_0/temp4[11] ,
         \MC_ARK_ARC_1_0/temp4[10] , \MC_ARK_ARC_1_0/temp4[9] ,
         \MC_ARK_ARC_1_0/temp4[8] , \MC_ARK_ARC_1_0/temp4[7] ,
         \MC_ARK_ARC_1_0/temp4[6] , \MC_ARK_ARC_1_0/temp4[5] ,
         \MC_ARK_ARC_1_0/temp4[4] , \MC_ARK_ARC_1_0/temp4[3] ,
         \MC_ARK_ARC_1_0/temp4[2] , \MC_ARK_ARC_1_0/temp4[1] ,
         \MC_ARK_ARC_1_0/temp4[0] , \MC_ARK_ARC_1_0/temp3[191] ,
         \MC_ARK_ARC_1_0/temp3[190] , \MC_ARK_ARC_1_0/temp3[189] ,
         \MC_ARK_ARC_1_0/temp3[188] , \MC_ARK_ARC_1_0/temp3[187] ,
         \MC_ARK_ARC_1_0/temp3[186] , \MC_ARK_ARC_1_0/temp3[185] ,
         \MC_ARK_ARC_1_0/temp3[184] , \MC_ARK_ARC_1_0/temp3[183] ,
         \MC_ARK_ARC_1_0/temp3[182] , \MC_ARK_ARC_1_0/temp3[181] ,
         \MC_ARK_ARC_1_0/temp3[180] , \MC_ARK_ARC_1_0/temp3[178] ,
         \MC_ARK_ARC_1_0/temp3[177] , \MC_ARK_ARC_1_0/temp3[174] ,
         \MC_ARK_ARC_1_0/temp3[173] , \MC_ARK_ARC_1_0/temp3[172] ,
         \MC_ARK_ARC_1_0/temp3[171] , \MC_ARK_ARC_1_0/temp3[170] ,
         \MC_ARK_ARC_1_0/temp3[169] , \MC_ARK_ARC_1_0/temp3[168] ,
         \MC_ARK_ARC_1_0/temp3[167] , \MC_ARK_ARC_1_0/temp3[165] ,
         \MC_ARK_ARC_1_0/temp3[163] , \MC_ARK_ARC_1_0/temp3[162] ,
         \MC_ARK_ARC_1_0/temp3[161] , \MC_ARK_ARC_1_0/temp3[160] ,
         \MC_ARK_ARC_1_0/temp3[159] , \MC_ARK_ARC_1_0/temp3[158] ,
         \MC_ARK_ARC_1_0/temp3[157] , \MC_ARK_ARC_1_0/temp3[156] ,
         \MC_ARK_ARC_1_0/temp3[154] , \MC_ARK_ARC_1_0/temp3[153] ,
         \MC_ARK_ARC_1_0/temp3[151] , \MC_ARK_ARC_1_0/temp3[150] ,
         \MC_ARK_ARC_1_0/temp3[149] , \MC_ARK_ARC_1_0/temp3[148] ,
         \MC_ARK_ARC_1_0/temp3[147] , \MC_ARK_ARC_1_0/temp3[145] ,
         \MC_ARK_ARC_1_0/temp3[144] , \MC_ARK_ARC_1_0/temp3[143] ,
         \MC_ARK_ARC_1_0/temp3[139] , \MC_ARK_ARC_1_0/temp3[138] ,
         \MC_ARK_ARC_1_0/temp3[137] , \MC_ARK_ARC_1_0/temp3[136] ,
         \MC_ARK_ARC_1_0/temp3[135] , \MC_ARK_ARC_1_0/temp3[133] ,
         \MC_ARK_ARC_1_0/temp3[130] , \MC_ARK_ARC_1_0/temp3[129] ,
         \MC_ARK_ARC_1_0/temp3[128] , \MC_ARK_ARC_1_0/temp3[127] ,
         \MC_ARK_ARC_1_0/temp3[126] , \MC_ARK_ARC_1_0/temp3[124] ,
         \MC_ARK_ARC_1_0/temp3[123] , \MC_ARK_ARC_1_0/temp3[122] ,
         \MC_ARK_ARC_1_0/temp3[121] , \MC_ARK_ARC_1_0/temp3[120] ,
         \MC_ARK_ARC_1_0/temp3[119] , \MC_ARK_ARC_1_0/temp3[118] ,
         \MC_ARK_ARC_1_0/temp3[115] , \MC_ARK_ARC_1_0/temp3[114] ,
         \MC_ARK_ARC_1_0/temp3[113] , \MC_ARK_ARC_1_0/temp3[112] ,
         \MC_ARK_ARC_1_0/temp3[111] , \MC_ARK_ARC_1_0/temp3[108] ,
         \MC_ARK_ARC_1_0/temp3[106] , \MC_ARK_ARC_1_0/temp3[104] ,
         \MC_ARK_ARC_1_0/temp3[103] , \MC_ARK_ARC_1_0/temp3[101] ,
         \MC_ARK_ARC_1_0/temp3[100] , \MC_ARK_ARC_1_0/temp3[96] ,
         \MC_ARK_ARC_1_0/temp3[94] , \MC_ARK_ARC_1_0/temp3[93] ,
         \MC_ARK_ARC_1_0/temp3[91] , \MC_ARK_ARC_1_0/temp3[90] ,
         \MC_ARK_ARC_1_0/temp3[88] , \MC_ARK_ARC_1_0/temp3[86] ,
         \MC_ARK_ARC_1_0/temp3[85] , \MC_ARK_ARC_1_0/temp3[84] ,
         \MC_ARK_ARC_1_0/temp3[83] , \MC_ARK_ARC_1_0/temp3[82] ,
         \MC_ARK_ARC_1_0/temp3[81] , \MC_ARK_ARC_1_0/temp3[80] ,
         \MC_ARK_ARC_1_0/temp3[78] , \MC_ARK_ARC_1_0/temp3[77] ,
         \MC_ARK_ARC_1_0/temp3[76] , \MC_ARK_ARC_1_0/temp3[73] ,
         \MC_ARK_ARC_1_0/temp3[72] , \MC_ARK_ARC_1_0/temp3[70] ,
         \MC_ARK_ARC_1_0/temp3[69] , \MC_ARK_ARC_1_0/temp3[68] ,
         \MC_ARK_ARC_1_0/temp3[67] , \MC_ARK_ARC_1_0/temp3[66] ,
         \MC_ARK_ARC_1_0/temp3[64] , \MC_ARK_ARC_1_0/temp3[62] ,
         \MC_ARK_ARC_1_0/temp3[61] , \MC_ARK_ARC_1_0/temp3[60] ,
         \MC_ARK_ARC_1_0/temp3[58] , \MC_ARK_ARC_1_0/temp3[55] ,
         \MC_ARK_ARC_1_0/temp3[54] , \MC_ARK_ARC_1_0/temp3[53] ,
         \MC_ARK_ARC_1_0/temp3[52] , \MC_ARK_ARC_1_0/temp3[49] ,
         \MC_ARK_ARC_1_0/temp3[48] , \MC_ARK_ARC_1_0/temp3[46] ,
         \MC_ARK_ARC_1_0/temp3[45] , \MC_ARK_ARC_1_0/temp3[44] ,
         \MC_ARK_ARC_1_0/temp3[42] , \MC_ARK_ARC_1_0/temp3[41] ,
         \MC_ARK_ARC_1_0/temp3[40] , \MC_ARK_ARC_1_0/temp3[39] ,
         \MC_ARK_ARC_1_0/temp3[37] , \MC_ARK_ARC_1_0/temp3[36] ,
         \MC_ARK_ARC_1_0/temp3[35] , \MC_ARK_ARC_1_0/temp3[33] ,
         \MC_ARK_ARC_1_0/temp3[31] , \MC_ARK_ARC_1_0/temp3[27] ,
         \MC_ARK_ARC_1_0/temp3[25] , \MC_ARK_ARC_1_0/temp3[24] ,
         \MC_ARK_ARC_1_0/temp3[23] , \MC_ARK_ARC_1_0/temp3[22] ,
         \MC_ARK_ARC_1_0/temp3[21] , \MC_ARK_ARC_1_0/temp3[19] ,
         \MC_ARK_ARC_1_0/temp3[18] , \MC_ARK_ARC_1_0/temp3[17] ,
         \MC_ARK_ARC_1_0/temp3[16] , \MC_ARK_ARC_1_0/temp3[15] ,
         \MC_ARK_ARC_1_0/temp3[14] , \MC_ARK_ARC_1_0/temp3[13] ,
         \MC_ARK_ARC_1_0/temp3[12] , \MC_ARK_ARC_1_0/temp3[10] ,
         \MC_ARK_ARC_1_0/temp3[8] , \MC_ARK_ARC_1_0/temp3[7] ,
         \MC_ARK_ARC_1_0/temp3[6] , \MC_ARK_ARC_1_0/temp3[5] ,
         \MC_ARK_ARC_1_0/temp3[4] , \MC_ARK_ARC_1_0/temp3[3] ,
         \MC_ARK_ARC_1_0/temp3[2] , \MC_ARK_ARC_1_0/temp3[1] ,
         \MC_ARK_ARC_1_0/temp3[0] , \MC_ARK_ARC_1_0/temp2[191] ,
         \MC_ARK_ARC_1_0/temp2[190] , \MC_ARK_ARC_1_0/temp2[187] ,
         \MC_ARK_ARC_1_0/temp2[186] , \MC_ARK_ARC_1_0/temp2[184] ,
         \MC_ARK_ARC_1_0/temp2[183] , \MC_ARK_ARC_1_0/temp2[182] ,
         \MC_ARK_ARC_1_0/temp2[181] , \MC_ARK_ARC_1_0/temp2[180] ,
         \MC_ARK_ARC_1_0/temp2[178] , \MC_ARK_ARC_1_0/temp2[177] ,
         \MC_ARK_ARC_1_0/temp2[176] , \MC_ARK_ARC_1_0/temp2[175] ,
         \MC_ARK_ARC_1_0/temp2[174] , \MC_ARK_ARC_1_0/temp2[172] ,
         \MC_ARK_ARC_1_0/temp2[170] , \MC_ARK_ARC_1_0/temp2[169] ,
         \MC_ARK_ARC_1_0/temp2[168] , \MC_ARK_ARC_1_0/temp2[166] ,
         \MC_ARK_ARC_1_0/temp2[165] , \MC_ARK_ARC_1_0/temp2[164] ,
         \MC_ARK_ARC_1_0/temp2[163] , \MC_ARK_ARC_1_0/temp2[162] ,
         \MC_ARK_ARC_1_0/temp2[159] , \MC_ARK_ARC_1_0/temp2[158] ,
         \MC_ARK_ARC_1_0/temp2[157] , \MC_ARK_ARC_1_0/temp2[154] ,
         \MC_ARK_ARC_1_0/temp2[151] , \MC_ARK_ARC_1_0/temp2[150] ,
         \MC_ARK_ARC_1_0/temp2[148] , \MC_ARK_ARC_1_0/temp2[147] ,
         \MC_ARK_ARC_1_0/temp2[145] , \MC_ARK_ARC_1_0/temp2[144] ,
         \MC_ARK_ARC_1_0/temp2[141] , \MC_ARK_ARC_1_0/temp2[139] ,
         \MC_ARK_ARC_1_0/temp2[138] , \MC_ARK_ARC_1_0/temp2[137] ,
         \MC_ARK_ARC_1_0/temp2[136] , \MC_ARK_ARC_1_0/temp2[133] ,
         \MC_ARK_ARC_1_0/temp2[132] , \MC_ARK_ARC_1_0/temp2[130] ,
         \MC_ARK_ARC_1_0/temp2[128] , \MC_ARK_ARC_1_0/temp2[127] ,
         \MC_ARK_ARC_1_0/temp2[126] , \MC_ARK_ARC_1_0/temp2[125] ,
         \MC_ARK_ARC_1_0/temp2[124] , \MC_ARK_ARC_1_0/temp2[122] ,
         \MC_ARK_ARC_1_0/temp2[121] , \MC_ARK_ARC_1_0/temp2[120] ,
         \MC_ARK_ARC_1_0/temp2[119] , \MC_ARK_ARC_1_0/temp2[118] ,
         \MC_ARK_ARC_1_0/temp2[117] , \MC_ARK_ARC_1_0/temp2[116] ,
         \MC_ARK_ARC_1_0/temp2[115] , \MC_ARK_ARC_1_0/temp2[114] ,
         \MC_ARK_ARC_1_0/temp2[112] , \MC_ARK_ARC_1_0/temp2[111] ,
         \MC_ARK_ARC_1_0/temp2[110] , \MC_ARK_ARC_1_0/temp2[109] ,
         \MC_ARK_ARC_1_0/temp2[108] , \MC_ARK_ARC_1_0/temp2[106] ,
         \MC_ARK_ARC_1_0/temp2[105] , \MC_ARK_ARC_1_0/temp2[103] ,
         \MC_ARK_ARC_1_0/temp2[101] , \MC_ARK_ARC_1_0/temp2[100] ,
         \MC_ARK_ARC_1_0/temp2[97] , \MC_ARK_ARC_1_0/temp2[96] ,
         \MC_ARK_ARC_1_0/temp2[95] , \MC_ARK_ARC_1_0/temp2[94] ,
         \MC_ARK_ARC_1_0/temp2[93] , \MC_ARK_ARC_1_0/temp2[91] ,
         \MC_ARK_ARC_1_0/temp2[90] , \MC_ARK_ARC_1_0/temp2[87] ,
         \MC_ARK_ARC_1_0/temp2[85] , \MC_ARK_ARC_1_0/temp2[84] ,
         \MC_ARK_ARC_1_0/temp2[83] , \MC_ARK_ARC_1_0/temp2[82] ,
         \MC_ARK_ARC_1_0/temp2[81] , \MC_ARK_ARC_1_0/temp2[79] ,
         \MC_ARK_ARC_1_0/temp2[78] , \MC_ARK_ARC_1_0/temp2[77] ,
         \MC_ARK_ARC_1_0/temp2[76] , \MC_ARK_ARC_1_0/temp2[73] ,
         \MC_ARK_ARC_1_0/temp2[72] , \MC_ARK_ARC_1_0/temp2[71] ,
         \MC_ARK_ARC_1_0/temp2[70] , \MC_ARK_ARC_1_0/temp2[69] ,
         \MC_ARK_ARC_1_0/temp2[67] , \MC_ARK_ARC_1_0/temp2[66] ,
         \MC_ARK_ARC_1_0/temp2[62] , \MC_ARK_ARC_1_0/temp2[61] ,
         \MC_ARK_ARC_1_0/temp2[60] , \MC_ARK_ARC_1_0/temp2[58] ,
         \MC_ARK_ARC_1_0/temp2[56] , \MC_ARK_ARC_1_0/temp2[54] ,
         \MC_ARK_ARC_1_0/temp2[53] , \MC_ARK_ARC_1_0/temp2[52] ,
         \MC_ARK_ARC_1_0/temp2[49] , \MC_ARK_ARC_1_0/temp2[48] ,
         \MC_ARK_ARC_1_0/temp2[47] , \MC_ARK_ARC_1_0/temp2[45] ,
         \MC_ARK_ARC_1_0/temp2[43] , \MC_ARK_ARC_1_0/temp2[42] ,
         \MC_ARK_ARC_1_0/temp2[40] , \MC_ARK_ARC_1_0/temp2[39] ,
         \MC_ARK_ARC_1_0/temp2[37] , \MC_ARK_ARC_1_0/temp2[36] ,
         \MC_ARK_ARC_1_0/temp2[33] , \MC_ARK_ARC_1_0/temp2[32] ,
         \MC_ARK_ARC_1_0/temp2[31] , \MC_ARK_ARC_1_0/temp2[29] ,
         \MC_ARK_ARC_1_0/temp2[28] , \MC_ARK_ARC_1_0/temp2[24] ,
         \MC_ARK_ARC_1_0/temp2[22] , \MC_ARK_ARC_1_0/temp2[19] ,
         \MC_ARK_ARC_1_0/temp2[18] , \MC_ARK_ARC_1_0/temp2[16] ,
         \MC_ARK_ARC_1_0/temp2[15] , \MC_ARK_ARC_1_0/temp2[14] ,
         \MC_ARK_ARC_1_0/temp2[13] , \MC_ARK_ARC_1_0/temp2[10] ,
         \MC_ARK_ARC_1_0/temp2[9] , \MC_ARK_ARC_1_0/temp2[7] ,
         \MC_ARK_ARC_1_0/temp2[6] , \MC_ARK_ARC_1_0/temp2[5] ,
         \MC_ARK_ARC_1_0/temp2[4] , \MC_ARK_ARC_1_0/temp2[1] ,
         \MC_ARK_ARC_1_0/temp2[0] , \MC_ARK_ARC_1_0/temp1[190] ,
         \MC_ARK_ARC_1_0/temp1[188] , \MC_ARK_ARC_1_0/temp1[187] ,
         \MC_ARK_ARC_1_0/temp1[186] , \MC_ARK_ARC_1_0/temp1[185] ,
         \MC_ARK_ARC_1_0/temp1[184] , \MC_ARK_ARC_1_0/temp1[182] ,
         \MC_ARK_ARC_1_0/temp1[181] , \MC_ARK_ARC_1_0/temp1[180] ,
         \MC_ARK_ARC_1_0/temp1[178] , \MC_ARK_ARC_1_0/temp1[177] ,
         \MC_ARK_ARC_1_0/temp1[175] , \MC_ARK_ARC_1_0/temp1[174] ,
         \MC_ARK_ARC_1_0/temp1[172] , \MC_ARK_ARC_1_0/temp1[170] ,
         \MC_ARK_ARC_1_0/temp1[169] , \MC_ARK_ARC_1_0/temp1[168] ,
         \MC_ARK_ARC_1_0/temp1[166] , \MC_ARK_ARC_1_0/temp1[163] ,
         \MC_ARK_ARC_1_0/temp1[162] , \MC_ARK_ARC_1_0/temp1[161] ,
         \MC_ARK_ARC_1_0/temp1[160] , \MC_ARK_ARC_1_0/temp1[158] ,
         \MC_ARK_ARC_1_0/temp1[157] , \MC_ARK_ARC_1_0/temp1[156] ,
         \MC_ARK_ARC_1_0/temp1[154] , \MC_ARK_ARC_1_0/temp1[151] ,
         \MC_ARK_ARC_1_0/temp1[148] , \MC_ARK_ARC_1_0/temp1[146] ,
         \MC_ARK_ARC_1_0/temp1[145] , \MC_ARK_ARC_1_0/temp1[144] ,
         \MC_ARK_ARC_1_0/temp1[143] , \MC_ARK_ARC_1_0/temp1[142] ,
         \MC_ARK_ARC_1_0/temp1[141] , \MC_ARK_ARC_1_0/temp1[139] ,
         \MC_ARK_ARC_1_0/temp1[138] , \MC_ARK_ARC_1_0/temp1[136] ,
         \MC_ARK_ARC_1_0/temp1[133] , \MC_ARK_ARC_1_0/temp1[131] ,
         \MC_ARK_ARC_1_0/temp1[130] , \MC_ARK_ARC_1_0/temp1[129] ,
         \MC_ARK_ARC_1_0/temp1[128] , \MC_ARK_ARC_1_0/temp1[127] ,
         \MC_ARK_ARC_1_0/temp1[126] , \MC_ARK_ARC_1_0/temp1[125] ,
         \MC_ARK_ARC_1_0/temp1[122] , \MC_ARK_ARC_1_0/temp1[121] ,
         \MC_ARK_ARC_1_0/temp1[120] , \MC_ARK_ARC_1_0/temp1[119] ,
         \MC_ARK_ARC_1_0/temp1[118] , \MC_ARK_ARC_1_0/temp1[116] ,
         \MC_ARK_ARC_1_0/temp1[115] , \MC_ARK_ARC_1_0/temp1[114] ,
         \MC_ARK_ARC_1_0/temp1[112] , \MC_ARK_ARC_1_0/temp1[111] ,
         \MC_ARK_ARC_1_0/temp1[110] , \MC_ARK_ARC_1_0/temp1[109] ,
         \MC_ARK_ARC_1_0/temp1[108] , \MC_ARK_ARC_1_0/temp1[106] ,
         \MC_ARK_ARC_1_0/temp1[105] , \MC_ARK_ARC_1_0/temp1[103] ,
         \MC_ARK_ARC_1_0/temp1[101] , \MC_ARK_ARC_1_0/temp1[100] ,
         \MC_ARK_ARC_1_0/temp1[99] , \MC_ARK_ARC_1_0/temp1[98] ,
         \MC_ARK_ARC_1_0/temp1[97] , \MC_ARK_ARC_1_0/temp1[96] ,
         \MC_ARK_ARC_1_0/temp1[94] , \MC_ARK_ARC_1_0/temp1[91] ,
         \MC_ARK_ARC_1_0/temp1[90] , \MC_ARK_ARC_1_0/temp1[89] ,
         \MC_ARK_ARC_1_0/temp1[88] , \MC_ARK_ARC_1_0/temp1[86] ,
         \MC_ARK_ARC_1_0/temp1[85] , \MC_ARK_ARC_1_0/temp1[84] ,
         \MC_ARK_ARC_1_0/temp1[83] , \MC_ARK_ARC_1_0/temp1[82] ,
         \MC_ARK_ARC_1_0/temp1[79] , \MC_ARK_ARC_1_0/temp1[78] ,
         \MC_ARK_ARC_1_0/temp1[77] , \MC_ARK_ARC_1_0/temp1[76] ,
         \MC_ARK_ARC_1_0/temp1[75] , \MC_ARK_ARC_1_0/temp1[74] ,
         \MC_ARK_ARC_1_0/temp1[73] , \MC_ARK_ARC_1_0/temp1[72] ,
         \MC_ARK_ARC_1_0/temp1[71] , \MC_ARK_ARC_1_0/temp1[70] ,
         \MC_ARK_ARC_1_0/temp1[69] , \MC_ARK_ARC_1_0/temp1[67] ,
         \MC_ARK_ARC_1_0/temp1[62] , \MC_ARK_ARC_1_0/temp1[60] ,
         \MC_ARK_ARC_1_0/temp1[58] , \MC_ARK_ARC_1_0/temp1[57] ,
         \MC_ARK_ARC_1_0/temp1[55] , \MC_ARK_ARC_1_0/temp1[54] ,
         \MC_ARK_ARC_1_0/temp1[53] , \MC_ARK_ARC_1_0/temp1[49] ,
         \MC_ARK_ARC_1_0/temp1[48] , \MC_ARK_ARC_1_0/temp1[46] ,
         \MC_ARK_ARC_1_0/temp1[45] , \MC_ARK_ARC_1_0/temp1[44] ,
         \MC_ARK_ARC_1_0/temp1[42] , \MC_ARK_ARC_1_0/temp1[41] ,
         \MC_ARK_ARC_1_0/temp1[37] , \MC_ARK_ARC_1_0/temp1[36] ,
         \MC_ARK_ARC_1_0/temp1[33] , \MC_ARK_ARC_1_0/temp1[32] ,
         \MC_ARK_ARC_1_0/temp1[31] , \MC_ARK_ARC_1_0/temp1[28] ,
         \MC_ARK_ARC_1_0/temp1[25] , \MC_ARK_ARC_1_0/temp1[24] ,
         \MC_ARK_ARC_1_0/temp1[23] , \MC_ARK_ARC_1_0/temp1[22] ,
         \MC_ARK_ARC_1_0/temp1[21] , \MC_ARK_ARC_1_0/temp1[19] ,
         \MC_ARK_ARC_1_0/temp1[18] , \MC_ARK_ARC_1_0/temp1[17] ,
         \MC_ARK_ARC_1_0/temp1[16] , \MC_ARK_ARC_1_0/temp1[15] ,
         \MC_ARK_ARC_1_0/temp1[14] , \MC_ARK_ARC_1_0/temp1[13] ,
         \MC_ARK_ARC_1_0/temp1[12] , \MC_ARK_ARC_1_0/temp1[10] ,
         \MC_ARK_ARC_1_0/temp1[8] , \MC_ARK_ARC_1_0/temp1[7] ,
         \MC_ARK_ARC_1_0/temp1[6] , \MC_ARK_ARC_1_0/temp1[5] ,
         \MC_ARK_ARC_1_0/temp1[4] , \MC_ARK_ARC_1_0/temp1[3] ,
         \MC_ARK_ARC_1_0/temp1[1] , \MC_ARK_ARC_1_0/buf_keyinput[92] ,
         \MC_ARK_ARC_1_0/buf_keyinput[71] , \MC_ARK_ARC_1_0/buf_keyinput[57] ,
         \MC_ARK_ARC_1_0/buf_datainput[173] ,
         \MC_ARK_ARC_1_0/buf_datainput[149] ,
         \MC_ARK_ARC_1_0/buf_datainput[139] ,
         \MC_ARK_ARC_1_0/buf_datainput[137] ,
         \MC_ARK_ARC_1_0/buf_datainput[113] ,
         \MC_ARK_ARC_1_0/buf_datainput[108] ,
         \MC_ARK_ARC_1_0/buf_datainput[102] ,
         \MC_ARK_ARC_1_0/buf_datainput[97] ,
         \MC_ARK_ARC_1_0/buf_datainput[84] ,
         \MC_ARK_ARC_1_0/buf_datainput[77] ,
         \MC_ARK_ARC_1_0/buf_datainput[75] ,
         \MC_ARK_ARC_1_0/buf_datainput[71] ,
         \MC_ARK_ARC_1_0/buf_datainput[70] ,
         \MC_ARK_ARC_1_0/buf_datainput[67] ,
         \MC_ARK_ARC_1_0/buf_datainput[64] ,
         \MC_ARK_ARC_1_0/buf_datainput[43] ,
         \MC_ARK_ARC_1_0/buf_datainput[41] ,
         \MC_ARK_ARC_1_0/buf_datainput[35] ,
         \MC_ARK_ARC_1_0/buf_datainput[31] , \MC_ARK_ARC_1_1/buf_output[191] ,
         \MC_ARK_ARC_1_1/buf_output[190] , \MC_ARK_ARC_1_1/buf_output[189] ,
         \MC_ARK_ARC_1_1/buf_output[188] , \MC_ARK_ARC_1_1/buf_output[187] ,
         \MC_ARK_ARC_1_1/buf_output[186] , \MC_ARK_ARC_1_1/buf_output[184] ,
         \MC_ARK_ARC_1_1/buf_output[183] , \MC_ARK_ARC_1_1/buf_output[182] ,
         \MC_ARK_ARC_1_1/buf_output[181] , \MC_ARK_ARC_1_1/buf_output[180] ,
         \MC_ARK_ARC_1_1/buf_output[179] , \MC_ARK_ARC_1_1/buf_output[178] ,
         \MC_ARK_ARC_1_1/buf_output[177] , \MC_ARK_ARC_1_1/buf_output[176] ,
         \MC_ARK_ARC_1_1/buf_output[175] , \MC_ARK_ARC_1_1/buf_output[174] ,
         \MC_ARK_ARC_1_1/buf_output[173] , \MC_ARK_ARC_1_1/buf_output[172] ,
         \MC_ARK_ARC_1_1/buf_output[171] , \MC_ARK_ARC_1_1/buf_output[170] ,
         \MC_ARK_ARC_1_1/buf_output[169] , \MC_ARK_ARC_1_1/buf_output[168] ,
         \MC_ARK_ARC_1_1/buf_output[167] , \MC_ARK_ARC_1_1/buf_output[166] ,
         \MC_ARK_ARC_1_1/buf_output[165] , \MC_ARK_ARC_1_1/buf_output[164] ,
         \MC_ARK_ARC_1_1/buf_output[163] , \MC_ARK_ARC_1_1/buf_output[162] ,
         \MC_ARK_ARC_1_1/buf_output[161] , \MC_ARK_ARC_1_1/buf_output[160] ,
         \MC_ARK_ARC_1_1/buf_output[159] , \MC_ARK_ARC_1_1/buf_output[158] ,
         \MC_ARK_ARC_1_1/buf_output[157] , \MC_ARK_ARC_1_1/buf_output[156] ,
         \MC_ARK_ARC_1_1/buf_output[155] , \MC_ARK_ARC_1_1/buf_output[154] ,
         \MC_ARK_ARC_1_1/buf_output[153] , \MC_ARK_ARC_1_1/buf_output[152] ,
         \MC_ARK_ARC_1_1/buf_output[151] , \MC_ARK_ARC_1_1/buf_output[150] ,
         \MC_ARK_ARC_1_1/buf_output[149] , \MC_ARK_ARC_1_1/buf_output[148] ,
         \MC_ARK_ARC_1_1/buf_output[147] , \MC_ARK_ARC_1_1/buf_output[146] ,
         \MC_ARK_ARC_1_1/buf_output[145] , \MC_ARK_ARC_1_1/buf_output[144] ,
         \MC_ARK_ARC_1_1/buf_output[143] , \MC_ARK_ARC_1_1/buf_output[142] ,
         \MC_ARK_ARC_1_1/buf_output[141] , \MC_ARK_ARC_1_1/buf_output[140] ,
         \MC_ARK_ARC_1_1/buf_output[139] , \MC_ARK_ARC_1_1/buf_output[138] ,
         \MC_ARK_ARC_1_1/buf_output[137] , \MC_ARK_ARC_1_1/buf_output[136] ,
         \MC_ARK_ARC_1_1/buf_output[135] , \MC_ARK_ARC_1_1/buf_output[134] ,
         \MC_ARK_ARC_1_1/buf_output[133] , \MC_ARK_ARC_1_1/buf_output[132] ,
         \MC_ARK_ARC_1_1/buf_output[131] , \MC_ARK_ARC_1_1/buf_output[130] ,
         \MC_ARK_ARC_1_1/buf_output[129] , \MC_ARK_ARC_1_1/buf_output[128] ,
         \MC_ARK_ARC_1_1/buf_output[127] , \MC_ARK_ARC_1_1/buf_output[126] ,
         \MC_ARK_ARC_1_1/buf_output[124] , \MC_ARK_ARC_1_1/buf_output[123] ,
         \MC_ARK_ARC_1_1/buf_output[122] , \MC_ARK_ARC_1_1/buf_output[121] ,
         \MC_ARK_ARC_1_1/buf_output[120] , \MC_ARK_ARC_1_1/buf_output[119] ,
         \MC_ARK_ARC_1_1/buf_output[118] , \MC_ARK_ARC_1_1/buf_output[117] ,
         \MC_ARK_ARC_1_1/buf_output[116] , \MC_ARK_ARC_1_1/buf_output[115] ,
         \MC_ARK_ARC_1_1/buf_output[114] , \MC_ARK_ARC_1_1/buf_output[113] ,
         \MC_ARK_ARC_1_1/buf_output[112] , \MC_ARK_ARC_1_1/buf_output[111] ,
         \MC_ARK_ARC_1_1/buf_output[110] , \MC_ARK_ARC_1_1/buf_output[109] ,
         \MC_ARK_ARC_1_1/buf_output[108] , \MC_ARK_ARC_1_1/buf_output[107] ,
         \MC_ARK_ARC_1_1/buf_output[106] , \MC_ARK_ARC_1_1/buf_output[105] ,
         \MC_ARK_ARC_1_1/buf_output[104] , \MC_ARK_ARC_1_1/buf_output[103] ,
         \MC_ARK_ARC_1_1/buf_output[102] , \MC_ARK_ARC_1_1/buf_output[101] ,
         \MC_ARK_ARC_1_1/buf_output[100] , \MC_ARK_ARC_1_1/buf_output[99] ,
         \MC_ARK_ARC_1_1/buf_output[98] , \MC_ARK_ARC_1_1/buf_output[97] ,
         \MC_ARK_ARC_1_1/buf_output[96] , \MC_ARK_ARC_1_1/buf_output[95] ,
         \MC_ARK_ARC_1_1/buf_output[94] , \MC_ARK_ARC_1_1/buf_output[93] ,
         \MC_ARK_ARC_1_1/buf_output[92] , \MC_ARK_ARC_1_1/buf_output[91] ,
         \MC_ARK_ARC_1_1/buf_output[90] , \MC_ARK_ARC_1_1/buf_output[89] ,
         \MC_ARK_ARC_1_1/buf_output[88] , \MC_ARK_ARC_1_1/buf_output[87] ,
         \MC_ARK_ARC_1_1/buf_output[86] , \MC_ARK_ARC_1_1/buf_output[85] ,
         \MC_ARK_ARC_1_1/buf_output[84] , \MC_ARK_ARC_1_1/buf_output[83] ,
         \MC_ARK_ARC_1_1/buf_output[82] , \MC_ARK_ARC_1_1/buf_output[81] ,
         \MC_ARK_ARC_1_1/buf_output[80] , \MC_ARK_ARC_1_1/buf_output[79] ,
         \MC_ARK_ARC_1_1/buf_output[78] , \MC_ARK_ARC_1_1/buf_output[77] ,
         \MC_ARK_ARC_1_1/buf_output[76] , \MC_ARK_ARC_1_1/buf_output[75] ,
         \MC_ARK_ARC_1_1/buf_output[74] , \MC_ARK_ARC_1_1/buf_output[73] ,
         \MC_ARK_ARC_1_1/buf_output[72] , \MC_ARK_ARC_1_1/buf_output[71] ,
         \MC_ARK_ARC_1_1/buf_output[70] , \MC_ARK_ARC_1_1/buf_output[69] ,
         \MC_ARK_ARC_1_1/buf_output[68] , \MC_ARK_ARC_1_1/buf_output[67] ,
         \MC_ARK_ARC_1_1/buf_output[66] , \MC_ARK_ARC_1_1/buf_output[65] ,
         \MC_ARK_ARC_1_1/buf_output[64] , \MC_ARK_ARC_1_1/buf_output[63] ,
         \MC_ARK_ARC_1_1/buf_output[62] , \MC_ARK_ARC_1_1/buf_output[61] ,
         \MC_ARK_ARC_1_1/buf_output[60] , \MC_ARK_ARC_1_1/buf_output[59] ,
         \MC_ARK_ARC_1_1/buf_output[58] , \MC_ARK_ARC_1_1/buf_output[57] ,
         \MC_ARK_ARC_1_1/buf_output[56] , \MC_ARK_ARC_1_1/buf_output[55] ,
         \MC_ARK_ARC_1_1/buf_output[53] , \MC_ARK_ARC_1_1/buf_output[52] ,
         \MC_ARK_ARC_1_1/buf_output[51] , \MC_ARK_ARC_1_1/buf_output[50] ,
         \MC_ARK_ARC_1_1/buf_output[49] , \MC_ARK_ARC_1_1/buf_output[48] ,
         \MC_ARK_ARC_1_1/buf_output[47] , \MC_ARK_ARC_1_1/buf_output[46] ,
         \MC_ARK_ARC_1_1/buf_output[45] , \MC_ARK_ARC_1_1/buf_output[44] ,
         \MC_ARK_ARC_1_1/buf_output[43] , \MC_ARK_ARC_1_1/buf_output[42] ,
         \MC_ARK_ARC_1_1/buf_output[41] , \MC_ARK_ARC_1_1/buf_output[40] ,
         \MC_ARK_ARC_1_1/buf_output[39] , \MC_ARK_ARC_1_1/buf_output[38] ,
         \MC_ARK_ARC_1_1/buf_output[37] , \MC_ARK_ARC_1_1/buf_output[36] ,
         \MC_ARK_ARC_1_1/buf_output[35] , \MC_ARK_ARC_1_1/buf_output[34] ,
         \MC_ARK_ARC_1_1/buf_output[33] , \MC_ARK_ARC_1_1/buf_output[32] ,
         \MC_ARK_ARC_1_1/buf_output[31] , \MC_ARK_ARC_1_1/buf_output[30] ,
         \MC_ARK_ARC_1_1/buf_output[29] , \MC_ARK_ARC_1_1/buf_output[28] ,
         \MC_ARK_ARC_1_1/buf_output[27] , \MC_ARK_ARC_1_1/buf_output[26] ,
         \MC_ARK_ARC_1_1/buf_output[25] , \MC_ARK_ARC_1_1/buf_output[24] ,
         \MC_ARK_ARC_1_1/buf_output[23] , \MC_ARK_ARC_1_1/buf_output[22] ,
         \MC_ARK_ARC_1_1/buf_output[21] , \MC_ARK_ARC_1_1/buf_output[20] ,
         \MC_ARK_ARC_1_1/buf_output[19] , \MC_ARK_ARC_1_1/buf_output[18] ,
         \MC_ARK_ARC_1_1/buf_output[17] , \MC_ARK_ARC_1_1/buf_output[16] ,
         \MC_ARK_ARC_1_1/buf_output[15] , \MC_ARK_ARC_1_1/buf_output[14] ,
         \MC_ARK_ARC_1_1/buf_output[13] , \MC_ARK_ARC_1_1/buf_output[12] ,
         \MC_ARK_ARC_1_1/buf_output[11] , \MC_ARK_ARC_1_1/buf_output[10] ,
         \MC_ARK_ARC_1_1/buf_output[8] , \MC_ARK_ARC_1_1/buf_output[7] ,
         \MC_ARK_ARC_1_1/buf_output[6] , \MC_ARK_ARC_1_1/buf_output[4] ,
         \MC_ARK_ARC_1_1/buf_output[3] , \MC_ARK_ARC_1_1/buf_output[2] ,
         \MC_ARK_ARC_1_1/buf_output[1] , \MC_ARK_ARC_1_1/buf_output[0] ,
         \MC_ARK_ARC_1_1/temp6[186] , \MC_ARK_ARC_1_1/temp6[185] ,
         \MC_ARK_ARC_1_1/temp6[183] , \MC_ARK_ARC_1_1/temp6[180] ,
         \MC_ARK_ARC_1_1/temp6[178] , \MC_ARK_ARC_1_1/temp6[177] ,
         \MC_ARK_ARC_1_1/temp6[175] , \MC_ARK_ARC_1_1/temp6[174] ,
         \MC_ARK_ARC_1_1/temp6[169] , \MC_ARK_ARC_1_1/temp6[164] ,
         \MC_ARK_ARC_1_1/temp6[163] , \MC_ARK_ARC_1_1/temp6[162] ,
         \MC_ARK_ARC_1_1/temp6[160] , \MC_ARK_ARC_1_1/temp6[158] ,
         \MC_ARK_ARC_1_1/temp6[157] , \MC_ARK_ARC_1_1/temp6[155] ,
         \MC_ARK_ARC_1_1/temp6[154] , \MC_ARK_ARC_1_1/temp6[153] ,
         \MC_ARK_ARC_1_1/temp6[152] , \MC_ARK_ARC_1_1/temp6[151] ,
         \MC_ARK_ARC_1_1/temp6[150] , \MC_ARK_ARC_1_1/temp6[148] ,
         \MC_ARK_ARC_1_1/temp6[145] , \MC_ARK_ARC_1_1/temp6[143] ,
         \MC_ARK_ARC_1_1/temp6[142] , \MC_ARK_ARC_1_1/temp6[140] ,
         \MC_ARK_ARC_1_1/temp6[139] , \MC_ARK_ARC_1_1/temp6[138] ,
         \MC_ARK_ARC_1_1/temp6[136] , \MC_ARK_ARC_1_1/temp6[135] ,
         \MC_ARK_ARC_1_1/temp6[129] , \MC_ARK_ARC_1_1/temp6[126] ,
         \MC_ARK_ARC_1_1/temp6[125] , \MC_ARK_ARC_1_1/temp6[124] ,
         \MC_ARK_ARC_1_1/temp6[119] , \MC_ARK_ARC_1_1/temp6[118] ,
         \MC_ARK_ARC_1_1/temp6[114] , \MC_ARK_ARC_1_1/temp6[111] ,
         \MC_ARK_ARC_1_1/temp6[110] , \MC_ARK_ARC_1_1/temp6[108] ,
         \MC_ARK_ARC_1_1/temp6[107] , \MC_ARK_ARC_1_1/temp6[106] ,
         \MC_ARK_ARC_1_1/temp6[105] , \MC_ARK_ARC_1_1/temp6[102] ,
         \MC_ARK_ARC_1_1/temp6[100] , \MC_ARK_ARC_1_1/temp6[99] ,
         \MC_ARK_ARC_1_1/temp6[98] , \MC_ARK_ARC_1_1/temp6[97] ,
         \MC_ARK_ARC_1_1/temp6[94] , \MC_ARK_ARC_1_1/temp6[92] ,
         \MC_ARK_ARC_1_1/temp6[89] , \MC_ARK_ARC_1_1/temp6[88] ,
         \MC_ARK_ARC_1_1/temp6[87] , \MC_ARK_ARC_1_1/temp6[86] ,
         \MC_ARK_ARC_1_1/temp6[85] , \MC_ARK_ARC_1_1/temp6[79] ,
         \MC_ARK_ARC_1_1/temp6[76] , \MC_ARK_ARC_1_1/temp6[72] ,
         \MC_ARK_ARC_1_1/temp6[70] , \MC_ARK_ARC_1_1/temp6[68] ,
         \MC_ARK_ARC_1_1/temp6[67] , \MC_ARK_ARC_1_1/temp6[66] ,
         \MC_ARK_ARC_1_1/temp6[65] , \MC_ARK_ARC_1_1/temp6[62] ,
         \MC_ARK_ARC_1_1/temp6[61] , \MC_ARK_ARC_1_1/temp6[58] ,
         \MC_ARK_ARC_1_1/temp6[53] , \MC_ARK_ARC_1_1/temp6[52] ,
         \MC_ARK_ARC_1_1/temp6[48] , \MC_ARK_ARC_1_1/temp6[46] ,
         \MC_ARK_ARC_1_1/temp6[40] , \MC_ARK_ARC_1_1/temp6[39] ,
         \MC_ARK_ARC_1_1/temp6[37] , \MC_ARK_ARC_1_1/temp6[36] ,
         \MC_ARK_ARC_1_1/temp6[35] , \MC_ARK_ARC_1_1/temp6[34] ,
         \MC_ARK_ARC_1_1/temp6[32] , \MC_ARK_ARC_1_1/temp6[30] ,
         \MC_ARK_ARC_1_1/temp6[28] , \MC_ARK_ARC_1_1/temp6[25] ,
         \MC_ARK_ARC_1_1/temp6[22] , \MC_ARK_ARC_1_1/temp6[21] ,
         \MC_ARK_ARC_1_1/temp6[20] , \MC_ARK_ARC_1_1/temp6[19] ,
         \MC_ARK_ARC_1_1/temp6[18] , \MC_ARK_ARC_1_1/temp6[16] ,
         \MC_ARK_ARC_1_1/temp6[15] , \MC_ARK_ARC_1_1/temp6[13] ,
         \MC_ARK_ARC_1_1/temp6[12] , \MC_ARK_ARC_1_1/temp6[11] ,
         \MC_ARK_ARC_1_1/temp6[9] , \MC_ARK_ARC_1_1/temp6[4] ,
         \MC_ARK_ARC_1_1/temp6[3] , \MC_ARK_ARC_1_1/temp6[1] ,
         \MC_ARK_ARC_1_1/temp6[0] , \MC_ARK_ARC_1_1/temp5[190] ,
         \MC_ARK_ARC_1_1/temp5[189] , \MC_ARK_ARC_1_1/temp5[184] ,
         \MC_ARK_ARC_1_1/temp5[181] , \MC_ARK_ARC_1_1/temp5[178] ,
         \MC_ARK_ARC_1_1/temp5[177] , \MC_ARK_ARC_1_1/temp5[174] ,
         \MC_ARK_ARC_1_1/temp5[171] , \MC_ARK_ARC_1_1/temp5[170] ,
         \MC_ARK_ARC_1_1/temp5[169] , \MC_ARK_ARC_1_1/temp5[166] ,
         \MC_ARK_ARC_1_1/temp5[163] , \MC_ARK_ARC_1_1/temp5[162] ,
         \MC_ARK_ARC_1_1/temp5[161] , \MC_ARK_ARC_1_1/temp5[156] ,
         \MC_ARK_ARC_1_1/temp5[155] , \MC_ARK_ARC_1_1/temp5[152] ,
         \MC_ARK_ARC_1_1/temp5[151] , \MC_ARK_ARC_1_1/temp5[150] ,
         \MC_ARK_ARC_1_1/temp5[146] , \MC_ARK_ARC_1_1/temp5[144] ,
         \MC_ARK_ARC_1_1/temp5[143] , \MC_ARK_ARC_1_1/temp5[142] ,
         \MC_ARK_ARC_1_1/temp5[139] , \MC_ARK_ARC_1_1/temp5[136] ,
         \MC_ARK_ARC_1_1/temp5[135] , \MC_ARK_ARC_1_1/temp5[133] ,
         \MC_ARK_ARC_1_1/temp5[131] , \MC_ARK_ARC_1_1/temp5[130] ,
         \MC_ARK_ARC_1_1/temp5[129] , \MC_ARK_ARC_1_1/temp5[126] ,
         \MC_ARK_ARC_1_1/temp5[125] , \MC_ARK_ARC_1_1/temp5[123] ,
         \MC_ARK_ARC_1_1/temp5[122] , \MC_ARK_ARC_1_1/temp5[119] ,
         \MC_ARK_ARC_1_1/temp5[118] , \MC_ARK_ARC_1_1/temp5[114] ,
         \MC_ARK_ARC_1_1/temp5[111] , \MC_ARK_ARC_1_1/temp5[108] ,
         \MC_ARK_ARC_1_1/temp5[105] , \MC_ARK_ARC_1_1/temp5[102] ,
         \MC_ARK_ARC_1_1/temp5[101] , \MC_ARK_ARC_1_1/temp5[100] ,
         \MC_ARK_ARC_1_1/temp5[99] , \MC_ARK_ARC_1_1/temp5[97] ,
         \MC_ARK_ARC_1_1/temp5[96] , \MC_ARK_ARC_1_1/temp5[94] ,
         \MC_ARK_ARC_1_1/temp5[93] , \MC_ARK_ARC_1_1/temp5[90] ,
         \MC_ARK_ARC_1_1/temp5[89] , \MC_ARK_ARC_1_1/temp5[87] ,
         \MC_ARK_ARC_1_1/temp5[85] , \MC_ARK_ARC_1_1/temp5[84] ,
         \MC_ARK_ARC_1_1/temp5[83] , \MC_ARK_ARC_1_1/temp5[80] ,
         \MC_ARK_ARC_1_1/temp5[79] , \MC_ARK_ARC_1_1/temp5[78] ,
         \MC_ARK_ARC_1_1/temp5[77] , \MC_ARK_ARC_1_1/temp5[76] ,
         \MC_ARK_ARC_1_1/temp5[74] , \MC_ARK_ARC_1_1/temp5[73] ,
         \MC_ARK_ARC_1_1/temp5[72] , \MC_ARK_ARC_1_1/temp5[70] ,
         \MC_ARK_ARC_1_1/temp5[68] , \MC_ARK_ARC_1_1/temp5[67] ,
         \MC_ARK_ARC_1_1/temp5[66] , \MC_ARK_ARC_1_1/temp5[65] ,
         \MC_ARK_ARC_1_1/temp5[64] , \MC_ARK_ARC_1_1/temp5[62] ,
         \MC_ARK_ARC_1_1/temp5[61] , \MC_ARK_ARC_1_1/temp5[60] ,
         \MC_ARK_ARC_1_1/temp5[58] , \MC_ARK_ARC_1_1/temp5[53] ,
         \MC_ARK_ARC_1_1/temp5[52] , \MC_ARK_ARC_1_1/temp5[48] ,
         \MC_ARK_ARC_1_1/temp5[46] , \MC_ARK_ARC_1_1/temp5[40] ,
         \MC_ARK_ARC_1_1/temp5[39] , \MC_ARK_ARC_1_1/temp5[36] ,
         \MC_ARK_ARC_1_1/temp5[34] , \MC_ARK_ARC_1_1/temp5[30] ,
         \MC_ARK_ARC_1_1/temp5[28] , \MC_ARK_ARC_1_1/temp5[24] ,
         \MC_ARK_ARC_1_1/temp5[22] , \MC_ARK_ARC_1_1/temp5[19] ,
         \MC_ARK_ARC_1_1/temp5[16] , \MC_ARK_ARC_1_1/temp5[13] ,
         \MC_ARK_ARC_1_1/temp5[12] , \MC_ARK_ARC_1_1/temp5[10] ,
         \MC_ARK_ARC_1_1/temp5[9] , \MC_ARK_ARC_1_1/temp5[8] ,
         \MC_ARK_ARC_1_1/temp5[6] , \MC_ARK_ARC_1_1/temp5[5] ,
         \MC_ARK_ARC_1_1/temp5[4] , \MC_ARK_ARC_1_1/temp5[2] ,
         \MC_ARK_ARC_1_1/temp5[1] , \MC_ARK_ARC_1_1/temp5[0] ,
         \MC_ARK_ARC_1_1/temp4[191] , \MC_ARK_ARC_1_1/temp4[190] ,
         \MC_ARK_ARC_1_1/temp4[189] , \MC_ARK_ARC_1_1/temp4[188] ,
         \MC_ARK_ARC_1_1/temp4[187] , \MC_ARK_ARC_1_1/temp4[186] ,
         \MC_ARK_ARC_1_1/temp4[185] , \MC_ARK_ARC_1_1/temp4[184] ,
         \MC_ARK_ARC_1_1/temp4[183] , \MC_ARK_ARC_1_1/temp4[182] ,
         \MC_ARK_ARC_1_1/temp4[181] , \MC_ARK_ARC_1_1/temp4[180] ,
         \MC_ARK_ARC_1_1/temp4[179] , \MC_ARK_ARC_1_1/temp4[178] ,
         \MC_ARK_ARC_1_1/temp4[177] , \MC_ARK_ARC_1_1/temp4[176] ,
         \MC_ARK_ARC_1_1/temp4[175] , \MC_ARK_ARC_1_1/temp4[174] ,
         \MC_ARK_ARC_1_1/temp4[173] , \MC_ARK_ARC_1_1/temp4[172] ,
         \MC_ARK_ARC_1_1/temp4[171] , \MC_ARK_ARC_1_1/temp4[170] ,
         \MC_ARK_ARC_1_1/temp4[169] , \MC_ARK_ARC_1_1/temp4[168] ,
         \MC_ARK_ARC_1_1/temp4[166] , \MC_ARK_ARC_1_1/temp4[164] ,
         \MC_ARK_ARC_1_1/temp4[163] , \MC_ARK_ARC_1_1/temp4[162] ,
         \MC_ARK_ARC_1_1/temp4[161] , \MC_ARK_ARC_1_1/temp4[160] ,
         \MC_ARK_ARC_1_1/temp4[159] , \MC_ARK_ARC_1_1/temp4[158] ,
         \MC_ARK_ARC_1_1/temp4[157] , \MC_ARK_ARC_1_1/temp4[156] ,
         \MC_ARK_ARC_1_1/temp4[155] , \MC_ARK_ARC_1_1/temp4[154] ,
         \MC_ARK_ARC_1_1/temp4[153] , \MC_ARK_ARC_1_1/temp4[152] ,
         \MC_ARK_ARC_1_1/temp4[151] , \MC_ARK_ARC_1_1/temp4[150] ,
         \MC_ARK_ARC_1_1/temp4[149] , \MC_ARK_ARC_1_1/temp4[148] ,
         \MC_ARK_ARC_1_1/temp4[146] , \MC_ARK_ARC_1_1/temp4[145] ,
         \MC_ARK_ARC_1_1/temp4[144] , \MC_ARK_ARC_1_1/temp4[143] ,
         \MC_ARK_ARC_1_1/temp4[142] , \MC_ARK_ARC_1_1/temp4[141] ,
         \MC_ARK_ARC_1_1/temp4[140] , \MC_ARK_ARC_1_1/temp4[139] ,
         \MC_ARK_ARC_1_1/temp4[138] , \MC_ARK_ARC_1_1/temp4[137] ,
         \MC_ARK_ARC_1_1/temp4[136] , \MC_ARK_ARC_1_1/temp4[133] ,
         \MC_ARK_ARC_1_1/temp4[132] , \MC_ARK_ARC_1_1/temp4[131] ,
         \MC_ARK_ARC_1_1/temp4[130] , \MC_ARK_ARC_1_1/temp4[129] ,
         \MC_ARK_ARC_1_1/temp4[128] , \MC_ARK_ARC_1_1/temp4[127] ,
         \MC_ARK_ARC_1_1/temp4[126] , \MC_ARK_ARC_1_1/temp4[125] ,
         \MC_ARK_ARC_1_1/temp4[124] , \MC_ARK_ARC_1_1/temp4[123] ,
         \MC_ARK_ARC_1_1/temp4[122] , \MC_ARK_ARC_1_1/temp4[121] ,
         \MC_ARK_ARC_1_1/temp4[120] , \MC_ARK_ARC_1_1/temp4[119] ,
         \MC_ARK_ARC_1_1/temp4[118] , \MC_ARK_ARC_1_1/temp4[117] ,
         \MC_ARK_ARC_1_1/temp4[115] , \MC_ARK_ARC_1_1/temp4[114] ,
         \MC_ARK_ARC_1_1/temp4[113] , \MC_ARK_ARC_1_1/temp4[112] ,
         \MC_ARK_ARC_1_1/temp4[111] , \MC_ARK_ARC_1_1/temp4[110] ,
         \MC_ARK_ARC_1_1/temp4[109] , \MC_ARK_ARC_1_1/temp4[108] ,
         \MC_ARK_ARC_1_1/temp4[106] , \MC_ARK_ARC_1_1/temp4[105] ,
         \MC_ARK_ARC_1_1/temp4[104] , \MC_ARK_ARC_1_1/temp4[103] ,
         \MC_ARK_ARC_1_1/temp4[101] , \MC_ARK_ARC_1_1/temp4[100] ,
         \MC_ARK_ARC_1_1/temp4[99] , \MC_ARK_ARC_1_1/temp4[97] ,
         \MC_ARK_ARC_1_1/temp4[96] , \MC_ARK_ARC_1_1/temp4[95] ,
         \MC_ARK_ARC_1_1/temp4[94] , \MC_ARK_ARC_1_1/temp4[93] ,
         \MC_ARK_ARC_1_1/temp4[92] , \MC_ARK_ARC_1_1/temp4[91] ,
         \MC_ARK_ARC_1_1/temp4[90] , \MC_ARK_ARC_1_1/temp4[89] ,
         \MC_ARK_ARC_1_1/temp4[88] , \MC_ARK_ARC_1_1/temp4[87] ,
         \MC_ARK_ARC_1_1/temp4[86] , \MC_ARK_ARC_1_1/temp4[85] ,
         \MC_ARK_ARC_1_1/temp4[84] , \MC_ARK_ARC_1_1/temp4[82] ,
         \MC_ARK_ARC_1_1/temp4[81] , \MC_ARK_ARC_1_1/temp4[79] ,
         \MC_ARK_ARC_1_1/temp4[78] , \MC_ARK_ARC_1_1/temp4[77] ,
         \MC_ARK_ARC_1_1/temp4[76] , \MC_ARK_ARC_1_1/temp4[75] ,
         \MC_ARK_ARC_1_1/temp4[74] , \MC_ARK_ARC_1_1/temp4[73] ,
         \MC_ARK_ARC_1_1/temp4[72] , \MC_ARK_ARC_1_1/temp4[71] ,
         \MC_ARK_ARC_1_1/temp4[70] , \MC_ARK_ARC_1_1/temp4[69] ,
         \MC_ARK_ARC_1_1/temp4[68] , \MC_ARK_ARC_1_1/temp4[67] ,
         \MC_ARK_ARC_1_1/temp4[65] , \MC_ARK_ARC_1_1/temp4[64] ,
         \MC_ARK_ARC_1_1/temp4[63] , \MC_ARK_ARC_1_1/temp4[62] ,
         \MC_ARK_ARC_1_1/temp4[61] , \MC_ARK_ARC_1_1/temp4[60] ,
         \MC_ARK_ARC_1_1/temp4[59] , \MC_ARK_ARC_1_1/temp4[58] ,
         \MC_ARK_ARC_1_1/temp4[57] , \MC_ARK_ARC_1_1/temp4[55] ,
         \MC_ARK_ARC_1_1/temp4[54] , \MC_ARK_ARC_1_1/temp4[53] ,
         \MC_ARK_ARC_1_1/temp4[52] , \MC_ARK_ARC_1_1/temp4[51] ,
         \MC_ARK_ARC_1_1/temp4[50] , \MC_ARK_ARC_1_1/temp4[49] ,
         \MC_ARK_ARC_1_1/temp4[48] , \MC_ARK_ARC_1_1/temp4[46] ,
         \MC_ARK_ARC_1_1/temp4[45] , \MC_ARK_ARC_1_1/temp4[43] ,
         \MC_ARK_ARC_1_1/temp4[42] , \MC_ARK_ARC_1_1/temp4[40] ,
         \MC_ARK_ARC_1_1/temp4[39] , \MC_ARK_ARC_1_1/temp4[37] ,
         \MC_ARK_ARC_1_1/temp4[36] , \MC_ARK_ARC_1_1/temp4[34] ,
         \MC_ARK_ARC_1_1/temp4[33] , \MC_ARK_ARC_1_1/temp4[31] ,
         \MC_ARK_ARC_1_1/temp4[30] , \MC_ARK_ARC_1_1/temp4[29] ,
         \MC_ARK_ARC_1_1/temp4[28] , \MC_ARK_ARC_1_1/temp4[27] ,
         \MC_ARK_ARC_1_1/temp4[26] , \MC_ARK_ARC_1_1/temp4[25] ,
         \MC_ARK_ARC_1_1/temp4[24] , \MC_ARK_ARC_1_1/temp4[23] ,
         \MC_ARK_ARC_1_1/temp4[22] , \MC_ARK_ARC_1_1/temp4[21] ,
         \MC_ARK_ARC_1_1/temp4[20] , \MC_ARK_ARC_1_1/temp4[19] ,
         \MC_ARK_ARC_1_1/temp4[18] , \MC_ARK_ARC_1_1/temp4[17] ,
         \MC_ARK_ARC_1_1/temp4[16] , \MC_ARK_ARC_1_1/temp4[15] ,
         \MC_ARK_ARC_1_1/temp4[13] , \MC_ARK_ARC_1_1/temp4[12] ,
         \MC_ARK_ARC_1_1/temp4[11] , \MC_ARK_ARC_1_1/temp4[10] ,
         \MC_ARK_ARC_1_1/temp4[9] , \MC_ARK_ARC_1_1/temp4[8] ,
         \MC_ARK_ARC_1_1/temp4[7] , \MC_ARK_ARC_1_1/temp4[6] ,
         \MC_ARK_ARC_1_1/temp4[5] , \MC_ARK_ARC_1_1/temp4[4] ,
         \MC_ARK_ARC_1_1/temp4[3] , \MC_ARK_ARC_1_1/temp4[2] ,
         \MC_ARK_ARC_1_1/temp4[1] , \MC_ARK_ARC_1_1/temp4[0] ,
         \MC_ARK_ARC_1_1/temp3[191] , \MC_ARK_ARC_1_1/temp3[190] ,
         \MC_ARK_ARC_1_1/temp3[189] , \MC_ARK_ARC_1_1/temp3[187] ,
         \MC_ARK_ARC_1_1/temp3[186] , \MC_ARK_ARC_1_1/temp3[185] ,
         \MC_ARK_ARC_1_1/temp3[184] , \MC_ARK_ARC_1_1/temp3[183] ,
         \MC_ARK_ARC_1_1/temp3[182] , \MC_ARK_ARC_1_1/temp3[181] ,
         \MC_ARK_ARC_1_1/temp3[180] , \MC_ARK_ARC_1_1/temp3[178] ,
         \MC_ARK_ARC_1_1/temp3[177] , \MC_ARK_ARC_1_1/temp3[176] ,
         \MC_ARK_ARC_1_1/temp3[175] , \MC_ARK_ARC_1_1/temp3[174] ,
         \MC_ARK_ARC_1_1/temp3[170] , \MC_ARK_ARC_1_1/temp3[169] ,
         \MC_ARK_ARC_1_1/temp3[168] , \MC_ARK_ARC_1_1/temp3[166] ,
         \MC_ARK_ARC_1_1/temp3[164] , \MC_ARK_ARC_1_1/temp3[163] ,
         \MC_ARK_ARC_1_1/temp3[161] , \MC_ARK_ARC_1_1/temp3[160] ,
         \MC_ARK_ARC_1_1/temp3[157] , \MC_ARK_ARC_1_1/temp3[156] ,
         \MC_ARK_ARC_1_1/temp3[155] , \MC_ARK_ARC_1_1/temp3[154] ,
         \MC_ARK_ARC_1_1/temp3[153] , \MC_ARK_ARC_1_1/temp3[151] ,
         \MC_ARK_ARC_1_1/temp3[150] , \MC_ARK_ARC_1_1/temp3[149] ,
         \MC_ARK_ARC_1_1/temp3[148] , \MC_ARK_ARC_1_1/temp3[146] ,
         \MC_ARK_ARC_1_1/temp3[145] , \MC_ARK_ARC_1_1/temp3[143] ,
         \MC_ARK_ARC_1_1/temp3[142] , \MC_ARK_ARC_1_1/temp3[141] ,
         \MC_ARK_ARC_1_1/temp3[140] , \MC_ARK_ARC_1_1/temp3[139] ,
         \MC_ARK_ARC_1_1/temp3[138] , \MC_ARK_ARC_1_1/temp3[137] ,
         \MC_ARK_ARC_1_1/temp3[136] , \MC_ARK_ARC_1_1/temp3[133] ,
         \MC_ARK_ARC_1_1/temp3[132] , \MC_ARK_ARC_1_1/temp3[131] ,
         \MC_ARK_ARC_1_1/temp3[130] , \MC_ARK_ARC_1_1/temp3[129] ,
         \MC_ARK_ARC_1_1/temp3[128] , \MC_ARK_ARC_1_1/temp3[127] ,
         \MC_ARK_ARC_1_1/temp3[126] , \MC_ARK_ARC_1_1/temp3[125] ,
         \MC_ARK_ARC_1_1/temp3[124] , \MC_ARK_ARC_1_1/temp3[123] ,
         \MC_ARK_ARC_1_1/temp3[121] , \MC_ARK_ARC_1_1/temp3[119] ,
         \MC_ARK_ARC_1_1/temp3[118] , \MC_ARK_ARC_1_1/temp3[117] ,
         \MC_ARK_ARC_1_1/temp3[114] , \MC_ARK_ARC_1_1/temp3[112] ,
         \MC_ARK_ARC_1_1/temp3[111] , \MC_ARK_ARC_1_1/temp3[110] ,
         \MC_ARK_ARC_1_1/temp3[108] , \MC_ARK_ARC_1_1/temp3[106] ,
         \MC_ARK_ARC_1_1/temp3[105] , \MC_ARK_ARC_1_1/temp3[103] ,
         \MC_ARK_ARC_1_1/temp3[100] , \MC_ARK_ARC_1_1/temp3[97] ,
         \MC_ARK_ARC_1_1/temp3[96] , \MC_ARK_ARC_1_1/temp3[94] ,
         \MC_ARK_ARC_1_1/temp3[92] , \MC_ARK_ARC_1_1/temp3[91] ,
         \MC_ARK_ARC_1_1/temp3[90] , \MC_ARK_ARC_1_1/temp3[89] ,
         \MC_ARK_ARC_1_1/temp3[87] , \MC_ARK_ARC_1_1/temp3[86] ,
         \MC_ARK_ARC_1_1/temp3[84] , \MC_ARK_ARC_1_1/temp3[82] ,
         \MC_ARK_ARC_1_1/temp3[81] , \MC_ARK_ARC_1_1/temp3[78] ,
         \MC_ARK_ARC_1_1/temp3[77] , \MC_ARK_ARC_1_1/temp3[76] ,
         \MC_ARK_ARC_1_1/temp3[75] , \MC_ARK_ARC_1_1/temp3[74] ,
         \MC_ARK_ARC_1_1/temp3[72] , \MC_ARK_ARC_1_1/temp3[70] ,
         \MC_ARK_ARC_1_1/temp3[69] , \MC_ARK_ARC_1_1/temp3[68] ,
         \MC_ARK_ARC_1_1/temp3[67] , \MC_ARK_ARC_1_1/temp3[65] ,
         \MC_ARK_ARC_1_1/temp3[64] , \MC_ARK_ARC_1_1/temp3[63] ,
         \MC_ARK_ARC_1_1/temp3[62] , \MC_ARK_ARC_1_1/temp3[61] ,
         \MC_ARK_ARC_1_1/temp3[60] , \MC_ARK_ARC_1_1/temp3[58] ,
         \MC_ARK_ARC_1_1/temp3[55] , \MC_ARK_ARC_1_1/temp3[54] ,
         \MC_ARK_ARC_1_1/temp3[53] , \MC_ARK_ARC_1_1/temp3[52] ,
         \MC_ARK_ARC_1_1/temp3[50] , \MC_ARK_ARC_1_1/temp3[49] ,
         \MC_ARK_ARC_1_1/temp3[48] , \MC_ARK_ARC_1_1/temp3[46] ,
         \MC_ARK_ARC_1_1/temp3[45] , \MC_ARK_ARC_1_1/temp3[43] ,
         \MC_ARK_ARC_1_1/temp3[42] , \MC_ARK_ARC_1_1/temp3[40] ,
         \MC_ARK_ARC_1_1/temp3[39] , \MC_ARK_ARC_1_1/temp3[37] ,
         \MC_ARK_ARC_1_1/temp3[36] , \MC_ARK_ARC_1_1/temp3[34] ,
         \MC_ARK_ARC_1_1/temp3[33] , \MC_ARK_ARC_1_1/temp3[30] ,
         \MC_ARK_ARC_1_1/temp3[28] , \MC_ARK_ARC_1_1/temp3[27] ,
         \MC_ARK_ARC_1_1/temp3[25] , \MC_ARK_ARC_1_1/temp3[24] ,
         \MC_ARK_ARC_1_1/temp3[23] , \MC_ARK_ARC_1_1/temp3[22] ,
         \MC_ARK_ARC_1_1/temp3[21] , \MC_ARK_ARC_1_1/temp3[20] ,
         \MC_ARK_ARC_1_1/temp3[19] , \MC_ARK_ARC_1_1/temp3[18] ,
         \MC_ARK_ARC_1_1/temp3[16] , \MC_ARK_ARC_1_1/temp3[13] ,
         \MC_ARK_ARC_1_1/temp3[11] , \MC_ARK_ARC_1_1/temp3[10] ,
         \MC_ARK_ARC_1_1/temp3[9] , \MC_ARK_ARC_1_1/temp3[8] ,
         \MC_ARK_ARC_1_1/temp3[7] , \MC_ARK_ARC_1_1/temp3[6] ,
         \MC_ARK_ARC_1_1/temp3[5] , \MC_ARK_ARC_1_1/temp3[4] ,
         \MC_ARK_ARC_1_1/temp3[2] , \MC_ARK_ARC_1_1/temp3[1] ,
         \MC_ARK_ARC_1_1/temp3[0] , \MC_ARK_ARC_1_1/temp2[190] ,
         \MC_ARK_ARC_1_1/temp2[189] , \MC_ARK_ARC_1_1/temp2[187] ,
         \MC_ARK_ARC_1_1/temp2[186] , \MC_ARK_ARC_1_1/temp2[185] ,
         \MC_ARK_ARC_1_1/temp2[184] , \MC_ARK_ARC_1_1/temp2[181] ,
         \MC_ARK_ARC_1_1/temp2[180] , \MC_ARK_ARC_1_1/temp2[178] ,
         \MC_ARK_ARC_1_1/temp2[177] , \MC_ARK_ARC_1_1/temp2[175] ,
         \MC_ARK_ARC_1_1/temp2[174] , \MC_ARK_ARC_1_1/temp2[169] ,
         \MC_ARK_ARC_1_1/temp2[168] , \MC_ARK_ARC_1_1/temp2[166] ,
         \MC_ARK_ARC_1_1/temp2[165] , \MC_ARK_ARC_1_1/temp2[164] ,
         \MC_ARK_ARC_1_1/temp2[163] , \MC_ARK_ARC_1_1/temp2[162] ,
         \MC_ARK_ARC_1_1/temp2[161] , \MC_ARK_ARC_1_1/temp2[160] ,
         \MC_ARK_ARC_1_1/temp2[159] , \MC_ARK_ARC_1_1/temp2[156] ,
         \MC_ARK_ARC_1_1/temp2[154] , \MC_ARK_ARC_1_1/temp2[153] ,
         \MC_ARK_ARC_1_1/temp2[152] , \MC_ARK_ARC_1_1/temp2[151] ,
         \MC_ARK_ARC_1_1/temp2[150] , \MC_ARK_ARC_1_1/temp2[148] ,
         \MC_ARK_ARC_1_1/temp2[145] , \MC_ARK_ARC_1_1/temp2[144] ,
         \MC_ARK_ARC_1_1/temp2[143] , \MC_ARK_ARC_1_1/temp2[142] ,
         \MC_ARK_ARC_1_1/temp2[141] , \MC_ARK_ARC_1_1/temp2[140] ,
         \MC_ARK_ARC_1_1/temp2[139] , \MC_ARK_ARC_1_1/temp2[136] ,
         \MC_ARK_ARC_1_1/temp2[133] , \MC_ARK_ARC_1_1/temp2[132] ,
         \MC_ARK_ARC_1_1/temp2[130] , \MC_ARK_ARC_1_1/temp2[128] ,
         \MC_ARK_ARC_1_1/temp2[127] , \MC_ARK_ARC_1_1/temp2[126] ,
         \MC_ARK_ARC_1_1/temp2[125] , \MC_ARK_ARC_1_1/temp2[124] ,
         \MC_ARK_ARC_1_1/temp2[119] , \MC_ARK_ARC_1_1/temp2[118] ,
         \MC_ARK_ARC_1_1/temp2[117] , \MC_ARK_ARC_1_1/temp2[114] ,
         \MC_ARK_ARC_1_1/temp2[112] , \MC_ARK_ARC_1_1/temp2[110] ,
         \MC_ARK_ARC_1_1/temp2[108] , \MC_ARK_ARC_1_1/temp2[106] ,
         \MC_ARK_ARC_1_1/temp2[105] , \MC_ARK_ARC_1_1/temp2[103] ,
         \MC_ARK_ARC_1_1/temp2[102] , \MC_ARK_ARC_1_1/temp2[100] ,
         \MC_ARK_ARC_1_1/temp2[99] , \MC_ARK_ARC_1_1/temp2[98] ,
         \MC_ARK_ARC_1_1/temp2[97] , \MC_ARK_ARC_1_1/temp2[96] ,
         \MC_ARK_ARC_1_1/temp2[94] , \MC_ARK_ARC_1_1/temp2[93] ,
         \MC_ARK_ARC_1_1/temp2[91] , \MC_ARK_ARC_1_1/temp2[90] ,
         \MC_ARK_ARC_1_1/temp2[88] , \MC_ARK_ARC_1_1/temp2[85] ,
         \MC_ARK_ARC_1_1/temp2[84] , \MC_ARK_ARC_1_1/temp2[81] ,
         \MC_ARK_ARC_1_1/temp2[79] , \MC_ARK_ARC_1_1/temp2[78] ,
         \MC_ARK_ARC_1_1/temp2[76] , \MC_ARK_ARC_1_1/temp2[75] ,
         \MC_ARK_ARC_1_1/temp2[73] , \MC_ARK_ARC_1_1/temp2[72] ,
         \MC_ARK_ARC_1_1/temp2[71] , \MC_ARK_ARC_1_1/temp2[70] ,
         \MC_ARK_ARC_1_1/temp2[68] , \MC_ARK_ARC_1_1/temp2[67] ,
         \MC_ARK_ARC_1_1/temp2[66] , \MC_ARK_ARC_1_1/temp2[64] ,
         \MC_ARK_ARC_1_1/temp2[63] , \MC_ARK_ARC_1_1/temp2[61] ,
         \MC_ARK_ARC_1_1/temp2[58] , \MC_ARK_ARC_1_1/temp2[57] ,
         \MC_ARK_ARC_1_1/temp2[54] , \MC_ARK_ARC_1_1/temp2[53] ,
         \MC_ARK_ARC_1_1/temp2[52] , \MC_ARK_ARC_1_1/temp2[51] ,
         \MC_ARK_ARC_1_1/temp2[49] , \MC_ARK_ARC_1_1/temp2[48] ,
         \MC_ARK_ARC_1_1/temp2[47] , \MC_ARK_ARC_1_1/temp2[46] ,
         \MC_ARK_ARC_1_1/temp2[45] , \MC_ARK_ARC_1_1/temp2[43] ,
         \MC_ARK_ARC_1_1/temp2[41] , \MC_ARK_ARC_1_1/temp2[40] ,
         \MC_ARK_ARC_1_1/temp2[39] , \MC_ARK_ARC_1_1/temp2[38] ,
         \MC_ARK_ARC_1_1/temp2[37] , \MC_ARK_ARC_1_1/temp2[36] ,
         \MC_ARK_ARC_1_1/temp2[34] , \MC_ARK_ARC_1_1/temp2[33] ,
         \MC_ARK_ARC_1_1/temp2[32] , \MC_ARK_ARC_1_1/temp2[30] ,
         \MC_ARK_ARC_1_1/temp2[25] , \MC_ARK_ARC_1_1/temp2[24] ,
         \MC_ARK_ARC_1_1/temp2[22] , \MC_ARK_ARC_1_1/temp2[19] ,
         \MC_ARK_ARC_1_1/temp2[18] , \MC_ARK_ARC_1_1/temp2[17] ,
         \MC_ARK_ARC_1_1/temp2[16] , \MC_ARK_ARC_1_1/temp2[15] ,
         \MC_ARK_ARC_1_1/temp2[13] , \MC_ARK_ARC_1_1/temp2[12] ,
         \MC_ARK_ARC_1_1/temp2[11] , \MC_ARK_ARC_1_1/temp2[10] ,
         \MC_ARK_ARC_1_1/temp2[9] , \MC_ARK_ARC_1_1/temp2[6] ,
         \MC_ARK_ARC_1_1/temp2[5] , \MC_ARK_ARC_1_1/temp2[4] ,
         \MC_ARK_ARC_1_1/temp2[3] , \MC_ARK_ARC_1_1/temp2[2] ,
         \MC_ARK_ARC_1_1/temp2[1] , \MC_ARK_ARC_1_1/temp1[190] ,
         \MC_ARK_ARC_1_1/temp1[189] , \MC_ARK_ARC_1_1/temp1[188] ,
         \MC_ARK_ARC_1_1/temp1[187] , \MC_ARK_ARC_1_1/temp1[186] ,
         \MC_ARK_ARC_1_1/temp1[184] , \MC_ARK_ARC_1_1/temp1[183] ,
         \MC_ARK_ARC_1_1/temp1[181] , \MC_ARK_ARC_1_1/temp1[180] ,
         \MC_ARK_ARC_1_1/temp1[179] , \MC_ARK_ARC_1_1/temp1[178] ,
         \MC_ARK_ARC_1_1/temp1[174] , \MC_ARK_ARC_1_1/temp1[169] ,
         \MC_ARK_ARC_1_1/temp1[168] , \MC_ARK_ARC_1_1/temp1[164] ,
         \MC_ARK_ARC_1_1/temp1[163] , \MC_ARK_ARC_1_1/temp1[162] ,
         \MC_ARK_ARC_1_1/temp1[160] , \MC_ARK_ARC_1_1/temp1[159] ,
         \MC_ARK_ARC_1_1/temp1[157] , \MC_ARK_ARC_1_1/temp1[155] ,
         \MC_ARK_ARC_1_1/temp1[153] , \MC_ARK_ARC_1_1/temp1[152] ,
         \MC_ARK_ARC_1_1/temp1[151] , \MC_ARK_ARC_1_1/temp1[150] ,
         \MC_ARK_ARC_1_1/temp1[145] , \MC_ARK_ARC_1_1/temp1[142] ,
         \MC_ARK_ARC_1_1/temp1[140] , \MC_ARK_ARC_1_1/temp1[139] ,
         \MC_ARK_ARC_1_1/temp1[138] , \MC_ARK_ARC_1_1/temp1[136] ,
         \MC_ARK_ARC_1_1/temp1[133] , \MC_ARK_ARC_1_1/temp1[132] ,
         \MC_ARK_ARC_1_1/temp1[130] , \MC_ARK_ARC_1_1/temp1[127] ,
         \MC_ARK_ARC_1_1/temp1[126] , \MC_ARK_ARC_1_1/temp1[124] ,
         \MC_ARK_ARC_1_1/temp1[122] , \MC_ARK_ARC_1_1/temp1[118] ,
         \MC_ARK_ARC_1_1/temp1[117] , \MC_ARK_ARC_1_1/temp1[115] ,
         \MC_ARK_ARC_1_1/temp1[112] , \MC_ARK_ARC_1_1/temp1[111] ,
         \MC_ARK_ARC_1_1/temp1[110] , \MC_ARK_ARC_1_1/temp1[109] ,
         \MC_ARK_ARC_1_1/temp1[108] , \MC_ARK_ARC_1_1/temp1[106] ,
         \MC_ARK_ARC_1_1/temp1[105] , \MC_ARK_ARC_1_1/temp1[104] ,
         \MC_ARK_ARC_1_1/temp1[103] , \MC_ARK_ARC_1_1/temp1[102] ,
         \MC_ARK_ARC_1_1/temp1[100] , \MC_ARK_ARC_1_1/temp1[99] ,
         \MC_ARK_ARC_1_1/temp1[97] , \MC_ARK_ARC_1_1/temp1[96] ,
         \MC_ARK_ARC_1_1/temp1[94] , \MC_ARK_ARC_1_1/temp1[92] ,
         \MC_ARK_ARC_1_1/temp1[91] , \MC_ARK_ARC_1_1/temp1[90] ,
         \MC_ARK_ARC_1_1/temp1[89] , \MC_ARK_ARC_1_1/temp1[87] ,
         \MC_ARK_ARC_1_1/temp1[86] , \MC_ARK_ARC_1_1/temp1[85] ,
         \MC_ARK_ARC_1_1/temp1[84] , \MC_ARK_ARC_1_1/temp1[82] ,
         \MC_ARK_ARC_1_1/temp1[77] , \MC_ARK_ARC_1_1/temp1[76] ,
         \MC_ARK_ARC_1_1/temp1[75] , \MC_ARK_ARC_1_1/temp1[74] ,
         \MC_ARK_ARC_1_1/temp1[73] , \MC_ARK_ARC_1_1/temp1[72] ,
         \MC_ARK_ARC_1_1/temp1[71] , \MC_ARK_ARC_1_1/temp1[70] ,
         \MC_ARK_ARC_1_1/temp1[69] , \MC_ARK_ARC_1_1/temp1[67] ,
         \MC_ARK_ARC_1_1/temp1[66] , \MC_ARK_ARC_1_1/temp1[65] ,
         \MC_ARK_ARC_1_1/temp1[64] , \MC_ARK_ARC_1_1/temp1[61] ,
         \MC_ARK_ARC_1_1/temp1[55] , \MC_ARK_ARC_1_1/temp1[54] ,
         \MC_ARK_ARC_1_1/temp1[52] , \MC_ARK_ARC_1_1/temp1[51] ,
         \MC_ARK_ARC_1_1/temp1[50] , \MC_ARK_ARC_1_1/temp1[49] ,
         \MC_ARK_ARC_1_1/temp1[48] , \MC_ARK_ARC_1_1/temp1[46] ,
         \MC_ARK_ARC_1_1/temp1[44] , \MC_ARK_ARC_1_1/temp1[43] ,
         \MC_ARK_ARC_1_1/temp1[42] , \MC_ARK_ARC_1_1/temp1[40] ,
         \MC_ARK_ARC_1_1/temp1[37] , \MC_ARK_ARC_1_1/temp1[36] ,
         \MC_ARK_ARC_1_1/temp1[34] , \MC_ARK_ARC_1_1/temp1[31] ,
         \MC_ARK_ARC_1_1/temp1[30] , \MC_ARK_ARC_1_1/temp1[28] ,
         \MC_ARK_ARC_1_1/temp1[27] , \MC_ARK_ARC_1_1/temp1[25] ,
         \MC_ARK_ARC_1_1/temp1[24] , \MC_ARK_ARC_1_1/temp1[22] ,
         \MC_ARK_ARC_1_1/temp1[19] , \MC_ARK_ARC_1_1/temp1[18] ,
         \MC_ARK_ARC_1_1/temp1[17] , \MC_ARK_ARC_1_1/temp1[16] ,
         \MC_ARK_ARC_1_1/temp1[15] , \MC_ARK_ARC_1_1/temp1[14] ,
         \MC_ARK_ARC_1_1/temp1[13] , \MC_ARK_ARC_1_1/temp1[12] ,
         \MC_ARK_ARC_1_1/temp1[11] , \MC_ARK_ARC_1_1/temp1[10] ,
         \MC_ARK_ARC_1_1/temp1[8] , \MC_ARK_ARC_1_1/temp1[6] ,
         \MC_ARK_ARC_1_1/temp1[5] , \MC_ARK_ARC_1_1/temp1[3] ,
         \MC_ARK_ARC_1_1/temp1[2] , \MC_ARK_ARC_1_1/temp1[1] ,
         \MC_ARK_ARC_1_1/buf_keyinput[148] ,
         \MC_ARK_ARC_1_1/buf_keyinput[119] ,
         \MC_ARK_ARC_1_1/buf_keyinput[111] ,
         \MC_ARK_ARC_1_1/buf_datainput[189] ,
         \MC_ARK_ARC_1_1/buf_datainput[188] ,
         \MC_ARK_ARC_1_1/buf_datainput[187] ,
         \MC_ARK_ARC_1_1/buf_datainput[182] ,
         \MC_ARK_ARC_1_1/buf_datainput[178] ,
         \MC_ARK_ARC_1_1/buf_datainput[177] ,
         \MC_ARK_ARC_1_1/buf_datainput[172] ,
         \MC_ARK_ARC_1_1/buf_datainput[168] ,
         \MC_ARK_ARC_1_1/buf_datainput[164] ,
         \MC_ARK_ARC_1_1/buf_datainput[163] ,
         \MC_ARK_ARC_1_1/buf_datainput[162] ,
         \MC_ARK_ARC_1_1/buf_datainput[152] ,
         \MC_ARK_ARC_1_1/buf_datainput[151] ,
         \MC_ARK_ARC_1_1/buf_datainput[150] ,
         \MC_ARK_ARC_1_1/buf_datainput[146] ,
         \MC_ARK_ARC_1_1/buf_datainput[145] ,
         \MC_ARK_ARC_1_1/buf_datainput[141] ,
         \MC_ARK_ARC_1_1/buf_datainput[125] ,
         \MC_ARK_ARC_1_1/buf_datainput[124] ,
         \MC_ARK_ARC_1_1/buf_datainput[122] ,
         \MC_ARK_ARC_1_1/buf_datainput[117] ,
         \MC_ARK_ARC_1_1/buf_datainput[110] ,
         \MC_ARK_ARC_1_1/buf_datainput[108] ,
         \MC_ARK_ARC_1_1/buf_datainput[103] ,
         \MC_ARK_ARC_1_1/buf_datainput[94] ,
         \MC_ARK_ARC_1_1/buf_datainput[84] ,
         \MC_ARK_ARC_1_1/buf_datainput[83] ,
         \MC_ARK_ARC_1_1/buf_datainput[76] ,
         \MC_ARK_ARC_1_1/buf_datainput[73] ,
         \MC_ARK_ARC_1_1/buf_datainput[72] ,
         \MC_ARK_ARC_1_1/buf_datainput[71] ,
         \MC_ARK_ARC_1_1/buf_datainput[62] ,
         \MC_ARK_ARC_1_1/buf_datainput[58] ,
         \MC_ARK_ARC_1_1/buf_datainput[50] ,
         \MC_ARK_ARC_1_1/buf_datainput[48] ,
         \MC_ARK_ARC_1_1/buf_datainput[45] ,
         \MC_ARK_ARC_1_1/buf_datainput[44] ,
         \MC_ARK_ARC_1_1/buf_datainput[38] ,
         \MC_ARK_ARC_1_1/buf_datainput[37] ,
         \MC_ARK_ARC_1_1/buf_datainput[36] ,
         \MC_ARK_ARC_1_1/buf_datainput[34] ,
         \MC_ARK_ARC_1_1/buf_datainput[32] ,
         \MC_ARK_ARC_1_1/buf_datainput[22] ,
         \MC_ARK_ARC_1_1/buf_datainput[21] ,
         \MC_ARK_ARC_1_1/buf_datainput[15] , \MC_ARK_ARC_1_1/buf_datainput[7] ,
         \MC_ARK_ARC_1_1/buf_datainput[4] , \MC_ARK_ARC_1_1/buf_datainput[3] ,
         \MC_ARK_ARC_1_1/buf_datainput[1] , \MC_ARK_ARC_1_1/buf_datainput[0] ,
         \MC_ARK_ARC_1_2/buf_output[190] , \MC_ARK_ARC_1_2/buf_output[189] ,
         \MC_ARK_ARC_1_2/buf_output[188] , \MC_ARK_ARC_1_2/buf_output[187] ,
         \MC_ARK_ARC_1_2/buf_output[186] , \MC_ARK_ARC_1_2/buf_output[185] ,
         \MC_ARK_ARC_1_2/buf_output[184] , \MC_ARK_ARC_1_2/buf_output[183] ,
         \MC_ARK_ARC_1_2/buf_output[182] , \MC_ARK_ARC_1_2/buf_output[181] ,
         \MC_ARK_ARC_1_2/buf_output[180] , \MC_ARK_ARC_1_2/buf_output[179] ,
         \MC_ARK_ARC_1_2/buf_output[178] , \MC_ARK_ARC_1_2/buf_output[177] ,
         \MC_ARK_ARC_1_2/buf_output[176] , \MC_ARK_ARC_1_2/buf_output[175] ,
         \MC_ARK_ARC_1_2/buf_output[174] , \MC_ARK_ARC_1_2/buf_output[173] ,
         \MC_ARK_ARC_1_2/buf_output[172] , \MC_ARK_ARC_1_2/buf_output[171] ,
         \MC_ARK_ARC_1_2/buf_output[170] , \MC_ARK_ARC_1_2/buf_output[169] ,
         \MC_ARK_ARC_1_2/buf_output[168] , \MC_ARK_ARC_1_2/buf_output[167] ,
         \MC_ARK_ARC_1_2/buf_output[166] , \MC_ARK_ARC_1_2/buf_output[164] ,
         \MC_ARK_ARC_1_2/buf_output[163] , \MC_ARK_ARC_1_2/buf_output[162] ,
         \MC_ARK_ARC_1_2/buf_output[160] , \MC_ARK_ARC_1_2/buf_output[159] ,
         \MC_ARK_ARC_1_2/buf_output[158] , \MC_ARK_ARC_1_2/buf_output[157] ,
         \MC_ARK_ARC_1_2/buf_output[156] , \MC_ARK_ARC_1_2/buf_output[155] ,
         \MC_ARK_ARC_1_2/buf_output[154] , \MC_ARK_ARC_1_2/buf_output[153] ,
         \MC_ARK_ARC_1_2/buf_output[152] , \MC_ARK_ARC_1_2/buf_output[151] ,
         \MC_ARK_ARC_1_2/buf_output[150] , \MC_ARK_ARC_1_2/buf_output[149] ,
         \MC_ARK_ARC_1_2/buf_output[148] , \MC_ARK_ARC_1_2/buf_output[147] ,
         \MC_ARK_ARC_1_2/buf_output[146] , \MC_ARK_ARC_1_2/buf_output[145] ,
         \MC_ARK_ARC_1_2/buf_output[144] , \MC_ARK_ARC_1_2/buf_output[143] ,
         \MC_ARK_ARC_1_2/buf_output[142] , \MC_ARK_ARC_1_2/buf_output[141] ,
         \MC_ARK_ARC_1_2/buf_output[140] , \MC_ARK_ARC_1_2/buf_output[139] ,
         \MC_ARK_ARC_1_2/buf_output[138] , \MC_ARK_ARC_1_2/buf_output[137] ,
         \MC_ARK_ARC_1_2/buf_output[136] , \MC_ARK_ARC_1_2/buf_output[135] ,
         \MC_ARK_ARC_1_2/buf_output[134] , \MC_ARK_ARC_1_2/buf_output[133] ,
         \MC_ARK_ARC_1_2/buf_output[132] , \MC_ARK_ARC_1_2/buf_output[131] ,
         \MC_ARK_ARC_1_2/buf_output[130] , \MC_ARK_ARC_1_2/buf_output[129] ,
         \MC_ARK_ARC_1_2/buf_output[128] , \MC_ARK_ARC_1_2/buf_output[127] ,
         \MC_ARK_ARC_1_2/buf_output[126] , \MC_ARK_ARC_1_2/buf_output[125] ,
         \MC_ARK_ARC_1_2/buf_output[124] , \MC_ARK_ARC_1_2/buf_output[123] ,
         \MC_ARK_ARC_1_2/buf_output[122] , \MC_ARK_ARC_1_2/buf_output[121] ,
         \MC_ARK_ARC_1_2/buf_output[120] , \MC_ARK_ARC_1_2/buf_output[119] ,
         \MC_ARK_ARC_1_2/buf_output[118] , \MC_ARK_ARC_1_2/buf_output[117] ,
         \MC_ARK_ARC_1_2/buf_output[116] , \MC_ARK_ARC_1_2/buf_output[115] ,
         \MC_ARK_ARC_1_2/buf_output[114] , \MC_ARK_ARC_1_2/buf_output[113] ,
         \MC_ARK_ARC_1_2/buf_output[112] , \MC_ARK_ARC_1_2/buf_output[111] ,
         \MC_ARK_ARC_1_2/buf_output[110] , \MC_ARK_ARC_1_2/buf_output[109] ,
         \MC_ARK_ARC_1_2/buf_output[108] , \MC_ARK_ARC_1_2/buf_output[107] ,
         \MC_ARK_ARC_1_2/buf_output[106] , \MC_ARK_ARC_1_2/buf_output[105] ,
         \MC_ARK_ARC_1_2/buf_output[104] , \MC_ARK_ARC_1_2/buf_output[103] ,
         \MC_ARK_ARC_1_2/buf_output[102] , \MC_ARK_ARC_1_2/buf_output[100] ,
         \MC_ARK_ARC_1_2/buf_output[99] , \MC_ARK_ARC_1_2/buf_output[98] ,
         \MC_ARK_ARC_1_2/buf_output[97] , \MC_ARK_ARC_1_2/buf_output[96] ,
         \MC_ARK_ARC_1_2/buf_output[95] , \MC_ARK_ARC_1_2/buf_output[94] ,
         \MC_ARK_ARC_1_2/buf_output[93] , \MC_ARK_ARC_1_2/buf_output[92] ,
         \MC_ARK_ARC_1_2/buf_output[91] , \MC_ARK_ARC_1_2/buf_output[90] ,
         \MC_ARK_ARC_1_2/buf_output[89] , \MC_ARK_ARC_1_2/buf_output[88] ,
         \MC_ARK_ARC_1_2/buf_output[87] , \MC_ARK_ARC_1_2/buf_output[86] ,
         \MC_ARK_ARC_1_2/buf_output[85] , \MC_ARK_ARC_1_2/buf_output[84] ,
         \MC_ARK_ARC_1_2/buf_output[83] , \MC_ARK_ARC_1_2/buf_output[82] ,
         \MC_ARK_ARC_1_2/buf_output[81] , \MC_ARK_ARC_1_2/buf_output[80] ,
         \MC_ARK_ARC_1_2/buf_output[79] , \MC_ARK_ARC_1_2/buf_output[78] ,
         \MC_ARK_ARC_1_2/buf_output[77] , \MC_ARK_ARC_1_2/buf_output[76] ,
         \MC_ARK_ARC_1_2/buf_output[75] , \MC_ARK_ARC_1_2/buf_output[74] ,
         \MC_ARK_ARC_1_2/buf_output[73] , \MC_ARK_ARC_1_2/buf_output[72] ,
         \MC_ARK_ARC_1_2/buf_output[71] , \MC_ARK_ARC_1_2/buf_output[70] ,
         \MC_ARK_ARC_1_2/buf_output[69] , \MC_ARK_ARC_1_2/buf_output[68] ,
         \MC_ARK_ARC_1_2/buf_output[67] , \MC_ARK_ARC_1_2/buf_output[66] ,
         \MC_ARK_ARC_1_2/buf_output[64] , \MC_ARK_ARC_1_2/buf_output[63] ,
         \MC_ARK_ARC_1_2/buf_output[62] , \MC_ARK_ARC_1_2/buf_output[61] ,
         \MC_ARK_ARC_1_2/buf_output[60] , \MC_ARK_ARC_1_2/buf_output[59] ,
         \MC_ARK_ARC_1_2/buf_output[58] , \MC_ARK_ARC_1_2/buf_output[57] ,
         \MC_ARK_ARC_1_2/buf_output[56] , \MC_ARK_ARC_1_2/buf_output[55] ,
         \MC_ARK_ARC_1_2/buf_output[54] , \MC_ARK_ARC_1_2/buf_output[53] ,
         \MC_ARK_ARC_1_2/buf_output[52] , \MC_ARK_ARC_1_2/buf_output[51] ,
         \MC_ARK_ARC_1_2/buf_output[50] , \MC_ARK_ARC_1_2/buf_output[49] ,
         \MC_ARK_ARC_1_2/buf_output[48] , \MC_ARK_ARC_1_2/buf_output[47] ,
         \MC_ARK_ARC_1_2/buf_output[46] , \MC_ARK_ARC_1_2/buf_output[45] ,
         \MC_ARK_ARC_1_2/buf_output[44] , \MC_ARK_ARC_1_2/buf_output[43] ,
         \MC_ARK_ARC_1_2/buf_output[42] , \MC_ARK_ARC_1_2/buf_output[41] ,
         \MC_ARK_ARC_1_2/buf_output[40] , \MC_ARK_ARC_1_2/buf_output[39] ,
         \MC_ARK_ARC_1_2/buf_output[38] , \MC_ARK_ARC_1_2/buf_output[37] ,
         \MC_ARK_ARC_1_2/buf_output[36] , \MC_ARK_ARC_1_2/buf_output[35] ,
         \MC_ARK_ARC_1_2/buf_output[34] , \MC_ARK_ARC_1_2/buf_output[33] ,
         \MC_ARK_ARC_1_2/buf_output[32] , \MC_ARK_ARC_1_2/buf_output[31] ,
         \MC_ARK_ARC_1_2/buf_output[30] , \MC_ARK_ARC_1_2/buf_output[29] ,
         \MC_ARK_ARC_1_2/buf_output[27] , \MC_ARK_ARC_1_2/buf_output[26] ,
         \MC_ARK_ARC_1_2/buf_output[25] , \MC_ARK_ARC_1_2/buf_output[24] ,
         \MC_ARK_ARC_1_2/buf_output[23] , \MC_ARK_ARC_1_2/buf_output[22] ,
         \MC_ARK_ARC_1_2/buf_output[21] , \MC_ARK_ARC_1_2/buf_output[20] ,
         \MC_ARK_ARC_1_2/buf_output[19] , \MC_ARK_ARC_1_2/buf_output[18] ,
         \MC_ARK_ARC_1_2/buf_output[16] , \MC_ARK_ARC_1_2/buf_output[15] ,
         \MC_ARK_ARC_1_2/buf_output[14] , \MC_ARK_ARC_1_2/buf_output[13] ,
         \MC_ARK_ARC_1_2/buf_output[12] , \MC_ARK_ARC_1_2/buf_output[11] ,
         \MC_ARK_ARC_1_2/buf_output[10] , \MC_ARK_ARC_1_2/buf_output[9] ,
         \MC_ARK_ARC_1_2/buf_output[8] , \MC_ARK_ARC_1_2/buf_output[7] ,
         \MC_ARK_ARC_1_2/buf_output[6] , \MC_ARK_ARC_1_2/buf_output[4] ,
         \MC_ARK_ARC_1_2/buf_output[3] , \MC_ARK_ARC_1_2/buf_output[2] ,
         \MC_ARK_ARC_1_2/buf_output[1] , \MC_ARK_ARC_1_2/buf_output[0] ,
         \MC_ARK_ARC_1_2/temp6[188] , \MC_ARK_ARC_1_2/temp6[185] ,
         \MC_ARK_ARC_1_2/temp6[184] , \MC_ARK_ARC_1_2/temp6[180] ,
         \MC_ARK_ARC_1_2/temp6[176] , \MC_ARK_ARC_1_2/temp6[174] ,
         \MC_ARK_ARC_1_2/temp6[173] , \MC_ARK_ARC_1_2/temp6[172] ,
         \MC_ARK_ARC_1_2/temp6[171] , \MC_ARK_ARC_1_2/temp6[170] ,
         \MC_ARK_ARC_1_2/temp6[169] , \MC_ARK_ARC_1_2/temp6[168] ,
         \MC_ARK_ARC_1_2/temp6[167] , \MC_ARK_ARC_1_2/temp6[166] ,
         \MC_ARK_ARC_1_2/temp6[165] , \MC_ARK_ARC_1_2/temp6[162] ,
         \MC_ARK_ARC_1_2/temp6[160] , \MC_ARK_ARC_1_2/temp6[159] ,
         \MC_ARK_ARC_1_2/temp6[156] , \MC_ARK_ARC_1_2/temp6[153] ,
         \MC_ARK_ARC_1_2/temp6[151] , \MC_ARK_ARC_1_2/temp6[150] ,
         \MC_ARK_ARC_1_2/temp6[148] , \MC_ARK_ARC_1_2/temp6[147] ,
         \MC_ARK_ARC_1_2/temp6[146] , \MC_ARK_ARC_1_2/temp6[144] ,
         \MC_ARK_ARC_1_2/temp6[143] , \MC_ARK_ARC_1_2/temp6[141] ,
         \MC_ARK_ARC_1_2/temp6[140] , \MC_ARK_ARC_1_2/temp6[139] ,
         \MC_ARK_ARC_1_2/temp6[138] , \MC_ARK_ARC_1_2/temp6[134] ,
         \MC_ARK_ARC_1_2/temp6[133] , \MC_ARK_ARC_1_2/temp6[132] ,
         \MC_ARK_ARC_1_2/temp6[131] , \MC_ARK_ARC_1_2/temp6[130] ,
         \MC_ARK_ARC_1_2/temp6[128] , \MC_ARK_ARC_1_2/temp6[127] ,
         \MC_ARK_ARC_1_2/temp6[126] , \MC_ARK_ARC_1_2/temp6[125] ,
         \MC_ARK_ARC_1_2/temp6[122] , \MC_ARK_ARC_1_2/temp6[121] ,
         \MC_ARK_ARC_1_2/temp6[120] , \MC_ARK_ARC_1_2/temp6[114] ,
         \MC_ARK_ARC_1_2/temp6[112] , \MC_ARK_ARC_1_2/temp6[110] ,
         \MC_ARK_ARC_1_2/temp6[109] , \MC_ARK_ARC_1_2/temp6[106] ,
         \MC_ARK_ARC_1_2/temp6[103] , \MC_ARK_ARC_1_2/temp6[95] ,
         \MC_ARK_ARC_1_2/temp6[94] , \MC_ARK_ARC_1_2/temp6[92] ,
         \MC_ARK_ARC_1_2/temp6[91] , \MC_ARK_ARC_1_2/temp6[90] ,
         \MC_ARK_ARC_1_2/temp6[84] , \MC_ARK_ARC_1_2/temp6[83] ,
         \MC_ARK_ARC_1_2/temp6[82] , \MC_ARK_ARC_1_2/temp6[80] ,
         \MC_ARK_ARC_1_2/temp6[79] , \MC_ARK_ARC_1_2/temp6[76] ,
         \MC_ARK_ARC_1_2/temp6[72] , \MC_ARK_ARC_1_2/temp6[70] ,
         \MC_ARK_ARC_1_2/temp6[65] , \MC_ARK_ARC_1_2/temp6[63] ,
         \MC_ARK_ARC_1_2/temp6[62] , \MC_ARK_ARC_1_2/temp6[61] ,
         \MC_ARK_ARC_1_2/temp6[52] , \MC_ARK_ARC_1_2/temp6[51] ,
         \MC_ARK_ARC_1_2/temp6[48] , \MC_ARK_ARC_1_2/temp6[46] ,
         \MC_ARK_ARC_1_2/temp6[42] , \MC_ARK_ARC_1_2/temp6[37] ,
         \MC_ARK_ARC_1_2/temp6[34] , \MC_ARK_ARC_1_2/temp6[33] ,
         \MC_ARK_ARC_1_2/temp6[31] , \MC_ARK_ARC_1_2/temp6[30] ,
         \MC_ARK_ARC_1_2/temp6[28] , \MC_ARK_ARC_1_2/temp6[27] ,
         \MC_ARK_ARC_1_2/temp6[25] , \MC_ARK_ARC_1_2/temp6[18] ,
         \MC_ARK_ARC_1_2/temp6[13] , \MC_ARK_ARC_1_2/temp6[11] ,
         \MC_ARK_ARC_1_2/temp6[5] , \MC_ARK_ARC_1_2/temp6[4] ,
         \MC_ARK_ARC_1_2/temp6[3] , \MC_ARK_ARC_1_2/temp5[191] ,
         \MC_ARK_ARC_1_2/temp5[190] , \MC_ARK_ARC_1_2/temp5[189] ,
         \MC_ARK_ARC_1_2/temp5[188] , \MC_ARK_ARC_1_2/temp5[187] ,
         \MC_ARK_ARC_1_2/temp5[184] , \MC_ARK_ARC_1_2/temp5[183] ,
         \MC_ARK_ARC_1_2/temp5[181] , \MC_ARK_ARC_1_2/temp5[177] ,
         \MC_ARK_ARC_1_2/temp5[176] , \MC_ARK_ARC_1_2/temp5[172] ,
         \MC_ARK_ARC_1_2/temp5[171] , \MC_ARK_ARC_1_2/temp5[170] ,
         \MC_ARK_ARC_1_2/temp5[165] , \MC_ARK_ARC_1_2/temp5[161] ,
         \MC_ARK_ARC_1_2/temp5[160] , \MC_ARK_ARC_1_2/temp5[159] ,
         \MC_ARK_ARC_1_2/temp5[157] , \MC_ARK_ARC_1_2/temp5[156] ,
         \MC_ARK_ARC_1_2/temp5[154] , \MC_ARK_ARC_1_2/temp5[151] ,
         \MC_ARK_ARC_1_2/temp5[150] , \MC_ARK_ARC_1_2/temp5[149] ,
         \MC_ARK_ARC_1_2/temp5[148] , \MC_ARK_ARC_1_2/temp5[147] ,
         \MC_ARK_ARC_1_2/temp5[144] , \MC_ARK_ARC_1_2/temp5[143] ,
         \MC_ARK_ARC_1_2/temp5[142] , \MC_ARK_ARC_1_2/temp5[141] ,
         \MC_ARK_ARC_1_2/temp5[140] , \MC_ARK_ARC_1_2/temp5[139] ,
         \MC_ARK_ARC_1_2/temp5[138] , \MC_ARK_ARC_1_2/temp5[135] ,
         \MC_ARK_ARC_1_2/temp5[134] , \MC_ARK_ARC_1_2/temp5[132] ,
         \MC_ARK_ARC_1_2/temp5[131] , \MC_ARK_ARC_1_2/temp5[130] ,
         \MC_ARK_ARC_1_2/temp5[129] , \MC_ARK_ARC_1_2/temp5[124] ,
         \MC_ARK_ARC_1_2/temp5[122] , \MC_ARK_ARC_1_2/temp5[120] ,
         \MC_ARK_ARC_1_2/temp5[118] , \MC_ARK_ARC_1_2/temp5[112] ,
         \MC_ARK_ARC_1_2/temp5[110] , \MC_ARK_ARC_1_2/temp5[108] ,
         \MC_ARK_ARC_1_2/temp5[102] , \MC_ARK_ARC_1_2/temp5[101] ,
         \MC_ARK_ARC_1_2/temp5[100] , \MC_ARK_ARC_1_2/temp5[99] ,
         \MC_ARK_ARC_1_2/temp5[97] , \MC_ARK_ARC_1_2/temp5[95] ,
         \MC_ARK_ARC_1_2/temp5[91] , \MC_ARK_ARC_1_2/temp5[90] ,
         \MC_ARK_ARC_1_2/temp5[86] , \MC_ARK_ARC_1_2/temp5[85] ,
         \MC_ARK_ARC_1_2/temp5[84] , \MC_ARK_ARC_1_2/temp5[83] ,
         \MC_ARK_ARC_1_2/temp5[82] , \MC_ARK_ARC_1_2/temp5[81] ,
         \MC_ARK_ARC_1_2/temp5[80] , \MC_ARK_ARC_1_2/temp5[79] ,
         \MC_ARK_ARC_1_2/temp5[77] , \MC_ARK_ARC_1_2/temp5[76] ,
         \MC_ARK_ARC_1_2/temp5[75] , \MC_ARK_ARC_1_2/temp5[74] ,
         \MC_ARK_ARC_1_2/temp5[73] , \MC_ARK_ARC_1_2/temp5[72] ,
         \MC_ARK_ARC_1_2/temp5[71] , \MC_ARK_ARC_1_2/temp5[69] ,
         \MC_ARK_ARC_1_2/temp5[68] , \MC_ARK_ARC_1_2/temp5[67] ,
         \MC_ARK_ARC_1_2/temp5[66] , \MC_ARK_ARC_1_2/temp5[64] ,
         \MC_ARK_ARC_1_2/temp5[61] , \MC_ARK_ARC_1_2/temp5[58] ,
         \MC_ARK_ARC_1_2/temp5[54] , \MC_ARK_ARC_1_2/temp5[53] ,
         \MC_ARK_ARC_1_2/temp5[52] , \MC_ARK_ARC_1_2/temp5[49] ,
         \MC_ARK_ARC_1_2/temp5[48] , \MC_ARK_ARC_1_2/temp5[47] ,
         \MC_ARK_ARC_1_2/temp5[45] , \MC_ARK_ARC_1_2/temp5[44] ,
         \MC_ARK_ARC_1_2/temp5[43] , \MC_ARK_ARC_1_2/temp5[42] ,
         \MC_ARK_ARC_1_2/temp5[37] , \MC_ARK_ARC_1_2/temp5[36] ,
         \MC_ARK_ARC_1_2/temp5[35] , \MC_ARK_ARC_1_2/temp5[34] ,
         \MC_ARK_ARC_1_2/temp5[31] , \MC_ARK_ARC_1_2/temp5[30] ,
         \MC_ARK_ARC_1_2/temp5[28] , \MC_ARK_ARC_1_2/temp5[27] ,
         \MC_ARK_ARC_1_2/temp5[25] , \MC_ARK_ARC_1_2/temp5[20] ,
         \MC_ARK_ARC_1_2/temp5[19] , \MC_ARK_ARC_1_2/temp5[17] ,
         \MC_ARK_ARC_1_2/temp5[16] , \MC_ARK_ARC_1_2/temp5[15] ,
         \MC_ARK_ARC_1_2/temp5[12] , \MC_ARK_ARC_1_2/temp5[10] ,
         \MC_ARK_ARC_1_2/temp5[8] , \MC_ARK_ARC_1_2/temp5[6] ,
         \MC_ARK_ARC_1_2/temp5[5] , \MC_ARK_ARC_1_2/temp5[4] ,
         \MC_ARK_ARC_1_2/temp5[3] , \MC_ARK_ARC_1_2/temp5[2] ,
         \MC_ARK_ARC_1_2/temp4[191] , \MC_ARK_ARC_1_2/temp4[190] ,
         \MC_ARK_ARC_1_2/temp4[189] , \MC_ARK_ARC_1_2/temp4[188] ,
         \MC_ARK_ARC_1_2/temp4[187] , \MC_ARK_ARC_1_2/temp4[186] ,
         \MC_ARK_ARC_1_2/temp4[185] , \MC_ARK_ARC_1_2/temp4[184] ,
         \MC_ARK_ARC_1_2/temp4[183] , \MC_ARK_ARC_1_2/temp4[182] ,
         \MC_ARK_ARC_1_2/temp4[181] , \MC_ARK_ARC_1_2/temp4[180] ,
         \MC_ARK_ARC_1_2/temp4[178] , \MC_ARK_ARC_1_2/temp4[177] ,
         \MC_ARK_ARC_1_2/temp4[175] , \MC_ARK_ARC_1_2/temp4[174] ,
         \MC_ARK_ARC_1_2/temp4[173] , \MC_ARK_ARC_1_2/temp4[172] ,
         \MC_ARK_ARC_1_2/temp4[171] , \MC_ARK_ARC_1_2/temp4[169] ,
         \MC_ARK_ARC_1_2/temp4[168] , \MC_ARK_ARC_1_2/temp4[167] ,
         \MC_ARK_ARC_1_2/temp4[166] , \MC_ARK_ARC_1_2/temp4[165] ,
         \MC_ARK_ARC_1_2/temp4[164] , \MC_ARK_ARC_1_2/temp4[163] ,
         \MC_ARK_ARC_1_2/temp4[162] , \MC_ARK_ARC_1_2/temp4[161] ,
         \MC_ARK_ARC_1_2/temp4[160] , \MC_ARK_ARC_1_2/temp4[159] ,
         \MC_ARK_ARC_1_2/temp4[158] , \MC_ARK_ARC_1_2/temp4[157] ,
         \MC_ARK_ARC_1_2/temp4[156] , \MC_ARK_ARC_1_2/temp4[154] ,
         \MC_ARK_ARC_1_2/temp4[152] , \MC_ARK_ARC_1_2/temp4[151] ,
         \MC_ARK_ARC_1_2/temp4[150] , \MC_ARK_ARC_1_2/temp4[149] ,
         \MC_ARK_ARC_1_2/temp4[148] , \MC_ARK_ARC_1_2/temp4[147] ,
         \MC_ARK_ARC_1_2/temp4[146] , \MC_ARK_ARC_1_2/temp4[145] ,
         \MC_ARK_ARC_1_2/temp4[144] , \MC_ARK_ARC_1_2/temp4[142] ,
         \MC_ARK_ARC_1_2/temp4[141] , \MC_ARK_ARC_1_2/temp4[140] ,
         \MC_ARK_ARC_1_2/temp4[138] , \MC_ARK_ARC_1_2/temp4[137] ,
         \MC_ARK_ARC_1_2/temp4[136] , \MC_ARK_ARC_1_2/temp4[135] ,
         \MC_ARK_ARC_1_2/temp4[134] , \MC_ARK_ARC_1_2/temp4[133] ,
         \MC_ARK_ARC_1_2/temp4[132] , \MC_ARK_ARC_1_2/temp4[131] ,
         \MC_ARK_ARC_1_2/temp4[130] , \MC_ARK_ARC_1_2/temp4[129] ,
         \MC_ARK_ARC_1_2/temp4[128] , \MC_ARK_ARC_1_2/temp4[127] ,
         \MC_ARK_ARC_1_2/temp4[126] , \MC_ARK_ARC_1_2/temp4[125] ,
         \MC_ARK_ARC_1_2/temp4[124] , \MC_ARK_ARC_1_2/temp4[123] ,
         \MC_ARK_ARC_1_2/temp4[122] , \MC_ARK_ARC_1_2/temp4[121] ,
         \MC_ARK_ARC_1_2/temp4[119] , \MC_ARK_ARC_1_2/temp4[118] ,
         \MC_ARK_ARC_1_2/temp4[117] , \MC_ARK_ARC_1_2/temp4[116] ,
         \MC_ARK_ARC_1_2/temp4[115] , \MC_ARK_ARC_1_2/temp4[114] ,
         \MC_ARK_ARC_1_2/temp4[113] , \MC_ARK_ARC_1_2/temp4[112] ,
         \MC_ARK_ARC_1_2/temp4[111] , \MC_ARK_ARC_1_2/temp4[109] ,
         \MC_ARK_ARC_1_2/temp4[108] , \MC_ARK_ARC_1_2/temp4[107] ,
         \MC_ARK_ARC_1_2/temp4[106] , \MC_ARK_ARC_1_2/temp4[105] ,
         \MC_ARK_ARC_1_2/temp4[104] , \MC_ARK_ARC_1_2/temp4[103] ,
         \MC_ARK_ARC_1_2/temp4[102] , \MC_ARK_ARC_1_2/temp4[101] ,
         \MC_ARK_ARC_1_2/temp4[100] , \MC_ARK_ARC_1_2/temp4[99] ,
         \MC_ARK_ARC_1_2/temp4[97] , \MC_ARK_ARC_1_2/temp4[96] ,
         \MC_ARK_ARC_1_2/temp4[95] , \MC_ARK_ARC_1_2/temp4[94] ,
         \MC_ARK_ARC_1_2/temp4[93] , \MC_ARK_ARC_1_2/temp4[91] ,
         \MC_ARK_ARC_1_2/temp4[90] , \MC_ARK_ARC_1_2/temp4[89] ,
         \MC_ARK_ARC_1_2/temp4[88] , \MC_ARK_ARC_1_2/temp4[87] ,
         \MC_ARK_ARC_1_2/temp4[86] , \MC_ARK_ARC_1_2/temp4[85] ,
         \MC_ARK_ARC_1_2/temp4[84] , \MC_ARK_ARC_1_2/temp4[83] ,
         \MC_ARK_ARC_1_2/temp4[82] , \MC_ARK_ARC_1_2/temp4[80] ,
         \MC_ARK_ARC_1_2/temp4[79] , \MC_ARK_ARC_1_2/temp4[78] ,
         \MC_ARK_ARC_1_2/temp4[77] , \MC_ARK_ARC_1_2/temp4[76] ,
         \MC_ARK_ARC_1_2/temp4[75] , \MC_ARK_ARC_1_2/temp4[73] ,
         \MC_ARK_ARC_1_2/temp4[72] , \MC_ARK_ARC_1_2/temp4[71] ,
         \MC_ARK_ARC_1_2/temp4[70] , \MC_ARK_ARC_1_2/temp4[69] ,
         \MC_ARK_ARC_1_2/temp4[68] , \MC_ARK_ARC_1_2/temp4[67] ,
         \MC_ARK_ARC_1_2/temp4[66] , \MC_ARK_ARC_1_2/temp4[64] ,
         \MC_ARK_ARC_1_2/temp4[63] , \MC_ARK_ARC_1_2/temp4[62] ,
         \MC_ARK_ARC_1_2/temp4[61] , \MC_ARK_ARC_1_2/temp4[60] ,
         \MC_ARK_ARC_1_2/temp4[58] , \MC_ARK_ARC_1_2/temp4[56] ,
         \MC_ARK_ARC_1_2/temp4[55] , \MC_ARK_ARC_1_2/temp4[54] ,
         \MC_ARK_ARC_1_2/temp4[53] , \MC_ARK_ARC_1_2/temp4[52] ,
         \MC_ARK_ARC_1_2/temp4[51] , \MC_ARK_ARC_1_2/temp4[50] ,
         \MC_ARK_ARC_1_2/temp4[49] , \MC_ARK_ARC_1_2/temp4[48] ,
         \MC_ARK_ARC_1_2/temp4[47] , \MC_ARK_ARC_1_2/temp4[46] ,
         \MC_ARK_ARC_1_2/temp4[45] , \MC_ARK_ARC_1_2/temp4[43] ,
         \MC_ARK_ARC_1_2/temp4[42] , \MC_ARK_ARC_1_2/temp4[40] ,
         \MC_ARK_ARC_1_2/temp4[39] , \MC_ARK_ARC_1_2/temp4[38] ,
         \MC_ARK_ARC_1_2/temp4[37] , \MC_ARK_ARC_1_2/temp4[36] ,
         \MC_ARK_ARC_1_2/temp4[35] , \MC_ARK_ARC_1_2/temp4[34] ,
         \MC_ARK_ARC_1_2/temp4[32] , \MC_ARK_ARC_1_2/temp4[31] ,
         \MC_ARK_ARC_1_2/temp4[30] , \MC_ARK_ARC_1_2/temp4[29] ,
         \MC_ARK_ARC_1_2/temp4[28] , \MC_ARK_ARC_1_2/temp4[27] ,
         \MC_ARK_ARC_1_2/temp4[26] , \MC_ARK_ARC_1_2/temp4[25] ,
         \MC_ARK_ARC_1_2/temp4[24] , \MC_ARK_ARC_1_2/temp4[22] ,
         \MC_ARK_ARC_1_2/temp4[21] , \MC_ARK_ARC_1_2/temp4[19] ,
         \MC_ARK_ARC_1_2/temp4[18] , \MC_ARK_ARC_1_2/temp4[16] ,
         \MC_ARK_ARC_1_2/temp4[15] , \MC_ARK_ARC_1_2/temp4[14] ,
         \MC_ARK_ARC_1_2/temp4[13] , \MC_ARK_ARC_1_2/temp4[12] ,
         \MC_ARK_ARC_1_2/temp4[11] , \MC_ARK_ARC_1_2/temp4[10] ,
         \MC_ARK_ARC_1_2/temp4[9] , \MC_ARK_ARC_1_2/temp4[8] ,
         \MC_ARK_ARC_1_2/temp4[7] , \MC_ARK_ARC_1_2/temp4[6] ,
         \MC_ARK_ARC_1_2/temp4[5] , \MC_ARK_ARC_1_2/temp4[4] ,
         \MC_ARK_ARC_1_2/temp4[3] , \MC_ARK_ARC_1_2/temp4[2] ,
         \MC_ARK_ARC_1_2/temp4[1] , \MC_ARK_ARC_1_2/temp4[0] ,
         \MC_ARK_ARC_1_2/temp3[190] , \MC_ARK_ARC_1_2/temp3[189] ,
         \MC_ARK_ARC_1_2/temp3[188] , \MC_ARK_ARC_1_2/temp3[187] ,
         \MC_ARK_ARC_1_2/temp3[186] , \MC_ARK_ARC_1_2/temp3[185] ,
         \MC_ARK_ARC_1_2/temp3[184] , \MC_ARK_ARC_1_2/temp3[182] ,
         \MC_ARK_ARC_1_2/temp3[177] , \MC_ARK_ARC_1_2/temp3[175] ,
         \MC_ARK_ARC_1_2/temp3[174] , \MC_ARK_ARC_1_2/temp3[173] ,
         \MC_ARK_ARC_1_2/temp3[172] , \MC_ARK_ARC_1_2/temp3[169] ,
         \MC_ARK_ARC_1_2/temp3[168] , \MC_ARK_ARC_1_2/temp3[167] ,
         \MC_ARK_ARC_1_2/temp3[166] , \MC_ARK_ARC_1_2/temp3[165] ,
         \MC_ARK_ARC_1_2/temp3[163] , \MC_ARK_ARC_1_2/temp3[161] ,
         \MC_ARK_ARC_1_2/temp3[160] , \MC_ARK_ARC_1_2/temp3[159] ,
         \MC_ARK_ARC_1_2/temp3[157] , \MC_ARK_ARC_1_2/temp3[156] ,
         \MC_ARK_ARC_1_2/temp3[154] , \MC_ARK_ARC_1_2/temp3[152] ,
         \MC_ARK_ARC_1_2/temp3[151] , \MC_ARK_ARC_1_2/temp3[150] ,
         \MC_ARK_ARC_1_2/temp3[149] , \MC_ARK_ARC_1_2/temp3[148] ,
         \MC_ARK_ARC_1_2/temp3[147] , \MC_ARK_ARC_1_2/temp3[146] ,
         \MC_ARK_ARC_1_2/temp3[145] , \MC_ARK_ARC_1_2/temp3[144] ,
         \MC_ARK_ARC_1_2/temp3[142] , \MC_ARK_ARC_1_2/temp3[141] ,
         \MC_ARK_ARC_1_2/temp3[138] , \MC_ARK_ARC_1_2/temp3[137] ,
         \MC_ARK_ARC_1_2/temp3[136] , \MC_ARK_ARC_1_2/temp3[135] ,
         \MC_ARK_ARC_1_2/temp3[134] , \MC_ARK_ARC_1_2/temp3[133] ,
         \MC_ARK_ARC_1_2/temp3[132] , \MC_ARK_ARC_1_2/temp3[131] ,
         \MC_ARK_ARC_1_2/temp3[130] , \MC_ARK_ARC_1_2/temp3[128] ,
         \MC_ARK_ARC_1_2/temp3[126] , \MC_ARK_ARC_1_2/temp3[125] ,
         \MC_ARK_ARC_1_2/temp3[124] , \MC_ARK_ARC_1_2/temp3[122] ,
         \MC_ARK_ARC_1_2/temp3[118] , \MC_ARK_ARC_1_2/temp3[117] ,
         \MC_ARK_ARC_1_2/temp3[116] , \MC_ARK_ARC_1_2/temp3[115] ,
         \MC_ARK_ARC_1_2/temp3[114] , \MC_ARK_ARC_1_2/temp3[112] ,
         \MC_ARK_ARC_1_2/temp3[109] , \MC_ARK_ARC_1_2/temp3[108] ,
         \MC_ARK_ARC_1_2/temp3[107] , \MC_ARK_ARC_1_2/temp3[106] ,
         \MC_ARK_ARC_1_2/temp3[105] , \MC_ARK_ARC_1_2/temp3[102] ,
         \MC_ARK_ARC_1_2/temp3[98] , \MC_ARK_ARC_1_2/temp3[97] ,
         \MC_ARK_ARC_1_2/temp3[96] , \MC_ARK_ARC_1_2/temp3[95] ,
         \MC_ARK_ARC_1_2/temp3[94] , \MC_ARK_ARC_1_2/temp3[93] ,
         \MC_ARK_ARC_1_2/temp3[91] , \MC_ARK_ARC_1_2/temp3[90] ,
         \MC_ARK_ARC_1_2/temp3[89] , \MC_ARK_ARC_1_2/temp3[88] ,
         \MC_ARK_ARC_1_2/temp3[86] , \MC_ARK_ARC_1_2/temp3[85] ,
         \MC_ARK_ARC_1_2/temp3[84] , \MC_ARK_ARC_1_2/temp3[83] ,
         \MC_ARK_ARC_1_2/temp3[82] , \MC_ARK_ARC_1_2/temp3[79] ,
         \MC_ARK_ARC_1_2/temp3[78] , \MC_ARK_ARC_1_2/temp3[77] ,
         \MC_ARK_ARC_1_2/temp3[76] , \MC_ARK_ARC_1_2/temp3[73] ,
         \MC_ARK_ARC_1_2/temp3[72] , \MC_ARK_ARC_1_2/temp3[71] ,
         \MC_ARK_ARC_1_2/temp3[70] , \MC_ARK_ARC_1_2/temp3[69] ,
         \MC_ARK_ARC_1_2/temp3[68] , \MC_ARK_ARC_1_2/temp3[66] ,
         \MC_ARK_ARC_1_2/temp3[64] , \MC_ARK_ARC_1_2/temp3[63] ,
         \MC_ARK_ARC_1_2/temp3[62] , \MC_ARK_ARC_1_2/temp3[61] ,
         \MC_ARK_ARC_1_2/temp3[60] , \MC_ARK_ARC_1_2/temp3[58] ,
         \MC_ARK_ARC_1_2/temp3[55] , \MC_ARK_ARC_1_2/temp3[53] ,
         \MC_ARK_ARC_1_2/temp3[52] , \MC_ARK_ARC_1_2/temp3[51] ,
         \MC_ARK_ARC_1_2/temp3[49] , \MC_ARK_ARC_1_2/temp3[47] ,
         \MC_ARK_ARC_1_2/temp3[46] , \MC_ARK_ARC_1_2/temp3[45] ,
         \MC_ARK_ARC_1_2/temp3[43] , \MC_ARK_ARC_1_2/temp3[42] ,
         \MC_ARK_ARC_1_2/temp3[40] , \MC_ARK_ARC_1_2/temp3[39] ,
         \MC_ARK_ARC_1_2/temp3[38] , \MC_ARK_ARC_1_2/temp3[37] ,
         \MC_ARK_ARC_1_2/temp3[36] , \MC_ARK_ARC_1_2/temp3[35] ,
         \MC_ARK_ARC_1_2/temp3[34] , \MC_ARK_ARC_1_2/temp3[32] ,
         \MC_ARK_ARC_1_2/temp3[31] , \MC_ARK_ARC_1_2/temp3[30] ,
         \MC_ARK_ARC_1_2/temp3[29] , \MC_ARK_ARC_1_2/temp3[27] ,
         \MC_ARK_ARC_1_2/temp3[26] , \MC_ARK_ARC_1_2/temp3[24] ,
         \MC_ARK_ARC_1_2/temp3[23] , \MC_ARK_ARC_1_2/temp3[22] ,
         \MC_ARK_ARC_1_2/temp3[21] , \MC_ARK_ARC_1_2/temp3[19] ,
         \MC_ARK_ARC_1_2/temp3[18] , \MC_ARK_ARC_1_2/temp3[17] ,
         \MC_ARK_ARC_1_2/temp3[16] , \MC_ARK_ARC_1_2/temp3[13] ,
         \MC_ARK_ARC_1_2/temp3[12] , \MC_ARK_ARC_1_2/temp3[11] ,
         \MC_ARK_ARC_1_2/temp3[10] , \MC_ARK_ARC_1_2/temp3[7] ,
         \MC_ARK_ARC_1_2/temp3[6] , \MC_ARK_ARC_1_2/temp3[5] ,
         \MC_ARK_ARC_1_2/temp3[4] , \MC_ARK_ARC_1_2/temp3[3] ,
         \MC_ARK_ARC_1_2/temp3[2] , \MC_ARK_ARC_1_2/temp3[1] ,
         \MC_ARK_ARC_1_2/temp3[0] , \MC_ARK_ARC_1_2/temp2[191] ,
         \MC_ARK_ARC_1_2/temp2[190] , \MC_ARK_ARC_1_2/temp2[188] ,
         \MC_ARK_ARC_1_2/temp2[187] , \MC_ARK_ARC_1_2/temp2[186] ,
         \MC_ARK_ARC_1_2/temp2[185] , \MC_ARK_ARC_1_2/temp2[181] ,
         \MC_ARK_ARC_1_2/temp2[180] , \MC_ARK_ARC_1_2/temp2[179] ,
         \MC_ARK_ARC_1_2/temp2[178] , \MC_ARK_ARC_1_2/temp2[177] ,
         \MC_ARK_ARC_1_2/temp2[176] , \MC_ARK_ARC_1_2/temp2[171] ,
         \MC_ARK_ARC_1_2/temp2[169] , \MC_ARK_ARC_1_2/temp2[168] ,
         \MC_ARK_ARC_1_2/temp2[166] , \MC_ARK_ARC_1_2/temp2[165] ,
         \MC_ARK_ARC_1_2/temp2[163] , \MC_ARK_ARC_1_2/temp2[162] ,
         \MC_ARK_ARC_1_2/temp2[160] , \MC_ARK_ARC_1_2/temp2[159] ,
         \MC_ARK_ARC_1_2/temp2[157] , \MC_ARK_ARC_1_2/temp2[156] ,
         \MC_ARK_ARC_1_2/temp2[153] , \MC_ARK_ARC_1_2/temp2[151] ,
         \MC_ARK_ARC_1_2/temp2[150] , \MC_ARK_ARC_1_2/temp2[149] ,
         \MC_ARK_ARC_1_2/temp2[148] , \MC_ARK_ARC_1_2/temp2[146] ,
         \MC_ARK_ARC_1_2/temp2[145] , \MC_ARK_ARC_1_2/temp2[143] ,
         \MC_ARK_ARC_1_2/temp2[142] , \MC_ARK_ARC_1_2/temp2[141] ,
         \MC_ARK_ARC_1_2/temp2[140] , \MC_ARK_ARC_1_2/temp2[138] ,
         \MC_ARK_ARC_1_2/temp2[136] , \MC_ARK_ARC_1_2/temp2[135] ,
         \MC_ARK_ARC_1_2/temp2[132] , \MC_ARK_ARC_1_2/temp2[131] ,
         \MC_ARK_ARC_1_2/temp2[130] , \MC_ARK_ARC_1_2/temp2[129] ,
         \MC_ARK_ARC_1_2/temp2[128] , \MC_ARK_ARC_1_2/temp2[127] ,
         \MC_ARK_ARC_1_2/temp2[126] , \MC_ARK_ARC_1_2/temp2[124] ,
         \MC_ARK_ARC_1_2/temp2[119] , \MC_ARK_ARC_1_2/temp2[118] ,
         \MC_ARK_ARC_1_2/temp2[116] , \MC_ARK_ARC_1_2/temp2[115] ,
         \MC_ARK_ARC_1_2/temp2[114] , \MC_ARK_ARC_1_2/temp2[112] ,
         \MC_ARK_ARC_1_2/temp2[111] , \MC_ARK_ARC_1_2/temp2[109] ,
         \MC_ARK_ARC_1_2/temp2[107] , \MC_ARK_ARC_1_2/temp2[106] ,
         \MC_ARK_ARC_1_2/temp2[104] , \MC_ARK_ARC_1_2/temp2[103] ,
         \MC_ARK_ARC_1_2/temp2[102] , \MC_ARK_ARC_1_2/temp2[100] ,
         \MC_ARK_ARC_1_2/temp2[98] , \MC_ARK_ARC_1_2/temp2[97] ,
         \MC_ARK_ARC_1_2/temp2[96] , \MC_ARK_ARC_1_2/temp2[95] ,
         \MC_ARK_ARC_1_2/temp2[94] , \MC_ARK_ARC_1_2/temp2[92] ,
         \MC_ARK_ARC_1_2/temp2[91] , \MC_ARK_ARC_1_2/temp2[90] ,
         \MC_ARK_ARC_1_2/temp2[88] , \MC_ARK_ARC_1_2/temp2[85] ,
         \MC_ARK_ARC_1_2/temp2[83] , \MC_ARK_ARC_1_2/temp2[82] ,
         \MC_ARK_ARC_1_2/temp2[81] , \MC_ARK_ARC_1_2/temp2[80] ,
         \MC_ARK_ARC_1_2/temp2[79] , \MC_ARK_ARC_1_2/temp2[78] ,
         \MC_ARK_ARC_1_2/temp2[77] , \MC_ARK_ARC_1_2/temp2[76] ,
         \MC_ARK_ARC_1_2/temp2[74] , \MC_ARK_ARC_1_2/temp2[73] ,
         \MC_ARK_ARC_1_2/temp2[72] , \MC_ARK_ARC_1_2/temp2[71] ,
         \MC_ARK_ARC_1_2/temp2[67] , \MC_ARK_ARC_1_2/temp2[66] ,
         \MC_ARK_ARC_1_2/temp2[64] , \MC_ARK_ARC_1_2/temp2[62] ,
         \MC_ARK_ARC_1_2/temp2[61] , \MC_ARK_ARC_1_2/temp2[60] ,
         \MC_ARK_ARC_1_2/temp2[58] , \MC_ARK_ARC_1_2/temp2[57] ,
         \MC_ARK_ARC_1_2/temp2[56] , \MC_ARK_ARC_1_2/temp2[55] ,
         \MC_ARK_ARC_1_2/temp2[54] , \MC_ARK_ARC_1_2/temp2[52] ,
         \MC_ARK_ARC_1_2/temp2[48] , \MC_ARK_ARC_1_2/temp2[47] ,
         \MC_ARK_ARC_1_2/temp2[46] , \MC_ARK_ARC_1_2/temp2[45] ,
         \MC_ARK_ARC_1_2/temp2[44] , \MC_ARK_ARC_1_2/temp2[42] ,
         \MC_ARK_ARC_1_2/temp2[40] , \MC_ARK_ARC_1_2/temp2[37] ,
         \MC_ARK_ARC_1_2/temp2[36] , \MC_ARK_ARC_1_2/temp2[32] ,
         \MC_ARK_ARC_1_2/temp2[31] , \MC_ARK_ARC_1_2/temp2[30] ,
         \MC_ARK_ARC_1_2/temp2[29] , \MC_ARK_ARC_1_2/temp2[27] ,
         \MC_ARK_ARC_1_2/temp2[25] , \MC_ARK_ARC_1_2/temp2[24] ,
         \MC_ARK_ARC_1_2/temp2[23] , \MC_ARK_ARC_1_2/temp2[21] ,
         \MC_ARK_ARC_1_2/temp2[20] , \MC_ARK_ARC_1_2/temp2[19] ,
         \MC_ARK_ARC_1_2/temp2[16] , \MC_ARK_ARC_1_2/temp2[13] ,
         \MC_ARK_ARC_1_2/temp2[12] , \MC_ARK_ARC_1_2/temp2[11] ,
         \MC_ARK_ARC_1_2/temp2[10] , \MC_ARK_ARC_1_2/temp2[9] ,
         \MC_ARK_ARC_1_2/temp2[7] , \MC_ARK_ARC_1_2/temp2[6] ,
         \MC_ARK_ARC_1_2/temp2[4] , \MC_ARK_ARC_1_2/temp2[3] ,
         \MC_ARK_ARC_1_2/temp2[1] , \MC_ARK_ARC_1_2/temp1[191] ,
         \MC_ARK_ARC_1_2/temp1[190] , \MC_ARK_ARC_1_2/temp1[189] ,
         \MC_ARK_ARC_1_2/temp1[188] , \MC_ARK_ARC_1_2/temp1[185] ,
         \MC_ARK_ARC_1_2/temp1[184] , \MC_ARK_ARC_1_2/temp1[182] ,
         \MC_ARK_ARC_1_2/temp1[181] , \MC_ARK_ARC_1_2/temp1[180] ,
         \MC_ARK_ARC_1_2/temp1[178] , \MC_ARK_ARC_1_2/temp1[176] ,
         \MC_ARK_ARC_1_2/temp1[175] , \MC_ARK_ARC_1_2/temp1[174] ,
         \MC_ARK_ARC_1_2/temp1[173] , \MC_ARK_ARC_1_2/temp1[168] ,
         \MC_ARK_ARC_1_2/temp1[167] , \MC_ARK_ARC_1_2/temp1[166] ,
         \MC_ARK_ARC_1_2/temp1[165] , \MC_ARK_ARC_1_2/temp1[163] ,
         \MC_ARK_ARC_1_2/temp1[161] , \MC_ARK_ARC_1_2/temp1[157] ,
         \MC_ARK_ARC_1_2/temp1[156] , \MC_ARK_ARC_1_2/temp1[153] ,
         \MC_ARK_ARC_1_2/temp1[151] , \MC_ARK_ARC_1_2/temp1[150] ,
         \MC_ARK_ARC_1_2/temp1[149] , \MC_ARK_ARC_1_2/temp1[148] ,
         \MC_ARK_ARC_1_2/temp1[145] , \MC_ARK_ARC_1_2/temp1[144] ,
         \MC_ARK_ARC_1_2/temp1[143] , \MC_ARK_ARC_1_2/temp1[142] ,
         \MC_ARK_ARC_1_2/temp1[141] , \MC_ARK_ARC_1_2/temp1[139] ,
         \MC_ARK_ARC_1_2/temp1[137] , \MC_ARK_ARC_1_2/temp1[136] ,
         \MC_ARK_ARC_1_2/temp1[135] , \MC_ARK_ARC_1_2/temp1[134] ,
         \MC_ARK_ARC_1_2/temp1[133] , \MC_ARK_ARC_1_2/temp1[132] ,
         \MC_ARK_ARC_1_2/temp1[130] , \MC_ARK_ARC_1_2/temp1[127] ,
         \MC_ARK_ARC_1_2/temp1[126] , \MC_ARK_ARC_1_2/temp1[125] ,
         \MC_ARK_ARC_1_2/temp1[123] , \MC_ARK_ARC_1_2/temp1[122] ,
         \MC_ARK_ARC_1_2/temp1[121] , \MC_ARK_ARC_1_2/temp1[120] ,
         \MC_ARK_ARC_1_2/temp1[118] , \MC_ARK_ARC_1_2/temp1[117] ,
         \MC_ARK_ARC_1_2/temp1[116] , \MC_ARK_ARC_1_2/temp1[114] ,
         \MC_ARK_ARC_1_2/temp1[112] , \MC_ARK_ARC_1_2/temp1[111] ,
         \MC_ARK_ARC_1_2/temp1[109] , \MC_ARK_ARC_1_2/temp1[108] ,
         \MC_ARK_ARC_1_2/temp1[106] , \MC_ARK_ARC_1_2/temp1[105] ,
         \MC_ARK_ARC_1_2/temp1[104] , \MC_ARK_ARC_1_2/temp1[103] ,
         \MC_ARK_ARC_1_2/temp1[102] , \MC_ARK_ARC_1_2/temp1[101] ,
         \MC_ARK_ARC_1_2/temp1[100] , \MC_ARK_ARC_1_2/temp1[97] ,
         \MC_ARK_ARC_1_2/temp1[96] , \MC_ARK_ARC_1_2/temp1[94] ,
         \MC_ARK_ARC_1_2/temp1[93] , \MC_ARK_ARC_1_2/temp1[91] ,
         \MC_ARK_ARC_1_2/temp1[88] , \MC_ARK_ARC_1_2/temp1[87] ,
         \MC_ARK_ARC_1_2/temp1[86] , \MC_ARK_ARC_1_2/temp1[84] ,
         \MC_ARK_ARC_1_2/temp1[83] , \MC_ARK_ARC_1_2/temp1[82] ,
         \MC_ARK_ARC_1_2/temp1[81] , \MC_ARK_ARC_1_2/temp1[79] ,
         \MC_ARK_ARC_1_2/temp1[78] , \MC_ARK_ARC_1_2/temp1[77] ,
         \MC_ARK_ARC_1_2/temp1[76] , \MC_ARK_ARC_1_2/temp1[73] ,
         \MC_ARK_ARC_1_2/temp1[72] , \MC_ARK_ARC_1_2/temp1[70] ,
         \MC_ARK_ARC_1_2/temp1[69] , \MC_ARK_ARC_1_2/temp1[67] ,
         \MC_ARK_ARC_1_2/temp1[66] , \MC_ARK_ARC_1_2/temp1[64] ,
         \MC_ARK_ARC_1_2/temp1[62] , \MC_ARK_ARC_1_2/temp1[61] ,
         \MC_ARK_ARC_1_2/temp1[59] , \MC_ARK_ARC_1_2/temp1[56] ,
         \MC_ARK_ARC_1_2/temp1[55] , \MC_ARK_ARC_1_2/temp1[54] ,
         \MC_ARK_ARC_1_2/temp1[52] , \MC_ARK_ARC_1_2/temp1[49] ,
         \MC_ARK_ARC_1_2/temp1[47] , \MC_ARK_ARC_1_2/temp1[46] ,
         \MC_ARK_ARC_1_2/temp1[45] , \MC_ARK_ARC_1_2/temp1[43] ,
         \MC_ARK_ARC_1_2/temp1[42] , \MC_ARK_ARC_1_2/temp1[40] ,
         \MC_ARK_ARC_1_2/temp1[38] , \MC_ARK_ARC_1_2/temp1[37] ,
         \MC_ARK_ARC_1_2/temp1[36] , \MC_ARK_ARC_1_2/temp1[34] ,
         \MC_ARK_ARC_1_2/temp1[31] , \MC_ARK_ARC_1_2/temp1[30] ,
         \MC_ARK_ARC_1_2/temp1[29] , \MC_ARK_ARC_1_2/temp1[27] ,
         \MC_ARK_ARC_1_2/temp1[25] , \MC_ARK_ARC_1_2/temp1[24] ,
         \MC_ARK_ARC_1_2/temp1[22] , \MC_ARK_ARC_1_2/temp1[21] ,
         \MC_ARK_ARC_1_2/temp1[19] , \MC_ARK_ARC_1_2/temp1[18] ,
         \MC_ARK_ARC_1_2/temp1[17] , \MC_ARK_ARC_1_2/temp1[16] ,
         \MC_ARK_ARC_1_2/temp1[15] , \MC_ARK_ARC_1_2/temp1[14] ,
         \MC_ARK_ARC_1_2/temp1[13] , \MC_ARK_ARC_1_2/temp1[12] ,
         \MC_ARK_ARC_1_2/temp1[6] , \MC_ARK_ARC_1_2/temp1[4] ,
         \MC_ARK_ARC_1_2/temp1[1] , \MC_ARK_ARC_1_2/temp1[0] ,
         \MC_ARK_ARC_1_2/buf_keyinput[79] ,
         \MC_ARK_ARC_1_2/buf_datainput[183] ,
         \MC_ARK_ARC_1_2/buf_datainput[181] ,
         \MC_ARK_ARC_1_2/buf_datainput[179] ,
         \MC_ARK_ARC_1_2/buf_datainput[172] ,
         \MC_ARK_ARC_1_2/buf_datainput[171] ,
         \MC_ARK_ARC_1_2/buf_datainput[164] ,
         \MC_ARK_ARC_1_2/buf_datainput[162] ,
         \MC_ARK_ARC_1_2/buf_datainput[151] ,
         \MC_ARK_ARC_1_2/buf_datainput[150] ,
         \MC_ARK_ARC_1_2/buf_datainput[147] ,
         \MC_ARK_ARC_1_2/buf_datainput[146] ,
         \MC_ARK_ARC_1_2/buf_datainput[143] ,
         \MC_ARK_ARC_1_2/buf_datainput[141] ,
         \MC_ARK_ARC_1_2/buf_datainput[133] ,
         \MC_ARK_ARC_1_2/buf_datainput[131] ,
         \MC_ARK_ARC_1_2/buf_datainput[124] ,
         \MC_ARK_ARC_1_2/buf_datainput[122] ,
         \MC_ARK_ARC_1_2/buf_datainput[121] ,
         \MC_ARK_ARC_1_2/buf_datainput[120] ,
         \MC_ARK_ARC_1_2/buf_datainput[115] ,
         \MC_ARK_ARC_1_2/buf_datainput[112] ,
         \MC_ARK_ARC_1_2/buf_datainput[110] ,
         \MC_ARK_ARC_1_2/buf_datainput[106] ,
         \MC_ARK_ARC_1_2/buf_datainput[100] ,
         \MC_ARK_ARC_1_2/buf_datainput[99] ,
         \MC_ARK_ARC_1_2/buf_datainput[98] ,
         \MC_ARK_ARC_1_2/buf_datainput[92] ,
         \MC_ARK_ARC_1_2/buf_datainput[89] ,
         \MC_ARK_ARC_1_2/buf_datainput[84] ,
         \MC_ARK_ARC_1_2/buf_datainput[79] ,
         \MC_ARK_ARC_1_2/buf_datainput[74] ,
         \MC_ARK_ARC_1_2/buf_datainput[70] ,
         \MC_ARK_ARC_1_2/buf_datainput[68] ,
         \MC_ARK_ARC_1_2/buf_datainput[65] ,
         \MC_ARK_ARC_1_2/buf_datainput[63] ,
         \MC_ARK_ARC_1_2/buf_datainput[61] ,
         \MC_ARK_ARC_1_2/buf_datainput[60] ,
         \MC_ARK_ARC_1_2/buf_datainput[56] ,
         \MC_ARK_ARC_1_2/buf_datainput[55] ,
         \MC_ARK_ARC_1_2/buf_datainput[52] ,
         \MC_ARK_ARC_1_2/buf_datainput[49] ,
         \MC_ARK_ARC_1_2/buf_datainput[45] ,
         \MC_ARK_ARC_1_2/buf_datainput[41] ,
         \MC_ARK_ARC_1_2/buf_datainput[40] ,
         \MC_ARK_ARC_1_2/buf_datainput[35] ,
         \MC_ARK_ARC_1_2/buf_datainput[29] ,
         \MC_ARK_ARC_1_2/buf_datainput[28] ,
         \MC_ARK_ARC_1_2/buf_datainput[25] ,
         \MC_ARK_ARC_1_2/buf_datainput[24] ,
         \MC_ARK_ARC_1_2/buf_datainput[23] ,
         \MC_ARK_ARC_1_2/buf_datainput[22] ,
         \MC_ARK_ARC_1_2/buf_datainput[14] ,
         \MC_ARK_ARC_1_2/buf_datainput[10] , \MC_ARK_ARC_1_2/buf_datainput[7] ,
         \MC_ARK_ARC_1_2/buf_datainput[3] , \MC_ARK_ARC_1_3/buf_output[191] ,
         \MC_ARK_ARC_1_3/buf_output[190] , \MC_ARK_ARC_1_3/buf_output[189] ,
         \MC_ARK_ARC_1_3/buf_output[188] , \MC_ARK_ARC_1_3/buf_output[187] ,
         \MC_ARK_ARC_1_3/buf_output[186] , \MC_ARK_ARC_1_3/buf_output[185] ,
         \MC_ARK_ARC_1_3/buf_output[184] , \MC_ARK_ARC_1_3/buf_output[183] ,
         \MC_ARK_ARC_1_3/buf_output[182] , \MC_ARK_ARC_1_3/buf_output[181] ,
         \MC_ARK_ARC_1_3/buf_output[180] , \MC_ARK_ARC_1_3/buf_output[179] ,
         \MC_ARK_ARC_1_3/buf_output[178] , \MC_ARK_ARC_1_3/buf_output[177] ,
         \MC_ARK_ARC_1_3/buf_output[176] , \MC_ARK_ARC_1_3/buf_output[175] ,
         \MC_ARK_ARC_1_3/buf_output[174] , \MC_ARK_ARC_1_3/buf_output[172] ,
         \MC_ARK_ARC_1_3/buf_output[171] , \MC_ARK_ARC_1_3/buf_output[170] ,
         \MC_ARK_ARC_1_3/buf_output[169] , \MC_ARK_ARC_1_3/buf_output[168] ,
         \MC_ARK_ARC_1_3/buf_output[167] , \MC_ARK_ARC_1_3/buf_output[166] ,
         \MC_ARK_ARC_1_3/buf_output[165] , \MC_ARK_ARC_1_3/buf_output[164] ,
         \MC_ARK_ARC_1_3/buf_output[163] , \MC_ARK_ARC_1_3/buf_output[162] ,
         \MC_ARK_ARC_1_3/buf_output[161] , \MC_ARK_ARC_1_3/buf_output[160] ,
         \MC_ARK_ARC_1_3/buf_output[159] , \MC_ARK_ARC_1_3/buf_output[158] ,
         \MC_ARK_ARC_1_3/buf_output[157] , \MC_ARK_ARC_1_3/buf_output[156] ,
         \MC_ARK_ARC_1_3/buf_output[155] , \MC_ARK_ARC_1_3/buf_output[154] ,
         \MC_ARK_ARC_1_3/buf_output[152] , \MC_ARK_ARC_1_3/buf_output[151] ,
         \MC_ARK_ARC_1_3/buf_output[150] , \MC_ARK_ARC_1_3/buf_output[149] ,
         \MC_ARK_ARC_1_3/buf_output[148] , \MC_ARK_ARC_1_3/buf_output[147] ,
         \MC_ARK_ARC_1_3/buf_output[146] , \MC_ARK_ARC_1_3/buf_output[145] ,
         \MC_ARK_ARC_1_3/buf_output[144] , \MC_ARK_ARC_1_3/buf_output[143] ,
         \MC_ARK_ARC_1_3/buf_output[142] , \MC_ARK_ARC_1_3/buf_output[139] ,
         \MC_ARK_ARC_1_3/buf_output[138] , \MC_ARK_ARC_1_3/buf_output[136] ,
         \MC_ARK_ARC_1_3/buf_output[135] , \MC_ARK_ARC_1_3/buf_output[134] ,
         \MC_ARK_ARC_1_3/buf_output[133] , \MC_ARK_ARC_1_3/buf_output[132] ,
         \MC_ARK_ARC_1_3/buf_output[131] , \MC_ARK_ARC_1_3/buf_output[130] ,
         \MC_ARK_ARC_1_3/buf_output[128] , \MC_ARK_ARC_1_3/buf_output[127] ,
         \MC_ARK_ARC_1_3/buf_output[126] , \MC_ARK_ARC_1_3/buf_output[125] ,
         \MC_ARK_ARC_1_3/buf_output[124] , \MC_ARK_ARC_1_3/buf_output[123] ,
         \MC_ARK_ARC_1_3/buf_output[122] , \MC_ARK_ARC_1_3/buf_output[121] ,
         \MC_ARK_ARC_1_3/buf_output[120] , \MC_ARK_ARC_1_3/buf_output[119] ,
         \MC_ARK_ARC_1_3/buf_output[118] , \MC_ARK_ARC_1_3/buf_output[117] ,
         \MC_ARK_ARC_1_3/buf_output[116] , \MC_ARK_ARC_1_3/buf_output[115] ,
         \MC_ARK_ARC_1_3/buf_output[114] , \MC_ARK_ARC_1_3/buf_output[113] ,
         \MC_ARK_ARC_1_3/buf_output[112] , \MC_ARK_ARC_1_3/buf_output[111] ,
         \MC_ARK_ARC_1_3/buf_output[110] , \MC_ARK_ARC_1_3/buf_output[109] ,
         \MC_ARK_ARC_1_3/buf_output[108] , \MC_ARK_ARC_1_3/buf_output[107] ,
         \MC_ARK_ARC_1_3/buf_output[106] , \MC_ARK_ARC_1_3/buf_output[104] ,
         \MC_ARK_ARC_1_3/buf_output[103] , \MC_ARK_ARC_1_3/buf_output[102] ,
         \MC_ARK_ARC_1_3/buf_output[101] , \MC_ARK_ARC_1_3/buf_output[100] ,
         \MC_ARK_ARC_1_3/buf_output[99] , \MC_ARK_ARC_1_3/buf_output[98] ,
         \MC_ARK_ARC_1_3/buf_output[97] , \MC_ARK_ARC_1_3/buf_output[96] ,
         \MC_ARK_ARC_1_3/buf_output[95] , \MC_ARK_ARC_1_3/buf_output[94] ,
         \MC_ARK_ARC_1_3/buf_output[93] , \MC_ARK_ARC_1_3/buf_output[92] ,
         \MC_ARK_ARC_1_3/buf_output[91] , \MC_ARK_ARC_1_3/buf_output[90] ,
         \MC_ARK_ARC_1_3/buf_output[89] , \MC_ARK_ARC_1_3/buf_output[88] ,
         \MC_ARK_ARC_1_3/buf_output[87] , \MC_ARK_ARC_1_3/buf_output[86] ,
         \MC_ARK_ARC_1_3/buf_output[85] , \MC_ARK_ARC_1_3/buf_output[84] ,
         \MC_ARK_ARC_1_3/buf_output[83] , \MC_ARK_ARC_1_3/buf_output[82] ,
         \MC_ARK_ARC_1_3/buf_output[81] , \MC_ARK_ARC_1_3/buf_output[80] ,
         \MC_ARK_ARC_1_3/buf_output[79] , \MC_ARK_ARC_1_3/buf_output[78] ,
         \MC_ARK_ARC_1_3/buf_output[77] , \MC_ARK_ARC_1_3/buf_output[76] ,
         \MC_ARK_ARC_1_3/buf_output[75] , \MC_ARK_ARC_1_3/buf_output[74] ,
         \MC_ARK_ARC_1_3/buf_output[73] , \MC_ARK_ARC_1_3/buf_output[72] ,
         \MC_ARK_ARC_1_3/buf_output[71] , \MC_ARK_ARC_1_3/buf_output[70] ,
         \MC_ARK_ARC_1_3/buf_output[69] , \MC_ARK_ARC_1_3/buf_output[68] ,
         \MC_ARK_ARC_1_3/buf_output[67] , \MC_ARK_ARC_1_3/buf_output[66] ,
         \MC_ARK_ARC_1_3/buf_output[64] , \MC_ARK_ARC_1_3/buf_output[63] ,
         \MC_ARK_ARC_1_3/buf_output[62] , \MC_ARK_ARC_1_3/buf_output[61] ,
         \MC_ARK_ARC_1_3/buf_output[60] , \MC_ARK_ARC_1_3/buf_output[59] ,
         \MC_ARK_ARC_1_3/buf_output[58] , \MC_ARK_ARC_1_3/buf_output[57] ,
         \MC_ARK_ARC_1_3/buf_output[56] , \MC_ARK_ARC_1_3/buf_output[55] ,
         \MC_ARK_ARC_1_3/buf_output[54] , \MC_ARK_ARC_1_3/buf_output[52] ,
         \MC_ARK_ARC_1_3/buf_output[51] , \MC_ARK_ARC_1_3/buf_output[50] ,
         \MC_ARK_ARC_1_3/buf_output[49] , \MC_ARK_ARC_1_3/buf_output[48] ,
         \MC_ARK_ARC_1_3/buf_output[47] , \MC_ARK_ARC_1_3/buf_output[46] ,
         \MC_ARK_ARC_1_3/buf_output[45] , \MC_ARK_ARC_1_3/buf_output[44] ,
         \MC_ARK_ARC_1_3/buf_output[43] , \MC_ARK_ARC_1_3/buf_output[42] ,
         \MC_ARK_ARC_1_3/buf_output[41] , \MC_ARK_ARC_1_3/buf_output[40] ,
         \MC_ARK_ARC_1_3/buf_output[39] , \MC_ARK_ARC_1_3/buf_output[38] ,
         \MC_ARK_ARC_1_3/buf_output[37] , \MC_ARK_ARC_1_3/buf_output[36] ,
         \MC_ARK_ARC_1_3/buf_output[35] , \MC_ARK_ARC_1_3/buf_output[34] ,
         \MC_ARK_ARC_1_3/buf_output[33] , \MC_ARK_ARC_1_3/buf_output[32] ,
         \MC_ARK_ARC_1_3/buf_output[31] , \MC_ARK_ARC_1_3/buf_output[30] ,
         \MC_ARK_ARC_1_3/buf_output[29] , \MC_ARK_ARC_1_3/buf_output[28] ,
         \MC_ARK_ARC_1_3/buf_output[27] , \MC_ARK_ARC_1_3/buf_output[26] ,
         \MC_ARK_ARC_1_3/buf_output[25] , \MC_ARK_ARC_1_3/buf_output[24] ,
         \MC_ARK_ARC_1_3/buf_output[23] , \MC_ARK_ARC_1_3/buf_output[22] ,
         \MC_ARK_ARC_1_3/buf_output[21] , \MC_ARK_ARC_1_3/buf_output[20] ,
         \MC_ARK_ARC_1_3/buf_output[19] , \MC_ARK_ARC_1_3/buf_output[18] ,
         \MC_ARK_ARC_1_3/buf_output[17] , \MC_ARK_ARC_1_3/buf_output[16] ,
         \MC_ARK_ARC_1_3/buf_output[15] , \MC_ARK_ARC_1_3/buf_output[14] ,
         \MC_ARK_ARC_1_3/buf_output[13] , \MC_ARK_ARC_1_3/buf_output[12] ,
         \MC_ARK_ARC_1_3/buf_output[10] , \MC_ARK_ARC_1_3/buf_output[9] ,
         \MC_ARK_ARC_1_3/buf_output[8] , \MC_ARK_ARC_1_3/buf_output[7] ,
         \MC_ARK_ARC_1_3/buf_output[6] , \MC_ARK_ARC_1_3/buf_output[4] ,
         \MC_ARK_ARC_1_3/buf_output[3] , \MC_ARK_ARC_1_3/buf_output[2] ,
         \MC_ARK_ARC_1_3/buf_output[1] , \MC_ARK_ARC_1_3/buf_output[0] ,
         \MC_ARK_ARC_1_3/temp6[190] , \MC_ARK_ARC_1_3/temp6[188] ,
         \MC_ARK_ARC_1_3/temp6[186] , \MC_ARK_ARC_1_3/temp6[184] ,
         \MC_ARK_ARC_1_3/temp6[175] , \MC_ARK_ARC_1_3/temp6[174] ,
         \MC_ARK_ARC_1_3/temp6[173] , \MC_ARK_ARC_1_3/temp6[171] ,
         \MC_ARK_ARC_1_3/temp6[169] , \MC_ARK_ARC_1_3/temp6[168] ,
         \MC_ARK_ARC_1_3/temp6[166] , \MC_ARK_ARC_1_3/temp6[165] ,
         \MC_ARK_ARC_1_3/temp6[164] , \MC_ARK_ARC_1_3/temp6[163] ,
         \MC_ARK_ARC_1_3/temp6[161] , \MC_ARK_ARC_1_3/temp6[160] ,
         \MC_ARK_ARC_1_3/temp6[157] , \MC_ARK_ARC_1_3/temp6[156] ,
         \MC_ARK_ARC_1_3/temp6[153] , \MC_ARK_ARC_1_3/temp6[151] ,
         \MC_ARK_ARC_1_3/temp6[150] , \MC_ARK_ARC_1_3/temp6[149] ,
         \MC_ARK_ARC_1_3/temp6[148] , \MC_ARK_ARC_1_3/temp6[146] ,
         \MC_ARK_ARC_1_3/temp6[145] , \MC_ARK_ARC_1_3/temp6[144] ,
         \MC_ARK_ARC_1_3/temp6[142] , \MC_ARK_ARC_1_3/temp6[139] ,
         \MC_ARK_ARC_1_3/temp6[138] , \MC_ARK_ARC_1_3/temp6[133] ,
         \MC_ARK_ARC_1_3/temp6[132] , \MC_ARK_ARC_1_3/temp6[130] ,
         \MC_ARK_ARC_1_3/temp6[129] , \MC_ARK_ARC_1_3/temp6[128] ,
         \MC_ARK_ARC_1_3/temp6[126] , \MC_ARK_ARC_1_3/temp6[123] ,
         \MC_ARK_ARC_1_3/temp6[121] , \MC_ARK_ARC_1_3/temp6[120] ,
         \MC_ARK_ARC_1_3/temp6[119] , \MC_ARK_ARC_1_3/temp6[116] ,
         \MC_ARK_ARC_1_3/temp6[113] , \MC_ARK_ARC_1_3/temp6[112] ,
         \MC_ARK_ARC_1_3/temp6[111] , \MC_ARK_ARC_1_3/temp6[108] ,
         \MC_ARK_ARC_1_3/temp6[106] , \MC_ARK_ARC_1_3/temp6[105] ,
         \MC_ARK_ARC_1_3/temp6[103] , \MC_ARK_ARC_1_3/temp6[101] ,
         \MC_ARK_ARC_1_3/temp6[97] , \MC_ARK_ARC_1_3/temp6[96] ,
         \MC_ARK_ARC_1_3/temp6[94] , \MC_ARK_ARC_1_3/temp6[93] ,
         \MC_ARK_ARC_1_3/temp6[92] , \MC_ARK_ARC_1_3/temp6[89] ,
         \MC_ARK_ARC_1_3/temp6[88] , \MC_ARK_ARC_1_3/temp6[85] ,
         \MC_ARK_ARC_1_3/temp6[84] , \MC_ARK_ARC_1_3/temp6[82] ,
         \MC_ARK_ARC_1_3/temp6[79] , \MC_ARK_ARC_1_3/temp6[78] ,
         \MC_ARK_ARC_1_3/temp6[76] , \MC_ARK_ARC_1_3/temp6[72] ,
         \MC_ARK_ARC_1_3/temp6[70] , \MC_ARK_ARC_1_3/temp6[68] ,
         \MC_ARK_ARC_1_3/temp6[66] , \MC_ARK_ARC_1_3/temp6[65] ,
         \MC_ARK_ARC_1_3/temp6[61] , \MC_ARK_ARC_1_3/temp6[57] ,
         \MC_ARK_ARC_1_3/temp6[52] , \MC_ARK_ARC_1_3/temp6[50] ,
         \MC_ARK_ARC_1_3/temp6[49] , \MC_ARK_ARC_1_3/temp6[48] ,
         \MC_ARK_ARC_1_3/temp6[46] , \MC_ARK_ARC_1_3/temp6[43] ,
         \MC_ARK_ARC_1_3/temp6[40] , \MC_ARK_ARC_1_3/temp6[34] ,
         \MC_ARK_ARC_1_3/temp6[31] , \MC_ARK_ARC_1_3/temp6[30] ,
         \MC_ARK_ARC_1_3/temp6[28] , \MC_ARK_ARC_1_3/temp6[25] ,
         \MC_ARK_ARC_1_3/temp6[24] , \MC_ARK_ARC_1_3/temp6[23] ,
         \MC_ARK_ARC_1_3/temp6[22] , \MC_ARK_ARC_1_3/temp6[19] ,
         \MC_ARK_ARC_1_3/temp6[15] , \MC_ARK_ARC_1_3/temp6[13] ,
         \MC_ARK_ARC_1_3/temp6[11] , \MC_ARK_ARC_1_3/temp6[9] ,
         \MC_ARK_ARC_1_3/temp6[8] , \MC_ARK_ARC_1_3/temp6[7] ,
         \MC_ARK_ARC_1_3/temp6[6] , \MC_ARK_ARC_1_3/temp6[5] ,
         \MC_ARK_ARC_1_3/temp6[4] , \MC_ARK_ARC_1_3/temp6[3] ,
         \MC_ARK_ARC_1_3/temp6[2] , \MC_ARK_ARC_1_3/temp6[1] ,
         \MC_ARK_ARC_1_3/temp5[188] , \MC_ARK_ARC_1_3/temp5[187] ,
         \MC_ARK_ARC_1_3/temp5[186] , \MC_ARK_ARC_1_3/temp5[181] ,
         \MC_ARK_ARC_1_3/temp5[179] , \MC_ARK_ARC_1_3/temp5[178] ,
         \MC_ARK_ARC_1_3/temp5[172] , \MC_ARK_ARC_1_3/temp5[169] ,
         \MC_ARK_ARC_1_3/temp5[168] , \MC_ARK_ARC_1_3/temp5[162] ,
         \MC_ARK_ARC_1_3/temp5[161] , \MC_ARK_ARC_1_3/temp5[160] ,
         \MC_ARK_ARC_1_3/temp5[159] , \MC_ARK_ARC_1_3/temp5[158] ,
         \MC_ARK_ARC_1_3/temp5[156] , \MC_ARK_ARC_1_3/temp5[153] ,
         \MC_ARK_ARC_1_3/temp5[152] , \MC_ARK_ARC_1_3/temp5[151] ,
         \MC_ARK_ARC_1_3/temp5[149] , \MC_ARK_ARC_1_3/temp5[148] ,
         \MC_ARK_ARC_1_3/temp5[146] , \MC_ARK_ARC_1_3/temp5[145] ,
         \MC_ARK_ARC_1_3/temp5[144] , \MC_ARK_ARC_1_3/temp5[142] ,
         \MC_ARK_ARC_1_3/temp5[140] , \MC_ARK_ARC_1_3/temp5[139] ,
         \MC_ARK_ARC_1_3/temp5[136] , \MC_ARK_ARC_1_3/temp5[131] ,
         \MC_ARK_ARC_1_3/temp5[128] , \MC_ARK_ARC_1_3/temp5[127] ,
         \MC_ARK_ARC_1_3/temp5[122] , \MC_ARK_ARC_1_3/temp5[121] ,
         \MC_ARK_ARC_1_3/temp5[120] , \MC_ARK_ARC_1_3/temp5[116] ,
         \MC_ARK_ARC_1_3/temp5[115] , \MC_ARK_ARC_1_3/temp5[112] ,
         \MC_ARK_ARC_1_3/temp5[111] , \MC_ARK_ARC_1_3/temp5[110] ,
         \MC_ARK_ARC_1_3/temp5[105] , \MC_ARK_ARC_1_3/temp5[104] ,
         \MC_ARK_ARC_1_3/temp5[100] , \MC_ARK_ARC_1_3/temp5[99] ,
         \MC_ARK_ARC_1_3/temp5[98] , \MC_ARK_ARC_1_3/temp5[97] ,
         \MC_ARK_ARC_1_3/temp5[96] , \MC_ARK_ARC_1_3/temp5[93] ,
         \MC_ARK_ARC_1_3/temp5[92] , \MC_ARK_ARC_1_3/temp5[88] ,
         \MC_ARK_ARC_1_3/temp5[86] , \MC_ARK_ARC_1_3/temp5[85] ,
         \MC_ARK_ARC_1_3/temp5[84] , \MC_ARK_ARC_1_3/temp5[83] ,
         \MC_ARK_ARC_1_3/temp5[82] , \MC_ARK_ARC_1_3/temp5[80] ,
         \MC_ARK_ARC_1_3/temp5[76] , \MC_ARK_ARC_1_3/temp5[75] ,
         \MC_ARK_ARC_1_3/temp5[71] , \MC_ARK_ARC_1_3/temp5[70] ,
         \MC_ARK_ARC_1_3/temp5[69] , \MC_ARK_ARC_1_3/temp5[68] ,
         \MC_ARK_ARC_1_3/temp5[66] , \MC_ARK_ARC_1_3/temp5[64] ,
         \MC_ARK_ARC_1_3/temp5[61] , \MC_ARK_ARC_1_3/temp5[60] ,
         \MC_ARK_ARC_1_3/temp5[58] , \MC_ARK_ARC_1_3/temp5[53] ,
         \MC_ARK_ARC_1_3/temp5[51] , \MC_ARK_ARC_1_3/temp5[50] ,
         \MC_ARK_ARC_1_3/temp5[49] , \MC_ARK_ARC_1_3/temp5[48] ,
         \MC_ARK_ARC_1_3/temp5[46] , \MC_ARK_ARC_1_3/temp5[44] ,
         \MC_ARK_ARC_1_3/temp5[40] , \MC_ARK_ARC_1_3/temp5[39] ,
         \MC_ARK_ARC_1_3/temp5[35] , \MC_ARK_ARC_1_3/temp5[34] ,
         \MC_ARK_ARC_1_3/temp5[33] , \MC_ARK_ARC_1_3/temp5[30] ,
         \MC_ARK_ARC_1_3/temp5[29] , \MC_ARK_ARC_1_3/temp5[26] ,
         \MC_ARK_ARC_1_3/temp5[23] , \MC_ARK_ARC_1_3/temp5[21] ,
         \MC_ARK_ARC_1_3/temp5[16] , \MC_ARK_ARC_1_3/temp5[13] ,
         \MC_ARK_ARC_1_3/temp5[12] , \MC_ARK_ARC_1_3/temp5[9] ,
         \MC_ARK_ARC_1_3/temp5[8] , \MC_ARK_ARC_1_3/temp5[7] ,
         \MC_ARK_ARC_1_3/temp5[6] , \MC_ARK_ARC_1_3/temp5[5] ,
         \MC_ARK_ARC_1_3/temp5[4] , \MC_ARK_ARC_1_3/temp5[2] ,
         \MC_ARK_ARC_1_3/temp5[0] , \MC_ARK_ARC_1_3/temp4[190] ,
         \MC_ARK_ARC_1_3/temp4[188] , \MC_ARK_ARC_1_3/temp4[187] ,
         \MC_ARK_ARC_1_3/temp4[186] , \MC_ARK_ARC_1_3/temp4[185] ,
         \MC_ARK_ARC_1_3/temp4[184] , \MC_ARK_ARC_1_3/temp4[182] ,
         \MC_ARK_ARC_1_3/temp4[181] , \MC_ARK_ARC_1_3/temp4[180] ,
         \MC_ARK_ARC_1_3/temp4[179] , \MC_ARK_ARC_1_3/temp4[178] ,
         \MC_ARK_ARC_1_3/temp4[177] , \MC_ARK_ARC_1_3/temp4[175] ,
         \MC_ARK_ARC_1_3/temp4[174] , \MC_ARK_ARC_1_3/temp4[173] ,
         \MC_ARK_ARC_1_3/temp4[172] , \MC_ARK_ARC_1_3/temp4[171] ,
         \MC_ARK_ARC_1_3/temp4[169] , \MC_ARK_ARC_1_3/temp4[168] ,
         \MC_ARK_ARC_1_3/temp4[167] , \MC_ARK_ARC_1_3/temp4[165] ,
         \MC_ARK_ARC_1_3/temp4[164] , \MC_ARK_ARC_1_3/temp4[163] ,
         \MC_ARK_ARC_1_3/temp4[162] , \MC_ARK_ARC_1_3/temp4[161] ,
         \MC_ARK_ARC_1_3/temp4[160] , \MC_ARK_ARC_1_3/temp4[159] ,
         \MC_ARK_ARC_1_3/temp4[158] , \MC_ARK_ARC_1_3/temp4[157] ,
         \MC_ARK_ARC_1_3/temp4[156] , \MC_ARK_ARC_1_3/temp4[154] ,
         \MC_ARK_ARC_1_3/temp4[153] , \MC_ARK_ARC_1_3/temp4[152] ,
         \MC_ARK_ARC_1_3/temp4[151] , \MC_ARK_ARC_1_3/temp4[150] ,
         \MC_ARK_ARC_1_3/temp4[149] , \MC_ARK_ARC_1_3/temp4[147] ,
         \MC_ARK_ARC_1_3/temp4[146] , \MC_ARK_ARC_1_3/temp4[145] ,
         \MC_ARK_ARC_1_3/temp4[144] , \MC_ARK_ARC_1_3/temp4[143] ,
         \MC_ARK_ARC_1_3/temp4[142] , \MC_ARK_ARC_1_3/temp4[141] ,
         \MC_ARK_ARC_1_3/temp4[140] , \MC_ARK_ARC_1_3/temp4[139] ,
         \MC_ARK_ARC_1_3/temp4[138] , \MC_ARK_ARC_1_3/temp4[136] ,
         \MC_ARK_ARC_1_3/temp4[135] , \MC_ARK_ARC_1_3/temp4[134] ,
         \MC_ARK_ARC_1_3/temp4[133] , \MC_ARK_ARC_1_3/temp4[132] ,
         \MC_ARK_ARC_1_3/temp4[131] , \MC_ARK_ARC_1_3/temp4[130] ,
         \MC_ARK_ARC_1_3/temp4[129] , \MC_ARK_ARC_1_3/temp4[128] ,
         \MC_ARK_ARC_1_3/temp4[127] , \MC_ARK_ARC_1_3/temp4[126] ,
         \MC_ARK_ARC_1_3/temp4[125] , \MC_ARK_ARC_1_3/temp4[124] ,
         \MC_ARK_ARC_1_3/temp4[123] , \MC_ARK_ARC_1_3/temp4[122] ,
         \MC_ARK_ARC_1_3/temp4[121] , \MC_ARK_ARC_1_3/temp4[120] ,
         \MC_ARK_ARC_1_3/temp4[118] , \MC_ARK_ARC_1_3/temp4[117] ,
         \MC_ARK_ARC_1_3/temp4[116] , \MC_ARK_ARC_1_3/temp4[115] ,
         \MC_ARK_ARC_1_3/temp4[113] , \MC_ARK_ARC_1_3/temp4[112] ,
         \MC_ARK_ARC_1_3/temp4[111] , \MC_ARK_ARC_1_3/temp4[110] ,
         \MC_ARK_ARC_1_3/temp4[109] , \MC_ARK_ARC_1_3/temp4[108] ,
         \MC_ARK_ARC_1_3/temp4[107] , \MC_ARK_ARC_1_3/temp4[106] ,
         \MC_ARK_ARC_1_3/temp4[105] , \MC_ARK_ARC_1_3/temp4[103] ,
         \MC_ARK_ARC_1_3/temp4[102] , \MC_ARK_ARC_1_3/temp4[101] ,
         \MC_ARK_ARC_1_3/temp4[100] , \MC_ARK_ARC_1_3/temp4[99] ,
         \MC_ARK_ARC_1_3/temp4[98] , \MC_ARK_ARC_1_3/temp4[97] ,
         \MC_ARK_ARC_1_3/temp4[96] , \MC_ARK_ARC_1_3/temp4[95] ,
         \MC_ARK_ARC_1_3/temp4[94] , \MC_ARK_ARC_1_3/temp4[93] ,
         \MC_ARK_ARC_1_3/temp4[92] , \MC_ARK_ARC_1_3/temp4[91] ,
         \MC_ARK_ARC_1_3/temp4[90] , \MC_ARK_ARC_1_3/temp4[89] ,
         \MC_ARK_ARC_1_3/temp4[88] , \MC_ARK_ARC_1_3/temp4[87] ,
         \MC_ARK_ARC_1_3/temp4[86] , \MC_ARK_ARC_1_3/temp4[85] ,
         \MC_ARK_ARC_1_3/temp4[84] , \MC_ARK_ARC_1_3/temp4[82] ,
         \MC_ARK_ARC_1_3/temp4[80] , \MC_ARK_ARC_1_3/temp4[79] ,
         \MC_ARK_ARC_1_3/temp4[78] , \MC_ARK_ARC_1_3/temp4[77] ,
         \MC_ARK_ARC_1_3/temp4[76] , \MC_ARK_ARC_1_3/temp4[75] ,
         \MC_ARK_ARC_1_3/temp4[74] , \MC_ARK_ARC_1_3/temp4[73] ,
         \MC_ARK_ARC_1_3/temp4[72] , \MC_ARK_ARC_1_3/temp4[71] ,
         \MC_ARK_ARC_1_3/temp4[70] , \MC_ARK_ARC_1_3/temp4[69] ,
         \MC_ARK_ARC_1_3/temp4[68] , \MC_ARK_ARC_1_3/temp4[67] ,
         \MC_ARK_ARC_1_3/temp4[66] , \MC_ARK_ARC_1_3/temp4[65] ,
         \MC_ARK_ARC_1_3/temp4[64] , \MC_ARK_ARC_1_3/temp4[63] ,
         \MC_ARK_ARC_1_3/temp4[62] , \MC_ARK_ARC_1_3/temp4[61] ,
         \MC_ARK_ARC_1_3/temp4[60] , \MC_ARK_ARC_1_3/temp4[59] ,
         \MC_ARK_ARC_1_3/temp4[58] , \MC_ARK_ARC_1_3/temp4[57] ,
         \MC_ARK_ARC_1_3/temp4[55] , \MC_ARK_ARC_1_3/temp4[53] ,
         \MC_ARK_ARC_1_3/temp4[52] , \MC_ARK_ARC_1_3/temp4[51] ,
         \MC_ARK_ARC_1_3/temp4[50] , \MC_ARK_ARC_1_3/temp4[49] ,
         \MC_ARK_ARC_1_3/temp4[48] , \MC_ARK_ARC_1_3/temp4[46] ,
         \MC_ARK_ARC_1_3/temp4[45] , \MC_ARK_ARC_1_3/temp4[44] ,
         \MC_ARK_ARC_1_3/temp4[43] , \MC_ARK_ARC_1_3/temp4[42] ,
         \MC_ARK_ARC_1_3/temp4[41] , \MC_ARK_ARC_1_3/temp4[40] ,
         \MC_ARK_ARC_1_3/temp4[39] , \MC_ARK_ARC_1_3/temp4[37] ,
         \MC_ARK_ARC_1_3/temp4[36] , \MC_ARK_ARC_1_3/temp4[34] ,
         \MC_ARK_ARC_1_3/temp4[33] , \MC_ARK_ARC_1_3/temp4[32] ,
         \MC_ARK_ARC_1_3/temp4[31] , \MC_ARK_ARC_1_3/temp4[30] ,
         \MC_ARK_ARC_1_3/temp4[29] , \MC_ARK_ARC_1_3/temp4[28] ,
         \MC_ARK_ARC_1_3/temp4[27] , \MC_ARK_ARC_1_3/temp4[26] ,
         \MC_ARK_ARC_1_3/temp4[25] , \MC_ARK_ARC_1_3/temp4[24] ,
         \MC_ARK_ARC_1_3/temp4[22] , \MC_ARK_ARC_1_3/temp4[21] ,
         \MC_ARK_ARC_1_3/temp4[20] , \MC_ARK_ARC_1_3/temp4[19] ,
         \MC_ARK_ARC_1_3/temp4[18] , \MC_ARK_ARC_1_3/temp4[17] ,
         \MC_ARK_ARC_1_3/temp4[16] , \MC_ARK_ARC_1_3/temp4[14] ,
         \MC_ARK_ARC_1_3/temp4[13] , \MC_ARK_ARC_1_3/temp4[12] ,
         \MC_ARK_ARC_1_3/temp4[11] , \MC_ARK_ARC_1_3/temp4[10] ,
         \MC_ARK_ARC_1_3/temp4[9] , \MC_ARK_ARC_1_3/temp4[8] ,
         \MC_ARK_ARC_1_3/temp4[7] , \MC_ARK_ARC_1_3/temp4[6] ,
         \MC_ARK_ARC_1_3/temp4[4] , \MC_ARK_ARC_1_3/temp4[3] ,
         \MC_ARK_ARC_1_3/temp4[2] , \MC_ARK_ARC_1_3/temp4[1] ,
         \MC_ARK_ARC_1_3/temp4[0] , \MC_ARK_ARC_1_3/temp3[190] ,
         \MC_ARK_ARC_1_3/temp3[187] , \MC_ARK_ARC_1_3/temp3[186] ,
         \MC_ARK_ARC_1_3/temp3[184] , \MC_ARK_ARC_1_3/temp3[182] ,
         \MC_ARK_ARC_1_3/temp3[181] , \MC_ARK_ARC_1_3/temp3[180] ,
         \MC_ARK_ARC_1_3/temp3[179] , \MC_ARK_ARC_1_3/temp3[178] ,
         \MC_ARK_ARC_1_3/temp3[173] , \MC_ARK_ARC_1_3/temp3[172] ,
         \MC_ARK_ARC_1_3/temp3[171] , \MC_ARK_ARC_1_3/temp3[169] ,
         \MC_ARK_ARC_1_3/temp3[168] , \MC_ARK_ARC_1_3/temp3[165] ,
         \MC_ARK_ARC_1_3/temp3[164] , \MC_ARK_ARC_1_3/temp3[163] ,
         \MC_ARK_ARC_1_3/temp3[162] , \MC_ARK_ARC_1_3/temp3[161] ,
         \MC_ARK_ARC_1_3/temp3[160] , \MC_ARK_ARC_1_3/temp3[159] ,
         \MC_ARK_ARC_1_3/temp3[158] , \MC_ARK_ARC_1_3/temp3[157] ,
         \MC_ARK_ARC_1_3/temp3[156] , \MC_ARK_ARC_1_3/temp3[154] ,
         \MC_ARK_ARC_1_3/temp3[151] , \MC_ARK_ARC_1_3/temp3[149] ,
         \MC_ARK_ARC_1_3/temp3[147] , \MC_ARK_ARC_1_3/temp3[146] ,
         \MC_ARK_ARC_1_3/temp3[145] , \MC_ARK_ARC_1_3/temp3[144] ,
         \MC_ARK_ARC_1_3/temp3[143] , \MC_ARK_ARC_1_3/temp3[142] ,
         \MC_ARK_ARC_1_3/temp3[140] , \MC_ARK_ARC_1_3/temp3[139] ,
         \MC_ARK_ARC_1_3/temp3[138] , \MC_ARK_ARC_1_3/temp3[136] ,
         \MC_ARK_ARC_1_3/temp3[133] , \MC_ARK_ARC_1_3/temp3[130] ,
         \MC_ARK_ARC_1_3/temp3[129] , \MC_ARK_ARC_1_3/temp3[128] ,
         \MC_ARK_ARC_1_3/temp3[127] , \MC_ARK_ARC_1_3/temp3[126] ,
         \MC_ARK_ARC_1_3/temp3[125] , \MC_ARK_ARC_1_3/temp3[123] ,
         \MC_ARK_ARC_1_3/temp3[122] , \MC_ARK_ARC_1_3/temp3[121] ,
         \MC_ARK_ARC_1_3/temp3[120] , \MC_ARK_ARC_1_3/temp3[118] ,
         \MC_ARK_ARC_1_3/temp3[116] , \MC_ARK_ARC_1_3/temp3[115] ,
         \MC_ARK_ARC_1_3/temp3[113] , \MC_ARK_ARC_1_3/temp3[112] ,
         \MC_ARK_ARC_1_3/temp3[111] , \MC_ARK_ARC_1_3/temp3[110] ,
         \MC_ARK_ARC_1_3/temp3[109] , \MC_ARK_ARC_1_3/temp3[108] ,
         \MC_ARK_ARC_1_3/temp3[105] , \MC_ARK_ARC_1_3/temp3[101] ,
         \MC_ARK_ARC_1_3/temp3[97] , \MC_ARK_ARC_1_3/temp3[96] ,
         \MC_ARK_ARC_1_3/temp3[94] , \MC_ARK_ARC_1_3/temp3[93] ,
         \MC_ARK_ARC_1_3/temp3[91] , \MC_ARK_ARC_1_3/temp3[90] ,
         \MC_ARK_ARC_1_3/temp3[89] , \MC_ARK_ARC_1_3/temp3[88] ,
         \MC_ARK_ARC_1_3/temp3[87] , \MC_ARK_ARC_1_3/temp3[86] ,
         \MC_ARK_ARC_1_3/temp3[85] , \MC_ARK_ARC_1_3/temp3[84] ,
         \MC_ARK_ARC_1_3/temp3[82] , \MC_ARK_ARC_1_3/temp3[80] ,
         \MC_ARK_ARC_1_3/temp3[79] , \MC_ARK_ARC_1_3/temp3[78] ,
         \MC_ARK_ARC_1_3/temp3[76] , \MC_ARK_ARC_1_3/temp3[75] ,
         \MC_ARK_ARC_1_3/temp3[73] , \MC_ARK_ARC_1_3/temp3[72] ,
         \MC_ARK_ARC_1_3/temp3[70] , \MC_ARK_ARC_1_3/temp3[69] ,
         \MC_ARK_ARC_1_3/temp3[68] , \MC_ARK_ARC_1_3/temp3[67] ,
         \MC_ARK_ARC_1_3/temp3[66] , \MC_ARK_ARC_1_3/temp3[65] ,
         \MC_ARK_ARC_1_3/temp3[64] , \MC_ARK_ARC_1_3/temp3[63] ,
         \MC_ARK_ARC_1_3/temp3[61] , \MC_ARK_ARC_1_3/temp3[60] ,
         \MC_ARK_ARC_1_3/temp3[58] , \MC_ARK_ARC_1_3/temp3[57] ,
         \MC_ARK_ARC_1_3/temp3[55] , \MC_ARK_ARC_1_3/temp3[53] ,
         \MC_ARK_ARC_1_3/temp3[52] , \MC_ARK_ARC_1_3/temp3[51] ,
         \MC_ARK_ARC_1_3/temp3[49] , \MC_ARK_ARC_1_3/temp3[48] ,
         \MC_ARK_ARC_1_3/temp3[47] , \MC_ARK_ARC_1_3/temp3[46] ,
         \MC_ARK_ARC_1_3/temp3[42] , \MC_ARK_ARC_1_3/temp3[40] ,
         \MC_ARK_ARC_1_3/temp3[39] , \MC_ARK_ARC_1_3/temp3[37] ,
         \MC_ARK_ARC_1_3/temp3[36] , \MC_ARK_ARC_1_3/temp3[34] ,
         \MC_ARK_ARC_1_3/temp3[32] , \MC_ARK_ARC_1_3/temp3[30] ,
         \MC_ARK_ARC_1_3/temp3[29] , \MC_ARK_ARC_1_3/temp3[28] ,
         \MC_ARK_ARC_1_3/temp3[27] , \MC_ARK_ARC_1_3/temp3[25] ,
         \MC_ARK_ARC_1_3/temp3[22] , \MC_ARK_ARC_1_3/temp3[21] ,
         \MC_ARK_ARC_1_3/temp3[18] , \MC_ARK_ARC_1_3/temp3[16] ,
         \MC_ARK_ARC_1_3/temp3[14] , \MC_ARK_ARC_1_3/temp3[12] ,
         \MC_ARK_ARC_1_3/temp3[11] , \MC_ARK_ARC_1_3/temp3[9] ,
         \MC_ARK_ARC_1_3/temp3[7] , \MC_ARK_ARC_1_3/temp3[6] ,
         \MC_ARK_ARC_1_3/temp3[4] , \MC_ARK_ARC_1_3/temp3[3] ,
         \MC_ARK_ARC_1_3/temp3[1] , \MC_ARK_ARC_1_3/temp3[0] ,
         \MC_ARK_ARC_1_3/temp2[190] , \MC_ARK_ARC_1_3/temp2[188] ,
         \MC_ARK_ARC_1_3/temp2[186] , \MC_ARK_ARC_1_3/temp2[179] ,
         \MC_ARK_ARC_1_3/temp2[178] , \MC_ARK_ARC_1_3/temp2[177] ,
         \MC_ARK_ARC_1_3/temp2[176] , \MC_ARK_ARC_1_3/temp2[175] ,
         \MC_ARK_ARC_1_3/temp2[173] , \MC_ARK_ARC_1_3/temp2[172] ,
         \MC_ARK_ARC_1_3/temp2[171] , \MC_ARK_ARC_1_3/temp2[169] ,
         \MC_ARK_ARC_1_3/temp2[168] , \MC_ARK_ARC_1_3/temp2[167] ,
         \MC_ARK_ARC_1_3/temp2[166] , \MC_ARK_ARC_1_3/temp2[165] ,
         \MC_ARK_ARC_1_3/temp2[161] , \MC_ARK_ARC_1_3/temp2[160] ,
         \MC_ARK_ARC_1_3/temp2[159] , \MC_ARK_ARC_1_3/temp2[157] ,
         \MC_ARK_ARC_1_3/temp2[156] , \MC_ARK_ARC_1_3/temp2[155] ,
         \MC_ARK_ARC_1_3/temp2[154] , \MC_ARK_ARC_1_3/temp2[152] ,
         \MC_ARK_ARC_1_3/temp2[150] , \MC_ARK_ARC_1_3/temp2[149] ,
         \MC_ARK_ARC_1_3/temp2[148] , \MC_ARK_ARC_1_3/temp2[144] ,
         \MC_ARK_ARC_1_3/temp2[142] , \MC_ARK_ARC_1_3/temp2[141] ,
         \MC_ARK_ARC_1_3/temp2[140] , \MC_ARK_ARC_1_3/temp2[139] ,
         \MC_ARK_ARC_1_3/temp2[135] , \MC_ARK_ARC_1_3/temp2[134] ,
         \MC_ARK_ARC_1_3/temp2[133] , \MC_ARK_ARC_1_3/temp2[132] ,
         \MC_ARK_ARC_1_3/temp2[130] , \MC_ARK_ARC_1_3/temp2[128] ,
         \MC_ARK_ARC_1_3/temp2[127] , \MC_ARK_ARC_1_3/temp2[126] ,
         \MC_ARK_ARC_1_3/temp2[125] , \MC_ARK_ARC_1_3/temp2[124] ,
         \MC_ARK_ARC_1_3/temp2[123] , \MC_ARK_ARC_1_3/temp2[122] ,
         \MC_ARK_ARC_1_3/temp2[121] , \MC_ARK_ARC_1_3/temp2[120] ,
         \MC_ARK_ARC_1_3/temp2[116] , \MC_ARK_ARC_1_3/temp2[114] ,
         \MC_ARK_ARC_1_3/temp2[113] , \MC_ARK_ARC_1_3/temp2[112] ,
         \MC_ARK_ARC_1_3/temp2[111] , \MC_ARK_ARC_1_3/temp2[110] ,
         \MC_ARK_ARC_1_3/temp2[109] , \MC_ARK_ARC_1_3/temp2[108] ,
         \MC_ARK_ARC_1_3/temp2[106] , \MC_ARK_ARC_1_3/temp2[105] ,
         \MC_ARK_ARC_1_3/temp2[104] , \MC_ARK_ARC_1_3/temp2[103] ,
         \MC_ARK_ARC_1_3/temp2[102] , \MC_ARK_ARC_1_3/temp2[101] ,
         \MC_ARK_ARC_1_3/temp2[99] , \MC_ARK_ARC_1_3/temp2[98] ,
         \MC_ARK_ARC_1_3/temp2[96] , \MC_ARK_ARC_1_3/temp2[94] ,
         \MC_ARK_ARC_1_3/temp2[93] , \MC_ARK_ARC_1_3/temp2[91] ,
         \MC_ARK_ARC_1_3/temp2[90] , \MC_ARK_ARC_1_3/temp2[88] ,
         \MC_ARK_ARC_1_3/temp2[87] , \MC_ARK_ARC_1_3/temp2[84] ,
         \MC_ARK_ARC_1_3/temp2[83] , \MC_ARK_ARC_1_3/temp2[82] ,
         \MC_ARK_ARC_1_3/temp2[78] , \MC_ARK_ARC_1_3/temp2[76] ,
         \MC_ARK_ARC_1_3/temp2[72] , \MC_ARK_ARC_1_3/temp2[71] ,
         \MC_ARK_ARC_1_3/temp2[70] , \MC_ARK_ARC_1_3/temp2[68] ,
         \MC_ARK_ARC_1_3/temp2[67] , \MC_ARK_ARC_1_3/temp2[66] ,
         \MC_ARK_ARC_1_3/temp2[65] , \MC_ARK_ARC_1_3/temp2[64] ,
         \MC_ARK_ARC_1_3/temp2[62] , \MC_ARK_ARC_1_3/temp2[61] ,
         \MC_ARK_ARC_1_3/temp2[58] , \MC_ARK_ARC_1_3/temp2[57] ,
         \MC_ARK_ARC_1_3/temp2[56] , \MC_ARK_ARC_1_3/temp2[55] ,
         \MC_ARK_ARC_1_3/temp2[54] , \MC_ARK_ARC_1_3/temp2[53] ,
         \MC_ARK_ARC_1_3/temp2[52] , \MC_ARK_ARC_1_3/temp2[50] ,
         \MC_ARK_ARC_1_3/temp2[49] , \MC_ARK_ARC_1_3/temp2[48] ,
         \MC_ARK_ARC_1_3/temp2[47] , \MC_ARK_ARC_1_3/temp2[46] ,
         \MC_ARK_ARC_1_3/temp2[43] , \MC_ARK_ARC_1_3/temp2[40] ,
         \MC_ARK_ARC_1_3/temp2[38] , \MC_ARK_ARC_1_3/temp2[36] ,
         \MC_ARK_ARC_1_3/temp2[34] , \MC_ARK_ARC_1_3/temp2[33] ,
         \MC_ARK_ARC_1_3/temp2[32] , \MC_ARK_ARC_1_3/temp2[30] ,
         \MC_ARK_ARC_1_3/temp2[25] , \MC_ARK_ARC_1_3/temp2[20] ,
         \MC_ARK_ARC_1_3/temp2[19] , \MC_ARK_ARC_1_3/temp2[18] ,
         \MC_ARK_ARC_1_3/temp2[17] , \MC_ARK_ARC_1_3/temp2[16] ,
         \MC_ARK_ARC_1_3/temp2[14] , \MC_ARK_ARC_1_3/temp2[13] ,
         \MC_ARK_ARC_1_3/temp2[12] , \MC_ARK_ARC_1_3/temp2[10] ,
         \MC_ARK_ARC_1_3/temp2[8] , \MC_ARK_ARC_1_3/temp2[6] ,
         \MC_ARK_ARC_1_3/temp2[5] , \MC_ARK_ARC_1_3/temp2[4] ,
         \MC_ARK_ARC_1_3/temp2[2] , \MC_ARK_ARC_1_3/temp2[1] ,
         \MC_ARK_ARC_1_3/temp2[0] , \MC_ARK_ARC_1_3/temp1[190] ,
         \MC_ARK_ARC_1_3/temp1[189] , \MC_ARK_ARC_1_3/temp1[188] ,
         \MC_ARK_ARC_1_3/temp1[187] , \MC_ARK_ARC_1_3/temp1[186] ,
         \MC_ARK_ARC_1_3/temp1[185] , \MC_ARK_ARC_1_3/temp1[184] ,
         \MC_ARK_ARC_1_3/temp1[181] , \MC_ARK_ARC_1_3/temp1[180] ,
         \MC_ARK_ARC_1_3/temp1[179] , \MC_ARK_ARC_1_3/temp1[178] ,
         \MC_ARK_ARC_1_3/temp1[177] , \MC_ARK_ARC_1_3/temp1[176] ,
         \MC_ARK_ARC_1_3/temp1[175] , \MC_ARK_ARC_1_3/temp1[174] ,
         \MC_ARK_ARC_1_3/temp1[173] , \MC_ARK_ARC_1_3/temp1[169] ,
         \MC_ARK_ARC_1_3/temp1[168] , \MC_ARK_ARC_1_3/temp1[167] ,
         \MC_ARK_ARC_1_3/temp1[166] , \MC_ARK_ARC_1_3/temp1[163] ,
         \MC_ARK_ARC_1_3/temp1[162] , \MC_ARK_ARC_1_3/temp1[161] ,
         \MC_ARK_ARC_1_3/temp1[160] , \MC_ARK_ARC_1_3/temp1[159] ,
         \MC_ARK_ARC_1_3/temp1[158] , \MC_ARK_ARC_1_3/temp1[157] ,
         \MC_ARK_ARC_1_3/temp1[156] , \MC_ARK_ARC_1_3/temp1[151] ,
         \MC_ARK_ARC_1_3/temp1[146] , \MC_ARK_ARC_1_3/temp1[145] ,
         \MC_ARK_ARC_1_3/temp1[144] , \MC_ARK_ARC_1_3/temp1[142] ,
         \MC_ARK_ARC_1_3/temp1[140] , \MC_ARK_ARC_1_3/temp1[139] ,
         \MC_ARK_ARC_1_3/temp1[136] , \MC_ARK_ARC_1_3/temp1[135] ,
         \MC_ARK_ARC_1_3/temp1[134] , \MC_ARK_ARC_1_3/temp1[133] ,
         \MC_ARK_ARC_1_3/temp1[130] , \MC_ARK_ARC_1_3/temp1[128] ,
         \MC_ARK_ARC_1_3/temp1[127] , \MC_ARK_ARC_1_3/temp1[126] ,
         \MC_ARK_ARC_1_3/temp1[125] , \MC_ARK_ARC_1_3/temp1[124] ,
         \MC_ARK_ARC_1_3/temp1[123] , \MC_ARK_ARC_1_3/temp1[121] ,
         \MC_ARK_ARC_1_3/temp1[119] , \MC_ARK_ARC_1_3/temp1[118] ,
         \MC_ARK_ARC_1_3/temp1[117] , \MC_ARK_ARC_1_3/temp1[116] ,
         \MC_ARK_ARC_1_3/temp1[115] , \MC_ARK_ARC_1_3/temp1[113] ,
         \MC_ARK_ARC_1_3/temp1[111] , \MC_ARK_ARC_1_3/temp1[109] ,
         \MC_ARK_ARC_1_3/temp1[108] , \MC_ARK_ARC_1_3/temp1[106] ,
         \MC_ARK_ARC_1_3/temp1[103] , \MC_ARK_ARC_1_3/temp1[102] ,
         \MC_ARK_ARC_1_3/temp1[101] , \MC_ARK_ARC_1_3/temp1[98] ,
         \MC_ARK_ARC_1_3/temp1[96] , \MC_ARK_ARC_1_3/temp1[92] ,
         \MC_ARK_ARC_1_3/temp1[90] , \MC_ARK_ARC_1_3/temp1[89] ,
         \MC_ARK_ARC_1_3/temp1[88] , \MC_ARK_ARC_1_3/temp1[87] ,
         \MC_ARK_ARC_1_3/temp1[86] , \MC_ARK_ARC_1_3/temp1[85] ,
         \MC_ARK_ARC_1_3/temp1[84] , \MC_ARK_ARC_1_3/temp1[83] ,
         \MC_ARK_ARC_1_3/temp1[82] , \MC_ARK_ARC_1_3/temp1[80] ,
         \MC_ARK_ARC_1_3/temp1[78] , \MC_ARK_ARC_1_3/temp1[77] ,
         \MC_ARK_ARC_1_3/temp1[76] , \MC_ARK_ARC_1_3/temp1[75] ,
         \MC_ARK_ARC_1_3/temp1[74] , \MC_ARK_ARC_1_3/temp1[72] ,
         \MC_ARK_ARC_1_3/temp1[69] , \MC_ARK_ARC_1_3/temp1[68] ,
         \MC_ARK_ARC_1_3/temp1[67] , \MC_ARK_ARC_1_3/temp1[66] ,
         \MC_ARK_ARC_1_3/temp1[65] , \MC_ARK_ARC_1_3/temp1[64] ,
         \MC_ARK_ARC_1_3/temp1[62] , \MC_ARK_ARC_1_3/temp1[61] ,
         \MC_ARK_ARC_1_3/temp1[60] , \MC_ARK_ARC_1_3/temp1[58] ,
         \MC_ARK_ARC_1_3/temp1[55] , \MC_ARK_ARC_1_3/temp1[54] ,
         \MC_ARK_ARC_1_3/temp1[53] , \MC_ARK_ARC_1_3/temp1[52] ,
         \MC_ARK_ARC_1_3/temp1[51] , \MC_ARK_ARC_1_3/temp1[49] ,
         \MC_ARK_ARC_1_3/temp1[48] , \MC_ARK_ARC_1_3/temp1[46] ,
         \MC_ARK_ARC_1_3/temp1[44] , \MC_ARK_ARC_1_3/temp1[43] ,
         \MC_ARK_ARC_1_3/temp1[42] , \MC_ARK_ARC_1_3/temp1[40] ,
         \MC_ARK_ARC_1_3/temp1[35] , \MC_ARK_ARC_1_3/temp1[34] ,
         \MC_ARK_ARC_1_3/temp1[32] , \MC_ARK_ARC_1_3/temp1[31] ,
         \MC_ARK_ARC_1_3/temp1[30] , \MC_ARK_ARC_1_3/temp1[28] ,
         \MC_ARK_ARC_1_3/temp1[27] , \MC_ARK_ARC_1_3/temp1[26] ,
         \MC_ARK_ARC_1_3/temp1[24] , \MC_ARK_ARC_1_3/temp1[21] ,
         \MC_ARK_ARC_1_3/temp1[16] , \MC_ARK_ARC_1_3/temp1[14] ,
         \MC_ARK_ARC_1_3/temp1[12] , \MC_ARK_ARC_1_3/temp1[10] ,
         \MC_ARK_ARC_1_3/temp1[9] , \MC_ARK_ARC_1_3/temp1[8] ,
         \MC_ARK_ARC_1_3/temp1[6] , \MC_ARK_ARC_1_3/temp1[4] ,
         \MC_ARK_ARC_1_3/temp1[3] , \MC_ARK_ARC_1_3/temp1[2] ,
         \MC_ARK_ARC_1_3/temp1[1] , \MC_ARK_ARC_1_3/temp1[0] ,
         \MC_ARK_ARC_1_3/buf_keyinput[183] ,
         \MC_ARK_ARC_1_3/buf_keyinput[132] ,
         \MC_ARK_ARC_1_3/buf_datainput[187] ,
         \MC_ARK_ARC_1_3/buf_datainput[184] ,
         \MC_ARK_ARC_1_3/buf_datainput[183] ,
         \MC_ARK_ARC_1_3/buf_datainput[182] ,
         \MC_ARK_ARC_1_3/buf_datainput[178] ,
         \MC_ARK_ARC_1_3/buf_datainput[177] ,
         \MC_ARK_ARC_1_3/buf_datainput[176] ,
         \MC_ARK_ARC_1_3/buf_datainput[170] ,
         \MC_ARK_ARC_1_3/buf_datainput[164] ,
         \MC_ARK_ARC_1_3/buf_datainput[159] ,
         \MC_ARK_ARC_1_3/buf_datainput[158] ,
         \MC_ARK_ARC_1_3/buf_datainput[157] ,
         \MC_ARK_ARC_1_3/buf_datainput[156] ,
         \MC_ARK_ARC_1_3/buf_datainput[155] ,
         \MC_ARK_ARC_1_3/buf_datainput[151] ,
         \MC_ARK_ARC_1_3/buf_datainput[147] ,
         \MC_ARK_ARC_1_3/buf_datainput[144] ,
         \MC_ARK_ARC_1_3/buf_datainput[143] ,
         \MC_ARK_ARC_1_3/buf_datainput[142] ,
         \MC_ARK_ARC_1_3/buf_datainput[141] ,
         \MC_ARK_ARC_1_3/buf_datainput[140] ,
         \MC_ARK_ARC_1_3/buf_datainput[133] ,
         \MC_ARK_ARC_1_3/buf_datainput[129] ,
         \MC_ARK_ARC_1_3/buf_datainput[128] ,
         \MC_ARK_ARC_1_3/buf_datainput[118] ,
         \MC_ARK_ARC_1_3/buf_datainput[116] ,
         \MC_ARK_ARC_1_3/buf_datainput[115] ,
         \MC_ARK_ARC_1_3/buf_datainput[109] ,
         \MC_ARK_ARC_1_3/buf_datainput[105] ,
         \MC_ARK_ARC_1_3/buf_datainput[102] ,
         \MC_ARK_ARC_1_3/buf_datainput[99] ,
         \MC_ARK_ARC_1_3/buf_datainput[96] ,
         \MC_ARK_ARC_1_3/buf_datainput[94] ,
         \MC_ARK_ARC_1_3/buf_datainput[80] ,
         \MC_ARK_ARC_1_3/buf_datainput[71] ,
         \MC_ARK_ARC_1_3/buf_datainput[69] ,
         \MC_ARK_ARC_1_3/buf_datainput[62] ,
         \MC_ARK_ARC_1_3/buf_datainput[53] ,
         \MC_ARK_ARC_1_3/buf_datainput[49] ,
         \MC_ARK_ARC_1_3/buf_datainput[46] ,
         \MC_ARK_ARC_1_3/buf_datainput[43] ,
         \MC_ARK_ARC_1_3/buf_datainput[39] ,
         \MC_ARK_ARC_1_3/buf_datainput[37] ,
         \MC_ARK_ARC_1_3/buf_datainput[32] ,
         \MC_ARK_ARC_1_3/buf_datainput[29] ,
         \MC_ARK_ARC_1_3/buf_datainput[24] ,
         \MC_ARK_ARC_1_3/buf_datainput[21] ,
         \MC_ARK_ARC_1_3/buf_datainput[20] ,
         \MC_ARK_ARC_1_3/buf_datainput[19] ,
         \MC_ARK_ARC_1_3/buf_datainput[15] , \MC_ARK_ARC_1_3/buf_datainput[7] ,
         \MC_ARK_ARC_1_3/buf_datainput[5] , \MC_ARK_ARC_1_3/buf_datainput[1] ,
         \MC_ARK_ARC_1_3/buf_datainput[0] , \MC_ARK_ARC_1_4/buf_output[191] ,
         \MC_ARK_ARC_1_4/buf_output[190] , \MC_ARK_ARC_1_4/buf_output[189] ,
         \MC_ARK_ARC_1_4/buf_output[188] , \MC_ARK_ARC_1_4/buf_output[187] ,
         \MC_ARK_ARC_1_4/buf_output[186] , \MC_ARK_ARC_1_4/buf_output[184] ,
         \MC_ARK_ARC_1_4/buf_output[183] , \MC_ARK_ARC_1_4/buf_output[182] ,
         \MC_ARK_ARC_1_4/buf_output[181] , \MC_ARK_ARC_1_4/buf_output[180] ,
         \MC_ARK_ARC_1_4/buf_output[178] , \MC_ARK_ARC_1_4/buf_output[177] ,
         \MC_ARK_ARC_1_4/buf_output[176] , \MC_ARK_ARC_1_4/buf_output[175] ,
         \MC_ARK_ARC_1_4/buf_output[174] , \MC_ARK_ARC_1_4/buf_output[172] ,
         \MC_ARK_ARC_1_4/buf_output[171] , \MC_ARK_ARC_1_4/buf_output[170] ,
         \MC_ARK_ARC_1_4/buf_output[169] , \MC_ARK_ARC_1_4/buf_output[168] ,
         \MC_ARK_ARC_1_4/buf_output[166] , \MC_ARK_ARC_1_4/buf_output[165] ,
         \MC_ARK_ARC_1_4/buf_output[164] , \MC_ARK_ARC_1_4/buf_output[163] ,
         \MC_ARK_ARC_1_4/buf_output[162] , \MC_ARK_ARC_1_4/buf_output[160] ,
         \MC_ARK_ARC_1_4/buf_output[159] , \MC_ARK_ARC_1_4/buf_output[158] ,
         \MC_ARK_ARC_1_4/buf_output[157] , \MC_ARK_ARC_1_4/buf_output[156] ,
         \MC_ARK_ARC_1_4/buf_output[154] , \MC_ARK_ARC_1_4/buf_output[153] ,
         \MC_ARK_ARC_1_4/buf_output[152] , \MC_ARK_ARC_1_4/buf_output[151] ,
         \MC_ARK_ARC_1_4/buf_output[150] , \MC_ARK_ARC_1_4/buf_output[148] ,
         \MC_ARK_ARC_1_4/buf_output[147] , \MC_ARK_ARC_1_4/buf_output[146] ,
         \MC_ARK_ARC_1_4/buf_output[145] , \MC_ARK_ARC_1_4/buf_output[144] ,
         \MC_ARK_ARC_1_4/buf_output[143] , \MC_ARK_ARC_1_4/buf_output[142] ,
         \MC_ARK_ARC_1_4/buf_output[141] , \MC_ARK_ARC_1_4/buf_output[140] ,
         \MC_ARK_ARC_1_4/buf_output[139] , \MC_ARK_ARC_1_4/buf_output[138] ,
         \MC_ARK_ARC_1_4/buf_output[136] , \MC_ARK_ARC_1_4/buf_output[135] ,
         \MC_ARK_ARC_1_4/buf_output[134] , \MC_ARK_ARC_1_4/buf_output[133] ,
         \MC_ARK_ARC_1_4/buf_output[132] , \MC_ARK_ARC_1_4/buf_output[131] ,
         \MC_ARK_ARC_1_4/buf_output[130] , \MC_ARK_ARC_1_4/buf_output[129] ,
         \MC_ARK_ARC_1_4/buf_output[128] , \MC_ARK_ARC_1_4/buf_output[127] ,
         \MC_ARK_ARC_1_4/buf_output[126] , \MC_ARK_ARC_1_4/buf_output[124] ,
         \MC_ARK_ARC_1_4/buf_output[123] , \MC_ARK_ARC_1_4/buf_output[122] ,
         \MC_ARK_ARC_1_4/buf_output[121] , \MC_ARK_ARC_1_4/buf_output[120] ,
         \MC_ARK_ARC_1_4/buf_output[119] , \MC_ARK_ARC_1_4/buf_output[118] ,
         \MC_ARK_ARC_1_4/buf_output[117] , \MC_ARK_ARC_1_4/buf_output[116] ,
         \MC_ARK_ARC_1_4/buf_output[115] , \MC_ARK_ARC_1_4/buf_output[114] ,
         \MC_ARK_ARC_1_4/buf_output[113] , \MC_ARK_ARC_1_4/buf_output[112] ,
         \MC_ARK_ARC_1_4/buf_output[111] , \MC_ARK_ARC_1_4/buf_output[110] ,
         \MC_ARK_ARC_1_4/buf_output[109] , \MC_ARK_ARC_1_4/buf_output[108] ,
         \MC_ARK_ARC_1_4/buf_output[106] , \MC_ARK_ARC_1_4/buf_output[105] ,
         \MC_ARK_ARC_1_4/buf_output[104] , \MC_ARK_ARC_1_4/buf_output[103] ,
         \MC_ARK_ARC_1_4/buf_output[102] , \MC_ARK_ARC_1_4/buf_output[101] ,
         \MC_ARK_ARC_1_4/buf_output[100] , \MC_ARK_ARC_1_4/buf_output[99] ,
         \MC_ARK_ARC_1_4/buf_output[98] , \MC_ARK_ARC_1_4/buf_output[97] ,
         \MC_ARK_ARC_1_4/buf_output[96] , \MC_ARK_ARC_1_4/buf_output[95] ,
         \MC_ARK_ARC_1_4/buf_output[94] , \MC_ARK_ARC_1_4/buf_output[93] ,
         \MC_ARK_ARC_1_4/buf_output[92] , \MC_ARK_ARC_1_4/buf_output[91] ,
         \MC_ARK_ARC_1_4/buf_output[90] , \MC_ARK_ARC_1_4/buf_output[88] ,
         \MC_ARK_ARC_1_4/buf_output[87] , \MC_ARK_ARC_1_4/buf_output[86] ,
         \MC_ARK_ARC_1_4/buf_output[85] , \MC_ARK_ARC_1_4/buf_output[84] ,
         \MC_ARK_ARC_1_4/buf_output[83] , \MC_ARK_ARC_1_4/buf_output[82] ,
         \MC_ARK_ARC_1_4/buf_output[81] , \MC_ARK_ARC_1_4/buf_output[79] ,
         \MC_ARK_ARC_1_4/buf_output[78] , \MC_ARK_ARC_1_4/buf_output[76] ,
         \MC_ARK_ARC_1_4/buf_output[75] , \MC_ARK_ARC_1_4/buf_output[74] ,
         \MC_ARK_ARC_1_4/buf_output[73] , \MC_ARK_ARC_1_4/buf_output[72] ,
         \MC_ARK_ARC_1_4/buf_output[71] , \MC_ARK_ARC_1_4/buf_output[70] ,
         \MC_ARK_ARC_1_4/buf_output[69] , \MC_ARK_ARC_1_4/buf_output[68] ,
         \MC_ARK_ARC_1_4/buf_output[67] , \MC_ARK_ARC_1_4/buf_output[66] ,
         \MC_ARK_ARC_1_4/buf_output[65] , \MC_ARK_ARC_1_4/buf_output[64] ,
         \MC_ARK_ARC_1_4/buf_output[63] , \MC_ARK_ARC_1_4/buf_output[62] ,
         \MC_ARK_ARC_1_4/buf_output[61] , \MC_ARK_ARC_1_4/buf_output[60] ,
         \MC_ARK_ARC_1_4/buf_output[58] , \MC_ARK_ARC_1_4/buf_output[57] ,
         \MC_ARK_ARC_1_4/buf_output[56] , \MC_ARK_ARC_1_4/buf_output[55] ,
         \MC_ARK_ARC_1_4/buf_output[54] , \MC_ARK_ARC_1_4/buf_output[52] ,
         \MC_ARK_ARC_1_4/buf_output[51] , \MC_ARK_ARC_1_4/buf_output[50] ,
         \MC_ARK_ARC_1_4/buf_output[49] , \MC_ARK_ARC_1_4/buf_output[48] ,
         \MC_ARK_ARC_1_4/buf_output[46] , \MC_ARK_ARC_1_4/buf_output[45] ,
         \MC_ARK_ARC_1_4/buf_output[44] , \MC_ARK_ARC_1_4/buf_output[43] ,
         \MC_ARK_ARC_1_4/buf_output[42] , \MC_ARK_ARC_1_4/buf_output[40] ,
         \MC_ARK_ARC_1_4/buf_output[39] , \MC_ARK_ARC_1_4/buf_output[38] ,
         \MC_ARK_ARC_1_4/buf_output[37] , \MC_ARK_ARC_1_4/buf_output[36] ,
         \MC_ARK_ARC_1_4/buf_output[34] , \MC_ARK_ARC_1_4/buf_output[33] ,
         \MC_ARK_ARC_1_4/buf_output[32] , \MC_ARK_ARC_1_4/buf_output[31] ,
         \MC_ARK_ARC_1_4/buf_output[30] , \MC_ARK_ARC_1_4/buf_output[29] ,
         \MC_ARK_ARC_1_4/buf_output[28] , \MC_ARK_ARC_1_4/buf_output[27] ,
         \MC_ARK_ARC_1_4/buf_output[26] , \MC_ARK_ARC_1_4/buf_output[25] ,
         \MC_ARK_ARC_1_4/buf_output[24] , \MC_ARK_ARC_1_4/buf_output[23] ,
         \MC_ARK_ARC_1_4/buf_output[22] , \MC_ARK_ARC_1_4/buf_output[21] ,
         \MC_ARK_ARC_1_4/buf_output[20] , \MC_ARK_ARC_1_4/buf_output[19] ,
         \MC_ARK_ARC_1_4/buf_output[18] , \MC_ARK_ARC_1_4/buf_output[17] ,
         \MC_ARK_ARC_1_4/buf_output[16] , \MC_ARK_ARC_1_4/buf_output[15] ,
         \MC_ARK_ARC_1_4/buf_output[14] , \MC_ARK_ARC_1_4/buf_output[13] ,
         \MC_ARK_ARC_1_4/buf_output[12] , \MC_ARK_ARC_1_4/buf_output[11] ,
         \MC_ARK_ARC_1_4/buf_output[10] , \MC_ARK_ARC_1_4/buf_output[9] ,
         \MC_ARK_ARC_1_4/buf_output[8] , \MC_ARK_ARC_1_4/buf_output[7] ,
         \MC_ARK_ARC_1_4/buf_output[6] , \MC_ARK_ARC_1_4/buf_output[4] ,
         \MC_ARK_ARC_1_4/buf_output[3] , \MC_ARK_ARC_1_4/buf_output[2] ,
         \MC_ARK_ARC_1_4/buf_output[1] , \MC_ARK_ARC_1_4/buf_output[0] ,
         \MC_ARK_ARC_1_4/temp6[190] , \MC_ARK_ARC_1_4/temp6[188] ,
         \MC_ARK_ARC_1_4/temp6[187] , \MC_ARK_ARC_1_4/temp6[185] ,
         \MC_ARK_ARC_1_4/temp6[181] , \MC_ARK_ARC_1_4/temp6[178] ,
         \MC_ARK_ARC_1_4/temp6[176] , \MC_ARK_ARC_1_4/temp6[175] ,
         \MC_ARK_ARC_1_4/temp6[174] , \MC_ARK_ARC_1_4/temp6[172] ,
         \MC_ARK_ARC_1_4/temp6[169] , \MC_ARK_ARC_1_4/temp6[168] ,
         \MC_ARK_ARC_1_4/temp6[167] , \MC_ARK_ARC_1_4/temp6[166] ,
         \MC_ARK_ARC_1_4/temp6[165] , \MC_ARK_ARC_1_4/temp6[164] ,
         \MC_ARK_ARC_1_4/temp6[162] , \MC_ARK_ARC_1_4/temp6[161] ,
         \MC_ARK_ARC_1_4/temp6[157] , \MC_ARK_ARC_1_4/temp6[156] ,
         \MC_ARK_ARC_1_4/temp6[154] , \MC_ARK_ARC_1_4/temp6[153] ,
         \MC_ARK_ARC_1_4/temp6[150] , \MC_ARK_ARC_1_4/temp6[148] ,
         \MC_ARK_ARC_1_4/temp6[146] , \MC_ARK_ARC_1_4/temp6[145] ,
         \MC_ARK_ARC_1_4/temp6[144] , \MC_ARK_ARC_1_4/temp6[143] ,
         \MC_ARK_ARC_1_4/temp6[142] , \MC_ARK_ARC_1_4/temp6[141] ,
         \MC_ARK_ARC_1_4/temp6[140] , \MC_ARK_ARC_1_4/temp6[136] ,
         \MC_ARK_ARC_1_4/temp6[135] , \MC_ARK_ARC_1_4/temp6[134] ,
         \MC_ARK_ARC_1_4/temp6[133] , \MC_ARK_ARC_1_4/temp6[132] ,
         \MC_ARK_ARC_1_4/temp6[131] , \MC_ARK_ARC_1_4/temp6[129] ,
         \MC_ARK_ARC_1_4/temp6[128] , \MC_ARK_ARC_1_4/temp6[127] ,
         \MC_ARK_ARC_1_4/temp6[125] , \MC_ARK_ARC_1_4/temp6[124] ,
         \MC_ARK_ARC_1_4/temp6[121] , \MC_ARK_ARC_1_4/temp6[118] ,
         \MC_ARK_ARC_1_4/temp6[117] , \MC_ARK_ARC_1_4/temp6[112] ,
         \MC_ARK_ARC_1_4/temp6[111] , \MC_ARK_ARC_1_4/temp6[108] ,
         \MC_ARK_ARC_1_4/temp6[104] , \MC_ARK_ARC_1_4/temp6[102] ,
         \MC_ARK_ARC_1_4/temp6[100] , \MC_ARK_ARC_1_4/temp6[99] ,
         \MC_ARK_ARC_1_4/temp6[98] , \MC_ARK_ARC_1_4/temp6[96] ,
         \MC_ARK_ARC_1_4/temp6[94] , \MC_ARK_ARC_1_4/temp6[92] ,
         \MC_ARK_ARC_1_4/temp6[91] , \MC_ARK_ARC_1_4/temp6[90] ,
         \MC_ARK_ARC_1_4/temp6[88] , \MC_ARK_ARC_1_4/temp6[85] ,
         \MC_ARK_ARC_1_4/temp6[84] , \MC_ARK_ARC_1_4/temp6[83] ,
         \MC_ARK_ARC_1_4/temp6[82] , \MC_ARK_ARC_1_4/temp6[81] ,
         \MC_ARK_ARC_1_4/temp6[79] , \MC_ARK_ARC_1_4/temp6[78] ,
         \MC_ARK_ARC_1_4/temp6[76] , \MC_ARK_ARC_1_4/temp6[72] ,
         \MC_ARK_ARC_1_4/temp6[70] , \MC_ARK_ARC_1_4/temp6[68] ,
         \MC_ARK_ARC_1_4/temp6[67] , \MC_ARK_ARC_1_4/temp6[66] ,
         \MC_ARK_ARC_1_4/temp6[64] , \MC_ARK_ARC_1_4/temp6[60] ,
         \MC_ARK_ARC_1_4/temp6[59] , \MC_ARK_ARC_1_4/temp6[57] ,
         \MC_ARK_ARC_1_4/temp6[54] , \MC_ARK_ARC_1_4/temp6[53] ,
         \MC_ARK_ARC_1_4/temp6[52] , \MC_ARK_ARC_1_4/temp6[51] ,
         \MC_ARK_ARC_1_4/temp6[50] , \MC_ARK_ARC_1_4/temp6[48] ,
         \MC_ARK_ARC_1_4/temp6[47] , \MC_ARK_ARC_1_4/temp6[45] ,
         \MC_ARK_ARC_1_4/temp6[43] , \MC_ARK_ARC_1_4/temp6[42] ,
         \MC_ARK_ARC_1_4/temp6[39] , \MC_ARK_ARC_1_4/temp6[38] ,
         \MC_ARK_ARC_1_4/temp6[37] , \MC_ARK_ARC_1_4/temp6[36] ,
         \MC_ARK_ARC_1_4/temp6[34] , \MC_ARK_ARC_1_4/temp6[33] ,
         \MC_ARK_ARC_1_4/temp6[32] , \MC_ARK_ARC_1_4/temp6[30] ,
         \MC_ARK_ARC_1_4/temp6[28] , \MC_ARK_ARC_1_4/temp6[23] ,
         \MC_ARK_ARC_1_4/temp6[18] , \MC_ARK_ARC_1_4/temp6[14] ,
         \MC_ARK_ARC_1_4/temp6[12] , \MC_ARK_ARC_1_4/temp6[11] ,
         \MC_ARK_ARC_1_4/temp6[10] , \MC_ARK_ARC_1_4/temp6[9] ,
         \MC_ARK_ARC_1_4/temp6[8] , \MC_ARK_ARC_1_4/temp6[5] ,
         \MC_ARK_ARC_1_4/temp6[4] , \MC_ARK_ARC_1_4/temp6[3] ,
         \MC_ARK_ARC_1_4/temp6[1] , \MC_ARK_ARC_1_4/temp5[187] ,
         \MC_ARK_ARC_1_4/temp5[185] , \MC_ARK_ARC_1_4/temp5[184] ,
         \MC_ARK_ARC_1_4/temp5[180] , \MC_ARK_ARC_1_4/temp5[179] ,
         \MC_ARK_ARC_1_4/temp5[178] , \MC_ARK_ARC_1_4/temp5[175] ,
         \MC_ARK_ARC_1_4/temp5[173] , \MC_ARK_ARC_1_4/temp5[172] ,
         \MC_ARK_ARC_1_4/temp5[171] , \MC_ARK_ARC_1_4/temp5[170] ,
         \MC_ARK_ARC_1_4/temp5[169] , \MC_ARK_ARC_1_4/temp5[168] ,
         \MC_ARK_ARC_1_4/temp5[167] , \MC_ARK_ARC_1_4/temp5[164] ,
         \MC_ARK_ARC_1_4/temp5[162] , \MC_ARK_ARC_1_4/temp5[160] ,
         \MC_ARK_ARC_1_4/temp5[159] , \MC_ARK_ARC_1_4/temp5[158] ,
         \MC_ARK_ARC_1_4/temp5[157] , \MC_ARK_ARC_1_4/temp5[156] ,
         \MC_ARK_ARC_1_4/temp5[154] , \MC_ARK_ARC_1_4/temp5[152] ,
         \MC_ARK_ARC_1_4/temp5[151] , \MC_ARK_ARC_1_4/temp5[150] ,
         \MC_ARK_ARC_1_4/temp5[148] , \MC_ARK_ARC_1_4/temp5[145] ,
         \MC_ARK_ARC_1_4/temp5[144] , \MC_ARK_ARC_1_4/temp5[143] ,
         \MC_ARK_ARC_1_4/temp5[142] , \MC_ARK_ARC_1_4/temp5[141] ,
         \MC_ARK_ARC_1_4/temp5[140] , \MC_ARK_ARC_1_4/temp5[138] ,
         \MC_ARK_ARC_1_4/temp5[137] , \MC_ARK_ARC_1_4/temp5[136] ,
         \MC_ARK_ARC_1_4/temp5[135] , \MC_ARK_ARC_1_4/temp5[133] ,
         \MC_ARK_ARC_1_4/temp5[132] , \MC_ARK_ARC_1_4/temp5[131] ,
         \MC_ARK_ARC_1_4/temp5[128] , \MC_ARK_ARC_1_4/temp5[126] ,
         \MC_ARK_ARC_1_4/temp5[125] , \MC_ARK_ARC_1_4/temp5[124] ,
         \MC_ARK_ARC_1_4/temp5[122] , \MC_ARK_ARC_1_4/temp5[121] ,
         \MC_ARK_ARC_1_4/temp5[120] , \MC_ARK_ARC_1_4/temp5[119] ,
         \MC_ARK_ARC_1_4/temp5[114] , \MC_ARK_ARC_1_4/temp5[112] ,
         \MC_ARK_ARC_1_4/temp5[111] , \MC_ARK_ARC_1_4/temp5[106] ,
         \MC_ARK_ARC_1_4/temp5[105] , \MC_ARK_ARC_1_4/temp5[104] ,
         \MC_ARK_ARC_1_4/temp5[102] , \MC_ARK_ARC_1_4/temp5[98] ,
         \MC_ARK_ARC_1_4/temp5[97] , \MC_ARK_ARC_1_4/temp5[96] ,
         \MC_ARK_ARC_1_4/temp5[94] , \MC_ARK_ARC_1_4/temp5[92] ,
         \MC_ARK_ARC_1_4/temp5[91] , \MC_ARK_ARC_1_4/temp5[90] ,
         \MC_ARK_ARC_1_4/temp5[89] , \MC_ARK_ARC_1_4/temp5[85] ,
         \MC_ARK_ARC_1_4/temp5[84] , \MC_ARK_ARC_1_4/temp5[83] ,
         \MC_ARK_ARC_1_4/temp5[82] , \MC_ARK_ARC_1_4/temp5[79] ,
         \MC_ARK_ARC_1_4/temp5[76] , \MC_ARK_ARC_1_4/temp5[73] ,
         \MC_ARK_ARC_1_4/temp5[71] , \MC_ARK_ARC_1_4/temp5[70] ,
         \MC_ARK_ARC_1_4/temp5[69] , \MC_ARK_ARC_1_4/temp5[68] ,
         \MC_ARK_ARC_1_4/temp5[67] , \MC_ARK_ARC_1_4/temp5[64] ,
         \MC_ARK_ARC_1_4/temp5[63] , \MC_ARK_ARC_1_4/temp5[61] ,
         \MC_ARK_ARC_1_4/temp5[59] , \MC_ARK_ARC_1_4/temp5[57] ,
         \MC_ARK_ARC_1_4/temp5[55] , \MC_ARK_ARC_1_4/temp5[53] ,
         \MC_ARK_ARC_1_4/temp5[52] , \MC_ARK_ARC_1_4/temp5[51] ,
         \MC_ARK_ARC_1_4/temp5[49] , \MC_ARK_ARC_1_4/temp5[47] ,
         \MC_ARK_ARC_1_4/temp5[46] , \MC_ARK_ARC_1_4/temp5[44] ,
         \MC_ARK_ARC_1_4/temp5[43] , \MC_ARK_ARC_1_4/temp5[40] ,
         \MC_ARK_ARC_1_4/temp5[37] , \MC_ARK_ARC_1_4/temp5[36] ,
         \MC_ARK_ARC_1_4/temp5[34] , \MC_ARK_ARC_1_4/temp5[32] ,
         \MC_ARK_ARC_1_4/temp5[31] , \MC_ARK_ARC_1_4/temp5[30] ,
         \MC_ARK_ARC_1_4/temp5[28] , \MC_ARK_ARC_1_4/temp5[27] ,
         \MC_ARK_ARC_1_4/temp5[26] , \MC_ARK_ARC_1_4/temp5[25] ,
         \MC_ARK_ARC_1_4/temp5[23] , \MC_ARK_ARC_1_4/temp5[22] ,
         \MC_ARK_ARC_1_4/temp5[21] , \MC_ARK_ARC_1_4/temp5[18] ,
         \MC_ARK_ARC_1_4/temp5[16] , \MC_ARK_ARC_1_4/temp5[14] ,
         \MC_ARK_ARC_1_4/temp5[13] , \MC_ARK_ARC_1_4/temp5[12] ,
         \MC_ARK_ARC_1_4/temp5[8] , \MC_ARK_ARC_1_4/temp5[5] ,
         \MC_ARK_ARC_1_4/temp5[4] , \MC_ARK_ARC_1_4/temp5[3] ,
         \MC_ARK_ARC_1_4/temp5[0] , \MC_ARK_ARC_1_4/temp4[191] ,
         \MC_ARK_ARC_1_4/temp4[190] , \MC_ARK_ARC_1_4/temp4[189] ,
         \MC_ARK_ARC_1_4/temp4[188] , \MC_ARK_ARC_1_4/temp4[187] ,
         \MC_ARK_ARC_1_4/temp4[186] , \MC_ARK_ARC_1_4/temp4[184] ,
         \MC_ARK_ARC_1_4/temp4[183] , \MC_ARK_ARC_1_4/temp4[182] ,
         \MC_ARK_ARC_1_4/temp4[181] , \MC_ARK_ARC_1_4/temp4[180] ,
         \MC_ARK_ARC_1_4/temp4[179] , \MC_ARK_ARC_1_4/temp4[178] ,
         \MC_ARK_ARC_1_4/temp4[177] , \MC_ARK_ARC_1_4/temp4[176] ,
         \MC_ARK_ARC_1_4/temp4[175] , \MC_ARK_ARC_1_4/temp4[174] ,
         \MC_ARK_ARC_1_4/temp4[172] , \MC_ARK_ARC_1_4/temp4[171] ,
         \MC_ARK_ARC_1_4/temp4[170] , \MC_ARK_ARC_1_4/temp4[169] ,
         \MC_ARK_ARC_1_4/temp4[168] , \MC_ARK_ARC_1_4/temp4[167] ,
         \MC_ARK_ARC_1_4/temp4[166] , \MC_ARK_ARC_1_4/temp4[165] ,
         \MC_ARK_ARC_1_4/temp4[164] , \MC_ARK_ARC_1_4/temp4[163] ,
         \MC_ARK_ARC_1_4/temp4[162] , \MC_ARK_ARC_1_4/temp4[161] ,
         \MC_ARK_ARC_1_4/temp4[160] , \MC_ARK_ARC_1_4/temp4[159] ,
         \MC_ARK_ARC_1_4/temp4[158] , \MC_ARK_ARC_1_4/temp4[157] ,
         \MC_ARK_ARC_1_4/temp4[156] , \MC_ARK_ARC_1_4/temp4[155] ,
         \MC_ARK_ARC_1_4/temp4[154] , \MC_ARK_ARC_1_4/temp4[153] ,
         \MC_ARK_ARC_1_4/temp4[152] , \MC_ARK_ARC_1_4/temp4[151] ,
         \MC_ARK_ARC_1_4/temp4[150] , \MC_ARK_ARC_1_4/temp4[149] ,
         \MC_ARK_ARC_1_4/temp4[148] , \MC_ARK_ARC_1_4/temp4[147] ,
         \MC_ARK_ARC_1_4/temp4[146] , \MC_ARK_ARC_1_4/temp4[145] ,
         \MC_ARK_ARC_1_4/temp4[144] , \MC_ARK_ARC_1_4/temp4[143] ,
         \MC_ARK_ARC_1_4/temp4[142] , \MC_ARK_ARC_1_4/temp4[141] ,
         \MC_ARK_ARC_1_4/temp4[140] , \MC_ARK_ARC_1_4/temp4[139] ,
         \MC_ARK_ARC_1_4/temp4[138] , \MC_ARK_ARC_1_4/temp4[137] ,
         \MC_ARK_ARC_1_4/temp4[136] , \MC_ARK_ARC_1_4/temp4[135] ,
         \MC_ARK_ARC_1_4/temp4[134] , \MC_ARK_ARC_1_4/temp4[133] ,
         \MC_ARK_ARC_1_4/temp4[132] , \MC_ARK_ARC_1_4/temp4[131] ,
         \MC_ARK_ARC_1_4/temp4[130] , \MC_ARK_ARC_1_4/temp4[129] ,
         \MC_ARK_ARC_1_4/temp4[128] , \MC_ARK_ARC_1_4/temp4[127] ,
         \MC_ARK_ARC_1_4/temp4[126] , \MC_ARK_ARC_1_4/temp4[125] ,
         \MC_ARK_ARC_1_4/temp4[123] , \MC_ARK_ARC_1_4/temp4[122] ,
         \MC_ARK_ARC_1_4/temp4[121] , \MC_ARK_ARC_1_4/temp4[120] ,
         \MC_ARK_ARC_1_4/temp4[119] , \MC_ARK_ARC_1_4/temp4[118] ,
         \MC_ARK_ARC_1_4/temp4[117] , \MC_ARK_ARC_1_4/temp4[116] ,
         \MC_ARK_ARC_1_4/temp4[115] , \MC_ARK_ARC_1_4/temp4[114] ,
         \MC_ARK_ARC_1_4/temp4[112] , \MC_ARK_ARC_1_4/temp4[111] ,
         \MC_ARK_ARC_1_4/temp4[110] , \MC_ARK_ARC_1_4/temp4[109] ,
         \MC_ARK_ARC_1_4/temp4[108] , \MC_ARK_ARC_1_4/temp4[107] ,
         \MC_ARK_ARC_1_4/temp4[106] , \MC_ARK_ARC_1_4/temp4[105] ,
         \MC_ARK_ARC_1_4/temp4[104] , \MC_ARK_ARC_1_4/temp4[103] ,
         \MC_ARK_ARC_1_4/temp4[102] , \MC_ARK_ARC_1_4/temp4[101] ,
         \MC_ARK_ARC_1_4/temp4[100] , \MC_ARK_ARC_1_4/temp4[99] ,
         \MC_ARK_ARC_1_4/temp4[98] , \MC_ARK_ARC_1_4/temp4[97] ,
         \MC_ARK_ARC_1_4/temp4[96] , \MC_ARK_ARC_1_4/temp4[95] ,
         \MC_ARK_ARC_1_4/temp4[94] , \MC_ARK_ARC_1_4/temp4[93] ,
         \MC_ARK_ARC_1_4/temp4[91] , \MC_ARK_ARC_1_4/temp4[90] ,
         \MC_ARK_ARC_1_4/temp4[89] , \MC_ARK_ARC_1_4/temp4[88] ,
         \MC_ARK_ARC_1_4/temp4[87] , \MC_ARK_ARC_1_4/temp4[86] ,
         \MC_ARK_ARC_1_4/temp4[85] , \MC_ARK_ARC_1_4/temp4[84] ,
         \MC_ARK_ARC_1_4/temp4[83] , \MC_ARK_ARC_1_4/temp4[82] ,
         \MC_ARK_ARC_1_4/temp4[81] , \MC_ARK_ARC_1_4/temp4[80] ,
         \MC_ARK_ARC_1_4/temp4[79] , \MC_ARK_ARC_1_4/temp4[78] ,
         \MC_ARK_ARC_1_4/temp4[77] , \MC_ARK_ARC_1_4/temp4[76] ,
         \MC_ARK_ARC_1_4/temp4[75] , \MC_ARK_ARC_1_4/temp4[74] ,
         \MC_ARK_ARC_1_4/temp4[73] , \MC_ARK_ARC_1_4/temp4[72] ,
         \MC_ARK_ARC_1_4/temp4[71] , \MC_ARK_ARC_1_4/temp4[70] ,
         \MC_ARK_ARC_1_4/temp4[69] , \MC_ARK_ARC_1_4/temp4[68] ,
         \MC_ARK_ARC_1_4/temp4[67] , \MC_ARK_ARC_1_4/temp4[66] ,
         \MC_ARK_ARC_1_4/temp4[65] , \MC_ARK_ARC_1_4/temp4[64] ,
         \MC_ARK_ARC_1_4/temp4[63] , \MC_ARK_ARC_1_4/temp4[62] ,
         \MC_ARK_ARC_1_4/temp4[61] , \MC_ARK_ARC_1_4/temp4[60] ,
         \MC_ARK_ARC_1_4/temp4[59] , \MC_ARK_ARC_1_4/temp4[58] ,
         \MC_ARK_ARC_1_4/temp4[57] , \MC_ARK_ARC_1_4/temp4[56] ,
         \MC_ARK_ARC_1_4/temp4[55] , \MC_ARK_ARC_1_4/temp4[54] ,
         \MC_ARK_ARC_1_4/temp4[53] , \MC_ARK_ARC_1_4/temp4[52] ,
         \MC_ARK_ARC_1_4/temp4[51] , \MC_ARK_ARC_1_4/temp4[50] ,
         \MC_ARK_ARC_1_4/temp4[49] , \MC_ARK_ARC_1_4/temp4[48] ,
         \MC_ARK_ARC_1_4/temp4[47] , \MC_ARK_ARC_1_4/temp4[46] ,
         \MC_ARK_ARC_1_4/temp4[45] , \MC_ARK_ARC_1_4/temp4[44] ,
         \MC_ARK_ARC_1_4/temp4[43] , \MC_ARK_ARC_1_4/temp4[42] ,
         \MC_ARK_ARC_1_4/temp4[41] , \MC_ARK_ARC_1_4/temp4[40] ,
         \MC_ARK_ARC_1_4/temp4[38] , \MC_ARK_ARC_1_4/temp4[37] ,
         \MC_ARK_ARC_1_4/temp4[36] , \MC_ARK_ARC_1_4/temp4[35] ,
         \MC_ARK_ARC_1_4/temp4[34] , \MC_ARK_ARC_1_4/temp4[32] ,
         \MC_ARK_ARC_1_4/temp4[31] , \MC_ARK_ARC_1_4/temp4[30] ,
         \MC_ARK_ARC_1_4/temp4[29] , \MC_ARK_ARC_1_4/temp4[28] ,
         \MC_ARK_ARC_1_4/temp4[27] , \MC_ARK_ARC_1_4/temp4[26] ,
         \MC_ARK_ARC_1_4/temp4[25] , \MC_ARK_ARC_1_4/temp4[24] ,
         \MC_ARK_ARC_1_4/temp4[23] , \MC_ARK_ARC_1_4/temp4[22] ,
         \MC_ARK_ARC_1_4/temp4[21] , \MC_ARK_ARC_1_4/temp4[20] ,
         \MC_ARK_ARC_1_4/temp4[19] , \MC_ARK_ARC_1_4/temp4[18] ,
         \MC_ARK_ARC_1_4/temp4[17] , \MC_ARK_ARC_1_4/temp4[16] ,
         \MC_ARK_ARC_1_4/temp4[15] , \MC_ARK_ARC_1_4/temp4[14] ,
         \MC_ARK_ARC_1_4/temp4[13] , \MC_ARK_ARC_1_4/temp4[12] ,
         \MC_ARK_ARC_1_4/temp4[10] , \MC_ARK_ARC_1_4/temp4[9] ,
         \MC_ARK_ARC_1_4/temp4[8] , \MC_ARK_ARC_1_4/temp4[7] ,
         \MC_ARK_ARC_1_4/temp4[6] , \MC_ARK_ARC_1_4/temp4[5] ,
         \MC_ARK_ARC_1_4/temp4[4] , \MC_ARK_ARC_1_4/temp4[3] ,
         \MC_ARK_ARC_1_4/temp4[2] , \MC_ARK_ARC_1_4/temp4[1] ,
         \MC_ARK_ARC_1_4/temp4[0] , \MC_ARK_ARC_1_4/temp3[191] ,
         \MC_ARK_ARC_1_4/temp3[190] , \MC_ARK_ARC_1_4/temp3[187] ,
         \MC_ARK_ARC_1_4/temp3[186] , \MC_ARK_ARC_1_4/temp3[184] ,
         \MC_ARK_ARC_1_4/temp3[182] , \MC_ARK_ARC_1_4/temp3[181] ,
         \MC_ARK_ARC_1_4/temp3[180] , \MC_ARK_ARC_1_4/temp3[178] ,
         \MC_ARK_ARC_1_4/temp3[177] , \MC_ARK_ARC_1_4/temp3[176] ,
         \MC_ARK_ARC_1_4/temp3[175] , \MC_ARK_ARC_1_4/temp3[174] ,
         \MC_ARK_ARC_1_4/temp3[172] , \MC_ARK_ARC_1_4/temp3[171] ,
         \MC_ARK_ARC_1_4/temp3[170] , \MC_ARK_ARC_1_4/temp3[169] ,
         \MC_ARK_ARC_1_4/temp3[167] , \MC_ARK_ARC_1_4/temp3[166] ,
         \MC_ARK_ARC_1_4/temp3[165] , \MC_ARK_ARC_1_4/temp3[164] ,
         \MC_ARK_ARC_1_4/temp3[163] , \MC_ARK_ARC_1_4/temp3[162] ,
         \MC_ARK_ARC_1_4/temp3[161] , \MC_ARK_ARC_1_4/temp3[160] ,
         \MC_ARK_ARC_1_4/temp3[159] , \MC_ARK_ARC_1_4/temp3[158] ,
         \MC_ARK_ARC_1_4/temp3[157] , \MC_ARK_ARC_1_4/temp3[156] ,
         \MC_ARK_ARC_1_4/temp3[155] , \MC_ARK_ARC_1_4/temp3[154] ,
         \MC_ARK_ARC_1_4/temp3[153] , \MC_ARK_ARC_1_4/temp3[151] ,
         \MC_ARK_ARC_1_4/temp3[150] , \MC_ARK_ARC_1_4/temp3[149] ,
         \MC_ARK_ARC_1_4/temp3[148] , \MC_ARK_ARC_1_4/temp3[146] ,
         \MC_ARK_ARC_1_4/temp3[145] , \MC_ARK_ARC_1_4/temp3[144] ,
         \MC_ARK_ARC_1_4/temp3[143] , \MC_ARK_ARC_1_4/temp3[142] ,
         \MC_ARK_ARC_1_4/temp3[141] , \MC_ARK_ARC_1_4/temp3[140] ,
         \MC_ARK_ARC_1_4/temp3[139] , \MC_ARK_ARC_1_4/temp3[138] ,
         \MC_ARK_ARC_1_4/temp3[137] , \MC_ARK_ARC_1_4/temp3[136] ,
         \MC_ARK_ARC_1_4/temp3[134] , \MC_ARK_ARC_1_4/temp3[133] ,
         \MC_ARK_ARC_1_4/temp3[132] , \MC_ARK_ARC_1_4/temp3[131] ,
         \MC_ARK_ARC_1_4/temp3[130] , \MC_ARK_ARC_1_4/temp3[129] ,
         \MC_ARK_ARC_1_4/temp3[128] , \MC_ARK_ARC_1_4/temp3[127] ,
         \MC_ARK_ARC_1_4/temp3[126] , \MC_ARK_ARC_1_4/temp3[125] ,
         \MC_ARK_ARC_1_4/temp3[123] , \MC_ARK_ARC_1_4/temp3[121] ,
         \MC_ARK_ARC_1_4/temp3[120] , \MC_ARK_ARC_1_4/temp3[119] ,
         \MC_ARK_ARC_1_4/temp3[118] , \MC_ARK_ARC_1_4/temp3[117] ,
         \MC_ARK_ARC_1_4/temp3[115] , \MC_ARK_ARC_1_4/temp3[114] ,
         \MC_ARK_ARC_1_4/temp3[112] , \MC_ARK_ARC_1_4/temp3[110] ,
         \MC_ARK_ARC_1_4/temp3[109] , \MC_ARK_ARC_1_4/temp3[107] ,
         \MC_ARK_ARC_1_4/temp3[106] , \MC_ARK_ARC_1_4/temp3[104] ,
         \MC_ARK_ARC_1_4/temp3[103] , \MC_ARK_ARC_1_4/temp3[102] ,
         \MC_ARK_ARC_1_4/temp3[100] , \MC_ARK_ARC_1_4/temp3[97] ,
         \MC_ARK_ARC_1_4/temp3[96] , \MC_ARK_ARC_1_4/temp3[94] ,
         \MC_ARK_ARC_1_4/temp3[91] , \MC_ARK_ARC_1_4/temp3[90] ,
         \MC_ARK_ARC_1_4/temp3[88] , \MC_ARK_ARC_1_4/temp3[86] ,
         \MC_ARK_ARC_1_4/temp3[85] , \MC_ARK_ARC_1_4/temp3[84] ,
         \MC_ARK_ARC_1_4/temp3[83] , \MC_ARK_ARC_1_4/temp3[79] ,
         \MC_ARK_ARC_1_4/temp3[78] , \MC_ARK_ARC_1_4/temp3[77] ,
         \MC_ARK_ARC_1_4/temp3[76] , \MC_ARK_ARC_1_4/temp3[73] ,
         \MC_ARK_ARC_1_4/temp3[72] , \MC_ARK_ARC_1_4/temp3[71] ,
         \MC_ARK_ARC_1_4/temp3[70] , \MC_ARK_ARC_1_4/temp3[69] ,
         \MC_ARK_ARC_1_4/temp3[67] , \MC_ARK_ARC_1_4/temp3[66] ,
         \MC_ARK_ARC_1_4/temp3[64] , \MC_ARK_ARC_1_4/temp3[63] ,
         \MC_ARK_ARC_1_4/temp3[61] , \MC_ARK_ARC_1_4/temp3[60] ,
         \MC_ARK_ARC_1_4/temp3[59] , \MC_ARK_ARC_1_4/temp3[58] ,
         \MC_ARK_ARC_1_4/temp3[57] , \MC_ARK_ARC_1_4/temp3[56] ,
         \MC_ARK_ARC_1_4/temp3[55] , \MC_ARK_ARC_1_4/temp3[54] ,
         \MC_ARK_ARC_1_4/temp3[53] , \MC_ARK_ARC_1_4/temp3[52] ,
         \MC_ARK_ARC_1_4/temp3[50] , \MC_ARK_ARC_1_4/temp3[49] ,
         \MC_ARK_ARC_1_4/temp3[48] , \MC_ARK_ARC_1_4/temp3[47] ,
         \MC_ARK_ARC_1_4/temp3[46] , \MC_ARK_ARC_1_4/temp3[45] ,
         \MC_ARK_ARC_1_4/temp3[43] , \MC_ARK_ARC_1_4/temp3[42] ,
         \MC_ARK_ARC_1_4/temp3[41] , \MC_ARK_ARC_1_4/temp3[37] ,
         \MC_ARK_ARC_1_4/temp3[36] , \MC_ARK_ARC_1_4/temp3[34] ,
         \MC_ARK_ARC_1_4/temp3[32] , \MC_ARK_ARC_1_4/temp3[31] ,
         \MC_ARK_ARC_1_4/temp3[30] , \MC_ARK_ARC_1_4/temp3[28] ,
         \MC_ARK_ARC_1_4/temp3[27] , \MC_ARK_ARC_1_4/temp3[26] ,
         \MC_ARK_ARC_1_4/temp3[25] , \MC_ARK_ARC_1_4/temp3[24] ,
         \MC_ARK_ARC_1_4/temp3[22] , \MC_ARK_ARC_1_4/temp3[19] ,
         \MC_ARK_ARC_1_4/temp3[18] , \MC_ARK_ARC_1_4/temp3[16] ,
         \MC_ARK_ARC_1_4/temp3[14] , \MC_ARK_ARC_1_4/temp3[13] ,
         \MC_ARK_ARC_1_4/temp3[12] , \MC_ARK_ARC_1_4/temp3[10] ,
         \MC_ARK_ARC_1_4/temp3[9] , \MC_ARK_ARC_1_4/temp3[8] ,
         \MC_ARK_ARC_1_4/temp3[7] , \MC_ARK_ARC_1_4/temp3[6] ,
         \MC_ARK_ARC_1_4/temp3[4] , \MC_ARK_ARC_1_4/temp3[3] ,
         \MC_ARK_ARC_1_4/temp3[1] , \MC_ARK_ARC_1_4/temp2[190] ,
         \MC_ARK_ARC_1_4/temp2[188] , \MC_ARK_ARC_1_4/temp2[187] ,
         \MC_ARK_ARC_1_4/temp2[186] , \MC_ARK_ARC_1_4/temp2[184] ,
         \MC_ARK_ARC_1_4/temp2[182] , \MC_ARK_ARC_1_4/temp2[181] ,
         \MC_ARK_ARC_1_4/temp2[180] , \MC_ARK_ARC_1_4/temp2[178] ,
         \MC_ARK_ARC_1_4/temp2[177] , \MC_ARK_ARC_1_4/temp2[175] ,
         \MC_ARK_ARC_1_4/temp2[174] , \MC_ARK_ARC_1_4/temp2[172] ,
         \MC_ARK_ARC_1_4/temp2[171] , \MC_ARK_ARC_1_4/temp2[170] ,
         \MC_ARK_ARC_1_4/temp2[169] , \MC_ARK_ARC_1_4/temp2[168] ,
         \MC_ARK_ARC_1_4/temp2[167] , \MC_ARK_ARC_1_4/temp2[166] ,
         \MC_ARK_ARC_1_4/temp2[165] , \MC_ARK_ARC_1_4/temp2[163] ,
         \MC_ARK_ARC_1_4/temp2[162] , \MC_ARK_ARC_1_4/temp2[161] ,
         \MC_ARK_ARC_1_4/temp2[160] , \MC_ARK_ARC_1_4/temp2[159] ,
         \MC_ARK_ARC_1_4/temp2[158] , \MC_ARK_ARC_1_4/temp2[157] ,
         \MC_ARK_ARC_1_4/temp2[156] , \MC_ARK_ARC_1_4/temp2[154] ,
         \MC_ARK_ARC_1_4/temp2[153] , \MC_ARK_ARC_1_4/temp2[151] ,
         \MC_ARK_ARC_1_4/temp2[148] , \MC_ARK_ARC_1_4/temp2[145] ,
         \MC_ARK_ARC_1_4/temp2[144] , \MC_ARK_ARC_1_4/temp2[143] ,
         \MC_ARK_ARC_1_4/temp2[142] , \MC_ARK_ARC_1_4/temp2[141] ,
         \MC_ARK_ARC_1_4/temp2[140] , \MC_ARK_ARC_1_4/temp2[138] ,
         \MC_ARK_ARC_1_4/temp2[137] , \MC_ARK_ARC_1_4/temp2[136] ,
         \MC_ARK_ARC_1_4/temp2[135] , \MC_ARK_ARC_1_4/temp2[134] ,
         \MC_ARK_ARC_1_4/temp2[132] , \MC_ARK_ARC_1_4/temp2[131] ,
         \MC_ARK_ARC_1_4/temp2[130] , \MC_ARK_ARC_1_4/temp2[128] ,
         \MC_ARK_ARC_1_4/temp2[126] , \MC_ARK_ARC_1_4/temp2[124] ,
         \MC_ARK_ARC_1_4/temp2[123] , \MC_ARK_ARC_1_4/temp2[121] ,
         \MC_ARK_ARC_1_4/temp2[120] , \MC_ARK_ARC_1_4/temp2[119] ,
         \MC_ARK_ARC_1_4/temp2[118] , \MC_ARK_ARC_1_4/temp2[115] ,
         \MC_ARK_ARC_1_4/temp2[112] , \MC_ARK_ARC_1_4/temp2[110] ,
         \MC_ARK_ARC_1_4/temp2[109] , \MC_ARK_ARC_1_4/temp2[108] ,
         \MC_ARK_ARC_1_4/temp2[106] , \MC_ARK_ARC_1_4/temp2[104] ,
         \MC_ARK_ARC_1_4/temp2[103] , \MC_ARK_ARC_1_4/temp2[100] ,
         \MC_ARK_ARC_1_4/temp2[98] , \MC_ARK_ARC_1_4/temp2[94] ,
         \MC_ARK_ARC_1_4/temp2[93] , \MC_ARK_ARC_1_4/temp2[91] ,
         \MC_ARK_ARC_1_4/temp2[90] , \MC_ARK_ARC_1_4/temp2[88] ,
         \MC_ARK_ARC_1_4/temp2[86] , \MC_ARK_ARC_1_4/temp2[85] ,
         \MC_ARK_ARC_1_4/temp2[84] , \MC_ARK_ARC_1_4/temp2[83] ,
         \MC_ARK_ARC_1_4/temp2[81] , \MC_ARK_ARC_1_4/temp2[80] ,
         \MC_ARK_ARC_1_4/temp2[79] , \MC_ARK_ARC_1_4/temp2[78] ,
         \MC_ARK_ARC_1_4/temp2[77] , \MC_ARK_ARC_1_4/temp2[76] ,
         \MC_ARK_ARC_1_4/temp2[73] , \MC_ARK_ARC_1_4/temp2[72] ,
         \MC_ARK_ARC_1_4/temp2[70] , \MC_ARK_ARC_1_4/temp2[67] ,
         \MC_ARK_ARC_1_4/temp2[66] , \MC_ARK_ARC_1_4/temp2[65] ,
         \MC_ARK_ARC_1_4/temp2[64] , \MC_ARK_ARC_1_4/temp2[63] ,
         \MC_ARK_ARC_1_4/temp2[61] , \MC_ARK_ARC_1_4/temp2[60] ,
         \MC_ARK_ARC_1_4/temp2[58] , \MC_ARK_ARC_1_4/temp2[57] ,
         \MC_ARK_ARC_1_4/temp2[55] , \MC_ARK_ARC_1_4/temp2[54] ,
         \MC_ARK_ARC_1_4/temp2[52] , \MC_ARK_ARC_1_4/temp2[51] ,
         \MC_ARK_ARC_1_4/temp2[49] , \MC_ARK_ARC_1_4/temp2[46] ,
         \MC_ARK_ARC_1_4/temp2[43] , \MC_ARK_ARC_1_4/temp2[42] ,
         \MC_ARK_ARC_1_4/temp2[37] , \MC_ARK_ARC_1_4/temp2[36] ,
         \MC_ARK_ARC_1_4/temp2[34] , \MC_ARK_ARC_1_4/temp2[31] ,
         \MC_ARK_ARC_1_4/temp2[30] , \MC_ARK_ARC_1_4/temp2[29] ,
         \MC_ARK_ARC_1_4/temp2[28] , \MC_ARK_ARC_1_4/temp2[26] ,
         \MC_ARK_ARC_1_4/temp2[24] , \MC_ARK_ARC_1_4/temp2[22] ,
         \MC_ARK_ARC_1_4/temp2[21] , \MC_ARK_ARC_1_4/temp2[18] ,
         \MC_ARK_ARC_1_4/temp2[16] , \MC_ARK_ARC_1_4/temp2[13] ,
         \MC_ARK_ARC_1_4/temp2[12] , \MC_ARK_ARC_1_4/temp2[10] ,
         \MC_ARK_ARC_1_4/temp2[9] , \MC_ARK_ARC_1_4/temp2[7] ,
         \MC_ARK_ARC_1_4/temp2[6] , \MC_ARK_ARC_1_4/temp2[4] ,
         \MC_ARK_ARC_1_4/temp1[190] , \MC_ARK_ARC_1_4/temp1[187] ,
         \MC_ARK_ARC_1_4/temp1[186] , \MC_ARK_ARC_1_4/temp1[184] ,
         \MC_ARK_ARC_1_4/temp1[183] , \MC_ARK_ARC_1_4/temp1[182] ,
         \MC_ARK_ARC_1_4/temp1[181] , \MC_ARK_ARC_1_4/temp1[180] ,
         \MC_ARK_ARC_1_4/temp1[178] , \MC_ARK_ARC_1_4/temp1[177] ,
         \MC_ARK_ARC_1_4/temp1[176] , \MC_ARK_ARC_1_4/temp1[175] ,
         \MC_ARK_ARC_1_4/temp1[174] , \MC_ARK_ARC_1_4/temp1[172] ,
         \MC_ARK_ARC_1_4/temp1[171] , \MC_ARK_ARC_1_4/temp1[169] ,
         \MC_ARK_ARC_1_4/temp1[168] , \MC_ARK_ARC_1_4/temp1[167] ,
         \MC_ARK_ARC_1_4/temp1[166] , \MC_ARK_ARC_1_4/temp1[165] ,
         \MC_ARK_ARC_1_4/temp1[164] , \MC_ARK_ARC_1_4/temp1[163] ,
         \MC_ARK_ARC_1_4/temp1[162] , \MC_ARK_ARC_1_4/temp1[161] ,
         \MC_ARK_ARC_1_4/temp1[160] , \MC_ARK_ARC_1_4/temp1[159] ,
         \MC_ARK_ARC_1_4/temp1[158] , \MC_ARK_ARC_1_4/temp1[157] ,
         \MC_ARK_ARC_1_4/temp1[156] , \MC_ARK_ARC_1_4/temp1[154] ,
         \MC_ARK_ARC_1_4/temp1[153] , \MC_ARK_ARC_1_4/temp1[151] ,
         \MC_ARK_ARC_1_4/temp1[150] , \MC_ARK_ARC_1_4/temp1[148] ,
         \MC_ARK_ARC_1_4/temp1[147] , \MC_ARK_ARC_1_4/temp1[145] ,
         \MC_ARK_ARC_1_4/temp1[144] , \MC_ARK_ARC_1_4/temp1[143] ,
         \MC_ARK_ARC_1_4/temp1[142] , \MC_ARK_ARC_1_4/temp1[141] ,
         \MC_ARK_ARC_1_4/temp1[140] , \MC_ARK_ARC_1_4/temp1[139] ,
         \MC_ARK_ARC_1_4/temp1[138] , \MC_ARK_ARC_1_4/temp1[137] ,
         \MC_ARK_ARC_1_4/temp1[136] , \MC_ARK_ARC_1_4/temp1[133] ,
         \MC_ARK_ARC_1_4/temp1[132] , \MC_ARK_ARC_1_4/temp1[128] ,
         \MC_ARK_ARC_1_4/temp1[127] , \MC_ARK_ARC_1_4/temp1[126] ,
         \MC_ARK_ARC_1_4/temp1[124] , \MC_ARK_ARC_1_4/temp1[123] ,
         \MC_ARK_ARC_1_4/temp1[121] , \MC_ARK_ARC_1_4/temp1[120] ,
         \MC_ARK_ARC_1_4/temp1[117] , \MC_ARK_ARC_1_4/temp1[115] ,
         \MC_ARK_ARC_1_4/temp1[112] , \MC_ARK_ARC_1_4/temp1[109] ,
         \MC_ARK_ARC_1_4/temp1[106] , \MC_ARK_ARC_1_4/temp1[103] ,
         \MC_ARK_ARC_1_4/temp1[102] , \MC_ARK_ARC_1_4/temp1[100] ,
         \MC_ARK_ARC_1_4/temp1[98] , \MC_ARK_ARC_1_4/temp1[96] ,
         \MC_ARK_ARC_1_4/temp1[94] , \MC_ARK_ARC_1_4/temp1[93] ,
         \MC_ARK_ARC_1_4/temp1[90] , \MC_ARK_ARC_1_4/temp1[86] ,
         \MC_ARK_ARC_1_4/temp1[85] , \MC_ARK_ARC_1_4/temp1[84] ,
         \MC_ARK_ARC_1_4/temp1[83] , \MC_ARK_ARC_1_4/temp1[82] ,
         \MC_ARK_ARC_1_4/temp1[80] , \MC_ARK_ARC_1_4/temp1[79] ,
         \MC_ARK_ARC_1_4/temp1[78] , \MC_ARK_ARC_1_4/temp1[77] ,
         \MC_ARK_ARC_1_4/temp1[76] , \MC_ARK_ARC_1_4/temp1[73] ,
         \MC_ARK_ARC_1_4/temp1[72] , \MC_ARK_ARC_1_4/temp1[71] ,
         \MC_ARK_ARC_1_4/temp1[70] , \MC_ARK_ARC_1_4/temp1[67] ,
         \MC_ARK_ARC_1_4/temp1[66] , \MC_ARK_ARC_1_4/temp1[64] ,
         \MC_ARK_ARC_1_4/temp1[63] , \MC_ARK_ARC_1_4/temp1[61] ,
         \MC_ARK_ARC_1_4/temp1[60] , \MC_ARK_ARC_1_4/temp1[58] ,
         \MC_ARK_ARC_1_4/temp1[57] , \MC_ARK_ARC_1_4/temp1[55] ,
         \MC_ARK_ARC_1_4/temp1[54] , \MC_ARK_ARC_1_4/temp1[52] ,
         \MC_ARK_ARC_1_4/temp1[51] , \MC_ARK_ARC_1_4/temp1[50] ,
         \MC_ARK_ARC_1_4/temp1[49] , \MC_ARK_ARC_1_4/temp1[46] ,
         \MC_ARK_ARC_1_4/temp1[45] , \MC_ARK_ARC_1_4/temp1[43] ,
         \MC_ARK_ARC_1_4/temp1[42] , \MC_ARK_ARC_1_4/temp1[41] ,
         \MC_ARK_ARC_1_4/temp1[39] , \MC_ARK_ARC_1_4/temp1[37] ,
         \MC_ARK_ARC_1_4/temp1[36] , \MC_ARK_ARC_1_4/temp1[35] ,
         \MC_ARK_ARC_1_4/temp1[34] , \MC_ARK_ARC_1_4/temp1[33] ,
         \MC_ARK_ARC_1_4/temp1[31] , \MC_ARK_ARC_1_4/temp1[30] ,
         \MC_ARK_ARC_1_4/temp1[29] , \MC_ARK_ARC_1_4/temp1[28] ,
         \MC_ARK_ARC_1_4/temp1[25] , \MC_ARK_ARC_1_4/temp1[24] ,
         \MC_ARK_ARC_1_4/temp1[22] , \MC_ARK_ARC_1_4/temp1[21] ,
         \MC_ARK_ARC_1_4/temp1[18] , \MC_ARK_ARC_1_4/temp1[17] ,
         \MC_ARK_ARC_1_4/temp1[16] , \MC_ARK_ARC_1_4/temp1[15] ,
         \MC_ARK_ARC_1_4/temp1[13] , \MC_ARK_ARC_1_4/temp1[12] ,
         \MC_ARK_ARC_1_4/temp1[10] , \MC_ARK_ARC_1_4/temp1[9] ,
         \MC_ARK_ARC_1_4/temp1[7] , \MC_ARK_ARC_1_4/temp1[4] ,
         \MC_ARK_ARC_1_4/temp1[2] , \MC_ARK_ARC_1_4/temp1[1] ,
         \MC_ARK_ARC_1_4/temp1[0] , \MC_ARK_ARC_1_4/buf_datainput[188] ,
         \MC_ARK_ARC_1_4/buf_datainput[184] ,
         \MC_ARK_ARC_1_4/buf_datainput[183] ,
         \MC_ARK_ARC_1_4/buf_datainput[177] ,
         \MC_ARK_ARC_1_4/buf_datainput[176] ,
         \MC_ARK_ARC_1_4/buf_datainput[173] ,
         \MC_ARK_ARC_1_4/buf_datainput[171] ,
         \MC_ARK_ARC_1_4/buf_datainput[170] ,
         \MC_ARK_ARC_1_4/buf_datainput[169] ,
         \MC_ARK_ARC_1_4/buf_datainput[168] ,
         \MC_ARK_ARC_1_4/buf_datainput[167] ,
         \MC_ARK_ARC_1_4/buf_datainput[165] ,
         \MC_ARK_ARC_1_4/buf_datainput[160] ,
         \MC_ARK_ARC_1_4/buf_datainput[154] ,
         \MC_ARK_ARC_1_4/buf_datainput[148] ,
         \MC_ARK_ARC_1_4/buf_datainput[141] ,
         \MC_ARK_ARC_1_4/buf_datainput[135] ,
         \MC_ARK_ARC_1_4/buf_datainput[132] ,
         \MC_ARK_ARC_1_4/buf_datainput[129] ,
         \MC_ARK_ARC_1_4/buf_datainput[120] ,
         \MC_ARK_ARC_1_4/buf_datainput[118] ,
         \MC_ARK_ARC_1_4/buf_datainput[117] ,
         \MC_ARK_ARC_1_4/buf_datainput[108] ,
         \MC_ARK_ARC_1_4/buf_datainput[97] ,
         \MC_ARK_ARC_1_4/buf_datainput[94] ,
         \MC_ARK_ARC_1_4/buf_datainput[93] ,
         \MC_ARK_ARC_1_4/buf_datainput[87] ,
         \MC_ARK_ARC_1_4/buf_datainput[86] ,
         \MC_ARK_ARC_1_4/buf_datainput[77] ,
         \MC_ARK_ARC_1_4/buf_datainput[76] ,
         \MC_ARK_ARC_1_4/buf_datainput[75] ,
         \MC_ARK_ARC_1_4/buf_datainput[73] ,
         \MC_ARK_ARC_1_4/buf_datainput[64] ,
         \MC_ARK_ARC_1_4/buf_datainput[63] ,
         \MC_ARK_ARC_1_4/buf_datainput[55] ,
         \MC_ARK_ARC_1_4/buf_datainput[54] ,
         \MC_ARK_ARC_1_4/buf_datainput[53] ,
         \MC_ARK_ARC_1_4/buf_datainput[45] ,
         \MC_ARK_ARC_1_4/buf_datainput[43] ,
         \MC_ARK_ARC_1_4/buf_datainput[39] ,
         \MC_ARK_ARC_1_4/buf_datainput[27] ,
         \MC_ARK_ARC_1_4/buf_datainput[23] ,
         \MC_ARK_ARC_1_4/buf_datainput[22] ,
         \MC_ARK_ARC_1_4/buf_datainput[18] ,
         \MC_ARK_ARC_1_4/buf_datainput[15] ,
         \MC_ARK_ARC_1_4/buf_datainput[12] , \MC_ARK_ARC_1_4/buf_datainput[9] ,
         \MC_ARK_ARC_1_4/buf_datainput[3] , \MC_ARK_ARC_1_4/buf_datainput[2] ,
         \SB1_0_0/buf_output[5] , \SB1_0_0/buf_output[4] ,
         \SB1_0_0/buf_output[2] , \SB1_0_0/i3[0] , \SB1_0_0/i1_5 ,
         \SB1_0_0/i1_7 , \SB1_0_0/i1[9] , \SB1_0_0/i0_0 , \SB1_0_0/i0_3 ,
         \SB1_0_0/i0_4 , \SB1_0_0/i0[10] , \SB1_0_0/i0[9] , \SB1_0_0/i0[8] ,
         \SB1_0_0/i0[7] , \SB1_0_0/i0[6] , \SB1_0_1/buf_output[5] ,
         \SB1_0_1/buf_output[4] , \SB1_0_1/buf_output[1] , \SB1_0_1/i3[0] ,
         \SB1_0_1/i1_5 , \SB1_0_1/i1_7 , \SB1_0_1/i1[9] , \SB1_0_1/i0_0 ,
         \SB1_0_1/i0_3 , \SB1_0_1/i0_4 , \SB1_0_1/i0[10] , \SB1_0_1/i0[9] ,
         \SB1_0_1/i0[8] , \SB1_0_1/i0[7] , \SB1_0_1/i0[6] ,
         \SB1_0_2/buf_output[2] , \SB1_0_2/buf_output[1] ,
         \SB1_0_2/buf_output[0] , \SB1_0_2/i3[0] , \SB1_0_2/i1_5 ,
         \SB1_0_2/i1_7 , \SB1_0_2/i1[9] , \SB1_0_2/i0_0 , \SB1_0_2/i0_3 ,
         \SB1_0_2/i0_4 , \SB1_0_2/i0[10] , \SB1_0_2/i0[9] , \SB1_0_2/i0[8] ,
         \SB1_0_2/i0[7] , \SB1_0_2/i0[6] , \SB1_0_3/buf_output[4] ,
         \SB1_0_3/buf_output[0] , \SB1_0_3/i3[0] , \SB1_0_3/i1_5 ,
         \SB1_0_3/i1_7 , \SB1_0_3/i1[9] , \SB1_0_3/i0_0 , \SB1_0_3/i0_3 ,
         \SB1_0_3/i0_4 , \SB1_0_3/i0[10] , \SB1_0_3/i0[9] , \SB1_0_3/i0[8] ,
         \SB1_0_3/i0[7] , \SB1_0_3/i0[6] , \SB1_0_4/buf_output[4] ,
         \SB1_0_4/i3[0] , \SB1_0_4/i1_5 , \SB1_0_4/i1_7 , \SB1_0_4/i1[9] ,
         \SB1_0_4/i0_0 , \SB1_0_4/i0_3 , \SB1_0_4/i0_4 , \SB1_0_4/i0[10] ,
         \SB1_0_4/i0[9] , \SB1_0_4/i0[8] , \SB1_0_4/i0[7] , \SB1_0_4/i0[6] ,
         \SB1_0_5/buf_output[5] , \SB1_0_5/buf_output[1] ,
         \SB1_0_5/buf_output[0] , \SB1_0_5/i3[0] , \SB1_0_5/i1_5 ,
         \SB1_0_5/i1_7 , \SB1_0_5/i1[9] , \SB1_0_5/i0_0 , \SB1_0_5/i0_3 ,
         \SB1_0_5/i0_4 , \SB1_0_5/i0[10] , \SB1_0_5/i0[9] , \SB1_0_5/i0[8] ,
         \SB1_0_5/i0[7] , \SB1_0_5/i0[6] , \SB1_0_6/buf_output[3] ,
         \SB1_0_6/i3[0] , \SB1_0_6/i1_5 , \SB1_0_6/i1_7 , \SB1_0_6/i1[9] ,
         \SB1_0_6/i0_0 , \SB1_0_6/i0_3 , \SB1_0_6/i0_4 , \SB1_0_6/i0[10] ,
         \SB1_0_6/i0[9] , \SB1_0_6/i0[8] , \SB1_0_6/i0[7] , \SB1_0_6/i0[6] ,
         \SB1_0_7/buf_output[3] , \SB1_0_7/buf_output[2] , \SB1_0_7/i3[0] ,
         \SB1_0_7/i1_5 , \SB1_0_7/i1_7 , \SB1_0_7/i1[9] , \SB1_0_7/i0_0 ,
         \SB1_0_7/i0_3 , \SB1_0_7/i0_4 , \SB1_0_7/i0[10] , \SB1_0_7/i0[9] ,
         \SB1_0_7/i0[8] , \SB1_0_7/i0[7] , \SB1_0_7/i0[6] ,
         \SB1_0_8/buf_output[4] , \SB1_0_8/buf_output[0] , \SB1_0_8/i3[0] ,
         \SB1_0_8/i1_5 , \SB1_0_8/i1_7 , \SB1_0_8/i1[9] , \SB1_0_8/i0_0 ,
         \SB1_0_8/i0_3 , \SB1_0_8/i0_4 , \SB1_0_8/i0[10] , \SB1_0_8/i0[9] ,
         \SB1_0_8/i0[8] , \SB1_0_8/i0[7] , \SB1_0_8/i0[6] ,
         \SB1_0_9/buf_output[5] , \SB1_0_9/buf_output[4] ,
         \SB1_0_9/buf_output[1] , \SB1_0_9/i3[0] , \SB1_0_9/i1_5 ,
         \SB1_0_9/i1_7 , \SB1_0_9/i1[9] , \SB1_0_9/i0_0 , \SB1_0_9/i0_3 ,
         \SB1_0_9/i0_4 , \SB1_0_9/i0[10] , \SB1_0_9/i0[9] , \SB1_0_9/i0[8] ,
         \SB1_0_9/i0[7] , \SB1_0_9/i0[6] , \SB1_0_10/buf_output[2] ,
         \SB1_0_10/buf_output[0] , \SB1_0_10/i3[0] , \SB1_0_10/i1_5 ,
         \SB1_0_10/i1_7 , \SB1_0_10/i1[9] , \SB1_0_10/i0_0 , \SB1_0_10/i0_3 ,
         \SB1_0_10/i0_4 , \SB1_0_10/i0[10] , \SB1_0_10/i0[9] ,
         \SB1_0_10/i0[8] , \SB1_0_10/i0[7] , \SB1_0_10/i0[6] ,
         \SB1_0_11/buf_output[3] , \SB1_0_11/buf_output[1] , \SB1_0_11/i3[0] ,
         \SB1_0_11/i1_5 , \SB1_0_11/i1_7 , \SB1_0_11/i1[9] , \SB1_0_11/i0_0 ,
         \SB1_0_11/i0_3 , \SB1_0_11/i0_4 , \SB1_0_11/i0[10] , \SB1_0_11/i0[9] ,
         \SB1_0_11/i0[8] , \SB1_0_11/i0[7] , \SB1_0_11/i0[6] ,
         \SB1_0_12/buf_output[5] , \SB1_0_12/buf_output[4] , \SB1_0_12/i3[0] ,
         \SB1_0_12/i1_5 , \SB1_0_12/i1_7 , \SB1_0_12/i1[9] , \SB1_0_12/i0_0 ,
         \SB1_0_12/i0_3 , \SB1_0_12/i0_4 , \SB1_0_12/i0[10] , \SB1_0_12/i0[9] ,
         \SB1_0_12/i0[8] , \SB1_0_12/i0[7] , \SB1_0_12/i0[6] ,
         \SB1_0_13/buf_output[4] , \SB1_0_13/buf_output[0] , \SB1_0_13/i3[0] ,
         \SB1_0_13/i1_5 , \SB1_0_13/i1_7 , \SB1_0_13/i1[9] , \SB1_0_13/i0_0 ,
         \SB1_0_13/i0_3 , \SB1_0_13/i0_4 , \SB1_0_13/i0[10] , \SB1_0_13/i0[9] ,
         \SB1_0_13/i0[8] , \SB1_0_13/i0[7] , \SB1_0_13/i0[6] ,
         \SB1_0_14/buf_output[5] , \SB1_0_14/buf_output[4] , \SB1_0_14/i3[0] ,
         \SB1_0_14/i1_5 , \SB1_0_14/i1_7 , \SB1_0_14/i1[9] , \SB1_0_14/i0_0 ,
         \SB1_0_14/i0_3 , \SB1_0_14/i0_4 , \SB1_0_14/i0[10] , \SB1_0_14/i0[9] ,
         \SB1_0_14/i0[8] , \SB1_0_14/i0[7] , \SB1_0_14/i0[6] ,
         \SB1_0_15/i3[0] , \SB1_0_15/i1_5 , \SB1_0_15/i1_7 , \SB1_0_15/i1[9] ,
         \SB1_0_15/i0_0 , \SB1_0_15/i0_3 , \SB1_0_15/i0_4 , \SB1_0_15/i0[10] ,
         \SB1_0_15/i0[9] , \SB1_0_15/i0[8] , \SB1_0_15/i0[7] ,
         \SB1_0_15/i0[6] , \SB1_0_16/buf_output[3] , \SB1_0_16/i3[0] ,
         \SB1_0_16/i1_5 , \SB1_0_16/i1_7 , \SB1_0_16/i1[9] , \SB1_0_16/i0_0 ,
         \SB1_0_16/i0_3 , \SB1_0_16/i0_4 , \SB1_0_16/i0[10] , \SB1_0_16/i0[9] ,
         \SB1_0_16/i0[8] , \SB1_0_16/i0[7] , \SB1_0_16/i0[6] ,
         \SB1_0_17/buf_output[2] , \SB1_0_17/i3[0] , \SB1_0_17/i1_5 ,
         \SB1_0_17/i1_7 , \SB1_0_17/i1[9] , \SB1_0_17/i0_0 , \SB1_0_17/i0_3 ,
         \SB1_0_17/i0_4 , \SB1_0_17/i0[10] , \SB1_0_17/i0[9] ,
         \SB1_0_17/i0[8] , \SB1_0_17/i0[7] , \SB1_0_17/i0[6] ,
         \SB1_0_18/buf_output[3] , \SB1_0_18/buf_output[2] ,
         \SB1_0_18/buf_output[0] , \SB1_0_18/i3[0] , \SB1_0_18/i1_5 ,
         \SB1_0_18/i1_7 , \SB1_0_18/i1[9] , \SB1_0_18/i0_3 , \SB1_0_18/i0_4 ,
         \SB1_0_18/i0[10] , \SB1_0_18/i0[9] , \SB1_0_18/i0[8] ,
         \SB1_0_18/i0[7] , \SB1_0_18/i0[6] , \SB1_0_19/buf_output[4] ,
         \SB1_0_19/buf_output[2] , \SB1_0_19/i3[0] , \SB1_0_19/i1_5 ,
         \SB1_0_19/i1_7 , \SB1_0_19/i1[9] , \SB1_0_19/i0_0 , \SB1_0_19/i0_3 ,
         \SB1_0_19/i0_4 , \SB1_0_19/i0[10] , \SB1_0_19/i0[9] ,
         \SB1_0_19/i0[8] , \SB1_0_19/i0[7] , \SB1_0_19/i0[6] ,
         \SB1_0_20/buf_output[5] , \SB1_0_20/buf_output[4] , \SB1_0_20/i3[0] ,
         \SB1_0_20/i1_5 , \SB1_0_20/i1_7 , \SB1_0_20/i1[9] , \SB1_0_20/i0_0 ,
         \SB1_0_20/i0_3 , \SB1_0_20/i0_4 , \SB1_0_20/i0[10] , \SB1_0_20/i0[9] ,
         \SB1_0_20/i0[8] , \SB1_0_20/i0[7] , \SB1_0_20/i0[6] ,
         \SB1_0_21/buf_output[4] , \SB1_0_21/buf_output[3] ,
         \SB1_0_21/buf_output[2] , \SB1_0_21/buf_output[1] , \SB1_0_21/i3[0] ,
         \SB1_0_21/i1_5 , \SB1_0_21/i1_7 , \SB1_0_21/i1[9] , \SB1_0_21/i0_0 ,
         \SB1_0_21/i0_3 , \SB1_0_21/i0_4 , \SB1_0_21/i0[10] , \SB1_0_21/i0[9] ,
         \SB1_0_21/i0[8] , \SB1_0_21/i0[7] , \SB1_0_21/i0[6] ,
         \SB1_0_22/buf_output[5] , \SB1_0_22/buf_output[4] ,
         \SB1_0_22/buf_output[3] , \SB1_0_22/buf_output[2] ,
         \SB1_0_22/buf_output[1] , \SB1_0_22/buf_output[0] , \SB1_0_22/i3[0] ,
         \SB1_0_22/i1_5 , \SB1_0_22/i1_7 , \SB1_0_22/i1[9] , \SB1_0_22/i0_0 ,
         \SB1_0_22/i0_3 , \SB1_0_22/i0_4 , \SB1_0_22/i0[10] , \SB1_0_22/i0[9] ,
         \SB1_0_22/i0[8] , \SB1_0_22/i0[7] , \SB1_0_22/i0[6] ,
         \SB1_0_23/buf_output[4] , \SB1_0_23/buf_output[1] , \SB1_0_23/i3[0] ,
         \SB1_0_23/i1_5 , \SB1_0_23/i1_7 , \SB1_0_23/i1[9] , \SB1_0_23/i0_0 ,
         \SB1_0_23/i0_3 , \SB1_0_23/i0_4 , \SB1_0_23/i0[10] , \SB1_0_23/i0[9] ,
         \SB1_0_23/i0[8] , \SB1_0_23/i0[7] , \SB1_0_23/i0[6] ,
         \SB1_0_24/buf_output[4] , \SB1_0_24/buf_output[3] ,
         \SB1_0_24/buf_output[2] , \SB1_0_24/i3[0] , \SB1_0_24/i1_5 ,
         \SB1_0_24/i1_7 , \SB1_0_24/i1[9] , \SB1_0_24/i0_0 , \SB1_0_24/i0_3 ,
         \SB1_0_24/i0_4 , \SB1_0_24/i0[10] , \SB1_0_24/i0[9] ,
         \SB1_0_24/i0[8] , \SB1_0_24/i0[7] , \SB1_0_24/i0[6] ,
         \SB1_0_25/buf_output[3] , \SB1_0_25/buf_output[1] ,
         \SB1_0_25/buf_output[0] , \SB1_0_25/i3[0] , \SB1_0_25/i1_5 ,
         \SB1_0_25/i1_7 , \SB1_0_25/i1[9] , \SB1_0_25/i0_0 , \SB1_0_25/i0_3 ,
         \SB1_0_25/i0_4 , \SB1_0_25/i0[10] , \SB1_0_25/i0[9] ,
         \SB1_0_25/i0[8] , \SB1_0_25/i0[7] , \SB1_0_25/i0[6] ,
         \SB1_0_26/buf_output[3] , \SB1_0_26/buf_output[1] , \SB1_0_26/i3[0] ,
         \SB1_0_26/i1_5 , \SB1_0_26/i1_7 , \SB1_0_26/i1[9] , \SB1_0_26/i0_0 ,
         \SB1_0_26/i0_3 , \SB1_0_26/i0_4 , \SB1_0_26/i0[10] , \SB1_0_26/i0[9] ,
         \SB1_0_26/i0[8] , \SB1_0_26/i0[7] , \SB1_0_26/i0[6] ,
         \SB1_0_27/buf_output[1] , \SB1_0_27/buf_output[0] , \SB1_0_27/i3[0] ,
         \SB1_0_27/i1_5 , \SB1_0_27/i1_7 , \SB1_0_27/i1[9] , \SB1_0_27/i0_0 ,
         \SB1_0_27/i0_3 , \SB1_0_27/i0_4 , \SB1_0_27/i0[10] , \SB1_0_27/i0[9] ,
         \SB1_0_27/i0[8] , \SB1_0_27/i0[7] , \SB1_0_27/i0[6] ,
         \SB1_0_28/buf_output[5] , \SB1_0_28/buf_output[4] ,
         \SB1_0_28/buf_output[3] , \SB1_0_28/buf_output[1] ,
         \SB1_0_28/buf_output[0] , \SB1_0_28/i3[0] , \SB1_0_28/i1_5 ,
         \SB1_0_28/i1_7 , \SB1_0_28/i1[9] , \SB1_0_28/i0_0 , \SB1_0_28/i0_3 ,
         \SB1_0_28/i0[10] , \SB1_0_28/i0[9] , \SB1_0_28/i0[8] ,
         \SB1_0_28/i0[7] , \SB1_0_28/i0[6] , \SB1_0_29/buf_output[5] ,
         \SB1_0_29/buf_output[2] , \SB1_0_29/buf_output[1] ,
         \SB1_0_29/buf_output[0] , \SB1_0_29/i3[0] , \SB1_0_29/i1_5 ,
         \SB1_0_29/i1_7 , \SB1_0_29/i1[9] , \SB1_0_29/i0_0 , \SB1_0_29/i0_3 ,
         \SB1_0_29/i0_4 , \SB1_0_29/i0[10] , \SB1_0_29/i0[9] ,
         \SB1_0_29/i0[8] , \SB1_0_29/i0[7] , \SB1_0_29/i0[6] ,
         \SB1_0_30/buf_output[5] , \SB1_0_30/buf_output[2] ,
         \SB1_0_30/buf_output[1] , \SB1_0_30/buf_output[0] , \SB1_0_30/i3[0] ,
         \SB1_0_30/i1_5 , \SB1_0_30/i1_7 , \SB1_0_30/i1[9] , \SB1_0_30/i0_0 ,
         \SB1_0_30/i0_3 , \SB1_0_30/i0_4 , \SB1_0_30/i0[10] , \SB1_0_30/i0[9] ,
         \SB1_0_30/i0[8] , \SB1_0_30/i0[7] , \SB1_0_30/i0[6] ,
         \SB1_0_31/buf_output[2] , \SB1_0_31/buf_output[1] , \SB1_0_31/i3[0] ,
         \SB1_0_31/i1_5 , \SB1_0_31/i1_7 , \SB1_0_31/i1[9] , \SB1_0_31/i0_0 ,
         \SB1_0_31/i0_3 , \SB1_0_31/i0_4 , \SB1_0_31/i0[10] , \SB1_0_31/i0[9] ,
         \SB1_0_31/i0[8] , \SB1_0_31/i0[7] , \SB1_0_31/i0[6] ,
         \SB2_0_0/buf_output[5] , \SB2_0_0/buf_output[4] ,
         \SB2_0_0/buf_output[3] , \SB2_0_0/buf_output[2] ,
         \SB2_0_0/buf_output[1] , \SB2_0_0/buf_output[0] , \SB2_0_0/i3[0] ,
         \SB2_0_0/i1_5 , \SB2_0_0/i1_7 , \SB2_0_0/i1[9] , \SB2_0_0/i0_0 ,
         \SB2_0_0/i0_3 , \SB2_0_0/i0[10] , \SB2_0_0/i0[9] , \SB2_0_0/i0[7] ,
         \SB2_0_0/i0[6] , \SB2_0_1/buf_output[5] , \SB2_0_1/buf_output[4] ,
         \SB2_0_1/buf_output[3] , \SB2_0_1/buf_output[2] ,
         \SB2_0_1/buf_output[1] , \SB2_0_1/buf_output[0] , \SB2_0_1/i1_5 ,
         \SB2_0_1/i1_7 , \SB2_0_1/i1[9] , \SB2_0_1/i0_0 , \SB2_0_1/i0_3 ,
         \SB2_0_1/i0_4 , \SB2_0_1/i0[10] , \SB2_0_1/i0[9] , \SB2_0_1/i0[8] ,
         \SB2_0_1/i0[7] , \SB2_0_1/i0[6] , \SB2_0_2/buf_output[5] ,
         \SB2_0_2/buf_output[4] , \SB2_0_2/buf_output[3] ,
         \SB2_0_2/buf_output[2] , \SB2_0_2/buf_output[1] ,
         \SB2_0_2/buf_output[0] , \SB2_0_2/i3[0] , \SB2_0_2/i1_5 ,
         \SB2_0_2/i1_7 , \SB2_0_2/i1[9] , \SB2_0_2/i0_0 , \SB2_0_2/i0_3 ,
         \SB2_0_2/i0[10] , \SB2_0_2/i0[9] , \SB2_0_2/i0[8] , \SB2_0_2/i0[7] ,
         \SB2_0_2/i0[6] , \SB2_0_3/buf_output[4] , \SB2_0_3/buf_output[3] ,
         \SB2_0_3/buf_output[2] , \SB2_0_3/buf_output[1] ,
         \SB2_0_3/buf_output[0] , \SB2_0_3/i3[0] , \SB2_0_3/i1_5 ,
         \SB2_0_3/i1_7 , \SB2_0_3/i1[9] , \SB2_0_3/i0_0 , \SB2_0_3/i0_3 ,
         \SB2_0_3/i0[10] , \SB2_0_3/i0[9] , \SB2_0_3/i0[8] , \SB2_0_3/i0[7] ,
         \SB2_0_3/i0[6] , \SB2_0_4/buf_output[5] , \SB2_0_4/buf_output[4] ,
         \SB2_0_4/buf_output[3] , \SB2_0_4/buf_output[2] ,
         \SB2_0_4/buf_output[1] , \SB2_0_4/buf_output[0] , \SB2_0_4/i1_5 ,
         \SB2_0_4/i1_7 , \SB2_0_4/i1[9] , \SB2_0_4/i0_0 , \SB2_0_4/i0_3 ,
         \SB2_0_4/i0[10] , \SB2_0_4/i0[9] , \SB2_0_4/i0[8] , \SB2_0_4/i0[7] ,
         \SB2_0_4/i0[6] , \SB2_0_5/buf_output[5] , \SB2_0_5/buf_output[4] ,
         \SB2_0_5/buf_output[3] , \SB2_0_5/buf_output[2] ,
         \SB2_0_5/buf_output[1] , \SB2_0_5/buf_output[0] , \SB2_0_5/i3[0] ,
         \SB2_0_5/i1_7 , \SB2_0_5/i1[9] , \SB2_0_5/i0_0 , \SB2_0_5/i0_3 ,
         \SB2_0_5/i0_4 , \SB2_0_5/i0[10] , \SB2_0_5/i0[9] , \SB2_0_5/i0[8] ,
         \SB2_0_5/i0[6] , \SB2_0_6/buf_output[5] , \SB2_0_6/buf_output[4] ,
         \SB2_0_6/buf_output[3] , \SB2_0_6/buf_output[2] ,
         \SB2_0_6/buf_output[1] , \SB2_0_6/buf_output[0] , \SB2_0_6/i3[0] ,
         \SB2_0_6/i1_5 , \SB2_0_6/i1_7 , \SB2_0_6/i1[9] , \SB2_0_6/i0_0 ,
         \SB2_0_6/i0_3 , \SB2_0_6/i0_4 , \SB2_0_6/i0[10] , \SB2_0_6/i0[9] ,
         \SB2_0_6/i0[8] , \SB2_0_6/i0[7] , \SB2_0_6/i0[6] ,
         \SB2_0_7/buf_output[4] , \SB2_0_7/buf_output[3] ,
         \SB2_0_7/buf_output[2] , \SB2_0_7/buf_output[1] ,
         \SB2_0_7/buf_output[0] , \SB2_0_7/i3[0] , \SB2_0_7/i1_5 ,
         \SB2_0_7/i1_7 , \SB2_0_7/i1[9] , \SB2_0_7/i0_0 , \SB2_0_7/i0_3 ,
         \SB2_0_7/i0[10] , \SB2_0_7/i0[9] , \SB2_0_7/i0[8] , \SB2_0_7/i0[7] ,
         \SB2_0_7/i0[6] , \SB2_0_8/buf_output[5] , \SB2_0_8/buf_output[4] ,
         \SB2_0_8/buf_output[3] , \SB2_0_8/buf_output[2] ,
         \SB2_0_8/buf_output[1] , \SB2_0_8/buf_output[0] , \SB2_0_8/i3[0] ,
         \SB2_0_8/i1_5 , \SB2_0_8/i1_7 , \SB2_0_8/i1[9] , \SB2_0_8/i0_0 ,
         \SB2_0_8/i0_3 , \SB2_0_8/i0[10] , \SB2_0_8/i0[9] , \SB2_0_8/i0[8] ,
         \SB2_0_8/i0[7] , \SB2_0_8/i0[6] , \SB2_0_9/buf_output[5] ,
         \SB2_0_9/buf_output[4] , \SB2_0_9/buf_output[3] ,
         \SB2_0_9/buf_output[2] , \SB2_0_9/buf_output[1] ,
         \SB2_0_9/buf_output[0] , \SB2_0_9/i3[0] , \SB2_0_9/i1_5 ,
         \SB2_0_9/i1_7 , \SB2_0_9/i1[9] , \SB2_0_9/i0_0 , \SB2_0_9/i0_3 ,
         \SB2_0_9/i0_4 , \SB2_0_9/i0[10] , \SB2_0_9/i0[9] , \SB2_0_9/i0[8] ,
         \SB2_0_9/i0[7] , \SB2_0_9/i0[6] , \SB2_0_10/buf_output[5] ,
         \SB2_0_10/buf_output[4] , \SB2_0_10/buf_output[3] ,
         \SB2_0_10/buf_output[2] , \SB2_0_10/buf_output[1] ,
         \SB2_0_10/buf_output[0] , \SB2_0_10/i3[0] , \SB2_0_10/i1_5 ,
         \SB2_0_10/i1_7 , \SB2_0_10/i1[9] , \SB2_0_10/i0_3 , \SB2_0_10/i0_4 ,
         \SB2_0_10/i0[10] , \SB2_0_10/i0[9] , \SB2_0_10/i0[8] ,
         \SB2_0_10/i0[6] , \SB2_0_11/buf_output[5] , \SB2_0_11/buf_output[4] ,
         \SB2_0_11/buf_output[3] , \SB2_0_11/buf_output[2] ,
         \SB2_0_11/buf_output[1] , \SB2_0_11/buf_output[0] , \SB2_0_11/i3[0] ,
         \SB2_0_11/i1_5 , \SB2_0_11/i1_7 , \SB2_0_11/i1[9] , \SB2_0_11/i0_0 ,
         \SB2_0_11/i0_3 , \SB2_0_11/i0_4 , \SB2_0_11/i0[10] , \SB2_0_11/i0[9] ,
         \SB2_0_11/i0[8] , \SB2_0_11/i0[7] , \SB2_0_11/i0[6] ,
         \SB2_0_12/buf_output[5] , \SB2_0_12/buf_output[4] ,
         \SB2_0_12/buf_output[3] , \SB2_0_12/buf_output[2] ,
         \SB2_0_12/buf_output[1] , \SB2_0_12/buf_output[0] , \SB2_0_12/i3[0] ,
         \SB2_0_12/i1_5 , \SB2_0_12/i1_7 , \SB2_0_12/i1[9] , \SB2_0_12/i0_0 ,
         \SB2_0_12/i0[10] , \SB2_0_12/i0[9] , \SB2_0_12/i0[8] ,
         \SB2_0_12/i0[7] , \SB2_0_12/i0[6] , \SB2_0_13/buf_output[5] ,
         \SB2_0_13/buf_output[4] , \SB2_0_13/buf_output[3] ,
         \SB2_0_13/buf_output[2] , \SB2_0_13/buf_output[1] ,
         \SB2_0_13/buf_output[0] , \SB2_0_13/i3[0] , \SB2_0_13/i1_5 ,
         \SB2_0_13/i1_7 , \SB2_0_13/i1[9] , \SB2_0_13/i0_0 , \SB2_0_13/i0_3 ,
         \SB2_0_13/i0[10] , \SB2_0_13/i0[9] , \SB2_0_13/i0[8] ,
         \SB2_0_13/i0[7] , \SB2_0_13/i0[6] , \SB2_0_14/buf_output[5] ,
         \SB2_0_14/buf_output[4] , \SB2_0_14/buf_output[3] ,
         \SB2_0_14/buf_output[2] , \SB2_0_14/buf_output[1] ,
         \SB2_0_14/buf_output[0] , \SB2_0_14/i3[0] , \SB2_0_14/i1_5 ,
         \SB2_0_14/i1_7 , \SB2_0_14/i1[9] , \SB2_0_14/i0_0 , \SB2_0_14/i0_3 ,
         \SB2_0_14/i0_4 , \SB2_0_14/i0[10] , \SB2_0_14/i0[9] ,
         \SB2_0_14/i0[8] , \SB2_0_14/i0[6] , \SB2_0_15/buf_output[5] ,
         \SB2_0_15/buf_output[4] , \SB2_0_15/buf_output[3] ,
         \SB2_0_15/buf_output[2] , \SB2_0_15/buf_output[0] , \SB2_0_15/i3[0] ,
         \SB2_0_15/i1_5 , \SB2_0_15/i1_7 , \SB2_0_15/i0_3 , \SB2_0_15/i0[10] ,
         \SB2_0_15/i0[9] , \SB2_0_15/i0[8] , \SB2_0_15/i0[7] ,
         \SB2_0_15/i0[6] , \SB2_0_16/buf_output[5] , \SB2_0_16/buf_output[4] ,
         \SB2_0_16/buf_output[3] , \SB2_0_16/buf_output[2] ,
         \SB2_0_16/buf_output[1] , \SB2_0_16/buf_output[0] , \SB2_0_16/i3[0] ,
         \SB2_0_16/i1_5 , \SB2_0_16/i1_7 , \SB2_0_16/i1[9] , \SB2_0_16/i0_0 ,
         \SB2_0_16/i0_3 , \SB2_0_16/i0[9] , \SB2_0_16/i0[8] , \SB2_0_16/i0[7] ,
         \SB2_0_16/i0[6] , \SB2_0_17/buf_output[5] , \SB2_0_17/buf_output[4] ,
         \SB2_0_17/buf_output[3] , \SB2_0_17/buf_output[2] ,
         \SB2_0_17/buf_output[1] , \SB2_0_17/buf_output[0] , \SB2_0_17/i3[0] ,
         \SB2_0_17/i1_5 , \SB2_0_17/i1_7 , \SB2_0_17/i1[9] , \SB2_0_17/i0_0 ,
         \SB2_0_17/i0_3 , \SB2_0_17/i0[10] , \SB2_0_17/i0[9] ,
         \SB2_0_17/i0[8] , \SB2_0_17/i0[7] , \SB2_0_17/i0[6] ,
         \SB2_0_18/buf_output[5] , \SB2_0_18/buf_output[4] ,
         \SB2_0_18/buf_output[3] , \SB2_0_18/buf_output[2] ,
         \SB2_0_18/buf_output[1] , \SB2_0_18/buf_output[0] , \SB2_0_18/i3[0] ,
         \SB2_0_18/i1_5 , \SB2_0_18/i1_7 , \SB2_0_18/i1[9] , \SB2_0_18/i0_0 ,
         \SB2_0_18/i0_3 , \SB2_0_18/i0[10] , \SB2_0_18/i0[9] ,
         \SB2_0_18/i0[8] , \SB2_0_18/i0[7] , \SB2_0_18/i0[6] ,
         \SB2_0_19/buf_output[5] , \SB2_0_19/buf_output[4] ,
         \SB2_0_19/buf_output[3] , \SB2_0_19/buf_output[2] ,
         \SB2_0_19/buf_output[1] , \SB2_0_19/buf_output[0] , \SB2_0_19/i3[0] ,
         \SB2_0_19/i1_5 , \SB2_0_19/i1_7 , \SB2_0_19/i1[9] , \SB2_0_19/i0_0 ,
         \SB2_0_19/i0[9] , \SB2_0_19/i0[8] , \SB2_0_19/i0[7] ,
         \SB2_0_19/i0[6] , \SB2_0_20/buf_output[5] , \SB2_0_20/buf_output[4] ,
         \SB2_0_20/buf_output[3] , \SB2_0_20/buf_output[2] ,
         \SB2_0_20/buf_output[1] , \SB2_0_20/buf_output[0] , \SB2_0_20/i3[0] ,
         \SB2_0_20/i1_5 , \SB2_0_20/i1_7 , \SB2_0_20/i1[9] , \SB2_0_20/i0_0 ,
         \SB2_0_20/i0_3 , \SB2_0_20/i0[10] , \SB2_0_20/i0[9] ,
         \SB2_0_20/i0[8] , \SB2_0_20/i0[7] , \SB2_0_20/i0[6] ,
         \SB2_0_21/buf_output[5] , \SB2_0_21/buf_output[4] ,
         \SB2_0_21/buf_output[3] , \SB2_0_21/buf_output[2] ,
         \SB2_0_21/buf_output[1] , \SB2_0_21/buf_output[0] , \SB2_0_21/i3[0] ,
         \SB2_0_21/i1_5 , \SB2_0_21/i1_7 , \SB2_0_21/i1[9] , \SB2_0_21/i0_0 ,
         \SB2_0_21/i0_3 , \SB2_0_21/i0_4 , \SB2_0_21/i0[10] , \SB2_0_21/i0[9] ,
         \SB2_0_21/i0[8] , \SB2_0_21/i0[7] , \SB2_0_21/i0[6] ,
         \SB2_0_22/buf_output[5] , \SB2_0_22/buf_output[4] ,
         \SB2_0_22/buf_output[3] , \SB2_0_22/buf_output[2] ,
         \SB2_0_22/buf_output[1] , \SB2_0_22/buf_output[0] , \SB2_0_22/i3[0] ,
         \SB2_0_22/i1_5 , \SB2_0_22/i1_7 , \SB2_0_22/i1[9] , \SB2_0_22/i0_0 ,
         \SB2_0_22/i0_3 , \SB2_0_22/i0[10] , \SB2_0_22/i0[9] ,
         \SB2_0_22/i0[8] , \SB2_0_22/i0[7] , \SB2_0_23/buf_output[5] ,
         \SB2_0_23/buf_output[4] , \SB2_0_23/buf_output[3] ,
         \SB2_0_23/buf_output[2] , \SB2_0_23/buf_output[1] ,
         \SB2_0_23/buf_output[0] , \SB2_0_23/i3[0] , \SB2_0_23/i1_5 ,
         \SB2_0_23/i1_7 , \SB2_0_23/i1[9] , \SB2_0_23/i0_0 , \SB2_0_23/i0_3 ,
         \SB2_0_23/i0[10] , \SB2_0_23/i0[9] , \SB2_0_23/i0[8] ,
         \SB2_0_23/i0[7] , \SB2_0_23/i0[6] , \SB2_0_24/buf_output[5] ,
         \SB2_0_24/buf_output[4] , \SB2_0_24/buf_output[3] ,
         \SB2_0_24/buf_output[2] , \SB2_0_24/buf_output[1] ,
         \SB2_0_24/buf_output[0] , \SB2_0_24/i3[0] , \SB2_0_24/i1_5 ,
         \SB2_0_24/i1_7 , \SB2_0_24/i1[9] , \SB2_0_24/i0_0 , \SB2_0_24/i0_3 ,
         \SB2_0_24/i0[10] , \SB2_0_24/i0[8] , \SB2_0_24/i0[7] ,
         \SB2_0_24/i0[6] , \SB2_0_25/buf_output[5] , \SB2_0_25/buf_output[4] ,
         \SB2_0_25/buf_output[3] , \SB2_0_25/buf_output[2] ,
         \SB2_0_25/buf_output[1] , \SB2_0_25/buf_output[0] , \SB2_0_25/i3[0] ,
         \SB2_0_25/i1_5 , \SB2_0_25/i1_7 , \SB2_0_25/i1[9] , \SB2_0_25/i0_0 ,
         \SB2_0_25/i0_3 , \SB2_0_25/i0_4 , \SB2_0_25/i0[10] , \SB2_0_25/i0[9] ,
         \SB2_0_25/i0[8] , \SB2_0_25/i0[6] , \SB2_0_26/buf_output[5] ,
         \SB2_0_26/buf_output[4] , \SB2_0_26/buf_output[3] ,
         \SB2_0_26/buf_output[2] , \SB2_0_26/buf_output[1] ,
         \SB2_0_26/buf_output[0] , \SB2_0_26/i3[0] , \SB2_0_26/i1_5 ,
         \SB2_0_26/i1_7 , \SB2_0_26/i1[9] , \SB2_0_26/i0_0 , \SB2_0_26/i0_3 ,
         \SB2_0_26/i0_4 , \SB2_0_26/i0[9] , \SB2_0_26/i0[8] , \SB2_0_26/i0[6] ,
         \SB2_0_27/buf_output[5] , \SB2_0_27/buf_output[4] ,
         \SB2_0_27/buf_output[3] , \SB2_0_27/buf_output[2] ,
         \SB2_0_27/buf_output[1] , \SB2_0_27/buf_output[0] , \SB2_0_27/i3[0] ,
         \SB2_0_27/i1_5 , \SB2_0_27/i1_7 , \SB2_0_27/i1[9] , \SB2_0_27/i0_0 ,
         \SB2_0_27/i0_3 , \SB2_0_27/i0[10] , \SB2_0_27/i0[9] ,
         \SB2_0_27/i0[8] , \SB2_0_27/i0[7] , \SB2_0_27/i0[6] ,
         \SB2_0_28/buf_output[5] , \SB2_0_28/buf_output[4] ,
         \SB2_0_28/buf_output[3] , \SB2_0_28/buf_output[2] ,
         \SB2_0_28/buf_output[1] , \SB2_0_28/buf_output[0] , \SB2_0_28/i3[0] ,
         \SB2_0_28/i1_5 , \SB2_0_28/i1_7 , \SB2_0_28/i1[9] , \SB2_0_28/i0_0 ,
         \SB2_0_28/i0_3 , \SB2_0_28/i0_4 , \SB2_0_28/i0[10] , \SB2_0_28/i0[9] ,
         \SB2_0_28/i0[8] , \SB2_0_28/i0[7] , \SB2_0_28/i0[6] ,
         \SB2_0_29/buf_output[5] , \SB2_0_29/buf_output[4] ,
         \SB2_0_29/buf_output[3] , \SB2_0_29/buf_output[2] ,
         \SB2_0_29/buf_output[1] , \SB2_0_29/buf_output[0] , \SB2_0_29/i3[0] ,
         \SB2_0_29/i1_5 , \SB2_0_29/i1_7 , \SB2_0_29/i1[9] , \SB2_0_29/i0_0 ,
         \SB2_0_29/i0_3 , \SB2_0_29/i0_4 , \SB2_0_29/i0[10] , \SB2_0_29/i0[9] ,
         \SB2_0_29/i0[8] , \SB2_0_29/i0[6] , \SB2_0_30/buf_output[5] ,
         \SB2_0_30/buf_output[4] , \SB2_0_30/buf_output[3] ,
         \SB2_0_30/buf_output[2] , \SB2_0_30/buf_output[1] ,
         \SB2_0_30/buf_output[0] , \SB2_0_30/i3[0] , \SB2_0_30/i1_5 ,
         \SB2_0_30/i1_7 , \SB2_0_30/i1[9] , \SB2_0_30/i0_0 , \SB2_0_30/i0_3 ,
         \SB2_0_30/i0_4 , \SB2_0_30/i0[10] , \SB2_0_30/i0[9] ,
         \SB2_0_30/i0[8] , \SB2_0_30/i0[7] , \SB2_0_30/i0[6] ,
         \SB2_0_31/buf_output[5] , \SB2_0_31/buf_output[4] ,
         \SB2_0_31/buf_output[3] , \SB2_0_31/buf_output[2] ,
         \SB2_0_31/buf_output[1] , \SB2_0_31/buf_output[0] , \SB2_0_31/i3[0] ,
         \SB2_0_31/i1_5 , \SB2_0_31/i1_7 , \SB2_0_31/i1[9] , \SB2_0_31/i0_0 ,
         \SB2_0_31/i0_3 , \SB2_0_31/i0[10] , \SB2_0_31/i0[9] ,
         \SB2_0_31/i0[8] , \SB2_0_31/i0[7] , \SB2_0_31/i0[6] ,
         \SB1_1_0/buf_output[5] , \SB1_1_0/buf_output[3] ,
         \SB1_1_0/buf_output[2] , \SB1_1_0/buf_output[1] ,
         \SB1_1_0/buf_output[0] , \SB1_1_0/i3[0] , \SB1_1_0/i1_5 ,
         \SB1_1_0/i1_7 , \SB1_1_0/i1[9] , \SB1_1_0/i0_0 , \SB1_1_0/i0_3 ,
         \SB1_1_0/i0_4 , \SB1_1_0/i0[10] , \SB1_1_0/i0[9] , \SB1_1_0/i0[8] ,
         \SB1_1_0/i0[7] , \SB1_1_0/i0[6] , \SB1_1_1/buf_output[5] ,
         \SB1_1_1/buf_output[3] , \SB1_1_1/buf_output[2] ,
         \SB1_1_1/buf_output[1] , \SB1_1_1/buf_output[0] , \SB1_1_1/i3[0] ,
         \SB1_1_1/i1_5 , \SB1_1_1/i1_7 , \SB1_1_1/i1[9] , \SB1_1_1/i0_0 ,
         \SB1_1_1/i0_3 , \SB1_1_1/i0_4 , \SB1_1_1/i0[10] , \SB1_1_1/i0[9] ,
         \SB1_1_1/i0[8] , \SB1_1_1/i0[7] , \SB1_1_1/i0[6] ,
         \SB1_1_2/buf_output[5] , \SB1_1_2/buf_output[4] ,
         \SB1_1_2/buf_output[3] , \SB1_1_2/buf_output[2] ,
         \SB1_1_2/buf_output[1] , \SB1_1_2/buf_output[0] , \SB1_1_2/i3[0] ,
         \SB1_1_2/i1_5 , \SB1_1_2/i1_7 , \SB1_1_2/i1[9] , \SB1_1_2/i0_0 ,
         \SB1_1_2/i0_3 , \SB1_1_2/i0_4 , \SB1_1_2/i0[10] , \SB1_1_2/i0[9] ,
         \SB1_1_2/i0[8] , \SB1_1_2/i0[7] , \SB1_1_2/i0[6] ,
         \SB1_1_3/buf_output[5] , \SB1_1_3/buf_output[3] ,
         \SB1_1_3/buf_output[2] , \SB1_1_3/buf_output[1] ,
         \SB1_1_3/buf_output[0] , \SB1_1_3/i3[0] , \SB1_1_3/i1_5 ,
         \SB1_1_3/i1_7 , \SB1_1_3/i1[9] , \SB1_1_3/i0_0 , \SB1_1_3/i0_3 ,
         \SB1_1_3/i0_4 , \SB1_1_3/i0[10] , \SB1_1_3/i0[9] , \SB1_1_3/i0[8] ,
         \SB1_1_3/i0[7] , \SB1_1_3/i0[6] , \SB1_1_4/buf_output[5] ,
         \SB1_1_4/buf_output[4] , \SB1_1_4/buf_output[3] ,
         \SB1_1_4/buf_output[2] , \SB1_1_4/buf_output[1] ,
         \SB1_1_4/buf_output[0] , \SB1_1_4/i3[0] , \SB1_1_4/i1_5 ,
         \SB1_1_4/i1_7 , \SB1_1_4/i1[9] , \SB1_1_4/i0_0 , \SB1_1_4/i0_3 ,
         \SB1_1_4/i0_4 , \SB1_1_4/i0[10] , \SB1_1_4/i0[9] , \SB1_1_4/i0[8] ,
         \SB1_1_4/i0[7] , \SB1_1_4/i0[6] , \SB1_1_5/buf_output[5] ,
         \SB1_1_5/buf_output[4] , \SB1_1_5/buf_output[3] ,
         \SB1_1_5/buf_output[2] , \SB1_1_5/buf_output[1] ,
         \SB1_1_5/buf_output[0] , \SB1_1_5/i3[0] , \SB1_1_5/i1_5 ,
         \SB1_1_5/i1_7 , \SB1_1_5/i1[9] , \SB1_1_5/i0_0 , \SB1_1_5/i0_3 ,
         \SB1_1_5/i0_4 , \SB1_1_5/i0[10] , \SB1_1_5/i0[9] , \SB1_1_5/i0[8] ,
         \SB1_1_5/i0[7] , \SB1_1_5/i0[6] , \SB1_1_6/buf_output[5] ,
         \SB1_1_6/buf_output[4] , \SB1_1_6/buf_output[3] ,
         \SB1_1_6/buf_output[2] , \SB1_1_6/buf_output[1] ,
         \SB1_1_6/buf_output[0] , \SB1_1_6/i3[0] , \SB1_1_6/i1_5 ,
         \SB1_1_6/i1_7 , \SB1_1_6/i1[9] , \SB1_1_6/i0_0 , \SB1_1_6/i0_3 ,
         \SB1_1_6/i0_4 , \SB1_1_6/i0[10] , \SB1_1_6/i0[9] , \SB1_1_6/i0[8] ,
         \SB1_1_6/i0[7] , \SB1_1_6/i0[6] , \SB1_1_7/buf_output[5] ,
         \SB1_1_7/buf_output[4] , \SB1_1_7/buf_output[3] ,
         \SB1_1_7/buf_output[2] , \SB1_1_7/buf_output[1] ,
         \SB1_1_7/buf_output[0] , \SB1_1_7/i3[0] , \SB1_1_7/i1_5 ,
         \SB1_1_7/i1_7 , \SB1_1_7/i1[9] , \SB1_1_7/i0_0 , \SB1_1_7/i0_3 ,
         \SB1_1_7/i0_4 , \SB1_1_7/i0[10] , \SB1_1_7/i0[9] , \SB1_1_7/i0[8] ,
         \SB1_1_7/i0[7] , \SB1_1_7/i0[6] , \SB1_1_8/buf_output[5] ,
         \SB1_1_8/buf_output[4] , \SB1_1_8/buf_output[3] ,
         \SB1_1_8/buf_output[2] , \SB1_1_8/buf_output[1] ,
         \SB1_1_8/buf_output[0] , \SB1_1_8/i3[0] , \SB1_1_8/i1_5 ,
         \SB1_1_8/i1_7 , \SB1_1_8/i1[9] , \SB1_1_8/i0_0 , \SB1_1_8/i0_3 ,
         \SB1_1_8/i0_4 , \SB1_1_8/i0[10] , \SB1_1_8/i0[9] , \SB1_1_8/i0[8] ,
         \SB1_1_8/i0[7] , \SB1_1_8/i0[6] , \SB1_1_9/buf_output[5] ,
         \SB1_1_9/buf_output[4] , \SB1_1_9/buf_output[3] ,
         \SB1_1_9/buf_output[1] , \SB1_1_9/buf_output[0] , \SB1_1_9/i3[0] ,
         \SB1_1_9/i1_5 , \SB1_1_9/i1_7 , \SB1_1_9/i1[9] , \SB1_1_9/i0_0 ,
         \SB1_1_9/i0_3 , \SB1_1_9/i0_4 , \SB1_1_9/i0[10] , \SB1_1_9/i0[9] ,
         \SB1_1_9/i0[8] , \SB1_1_9/i0[7] , \SB1_1_9/i0[6] ,
         \SB1_1_10/buf_output[5] , \SB1_1_10/buf_output[4] ,
         \SB1_1_10/buf_output[3] , \SB1_1_10/buf_output[2] ,
         \SB1_1_10/buf_output[1] , \SB1_1_10/buf_output[0] , \SB1_1_10/i3[0] ,
         \SB1_1_10/i1_5 , \SB1_1_10/i1_7 , \SB1_1_10/i1[9] , \SB1_1_10/i0_0 ,
         \SB1_1_10/i0_3 , \SB1_1_10/i0_4 , \SB1_1_10/i0[10] , \SB1_1_10/i0[9] ,
         \SB1_1_10/i0[8] , \SB1_1_10/i0[7] , \SB1_1_10/i0[6] ,
         \SB1_1_11/buf_output[5] , \SB1_1_11/buf_output[4] ,
         \SB1_1_11/buf_output[3] , \SB1_1_11/buf_output[2] ,
         \SB1_1_11/buf_output[1] , \SB1_1_11/buf_output[0] , \SB1_1_11/i3[0] ,
         \SB1_1_11/i1_5 , \SB1_1_11/i1_7 , \SB1_1_11/i1[9] , \SB1_1_11/i0_0 ,
         \SB1_1_11/i0_3 , \SB1_1_11/i0_4 , \SB1_1_11/i0[10] , \SB1_1_11/i0[9] ,
         \SB1_1_11/i0[8] , \SB1_1_11/i0[7] , \SB1_1_11/i0[6] ,
         \SB1_1_12/buf_output[5] , \SB1_1_12/buf_output[4] ,
         \SB1_1_12/buf_output[3] , \SB1_1_12/buf_output[2] ,
         \SB1_1_12/buf_output[1] , \SB1_1_12/buf_output[0] , \SB1_1_12/i3[0] ,
         \SB1_1_12/i1_5 , \SB1_1_12/i1_7 , \SB1_1_12/i1[9] , \SB1_1_12/i0_0 ,
         \SB1_1_12/i0_3 , \SB1_1_12/i0_4 , \SB1_1_12/i0[10] , \SB1_1_12/i0[9] ,
         \SB1_1_12/i0[8] , \SB1_1_12/i0[7] , \SB1_1_12/i0[6] ,
         \SB1_1_13/buf_output[5] , \SB1_1_13/buf_output[4] ,
         \SB1_1_13/buf_output[3] , \SB1_1_13/buf_output[2] ,
         \SB1_1_13/buf_output[1] , \SB1_1_13/buf_output[0] , \SB1_1_13/i3[0] ,
         \SB1_1_13/i1_5 , \SB1_1_13/i1_7 , \SB1_1_13/i1[9] , \SB1_1_13/i0_0 ,
         \SB1_1_13/i0_3 , \SB1_1_13/i0_4 , \SB1_1_13/i0[10] , \SB1_1_13/i0[9] ,
         \SB1_1_13/i0[8] , \SB1_1_13/i0[7] , \SB1_1_13/i0[6] ,
         \SB1_1_14/buf_output[5] , \SB1_1_14/buf_output[4] ,
         \SB1_1_14/buf_output[3] , \SB1_1_14/buf_output[2] ,
         \SB1_1_14/buf_output[1] , \SB1_1_14/buf_output[0] , \SB1_1_14/i3[0] ,
         \SB1_1_14/i1_5 , \SB1_1_14/i1_7 , \SB1_1_14/i1[9] , \SB1_1_14/i0_0 ,
         \SB1_1_14/i0_3 , \SB1_1_14/i0_4 , \SB1_1_14/i0[10] , \SB1_1_14/i0[9] ,
         \SB1_1_14/i0[8] , \SB1_1_14/i0[7] , \SB1_1_14/i0[6] ,
         \SB1_1_15/buf_output[5] , \SB1_1_15/buf_output[4] ,
         \SB1_1_15/buf_output[2] , \SB1_1_15/buf_output[1] ,
         \SB1_1_15/buf_output[0] , \SB1_1_15/i3[0] , \SB1_1_15/i1_5 ,
         \SB1_1_15/i1_7 , \SB1_1_15/i1[9] , \SB1_1_15/i0_0 , \SB1_1_15/i0_3 ,
         \SB1_1_15/i0_4 , \SB1_1_15/i0[10] , \SB1_1_15/i0[9] ,
         \SB1_1_15/i0[8] , \SB1_1_15/i0[7] , \SB1_1_15/i0[6] ,
         \SB1_1_16/buf_output[5] , \SB1_1_16/buf_output[4] ,
         \SB1_1_16/buf_output[3] , \SB1_1_16/buf_output[2] ,
         \SB1_1_16/buf_output[1] , \SB1_1_16/buf_output[0] , \SB1_1_16/i3[0] ,
         \SB1_1_16/i1_5 , \SB1_1_16/i1_7 , \SB1_1_16/i1[9] , \SB1_1_16/i0_0 ,
         \SB1_1_16/i0_3 , \SB1_1_16/i0_4 , \SB1_1_16/i0[10] , \SB1_1_16/i0[9] ,
         \SB1_1_16/i0[8] , \SB1_1_16/i0[7] , \SB1_1_16/i0[6] ,
         \SB1_1_17/buf_output[5] , \SB1_1_17/buf_output[4] ,
         \SB1_1_17/buf_output[3] , \SB1_1_17/buf_output[2] ,
         \SB1_1_17/buf_output[1] , \SB1_1_17/buf_output[0] , \SB1_1_17/i3[0] ,
         \SB1_1_17/i1_5 , \SB1_1_17/i1_7 , \SB1_1_17/i1[9] , \SB1_1_17/i0_0 ,
         \SB1_1_17/i0_3 , \SB1_1_17/i0_4 , \SB1_1_17/i0[10] , \SB1_1_17/i0[9] ,
         \SB1_1_17/i0[8] , \SB1_1_17/i0[7] , \SB1_1_17/i0[6] ,
         \SB1_1_18/buf_output[5] , \SB1_1_18/buf_output[4] ,
         \SB1_1_18/buf_output[3] , \SB1_1_18/buf_output[2] ,
         \SB1_1_18/buf_output[1] , \SB1_1_18/buf_output[0] , \SB1_1_18/i3[0] ,
         \SB1_1_18/i1_5 , \SB1_1_18/i1_7 , \SB1_1_18/i1[9] , \SB1_1_18/i0_0 ,
         \SB1_1_18/i0_3 , \SB1_1_18/i0_4 , \SB1_1_18/i0[10] , \SB1_1_18/i0[9] ,
         \SB1_1_18/i0[8] , \SB1_1_18/i0[7] , \SB1_1_18/i0[6] ,
         \SB1_1_19/buf_output[5] , \SB1_1_19/buf_output[4] ,
         \SB1_1_19/buf_output[3] , \SB1_1_19/buf_output[2] ,
         \SB1_1_19/buf_output[1] , \SB1_1_19/buf_output[0] , \SB1_1_19/i3[0] ,
         \SB1_1_19/i1_5 , \SB1_1_19/i1_7 , \SB1_1_19/i1[9] , \SB1_1_19/i0_0 ,
         \SB1_1_19/i0_3 , \SB1_1_19/i0_4 , \SB1_1_19/i0[10] , \SB1_1_19/i0[9] ,
         \SB1_1_19/i0[8] , \SB1_1_19/i0[7] , \SB1_1_19/i0[6] ,
         \SB1_1_20/buf_output[5] , \SB1_1_20/buf_output[3] ,
         \SB1_1_20/buf_output[2] , \SB1_1_20/buf_output[1] ,
         \SB1_1_20/buf_output[0] , \SB1_1_20/i3[0] , \SB1_1_20/i1_5 ,
         \SB1_1_20/i1_7 , \SB1_1_20/i1[9] , \SB1_1_20/i0_0 , \SB1_1_20/i0_3 ,
         \SB1_1_20/i0_4 , \SB1_1_20/i0[10] , \SB1_1_20/i0[9] ,
         \SB1_1_20/i0[8] , \SB1_1_20/i0[7] , \SB1_1_20/i0[6] ,
         \SB1_1_21/buf_output[5] , \SB1_1_21/buf_output[3] ,
         \SB1_1_21/buf_output[2] , \SB1_1_21/buf_output[1] ,
         \SB1_1_21/buf_output[0] , \SB1_1_21/i3[0] , \SB1_1_21/i1_5 ,
         \SB1_1_21/i1_7 , \SB1_1_21/i1[9] , \SB1_1_21/i0_0 , \SB1_1_21/i0_3 ,
         \SB1_1_21/i0_4 , \SB1_1_21/i0[10] , \SB1_1_21/i0[9] ,
         \SB1_1_21/i0[8] , \SB1_1_21/i0[7] , \SB1_1_21/i0[6] ,
         \SB1_1_22/buf_output[5] , \SB1_1_22/buf_output[4] ,
         \SB1_1_22/buf_output[3] , \SB1_1_22/buf_output[2] ,
         \SB1_1_22/buf_output[1] , \SB1_1_22/buf_output[0] , \SB1_1_22/i3[0] ,
         \SB1_1_22/i1_5 , \SB1_1_22/i1_7 , \SB1_1_22/i1[9] , \SB1_1_22/i0_0 ,
         \SB1_1_22/i0_3 , \SB1_1_22/i0_4 , \SB1_1_22/i0[10] , \SB1_1_22/i0[9] ,
         \SB1_1_22/i0[8] , \SB1_1_22/i0[7] , \SB1_1_22/i0[6] ,
         \SB1_1_23/buf_output[5] , \SB1_1_23/buf_output[3] ,
         \SB1_1_23/buf_output[2] , \SB1_1_23/buf_output[1] ,
         \SB1_1_23/buf_output[0] , \SB1_1_23/i3[0] , \SB1_1_23/i1_5 ,
         \SB1_1_23/i1_7 , \SB1_1_23/i1[9] , \SB1_1_23/i0_0 , \SB1_1_23/i0_3 ,
         \SB1_1_23/i0_4 , \SB1_1_23/i0[10] , \SB1_1_23/i0[9] ,
         \SB1_1_23/i0[8] , \SB1_1_23/i0[7] , \SB1_1_23/i0[6] ,
         \SB1_1_24/buf_output[5] , \SB1_1_24/buf_output[4] ,
         \SB1_1_24/buf_output[3] , \SB1_1_24/buf_output[2] ,
         \SB1_1_24/buf_output[1] , \SB1_1_24/buf_output[0] , \SB1_1_24/i3[0] ,
         \SB1_1_24/i1_5 , \SB1_1_24/i1_7 , \SB1_1_24/i1[9] , \SB1_1_24/i0_0 ,
         \SB1_1_24/i0_4 , \SB1_1_24/i0[10] , \SB1_1_24/i0[9] ,
         \SB1_1_24/i0[8] , \SB1_1_24/i0[7] , \SB1_1_24/i0[6] ,
         \SB1_1_25/buf_output[5] , \SB1_1_25/buf_output[4] ,
         \SB1_1_25/buf_output[3] , \SB1_1_25/buf_output[2] ,
         \SB1_1_25/buf_output[1] , \SB1_1_25/buf_output[0] , \SB1_1_25/i3[0] ,
         \SB1_1_25/i1_5 , \SB1_1_25/i1_7 , \SB1_1_25/i1[9] , \SB1_1_25/i0_0 ,
         \SB1_1_25/i0_3 , \SB1_1_25/i0_4 , \SB1_1_25/i0[10] , \SB1_1_25/i0[9] ,
         \SB1_1_25/i0[8] , \SB1_1_25/i0[7] , \SB1_1_25/i0[6] ,
         \SB1_1_26/buf_output[5] , \SB1_1_26/buf_output[4] ,
         \SB1_1_26/buf_output[3] , \SB1_1_26/buf_output[2] ,
         \SB1_1_26/buf_output[1] , \SB1_1_26/buf_output[0] , \SB1_1_26/i3[0] ,
         \SB1_1_26/i1_5 , \SB1_1_26/i1_7 , \SB1_1_26/i1[9] , \SB1_1_26/i0_0 ,
         \SB1_1_26/i0_3 , \SB1_1_26/i0_4 , \SB1_1_26/i0[10] , \SB1_1_26/i0[9] ,
         \SB1_1_26/i0[8] , \SB1_1_26/i0[7] , \SB1_1_26/i0[6] ,
         \SB1_1_27/buf_output[5] , \SB1_1_27/buf_output[4] ,
         \SB1_1_27/buf_output[3] , \SB1_1_27/buf_output[2] ,
         \SB1_1_27/buf_output[1] , \SB1_1_27/buf_output[0] , \SB1_1_27/i3[0] ,
         \SB1_1_27/i1_5 , \SB1_1_27/i1_7 , \SB1_1_27/i1[9] , \SB1_1_27/i0_0 ,
         \SB1_1_27/i0_3 , \SB1_1_27/i0_4 , \SB1_1_27/i0[10] , \SB1_1_27/i0[9] ,
         \SB1_1_27/i0[8] , \SB1_1_27/i0[7] , \SB1_1_27/i0[6] ,
         \SB1_1_28/buf_output[5] , \SB1_1_28/buf_output[4] ,
         \SB1_1_28/buf_output[3] , \SB1_1_28/buf_output[2] ,
         \SB1_1_28/buf_output[1] , \SB1_1_28/buf_output[0] , \SB1_1_28/i3[0] ,
         \SB1_1_28/i1_5 , \SB1_1_28/i1_7 , \SB1_1_28/i1[9] , \SB1_1_28/i0_0 ,
         \SB1_1_28/i0_3 , \SB1_1_28/i0_4 , \SB1_1_28/i0[10] , \SB1_1_28/i0[9] ,
         \SB1_1_28/i0[8] , \SB1_1_28/i0[7] , \SB1_1_28/i0[6] ,
         \SB1_1_29/buf_output[5] , \SB1_1_29/buf_output[4] ,
         \SB1_1_29/buf_output[3] , \SB1_1_29/buf_output[2] ,
         \SB1_1_29/buf_output[1] , \SB1_1_29/buf_output[0] , \SB1_1_29/i3[0] ,
         \SB1_1_29/i1_5 , \SB1_1_29/i1_7 , \SB1_1_29/i1[9] , \SB1_1_29/i0_0 ,
         \SB1_1_29/i0_3 , \SB1_1_29/i0_4 , \SB1_1_29/i0[10] , \SB1_1_29/i0[9] ,
         \SB1_1_29/i0[8] , \SB1_1_29/i0[7] , \SB1_1_29/i0[6] ,
         \SB1_1_30/buf_output[5] , \SB1_1_30/buf_output[3] ,
         \SB1_1_30/buf_output[2] , \SB1_1_30/buf_output[1] ,
         \SB1_1_30/buf_output[0] , \SB1_1_30/i3[0] , \SB1_1_30/i1_5 ,
         \SB1_1_30/i1_7 , \SB1_1_30/i1[9] , \SB1_1_30/i0_0 , \SB1_1_30/i0_3 ,
         \SB1_1_30/i0_4 , \SB1_1_30/i0[10] , \SB1_1_30/i0[9] ,
         \SB1_1_30/i0[8] , \SB1_1_30/i0[7] , \SB1_1_30/i0[6] ,
         \SB1_1_31/buf_output[5] , \SB1_1_31/buf_output[4] ,
         \SB1_1_31/buf_output[3] , \SB1_1_31/buf_output[2] ,
         \SB1_1_31/buf_output[1] , \SB1_1_31/buf_output[0] , \SB1_1_31/i3[0] ,
         \SB1_1_31/i1_5 , \SB1_1_31/i1_7 , \SB1_1_31/i1[9] , \SB1_1_31/i0_0 ,
         \SB1_1_31/i0_3 , \SB1_1_31/i0_4 , \SB1_1_31/i0[10] , \SB1_1_31/i0[9] ,
         \SB1_1_31/i0[8] , \SB1_1_31/i0[7] , \SB1_1_31/i0[6] ,
         \SB2_1_0/buf_output[5] , \SB2_1_0/buf_output[4] ,
         \SB2_1_0/buf_output[3] , \SB2_1_0/buf_output[2] ,
         \SB2_1_0/buf_output[1] , \SB2_1_0/buf_output[0] , \SB2_1_0/i3[0] ,
         \SB2_1_0/i1_5 , \SB2_1_0/i1_7 , \SB2_1_0/i1[9] , \SB2_1_0/i0_0 ,
         \SB2_1_0/i0_3 , \SB2_1_0/i0[10] , \SB2_1_0/i0[9] , \SB2_1_0/i0[8] ,
         \SB2_1_0/i0[7] , \SB2_1_0/i0[6] , \SB2_1_1/buf_output[5] ,
         \SB2_1_1/buf_output[4] , \SB2_1_1/buf_output[3] ,
         \SB2_1_1/buf_output[0] , \SB2_1_1/i3[0] , \SB2_1_1/i1_5 ,
         \SB2_1_1/i1_7 , \SB2_1_1/i1[9] , \SB2_1_1/i0_0 , \SB2_1_1/i0_3 ,
         \SB2_1_1/i0_4 , \SB2_1_1/i0[10] , \SB2_1_1/i0[9] , \SB2_1_1/i0[8] ,
         \SB2_1_1/i0[7] , \SB2_1_1/i0[6] , \SB2_1_2/buf_output[5] ,
         \SB2_1_2/buf_output[4] , \SB2_1_2/buf_output[3] ,
         \SB2_1_2/buf_output[2] , \SB2_1_2/buf_output[1] ,
         \SB2_1_2/buf_output[0] , \SB2_1_2/i3[0] , \SB2_1_2/i1_5 ,
         \SB2_1_2/i1_7 , \SB2_1_2/i1[9] , \SB2_1_2/i0_0 , \SB2_1_2/i0_3 ,
         \SB2_1_2/i0_4 , \SB2_1_2/i0[10] , \SB2_1_2/i0[9] , \SB2_1_2/i0[8] ,
         \SB2_1_2/i0[7] , \SB2_1_2/i0[6] , \SB2_1_3/buf_output[5] ,
         \SB2_1_3/buf_output[4] , \SB2_1_3/buf_output[3] ,
         \SB2_1_3/buf_output[2] , \SB2_1_3/buf_output[1] ,
         \SB2_1_3/buf_output[0] , \SB2_1_3/i3[0] , \SB2_1_3/i1_5 ,
         \SB2_1_3/i1_7 , \SB2_1_3/i1[9] , \SB2_1_3/i0_0 , \SB2_1_3/i0_3 ,
         \SB2_1_3/i0_4 , \SB2_1_3/i0[10] , \SB2_1_3/i0[9] , \SB2_1_3/i0[8] ,
         \SB2_1_3/i0[7] , \SB2_1_3/i0[6] , \SB2_1_4/buf_output[5] ,
         \SB2_1_4/buf_output[3] , \SB2_1_4/buf_output[2] ,
         \SB2_1_4/buf_output[1] , \SB2_1_4/buf_output[0] , \SB2_1_4/i3[0] ,
         \SB2_1_4/i1_5 , \SB2_1_4/i1_7 , \SB2_1_4/i1[9] , \SB2_1_4/i0_0 ,
         \SB2_1_4/i0_3 , \SB2_1_4/i0_4 , \SB2_1_4/i0[10] , \SB2_1_4/i0[9] ,
         \SB2_1_4/i0[8] , \SB2_1_4/i0[7] , \SB2_1_5/buf_output[5] ,
         \SB2_1_5/buf_output[4] , \SB2_1_5/buf_output[3] ,
         \SB2_1_5/buf_output[2] , \SB2_1_5/buf_output[1] ,
         \SB2_1_5/buf_output[0] , \SB2_1_5/i3[0] , \SB2_1_5/i1_5 ,
         \SB2_1_5/i1_7 , \SB2_1_5/i1[9] , \SB2_1_5/i0_0 , \SB2_1_5/i0_3 ,
         \SB2_1_5/i0_4 , \SB2_1_5/i0[10] , \SB2_1_5/i0[9] , \SB2_1_5/i0[8] ,
         \SB2_1_5/i0[7] , \SB2_1_5/i0[6] , \SB2_1_6/buf_output[5] ,
         \SB2_1_6/buf_output[4] , \SB2_1_6/buf_output[3] ,
         \SB2_1_6/buf_output[2] , \SB2_1_6/buf_output[1] ,
         \SB2_1_6/buf_output[0] , \SB2_1_6/i3[0] , \SB2_1_6/i1_5 ,
         \SB2_1_6/i1_7 , \SB2_1_6/i1[9] , \SB2_1_6/i0_0 , \SB2_1_6/i0_3 ,
         \SB2_1_6/i0_4 , \SB2_1_6/i0[10] , \SB2_1_6/i0[9] , \SB2_1_6/i0[8] ,
         \SB2_1_6/i0[7] , \SB2_1_6/i0[6] , \SB2_1_7/buf_output[5] ,
         \SB2_1_7/buf_output[4] , \SB2_1_7/buf_output[3] ,
         \SB2_1_7/buf_output[2] , \SB2_1_7/buf_output[1] ,
         \SB2_1_7/buf_output[0] , \SB2_1_7/i3[0] , \SB2_1_7/i1_5 ,
         \SB2_1_7/i1_7 , \SB2_1_7/i1[9] , \SB2_1_7/i0_0 , \SB2_1_7/i0_3 ,
         \SB2_1_7/i0_4 , \SB2_1_7/i0[10] , \SB2_1_7/i0[9] , \SB2_1_7/i0[8] ,
         \SB2_1_7/i0[7] , \SB2_1_7/i0[6] , \SB2_1_8/buf_output[5] ,
         \SB2_1_8/buf_output[4] , \SB2_1_8/buf_output[3] ,
         \SB2_1_8/buf_output[2] , \SB2_1_8/buf_output[1] ,
         \SB2_1_8/buf_output[0] , \SB2_1_8/i3[0] , \SB2_1_8/i1_5 ,
         \SB2_1_8/i1_7 , \SB2_1_8/i1[9] , \SB2_1_8/i0_0 , \SB2_1_8/i0_3 ,
         \SB2_1_8/i0_4 , \SB2_1_8/i0[10] , \SB2_1_8/i0[9] , \SB2_1_8/i0[8] ,
         \SB2_1_8/i0[7] , \SB2_1_8/i0[6] , \SB2_1_9/buf_output[5] ,
         \SB2_1_9/buf_output[4] , \SB2_1_9/buf_output[3] ,
         \SB2_1_9/buf_output[2] , \SB2_1_9/buf_output[1] ,
         \SB2_1_9/buf_output[0] , \SB2_1_9/i3[0] , \SB2_1_9/i1_5 ,
         \SB2_1_9/i1_7 , \SB2_1_9/i1[9] , \SB2_1_9/i0_0 , \SB2_1_9/i0_3 ,
         \SB2_1_9/i0_4 , \SB2_1_9/i0[10] , \SB2_1_9/i0[9] , \SB2_1_9/i0[8] ,
         \SB2_1_9/i0[7] , \SB2_1_9/i0[6] , \SB2_1_10/buf_output[5] ,
         \SB2_1_10/buf_output[4] , \SB2_1_10/buf_output[3] ,
         \SB2_1_10/buf_output[2] , \SB2_1_10/buf_output[1] ,
         \SB2_1_10/buf_output[0] , \SB2_1_10/i3[0] , \SB2_1_10/i1_5 ,
         \SB2_1_10/i1_7 , \SB2_1_10/i1[9] , \SB2_1_10/i0_0 , \SB2_1_10/i0_3 ,
         \SB2_1_10/i0_4 , \SB2_1_10/i0[10] , \SB2_1_10/i0[9] ,
         \SB2_1_10/i0[8] , \SB2_1_10/i0[7] , \SB2_1_10/i0[6] ,
         \SB2_1_11/buf_output[5] , \SB2_1_11/buf_output[4] ,
         \SB2_1_11/buf_output[3] , \SB2_1_11/buf_output[2] ,
         \SB2_1_11/buf_output[1] , \SB2_1_11/buf_output[0] , \SB2_1_11/i3[0] ,
         \SB2_1_11/i1_5 , \SB2_1_11/i1_7 , \SB2_1_11/i1[9] , \SB2_1_11/i0_0 ,
         \SB2_1_11/i0_3 , \SB2_1_11/i0_4 , \SB2_1_11/i0[10] , \SB2_1_11/i0[9] ,
         \SB2_1_11/i0[8] , \SB2_1_11/i0[7] , \SB2_1_11/i0[6] ,
         \SB2_1_12/buf_output[5] , \SB2_1_12/buf_output[4] ,
         \SB2_1_12/buf_output[3] , \SB2_1_12/buf_output[2] ,
         \SB2_1_12/buf_output[1] , \SB2_1_12/buf_output[0] , \SB2_1_12/i3[0] ,
         \SB2_1_12/i1_5 , \SB2_1_12/i1_7 , \SB2_1_12/i1[9] , \SB2_1_12/i0_0 ,
         \SB2_1_12/i0_3 , \SB2_1_12/i0_4 , \SB2_1_12/i0[10] , \SB2_1_12/i0[9] ,
         \SB2_1_12/i0[8] , \SB2_1_12/i0[7] , \SB2_1_12/i0[6] ,
         \SB2_1_13/buf_output[5] , \SB2_1_13/buf_output[4] ,
         \SB2_1_13/buf_output[3] , \SB2_1_13/buf_output[2] ,
         \SB2_1_13/buf_output[1] , \SB2_1_13/buf_output[0] , \SB2_1_13/i3[0] ,
         \SB2_1_13/i1_5 , \SB2_1_13/i1_7 , \SB2_1_13/i1[9] , \SB2_1_13/i0_0 ,
         \SB2_1_13/i0_3 , \SB2_1_13/i0_4 , \SB2_1_13/i0[10] , \SB2_1_13/i0[9] ,
         \SB2_1_13/i0[8] , \SB2_1_13/i0[7] , \SB2_1_13/i0[6] ,
         \SB2_1_14/buf_output[5] , \SB2_1_14/buf_output[4] ,
         \SB2_1_14/buf_output[3] , \SB2_1_14/buf_output[2] ,
         \SB2_1_14/buf_output[1] , \SB2_1_14/buf_output[0] , \SB2_1_14/i3[0] ,
         \SB2_1_14/i1_5 , \SB2_1_14/i1_7 , \SB2_1_14/i1[9] , \SB2_1_14/i0_0 ,
         \SB2_1_14/i0_3 , \SB2_1_14/i0_4 , \SB2_1_14/i0[10] , \SB2_1_14/i0[9] ,
         \SB2_1_14/i0[8] , \SB2_1_14/i0[7] , \SB2_1_14/i0[6] ,
         \SB2_1_15/buf_output[5] , \SB2_1_15/buf_output[4] ,
         \SB2_1_15/buf_output[3] , \SB2_1_15/buf_output[2] ,
         \SB2_1_15/buf_output[1] , \SB2_1_15/buf_output[0] , \SB2_1_15/i3[0] ,
         \SB2_1_15/i1_5 , \SB2_1_15/i1_7 , \SB2_1_15/i1[9] , \SB2_1_15/i0_0 ,
         \SB2_1_15/i0_3 , \SB2_1_15/i0_4 , \SB2_1_15/i0[10] , \SB2_1_15/i0[9] ,
         \SB2_1_15/i0[8] , \SB2_1_15/i0[7] , \SB2_1_15/i0[6] ,
         \SB2_1_16/buf_output[5] , \SB2_1_16/buf_output[4] ,
         \SB2_1_16/buf_output[3] , \SB2_1_16/buf_output[2] ,
         \SB2_1_16/buf_output[1] , \SB2_1_16/buf_output[0] , \SB2_1_16/i3[0] ,
         \SB2_1_16/i1_5 , \SB2_1_16/i1_7 , \SB2_1_16/i1[9] , \SB2_1_16/i0_0 ,
         \SB2_1_16/i0_3 , \SB2_1_16/i0_4 , \SB2_1_16/i0[10] , \SB2_1_16/i0[9] ,
         \SB2_1_16/i0[8] , \SB2_1_16/i0[7] , \SB2_1_16/i0[6] ,
         \SB2_1_17/buf_output[5] , \SB2_1_17/buf_output[4] ,
         \SB2_1_17/buf_output[3] , \SB2_1_17/buf_output[2] ,
         \SB2_1_17/buf_output[1] , \SB2_1_17/buf_output[0] , \SB2_1_17/i3[0] ,
         \SB2_1_17/i1_7 , \SB2_1_17/i1[9] , \SB2_1_17/i0_0 , \SB2_1_17/i0_3 ,
         \SB2_1_17/i0_4 , \SB2_1_17/i0[10] , \SB2_1_17/i0[9] ,
         \SB2_1_17/i0[8] , \SB2_1_17/i0[7] , \SB2_1_17/i0[6] ,
         \SB2_1_18/buf_output[5] , \SB2_1_18/buf_output[4] ,
         \SB2_1_18/buf_output[3] , \SB2_1_18/buf_output[2] ,
         \SB2_1_18/buf_output[1] , \SB2_1_18/buf_output[0] , \SB2_1_18/i3[0] ,
         \SB2_1_18/i1_5 , \SB2_1_18/i1_7 , \SB2_1_18/i1[9] , \SB2_1_18/i0_0 ,
         \SB2_1_18/i0_3 , \SB2_1_18/i0_4 , \SB2_1_18/i0[10] , \SB2_1_18/i0[9] ,
         \SB2_1_18/i0[8] , \SB2_1_18/i0[7] , \SB2_1_18/i0[6] ,
         \SB2_1_19/buf_output[5] , \SB2_1_19/buf_output[4] ,
         \SB2_1_19/buf_output[3] , \SB2_1_19/buf_output[2] ,
         \SB2_1_19/buf_output[1] , \SB2_1_19/buf_output[0] , \SB2_1_19/i3[0] ,
         \SB2_1_19/i1_5 , \SB2_1_19/i1_7 , \SB2_1_19/i1[9] , \SB2_1_19/i0_0 ,
         \SB2_1_19/i0_3 , \SB2_1_19/i0_4 , \SB2_1_19/i0[10] , \SB2_1_19/i0[9] ,
         \SB2_1_19/i0[8] , \SB2_1_19/i0[7] , \SB2_1_19/i0[6] ,
         \SB2_1_20/buf_output[5] , \SB2_1_20/buf_output[4] ,
         \SB2_1_20/buf_output[3] , \SB2_1_20/buf_output[2] ,
         \SB2_1_20/buf_output[1] , \SB2_1_20/buf_output[0] , \SB2_1_20/i3[0] ,
         \SB2_1_20/i1_5 , \SB2_1_20/i1_7 , \SB2_1_20/i1[9] , \SB2_1_20/i0_0 ,
         \SB2_1_20/i0_3 , \SB2_1_20/i0_4 , \SB2_1_20/i0[10] , \SB2_1_20/i0[9] ,
         \SB2_1_20/i0[8] , \SB2_1_20/i0[7] , \SB2_1_20/i0[6] ,
         \SB2_1_21/buf_output[5] , \SB2_1_21/buf_output[4] ,
         \SB2_1_21/buf_output[3] , \SB2_1_21/buf_output[2] ,
         \SB2_1_21/buf_output[1] , \SB2_1_21/buf_output[0] , \SB2_1_21/i3[0] ,
         \SB2_1_21/i1_5 , \SB2_1_21/i1_7 , \SB2_1_21/i1[9] , \SB2_1_21/i0_0 ,
         \SB2_1_21/i0_3 , \SB2_1_21/i0_4 , \SB2_1_21/i0[10] , \SB2_1_21/i0[9] ,
         \SB2_1_21/i0[8] , \SB2_1_21/i0[7] , \SB2_1_21/i0[6] ,
         \SB2_1_22/buf_output[5] , \SB2_1_22/buf_output[4] ,
         \SB2_1_22/buf_output[3] , \SB2_1_22/buf_output[2] ,
         \SB2_1_22/buf_output[1] , \SB2_1_22/buf_output[0] , \SB2_1_22/i3[0] ,
         \SB2_1_22/i1_5 , \SB2_1_22/i1_7 , \SB2_1_22/i1[9] , \SB2_1_22/i0_0 ,
         \SB2_1_22/i0_3 , \SB2_1_22/i0_4 , \SB2_1_22/i0[10] , \SB2_1_22/i0[9] ,
         \SB2_1_22/i0[7] , \SB2_1_22/i0[6] , \SB2_1_23/buf_output[5] ,
         \SB2_1_23/buf_output[4] , \SB2_1_23/buf_output[3] ,
         \SB2_1_23/buf_output[2] , \SB2_1_23/buf_output[1] ,
         \SB2_1_23/buf_output[0] , \SB2_1_23/i3[0] , \SB2_1_23/i1_5 ,
         \SB2_1_23/i1_7 , \SB2_1_23/i1[9] , \SB2_1_23/i0_0 , \SB2_1_23/i0_3 ,
         \SB2_1_23/i0_4 , \SB2_1_23/i0[10] , \SB2_1_23/i0[9] ,
         \SB2_1_23/i0[8] , \SB2_1_23/i0[7] , \SB2_1_23/i0[6] ,
         \SB2_1_24/buf_output[5] , \SB2_1_24/buf_output[4] ,
         \SB2_1_24/buf_output[3] , \SB2_1_24/buf_output[2] ,
         \SB2_1_24/buf_output[1] , \SB2_1_24/buf_output[0] , \SB2_1_24/i3[0] ,
         \SB2_1_24/i1_5 , \SB2_1_24/i1_7 , \SB2_1_24/i1[9] , \SB2_1_24/i0_0 ,
         \SB2_1_24/i0_3 , \SB2_1_24/i0_4 , \SB2_1_24/i0[10] , \SB2_1_24/i0[9] ,
         \SB2_1_24/i0[8] , \SB2_1_24/i0[7] , \SB2_1_24/i0[6] ,
         \SB2_1_25/buf_output[5] , \SB2_1_25/buf_output[4] ,
         \SB2_1_25/buf_output[3] , \SB2_1_25/buf_output[2] ,
         \SB2_1_25/buf_output[1] , \SB2_1_25/buf_output[0] , \SB2_1_25/i3[0] ,
         \SB2_1_25/i1_5 , \SB2_1_25/i1_7 , \SB2_1_25/i1[9] , \SB2_1_25/i0_0 ,
         \SB2_1_25/i0_3 , \SB2_1_25/i0_4 , \SB2_1_25/i0[9] , \SB2_1_25/i0[7] ,
         \SB2_1_25/i0[6] , \SB2_1_26/buf_output[5] , \SB2_1_26/buf_output[4] ,
         \SB2_1_26/buf_output[3] , \SB2_1_26/buf_output[2] ,
         \SB2_1_26/buf_output[1] , \SB2_1_26/buf_output[0] , \SB2_1_26/i3[0] ,
         \SB2_1_26/i1_5 , \SB2_1_26/i1_7 , \SB2_1_26/i1[9] , \SB2_1_26/i0_0 ,
         \SB2_1_26/i0_3 , \SB2_1_26/i0_4 , \SB2_1_26/i0[10] , \SB2_1_26/i0[9] ,
         \SB2_1_26/i0[8] , \SB2_1_26/i0[7] , \SB2_1_26/i0[6] ,
         \SB2_1_27/buf_output[5] , \SB2_1_27/buf_output[4] ,
         \SB2_1_27/buf_output[3] , \SB2_1_27/buf_output[2] ,
         \SB2_1_27/buf_output[1] , \SB2_1_27/buf_output[0] , \SB2_1_27/i3[0] ,
         \SB2_1_27/i1_5 , \SB2_1_27/i1_7 , \SB2_1_27/i1[9] , \SB2_1_27/i0_3 ,
         \SB2_1_27/i0_4 , \SB2_1_27/i0[10] , \SB2_1_27/i0[9] ,
         \SB2_1_27/i0[8] , \SB2_1_27/i0[7] , \SB2_1_27/i0[6] ,
         \SB2_1_28/buf_output[5] , \SB2_1_28/buf_output[4] ,
         \SB2_1_28/buf_output[3] , \SB2_1_28/buf_output[2] ,
         \SB2_1_28/buf_output[1] , \SB2_1_28/buf_output[0] , \SB2_1_28/i3[0] ,
         \SB2_1_28/i1_5 , \SB2_1_28/i1_7 , \SB2_1_28/i1[9] , \SB2_1_28/i0_0 ,
         \SB2_1_28/i0_3 , \SB2_1_28/i0_4 , \SB2_1_28/i0[10] , \SB2_1_28/i0[9] ,
         \SB2_1_28/i0[8] , \SB2_1_28/i0[7] , \SB2_1_28/i0[6] ,
         \SB2_1_29/buf_output[5] , \SB2_1_29/buf_output[4] ,
         \SB2_1_29/buf_output[3] , \SB2_1_29/buf_output[2] ,
         \SB2_1_29/buf_output[1] , \SB2_1_29/buf_output[0] , \SB2_1_29/i3[0] ,
         \SB2_1_29/i1_5 , \SB2_1_29/i1_7 , \SB2_1_29/i1[9] , \SB2_1_29/i0_0 ,
         \SB2_1_29/i0_3 , \SB2_1_29/i0_4 , \SB2_1_29/i0[10] , \SB2_1_29/i0[9] ,
         \SB2_1_29/i0[8] , \SB2_1_29/i0[6] , \SB2_1_30/buf_output[5] ,
         \SB2_1_30/buf_output[4] , \SB2_1_30/buf_output[3] ,
         \SB2_1_30/buf_output[2] , \SB2_1_30/buf_output[1] ,
         \SB2_1_30/buf_output[0] , \SB2_1_30/i3[0] , \SB2_1_30/i1_5 ,
         \SB2_1_30/i1_7 , \SB2_1_30/i1[9] , \SB2_1_30/i0_0 , \SB2_1_30/i0_3 ,
         \SB2_1_30/i0_4 , \SB2_1_30/i0[10] , \SB2_1_30/i0[9] ,
         \SB2_1_30/i0[8] , \SB2_1_30/i0[7] , \SB2_1_30/i0[6] ,
         \SB2_1_31/buf_output[5] , \SB2_1_31/buf_output[4] ,
         \SB2_1_31/buf_output[3] , \SB2_1_31/buf_output[2] ,
         \SB2_1_31/buf_output[1] , \SB2_1_31/buf_output[0] , \SB2_1_31/i3[0] ,
         \SB2_1_31/i1_5 , \SB2_1_31/i1_7 , \SB2_1_31/i1[9] , \SB2_1_31/i0_0 ,
         \SB2_1_31/i0_3 , \SB2_1_31/i0_4 , \SB2_1_31/i0[10] , \SB2_1_31/i0[9] ,
         \SB2_1_31/i0[8] , \SB2_1_31/i0[7] , \SB2_1_31/i0[6] ,
         \SB1_2_0/buf_output[5] , \SB1_2_0/buf_output[4] ,
         \SB1_2_0/buf_output[3] , \SB1_2_0/buf_output[2] ,
         \SB1_2_0/buf_output[1] , \SB1_2_0/buf_output[0] , \SB1_2_0/i3[0] ,
         \SB1_2_0/i1_5 , \SB1_2_0/i1_7 , \SB1_2_0/i1[9] , \SB1_2_0/i0_0 ,
         \SB1_2_0/i0_4 , \SB1_2_0/i0[10] , \SB1_2_0/i0[9] , \SB1_2_0/i0[8] ,
         \SB1_2_0/i0[7] , \SB1_2_0/i0[6] , \SB1_2_1/buf_output[5] ,
         \SB1_2_1/buf_output[3] , \SB1_2_1/buf_output[2] ,
         \SB1_2_1/buf_output[1] , \SB1_2_1/buf_output[0] , \SB1_2_1/i3[0] ,
         \SB1_2_1/i1_5 , \SB1_2_1/i1_7 , \SB1_2_1/i1[9] , \SB1_2_1/i0_0 ,
         \SB1_2_1/i0_3 , \SB1_2_1/i0_4 , \SB1_2_1/i0[10] , \SB1_2_1/i0[9] ,
         \SB1_2_1/i0[8] , \SB1_2_1/i0[7] , \SB1_2_1/i0[6] ,
         \SB1_2_2/buf_output[5] , \SB1_2_2/buf_output[4] ,
         \SB1_2_2/buf_output[3] , \SB1_2_2/buf_output[2] ,
         \SB1_2_2/buf_output[1] , \SB1_2_2/buf_output[0] , \SB1_2_2/i3[0] ,
         \SB1_2_2/i1_5 , \SB1_2_2/i1_7 , \SB1_2_2/i1[9] , \SB1_2_2/i0_0 ,
         \SB1_2_2/i0_3 , \SB1_2_2/i0_4 , \SB1_2_2/i0[10] , \SB1_2_2/i0[9] ,
         \SB1_2_2/i0[8] , \SB1_2_2/i0[7] , \SB1_2_2/i0[6] ,
         \SB1_2_3/buf_output[5] , \SB1_2_3/buf_output[4] ,
         \SB1_2_3/buf_output[3] , \SB1_2_3/buf_output[2] ,
         \SB1_2_3/buf_output[1] , \SB1_2_3/buf_output[0] , \SB1_2_3/i3[0] ,
         \SB1_2_3/i1_5 , \SB1_2_3/i1_7 , \SB1_2_3/i1[9] , \SB1_2_3/i0_0 ,
         \SB1_2_3/i0_3 , \SB1_2_3/i0_4 , \SB1_2_3/i0[10] , \SB1_2_3/i0[9] ,
         \SB1_2_3/i0[8] , \SB1_2_3/i0[7] , \SB1_2_3/i0[6] ,
         \SB1_2_4/buf_output[5] , \SB1_2_4/buf_output[4] ,
         \SB1_2_4/buf_output[3] , \SB1_2_4/buf_output[2] ,
         \SB1_2_4/buf_output[1] , \SB1_2_4/buf_output[0] , \SB1_2_4/i3[0] ,
         \SB1_2_4/i1_5 , \SB1_2_4/i1_7 , \SB1_2_4/i1[9] , \SB1_2_4/i0_0 ,
         \SB1_2_4/i0_3 , \SB1_2_4/i0_4 , \SB1_2_4/i0[10] , \SB1_2_4/i0[9] ,
         \SB1_2_4/i0[8] , \SB1_2_4/i0[7] , \SB1_2_4/i0[6] ,
         \SB1_2_5/buf_output[5] , \SB1_2_5/buf_output[3] ,
         \SB1_2_5/buf_output[2] , \SB1_2_5/buf_output[1] ,
         \SB1_2_5/buf_output[0] , \SB1_2_5/i3[0] , \SB1_2_5/i1_5 ,
         \SB1_2_5/i1_7 , \SB1_2_5/i1[9] , \SB1_2_5/i0_0 , \SB1_2_5/i0_3 ,
         \SB1_2_5/i0_4 , \SB1_2_5/i0[10] , \SB1_2_5/i0[9] , \SB1_2_5/i0[8] ,
         \SB1_2_5/i0[7] , \SB1_2_5/i0[6] , \SB1_2_6/buf_output[5] ,
         \SB1_2_6/buf_output[4] , \SB1_2_6/buf_output[3] ,
         \SB1_2_6/buf_output[2] , \SB1_2_6/buf_output[1] ,
         \SB1_2_6/buf_output[0] , \SB1_2_6/i3[0] , \SB1_2_6/i1_5 ,
         \SB1_2_6/i1_7 , \SB1_2_6/i1[9] , \SB1_2_6/i0_0 , \SB1_2_6/i0_3 ,
         \SB1_2_6/i0_4 , \SB1_2_6/i0[10] , \SB1_2_6/i0[9] , \SB1_2_6/i0[8] ,
         \SB1_2_6/i0[7] , \SB1_2_6/i0[6] , \SB1_2_7/buf_output[5] ,
         \SB1_2_7/buf_output[4] , \SB1_2_7/buf_output[3] ,
         \SB1_2_7/buf_output[2] , \SB1_2_7/buf_output[1] ,
         \SB1_2_7/buf_output[0] , \SB1_2_7/i3[0] , \SB1_2_7/i1_5 ,
         \SB1_2_7/i1_7 , \SB1_2_7/i1[9] , \SB1_2_7/i0_0 , \SB1_2_7/i0_4 ,
         \SB1_2_7/i0[10] , \SB1_2_7/i0[9] , \SB1_2_7/i0[7] , \SB1_2_7/i0[6] ,
         \SB1_2_8/buf_output[5] , \SB1_2_8/buf_output[4] ,
         \SB1_2_8/buf_output[3] , \SB1_2_8/buf_output[2] ,
         \SB1_2_8/buf_output[1] , \SB1_2_8/buf_output[0] , \SB1_2_8/i3[0] ,
         \SB1_2_8/i1_5 , \SB1_2_8/i1_7 , \SB1_2_8/i1[9] , \SB1_2_8/i0_0 ,
         \SB1_2_8/i0_3 , \SB1_2_8/i0_4 , \SB1_2_8/i0[10] , \SB1_2_8/i0[9] ,
         \SB1_2_8/i0[8] , \SB1_2_8/i0[7] , \SB1_2_8/i0[6] ,
         \SB1_2_9/buf_output[5] , \SB1_2_9/buf_output[4] ,
         \SB1_2_9/buf_output[3] , \SB1_2_9/buf_output[2] ,
         \SB1_2_9/buf_output[1] , \SB1_2_9/buf_output[0] , \SB1_2_9/i3[0] ,
         \SB1_2_9/i1_5 , \SB1_2_9/i1_7 , \SB1_2_9/i1[9] , \SB1_2_9/i0_0 ,
         \SB1_2_9/i0_3 , \SB1_2_9/i0_4 , \SB1_2_9/i0[10] , \SB1_2_9/i0[9] ,
         \SB1_2_9/i0[8] , \SB1_2_9/i0[7] , \SB1_2_9/i0[6] ,
         \SB1_2_10/buf_output[4] , \SB1_2_10/buf_output[3] ,
         \SB1_2_10/buf_output[2] , \SB1_2_10/buf_output[1] ,
         \SB1_2_10/buf_output[0] , \SB1_2_10/i3[0] , \SB1_2_10/i1_5 ,
         \SB1_2_10/i1_7 , \SB1_2_10/i1[9] , \SB1_2_10/i0_0 , \SB1_2_10/i0_3 ,
         \SB1_2_10/i0_4 , \SB1_2_10/i0[10] , \SB1_2_10/i0[9] ,
         \SB1_2_10/i0[8] , \SB1_2_10/i0[7] , \SB1_2_10/i0[6] ,
         \SB1_2_11/buf_output[5] , \SB1_2_11/buf_output[4] ,
         \SB1_2_11/buf_output[3] , \SB1_2_11/buf_output[2] ,
         \SB1_2_11/buf_output[1] , \SB1_2_11/buf_output[0] , \SB1_2_11/i3[0] ,
         \SB1_2_11/i1_5 , \SB1_2_11/i1_7 , \SB1_2_11/i1[9] , \SB1_2_11/i0_0 ,
         \SB1_2_11/i0_3 , \SB1_2_11/i0_4 , \SB1_2_11/i0[10] , \SB1_2_11/i0[9] ,
         \SB1_2_11/i0[8] , \SB1_2_11/i0[7] , \SB1_2_11/i0[6] ,
         \SB1_2_12/buf_output[5] , \SB1_2_12/buf_output[4] ,
         \SB1_2_12/buf_output[3] , \SB1_2_12/buf_output[2] ,
         \SB1_2_12/buf_output[1] , \SB1_2_12/buf_output[0] , \SB1_2_12/i3[0] ,
         \SB1_2_12/i1_5 , \SB1_2_12/i1_7 , \SB1_2_12/i1[9] , \SB1_2_12/i0_4 ,
         \SB1_2_12/i0[10] , \SB1_2_12/i0[9] , \SB1_2_12/i0[8] ,
         \SB1_2_12/i0[7] , \SB1_2_12/i0[6] , \SB1_2_13/buf_output[5] ,
         \SB1_2_13/buf_output[4] , \SB1_2_13/buf_output[3] ,
         \SB1_2_13/buf_output[2] , \SB1_2_13/buf_output[1] ,
         \SB1_2_13/buf_output[0] , \SB1_2_13/i3[0] , \SB1_2_13/i1_5 ,
         \SB1_2_13/i1_7 , \SB1_2_13/i1[9] , \SB1_2_13/i0_0 , \SB1_2_13/i0_3 ,
         \SB1_2_13/i0_4 , \SB1_2_13/i0[10] , \SB1_2_13/i0[9] ,
         \SB1_2_13/i0[8] , \SB1_2_13/i0[7] , \SB1_2_13/i0[6] ,
         \SB1_2_14/buf_output[5] , \SB1_2_14/buf_output[4] ,
         \SB1_2_14/buf_output[3] , \SB1_2_14/buf_output[2] ,
         \SB1_2_14/buf_output[1] , \SB1_2_14/buf_output[0] , \SB1_2_14/i3[0] ,
         \SB1_2_14/i1_5 , \SB1_2_14/i1_7 , \SB1_2_14/i1[9] , \SB1_2_14/i0_0 ,
         \SB1_2_14/i0_4 , \SB1_2_14/i0[10] , \SB1_2_14/i0[9] ,
         \SB1_2_14/i0[8] , \SB1_2_14/i0[7] , \SB1_2_14/i0[6] ,
         \SB1_2_15/buf_output[5] , \SB1_2_15/buf_output[4] ,
         \SB1_2_15/buf_output[3] , \SB1_2_15/buf_output[2] ,
         \SB1_2_15/buf_output[0] , \SB1_2_15/i3[0] , \SB1_2_15/i1_5 ,
         \SB1_2_15/i1_7 , \SB1_2_15/i1[9] , \SB1_2_15/i0_0 , \SB1_2_15/i0_4 ,
         \SB1_2_15/i0[10] , \SB1_2_15/i0[9] , \SB1_2_15/i0[8] ,
         \SB1_2_15/i0[7] , \SB1_2_15/i0[6] , \SB1_2_16/buf_output[5] ,
         \SB1_2_16/buf_output[4] , \SB1_2_16/buf_output[3] ,
         \SB1_2_16/buf_output[2] , \SB1_2_16/buf_output[1] ,
         \SB1_2_16/buf_output[0] , \SB1_2_16/i3[0] , \SB1_2_16/i1_5 ,
         \SB1_2_16/i1_7 , \SB1_2_16/i1[9] , \SB1_2_16/i0_0 , \SB1_2_16/i0_3 ,
         \SB1_2_16/i0_4 , \SB1_2_16/i0[10] , \SB1_2_16/i0[9] ,
         \SB1_2_16/i0[8] , \SB1_2_16/i0[7] , \SB1_2_16/i0[6] ,
         \SB1_2_17/buf_output[5] , \SB1_2_17/buf_output[4] ,
         \SB1_2_17/buf_output[3] , \SB1_2_17/buf_output[2] ,
         \SB1_2_17/buf_output[1] , \SB1_2_17/buf_output[0] , \SB1_2_17/i3[0] ,
         \SB1_2_17/i1_5 , \SB1_2_17/i1_7 , \SB1_2_17/i1[9] , \SB1_2_17/i0_0 ,
         \SB1_2_17/i0_3 , \SB1_2_17/i0_4 , \SB1_2_17/i0[10] , \SB1_2_17/i0[9] ,
         \SB1_2_17/i0[8] , \SB1_2_17/i0[7] , \SB1_2_17/i0[6] ,
         \SB1_2_18/buf_output[5] , \SB1_2_18/buf_output[4] ,
         \SB1_2_18/buf_output[3] , \SB1_2_18/buf_output[2] ,
         \SB1_2_18/buf_output[1] , \SB1_2_18/buf_output[0] , \SB1_2_18/i3[0] ,
         \SB1_2_18/i1_5 , \SB1_2_18/i1_7 , \SB1_2_18/i1[9] , \SB1_2_18/i0_0 ,
         \SB1_2_18/i0_3 , \SB1_2_18/i0_4 , \SB1_2_18/i0[10] , \SB1_2_18/i0[9] ,
         \SB1_2_18/i0[8] , \SB1_2_18/i0[7] , \SB1_2_18/i0[6] ,
         \SB1_2_19/buf_output[5] , \SB1_2_19/buf_output[3] ,
         \SB1_2_19/buf_output[2] , \SB1_2_19/buf_output[0] , \SB1_2_19/i3[0] ,
         \SB1_2_19/i1_5 , \SB1_2_19/i1_7 , \SB1_2_19/i1[9] , \SB1_2_19/i0_0 ,
         \SB1_2_19/i0_3 , \SB1_2_19/i0_4 , \SB1_2_19/i0[10] , \SB1_2_19/i0[9] ,
         \SB1_2_19/i0[8] , \SB1_2_19/i0[7] , \SB1_2_19/i0[6] ,
         \SB1_2_20/buf_output[5] , \SB1_2_20/buf_output[4] ,
         \SB1_2_20/buf_output[3] , \SB1_2_20/buf_output[2] ,
         \SB1_2_20/buf_output[1] , \SB1_2_20/buf_output[0] , \SB1_2_20/i3[0] ,
         \SB1_2_20/i1_5 , \SB1_2_20/i1_7 , \SB1_2_20/i1[9] , \SB1_2_20/i0_0 ,
         \SB1_2_20/i0_3 , \SB1_2_20/i0_4 , \SB1_2_20/i0[10] , \SB1_2_20/i0[9] ,
         \SB1_2_20/i0[8] , \SB1_2_20/i0[7] , \SB1_2_20/i0[6] ,
         \SB1_2_21/buf_output[5] , \SB1_2_21/buf_output[4] ,
         \SB1_2_21/buf_output[3] , \SB1_2_21/buf_output[2] ,
         \SB1_2_21/buf_output[1] , \SB1_2_21/buf_output[0] , \SB1_2_21/i3[0] ,
         \SB1_2_21/i1_5 , \SB1_2_21/i1_7 , \SB1_2_21/i1[9] , \SB1_2_21/i0_0 ,
         \SB1_2_21/i0_3 , \SB1_2_21/i0_4 , \SB1_2_21/i0[10] , \SB1_2_21/i0[9] ,
         \SB1_2_21/i0[8] , \SB1_2_21/i0[7] , \SB1_2_21/i0[6] ,
         \SB1_2_22/buf_output[5] , \SB1_2_22/buf_output[4] ,
         \SB1_2_22/buf_output[3] , \SB1_2_22/buf_output[2] ,
         \SB1_2_22/buf_output[1] , \SB1_2_22/buf_output[0] , \SB1_2_22/i3[0] ,
         \SB1_2_22/i1_5 , \SB1_2_22/i1_7 , \SB1_2_22/i1[9] , \SB1_2_22/i0_0 ,
         \SB1_2_22/i0_4 , \SB1_2_22/i0[10] , \SB1_2_22/i0[9] ,
         \SB1_2_22/i0[8] , \SB1_2_22/i0[7] , \SB1_2_22/i0[6] ,
         \SB1_2_23/buf_output[5] , \SB1_2_23/buf_output[4] ,
         \SB1_2_23/buf_output[3] , \SB1_2_23/buf_output[2] ,
         \SB1_2_23/buf_output[1] , \SB1_2_23/buf_output[0] , \SB1_2_23/i3[0] ,
         \SB1_2_23/i1_5 , \SB1_2_23/i1_7 , \SB1_2_23/i1[9] , \SB1_2_23/i0_0 ,
         \SB1_2_23/i0_3 , \SB1_2_23/i0_4 , \SB1_2_23/i0[10] , \SB1_2_23/i0[9] ,
         \SB1_2_23/i0[8] , \SB1_2_23/i0[7] , \SB1_2_23/i0[6] ,
         \SB1_2_24/buf_output[5] , \SB1_2_24/buf_output[3] ,
         \SB1_2_24/buf_output[2] , \SB1_2_24/buf_output[1] ,
         \SB1_2_24/buf_output[0] , \SB1_2_24/i3[0] , \SB1_2_24/i1_5 ,
         \SB1_2_24/i1_7 , \SB1_2_24/i1[9] , \SB1_2_24/i0_0 , \SB1_2_24/i0_3 ,
         \SB1_2_24/i0_4 , \SB1_2_24/i0[10] , \SB1_2_24/i0[9] ,
         \SB1_2_24/i0[8] , \SB1_2_24/i0[7] , \SB1_2_24/i0[6] ,
         \SB1_2_25/buf_output[5] , \SB1_2_25/buf_output[4] ,
         \SB1_2_25/buf_output[3] , \SB1_2_25/buf_output[2] ,
         \SB1_2_25/buf_output[1] , \SB1_2_25/buf_output[0] , \SB1_2_25/i3[0] ,
         \SB1_2_25/i1_5 , \SB1_2_25/i1_7 , \SB1_2_25/i1[9] , \SB1_2_25/i0_0 ,
         \SB1_2_25/i0_3 , \SB1_2_25/i0_4 , \SB1_2_25/i0[10] , \SB1_2_25/i0[9] ,
         \SB1_2_25/i0[8] , \SB1_2_25/i0[7] , \SB1_2_25/i0[6] ,
         \SB1_2_26/buf_output[5] , \SB1_2_26/buf_output[4] ,
         \SB1_2_26/buf_output[3] , \SB1_2_26/buf_output[2] ,
         \SB1_2_26/buf_output[1] , \SB1_2_26/buf_output[0] , \SB1_2_26/i3[0] ,
         \SB1_2_26/i1_5 , \SB1_2_26/i1_7 , \SB1_2_26/i1[9] , \SB1_2_26/i0_0 ,
         \SB1_2_26/i0_3 , \SB1_2_26/i0_4 , \SB1_2_26/i0[10] , \SB1_2_26/i0[9] ,
         \SB1_2_26/i0[8] , \SB1_2_26/i0[7] , \SB1_2_26/i0[6] ,
         \SB1_2_27/buf_output[5] , \SB1_2_27/buf_output[3] ,
         \SB1_2_27/buf_output[2] , \SB1_2_27/buf_output[1] ,
         \SB1_2_27/buf_output[0] , \SB1_2_27/i3[0] , \SB1_2_27/i1_5 ,
         \SB1_2_27/i1_7 , \SB1_2_27/i1[9] , \SB1_2_27/i0_0 , \SB1_2_27/i0_3 ,
         \SB1_2_27/i0_4 , \SB1_2_27/i0[10] , \SB1_2_27/i0[9] ,
         \SB1_2_27/i0[8] , \SB1_2_27/i0[7] , \SB1_2_27/i0[6] ,
         \SB1_2_28/buf_output[5] , \SB1_2_28/buf_output[4] ,
         \SB1_2_28/buf_output[3] , \SB1_2_28/buf_output[2] ,
         \SB1_2_28/buf_output[1] , \SB1_2_28/buf_output[0] , \SB1_2_28/i3[0] ,
         \SB1_2_28/i1_5 , \SB1_2_28/i1_7 , \SB1_2_28/i1[9] , \SB1_2_28/i0_0 ,
         \SB1_2_28/i0_3 , \SB1_2_28/i0_4 , \SB1_2_28/i0[10] , \SB1_2_28/i0[9] ,
         \SB1_2_28/i0[8] , \SB1_2_28/i0[7] , \SB1_2_28/i0[6] ,
         \SB1_2_29/buf_output[5] , \SB1_2_29/buf_output[4] ,
         \SB1_2_29/buf_output[3] , \SB1_2_29/buf_output[2] ,
         \SB1_2_29/buf_output[1] , \SB1_2_29/buf_output[0] , \SB1_2_29/i3[0] ,
         \SB1_2_29/i1_5 , \SB1_2_29/i1_7 , \SB1_2_29/i1[9] , \SB1_2_29/i0_0 ,
         \SB1_2_29/i0_4 , \SB1_2_29/i0[10] , \SB1_2_29/i0[9] ,
         \SB1_2_29/i0[8] , \SB1_2_29/i0[7] , \SB1_2_29/i0[6] ,
         \SB1_2_30/buf_output[5] , \SB1_2_30/buf_output[4] ,
         \SB1_2_30/buf_output[3] , \SB1_2_30/buf_output[2] ,
         \SB1_2_30/buf_output[1] , \SB1_2_30/buf_output[0] , \SB1_2_30/i3[0] ,
         \SB1_2_30/i1_5 , \SB1_2_30/i1_7 , \SB1_2_30/i1[9] , \SB1_2_30/i0_0 ,
         \SB1_2_30/i0_3 , \SB1_2_30/i0_4 , \SB1_2_30/i0[10] , \SB1_2_30/i0[9] ,
         \SB1_2_30/i0[8] , \SB1_2_30/i0[7] , \SB1_2_30/i0[6] ,
         \SB1_2_31/buf_output[5] , \SB1_2_31/buf_output[4] ,
         \SB1_2_31/buf_output[3] , \SB1_2_31/buf_output[2] ,
         \SB1_2_31/buf_output[1] , \SB1_2_31/buf_output[0] , \SB1_2_31/i3[0] ,
         \SB1_2_31/i1_5 , \SB1_2_31/i1_7 , \SB1_2_31/i1[9] , \SB1_2_31/i0_0 ,
         \SB1_2_31/i0_3 , \SB1_2_31/i0_4 , \SB1_2_31/i0[10] , \SB1_2_31/i0[9] ,
         \SB1_2_31/i0[8] , \SB1_2_31/i0[7] , \SB1_2_31/i0[6] ,
         \SB2_2_0/buf_output[5] , \SB2_2_0/buf_output[4] ,
         \SB2_2_0/buf_output[3] , \SB2_2_0/buf_output[2] ,
         \SB2_2_0/buf_output[1] , \SB2_2_0/buf_output[0] , \SB2_2_0/i3[0] ,
         \SB2_2_0/i1_5 , \SB2_2_0/i1_7 , \SB2_2_0/i1[9] , \SB2_2_0/i0_0 ,
         \SB2_2_0/i0_3 , \SB2_2_0/i0[10] , \SB2_2_0/i0[9] , \SB2_2_0/i0[8] ,
         \SB2_2_0/i0[7] , \SB2_2_0/i0[6] , \SB2_2_1/buf_output[5] ,
         \SB2_2_1/buf_output[4] , \SB2_2_1/buf_output[3] ,
         \SB2_2_1/buf_output[2] , \SB2_2_1/buf_output[1] ,
         \SB2_2_1/buf_output[0] , \SB2_2_1/i3[0] , \SB2_2_1/i1_5 ,
         \SB2_2_1/i1_7 , \SB2_2_1/i1[9] , \SB2_2_1/i0_0 , \SB2_2_1/i0_3 ,
         \SB2_2_1/i0[10] , \SB2_2_1/i0[9] , \SB2_2_1/i0[8] , \SB2_2_1/i0[6] ,
         \SB2_2_2/buf_output[5] , \SB2_2_2/buf_output[4] ,
         \SB2_2_2/buf_output[3] , \SB2_2_2/buf_output[2] ,
         \SB2_2_2/buf_output[1] , \SB2_2_2/buf_output[0] , \SB2_2_2/i3[0] ,
         \SB2_2_2/i1_5 , \SB2_2_2/i1_7 , \SB2_2_2/i0_0 , \SB2_2_2/i0_3 ,
         \SB2_2_2/i0_4 , \SB2_2_2/i0[10] , \SB2_2_2/i0[9] , \SB2_2_2/i0[8] ,
         \SB2_2_2/i0[7] , \SB2_2_2/i0[6] , \SB2_2_3/buf_output[5] ,
         \SB2_2_3/buf_output[4] , \SB2_2_3/buf_output[3] ,
         \SB2_2_3/buf_output[2] , \SB2_2_3/buf_output[1] ,
         \SB2_2_3/buf_output[0] , \SB2_2_3/i3[0] , \SB2_2_3/i1_7 ,
         \SB2_2_3/i1[9] , \SB2_2_3/i0_0 , \SB2_2_3/i0_3 , \SB2_2_3/i0_4 ,
         \SB2_2_3/i0[10] , \SB2_2_3/i0[9] , \SB2_2_3/i0[7] , \SB2_2_3/i0[6] ,
         \SB2_2_4/buf_output[5] , \SB2_2_4/buf_output[4] ,
         \SB2_2_4/buf_output[3] , \SB2_2_4/buf_output[2] ,
         \SB2_2_4/buf_output[1] , \SB2_2_4/buf_output[0] , \SB2_2_4/i3[0] ,
         \SB2_2_4/i1_5 , \SB2_2_4/i1_7 , \SB2_2_4/i1[9] , \SB2_2_4/i0_0 ,
         \SB2_2_4/i0_3 , \SB2_2_4/i0_4 , \SB2_2_4/i0[10] , \SB2_2_4/i0[9] ,
         \SB2_2_4/i0[8] , \SB2_2_4/i0[7] , \SB2_2_4/i0[6] ,
         \SB2_2_5/buf_output[5] , \SB2_2_5/buf_output[4] ,
         \SB2_2_5/buf_output[3] , \SB2_2_5/buf_output[2] ,
         \SB2_2_5/buf_output[1] , \SB2_2_5/buf_output[0] , \SB2_2_5/i3[0] ,
         \SB2_2_5/i1_5 , \SB2_2_5/i1_7 , \SB2_2_5/i1[9] , \SB2_2_5/i0_0 ,
         \SB2_2_5/i0_3 , \SB2_2_5/i0_4 , \SB2_2_5/i0[10] , \SB2_2_5/i0[9] ,
         \SB2_2_5/i0[8] , \SB2_2_5/i0[7] , \SB2_2_5/i0[6] ,
         \SB2_2_6/buf_output[5] , \SB2_2_6/buf_output[4] ,
         \SB2_2_6/buf_output[3] , \SB2_2_6/buf_output[2] ,
         \SB2_2_6/buf_output[1] , \SB2_2_6/buf_output[0] , \SB2_2_6/i3[0] ,
         \SB2_2_6/i1_5 , \SB2_2_6/i1_7 , \SB2_2_6/i1[9] , \SB2_2_6/i0_0 ,
         \SB2_2_6/i0_3 , \SB2_2_6/i0_4 , \SB2_2_6/i0[10] , \SB2_2_6/i0[9] ,
         \SB2_2_6/i0[8] , \SB2_2_6/i0[7] , \SB2_2_6/i0[6] ,
         \SB2_2_7/buf_output[5] , \SB2_2_7/buf_output[4] ,
         \SB2_2_7/buf_output[3] , \SB2_2_7/buf_output[2] ,
         \SB2_2_7/buf_output[1] , \SB2_2_7/buf_output[0] , \SB2_2_7/i3[0] ,
         \SB2_2_7/i1_5 , \SB2_2_7/i1_7 , \SB2_2_7/i1[9] , \SB2_2_7/i0_0 ,
         \SB2_2_7/i0_3 , \SB2_2_7/i0_4 , \SB2_2_7/i0[10] , \SB2_2_7/i0[9] ,
         \SB2_2_7/i0[8] , \SB2_2_7/i0[7] , \SB2_2_7/i0[6] ,
         \SB2_2_8/buf_output[5] , \SB2_2_8/buf_output[4] ,
         \SB2_2_8/buf_output[3] , \SB2_2_8/buf_output[2] ,
         \SB2_2_8/buf_output[1] , \SB2_2_8/buf_output[0] , \SB2_2_8/i3[0] ,
         \SB2_2_8/i1_5 , \SB2_2_8/i1_7 , \SB2_2_8/i1[9] , \SB2_2_8/i0_0 ,
         \SB2_2_8/i0_3 , \SB2_2_8/i0_4 , \SB2_2_8/i0[10] , \SB2_2_8/i0[9] ,
         \SB2_2_8/i0[8] , \SB2_2_8/i0[7] , \SB2_2_8/i0[6] ,
         \SB2_2_9/buf_output[5] , \SB2_2_9/buf_output[4] ,
         \SB2_2_9/buf_output[3] , \SB2_2_9/buf_output[2] ,
         \SB2_2_9/buf_output[0] , \SB2_2_9/i3[0] , \SB2_2_9/i1_5 ,
         \SB2_2_9/i1_7 , \SB2_2_9/i1[9] , \SB2_2_9/i0_0 , \SB2_2_9/i0_3 ,
         \SB2_2_9/i0_4 , \SB2_2_9/i0[10] , \SB2_2_9/i0[9] , \SB2_2_9/i0[8] ,
         \SB2_2_9/i0[7] , \SB2_2_9/i0[6] , \SB2_2_10/buf_output[5] ,
         \SB2_2_10/buf_output[4] , \SB2_2_10/buf_output[3] ,
         \SB2_2_10/buf_output[2] , \SB2_2_10/buf_output[1] ,
         \SB2_2_10/buf_output[0] , \SB2_2_10/i3[0] , \SB2_2_10/i1_7 ,
         \SB2_2_10/i1[9] , \SB2_2_10/i0_0 , \SB2_2_10/i0_3 , \SB2_2_10/i0_4 ,
         \SB2_2_10/i0[10] , \SB2_2_10/i0[9] , \SB2_2_10/i0[8] ,
         \SB2_2_10/i0[7] , \SB2_2_10/i0[6] , \SB2_2_11/buf_output[5] ,
         \SB2_2_11/buf_output[4] , \SB2_2_11/buf_output[3] ,
         \SB2_2_11/buf_output[2] , \SB2_2_11/buf_output[1] ,
         \SB2_2_11/buf_output[0] , \SB2_2_11/i3[0] , \SB2_2_11/i1_5 ,
         \SB2_2_11/i1_7 , \SB2_2_11/i1[9] , \SB2_2_11/i0_0 , \SB2_2_11/i0_3 ,
         \SB2_2_11/i0_4 , \SB2_2_11/i0[10] , \SB2_2_11/i0[9] ,
         \SB2_2_11/i0[8] , \SB2_2_11/i0[7] , \SB2_2_11/i0[6] ,
         \SB2_2_12/buf_output[5] , \SB2_2_12/buf_output[4] ,
         \SB2_2_12/buf_output[3] , \SB2_2_12/buf_output[2] ,
         \SB2_2_12/buf_output[1] , \SB2_2_12/buf_output[0] , \SB2_2_12/i3[0] ,
         \SB2_2_12/i1_5 , \SB2_2_12/i1_7 , \SB2_2_12/i1[9] , \SB2_2_12/i0_0 ,
         \SB2_2_12/i0_3 , \SB2_2_12/i0_4 , \SB2_2_12/i0[10] , \SB2_2_12/i0[9] ,
         \SB2_2_12/i0[8] , \SB2_2_12/i0[7] , \SB2_2_12/i0[6] ,
         \SB2_2_13/buf_output[5] , \SB2_2_13/buf_output[4] ,
         \SB2_2_13/buf_output[3] , \SB2_2_13/buf_output[2] ,
         \SB2_2_13/buf_output[1] , \SB2_2_13/buf_output[0] , \SB2_2_13/i3[0] ,
         \SB2_2_13/i1_5 , \SB2_2_13/i1_7 , \SB2_2_13/i1[9] , \SB2_2_13/i0_0 ,
         \SB2_2_13/i0_3 , \SB2_2_13/i0_4 , \SB2_2_13/i0[10] , \SB2_2_13/i0[9] ,
         \SB2_2_13/i0[8] , \SB2_2_13/i0[7] , \SB2_2_13/i0[6] ,
         \SB2_2_14/buf_output[5] , \SB2_2_14/buf_output[4] ,
         \SB2_2_14/buf_output[3] , \SB2_2_14/buf_output[2] ,
         \SB2_2_14/buf_output[1] , \SB2_2_14/buf_output[0] , \SB2_2_14/i3[0] ,
         \SB2_2_14/i1_5 , \SB2_2_14/i1_7 , \SB2_2_14/i1[9] , \SB2_2_14/i0_0 ,
         \SB2_2_14/i0_3 , \SB2_2_14/i0_4 , \SB2_2_14/i0[10] , \SB2_2_14/i0[9] ,
         \SB2_2_14/i0[8] , \SB2_2_14/i0[7] , \SB2_2_14/i0[6] ,
         \SB2_2_15/buf_output[5] , \SB2_2_15/buf_output[4] ,
         \SB2_2_15/buf_output[3] , \SB2_2_15/buf_output[2] ,
         \SB2_2_15/buf_output[1] , \SB2_2_15/buf_output[0] , \SB2_2_15/i3[0] ,
         \SB2_2_15/i1_5 , \SB2_2_15/i1_7 , \SB2_2_15/i1[9] , \SB2_2_15/i0_0 ,
         \SB2_2_15/i0_3 , \SB2_2_15/i0_4 , \SB2_2_15/i0[10] , \SB2_2_15/i0[9] ,
         \SB2_2_15/i0[8] , \SB2_2_15/i0[7] , \SB2_2_15/i0[6] ,
         \SB2_2_16/buf_output[5] , \SB2_2_16/buf_output[4] ,
         \SB2_2_16/buf_output[3] , \SB2_2_16/buf_output[2] ,
         \SB2_2_16/buf_output[1] , \SB2_2_16/buf_output[0] , \SB2_2_16/i3[0] ,
         \SB2_2_16/i1_5 , \SB2_2_16/i1_7 , \SB2_2_16/i1[9] , \SB2_2_16/i0_0 ,
         \SB2_2_16/i0_3 , \SB2_2_16/i0_4 , \SB2_2_16/i0[10] , \SB2_2_16/i0[9] ,
         \SB2_2_16/i0[8] , \SB2_2_16/i0[7] , \SB2_2_16/i0[6] ,
         \SB2_2_17/buf_output[5] , \SB2_2_17/buf_output[4] ,
         \SB2_2_17/buf_output[3] , \SB2_2_17/buf_output[2] ,
         \SB2_2_17/buf_output[1] , \SB2_2_17/buf_output[0] , \SB2_2_17/i3[0] ,
         \SB2_2_17/i1_5 , \SB2_2_17/i1_7 , \SB2_2_17/i1[9] , \SB2_2_17/i0_0 ,
         \SB2_2_17/i0_3 , \SB2_2_17/i0[10] , \SB2_2_17/i0[9] ,
         \SB2_2_17/i0[8] , \SB2_2_17/i0[7] , \SB2_2_17/i0[6] ,
         \SB2_2_18/buf_output[5] , \SB2_2_18/buf_output[4] ,
         \SB2_2_18/buf_output[3] , \SB2_2_18/buf_output[2] ,
         \SB2_2_18/buf_output[1] , \SB2_2_18/buf_output[0] , \SB2_2_18/i3[0] ,
         \SB2_2_18/i1_5 , \SB2_2_18/i1_7 , \SB2_2_18/i1[9] , \SB2_2_18/i0_0 ,
         \SB2_2_18/i0_3 , \SB2_2_18/i0_4 , \SB2_2_18/i0[10] , \SB2_2_18/i0[9] ,
         \SB2_2_18/i0[8] , \SB2_2_18/i0[6] , \SB2_2_19/buf_output[5] ,
         \SB2_2_19/buf_output[4] , \SB2_2_19/buf_output[3] ,
         \SB2_2_19/buf_output[2] , \SB2_2_19/buf_output[1] ,
         \SB2_2_19/buf_output[0] , \SB2_2_19/i3[0] , \SB2_2_19/i1_5 ,
         \SB2_2_19/i1_7 , \SB2_2_19/i1[9] , \SB2_2_19/i0_0 , \SB2_2_19/i0_3 ,
         \SB2_2_19/i0_4 , \SB2_2_19/i0[10] , \SB2_2_19/i0[9] ,
         \SB2_2_19/i0[8] , \SB2_2_19/i0[7] , \SB2_2_19/i0[6] ,
         \SB2_2_20/buf_output[5] , \SB2_2_20/buf_output[4] ,
         \SB2_2_20/buf_output[3] , \SB2_2_20/buf_output[2] ,
         \SB2_2_20/buf_output[1] , \SB2_2_20/buf_output[0] , \SB2_2_20/i3[0] ,
         \SB2_2_20/i1_5 , \SB2_2_20/i1_7 , \SB2_2_20/i1[9] , \SB2_2_20/i0_0 ,
         \SB2_2_20/i0_3 , \SB2_2_20/i0_4 , \SB2_2_20/i0[10] , \SB2_2_20/i0[9] ,
         \SB2_2_20/i0[8] , \SB2_2_20/i0[7] , \SB2_2_20/i0[6] ,
         \SB2_2_21/buf_output[5] , \SB2_2_21/buf_output[4] ,
         \SB2_2_21/buf_output[3] , \SB2_2_21/buf_output[2] ,
         \SB2_2_21/buf_output[1] , \SB2_2_21/buf_output[0] , \SB2_2_21/i3[0] ,
         \SB2_2_21/i1_5 , \SB2_2_21/i1_7 , \SB2_2_21/i1[9] , \SB2_2_21/i0_0 ,
         \SB2_2_21/i0_3 , \SB2_2_21/i0[10] , \SB2_2_21/i0[9] ,
         \SB2_2_21/i0[8] , \SB2_2_21/i0[6] , \SB2_2_22/buf_output[5] ,
         \SB2_2_22/buf_output[4] , \SB2_2_22/buf_output[3] ,
         \SB2_2_22/buf_output[2] , \SB2_2_22/buf_output[1] ,
         \SB2_2_22/buf_output[0] , \SB2_2_22/i3[0] , \SB2_2_22/i1_5 ,
         \SB2_2_22/i1_7 , \SB2_2_22/i1[9] , \SB2_2_22/i0_0 , \SB2_2_22/i0_3 ,
         \SB2_2_22/i0_4 , \SB2_2_22/i0[10] , \SB2_2_22/i0[9] ,
         \SB2_2_22/i0[8] , \SB2_2_22/i0[7] , \SB2_2_22/i0[6] ,
         \SB2_2_23/buf_output[5] , \SB2_2_23/buf_output[4] ,
         \SB2_2_23/buf_output[3] , \SB2_2_23/buf_output[2] ,
         \SB2_2_23/buf_output[1] , \SB2_2_23/buf_output[0] , \SB2_2_23/i3[0] ,
         \SB2_2_23/i1_5 , \SB2_2_23/i1_7 , \SB2_2_23/i1[9] , \SB2_2_23/i0_0 ,
         \SB2_2_23/i0_3 , \SB2_2_23/i0_4 , \SB2_2_23/i0[10] , \SB2_2_23/i0[9] ,
         \SB2_2_23/i0[8] , \SB2_2_23/i0[7] , \SB2_2_23/i0[6] ,
         \SB2_2_24/buf_output[5] , \SB2_2_24/buf_output[4] ,
         \SB2_2_24/buf_output[3] , \SB2_2_24/buf_output[2] ,
         \SB2_2_24/buf_output[1] , \SB2_2_24/buf_output[0] , \SB2_2_24/i3[0] ,
         \SB2_2_24/i1_5 , \SB2_2_24/i1_7 , \SB2_2_24/i1[9] , \SB2_2_24/i0_0 ,
         \SB2_2_24/i0_3 , \SB2_2_24/i0_4 , \SB2_2_24/i0[10] , \SB2_2_24/i0[9] ,
         \SB2_2_24/i0[8] , \SB2_2_24/i0[7] , \SB2_2_24/i0[6] ,
         \SB2_2_25/buf_output[5] , \SB2_2_25/buf_output[4] ,
         \SB2_2_25/buf_output[3] , \SB2_2_25/buf_output[2] ,
         \SB2_2_25/buf_output[1] , \SB2_2_25/buf_output[0] , \SB2_2_25/i3[0] ,
         \SB2_2_25/i1_5 , \SB2_2_25/i1_7 , \SB2_2_25/i1[9] , \SB2_2_25/i0_0 ,
         \SB2_2_25/i0_3 , \SB2_2_25/i0_4 , \SB2_2_25/i0[10] , \SB2_2_25/i0[9] ,
         \SB2_2_25/i0[8] , \SB2_2_25/i0[7] , \SB2_2_25/i0[6] ,
         \SB2_2_26/buf_output[5] , \SB2_2_26/buf_output[4] ,
         \SB2_2_26/buf_output[3] , \SB2_2_26/buf_output[2] ,
         \SB2_2_26/buf_output[1] , \SB2_2_26/buf_output[0] , \SB2_2_26/i3[0] ,
         \SB2_2_26/i1_5 , \SB2_2_26/i1_7 , \SB2_2_26/i1[9] , \SB2_2_26/i0_0 ,
         \SB2_2_26/i0_3 , \SB2_2_26/i0_4 , \SB2_2_26/i0[10] , \SB2_2_26/i0[9] ,
         \SB2_2_26/i0[8] , \SB2_2_26/i0[7] , \SB2_2_26/i0[6] ,
         \SB2_2_27/buf_output[5] , \SB2_2_27/buf_output[4] ,
         \SB2_2_27/buf_output[3] , \SB2_2_27/buf_output[2] ,
         \SB2_2_27/buf_output[1] , \SB2_2_27/buf_output[0] , \SB2_2_27/i3[0] ,
         \SB2_2_27/i1_5 , \SB2_2_27/i1_7 , \SB2_2_27/i1[9] , \SB2_2_27/i0_0 ,
         \SB2_2_27/i0_3 , \SB2_2_27/i0_4 , \SB2_2_27/i0[10] , \SB2_2_27/i0[9] ,
         \SB2_2_27/i0[8] , \SB2_2_27/i0[7] , \SB2_2_27/i0[6] ,
         \SB2_2_28/buf_output[5] , \SB2_2_28/buf_output[4] ,
         \SB2_2_28/buf_output[3] , \SB2_2_28/buf_output[2] ,
         \SB2_2_28/buf_output[1] , \SB2_2_28/buf_output[0] , \SB2_2_28/i3[0] ,
         \SB2_2_28/i1_5 , \SB2_2_28/i1_7 , \SB2_2_28/i1[9] , \SB2_2_28/i0_0 ,
         \SB2_2_28/i0_3 , \SB2_2_28/i0_4 , \SB2_2_28/i0[10] , \SB2_2_28/i0[9] ,
         \SB2_2_28/i0[8] , \SB2_2_28/i0[7] , \SB2_2_28/i0[6] ,
         \SB2_2_29/buf_output[5] , \SB2_2_29/buf_output[4] ,
         \SB2_2_29/buf_output[3] , \SB2_2_29/buf_output[2] ,
         \SB2_2_29/buf_output[1] , \SB2_2_29/buf_output[0] , \SB2_2_29/i3[0] ,
         \SB2_2_29/i1_5 , \SB2_2_29/i1_7 , \SB2_2_29/i1[9] , \SB2_2_29/i0_0 ,
         \SB2_2_29/i0_3 , \SB2_2_29/i0_4 , \SB2_2_29/i0[10] , \SB2_2_29/i0[9] ,
         \SB2_2_29/i0[8] , \SB2_2_29/i0[7] , \SB2_2_29/i0[6] ,
         \SB2_2_30/buf_output[5] , \SB2_2_30/buf_output[4] ,
         \SB2_2_30/buf_output[3] , \SB2_2_30/buf_output[2] ,
         \SB2_2_30/buf_output[1] , \SB2_2_30/buf_output[0] , \SB2_2_30/i3[0] ,
         \SB2_2_30/i1_5 , \SB2_2_30/i1_7 , \SB2_2_30/i1[9] , \SB2_2_30/i0_0 ,
         \SB2_2_30/i0_3 , \SB2_2_30/i0_4 , \SB2_2_30/i0[10] , \SB2_2_30/i0[9] ,
         \SB2_2_30/i0[8] , \SB2_2_30/i0[7] , \SB2_2_30/i0[6] ,
         \SB2_2_31/buf_output[5] , \SB2_2_31/buf_output[4] ,
         \SB2_2_31/buf_output[3] , \SB2_2_31/buf_output[2] ,
         \SB2_2_31/buf_output[1] , \SB2_2_31/buf_output[0] , \SB2_2_31/i3[0] ,
         \SB2_2_31/i1_5 , \SB2_2_31/i1_7 , \SB2_2_31/i1[9] , \SB2_2_31/i0_0 ,
         \SB2_2_31/i0_3 , \SB2_2_31/i0_4 , \SB2_2_31/i0[10] , \SB2_2_31/i0[9] ,
         \SB2_2_31/i0[8] , \SB2_2_31/i0[7] , \SB2_2_31/i0[6] ,
         \SB1_3_0/buf_output[5] , \SB1_3_0/buf_output[4] ,
         \SB1_3_0/buf_output[3] , \SB1_3_0/buf_output[2] ,
         \SB1_3_0/buf_output[1] , \SB1_3_0/buf_output[0] , \SB1_3_0/i3[0] ,
         \SB1_3_0/i1_5 , \SB1_3_0/i1_7 , \SB1_3_0/i1[9] , \SB1_3_0/i0_0 ,
         \SB1_3_0/i0_3 , \SB1_3_0/i0_4 , \SB1_3_0/i0[10] , \SB1_3_0/i0[9] ,
         \SB1_3_0/i0[8] , \SB1_3_0/i0[7] , \SB1_3_0/i0[6] ,
         \SB1_3_1/buf_output[5] , \SB1_3_1/buf_output[4] ,
         \SB1_3_1/buf_output[3] , \SB1_3_1/buf_output[2] ,
         \SB1_3_1/buf_output[1] , \SB1_3_1/buf_output[0] , \SB1_3_1/i3[0] ,
         \SB1_3_1/i1_5 , \SB1_3_1/i1_7 , \SB1_3_1/i1[9] , \SB1_3_1/i0_0 ,
         \SB1_3_1/i0_3 , \SB1_3_1/i0_4 , \SB1_3_1/i0[10] , \SB1_3_1/i0[9] ,
         \SB1_3_1/i0[8] , \SB1_3_1/i0[7] , \SB1_3_1/i0[6] ,
         \SB1_3_2/buf_output[5] , \SB1_3_2/buf_output[4] ,
         \SB1_3_2/buf_output[3] , \SB1_3_2/buf_output[2] ,
         \SB1_3_2/buf_output[1] , \SB1_3_2/buf_output[0] , \SB1_3_2/i3[0] ,
         \SB1_3_2/i1_5 , \SB1_3_2/i1_7 , \SB1_3_2/i1[9] , \SB1_3_2/i0_0 ,
         \SB1_3_2/i0_3 , \SB1_3_2/i0_4 , \SB1_3_2/i0[10] , \SB1_3_2/i0[9] ,
         \SB1_3_2/i0[8] , \SB1_3_2/i0[7] , \SB1_3_2/i0[6] ,
         \SB1_3_3/buf_output[5] , \SB1_3_3/buf_output[4] ,
         \SB1_3_3/buf_output[3] , \SB1_3_3/buf_output[2] ,
         \SB1_3_3/buf_output[1] , \SB1_3_3/buf_output[0] , \SB1_3_3/i3[0] ,
         \SB1_3_3/i1_5 , \SB1_3_3/i1_7 , \SB1_3_3/i1[9] , \SB1_3_3/i0_0 ,
         \SB1_3_3/i0_3 , \SB1_3_3/i0_4 , \SB1_3_3/i0[10] , \SB1_3_3/i0[9] ,
         \SB1_3_3/i0[8] , \SB1_3_3/i0[7] , \SB1_3_3/i0[6] ,
         \SB1_3_4/buf_output[5] , \SB1_3_4/buf_output[4] ,
         \SB1_3_4/buf_output[3] , \SB1_3_4/buf_output[2] ,
         \SB1_3_4/buf_output[1] , \SB1_3_4/buf_output[0] , \SB1_3_4/i3[0] ,
         \SB1_3_4/i1_5 , \SB1_3_4/i1_7 , \SB1_3_4/i1[9] , \SB1_3_4/i0_0 ,
         \SB1_3_4/i0_4 , \SB1_3_4/i0[10] , \SB1_3_4/i0[9] , \SB1_3_4/i0[8] ,
         \SB1_3_4/i0[7] , \SB1_3_4/i0[6] , \SB1_3_5/buf_output[5] ,
         \SB1_3_5/buf_output[3] , \SB1_3_5/buf_output[2] ,
         \SB1_3_5/buf_output[1] , \SB1_3_5/buf_output[0] , \SB1_3_5/i3[0] ,
         \SB1_3_5/i1_5 , \SB1_3_5/i1_7 , \SB1_3_5/i1[9] , \SB1_3_5/i0_0 ,
         \SB1_3_5/i0_3 , \SB1_3_5/i0_4 , \SB1_3_5/i0[10] , \SB1_3_5/i0[9] ,
         \SB1_3_5/i0[8] , \SB1_3_5/i0[7] , \SB1_3_5/i0[6] ,
         \SB1_3_6/buf_output[5] , \SB1_3_6/buf_output[3] ,
         \SB1_3_6/buf_output[2] , \SB1_3_6/buf_output[1] ,
         \SB1_3_6/buf_output[0] , \SB1_3_6/i3[0] , \SB1_3_6/i1_5 ,
         \SB1_3_6/i1_7 , \SB1_3_6/i1[9] , \SB1_3_6/i0_0 , \SB1_3_6/i0_3 ,
         \SB1_3_6/i0_4 , \SB1_3_6/i0[10] , \SB1_3_6/i0[9] , \SB1_3_6/i0[8] ,
         \SB1_3_6/i0[7] , \SB1_3_6/i0[6] , \SB1_3_7/buf_output[5] ,
         \SB1_3_7/buf_output[4] , \SB1_3_7/buf_output[3] ,
         \SB1_3_7/buf_output[2] , \SB1_3_7/buf_output[1] ,
         \SB1_3_7/buf_output[0] , \SB1_3_7/i3[0] , \SB1_3_7/i1_5 ,
         \SB1_3_7/i1_7 , \SB1_3_7/i1[9] , \SB1_3_7/i0_0 , \SB1_3_7/i0_3 ,
         \SB1_3_7/i0_4 , \SB1_3_7/i0[10] , \SB1_3_7/i0[9] , \SB1_3_7/i0[8] ,
         \SB1_3_7/i0[7] , \SB1_3_7/i0[6] , \SB1_3_8/buf_output[3] ,
         \SB1_3_8/buf_output[2] , \SB1_3_8/buf_output[1] ,
         \SB1_3_8/buf_output[0] , \SB1_3_8/i3[0] , \SB1_3_8/i1_5 ,
         \SB1_3_8/i1_7 , \SB1_3_8/i1[9] , \SB1_3_8/i0_0 , \SB1_3_8/i0_3 ,
         \SB1_3_8/i0_4 , \SB1_3_8/i0[10] , \SB1_3_8/i0[9] , \SB1_3_8/i0[8] ,
         \SB1_3_8/i0[7] , \SB1_3_8/i0[6] , \SB1_3_9/buf_output[5] ,
         \SB1_3_9/buf_output[4] , \SB1_3_9/buf_output[3] ,
         \SB1_3_9/buf_output[2] , \SB1_3_9/buf_output[1] ,
         \SB1_3_9/buf_output[0] , \SB1_3_9/i3[0] , \SB1_3_9/i1_5 ,
         \SB1_3_9/i1_7 , \SB1_3_9/i1[9] , \SB1_3_9/i0_0 , \SB1_3_9/i0_3 ,
         \SB1_3_9/i0_4 , \SB1_3_9/i0[10] , \SB1_3_9/i0[8] , \SB1_3_9/i0[7] ,
         \SB1_3_9/i0[6] , \SB1_3_10/buf_output[5] , \SB1_3_10/buf_output[4] ,
         \SB1_3_10/buf_output[3] , \SB1_3_10/buf_output[2] ,
         \SB1_3_10/buf_output[1] , \SB1_3_10/buf_output[0] , \SB1_3_10/i3[0] ,
         \SB1_3_10/i1_5 , \SB1_3_10/i1_7 , \SB1_3_10/i1[9] , \SB1_3_10/i0_0 ,
         \SB1_3_10/i0_3 , \SB1_3_10/i0_4 , \SB1_3_10/i0[10] , \SB1_3_10/i0[9] ,
         \SB1_3_10/i0[8] , \SB1_3_10/i0[7] , \SB1_3_10/i0[6] ,
         \SB1_3_11/buf_output[5] , \SB1_3_11/buf_output[3] ,
         \SB1_3_11/buf_output[2] , \SB1_3_11/buf_output[1] ,
         \SB1_3_11/buf_output[0] , \SB1_3_11/i3[0] , \SB1_3_11/i1_5 ,
         \SB1_3_11/i1_7 , \SB1_3_11/i1[9] , \SB1_3_11/i0_0 , \SB1_3_11/i0_3 ,
         \SB1_3_11/i0_4 , \SB1_3_11/i0[10] , \SB1_3_11/i0[9] ,
         \SB1_3_11/i0[8] , \SB1_3_11/i0[7] , \SB1_3_11/i0[6] ,
         \SB1_3_12/buf_output[5] , \SB1_3_12/buf_output[4] ,
         \SB1_3_12/buf_output[3] , \SB1_3_12/buf_output[2] ,
         \SB1_3_12/buf_output[1] , \SB1_3_12/buf_output[0] , \SB1_3_12/i3[0] ,
         \SB1_3_12/i1_5 , \SB1_3_12/i1_7 , \SB1_3_12/i1[9] , \SB1_3_12/i0_0 ,
         \SB1_3_12/i0_3 , \SB1_3_12/i0_4 , \SB1_3_12/i0[10] , \SB1_3_12/i0[9] ,
         \SB1_3_12/i0[8] , \SB1_3_12/i0[7] , \SB1_3_12/i0[6] ,
         \SB1_3_13/buf_output[5] , \SB1_3_13/buf_output[3] ,
         \SB1_3_13/buf_output[2] , \SB1_3_13/buf_output[1] ,
         \SB1_3_13/buf_output[0] , \SB1_3_13/i3[0] , \SB1_3_13/i1_5 ,
         \SB1_3_13/i1_7 , \SB1_3_13/i1[9] , \SB1_3_13/i0_0 , \SB1_3_13/i0_3 ,
         \SB1_3_13/i0_4 , \SB1_3_13/i0[10] , \SB1_3_13/i0[9] ,
         \SB1_3_13/i0[8] , \SB1_3_13/i0[7] , \SB1_3_13/i0[6] ,
         \SB1_3_14/buf_output[5] , \SB1_3_14/buf_output[3] ,
         \SB1_3_14/buf_output[2] , \SB1_3_14/buf_output[1] ,
         \SB1_3_14/buf_output[0] , \SB1_3_14/i3[0] , \SB1_3_14/i1_5 ,
         \SB1_3_14/i1_7 , \SB1_3_14/i1[9] , \SB1_3_14/i0_0 , \SB1_3_14/i0_4 ,
         \SB1_3_14/i0[10] , \SB1_3_14/i0[9] , \SB1_3_14/i0[8] ,
         \SB1_3_14/i0[7] , \SB1_3_14/i0[6] , \SB1_3_15/buf_output[5] ,
         \SB1_3_15/buf_output[4] , \SB1_3_15/buf_output[3] ,
         \SB1_3_15/buf_output[2] , \SB1_3_15/buf_output[1] ,
         \SB1_3_15/buf_output[0] , \SB1_3_15/i3[0] , \SB1_3_15/i1_5 ,
         \SB1_3_15/i1_7 , \SB1_3_15/i1[9] , \SB1_3_15/i0_0 , \SB1_3_15/i0_3 ,
         \SB1_3_15/i0_4 , \SB1_3_15/i0[10] , \SB1_3_15/i0[9] ,
         \SB1_3_15/i0[8] , \SB1_3_15/i0[7] , \SB1_3_15/i0[6] ,
         \SB1_3_16/buf_output[5] , \SB1_3_16/buf_output[4] ,
         \SB1_3_16/buf_output[3] , \SB1_3_16/buf_output[2] ,
         \SB1_3_16/buf_output[1] , \SB1_3_16/buf_output[0] , \SB1_3_16/i3[0] ,
         \SB1_3_16/i1_5 , \SB1_3_16/i1_7 , \SB1_3_16/i1[9] , \SB1_3_16/i0_0 ,
         \SB1_3_16/i0_3 , \SB1_3_16/i0_4 , \SB1_3_16/i0[10] , \SB1_3_16/i0[8] ,
         \SB1_3_16/i0[7] , \SB1_3_16/i0[6] , \SB1_3_17/buf_output[5] ,
         \SB1_3_17/buf_output[4] , \SB1_3_17/buf_output[3] ,
         \SB1_3_17/buf_output[2] , \SB1_3_17/buf_output[1] ,
         \SB1_3_17/buf_output[0] , \SB1_3_17/i3[0] , \SB1_3_17/i1_5 ,
         \SB1_3_17/i1_7 , \SB1_3_17/i1[9] , \SB1_3_17/i0_0 , \SB1_3_17/i0_3 ,
         \SB1_3_17/i0_4 , \SB1_3_17/i0[10] , \SB1_3_17/i0[9] ,
         \SB1_3_17/i0[8] , \SB1_3_17/i0[7] , \SB1_3_17/i0[6] ,
         \SB1_3_18/buf_output[5] , \SB1_3_18/buf_output[4] ,
         \SB1_3_18/buf_output[3] , \SB1_3_18/buf_output[2] ,
         \SB1_3_18/buf_output[1] , \SB1_3_18/buf_output[0] , \SB1_3_18/i3[0] ,
         \SB1_3_18/i1_5 , \SB1_3_18/i1_7 , \SB1_3_18/i1[9] , \SB1_3_18/i0_0 ,
         \SB1_3_18/i0_3 , \SB1_3_18/i0_4 , \SB1_3_18/i0[10] , \SB1_3_18/i0[9] ,
         \SB1_3_18/i0[8] , \SB1_3_18/i0[7] , \SB1_3_18/i0[6] ,
         \SB1_3_19/buf_output[5] , \SB1_3_19/buf_output[4] ,
         \SB1_3_19/buf_output[3] , \SB1_3_19/buf_output[2] ,
         \SB1_3_19/buf_output[1] , \SB1_3_19/buf_output[0] , \SB1_3_19/i3[0] ,
         \SB1_3_19/i1_5 , \SB1_3_19/i1_7 , \SB1_3_19/i1[9] , \SB1_3_19/i0_0 ,
         \SB1_3_19/i0_3 , \SB1_3_19/i0_4 , \SB1_3_19/i0[10] , \SB1_3_19/i0[9] ,
         \SB1_3_19/i0[8] , \SB1_3_19/i0[7] , \SB1_3_19/i0[6] ,
         \SB1_3_20/buf_output[5] , \SB1_3_20/buf_output[4] ,
         \SB1_3_20/buf_output[3] , \SB1_3_20/buf_output[2] ,
         \SB1_3_20/buf_output[1] , \SB1_3_20/buf_output[0] , \SB1_3_20/i3[0] ,
         \SB1_3_20/i1_5 , \SB1_3_20/i1_7 , \SB1_3_20/i1[9] , \SB1_3_20/i0_0 ,
         \SB1_3_20/i0_3 , \SB1_3_20/i0_4 , \SB1_3_20/i0[10] , \SB1_3_20/i0[9] ,
         \SB1_3_20/i0[8] , \SB1_3_20/i0[7] , \SB1_3_20/i0[6] ,
         \SB1_3_21/buf_output[5] , \SB1_3_21/buf_output[3] ,
         \SB1_3_21/buf_output[2] , \SB1_3_21/buf_output[1] ,
         \SB1_3_21/buf_output[0] , \SB1_3_21/i3[0] , \SB1_3_21/i1_5 ,
         \SB1_3_21/i1_7 , \SB1_3_21/i1[9] , \SB1_3_21/i0_0 , \SB1_3_21/i0_3 ,
         \SB1_3_21/i0_4 , \SB1_3_21/i0[10] , \SB1_3_21/i0[9] ,
         \SB1_3_21/i0[8] , \SB1_3_21/i0[7] , \SB1_3_21/i0[6] ,
         \SB1_3_22/buf_output[5] , \SB1_3_22/buf_output[3] ,
         \SB1_3_22/buf_output[2] , \SB1_3_22/buf_output[1] ,
         \SB1_3_22/buf_output[0] , \SB1_3_22/i3[0] , \SB1_3_22/i1_5 ,
         \SB1_3_22/i1_7 , \SB1_3_22/i1[9] , \SB1_3_22/i0_0 , \SB1_3_22/i0_3 ,
         \SB1_3_22/i0_4 , \SB1_3_22/i0[10] , \SB1_3_22/i0[9] ,
         \SB1_3_22/i0[8] , \SB1_3_22/i0[7] , \SB1_3_22/i0[6] ,
         \SB1_3_23/buf_output[5] , \SB1_3_23/buf_output[3] ,
         \SB1_3_23/buf_output[2] , \SB1_3_23/buf_output[1] ,
         \SB1_3_23/buf_output[0] , \SB1_3_23/i3[0] , \SB1_3_23/i1_5 ,
         \SB1_3_23/i1_7 , \SB1_3_23/i1[9] , \SB1_3_23/i0_0 , \SB1_3_23/i0_3 ,
         \SB1_3_23/i0_4 , \SB1_3_23/i0[10] , \SB1_3_23/i0[9] ,
         \SB1_3_23/i0[8] , \SB1_3_23/i0[7] , \SB1_3_23/i0[6] ,
         \SB1_3_24/buf_output[5] , \SB1_3_24/buf_output[4] ,
         \SB1_3_24/buf_output[3] , \SB1_3_24/buf_output[2] ,
         \SB1_3_24/buf_output[1] , \SB1_3_24/buf_output[0] , \SB1_3_24/i3[0] ,
         \SB1_3_24/i1_5 , \SB1_3_24/i1_7 , \SB1_3_24/i1[9] , \SB1_3_24/i0_0 ,
         \SB1_3_24/i0_3 , \SB1_3_24/i0_4 , \SB1_3_24/i0[10] , \SB1_3_24/i0[9] ,
         \SB1_3_24/i0[8] , \SB1_3_24/i0[7] , \SB1_3_24/i0[6] ,
         \SB1_3_25/buf_output[5] , \SB1_3_25/buf_output[4] ,
         \SB1_3_25/buf_output[3] , \SB1_3_25/buf_output[2] ,
         \SB1_3_25/buf_output[1] , \SB1_3_25/buf_output[0] , \SB1_3_25/i3[0] ,
         \SB1_3_25/i1_5 , \SB1_3_25/i1_7 , \SB1_3_25/i1[9] , \SB1_3_25/i0_0 ,
         \SB1_3_25/i0_3 , \SB1_3_25/i0_4 , \SB1_3_25/i0[10] , \SB1_3_25/i0[9] ,
         \SB1_3_25/i0[8] , \SB1_3_25/i0[7] , \SB1_3_25/i0[6] ,
         \SB1_3_26/buf_output[5] , \SB1_3_26/buf_output[4] ,
         \SB1_3_26/buf_output[3] , \SB1_3_26/buf_output[2] ,
         \SB1_3_26/buf_output[1] , \SB1_3_26/buf_output[0] , \SB1_3_26/i3[0] ,
         \SB1_3_26/i1_5 , \SB1_3_26/i1_7 , \SB1_3_26/i1[9] , \SB1_3_26/i0_0 ,
         \SB1_3_26/i0_3 , \SB1_3_26/i0_4 , \SB1_3_26/i0[10] , \SB1_3_26/i0[9] ,
         \SB1_3_26/i0[8] , \SB1_3_26/i0[7] , \SB1_3_26/i0[6] ,
         \SB1_3_27/buf_output[5] , \SB1_3_27/buf_output[3] ,
         \SB1_3_27/buf_output[2] , \SB1_3_27/buf_output[1] ,
         \SB1_3_27/buf_output[0] , \SB1_3_27/i3[0] , \SB1_3_27/i1_5 ,
         \SB1_3_27/i1_7 , \SB1_3_27/i1[9] , \SB1_3_27/i0_0 , \SB1_3_27/i0_3 ,
         \SB1_3_27/i0_4 , \SB1_3_27/i0[10] , \SB1_3_27/i0[9] ,
         \SB1_3_27/i0[8] , \SB1_3_27/i0[7] , \SB1_3_27/i0[6] ,
         \SB1_3_28/buf_output[5] , \SB1_3_28/buf_output[4] ,
         \SB1_3_28/buf_output[3] , \SB1_3_28/buf_output[2] ,
         \SB1_3_28/buf_output[1] , \SB1_3_28/buf_output[0] , \SB1_3_28/i3[0] ,
         \SB1_3_28/i1_5 , \SB1_3_28/i1_7 , \SB1_3_28/i1[9] , \SB1_3_28/i0_0 ,
         \SB1_3_28/i0_3 , \SB1_3_28/i0_4 , \SB1_3_28/i0[10] , \SB1_3_28/i0[9] ,
         \SB1_3_28/i0[8] , \SB1_3_28/i0[7] , \SB1_3_28/i0[6] ,
         \SB1_3_29/buf_output[5] , \SB1_3_29/buf_output[4] ,
         \SB1_3_29/buf_output[3] , \SB1_3_29/buf_output[2] ,
         \SB1_3_29/buf_output[1] , \SB1_3_29/buf_output[0] , \SB1_3_29/i3[0] ,
         \SB1_3_29/i1_5 , \SB1_3_29/i1_7 , \SB1_3_29/i1[9] , \SB1_3_29/i0_0 ,
         \SB1_3_29/i0_3 , \SB1_3_29/i0_4 , \SB1_3_29/i0[10] , \SB1_3_29/i0[9] ,
         \SB1_3_29/i0[8] , \SB1_3_29/i0[7] , \SB1_3_29/i0[6] ,
         \SB1_3_30/buf_output[5] , \SB1_3_30/buf_output[3] ,
         \SB1_3_30/buf_output[2] , \SB1_3_30/buf_output[1] ,
         \SB1_3_30/buf_output[0] , \SB1_3_30/i3[0] , \SB1_3_30/i1_5 ,
         \SB1_3_30/i1_7 , \SB1_3_30/i1[9] , \SB1_3_30/i0_0 , \SB1_3_30/i0_3 ,
         \SB1_3_30/i0_4 , \SB1_3_30/i0[10] , \SB1_3_30/i0[9] ,
         \SB1_3_30/i0[8] , \SB1_3_30/i0[7] , \SB1_3_30/i0[6] ,
         \SB1_3_31/buf_output[5] , \SB1_3_31/buf_output[4] ,
         \SB1_3_31/buf_output[3] , \SB1_3_31/buf_output[2] ,
         \SB1_3_31/buf_output[1] , \SB1_3_31/buf_output[0] , \SB1_3_31/i3[0] ,
         \SB1_3_31/i1_5 , \SB1_3_31/i1_7 , \SB1_3_31/i1[9] , \SB1_3_31/i0_0 ,
         \SB1_3_31/i0_3 , \SB1_3_31/i0_4 , \SB1_3_31/i0[10] , \SB1_3_31/i0[9] ,
         \SB1_3_31/i0[7] , \SB1_3_31/i0[6] , \SB2_3_0/buf_output[5] ,
         \SB2_3_0/buf_output[4] , \SB2_3_0/buf_output[3] ,
         \SB2_3_0/buf_output[2] , \SB2_3_0/buf_output[1] ,
         \SB2_3_0/buf_output[0] , \SB2_3_0/i3[0] , \SB2_3_0/i1_5 ,
         \SB2_3_0/i1_7 , \SB2_3_0/i1[9] , \SB2_3_0/i0_0 , \SB2_3_0/i0_3 ,
         \SB2_3_0/i0_4 , \SB2_3_0/i0[10] , \SB2_3_0/i0[9] , \SB2_3_0/i0[8] ,
         \SB2_3_0/i0[7] , \SB2_3_0/i0[6] , \SB2_3_1/buf_output[5] ,
         \SB2_3_1/buf_output[4] , \SB2_3_1/buf_output[3] ,
         \SB2_3_1/buf_output[2] , \SB2_3_1/buf_output[1] ,
         \SB2_3_1/buf_output[0] , \SB2_3_1/i3[0] , \SB2_3_1/i1_5 ,
         \SB2_3_1/i1_7 , \SB2_3_1/i1[9] , \SB2_3_1/i0_0 , \SB2_3_1/i0_3 ,
         \SB2_3_1/i0_4 , \SB2_3_1/i0[10] , \SB2_3_1/i0[9] , \SB2_3_1/i0[8] ,
         \SB2_3_1/i0[7] , \SB2_3_1/i0[6] , \SB2_3_2/buf_output[5] ,
         \SB2_3_2/buf_output[4] , \SB2_3_2/buf_output[3] ,
         \SB2_3_2/buf_output[2] , \SB2_3_2/buf_output[1] ,
         \SB2_3_2/buf_output[0] , \SB2_3_2/i3[0] , \SB2_3_2/i1_5 ,
         \SB2_3_2/i1_7 , \SB2_3_2/i1[9] , \SB2_3_2/i0_0 , \SB2_3_2/i0_3 ,
         \SB2_3_2/i0_4 , \SB2_3_2/i0[10] , \SB2_3_2/i0[9] , \SB2_3_2/i0[8] ,
         \SB2_3_2/i0[7] , \SB2_3_2/i0[6] , \SB2_3_3/buf_output[5] ,
         \SB2_3_3/buf_output[4] , \SB2_3_3/buf_output[3] ,
         \SB2_3_3/buf_output[2] , \SB2_3_3/buf_output[1] ,
         \SB2_3_3/buf_output[0] , \SB2_3_3/i3[0] , \SB2_3_3/i1_5 ,
         \SB2_3_3/i1_7 , \SB2_3_3/i1[9] , \SB2_3_3/i0_0 , \SB2_3_3/i0_3 ,
         \SB2_3_3/i0_4 , \SB2_3_3/i0[10] , \SB2_3_3/i0[9] , \SB2_3_3/i0[8] ,
         \SB2_3_3/i0[7] , \SB2_3_3/i0[6] , \SB2_3_4/buf_output[5] ,
         \SB2_3_4/buf_output[4] , \SB2_3_4/buf_output[3] ,
         \SB2_3_4/buf_output[2] , \SB2_3_4/buf_output[1] ,
         \SB2_3_4/buf_output[0] , \SB2_3_4/i3[0] , \SB2_3_4/i1_5 ,
         \SB2_3_4/i1_7 , \SB2_3_4/i1[9] , \SB2_3_4/i0_0 , \SB2_3_4/i0_3 ,
         \SB2_3_4/i0_4 , \SB2_3_4/i0[10] , \SB2_3_4/i0[9] , \SB2_3_4/i0[8] ,
         \SB2_3_4/i0[7] , \SB2_3_4/i0[6] , \SB2_3_5/buf_output[5] ,
         \SB2_3_5/buf_output[4] , \SB2_3_5/buf_output[3] ,
         \SB2_3_5/buf_output[2] , \SB2_3_5/buf_output[1] ,
         \SB2_3_5/buf_output[0] , \SB2_3_5/i3[0] , \SB2_3_5/i1_5 ,
         \SB2_3_5/i1_7 , \SB2_3_5/i1[9] , \SB2_3_5/i0_0 , \SB2_3_5/i0_3 ,
         \SB2_3_5/i0_4 , \SB2_3_5/i0[10] , \SB2_3_5/i0[9] , \SB2_3_5/i0[8] ,
         \SB2_3_5/i0[7] , \SB2_3_5/i0[6] , \SB2_3_6/buf_output[5] ,
         \SB2_3_6/buf_output[4] , \SB2_3_6/buf_output[3] ,
         \SB2_3_6/buf_output[2] , \SB2_3_6/buf_output[1] ,
         \SB2_3_6/buf_output[0] , \SB2_3_6/i3[0] , \SB2_3_6/i1_5 ,
         \SB2_3_6/i1_7 , \SB2_3_6/i1[9] , \SB2_3_6/i0_0 , \SB2_3_6/i0_3 ,
         \SB2_3_6/i0_4 , \SB2_3_6/i0[10] , \SB2_3_6/i0[9] , \SB2_3_6/i0[8] ,
         \SB2_3_6/i0[7] , \SB2_3_6/i0[6] , \SB2_3_7/buf_output[5] ,
         \SB2_3_7/buf_output[4] , \SB2_3_7/buf_output[3] ,
         \SB2_3_7/buf_output[2] , \SB2_3_7/buf_output[1] ,
         \SB2_3_7/buf_output[0] , \SB2_3_7/i3[0] , \SB2_3_7/i1_5 ,
         \SB2_3_7/i1_7 , \SB2_3_7/i1[9] , \SB2_3_7/i0_0 , \SB2_3_7/i0_3 ,
         \SB2_3_7/i0_4 , \SB2_3_7/i0[10] , \SB2_3_7/i0[9] , \SB2_3_7/i0[8] ,
         \SB2_3_7/i0[7] , \SB2_3_7/i0[6] , \SB2_3_8/buf_output[5] ,
         \SB2_3_8/buf_output[4] , \SB2_3_8/buf_output[3] ,
         \SB2_3_8/buf_output[2] , \SB2_3_8/buf_output[1] ,
         \SB2_3_8/buf_output[0] , \SB2_3_8/i3[0] , \SB2_3_8/i1_5 ,
         \SB2_3_8/i1_7 , \SB2_3_8/i1[9] , \SB2_3_8/i0_0 , \SB2_3_8/i0_3 ,
         \SB2_3_8/i0_4 , \SB2_3_8/i0[10] , \SB2_3_8/i0[9] , \SB2_3_8/i0[8] ,
         \SB2_3_8/i0[7] , \SB2_3_8/i0[6] , \SB2_3_9/buf_output[5] ,
         \SB2_3_9/buf_output[4] , \SB2_3_9/buf_output[3] ,
         \SB2_3_9/buf_output[2] , \SB2_3_9/buf_output[1] ,
         \SB2_3_9/buf_output[0] , \SB2_3_9/i3[0] , \SB2_3_9/i1_5 ,
         \SB2_3_9/i1_7 , \SB2_3_9/i1[9] , \SB2_3_9/i0_0 , \SB2_3_9/i0_3 ,
         \SB2_3_9/i0[10] , \SB2_3_9/i0[9] , \SB2_3_9/i0[8] , \SB2_3_9/i0[6] ,
         \SB2_3_10/buf_output[5] , \SB2_3_10/buf_output[4] ,
         \SB2_3_10/buf_output[3] , \SB2_3_10/buf_output[2] ,
         \SB2_3_10/buf_output[1] , \SB2_3_10/buf_output[0] , \SB2_3_10/i3[0] ,
         \SB2_3_10/i1_5 , \SB2_3_10/i1_7 , \SB2_3_10/i1[9] , \SB2_3_10/i0_0 ,
         \SB2_3_10/i0_3 , \SB2_3_10/i0_4 , \SB2_3_10/i0[10] , \SB2_3_10/i0[9] ,
         \SB2_3_10/i0[8] , \SB2_3_10/i0[7] , \SB2_3_10/i0[6] ,
         \SB2_3_11/buf_output[5] , \SB2_3_11/buf_output[4] ,
         \SB2_3_11/buf_output[3] , \SB2_3_11/buf_output[2] ,
         \SB2_3_11/buf_output[1] , \SB2_3_11/buf_output[0] , \SB2_3_11/i3[0] ,
         \SB2_3_11/i1_5 , \SB2_3_11/i1_7 , \SB2_3_11/i1[9] , \SB2_3_11/i0_0 ,
         \SB2_3_11/i0_3 , \SB2_3_11/i0_4 , \SB2_3_11/i0[10] , \SB2_3_11/i0[9] ,
         \SB2_3_11/i0[8] , \SB2_3_11/i0[7] , \SB2_3_11/i0[6] ,
         \SB2_3_12/buf_output[5] , \SB2_3_12/buf_output[4] ,
         \SB2_3_12/buf_output[3] , \SB2_3_12/buf_output[2] ,
         \SB2_3_12/buf_output[1] , \SB2_3_12/buf_output[0] , \SB2_3_12/i3[0] ,
         \SB2_3_12/i1_5 , \SB2_3_12/i1_7 , \SB2_3_12/i1[9] , \SB2_3_12/i0_0 ,
         \SB2_3_12/i0_3 , \SB2_3_12/i0[10] , \SB2_3_12/i0[9] ,
         \SB2_3_12/i0[8] , \SB2_3_12/i0[6] , \SB2_3_13/buf_output[5] ,
         \SB2_3_13/buf_output[4] , \SB2_3_13/buf_output[2] ,
         \SB2_3_13/buf_output[1] , \SB2_3_13/buf_output[0] , \SB2_3_13/i3[0] ,
         \SB2_3_13/i1_5 , \SB2_3_13/i1_7 , \SB2_3_13/i1[9] , \SB2_3_13/i0_0 ,
         \SB2_3_13/i0_3 , \SB2_3_13/i0_4 , \SB2_3_13/i0[10] , \SB2_3_13/i0[9] ,
         \SB2_3_13/i0[8] , \SB2_3_13/i0[7] , \SB2_3_13/i0[6] ,
         \SB2_3_14/buf_output[5] , \SB2_3_14/buf_output[4] ,
         \SB2_3_14/buf_output[3] , \SB2_3_14/buf_output[2] ,
         \SB2_3_14/buf_output[1] , \SB2_3_14/buf_output[0] , \SB2_3_14/i3[0] ,
         \SB2_3_14/i1_5 , \SB2_3_14/i1_7 , \SB2_3_14/i1[9] , \SB2_3_14/i0_0 ,
         \SB2_3_14/i0_3 , \SB2_3_14/i0_4 , \SB2_3_14/i0[10] , \SB2_3_14/i0[9] ,
         \SB2_3_14/i0[8] , \SB2_3_14/i0[7] , \SB2_3_14/i0[6] ,
         \SB2_3_15/buf_output[5] , \SB2_3_15/buf_output[4] ,
         \SB2_3_15/buf_output[3] , \SB2_3_15/buf_output[2] ,
         \SB2_3_15/buf_output[1] , \SB2_3_15/buf_output[0] , \SB2_3_15/i3[0] ,
         \SB2_3_15/i1_5 , \SB2_3_15/i1_7 , \SB2_3_15/i1[9] , \SB2_3_15/i0_0 ,
         \SB2_3_15/i0_3 , \SB2_3_15/i0_4 , \SB2_3_15/i0[10] , \SB2_3_15/i0[9] ,
         \SB2_3_15/i0[8] , \SB2_3_15/i0[7] , \SB2_3_15/i0[6] ,
         \SB2_3_16/buf_output[5] , \SB2_3_16/buf_output[4] ,
         \SB2_3_16/buf_output[3] , \SB2_3_16/buf_output[2] ,
         \SB2_3_16/buf_output[1] , \SB2_3_16/buf_output[0] , \SB2_3_16/i3[0] ,
         \SB2_3_16/i1_7 , \SB2_3_16/i1[9] , \SB2_3_16/i0_0 , \SB2_3_16/i0_3 ,
         \SB2_3_16/i0_4 , \SB2_3_16/i0[10] , \SB2_3_16/i0[9] ,
         \SB2_3_16/i0[8] , \SB2_3_16/i0[7] , \SB2_3_16/i0[6] ,
         \SB2_3_17/buf_output[5] , \SB2_3_17/buf_output[4] ,
         \SB2_3_17/buf_output[3] , \SB2_3_17/buf_output[2] ,
         \SB2_3_17/buf_output[1] , \SB2_3_17/buf_output[0] , \SB2_3_17/i3[0] ,
         \SB2_3_17/i1_5 , \SB2_3_17/i1_7 , \SB2_3_17/i1[9] , \SB2_3_17/i0_0 ,
         \SB2_3_17/i0_3 , \SB2_3_17/i0_4 , \SB2_3_17/i0[10] , \SB2_3_17/i0[9] ,
         \SB2_3_17/i0[8] , \SB2_3_17/i0[7] , \SB2_3_17/i0[6] ,
         \SB2_3_18/buf_output[5] , \SB2_3_18/buf_output[4] ,
         \SB2_3_18/buf_output[3] , \SB2_3_18/buf_output[2] ,
         \SB2_3_18/buf_output[1] , \SB2_3_18/buf_output[0] , \SB2_3_18/i3[0] ,
         \SB2_3_18/i1_5 , \SB2_3_18/i1_7 , \SB2_3_18/i1[9] , \SB2_3_18/i0_0 ,
         \SB2_3_18/i0_3 , \SB2_3_18/i0_4 , \SB2_3_18/i0[10] , \SB2_3_18/i0[9] ,
         \SB2_3_18/i0[8] , \SB2_3_18/i0[7] , \SB2_3_18/i0[6] ,
         \SB2_3_19/buf_output[5] , \SB2_3_19/buf_output[4] ,
         \SB2_3_19/buf_output[3] , \SB2_3_19/buf_output[2] ,
         \SB2_3_19/buf_output[1] , \SB2_3_19/buf_output[0] , \SB2_3_19/i3[0] ,
         \SB2_3_19/i1_5 , \SB2_3_19/i1_7 , \SB2_3_19/i1[9] , \SB2_3_19/i0_0 ,
         \SB2_3_19/i0_3 , \SB2_3_19/i0[10] , \SB2_3_19/i0[9] ,
         \SB2_3_19/i0[8] , \SB2_3_19/i0[7] , \SB2_3_19/i0[6] ,
         \SB2_3_20/buf_output[5] , \SB2_3_20/buf_output[4] ,
         \SB2_3_20/buf_output[3] , \SB2_3_20/buf_output[2] ,
         \SB2_3_20/buf_output[0] , \SB2_3_20/i3[0] , \SB2_3_20/i1_7 ,
         \SB2_3_20/i1[9] , \SB2_3_20/i0_0 , \SB2_3_20/i0_3 , \SB2_3_20/i0[10] ,
         \SB2_3_20/i0[9] , \SB2_3_20/i0[8] , \SB2_3_20/i0[7] ,
         \SB2_3_20/i0[6] , \SB2_3_21/buf_output[5] , \SB2_3_21/buf_output[4] ,
         \SB2_3_21/buf_output[3] , \SB2_3_21/buf_output[2] ,
         \SB2_3_21/buf_output[1] , \SB2_3_21/buf_output[0] , \SB2_3_21/i3[0] ,
         \SB2_3_21/i1_5 , \SB2_3_21/i1_7 , \SB2_3_21/i1[9] , \SB2_3_21/i0_0 ,
         \SB2_3_21/i0_3 , \SB2_3_21/i0[10] , \SB2_3_21/i0[9] ,
         \SB2_3_21/i0[8] , \SB2_3_21/i0[6] , \SB2_3_22/buf_output[5] ,
         \SB2_3_22/buf_output[4] , \SB2_3_22/buf_output[3] ,
         \SB2_3_22/buf_output[2] , \SB2_3_22/buf_output[1] ,
         \SB2_3_22/buf_output[0] , \SB2_3_22/i3[0] , \SB2_3_22/i1_5 ,
         \SB2_3_22/i1_7 , \SB2_3_22/i1[9] , \SB2_3_22/i0_0 , \SB2_3_22/i0_3 ,
         \SB2_3_22/i0[10] , \SB2_3_22/i0[9] , \SB2_3_22/i0[8] ,
         \SB2_3_22/i0[6] , \SB2_3_23/buf_output[5] , \SB2_3_23/buf_output[4] ,
         \SB2_3_23/buf_output[3] , \SB2_3_23/buf_output[2] ,
         \SB2_3_23/buf_output[1] , \SB2_3_23/buf_output[0] , \SB2_3_23/i3[0] ,
         \SB2_3_23/i1_5 , \SB2_3_23/i1_7 , \SB2_3_23/i1[9] , \SB2_3_23/i0_0 ,
         \SB2_3_23/i0_3 , \SB2_3_23/i0_4 , \SB2_3_23/i0[10] , \SB2_3_23/i0[9] ,
         \SB2_3_23/i0[8] , \SB2_3_23/i0[7] , \SB2_3_23/i0[6] ,
         \SB2_3_24/buf_output[5] , \SB2_3_24/buf_output[4] ,
         \SB2_3_24/buf_output[3] , \SB2_3_24/buf_output[2] ,
         \SB2_3_24/buf_output[1] , \SB2_3_24/buf_output[0] , \SB2_3_24/i3[0] ,
         \SB2_3_24/i1_5 , \SB2_3_24/i1_7 , \SB2_3_24/i1[9] , \SB2_3_24/i0_0 ,
         \SB2_3_24/i0_3 , \SB2_3_24/i0_4 , \SB2_3_24/i0[10] , \SB2_3_24/i0[9] ,
         \SB2_3_24/i0[8] , \SB2_3_24/i0[7] , \SB2_3_24/i0[6] ,
         \SB2_3_25/buf_output[5] , \SB2_3_25/buf_output[4] ,
         \SB2_3_25/buf_output[3] , \SB2_3_25/buf_output[2] ,
         \SB2_3_25/buf_output[1] , \SB2_3_25/buf_output[0] , \SB2_3_25/i3[0] ,
         \SB2_3_25/i1_5 , \SB2_3_25/i1_7 , \SB2_3_25/i1[9] , \SB2_3_25/i0_0 ,
         \SB2_3_25/i0_3 , \SB2_3_25/i0_4 , \SB2_3_25/i0[10] , \SB2_3_25/i0[8] ,
         \SB2_3_25/i0[7] , \SB2_3_25/i0[6] , \SB2_3_26/buf_output[5] ,
         \SB2_3_26/buf_output[4] , \SB2_3_26/buf_output[3] ,
         \SB2_3_26/buf_output[2] , \SB2_3_26/buf_output[1] ,
         \SB2_3_26/buf_output[0] , \SB2_3_26/i3[0] , \SB2_3_26/i1_5 ,
         \SB2_3_26/i1_7 , \SB2_3_26/i1[9] , \SB2_3_26/i0_0 , \SB2_3_26/i0_3 ,
         \SB2_3_26/i0_4 , \SB2_3_26/i0[10] , \SB2_3_26/i0[9] ,
         \SB2_3_26/i0[8] , \SB2_3_26/i0[6] , \SB2_3_27/buf_output[5] ,
         \SB2_3_27/buf_output[4] , \SB2_3_27/buf_output[3] ,
         \SB2_3_27/buf_output[2] , \SB2_3_27/buf_output[1] ,
         \SB2_3_27/buf_output[0] , \SB2_3_27/i3[0] , \SB2_3_27/i1_5 ,
         \SB2_3_27/i1_7 , \SB2_3_27/i1[9] , \SB2_3_27/i0_0 , \SB2_3_27/i0_3 ,
         \SB2_3_27/i0_4 , \SB2_3_27/i0[10] , \SB2_3_27/i0[9] ,
         \SB2_3_27/i0[8] , \SB2_3_27/i0[7] , \SB2_3_27/i0[6] ,
         \SB2_3_28/buf_output[5] , \SB2_3_28/buf_output[4] ,
         \SB2_3_28/buf_output[3] , \SB2_3_28/buf_output[2] ,
         \SB2_3_28/buf_output[1] , \SB2_3_28/buf_output[0] , \SB2_3_28/i3[0] ,
         \SB2_3_28/i1_5 , \SB2_3_28/i1_7 , \SB2_3_28/i1[9] , \SB2_3_28/i0_0 ,
         \SB2_3_28/i0_3 , \SB2_3_28/i0[10] , \SB2_3_28/i0[9] ,
         \SB2_3_28/i0[8] , \SB2_3_28/i0[6] , \SB2_3_29/buf_output[5] ,
         \SB2_3_29/buf_output[4] , \SB2_3_29/buf_output[3] ,
         \SB2_3_29/buf_output[2] , \SB2_3_29/buf_output[1] ,
         \SB2_3_29/buf_output[0] , \SB2_3_29/i3[0] , \SB2_3_29/i1_5 ,
         \SB2_3_29/i1_7 , \SB2_3_29/i1[9] , \SB2_3_29/i0_0 , \SB2_3_29/i0_3 ,
         \SB2_3_29/i0_4 , \SB2_3_29/i0[10] , \SB2_3_29/i0[9] ,
         \SB2_3_29/i0[8] , \SB2_3_30/buf_output[5] , \SB2_3_30/buf_output[4] ,
         \SB2_3_30/buf_output[3] , \SB2_3_30/buf_output[2] ,
         \SB2_3_30/buf_output[1] , \SB2_3_30/buf_output[0] , \SB2_3_30/i3[0] ,
         \SB2_3_30/i1_5 , \SB2_3_30/i1_7 , \SB2_3_30/i1[9] , \SB2_3_30/i0_0 ,
         \SB2_3_30/i0_3 , \SB2_3_30/i0_4 , \SB2_3_30/i0[10] , \SB2_3_30/i0[9] ,
         \SB2_3_30/i0[8] , \SB2_3_30/i0[7] , \SB2_3_30/i0[6] ,
         \SB2_3_31/buf_output[5] , \SB2_3_31/buf_output[4] ,
         \SB2_3_31/buf_output[3] , \SB2_3_31/buf_output[2] ,
         \SB2_3_31/buf_output[1] , \SB2_3_31/buf_output[0] , \SB2_3_31/i3[0] ,
         \SB2_3_31/i1_5 , \SB2_3_31/i1_7 , \SB2_3_31/i1[9] , \SB2_3_31/i0_0 ,
         \SB2_3_31/i0_3 , \SB2_3_31/i0_4 , \SB2_3_31/i0[10] , \SB2_3_31/i0[9] ,
         \SB2_3_31/i0[8] , \SB2_3_31/i0[7] , \SB2_3_31/i0[6] ,
         \SB1_4_0/buf_output[5] , \SB1_4_0/buf_output[4] ,
         \SB1_4_0/buf_output[3] , \SB1_4_0/buf_output[2] ,
         \SB1_4_0/buf_output[1] , \SB1_4_0/buf_output[0] , \SB1_4_0/i3[0] ,
         \SB1_4_0/i1_5 , \SB1_4_0/i1_7 , \SB1_4_0/i1[9] , \SB1_4_0/i0_0 ,
         \SB1_4_0/i0_3 , \SB1_4_0/i0_4 , \SB1_4_0/i0[10] , \SB1_4_0/i0[9] ,
         \SB1_4_0/i0[8] , \SB1_4_0/i0[7] , \SB1_4_0/i0[6] ,
         \SB1_4_1/buf_output[5] , \SB1_4_1/buf_output[4] ,
         \SB1_4_1/buf_output[3] , \SB1_4_1/buf_output[2] ,
         \SB1_4_1/buf_output[1] , \SB1_4_1/buf_output[0] , \SB1_4_1/i3[0] ,
         \SB1_4_1/i1_5 , \SB1_4_1/i1_7 , \SB1_4_1/i1[9] , \SB1_4_1/i0_0 ,
         \SB1_4_1/i0_3 , \SB1_4_1/i0_4 , \SB1_4_1/i0[10] , \SB1_4_1/i0[9] ,
         \SB1_4_1/i0[8] , \SB1_4_1/i0[7] , \SB1_4_1/i0[6] ,
         \SB1_4_2/buf_output[5] , \SB1_4_2/buf_output[3] ,
         \SB1_4_2/buf_output[2] , \SB1_4_2/buf_output[1] ,
         \SB1_4_2/buf_output[0] , \SB1_4_2/i3[0] , \SB1_4_2/i1_5 ,
         \SB1_4_2/i1_7 , \SB1_4_2/i1[9] , \SB1_4_2/i0_0 , \SB1_4_2/i0_3 ,
         \SB1_4_2/i0_4 , \SB1_4_2/i0[10] , \SB1_4_2/i0[9] , \SB1_4_2/i0[8] ,
         \SB1_4_2/i0[7] , \SB1_4_2/i0[6] , \SB1_4_3/buf_output[5] ,
         \SB1_4_3/buf_output[4] , \SB1_4_3/buf_output[3] ,
         \SB1_4_3/buf_output[1] , \SB1_4_3/buf_output[0] , \SB1_4_3/i3[0] ,
         \SB1_4_3/i1_5 , \SB1_4_3/i1_7 , \SB1_4_3/i1[9] , \SB1_4_3/i0_0 ,
         \SB1_4_3/i0_3 , \SB1_4_3/i0_4 , \SB1_4_3/i0[10] , \SB1_4_3/i0[9] ,
         \SB1_4_3/i0[8] , \SB1_4_3/i0[7] , \SB1_4_3/i0[6] ,
         \SB1_4_4/buf_output[5] , \SB1_4_4/buf_output[4] ,
         \SB1_4_4/buf_output[3] , \SB1_4_4/buf_output[2] ,
         \SB1_4_4/buf_output[1] , \SB1_4_4/buf_output[0] , \SB1_4_4/i3[0] ,
         \SB1_4_4/i1_5 , \SB1_4_4/i1_7 , \SB1_4_4/i1[9] , \SB1_4_4/i0_0 ,
         \SB1_4_4/i0_3 , \SB1_4_4/i0_4 , \SB1_4_4/i0[10] , \SB1_4_4/i0[9] ,
         \SB1_4_4/i0[8] , \SB1_4_4/i0[7] , \SB1_4_4/i0[6] ,
         \SB1_4_5/buf_output[5] , \SB1_4_5/buf_output[4] ,
         \SB1_4_5/buf_output[3] , \SB1_4_5/buf_output[2] ,
         \SB1_4_5/buf_output[1] , \SB1_4_5/buf_output[0] , \SB1_4_5/i3[0] ,
         \SB1_4_5/i1_5 , \SB1_4_5/i1_7 , \SB1_4_5/i1[9] , \SB1_4_5/i0_0 ,
         \SB1_4_5/i0_3 , \SB1_4_5/i0_4 , \SB1_4_5/i0[10] , \SB1_4_5/i0[9] ,
         \SB1_4_5/i0[8] , \SB1_4_5/i0[7] , \SB1_4_5/i0[6] ,
         \SB1_4_6/buf_output[5] , \SB1_4_6/buf_output[4] ,
         \SB1_4_6/buf_output[3] , \SB1_4_6/buf_output[2] ,
         \SB1_4_6/buf_output[1] , \SB1_4_6/buf_output[0] , \SB1_4_6/i3[0] ,
         \SB1_4_6/i1_5 , \SB1_4_6/i1_7 , \SB1_4_6/i1[9] , \SB1_4_6/i0_0 ,
         \SB1_4_6/i0_4 , \SB1_4_6/i0[10] , \SB1_4_6/i0[9] , \SB1_4_6/i0[8] ,
         \SB1_4_6/i0[7] , \SB1_4_6/i0[6] , \SB1_4_7/buf_output[5] ,
         \SB1_4_7/buf_output[4] , \SB1_4_7/buf_output[3] ,
         \SB1_4_7/buf_output[2] , \SB1_4_7/buf_output[1] ,
         \SB1_4_7/buf_output[0] , \SB1_4_7/i3[0] , \SB1_4_7/i1_5 ,
         \SB1_4_7/i1_7 , \SB1_4_7/i1[9] , \SB1_4_7/i0_0 , \SB1_4_7/i0_3 ,
         \SB1_4_7/i0_4 , \SB1_4_7/i0[10] , \SB1_4_7/i0[9] , \SB1_4_7/i0[8] ,
         \SB1_4_7/i0[7] , \SB1_4_7/i0[6] , \SB1_4_8/buf_output[5] ,
         \SB1_4_8/buf_output[4] , \SB1_4_8/buf_output[3] ,
         \SB1_4_8/buf_output[2] , \SB1_4_8/buf_output[1] ,
         \SB1_4_8/buf_output[0] , \SB1_4_8/i3[0] , \SB1_4_8/i1_5 ,
         \SB1_4_8/i1_7 , \SB1_4_8/i1[9] , \SB1_4_8/i0_0 , \SB1_4_8/i0_3 ,
         \SB1_4_8/i0_4 , \SB1_4_8/i0[10] , \SB1_4_8/i0[9] , \SB1_4_8/i0[8] ,
         \SB1_4_8/i0[7] , \SB1_4_8/i0[6] , \SB1_4_9/buf_output[5] ,
         \SB1_4_9/buf_output[3] , \SB1_4_9/buf_output[2] ,
         \SB1_4_9/buf_output[1] , \SB1_4_9/buf_output[0] , \SB1_4_9/i3[0] ,
         \SB1_4_9/i1_5 , \SB1_4_9/i1_7 , \SB1_4_9/i1[9] , \SB1_4_9/i0_0 ,
         \SB1_4_9/i0_3 , \SB1_4_9/i0_4 , \SB1_4_9/i0[10] , \SB1_4_9/i0[9] ,
         \SB1_4_9/i0[8] , \SB1_4_9/i0[7] , \SB1_4_9/i0[6] ,
         \SB1_4_10/buf_output[5] , \SB1_4_10/buf_output[4] ,
         \SB1_4_10/buf_output[3] , \SB1_4_10/buf_output[2] ,
         \SB1_4_10/buf_output[1] , \SB1_4_10/buf_output[0] , \SB1_4_10/i3[0] ,
         \SB1_4_10/i1_5 , \SB1_4_10/i1_7 , \SB1_4_10/i1[9] , \SB1_4_10/i0_0 ,
         \SB1_4_10/i0_4 , \SB1_4_10/i0[10] , \SB1_4_10/i0[9] ,
         \SB1_4_10/i0[8] , \SB1_4_10/i0[7] , \SB1_4_10/i0[6] ,
         \SB1_4_11/buf_output[5] , \SB1_4_11/buf_output[4] ,
         \SB1_4_11/buf_output[3] , \SB1_4_11/buf_output[2] ,
         \SB1_4_11/buf_output[1] , \SB1_4_11/buf_output[0] , \SB1_4_11/i3[0] ,
         \SB1_4_11/i1_5 , \SB1_4_11/i1_7 , \SB1_4_11/i1[9] , \SB1_4_11/i0_0 ,
         \SB1_4_11/i0_3 , \SB1_4_11/i0_4 , \SB1_4_11/i0[10] , \SB1_4_11/i0[9] ,
         \SB1_4_11/i0[8] , \SB1_4_11/i0[7] , \SB1_4_11/i0[6] ,
         \SB1_4_12/buf_output[5] , \SB1_4_12/buf_output[4] ,
         \SB1_4_12/buf_output[3] , \SB1_4_12/buf_output[2] ,
         \SB1_4_12/buf_output[1] , \SB1_4_12/buf_output[0] , \SB1_4_12/i3[0] ,
         \SB1_4_12/i1_5 , \SB1_4_12/i1_7 , \SB1_4_12/i1[9] , \SB1_4_12/i0_0 ,
         \SB1_4_12/i0_4 , \SB1_4_12/i0[10] , \SB1_4_12/i0[9] ,
         \SB1_4_12/i0[8] , \SB1_4_12/i0[7] , \SB1_4_12/i0[6] ,
         \SB1_4_13/buf_output[5] , \SB1_4_13/buf_output[4] ,
         \SB1_4_13/buf_output[3] , \SB1_4_13/buf_output[2] ,
         \SB1_4_13/buf_output[1] , \SB1_4_13/buf_output[0] , \SB1_4_13/i3[0] ,
         \SB1_4_13/i1_5 , \SB1_4_13/i1_7 , \SB1_4_13/i1[9] , \SB1_4_13/i0_0 ,
         \SB1_4_13/i0_3 , \SB1_4_13/i0_4 , \SB1_4_13/i0[10] , \SB1_4_13/i0[9] ,
         \SB1_4_13/i0[8] , \SB1_4_13/i0[7] , \SB1_4_13/i0[6] ,
         \SB1_4_14/buf_output[5] , \SB1_4_14/buf_output[4] ,
         \SB1_4_14/buf_output[3] , \SB1_4_14/buf_output[2] ,
         \SB1_4_14/buf_output[0] , \SB1_4_14/i3[0] , \SB1_4_14/i1_5 ,
         \SB1_4_14/i1_7 , \SB1_4_14/i1[9] , \SB1_4_14/i0_0 , \SB1_4_14/i0_3 ,
         \SB1_4_14/i0_4 , \SB1_4_14/i0[10] , \SB1_4_14/i0[9] ,
         \SB1_4_14/i0[8] , \SB1_4_14/i0[7] , \SB1_4_14/i0[6] ,
         \SB1_4_15/buf_output[5] , \SB1_4_15/buf_output[4] ,
         \SB1_4_15/buf_output[3] , \SB1_4_15/buf_output[2] ,
         \SB1_4_15/buf_output[1] , \SB1_4_15/buf_output[0] , \SB1_4_15/i3[0] ,
         \SB1_4_15/i1_5 , \SB1_4_15/i1_7 , \SB1_4_15/i1[9] , \SB1_4_15/i0_0 ,
         \SB1_4_15/i0_3 , \SB1_4_15/i0_4 , \SB1_4_15/i0[10] , \SB1_4_15/i0[9] ,
         \SB1_4_15/i0[8] , \SB1_4_15/i0[7] , \SB1_4_15/i0[6] ,
         \SB1_4_16/buf_output[5] , \SB1_4_16/buf_output[4] ,
         \SB1_4_16/buf_output[3] , \SB1_4_16/buf_output[2] ,
         \SB1_4_16/buf_output[1] , \SB1_4_16/buf_output[0] , \SB1_4_16/i3[0] ,
         \SB1_4_16/i1_5 , \SB1_4_16/i1_7 , \SB1_4_16/i1[9] , \SB1_4_16/i0_0 ,
         \SB1_4_16/i0_3 , \SB1_4_16/i0_4 , \SB1_4_16/i0[10] , \SB1_4_16/i0[9] ,
         \SB1_4_16/i0[8] , \SB1_4_16/i0[7] , \SB1_4_16/i0[6] ,
         \SB1_4_17/buf_output[5] , \SB1_4_17/buf_output[4] ,
         \SB1_4_17/buf_output[3] , \SB1_4_17/buf_output[2] ,
         \SB1_4_17/buf_output[1] , \SB1_4_17/buf_output[0] , \SB1_4_17/i3[0] ,
         \SB1_4_17/i1_5 , \SB1_4_17/i1_7 , \SB1_4_17/i1[9] , \SB1_4_17/i0_0 ,
         \SB1_4_17/i0_3 , \SB1_4_17/i0_4 , \SB1_4_17/i0[10] , \SB1_4_17/i0[9] ,
         \SB1_4_17/i0[8] , \SB1_4_17/i0[7] , \SB1_4_17/i0[6] ,
         \SB1_4_18/buf_output[5] , \SB1_4_18/buf_output[4] ,
         \SB1_4_18/buf_output[3] , \SB1_4_18/buf_output[2] ,
         \SB1_4_18/buf_output[1] , \SB1_4_18/buf_output[0] , \SB1_4_18/i3[0] ,
         \SB1_4_18/i1_5 , \SB1_4_18/i1_7 , \SB1_4_18/i1[9] , \SB1_4_18/i0_0 ,
         \SB1_4_18/i0_3 , \SB1_4_18/i0_4 , \SB1_4_18/i0[10] , \SB1_4_18/i0[9] ,
         \SB1_4_18/i0[8] , \SB1_4_18/i0[7] , \SB1_4_18/i0[6] ,
         \SB1_4_19/buf_output[5] , \SB1_4_19/buf_output[4] ,
         \SB1_4_19/buf_output[3] , \SB1_4_19/buf_output[2] ,
         \SB1_4_19/buf_output[1] , \SB1_4_19/buf_output[0] , \SB1_4_19/i3[0] ,
         \SB1_4_19/i1_5 , \SB1_4_19/i1_7 , \SB1_4_19/i1[9] , \SB1_4_19/i0_0 ,
         \SB1_4_19/i0_3 , \SB1_4_19/i0_4 , \SB1_4_19/i0[10] , \SB1_4_19/i0[9] ,
         \SB1_4_19/i0[8] , \SB1_4_19/i0[7] , \SB1_4_19/i0[6] ,
         \SB1_4_20/buf_output[5] , \SB1_4_20/buf_output[4] ,
         \SB1_4_20/buf_output[3] , \SB1_4_20/buf_output[2] ,
         \SB1_4_20/buf_output[1] , \SB1_4_20/buf_output[0] , \SB1_4_20/i3[0] ,
         \SB1_4_20/i1_5 , \SB1_4_20/i1_7 , \SB1_4_20/i1[9] , \SB1_4_20/i0_0 ,
         \SB1_4_20/i0_3 , \SB1_4_20/i0_4 , \SB1_4_20/i0[10] , \SB1_4_20/i0[9] ,
         \SB1_4_20/i0[8] , \SB1_4_20/i0[7] , \SB1_4_20/i0[6] ,
         \SB1_4_21/buf_output[5] , \SB1_4_21/buf_output[3] ,
         \SB1_4_21/buf_output[2] , \SB1_4_21/buf_output[1] ,
         \SB1_4_21/buf_output[0] , \SB1_4_21/i3[0] , \SB1_4_21/i1_5 ,
         \SB1_4_21/i1_7 , \SB1_4_21/i1[9] , \SB1_4_21/i0_0 , \SB1_4_21/i0_3 ,
         \SB1_4_21/i0_4 , \SB1_4_21/i0[10] , \SB1_4_21/i0[9] ,
         \SB1_4_21/i0[8] , \SB1_4_21/i0[7] , \SB1_4_21/i0[6] ,
         \SB1_4_22/buf_output[5] , \SB1_4_22/buf_output[4] ,
         \SB1_4_22/buf_output[3] , \SB1_4_22/buf_output[2] ,
         \SB1_4_22/buf_output[1] , \SB1_4_22/buf_output[0] , \SB1_4_22/i3[0] ,
         \SB1_4_22/i1_5 , \SB1_4_22/i1_7 , \SB1_4_22/i1[9] , \SB1_4_22/i0_0 ,
         \SB1_4_22/i0_4 , \SB1_4_22/i0[10] , \SB1_4_22/i0[9] ,
         \SB1_4_22/i0[8] , \SB1_4_22/i0[7] , \SB1_4_22/i0[6] ,
         \SB1_4_23/buf_output[5] , \SB1_4_23/buf_output[4] ,
         \SB1_4_23/buf_output[3] , \SB1_4_23/buf_output[2] ,
         \SB1_4_23/buf_output[1] , \SB1_4_23/buf_output[0] , \SB1_4_23/i3[0] ,
         \SB1_4_23/i1_5 , \SB1_4_23/i1_7 , \SB1_4_23/i1[9] , \SB1_4_23/i0_0 ,
         \SB1_4_23/i0_3 , \SB1_4_23/i0_4 , \SB1_4_23/i0[10] , \SB1_4_23/i0[9] ,
         \SB1_4_23/i0[8] , \SB1_4_23/i0[7] , \SB1_4_23/i0[6] ,
         \SB1_4_24/buf_output[5] , \SB1_4_24/buf_output[4] ,
         \SB1_4_24/buf_output[3] , \SB1_4_24/buf_output[2] ,
         \SB1_4_24/buf_output[1] , \SB1_4_24/buf_output[0] , \SB1_4_24/i3[0] ,
         \SB1_4_24/i1_5 , \SB1_4_24/i1_7 , \SB1_4_24/i1[9] , \SB1_4_24/i0_0 ,
         \SB1_4_24/i0_3 , \SB1_4_24/i0_4 , \SB1_4_24/i0[10] , \SB1_4_24/i0[9] ,
         \SB1_4_24/i0[8] , \SB1_4_24/i0[7] , \SB1_4_24/i0[6] ,
         \SB1_4_25/buf_output[5] , \SB1_4_25/buf_output[4] ,
         \SB1_4_25/buf_output[3] , \SB1_4_25/buf_output[2] ,
         \SB1_4_25/buf_output[1] , \SB1_4_25/buf_output[0] , \SB1_4_25/i3[0] ,
         \SB1_4_25/i1_5 , \SB1_4_25/i1_7 , \SB1_4_25/i1[9] , \SB1_4_25/i0_0 ,
         \SB1_4_25/i0_3 , \SB1_4_25/i0_4 , \SB1_4_25/i0[10] , \SB1_4_25/i0[9] ,
         \SB1_4_25/i0[8] , \SB1_4_25/i0[7] , \SB1_4_25/i0[6] ,
         \SB1_4_26/buf_output[5] , \SB1_4_26/buf_output[4] ,
         \SB1_4_26/buf_output[3] , \SB1_4_26/buf_output[2] ,
         \SB1_4_26/buf_output[1] , \SB1_4_26/buf_output[0] , \SB1_4_26/i3[0] ,
         \SB1_4_26/i1_5 , \SB1_4_26/i1_7 , \SB1_4_26/i1[9] , \SB1_4_26/i0_0 ,
         \SB1_4_26/i0_3 , \SB1_4_26/i0_4 , \SB1_4_26/i0[10] , \SB1_4_26/i0[9] ,
         \SB1_4_26/i0[8] , \SB1_4_26/i0[7] , \SB1_4_26/i0[6] ,
         \SB1_4_27/buf_output[5] , \SB1_4_27/buf_output[4] ,
         \SB1_4_27/buf_output[3] , \SB1_4_27/buf_output[2] ,
         \SB1_4_27/buf_output[1] , \SB1_4_27/buf_output[0] , \SB1_4_27/i3[0] ,
         \SB1_4_27/i1_5 , \SB1_4_27/i1_7 , \SB1_4_27/i1[9] , \SB1_4_27/i0_3 ,
         \SB1_4_27/i0_4 , \SB1_4_27/i0[10] , \SB1_4_27/i0[9] ,
         \SB1_4_27/i0[8] , \SB1_4_27/i0[7] , \SB1_4_27/i0[6] ,
         \SB1_4_28/buf_output[5] , \SB1_4_28/buf_output[4] ,
         \SB1_4_28/buf_output[3] , \SB1_4_28/buf_output[2] ,
         \SB1_4_28/buf_output[1] , \SB1_4_28/buf_output[0] , \SB1_4_28/i3[0] ,
         \SB1_4_28/i1_5 , \SB1_4_28/i1_7 , \SB1_4_28/i1[9] , \SB1_4_28/i0_0 ,
         \SB1_4_28/i0_3 , \SB1_4_28/i0_4 , \SB1_4_28/i0[10] , \SB1_4_28/i0[9] ,
         \SB1_4_28/i0[8] , \SB1_4_28/i0[7] , \SB1_4_28/i0[6] ,
         \SB1_4_29/buf_output[5] , \SB1_4_29/buf_output[4] ,
         \SB1_4_29/buf_output[3] , \SB1_4_29/buf_output[2] ,
         \SB1_4_29/buf_output[1] , \SB1_4_29/buf_output[0] , \SB1_4_29/i3[0] ,
         \SB1_4_29/i1_5 , \SB1_4_29/i1_7 , \SB1_4_29/i1[9] , \SB1_4_29/i0_0 ,
         \SB1_4_29/i0_4 , \SB1_4_29/i0[10] , \SB1_4_29/i0[9] ,
         \SB1_4_29/i0[8] , \SB1_4_29/i0[7] , \SB1_4_29/i0[6] ,
         \SB1_4_30/buf_output[5] , \SB1_4_30/buf_output[4] ,
         \SB1_4_30/buf_output[3] , \SB1_4_30/buf_output[2] ,
         \SB1_4_30/buf_output[1] , \SB1_4_30/buf_output[0] , \SB1_4_30/i3[0] ,
         \SB1_4_30/i1_5 , \SB1_4_30/i1_7 , \SB1_4_30/i1[9] , \SB1_4_30/i0_0 ,
         \SB1_4_30/i0_3 , \SB1_4_30/i0_4 , \SB1_4_30/i0[10] , \SB1_4_30/i0[9] ,
         \SB1_4_30/i0[8] , \SB1_4_30/i0[7] , \SB1_4_30/i0[6] ,
         \SB1_4_31/buf_output[5] , \SB1_4_31/buf_output[4] ,
         \SB1_4_31/buf_output[3] , \SB1_4_31/buf_output[2] ,
         \SB1_4_31/buf_output[1] , \SB1_4_31/buf_output[0] , \SB1_4_31/i3[0] ,
         \SB1_4_31/i1_5 , \SB1_4_31/i1_7 , \SB1_4_31/i1[9] , \SB1_4_31/i0_0 ,
         \SB1_4_31/i0_3 , \SB1_4_31/i0_4 , \SB1_4_31/i0[10] , \SB1_4_31/i0[9] ,
         \SB1_4_31/i0[8] , \SB1_4_31/i0[7] , \SB1_4_31/i0[6] ,
         \SB2_4_0/buf_output[5] , \SB2_4_0/buf_output[4] ,
         \SB2_4_0/buf_output[3] , \SB2_4_0/buf_output[2] ,
         \SB2_4_0/buf_output[1] , \SB2_4_0/buf_output[0] , \SB2_4_0/i3[0] ,
         \SB2_4_0/i1_7 , \SB2_4_0/i1[9] , \SB2_4_0/i0_0 , \SB2_4_0/i0_3 ,
         \SB2_4_0/i0_4 , \SB2_4_0/i0[10] , \SB2_4_0/i0[9] , \SB2_4_0/i0[8] ,
         \SB2_4_0/i0[7] , \SB2_4_0/i0[6] , \SB2_4_1/buf_output[5] ,
         \SB2_4_1/buf_output[4] , \SB2_4_1/buf_output[3] ,
         \SB2_4_1/buf_output[2] , \SB2_4_1/buf_output[1] ,
         \SB2_4_1/buf_output[0] , \SB2_4_1/i3[0] , \SB2_4_1/i1_7 ,
         \SB2_4_1/i1[9] , \SB2_4_1/i0_0 , \SB2_4_1/i0_3 , \SB2_4_1/i0_4 ,
         \SB2_4_1/i0[10] , \SB2_4_1/i0[9] , \SB2_4_1/i0[8] , \SB2_4_1/i0[6] ,
         \SB2_4_2/buf_output[5] , \SB2_4_2/buf_output[4] ,
         \SB2_4_2/buf_output[3] , \SB2_4_2/buf_output[2] ,
         \SB2_4_2/buf_output[1] , \SB2_4_2/buf_output[0] , \SB2_4_2/i3[0] ,
         \SB2_4_2/i1_5 , \SB2_4_2/i1_7 , \SB2_4_2/i1[9] , \SB2_4_2/i0_0 ,
         \SB2_4_2/i0_3 , \SB2_4_2/i0_4 , \SB2_4_2/i0[10] , \SB2_4_2/i0[9] ,
         \SB2_4_2/i0[8] , \SB2_4_2/i0[7] , \SB2_4_2/i0[6] ,
         \SB2_4_3/buf_output[5] , \SB2_4_3/buf_output[4] ,
         \SB2_4_3/buf_output[3] , \SB2_4_3/buf_output[2] ,
         \SB2_4_3/buf_output[1] , \SB2_4_3/buf_output[0] , \SB2_4_3/i3[0] ,
         \SB2_4_3/i1_7 , \SB2_4_3/i1[9] , \SB2_4_3/i0_0 , \SB2_4_3/i0_3 ,
         \SB2_4_3/i0_4 , \SB2_4_3/i0[10] , \SB2_4_3/i0[9] , \SB2_4_3/i0[8] ,
         \SB2_4_3/i0[7] , \SB2_4_3/i0[6] , \SB2_4_4/buf_output[5] ,
         \SB2_4_4/buf_output[4] , \SB2_4_4/buf_output[3] ,
         \SB2_4_4/buf_output[2] , \SB2_4_4/buf_output[1] ,
         \SB2_4_4/buf_output[0] , \SB2_4_4/i3[0] , \SB2_4_4/i1_5 ,
         \SB2_4_4/i1_7 , \SB2_4_4/i1[9] , \SB2_4_4/i0_0 , \SB2_4_4/i0_3 ,
         \SB2_4_4/i0_4 , \SB2_4_4/i0[10] , \SB2_4_4/i0[9] , \SB2_4_4/i0[8] ,
         \SB2_4_4/i0[7] , \SB2_4_4/i0[6] , \SB2_4_5/buf_output[5] ,
         \SB2_4_5/buf_output[4] , \SB2_4_5/buf_output[3] ,
         \SB2_4_5/buf_output[2] , \SB2_4_5/buf_output[1] ,
         \SB2_4_5/buf_output[0] , \SB2_4_5/i3[0] , \SB2_4_5/i1_5 ,
         \SB2_4_5/i1_7 , \SB2_4_5/i1[9] , \SB2_4_5/i0_0 , \SB2_4_5/i0_3 ,
         \SB2_4_5/i0[10] , \SB2_4_5/i0[9] , \SB2_4_5/i0[8] , \SB2_4_5/i0[7] ,
         \SB2_4_5/i0[6] , \SB2_4_6/buf_output[5] , \SB2_4_6/buf_output[4] ,
         \SB2_4_6/buf_output[3] , \SB2_4_6/buf_output[2] ,
         \SB2_4_6/buf_output[0] , \SB2_4_6/i3[0] , \SB2_4_6/i1_5 ,
         \SB2_4_6/i1_7 , \SB2_4_6/i1[9] , \SB2_4_6/i0_0 , \SB2_4_6/i0_3 ,
         \SB2_4_6/i0_4 , \SB2_4_6/i0[10] , \SB2_4_6/i0[9] , \SB2_4_6/i0[8] ,
         \SB2_4_6/i0[7] , \SB2_4_6/i0[6] , \SB2_4_7/buf_output[5] ,
         \SB2_4_7/buf_output[4] , \SB2_4_7/buf_output[3] ,
         \SB2_4_7/buf_output[2] , \SB2_4_7/buf_output[1] ,
         \SB2_4_7/buf_output[0] , \SB2_4_7/i3[0] , \SB2_4_7/i1_5 ,
         \SB2_4_7/i1_7 , \SB2_4_7/i1[9] , \SB2_4_7/i0_0 , \SB2_4_7/i0_3 ,
         \SB2_4_7/i0[10] , \SB2_4_7/i0[9] , \SB2_4_7/i0[8] , \SB2_4_7/i0[7] ,
         \SB2_4_7/i0[6] , \SB2_4_8/buf_output[5] , \SB2_4_8/buf_output[4] ,
         \SB2_4_8/buf_output[3] , \SB2_4_8/buf_output[2] ,
         \SB2_4_8/buf_output[1] , \SB2_4_8/buf_output[0] , \SB2_4_8/i3[0] ,
         \SB2_4_8/i1_5 , \SB2_4_8/i1_7 , \SB2_4_8/i1[9] , \SB2_4_8/i0_0 ,
         \SB2_4_8/i0_3 , \SB2_4_8/i0[10] , \SB2_4_8/i0[9] , \SB2_4_8/i0[8] ,
         \SB2_4_8/i0[7] , \SB2_4_8/i0[6] , \SB2_4_9/buf_output[5] ,
         \SB2_4_9/buf_output[4] , \SB2_4_9/buf_output[3] ,
         \SB2_4_9/buf_output[2] , \SB2_4_9/buf_output[1] ,
         \SB2_4_9/buf_output[0] , \SB2_4_9/i3[0] , \SB2_4_9/i1_5 ,
         \SB2_4_9/i1_7 , \SB2_4_9/i1[9] , \SB2_4_9/i0_0 , \SB2_4_9/i0_3 ,
         \SB2_4_9/i0_4 , \SB2_4_9/i0[10] , \SB2_4_9/i0[9] , \SB2_4_9/i0[8] ,
         \SB2_4_9/i0[7] , \SB2_4_9/i0[6] , \SB2_4_10/buf_output[5] ,
         \SB2_4_10/buf_output[4] , \SB2_4_10/buf_output[3] ,
         \SB2_4_10/buf_output[2] , \SB2_4_10/buf_output[1] ,
         \SB2_4_10/buf_output[0] , \SB2_4_10/i3[0] , \SB2_4_10/i1_7 ,
         \SB2_4_10/i1[9] , \SB2_4_10/i0_0 , \SB2_4_10/i0_3 , \SB2_4_10/i0_4 ,
         \SB2_4_10/i0[10] , \SB2_4_10/i0[9] , \SB2_4_10/i0[8] ,
         \SB2_4_10/i0[7] , \SB2_4_10/i0[6] , \SB2_4_11/buf_output[5] ,
         \SB2_4_11/buf_output[4] , \SB2_4_11/buf_output[3] ,
         \SB2_4_11/buf_output[2] , \SB2_4_11/buf_output[1] ,
         \SB2_4_11/buf_output[0] , \SB2_4_11/i3[0] , \SB2_4_11/i1_5 ,
         \SB2_4_11/i1_7 , \SB2_4_11/i1[9] , \SB2_4_11/i0_0 , \SB2_4_11/i0_3 ,
         \SB2_4_11/i0_4 , \SB2_4_11/i0[10] , \SB2_4_11/i0[9] ,
         \SB2_4_11/i0[8] , \SB2_4_11/i0[7] , \SB2_4_11/i0[6] ,
         \SB2_4_12/buf_output[5] , \SB2_4_12/buf_output[4] ,
         \SB2_4_12/buf_output[3] , \SB2_4_12/buf_output[2] ,
         \SB2_4_12/buf_output[1] , \SB2_4_12/buf_output[0] , \SB2_4_12/i3[0] ,
         \SB2_4_12/i1_5 , \SB2_4_12/i1_7 , \SB2_4_12/i1[9] , \SB2_4_12/i0_0 ,
         \SB2_4_12/i0_3 , \SB2_4_12/i0_4 , \SB2_4_12/i0[10] , \SB2_4_12/i0[9] ,
         \SB2_4_12/i0[8] , \SB2_4_12/i0[7] , \SB2_4_12/i0[6] ,
         \SB2_4_13/buf_output[5] , \SB2_4_13/buf_output[4] ,
         \SB2_4_13/buf_output[3] , \SB2_4_13/buf_output[2] ,
         \SB2_4_13/buf_output[1] , \SB2_4_13/buf_output[0] , \SB2_4_13/i3[0] ,
         \SB2_4_13/i1_5 , \SB2_4_13/i1_7 , \SB2_4_13/i1[9] , \SB2_4_13/i0_0 ,
         \SB2_4_13/i0_3 , \SB2_4_13/i0_4 , \SB2_4_13/i0[10] , \SB2_4_13/i0[9] ,
         \SB2_4_13/i0[8] , \SB2_4_13/i0[7] , \SB2_4_13/i0[6] ,
         \SB2_4_14/buf_output[5] , \SB2_4_14/buf_output[4] ,
         \SB2_4_14/buf_output[3] , \SB2_4_14/buf_output[2] ,
         \SB2_4_14/buf_output[1] , \SB2_4_14/buf_output[0] , \SB2_4_14/i3[0] ,
         \SB2_4_14/i1_5 , \SB2_4_14/i1_7 , \SB2_4_14/i1[9] , \SB2_4_14/i0_0 ,
         \SB2_4_14/i0_3 , \SB2_4_14/i0_4 , \SB2_4_14/i0[10] , \SB2_4_14/i0[9] ,
         \SB2_4_14/i0[8] , \SB2_4_14/i0[7] , \SB2_4_14/i0[6] ,
         \SB2_4_15/buf_output[5] , \SB2_4_15/buf_output[4] ,
         \SB2_4_15/buf_output[3] , \SB2_4_15/buf_output[1] ,
         \SB2_4_15/buf_output[0] , \SB2_4_15/i3[0] , \SB2_4_15/i1_5 ,
         \SB2_4_15/i1_7 , \SB2_4_15/i1[9] , \SB2_4_15/i0_0 , \SB2_4_15/i0_3 ,
         \SB2_4_15/i0_4 , \SB2_4_15/i0[10] , \SB2_4_15/i0[9] ,
         \SB2_4_15/i0[8] , \SB2_4_15/i0[7] , \SB2_4_15/i0[6] ,
         \SB2_4_16/buf_output[5] , \SB2_4_16/buf_output[4] ,
         \SB2_4_16/buf_output[3] , \SB2_4_16/buf_output[2] ,
         \SB2_4_16/buf_output[1] , \SB2_4_16/buf_output[0] , \SB2_4_16/i3[0] ,
         \SB2_4_16/i1_5 , \SB2_4_16/i1_7 , \SB2_4_16/i1[9] , \SB2_4_16/i0_0 ,
         \SB2_4_16/i0_3 , \SB2_4_16/i0_4 , \SB2_4_16/i0[10] , \SB2_4_16/i0[9] ,
         \SB2_4_16/i0[8] , \SB2_4_16/i0[7] , \SB2_4_16/i0[6] ,
         \SB2_4_17/buf_output[5] , \SB2_4_17/buf_output[4] ,
         \SB2_4_17/buf_output[3] , \SB2_4_17/buf_output[2] ,
         \SB2_4_17/buf_output[0] , \SB2_4_17/i3[0] , \SB2_4_17/i1_5 ,
         \SB2_4_17/i1_7 , \SB2_4_17/i1[9] , \SB2_4_17/i0_0 , \SB2_4_17/i0_3 ,
         \SB2_4_17/i0_4 , \SB2_4_17/i0[10] , \SB2_4_17/i0[9] ,
         \SB2_4_17/i0[8] , \SB2_4_17/i0[7] , \SB2_4_17/i0[6] ,
         \SB2_4_18/buf_output[5] , \SB2_4_18/buf_output[4] ,
         \SB2_4_18/buf_output[3] , \SB2_4_18/buf_output[2] ,
         \SB2_4_18/buf_output[1] , \SB2_4_18/buf_output[0] , \SB2_4_18/i3[0] ,
         \SB2_4_18/i1_5 , \SB2_4_18/i1_7 , \SB2_4_18/i1[9] , \SB2_4_18/i0_0 ,
         \SB2_4_18/i0_3 , \SB2_4_18/i0_4 , \SB2_4_18/i0[10] , \SB2_4_18/i0[9] ,
         \SB2_4_18/i0[8] , \SB2_4_18/i0[7] , \SB2_4_18/i0[6] ,
         \SB2_4_19/buf_output[5] , \SB2_4_19/buf_output[4] ,
         \SB2_4_19/buf_output[3] , \SB2_4_19/buf_output[2] ,
         \SB2_4_19/buf_output[1] , \SB2_4_19/buf_output[0] , \SB2_4_19/i3[0] ,
         \SB2_4_19/i1_5 , \SB2_4_19/i1_7 , \SB2_4_19/i1[9] , \SB2_4_19/i0_0 ,
         \SB2_4_19/i0_3 , \SB2_4_19/i0_4 , \SB2_4_19/i0[10] , \SB2_4_19/i0[9] ,
         \SB2_4_19/i0[8] , \SB2_4_19/i0[7] , \SB2_4_19/i0[6] ,
         \SB2_4_20/buf_output[5] , \SB2_4_20/buf_output[4] ,
         \SB2_4_20/buf_output[3] , \SB2_4_20/buf_output[2] ,
         \SB2_4_20/buf_output[1] , \SB2_4_20/buf_output[0] , \SB2_4_20/i3[0] ,
         \SB2_4_20/i1_5 , \SB2_4_20/i1_7 , \SB2_4_20/i1[9] , \SB2_4_20/i0_0 ,
         \SB2_4_20/i0_3 , \SB2_4_20/i0_4 , \SB2_4_20/i0[10] , \SB2_4_20/i0[9] ,
         \SB2_4_20/i0[8] , \SB2_4_20/i0[7] , \SB2_4_20/i0[6] ,
         \SB2_4_21/buf_output[5] , \SB2_4_21/buf_output[4] ,
         \SB2_4_21/buf_output[3] , \SB2_4_21/buf_output[2] ,
         \SB2_4_21/buf_output[1] , \SB2_4_21/buf_output[0] , \SB2_4_21/i3[0] ,
         \SB2_4_21/i1_5 , \SB2_4_21/i1_7 , \SB2_4_21/i1[9] , \SB2_4_21/i0_0 ,
         \SB2_4_21/i0_3 , \SB2_4_21/i0_4 , \SB2_4_21/i0[10] , \SB2_4_21/i0[9] ,
         \SB2_4_21/i0[8] , \SB2_4_21/i0[7] , \SB2_4_21/i0[6] ,
         \SB2_4_22/buf_output[5] , \SB2_4_22/buf_output[4] ,
         \SB2_4_22/buf_output[3] , \SB2_4_22/buf_output[2] ,
         \SB2_4_22/buf_output[1] , \SB2_4_22/buf_output[0] , \SB2_4_22/i3[0] ,
         \SB2_4_22/i1_5 , \SB2_4_22/i1_7 , \SB2_4_22/i1[9] , \SB2_4_22/i0_0 ,
         \SB2_4_22/i0_3 , \SB2_4_22/i0_4 , \SB2_4_22/i0[10] , \SB2_4_22/i0[9] ,
         \SB2_4_22/i0[8] , \SB2_4_22/i0[7] , \SB2_4_22/i0[6] ,
         \SB2_4_23/buf_output[5] , \SB2_4_23/buf_output[4] ,
         \SB2_4_23/buf_output[3] , \SB2_4_23/buf_output[2] ,
         \SB2_4_23/buf_output[1] , \SB2_4_23/buf_output[0] , \SB2_4_23/i3[0] ,
         \SB2_4_23/i1_5 , \SB2_4_23/i1_7 , \SB2_4_23/i1[9] , \SB2_4_23/i0_0 ,
         \SB2_4_23/i0_3 , \SB2_4_23/i0_4 , \SB2_4_23/i0[10] , \SB2_4_23/i0[9] ,
         \SB2_4_23/i0[8] , \SB2_4_23/i0[7] , \SB2_4_23/i0[6] ,
         \SB2_4_24/buf_output[5] , \SB2_4_24/buf_output[4] ,
         \SB2_4_24/buf_output[3] , \SB2_4_24/buf_output[2] ,
         \SB2_4_24/buf_output[1] , \SB2_4_24/buf_output[0] , \SB2_4_24/i3[0] ,
         \SB2_4_24/i1_7 , \SB2_4_24/i0_0 , \SB2_4_24/i0_3 , \SB2_4_24/i0_4 ,
         \SB2_4_24/i0[10] , \SB2_4_24/i0[9] , \SB2_4_24/i0[8] ,
         \SB2_4_24/i0[7] , \SB2_4_24/i0[6] , \SB2_4_25/buf_output[5] ,
         \SB2_4_25/buf_output[4] , \SB2_4_25/buf_output[3] ,
         \SB2_4_25/buf_output[2] , \SB2_4_25/buf_output[1] ,
         \SB2_4_25/buf_output[0] , \SB2_4_25/i3[0] , \SB2_4_25/i1_5 ,
         \SB2_4_25/i1_7 , \SB2_4_25/i1[9] , \SB2_4_25/i0_0 , \SB2_4_25/i0_3 ,
         \SB2_4_25/i0_4 , \SB2_4_25/i0[10] , \SB2_4_25/i0[9] ,
         \SB2_4_25/i0[8] , \SB2_4_25/i0[7] , \SB2_4_25/i0[6] ,
         \SB2_4_26/buf_output[5] , \SB2_4_26/buf_output[4] ,
         \SB2_4_26/buf_output[3] , \SB2_4_26/buf_output[2] ,
         \SB2_4_26/buf_output[1] , \SB2_4_26/buf_output[0] , \SB2_4_26/i3[0] ,
         \SB2_4_26/i1_5 , \SB2_4_26/i1_7 , \SB2_4_26/i1[9] , \SB2_4_26/i0_0 ,
         \SB2_4_26/i0_3 , \SB2_4_26/i0_4 , \SB2_4_26/i0[10] , \SB2_4_26/i0[9] ,
         \SB2_4_26/i0[8] , \SB2_4_26/i0[7] , \SB2_4_26/i0[6] ,
         \SB2_4_27/buf_output[5] , \SB2_4_27/buf_output[4] ,
         \SB2_4_27/buf_output[3] , \SB2_4_27/buf_output[2] ,
         \SB2_4_27/buf_output[1] , \SB2_4_27/buf_output[0] , \SB2_4_27/i3[0] ,
         \SB2_4_27/i1_5 , \SB2_4_27/i1_7 , \SB2_4_27/i1[9] , \SB2_4_27/i0_0 ,
         \SB2_4_27/i0_3 , \SB2_4_27/i0_4 , \SB2_4_27/i0[10] , \SB2_4_27/i0[9] ,
         \SB2_4_27/i0[8] , \SB2_4_27/i0[7] , \SB2_4_27/i0[6] ,
         \SB2_4_28/buf_output[5] , \SB2_4_28/buf_output[4] ,
         \SB2_4_28/buf_output[3] , \SB2_4_28/buf_output[2] ,
         \SB2_4_28/buf_output[1] , \SB2_4_28/buf_output[0] , \SB2_4_28/i3[0] ,
         \SB2_4_28/i1_5 , \SB2_4_28/i1_7 , \SB2_4_28/i1[9] , \SB2_4_28/i0_0 ,
         \SB2_4_28/i0_3 , \SB2_4_28/i0_4 , \SB2_4_28/i0[10] , \SB2_4_28/i0[9] ,
         \SB2_4_28/i0[7] , \SB2_4_28/i0[6] , \SB2_4_29/buf_output[5] ,
         \SB2_4_29/buf_output[4] , \SB2_4_29/buf_output[3] ,
         \SB2_4_29/buf_output[2] , \SB2_4_29/buf_output[1] ,
         \SB2_4_29/buf_output[0] , \SB2_4_29/i3[0] , \SB2_4_29/i1_5 ,
         \SB2_4_29/i1_7 , \SB2_4_29/i1[9] , \SB2_4_29/i0_0 , \SB2_4_29/i0_3 ,
         \SB2_4_29/i0_4 , \SB2_4_29/i0[10] , \SB2_4_29/i0[9] ,
         \SB2_4_29/i0[8] , \SB2_4_29/i0[7] , \SB2_4_29/i0[6] ,
         \SB2_4_30/buf_output[5] , \SB2_4_30/buf_output[4] ,
         \SB2_4_30/buf_output[3] , \SB2_4_30/buf_output[2] ,
         \SB2_4_30/buf_output[1] , \SB2_4_30/buf_output[0] , \SB2_4_30/i1_5 ,
         \SB2_4_30/i1_7 , \SB2_4_30/i1[9] , \SB2_4_30/i0_0 , \SB2_4_30/i0_3 ,
         \SB2_4_30/i0[10] , \SB2_4_30/i0[9] , \SB2_4_30/i0[8] ,
         \SB2_4_30/i0[6] , \SB2_4_31/buf_output[5] , \SB2_4_31/buf_output[4] ,
         \SB2_4_31/buf_output[3] , \SB2_4_31/buf_output[2] ,
         \SB2_4_31/buf_output[1] , \SB2_4_31/buf_output[0] , \SB2_4_31/i3[0] ,
         \SB2_4_31/i1_5 , \SB2_4_31/i1_7 , \SB2_4_31/i1[9] , \SB2_4_31/i0_0 ,
         \SB2_4_31/i0_3 , \SB2_4_31/i0_4 , \SB2_4_31/i0[10] , \SB2_4_31/i0[9] ,
         \SB2_4_31/i0[8] , \SB2_4_31/i0[7] , \SB2_4_31/i0[6] ,
         \SB3_0/buf_output[5] , \SB3_0/buf_output[4] , \SB3_0/buf_output[3] ,
         \SB3_0/buf_output[2] , \SB3_0/buf_output[1] , \SB3_0/buf_output[0] ,
         \SB3_0/i3[0] , \SB3_0/i1_5 , \SB3_0/i1_7 , \SB3_0/i1[9] ,
         \SB3_0/i0_0 , \SB3_0/i0_3 , \SB3_0/i0_4 , \SB3_0/i0[10] ,
         \SB3_0/i0[9] , \SB3_0/i0[8] , \SB3_0/i0[7] , \SB3_0/i0[6] ,
         \SB3_1/buf_output[4] , \SB3_1/buf_output[3] , \SB3_1/buf_output[1] ,
         \SB3_1/buf_output[0] , \SB3_1/i3[0] , \SB3_1/i1_5 , \SB3_1/i1_7 ,
         \SB3_1/i1[9] , \SB3_1/i0_0 , \SB3_1/i0_3 , \SB3_1/i0_4 ,
         \SB3_1/i0[10] , \SB3_1/i0[9] , \SB3_1/i0[8] , \SB3_1/i0[7] ,
         \SB3_1/i0[6] , \SB3_2/buf_output[5] , \SB3_2/buf_output[4] ,
         \SB3_2/buf_output[3] , \SB3_2/buf_output[2] , \SB3_2/buf_output[1] ,
         \SB3_2/buf_output[0] , \SB3_2/i3[0] , \SB3_2/i1_5 , \SB3_2/i1_7 ,
         \SB3_2/i1[9] , \SB3_2/i0_0 , \SB3_2/i0_3 , \SB3_2/i0_4 ,
         \SB3_2/i0[10] , \SB3_2/i0[9] , \SB3_2/i0[8] , \SB3_2/i0[7] ,
         \SB3_2/i0[6] , \SB3_3/buf_output[5] , \SB3_3/buf_output[4] ,
         \SB3_3/buf_output[3] , \SB3_3/buf_output[2] , \SB3_3/buf_output[1] ,
         \SB3_3/buf_output[0] , \SB3_3/i3[0] , \SB3_3/i1_5 , \SB3_3/i1_7 ,
         \SB3_3/i1[9] , \SB3_3/i0_0 , \SB3_3/i0_3 , \SB3_3/i0_4 ,
         \SB3_3/i0[10] , \SB3_3/i0[9] , \SB3_3/i0[8] , \SB3_3/i0[7] ,
         \SB3_3/i0[6] , \SB3_4/buf_output[5] , \SB3_4/buf_output[4] ,
         \SB3_4/buf_output[3] , \SB3_4/buf_output[2] , \SB3_4/buf_output[1] ,
         \SB3_4/buf_output[0] , \SB3_4/i3[0] , \SB3_4/i1_5 , \SB3_4/i1_7 ,
         \SB3_4/i1[9] , \SB3_4/i0_0 , \SB3_4/i0_3 , \SB3_4/i0_4 ,
         \SB3_4/i0[10] , \SB3_4/i0[9] , \SB3_4/i0[8] , \SB3_4/i0[7] ,
         \SB3_4/i0[6] , \SB3_5/buf_output[5] , \SB3_5/buf_output[4] ,
         \SB3_5/buf_output[2] , \SB3_5/buf_output[1] , \SB3_5/buf_output[0] ,
         \SB3_5/i3[0] , \SB3_5/i1_5 , \SB3_5/i1_7 , \SB3_5/i1[9] ,
         \SB3_5/i0_0 , \SB3_5/i0_3 , \SB3_5/i0_4 , \SB3_5/i0[10] ,
         \SB3_5/i0[9] , \SB3_5/i0[8] , \SB3_5/i0[7] , \SB3_5/i0[6] ,
         \SB3_6/buf_output[5] , \SB3_6/buf_output[4] , \SB3_6/buf_output[3] ,
         \SB3_6/buf_output[2] , \SB3_6/buf_output[1] , \SB3_6/buf_output[0] ,
         \SB3_6/i3[0] , \SB3_6/i1_5 , \SB3_6/i1_7 , \SB3_6/i1[9] ,
         \SB3_6/i0_0 , \SB3_6/i0_3 , \SB3_6/i0_4 , \SB3_6/i0[10] ,
         \SB3_6/i0[9] , \SB3_6/i0[8] , \SB3_6/i0[7] , \SB3_6/i0[6] ,
         \SB3_7/buf_output[4] , \SB3_7/buf_output[3] , \SB3_7/buf_output[2] ,
         \SB3_7/buf_output[1] , \SB3_7/buf_output[0] , \SB3_7/i3[0] ,
         \SB3_7/i1_5 , \SB3_7/i1_7 , \SB3_7/i1[9] , \SB3_7/i0_0 , \SB3_7/i0_3 ,
         \SB3_7/i0_4 , \SB3_7/i0[10] , \SB3_7/i0[9] , \SB3_7/i0[8] ,
         \SB3_7/i0[7] , \SB3_7/i0[6] , \SB3_8/buf_output[5] ,
         \SB3_8/buf_output[4] , \SB3_8/buf_output[3] , \SB3_8/buf_output[2] ,
         \SB3_8/buf_output[1] , \SB3_8/buf_output[0] , \SB3_8/i3[0] ,
         \SB3_8/i1_5 , \SB3_8/i1_7 , \SB3_8/i1[9] , \SB3_8/i0_0 , \SB3_8/i0_3 ,
         \SB3_8/i0_4 , \SB3_8/i0[10] , \SB3_8/i0[9] , \SB3_8/i0[8] ,
         \SB3_8/i0[7] , \SB3_8/i0[6] , \SB3_9/buf_output[5] ,
         \SB3_9/buf_output[4] , \SB3_9/buf_output[3] , \SB3_9/buf_output[2] ,
         \SB3_9/buf_output[1] , \SB3_9/buf_output[0] , \SB3_9/i3[0] ,
         \SB3_9/i1_5 , \SB3_9/i1_7 , \SB3_9/i1[9] , \SB3_9/i0_0 , \SB3_9/i0_3 ,
         \SB3_9/i0_4 , \SB3_9/i0[10] , \SB3_9/i0[9] , \SB3_9/i0[8] ,
         \SB3_9/i0[7] , \SB3_9/i0[6] , \SB3_10/buf_output[5] ,
         \SB3_10/buf_output[4] , \SB3_10/buf_output[3] ,
         \SB3_10/buf_output[2] , \SB3_10/buf_output[1] ,
         \SB3_10/buf_output[0] , \SB3_10/i3[0] , \SB3_10/i1_5 , \SB3_10/i1_7 ,
         \SB3_10/i1[9] , \SB3_10/i0_0 , \SB3_10/i0_3 , \SB3_10/i0_4 ,
         \SB3_10/i0[10] , \SB3_10/i0[9] , \SB3_10/i0[8] , \SB3_10/i0[7] ,
         \SB3_10/i0[6] , \SB3_11/buf_output[5] , \SB3_11/buf_output[4] ,
         \SB3_11/buf_output[1] , \SB3_11/buf_output[0] , \SB3_11/i3[0] ,
         \SB3_11/i1_5 , \SB3_11/i1_7 , \SB3_11/i1[9] , \SB3_11/i0_0 ,
         \SB3_11/i0_3 , \SB3_11/i0_4 , \SB3_11/i0[10] , \SB3_11/i0[9] ,
         \SB3_11/i0[8] , \SB3_11/i0[7] , \SB3_11/i0[6] ,
         \SB3_12/buf_output[5] , \SB3_12/buf_output[4] ,
         \SB3_12/buf_output[3] , \SB3_12/buf_output[2] ,
         \SB3_12/buf_output[1] , \SB3_12/buf_output[0] , \SB3_12/i3[0] ,
         \SB3_12/i1_5 , \SB3_12/i1_7 , \SB3_12/i1[9] , \SB3_12/i0_0 ,
         \SB3_12/i0_4 , \SB3_12/i0[10] , \SB3_12/i0[9] , \SB3_12/i0[8] ,
         \SB3_12/i0[7] , \SB3_12/i0[6] , \SB3_13/buf_output[5] ,
         \SB3_13/buf_output[4] , \SB3_13/buf_output[3] ,
         \SB3_13/buf_output[1] , \SB3_13/buf_output[0] , \SB3_13/i3[0] ,
         \SB3_13/i1_5 , \SB3_13/i1_7 , \SB3_13/i1[9] , \SB3_13/i0_0 ,
         \SB3_13/i0_3 , \SB3_13/i0_4 , \SB3_13/i0[10] , \SB3_13/i0[9] ,
         \SB3_13/i0[8] , \SB3_13/i0[7] , \SB3_13/i0[6] ,
         \SB3_14/buf_output[5] , \SB3_14/buf_output[4] ,
         \SB3_14/buf_output[3] , \SB3_14/buf_output[2] ,
         \SB3_14/buf_output[1] , \SB3_14/buf_output[0] , \SB3_14/i3[0] ,
         \SB3_14/i1_5 , \SB3_14/i1_7 , \SB3_14/i1[9] , \SB3_14/i0_0 ,
         \SB3_14/i0_3 , \SB3_14/i0_4 , \SB3_14/i0[10] , \SB3_14/i0[9] ,
         \SB3_14/i0[8] , \SB3_14/i0[7] , \SB3_14/i0[6] ,
         \SB3_15/buf_output[5] , \SB3_15/buf_output[4] ,
         \SB3_15/buf_output[3] , \SB3_15/buf_output[2] ,
         \SB3_15/buf_output[1] , \SB3_15/buf_output[0] , \SB3_15/i3[0] ,
         \SB3_15/i1_5 , \SB3_15/i1_7 , \SB3_15/i1[9] , \SB3_15/i0_0 ,
         \SB3_15/i0_3 , \SB3_15/i0_4 , \SB3_15/i0[10] , \SB3_15/i0[9] ,
         \SB3_15/i0[8] , \SB3_15/i0[7] , \SB3_15/i0[6] ,
         \SB3_16/buf_output[5] , \SB3_16/buf_output[4] ,
         \SB3_16/buf_output[3] , \SB3_16/buf_output[2] ,
         \SB3_16/buf_output[1] , \SB3_16/buf_output[0] , \SB3_16/i3[0] ,
         \SB3_16/i1_5 , \SB3_16/i1_7 , \SB3_16/i1[9] , \SB3_16/i0_0 ,
         \SB3_16/i0_3 , \SB3_16/i0_4 , \SB3_16/i0[10] , \SB3_16/i0[9] ,
         \SB3_16/i0[8] , \SB3_16/i0[7] , \SB3_16/i0[6] ,
         \SB3_17/buf_output[5] , \SB3_17/buf_output[4] ,
         \SB3_17/buf_output[3] , \SB3_17/buf_output[2] ,
         \SB3_17/buf_output[1] , \SB3_17/buf_output[0] , \SB3_17/i3[0] ,
         \SB3_17/i1_5 , \SB3_17/i1_7 , \SB3_17/i1[9] , \SB3_17/i0_0 ,
         \SB3_17/i0_3 , \SB3_17/i0_4 , \SB3_17/i0[10] , \SB3_17/i0[9] ,
         \SB3_17/i0[8] , \SB3_17/i0[7] , \SB3_17/i0[6] ,
         \SB3_18/buf_output[5] , \SB3_18/buf_output[4] ,
         \SB3_18/buf_output[3] , \SB3_18/buf_output[2] ,
         \SB3_18/buf_output[1] , \SB3_18/buf_output[0] , \SB3_18/i3[0] ,
         \SB3_18/i1_5 , \SB3_18/i1_7 , \SB3_18/i1[9] , \SB3_18/i0_0 ,
         \SB3_18/i0_3 , \SB3_18/i0_4 , \SB3_18/i0[10] , \SB3_18/i0[9] ,
         \SB3_18/i0[8] , \SB3_18/i0[7] , \SB3_18/i0[6] ,
         \SB3_19/buf_output[5] , \SB3_19/buf_output[4] ,
         \SB3_19/buf_output[2] , \SB3_19/buf_output[1] ,
         \SB3_19/buf_output[0] , \SB3_19/i3[0] , \SB3_19/i1_5 , \SB3_19/i1_7 ,
         \SB3_19/i1[9] , \SB3_19/i0_0 , \SB3_19/i0_3 , \SB3_19/i0_4 ,
         \SB3_19/i0[10] , \SB3_19/i0[9] , \SB3_19/i0[8] , \SB3_19/i0[7] ,
         \SB3_19/i0[6] , \SB3_20/buf_output[5] , \SB3_20/buf_output[4] ,
         \SB3_20/buf_output[3] , \SB3_20/buf_output[2] ,
         \SB3_20/buf_output[1] , \SB3_20/buf_output[0] , \SB3_20/i3[0] ,
         \SB3_20/i1_5 , \SB3_20/i1_7 , \SB3_20/i1[9] , \SB3_20/i0_0 ,
         \SB3_20/i0_3 , \SB3_20/i0_4 , \SB3_20/i0[10] , \SB3_20/i0[9] ,
         \SB3_20/i0[8] , \SB3_20/i0[7] , \SB3_20/i0[6] ,
         \SB3_21/buf_output[5] , \SB3_21/buf_output[4] ,
         \SB3_21/buf_output[3] , \SB3_21/buf_output[1] ,
         \SB3_21/buf_output[0] , \SB3_21/i3[0] , \SB3_21/i1_7 , \SB3_21/i1[9] ,
         \SB3_21/i0_0 , \SB3_21/i0_3 , \SB3_21/i0_4 , \SB3_21/i0[10] ,
         \SB3_21/i0[9] , \SB3_21/i0[8] , \SB3_21/i0[7] , \SB3_21/i0[6] ,
         \SB3_22/buf_output[5] , \SB3_22/buf_output[4] ,
         \SB3_22/buf_output[3] , \SB3_22/buf_output[2] ,
         \SB3_22/buf_output[1] , \SB3_22/buf_output[0] , \SB3_22/i3[0] ,
         \SB3_22/i1_5 , \SB3_22/i1_7 , \SB3_22/i1[9] , \SB3_22/i0_0 ,
         \SB3_22/i0_3 , \SB3_22/i0_4 , \SB3_22/i0[10] , \SB3_22/i0[9] ,
         \SB3_22/i0[8] , \SB3_22/i0[7] , \SB3_22/i0[6] ,
         \SB3_23/buf_output[5] , \SB3_23/buf_output[4] ,
         \SB3_23/buf_output[3] , \SB3_23/buf_output[2] ,
         \SB3_23/buf_output[0] , \SB3_23/i3[0] , \SB3_23/i1_5 , \SB3_23/i1_7 ,
         \SB3_23/i1[9] , \SB3_23/i0_0 , \SB3_23/i0_3 , \SB3_23/i0_4 ,
         \SB3_23/i0[10] , \SB3_23/i0[9] , \SB3_23/i0[8] , \SB3_23/i0[7] ,
         \SB3_23/i0[6] , \SB3_24/buf_output[5] , \SB3_24/buf_output[4] ,
         \SB3_24/buf_output[3] , \SB3_24/buf_output[2] ,
         \SB3_24/buf_output[1] , \SB3_24/buf_output[0] , \SB3_24/i3[0] ,
         \SB3_24/i1_5 , \SB3_24/i1_7 , \SB3_24/i1[9] , \SB3_24/i0_0 ,
         \SB3_24/i0_3 , \SB3_24/i0_4 , \SB3_24/i0[10] , \SB3_24/i0[9] ,
         \SB3_24/i0[8] , \SB3_24/i0[7] , \SB3_24/i0[6] ,
         \SB3_25/buf_output[5] , \SB3_25/buf_output[4] ,
         \SB3_25/buf_output[2] , \SB3_25/buf_output[1] ,
         \SB3_25/buf_output[0] , \SB3_25/i3[0] , \SB3_25/i1_5 , \SB3_25/i1_7 ,
         \SB3_25/i1[9] , \SB3_25/i0_0 , \SB3_25/i0_3 , \SB3_25/i0_4 ,
         \SB3_25/i0[10] , \SB3_25/i0[9] , \SB3_25/i0[8] , \SB3_25/i0[7] ,
         \SB3_25/i0[6] , \SB3_26/buf_output[5] , \SB3_26/buf_output[4] ,
         \SB3_26/buf_output[3] , \SB3_26/buf_output[2] ,
         \SB3_26/buf_output[1] , \SB3_26/buf_output[0] , \SB3_26/i3[0] ,
         \SB3_26/i1_5 , \SB3_26/i1_7 , \SB3_26/i1[9] , \SB3_26/i0_0 ,
         \SB3_26/i0_3 , \SB3_26/i0_4 , \SB3_26/i0[10] , \SB3_26/i0[9] ,
         \SB3_26/i0[8] , \SB3_26/i0[7] , \SB3_26/i0[6] ,
         \SB3_27/buf_output[5] , \SB3_27/buf_output[4] ,
         \SB3_27/buf_output[3] , \SB3_27/buf_output[2] ,
         \SB3_27/buf_output[1] , \SB3_27/buf_output[0] , \SB3_27/i3[0] ,
         \SB3_27/i1_5 , \SB3_27/i1_7 , \SB3_27/i1[9] , \SB3_27/i0_0 ,
         \SB3_27/i0_3 , \SB3_27/i0_4 , \SB3_27/i0[10] , \SB3_27/i0[9] ,
         \SB3_27/i0[8] , \SB3_27/i0[7] , \SB3_27/i0[6] ,
         \SB3_28/buf_output[5] , \SB3_28/buf_output[4] ,
         \SB3_28/buf_output[2] , \SB3_28/buf_output[1] ,
         \SB3_28/buf_output[0] , \SB3_28/i3[0] , \SB3_28/i1_5 , \SB3_28/i1_7 ,
         \SB3_28/i1[9] , \SB3_28/i0_0 , \SB3_28/i0_3 , \SB3_28/i0_4 ,
         \SB3_28/i0[10] , \SB3_28/i0[9] , \SB3_28/i0[8] , \SB3_28/i0[7] ,
         \SB3_28/i0[6] , \SB3_29/buf_output[5] , \SB3_29/buf_output[4] ,
         \SB3_29/buf_output[3] , \SB3_29/buf_output[2] ,
         \SB3_29/buf_output[1] , \SB3_29/buf_output[0] , \SB3_29/i3[0] ,
         \SB3_29/i1_5 , \SB3_29/i1_7 , \SB3_29/i1[9] , \SB3_29/i0_0 ,
         \SB3_29/i0_4 , \SB3_29/i0[10] , \SB3_29/i0[9] , \SB3_29/i0[8] ,
         \SB3_29/i0[7] , \SB3_29/i0[6] , \SB3_30/buf_output[5] ,
         \SB3_30/buf_output[4] , \SB3_30/buf_output[3] ,
         \SB3_30/buf_output[2] , \SB3_30/buf_output[1] , \SB3_30/i3[0] ,
         \SB3_30/i1_5 , \SB3_30/i1_7 , \SB3_30/i1[9] , \SB3_30/i0_0 ,
         \SB3_30/i0_3 , \SB3_30/i0_4 , \SB3_30/i0[10] , \SB3_30/i0[9] ,
         \SB3_30/i0[8] , \SB3_30/i0[7] , \SB3_30/i0[6] ,
         \SB3_31/buf_output[5] , \SB3_31/buf_output[4] ,
         \SB3_31/buf_output[3] , \SB3_31/buf_output[2] ,
         \SB3_31/buf_output[1] , \SB3_31/buf_output[0] , \SB3_31/i3[0] ,
         \SB3_31/i1_5 , \SB3_31/i1_7 , \SB3_31/i1[9] , \SB3_31/i0_0 ,
         \SB3_31/i0_3 , \SB3_31/i0_4 , \SB3_31/i0[10] , \SB3_31/i0[9] ,
         \SB3_31/i0[8] , \SB3_31/i0[7] , \SB3_31/i0[6] , \SB4_0/i3[0] ,
         \SB4_0/i1_5 , \SB4_0/i1_7 , \SB4_0/i1[9] , \SB4_0/i0_0 , \SB4_0/i0_3 ,
         \SB4_0/i0_4 , \SB4_0/i0[10] , \SB4_0/i0[9] , \SB4_0/i0[8] ,
         \SB4_0/i0[7] , \SB4_0/i0[6] , \SB4_1/i3[0] , \SB4_1/i1_7 ,
         \SB4_1/i1[9] , \SB4_1/i0_0 , \SB4_1/i0_3 , \SB4_1/i0_4 ,
         \SB4_1/i0[10] , \SB4_1/i0[9] , \SB4_1/i0[8] , \SB4_1/i0[7] ,
         \SB4_1/i0[6] , \SB4_2/i3[0] , \SB4_2/i1_5 , \SB4_2/i1_7 ,
         \SB4_2/i1[9] , \SB4_2/i0_0 , \SB4_2/i0_3 , \SB4_2/i0_4 ,
         \SB4_2/i0[10] , \SB4_2/i0[9] , \SB4_2/i0[8] , \SB4_2/i0[7] ,
         \SB4_2/i0[6] , \SB4_3/i3[0] , \SB4_3/i1_5 , \SB4_3/i1_7 ,
         \SB4_3/i1[9] , \SB4_3/i0_0 , \SB4_3/i0_3 , \SB4_3/i0_4 ,
         \SB4_3/i0[10] , \SB4_3/i0[9] , \SB4_3/i0[8] , \SB4_3/i0[7] ,
         \SB4_3/i0[6] , \SB4_4/i3[0] , \SB4_4/i1_5 , \SB4_4/i1_7 ,
         \SB4_4/i1[9] , \SB4_4/i0_0 , \SB4_4/i0_3 , \SB4_4/i0_4 ,
         \SB4_4/i0[10] , \SB4_4/i0[9] , \SB4_4/i0[8] , \SB4_4/i0[7] ,
         \SB4_4/i0[6] , \SB4_5/i3[0] , \SB4_5/i1_5 , \SB4_5/i1_7 ,
         \SB4_5/i1[9] , \SB4_5/i0_0 , \SB4_5/i0_3 , \SB4_5/i0_4 ,
         \SB4_5/i0[10] , \SB4_5/i0[9] , \SB4_5/i0[8] , \SB4_5/i0[7] ,
         \SB4_5/i0[6] , \SB4_6/i3[0] , \SB4_6/i1_5 , \SB4_6/i1_7 ,
         \SB4_6/i1[9] , \SB4_6/i0_0 , \SB4_6/i0_3 , \SB4_6/i0_4 ,
         \SB4_6/i0[10] , \SB4_6/i0[9] , \SB4_6/i0[8] , \SB4_6/i0[7] ,
         \SB4_6/i0[6] , \SB4_7/i3[0] , \SB4_7/i1_5 , \SB4_7/i1_7 ,
         \SB4_7/i1[9] , \SB4_7/i0_0 , \SB4_7/i0_3 , \SB4_7/i0_4 ,
         \SB4_7/i0[9] , \SB4_7/i0[7] , \SB4_7/i0[6] , \SB4_8/i3[0] ,
         \SB4_8/i1_5 , \SB4_8/i1_7 , \SB4_8/i0_0 , \SB4_8/i0_3 , \SB4_8/i0_4 ,
         \SB4_8/i0[10] , \SB4_8/i0[9] , \SB4_8/i0[8] , \SB4_8/i0[7] ,
         \SB4_8/i0[6] , \SB4_9/i3[0] , \SB4_9/i1_5 , \SB4_9/i1_7 ,
         \SB4_9/i1[9] , \SB4_9/i0_0 , \SB4_9/i0_3 , \SB4_9/i0[10] ,
         \SB4_9/i0[9] , \SB4_9/i0[7] , \SB4_9/i0[6] , \SB4_10/i3[0] ,
         \SB4_10/i1_5 , \SB4_10/i1_7 , \SB4_10/i1[9] , \SB4_10/i0_0 ,
         \SB4_10/i0_3 , \SB4_10/i0_4 , \SB4_10/i0[10] , \SB4_10/i0[9] ,
         \SB4_10/i0[8] , \SB4_10/i0[7] , \SB4_10/i0[6] , \SB4_11/i3[0] ,
         \SB4_11/i1_5 , \SB4_11/i1_7 , \SB4_11/i1[9] , \SB4_11/i0_0 ,
         \SB4_11/i0_3 , \SB4_11/i0_4 , \SB4_11/i0[10] , \SB4_11/i0[9] ,
         \SB4_11/i0[8] , \SB4_11/i0[7] , \SB4_11/i0[6] , \SB4_12/i3[0] ,
         \SB4_12/i1_5 , \SB4_12/i1_7 , \SB4_12/i1[9] , \SB4_12/i0_0 ,
         \SB4_12/i0_3 , \SB4_12/i0_4 , \SB4_12/i0[10] , \SB4_12/i0[9] ,
         \SB4_12/i0[8] , \SB4_12/i0[7] , \SB4_12/i0[6] , \SB4_13/i3[0] ,
         \SB4_13/i1_7 , \SB4_13/i1[9] , \SB4_13/i0_0 , \SB4_13/i0_3 ,
         \SB4_13/i0_4 , \SB4_13/i0[9] , \SB4_13/i0[7] , \SB4_13/i0[6] ,
         \SB4_14/i3[0] , \SB4_14/i1_7 , \SB4_14/i1[9] , \SB4_14/i0_0 ,
         \SB4_14/i0_3 , \SB4_14/i0_4 , \SB4_14/i0[10] , \SB4_14/i0[9] ,
         \SB4_14/i0[8] , \SB4_14/i0[7] , \SB4_14/i0[6] , \SB4_15/i3[0] ,
         \SB4_15/i1_5 , \SB4_15/i1_7 , \SB4_15/i1[9] , \SB4_15/i0_0 ,
         \SB4_15/i0_3 , \SB4_15/i0_4 , \SB4_15/i0[9] , \SB4_15/i0[7] ,
         \SB4_15/i0[6] , \SB4_16/i3[0] , \SB4_16/i1_5 , \SB4_16/i1_7 ,
         \SB4_16/i1[9] , \SB4_16/i0_0 , \SB4_16/i0_3 , \SB4_16/i0_4 ,
         \SB4_16/i0[10] , \SB4_16/i0[9] , \SB4_16/i0[8] , \SB4_16/i0[7] ,
         \SB4_16/i0[6] , \SB4_17/i3[0] , \SB4_17/i1_7 , \SB4_17/i1[9] ,
         \SB4_17/i0_0 , \SB4_17/i0_3 , \SB4_17/i0_4 , \SB4_17/i0[10] ,
         \SB4_17/i0[9] , \SB4_17/i0[7] , \SB4_17/i0[6] , \SB4_18/i3[0] ,
         \SB4_18/i1_5 , \SB4_18/i1_7 , \SB4_18/i0_0 , \SB4_18/i0_3 ,
         \SB4_18/i0_4 , \SB4_18/i0[10] , \SB4_18/i0[9] , \SB4_18/i0[8] ,
         \SB4_18/i0[7] , \SB4_18/i0[6] , \SB4_19/i3[0] , \SB4_19/i1_7 ,
         \SB4_19/i1[9] , \SB4_19/i0_0 , \SB4_19/i0_3 , \SB4_19/i0_4 ,
         \SB4_19/i0[10] , \SB4_19/i0[9] , \SB4_19/i0[8] , \SB4_19/i0[7] ,
         \SB4_19/i0[6] , \SB4_20/i3[0] , \SB4_20/i1_5 , \SB4_20/i1_7 ,
         \SB4_20/i1[9] , \SB4_20/i0_0 , \SB4_20/i0_3 , \SB4_20/i0_4 ,
         \SB4_20/i0[10] , \SB4_20/i0[9] , \SB4_20/i0[8] , \SB4_20/i0[7] ,
         \SB4_20/i0[6] , \SB4_21/i3[0] , \SB4_21/i1_5 , \SB4_21/i1_7 ,
         \SB4_21/i0_3 , \SB4_21/i0_4 , \SB4_21/i0[10] , \SB4_21/i0[9] ,
         \SB4_21/i0[8] , \SB4_21/i0[7] , \SB4_21/i0[6] , \SB4_22/i3[0] ,
         \SB4_22/i1_5 , \SB4_22/i1_7 , \SB4_22/i1[9] , \SB4_22/i0_0 ,
         \SB4_22/i0_3 , \SB4_22/i0_4 , \SB4_22/i0[10] , \SB4_22/i0[9] ,
         \SB4_22/i0[8] , \SB4_22/i0[7] , \SB4_22/i0[6] , \SB4_23/i3[0] ,
         \SB4_23/i1_5 , \SB4_23/i1_7 , \SB4_23/i1[9] , \SB4_23/i0_0 ,
         \SB4_23/i0_3 , \SB4_23/i0_4 , \SB4_23/i0[10] , \SB4_23/i0[9] ,
         \SB4_23/i0[7] , \SB4_23/i0[6] , \SB4_24/i3[0] , \SB4_24/i1_5 ,
         \SB4_24/i1_7 , \SB4_24/i1[9] , \SB4_24/i0_0 , \SB4_24/i0_3 ,
         \SB4_24/i0_4 , \SB4_24/i0[9] , \SB4_24/i0[7] , \SB4_24/i0[6] ,
         \SB4_25/i1_5 , \SB4_25/i1_7 , \SB4_25/i1[9] , \SB4_25/i0_0 ,
         \SB4_25/i0_3 , \SB4_25/i0_4 , \SB4_25/i0[10] , \SB4_25/i0[8] ,
         \SB4_25/i0[7] , \SB4_25/i0[6] , \SB4_26/i3[0] , \SB4_26/i1_5 ,
         \SB4_26/i1_7 , \SB4_26/i0_3 , \SB4_26/i0_4 , \SB4_26/i0[10] ,
         \SB4_26/i0[9] , \SB4_26/i0[7] , \SB4_26/i0[6] , \SB4_27/i3[0] ,
         \SB4_27/i1_5 , \SB4_27/i1_7 , \SB4_27/i1[9] , \SB4_27/i0_0 ,
         \SB4_27/i0_3 , \SB4_27/i0_4 , \SB4_27/i0[10] , \SB4_27/i0[9] ,
         \SB4_27/i0[8] , \SB4_27/i0[7] , \SB4_27/i0[6] , \SB4_28/i3[0] ,
         \SB4_28/i1_5 , \SB4_28/i1_7 , \SB4_28/i1[9] , \SB4_28/i0_0 ,
         \SB4_28/i0_3 , \SB4_28/i0_4 , \SB4_28/i0[10] , \SB4_28/i0[9] ,
         \SB4_28/i0[8] , \SB4_28/i0[7] , \SB4_28/i0[6] , \SB4_29/i3[0] ,
         \SB4_29/i1_5 , \SB4_29/i1_7 , \SB4_29/i1[9] , \SB4_29/i0_0 ,
         \SB4_29/i0_3 , \SB4_29/i0_4 , \SB4_29/i0[10] , \SB4_29/i0[9] ,
         \SB4_29/i0[8] , \SB4_29/i0[7] , \SB4_29/i0[6] , \SB4_30/i3[0] ,
         \SB4_30/i1_5 , \SB4_30/i1_7 , \SB4_30/i0_0 , \SB4_30/i0_3 ,
         \SB4_30/i0_4 , \SB4_30/i0[10] , \SB4_30/i0[9] , \SB4_30/i0[8] ,
         \SB4_30/i0[7] , \SB4_30/i0[6] , \SB4_31/i3[0] , \SB4_31/i1_5 ,
         \SB4_31/i1_7 , \SB4_31/i1[9] , \SB4_31/i0_0 , \SB4_31/i0_3 ,
         \SB4_31/i0_4 , \SB4_31/i0[10] , \SB4_31/i0[9] , \SB4_31/i0[8] ,
         \SB4_31/i0[7] , \SB4_31/i0[6] ,
         \SB1_0_0/Component_Function_2/NAND4_in[0] ,
         \SB1_0_0/Component_Function_3/NAND4_in[3] ,
         \SB1_0_0/Component_Function_3/NAND4_in[0] ,
         \SB1_0_0/Component_Function_4/NAND4_in[1] ,
         \SB1_0_0/Component_Function_4/NAND4_in[0] ,
         \SB1_0_1/Component_Function_2/NAND4_in[2] ,
         \SB1_0_1/Component_Function_2/NAND4_in[1] ,
         \SB1_0_1/Component_Function_2/NAND4_in[0] ,
         \SB1_0_1/Component_Function_3/NAND4_in[3] ,
         \SB1_0_1/Component_Function_3/NAND4_in[2] ,
         \SB1_0_1/Component_Function_3/NAND4_in[1] ,
         \SB1_0_1/Component_Function_3/NAND4_in[0] ,
         \SB1_0_1/Component_Function_4/NAND4_in[2] ,
         \SB1_0_1/Component_Function_4/NAND4_in[1] ,
         \SB1_0_1/Component_Function_4/NAND4_in[0] ,
         \SB1_0_2/Component_Function_2/NAND4_in[2] ,
         \SB1_0_2/Component_Function_2/NAND4_in[1] ,
         \SB1_0_2/Component_Function_2/NAND4_in[0] ,
         \SB1_0_2/Component_Function_3/NAND4_in[3] ,
         \SB1_0_2/Component_Function_3/NAND4_in[1] ,
         \SB1_0_2/Component_Function_3/NAND4_in[0] ,
         \SB1_0_2/Component_Function_4/NAND4_in[3] ,
         \SB1_0_2/Component_Function_4/NAND4_in[2] ,
         \SB1_0_2/Component_Function_4/NAND4_in[1] ,
         \SB1_0_2/Component_Function_4/NAND4_in[0] ,
         \SB1_0_3/Component_Function_2/NAND4_in[3] ,
         \SB1_0_3/Component_Function_2/NAND4_in[2] ,
         \SB1_0_3/Component_Function_3/NAND4_in[3] ,
         \SB1_0_3/Component_Function_3/NAND4_in[0] ,
         \SB1_0_3/Component_Function_4/NAND4_in[3] ,
         \SB1_0_3/Component_Function_4/NAND4_in[2] ,
         \SB1_0_3/Component_Function_4/NAND4_in[1] ,
         \SB1_0_3/Component_Function_4/NAND4_in[0] ,
         \SB1_0_4/Component_Function_2/NAND4_in[2] ,
         \SB1_0_4/Component_Function_2/NAND4_in[1] ,
         \SB1_0_4/Component_Function_3/NAND4_in[3] ,
         \SB1_0_4/Component_Function_3/NAND4_in[1] ,
         \SB1_0_4/Component_Function_3/NAND4_in[0] ,
         \SB1_0_4/Component_Function_4/NAND4_in[2] ,
         \SB1_0_4/Component_Function_4/NAND4_in[1] ,
         \SB1_0_4/Component_Function_4/NAND4_in[0] ,
         \SB1_0_5/Component_Function_2/NAND4_in[2] ,
         \SB1_0_5/Component_Function_2/NAND4_in[0] ,
         \SB1_0_5/Component_Function_3/NAND4_in[3] ,
         \SB1_0_5/Component_Function_3/NAND4_in[1] ,
         \SB1_0_5/Component_Function_3/NAND4_in[0] ,
         \SB1_0_5/Component_Function_4/NAND4_in[3] ,
         \SB1_0_5/Component_Function_4/NAND4_in[1] ,
         \SB1_0_5/Component_Function_4/NAND4_in[0] ,
         \SB1_0_6/Component_Function_2/NAND4_in[2] ,
         \SB1_0_6/Component_Function_3/NAND4_in[3] ,
         \SB1_0_6/Component_Function_3/NAND4_in[2] ,
         \SB1_0_6/Component_Function_3/NAND4_in[1] ,
         \SB1_0_6/Component_Function_3/NAND4_in[0] ,
         \SB1_0_6/Component_Function_4/NAND4_in[3] ,
         \SB1_0_6/Component_Function_4/NAND4_in[1] ,
         \SB1_0_7/Component_Function_2/NAND4_in[2] ,
         \SB1_0_7/Component_Function_2/NAND4_in[1] ,
         \SB1_0_7/Component_Function_2/NAND4_in[0] ,
         \SB1_0_7/Component_Function_3/NAND4_in[3] ,
         \SB1_0_7/Component_Function_3/NAND4_in[2] ,
         \SB1_0_7/Component_Function_3/NAND4_in[1] ,
         \SB1_0_7/Component_Function_3/NAND4_in[0] ,
         \SB1_0_7/Component_Function_4/NAND4_in[3] ,
         \SB1_0_7/Component_Function_4/NAND4_in[1] ,
         \SB1_0_7/Component_Function_4/NAND4_in[0] ,
         \SB1_0_8/Component_Function_2/NAND4_in[2] ,
         \SB1_0_8/Component_Function_2/NAND4_in[1] ,
         \SB1_0_8/Component_Function_3/NAND4_in[3] ,
         \SB1_0_8/Component_Function_3/NAND4_in[1] ,
         \SB1_0_8/Component_Function_4/NAND4_in[3] ,
         \SB1_0_8/Component_Function_4/NAND4_in[1] ,
         \SB1_0_8/Component_Function_4/NAND4_in[0] ,
         \SB1_0_9/Component_Function_2/NAND4_in[2] ,
         \SB1_0_9/Component_Function_2/NAND4_in[1] ,
         \SB1_0_9/Component_Function_2/NAND4_in[0] ,
         \SB1_0_9/Component_Function_3/NAND4_in[3] ,
         \SB1_0_9/Component_Function_3/NAND4_in[1] ,
         \SB1_0_9/Component_Function_3/NAND4_in[0] ,
         \SB1_0_9/Component_Function_4/NAND4_in[3] ,
         \SB1_0_9/Component_Function_4/NAND4_in[2] ,
         \SB1_0_9/Component_Function_4/NAND4_in[1] ,
         \SB1_0_9/Component_Function_4/NAND4_in[0] ,
         \SB1_0_10/Component_Function_2/NAND4_in[2] ,
         \SB1_0_10/Component_Function_3/NAND4_in[2] ,
         \SB1_0_10/Component_Function_4/NAND4_in[2] ,
         \SB1_0_10/Component_Function_4/NAND4_in[0] ,
         \SB1_0_11/Component_Function_2/NAND4_in[2] ,
         \SB1_0_11/Component_Function_3/NAND4_in[3] ,
         \SB1_0_11/Component_Function_3/NAND4_in[1] ,
         \SB1_0_11/Component_Function_3/NAND4_in[0] ,
         \SB1_0_11/Component_Function_4/NAND4_in[3] ,
         \SB1_0_11/Component_Function_4/NAND4_in[2] ,
         \SB1_0_11/Component_Function_4/NAND4_in[1] ,
         \SB1_0_12/Component_Function_2/NAND4_in[2] ,
         \SB1_0_12/Component_Function_3/NAND4_in[3] ,
         \SB1_0_12/Component_Function_3/NAND4_in[1] ,
         \SB1_0_12/Component_Function_3/NAND4_in[0] ,
         \SB1_0_12/Component_Function_4/NAND4_in[3] ,
         \SB1_0_12/Component_Function_4/NAND4_in[2] ,
         \SB1_0_12/Component_Function_4/NAND4_in[1] ,
         \SB1_0_12/Component_Function_4/NAND4_in[0] ,
         \SB1_0_13/Component_Function_2/NAND4_in[3] ,
         \SB1_0_13/Component_Function_2/NAND4_in[2] ,
         \SB1_0_13/Component_Function_2/NAND4_in[1] ,
         \SB1_0_13/Component_Function_2/NAND4_in[0] ,
         \SB1_0_13/Component_Function_3/NAND4_in[3] ,
         \SB1_0_13/Component_Function_3/NAND4_in[2] ,
         \SB1_0_13/Component_Function_3/NAND4_in[1] ,
         \SB1_0_13/Component_Function_3/NAND4_in[0] ,
         \SB1_0_13/Component_Function_4/NAND4_in[3] ,
         \SB1_0_13/Component_Function_4/NAND4_in[1] ,
         \SB1_0_13/Component_Function_4/NAND4_in[0] ,
         \SB1_0_14/Component_Function_2/NAND4_in[1] ,
         \SB1_0_14/Component_Function_2/NAND4_in[0] ,
         \SB1_0_14/Component_Function_3/NAND4_in[3] ,
         \SB1_0_14/Component_Function_3/NAND4_in[2] ,
         \SB1_0_14/Component_Function_3/NAND4_in[1] ,
         \SB1_0_14/Component_Function_4/NAND4_in[3] ,
         \SB1_0_14/Component_Function_4/NAND4_in[1] ,
         \SB1_0_14/Component_Function_4/NAND4_in[0] ,
         \SB1_0_15/Component_Function_2/NAND4_in[2] ,
         \SB1_0_15/Component_Function_2/NAND4_in[0] ,
         \SB1_0_15/Component_Function_3/NAND4_in[3] ,
         \SB1_0_15/Component_Function_3/NAND4_in[2] ,
         \SB1_0_15/Component_Function_3/NAND4_in[1] ,
         \SB1_0_15/Component_Function_4/NAND4_in[3] ,
         \SB1_0_15/Component_Function_4/NAND4_in[1] ,
         \SB1_0_15/Component_Function_4/NAND4_in[0] ,
         \SB1_0_16/Component_Function_2/NAND4_in[3] ,
         \SB1_0_16/Component_Function_2/NAND4_in[1] ,
         \SB1_0_16/Component_Function_3/NAND4_in[3] ,
         \SB1_0_16/Component_Function_3/NAND4_in[2] ,
         \SB1_0_16/Component_Function_3/NAND4_in[1] ,
         \SB1_0_16/Component_Function_3/NAND4_in[0] ,
         \SB1_0_16/Component_Function_4/NAND4_in[3] ,
         \SB1_0_16/Component_Function_4/NAND4_in[1] ,
         \SB1_0_16/Component_Function_4/NAND4_in[0] ,
         \SB1_0_17/Component_Function_2/NAND4_in[2] ,
         \SB1_0_17/Component_Function_3/NAND4_in[3] ,
         \SB1_0_17/Component_Function_3/NAND4_in[1] ,
         \SB1_0_17/Component_Function_3/NAND4_in[0] ,
         \SB1_0_17/Component_Function_4/NAND4_in[3] ,
         \SB1_0_17/Component_Function_4/NAND4_in[1] ,
         \SB1_0_17/Component_Function_4/NAND4_in[0] ,
         \SB1_0_18/Component_Function_2/NAND4_in[2] ,
         \SB1_0_18/Component_Function_2/NAND4_in[1] ,
         \SB1_0_18/Component_Function_2/NAND4_in[0] ,
         \SB1_0_18/Component_Function_3/NAND4_in[3] ,
         \SB1_0_18/Component_Function_3/NAND4_in[1] ,
         \SB1_0_18/Component_Function_3/NAND4_in[0] ,
         \SB1_0_18/Component_Function_4/NAND4_in[3] ,
         \SB1_0_18/Component_Function_4/NAND4_in[2] ,
         \SB1_0_18/Component_Function_4/NAND4_in[1] ,
         \SB1_0_19/Component_Function_2/NAND4_in[2] ,
         \SB1_0_19/Component_Function_2/NAND4_in[0] ,
         \SB1_0_19/Component_Function_3/NAND4_in[3] ,
         \SB1_0_19/Component_Function_3/NAND4_in[2] ,
         \SB1_0_19/Component_Function_3/NAND4_in[1] ,
         \SB1_0_19/Component_Function_4/NAND4_in[1] ,
         \SB1_0_19/Component_Function_4/NAND4_in[0] ,
         \SB1_0_20/Component_Function_2/NAND4_in[3] ,
         \SB1_0_20/Component_Function_2/NAND4_in[2] ,
         \SB1_0_20/Component_Function_2/NAND4_in[1] ,
         \SB1_0_20/Component_Function_2/NAND4_in[0] ,
         \SB1_0_20/Component_Function_3/NAND4_in[3] ,
         \SB1_0_20/Component_Function_3/NAND4_in[2] ,
         \SB1_0_20/Component_Function_3/NAND4_in[1] ,
         \SB1_0_20/Component_Function_4/NAND4_in[3] ,
         \SB1_0_20/Component_Function_4/NAND4_in[1] ,
         \SB1_0_20/Component_Function_4/NAND4_in[0] ,
         \SB1_0_21/Component_Function_2/NAND4_in[2] ,
         \SB1_0_21/Component_Function_2/NAND4_in[1] ,
         \SB1_0_21/Component_Function_3/NAND4_in[3] ,
         \SB1_0_21/Component_Function_3/NAND4_in[2] ,
         \SB1_0_21/Component_Function_3/NAND4_in[1] ,
         \SB1_0_21/Component_Function_3/NAND4_in[0] ,
         \SB1_0_21/Component_Function_4/NAND4_in[3] ,
         \SB1_0_21/Component_Function_4/NAND4_in[1] ,
         \SB1_0_22/Component_Function_2/NAND4_in[3] ,
         \SB1_0_22/Component_Function_2/NAND4_in[2] ,
         \SB1_0_22/Component_Function_2/NAND4_in[1] ,
         \SB1_0_22/Component_Function_2/NAND4_in[0] ,
         \SB1_0_22/Component_Function_3/NAND4_in[3] ,
         \SB1_0_22/Component_Function_3/NAND4_in[2] ,
         \SB1_0_22/Component_Function_3/NAND4_in[1] ,
         \SB1_0_22/Component_Function_3/NAND4_in[0] ,
         \SB1_0_22/Component_Function_4/NAND4_in[3] ,
         \SB1_0_22/Component_Function_4/NAND4_in[2] ,
         \SB1_0_22/Component_Function_4/NAND4_in[1] ,
         \SB1_0_22/Component_Function_4/NAND4_in[0] ,
         \SB1_0_23/Component_Function_2/NAND4_in[3] ,
         \SB1_0_23/Component_Function_2/NAND4_in[2] ,
         \SB1_0_23/Component_Function_2/NAND4_in[1] ,
         \SB1_0_23/Component_Function_2/NAND4_in[0] ,
         \SB1_0_23/Component_Function_3/NAND4_in[3] ,
         \SB1_0_23/Component_Function_3/NAND4_in[2] ,
         \SB1_0_23/Component_Function_3/NAND4_in[1] ,
         \SB1_0_23/Component_Function_3/NAND4_in[0] ,
         \SB1_0_23/Component_Function_4/NAND4_in[3] ,
         \SB1_0_23/Component_Function_4/NAND4_in[2] ,
         \SB1_0_23/Component_Function_4/NAND4_in[1] ,
         \SB1_0_23/Component_Function_4/NAND4_in[0] ,
         \SB1_0_24/Component_Function_2/NAND4_in[1] ,
         \SB1_0_24/Component_Function_3/NAND4_in[2] ,
         \SB1_0_24/Component_Function_3/NAND4_in[1] ,
         \SB1_0_24/Component_Function_3/NAND4_in[0] ,
         \SB1_0_24/Component_Function_4/NAND4_in[2] ,
         \SB1_0_24/Component_Function_4/NAND4_in[1] ,
         \SB1_0_24/Component_Function_4/NAND4_in[0] ,
         \SB1_0_25/Component_Function_2/NAND4_in[3] ,
         \SB1_0_25/Component_Function_2/NAND4_in[0] ,
         \SB1_0_25/Component_Function_3/NAND4_in[3] ,
         \SB1_0_25/Component_Function_3/NAND4_in[1] ,
         \SB1_0_25/Component_Function_3/NAND4_in[0] ,
         \SB1_0_25/Component_Function_4/NAND4_in[3] ,
         \SB1_0_25/Component_Function_4/NAND4_in[1] ,
         \SB1_0_25/Component_Function_4/NAND4_in[0] ,
         \SB1_0_26/Component_Function_2/NAND4_in[3] ,
         \SB1_0_26/Component_Function_2/NAND4_in[1] ,
         \SB1_0_26/Component_Function_2/NAND4_in[0] ,
         \SB1_0_26/Component_Function_3/NAND4_in[2] ,
         \SB1_0_26/Component_Function_3/NAND4_in[1] ,
         \SB1_0_26/Component_Function_3/NAND4_in[0] ,
         \SB1_0_26/Component_Function_4/NAND4_in[3] ,
         \SB1_0_26/Component_Function_4/NAND4_in[2] ,
         \SB1_0_26/Component_Function_4/NAND4_in[1] ,
         \SB1_0_27/Component_Function_2/NAND4_in[3] ,
         \SB1_0_27/Component_Function_2/NAND4_in[1] ,
         \SB1_0_27/Component_Function_2/NAND4_in[0] ,
         \SB1_0_27/Component_Function_3/NAND4_in[3] ,
         \SB1_0_27/Component_Function_3/NAND4_in[2] ,
         \SB1_0_27/Component_Function_3/NAND4_in[1] ,
         \SB1_0_27/Component_Function_3/NAND4_in[0] ,
         \SB1_0_27/Component_Function_4/NAND4_in[3] ,
         \SB1_0_27/Component_Function_4/NAND4_in[2] ,
         \SB1_0_27/Component_Function_4/NAND4_in[1] ,
         \SB1_0_28/Component_Function_2/NAND4_in[3] ,
         \SB1_0_28/Component_Function_2/NAND4_in[2] ,
         \SB1_0_28/Component_Function_2/NAND4_in[1] ,
         \SB1_0_28/Component_Function_2/NAND4_in[0] ,
         \SB1_0_28/Component_Function_3/NAND4_in[3] ,
         \SB1_0_28/Component_Function_3/NAND4_in[1] ,
         \SB1_0_28/Component_Function_3/NAND4_in[0] ,
         \SB1_0_28/Component_Function_4/NAND4_in[2] ,
         \SB1_0_28/Component_Function_4/NAND4_in[1] ,
         \SB1_0_28/Component_Function_4/NAND4_in[0] ,
         \SB1_0_29/Component_Function_2/NAND4_in[2] ,
         \SB1_0_29/Component_Function_2/NAND4_in[0] ,
         \SB1_0_29/Component_Function_3/NAND4_in[3] ,
         \SB1_0_29/Component_Function_3/NAND4_in[2] ,
         \SB1_0_29/Component_Function_3/NAND4_in[1] ,
         \SB1_0_29/Component_Function_3/NAND4_in[0] ,
         \SB1_0_29/Component_Function_4/NAND4_in[2] ,
         \SB1_0_29/Component_Function_4/NAND4_in[1] ,
         \SB1_0_29/Component_Function_4/NAND4_in[0] ,
         \SB1_0_30/Component_Function_2/NAND4_in[2] ,
         \SB1_0_30/Component_Function_2/NAND4_in[0] ,
         \SB1_0_30/Component_Function_3/NAND4_in[3] ,
         \SB1_0_30/Component_Function_3/NAND4_in[2] ,
         \SB1_0_30/Component_Function_4/NAND4_in[3] ,
         \SB1_0_30/Component_Function_4/NAND4_in[2] ,
         \SB1_0_30/Component_Function_4/NAND4_in[0] ,
         \SB1_0_31/Component_Function_2/NAND4_in[3] ,
         \SB1_0_31/Component_Function_2/NAND4_in[2] ,
         \SB1_0_31/Component_Function_2/NAND4_in[1] ,
         \SB1_0_31/Component_Function_2/NAND4_in[0] ,
         \SB1_0_31/Component_Function_3/NAND4_in[3] ,
         \SB1_0_31/Component_Function_3/NAND4_in[1] ,
         \SB1_0_31/Component_Function_4/NAND4_in[3] ,
         \SB1_0_31/Component_Function_4/NAND4_in[1] ,
         \SB1_0_31/Component_Function_4/NAND4_in[0] ,
         \SB2_0_0/Component_Function_2/NAND4_in[3] ,
         \SB2_0_0/Component_Function_2/NAND4_in[2] ,
         \SB2_0_0/Component_Function_2/NAND4_in[0] ,
         \SB2_0_0/Component_Function_3/NAND4_in[2] ,
         \SB2_0_0/Component_Function_3/NAND4_in[1] ,
         \SB2_0_0/Component_Function_3/NAND4_in[0] ,
         \SB2_0_0/Component_Function_4/NAND4_in[3] ,
         \SB2_0_0/Component_Function_4/NAND4_in[1] ,
         \SB2_0_0/Component_Function_4/NAND4_in[0] ,
         \SB2_0_1/Component_Function_2/NAND4_in[1] ,
         \SB2_0_1/Component_Function_2/NAND4_in[0] ,
         \SB2_0_1/Component_Function_3/NAND4_in[2] ,
         \SB2_0_1/Component_Function_3/NAND4_in[1] ,
         \SB2_0_1/Component_Function_3/NAND4_in[0] ,
         \SB2_0_1/Component_Function_4/NAND4_in[3] ,
         \SB2_0_1/Component_Function_4/NAND4_in[2] ,
         \SB2_0_1/Component_Function_4/NAND4_in[1] ,
         \SB2_0_1/Component_Function_4/NAND4_in[0] ,
         \SB2_0_2/Component_Function_2/NAND4_in[2] ,
         \SB2_0_2/Component_Function_2/NAND4_in[1] ,
         \SB2_0_2/Component_Function_2/NAND4_in[0] ,
         \SB2_0_2/Component_Function_3/NAND4_in[3] ,
         \SB2_0_2/Component_Function_3/NAND4_in[2] ,
         \SB2_0_2/Component_Function_3/NAND4_in[1] ,
         \SB2_0_2/Component_Function_3/NAND4_in[0] ,
         \SB2_0_2/Component_Function_4/NAND4_in[3] ,
         \SB2_0_2/Component_Function_4/NAND4_in[2] ,
         \SB2_0_2/Component_Function_4/NAND4_in[1] ,
         \SB2_0_2/Component_Function_4/NAND4_in[0] ,
         \SB2_0_3/Component_Function_2/NAND4_in[2] ,
         \SB2_0_3/Component_Function_2/NAND4_in[1] ,
         \SB2_0_3/Component_Function_2/NAND4_in[0] ,
         \SB2_0_3/Component_Function_3/NAND4_in[3] ,
         \SB2_0_3/Component_Function_3/NAND4_in[0] ,
         \SB2_0_3/Component_Function_4/NAND4_in[3] ,
         \SB2_0_3/Component_Function_4/NAND4_in[1] ,
         \SB2_0_3/Component_Function_4/NAND4_in[0] ,
         \SB2_0_4/Component_Function_2/NAND4_in[2] ,
         \SB2_0_4/Component_Function_2/NAND4_in[0] ,
         \SB2_0_4/Component_Function_3/NAND4_in[2] ,
         \SB2_0_4/Component_Function_3/NAND4_in[0] ,
         \SB2_0_4/Component_Function_4/NAND4_in[1] ,
         \SB2_0_5/Component_Function_2/NAND4_in[3] ,
         \SB2_0_5/Component_Function_2/NAND4_in[1] ,
         \SB2_0_5/Component_Function_2/NAND4_in[0] ,
         \SB2_0_5/Component_Function_3/NAND4_in[3] ,
         \SB2_0_5/Component_Function_3/NAND4_in[2] ,
         \SB2_0_5/Component_Function_3/NAND4_in[1] ,
         \SB2_0_5/Component_Function_3/NAND4_in[0] ,
         \SB2_0_5/Component_Function_4/NAND4_in[3] ,
         \SB2_0_5/Component_Function_4/NAND4_in[1] ,
         \SB2_0_5/Component_Function_4/NAND4_in[0] ,
         \SB2_0_6/Component_Function_2/NAND4_in[3] ,
         \SB2_0_6/Component_Function_2/NAND4_in[2] ,
         \SB2_0_6/Component_Function_2/NAND4_in[1] ,
         \SB2_0_6/Component_Function_2/NAND4_in[0] ,
         \SB2_0_6/Component_Function_3/NAND4_in[3] ,
         \SB2_0_6/Component_Function_3/NAND4_in[2] ,
         \SB2_0_6/Component_Function_3/NAND4_in[1] ,
         \SB2_0_6/Component_Function_3/NAND4_in[0] ,
         \SB2_0_6/Component_Function_4/NAND4_in[2] ,
         \SB2_0_6/Component_Function_4/NAND4_in[1] ,
         \SB2_0_6/Component_Function_4/NAND4_in[0] ,
         \SB2_0_7/Component_Function_2/NAND4_in[2] ,
         \SB2_0_7/Component_Function_2/NAND4_in[1] ,
         \SB2_0_7/Component_Function_3/NAND4_in[3] ,
         \SB2_0_7/Component_Function_3/NAND4_in[2] ,
         \SB2_0_7/Component_Function_3/NAND4_in[1] ,
         \SB2_0_7/Component_Function_3/NAND4_in[0] ,
         \SB2_0_7/Component_Function_4/NAND4_in[3] ,
         \SB2_0_7/Component_Function_4/NAND4_in[2] ,
         \SB2_0_7/Component_Function_4/NAND4_in[1] ,
         \SB2_0_7/Component_Function_4/NAND4_in[0] ,
         \SB2_0_8/Component_Function_2/NAND4_in[3] ,
         \SB2_0_8/Component_Function_2/NAND4_in[2] ,
         \SB2_0_8/Component_Function_2/NAND4_in[1] ,
         \SB2_0_8/Component_Function_2/NAND4_in[0] ,
         \SB2_0_8/Component_Function_3/NAND4_in[2] ,
         \SB2_0_8/Component_Function_3/NAND4_in[1] ,
         \SB2_0_8/Component_Function_3/NAND4_in[0] ,
         \SB2_0_8/Component_Function_4/NAND4_in[3] ,
         \SB2_0_8/Component_Function_4/NAND4_in[2] ,
         \SB2_0_8/Component_Function_4/NAND4_in[1] ,
         \SB2_0_9/Component_Function_2/NAND4_in[3] ,
         \SB2_0_9/Component_Function_2/NAND4_in[1] ,
         \SB2_0_9/Component_Function_2/NAND4_in[0] ,
         \SB2_0_9/Component_Function_3/NAND4_in[3] ,
         \SB2_0_9/Component_Function_3/NAND4_in[1] ,
         \SB2_0_9/Component_Function_3/NAND4_in[0] ,
         \SB2_0_9/Component_Function_4/NAND4_in[3] ,
         \SB2_0_9/Component_Function_4/NAND4_in[1] ,
         \SB2_0_9/Component_Function_4/NAND4_in[0] ,
         \SB2_0_10/Component_Function_2/NAND4_in[3] ,
         \SB2_0_10/Component_Function_2/NAND4_in[2] ,
         \SB2_0_10/Component_Function_2/NAND4_in[0] ,
         \SB2_0_10/Component_Function_3/NAND4_in[3] ,
         \SB2_0_10/Component_Function_3/NAND4_in[2] ,
         \SB2_0_10/Component_Function_3/NAND4_in[1] ,
         \SB2_0_10/Component_Function_3/NAND4_in[0] ,
         \SB2_0_10/Component_Function_4/NAND4_in[2] ,
         \SB2_0_10/Component_Function_4/NAND4_in[1] ,
         \SB2_0_10/Component_Function_4/NAND4_in[0] ,
         \SB2_0_11/Component_Function_2/NAND4_in[3] ,
         \SB2_0_11/Component_Function_2/NAND4_in[2] ,
         \SB2_0_11/Component_Function_2/NAND4_in[0] ,
         \SB2_0_11/Component_Function_3/NAND4_in[3] ,
         \SB2_0_11/Component_Function_3/NAND4_in[1] ,
         \SB2_0_11/Component_Function_3/NAND4_in[0] ,
         \SB2_0_11/Component_Function_4/NAND4_in[3] ,
         \SB2_0_11/Component_Function_4/NAND4_in[0] ,
         \SB2_0_12/Component_Function_2/NAND4_in[2] ,
         \SB2_0_12/Component_Function_3/NAND4_in[3] ,
         \SB2_0_12/Component_Function_3/NAND4_in[2] ,
         \SB2_0_12/Component_Function_3/NAND4_in[1] ,
         \SB2_0_12/Component_Function_3/NAND4_in[0] ,
         \SB2_0_12/Component_Function_4/NAND4_in[2] ,
         \SB2_0_12/Component_Function_4/NAND4_in[1] ,
         \SB2_0_12/Component_Function_4/NAND4_in[0] ,
         \SB2_0_13/Component_Function_2/NAND4_in[3] ,
         \SB2_0_13/Component_Function_2/NAND4_in[2] ,
         \SB2_0_13/Component_Function_2/NAND4_in[1] ,
         \SB2_0_13/Component_Function_2/NAND4_in[0] ,
         \SB2_0_13/Component_Function_3/NAND4_in[2] ,
         \SB2_0_13/Component_Function_3/NAND4_in[0] ,
         \SB2_0_13/Component_Function_4/NAND4_in[3] ,
         \SB2_0_13/Component_Function_4/NAND4_in[1] ,
         \SB2_0_13/Component_Function_4/NAND4_in[0] ,
         \SB2_0_14/Component_Function_2/NAND4_in[2] ,
         \SB2_0_14/Component_Function_2/NAND4_in[1] ,
         \SB2_0_14/Component_Function_2/NAND4_in[0] ,
         \SB2_0_14/Component_Function_3/NAND4_in[3] ,
         \SB2_0_14/Component_Function_3/NAND4_in[1] ,
         \SB2_0_14/Component_Function_3/NAND4_in[0] ,
         \SB2_0_14/Component_Function_4/NAND4_in[3] ,
         \SB2_0_14/Component_Function_4/NAND4_in[1] ,
         \SB2_0_14/Component_Function_4/NAND4_in[0] ,
         \SB2_0_15/Component_Function_2/NAND4_in[3] ,
         \SB2_0_15/Component_Function_2/NAND4_in[1] ,
         \SB2_0_15/Component_Function_2/NAND4_in[0] ,
         \SB2_0_15/Component_Function_3/NAND4_in[3] ,
         \SB2_0_15/Component_Function_3/NAND4_in[2] ,
         \SB2_0_15/Component_Function_4/NAND4_in[3] ,
         \SB2_0_15/Component_Function_4/NAND4_in[1] ,
         \SB2_0_15/Component_Function_4/NAND4_in[0] ,
         \SB2_0_16/Component_Function_2/NAND4_in[0] ,
         \SB2_0_16/Component_Function_3/NAND4_in[3] ,
         \SB2_0_16/Component_Function_3/NAND4_in[2] ,
         \SB2_0_16/Component_Function_3/NAND4_in[0] ,
         \SB2_0_16/Component_Function_4/NAND4_in[3] ,
         \SB2_0_16/Component_Function_4/NAND4_in[1] ,
         \SB2_0_16/Component_Function_4/NAND4_in[0] ,
         \SB2_0_17/Component_Function_2/NAND4_in[2] ,
         \SB2_0_17/Component_Function_2/NAND4_in[0] ,
         \SB2_0_17/Component_Function_3/NAND4_in[3] ,
         \SB2_0_17/Component_Function_3/NAND4_in[0] ,
         \SB2_0_17/Component_Function_4/NAND4_in[3] ,
         \SB2_0_17/Component_Function_4/NAND4_in[2] ,
         \SB2_0_17/Component_Function_4/NAND4_in[1] ,
         \SB2_0_17/Component_Function_4/NAND4_in[0] ,
         \SB2_0_18/Component_Function_2/NAND4_in[0] ,
         \SB2_0_18/Component_Function_3/NAND4_in[3] ,
         \SB2_0_18/Component_Function_3/NAND4_in[1] ,
         \SB2_0_18/Component_Function_3/NAND4_in[0] ,
         \SB2_0_18/Component_Function_4/NAND4_in[3] ,
         \SB2_0_18/Component_Function_4/NAND4_in[1] ,
         \SB2_0_18/Component_Function_4/NAND4_in[0] ,
         \SB2_0_19/Component_Function_2/NAND4_in[3] ,
         \SB2_0_19/Component_Function_2/NAND4_in[2] ,
         \SB2_0_19/Component_Function_2/NAND4_in[1] ,
         \SB2_0_19/Component_Function_2/NAND4_in[0] ,
         \SB2_0_19/Component_Function_3/NAND4_in[3] ,
         \SB2_0_19/Component_Function_3/NAND4_in[2] ,
         \SB2_0_19/Component_Function_3/NAND4_in[1] ,
         \SB2_0_19/Component_Function_3/NAND4_in[0] ,
         \SB2_0_19/Component_Function_4/NAND4_in[3] ,
         \SB2_0_19/Component_Function_4/NAND4_in[0] ,
         \SB2_0_20/Component_Function_2/NAND4_in[3] ,
         \SB2_0_20/Component_Function_2/NAND4_in[2] ,
         \SB2_0_20/Component_Function_2/NAND4_in[1] ,
         \SB2_0_20/Component_Function_2/NAND4_in[0] ,
         \SB2_0_20/Component_Function_3/NAND4_in[3] ,
         \SB2_0_20/Component_Function_3/NAND4_in[2] ,
         \SB2_0_20/Component_Function_3/NAND4_in[1] ,
         \SB2_0_20/Component_Function_3/NAND4_in[0] ,
         \SB2_0_20/Component_Function_4/NAND4_in[3] ,
         \SB2_0_20/Component_Function_4/NAND4_in[2] ,
         \SB2_0_20/Component_Function_4/NAND4_in[1] ,
         \SB2_0_20/Component_Function_4/NAND4_in[0] ,
         \SB2_0_21/Component_Function_2/NAND4_in[2] ,
         \SB2_0_21/Component_Function_2/NAND4_in[1] ,
         \SB2_0_21/Component_Function_2/NAND4_in[0] ,
         \SB2_0_21/Component_Function_3/NAND4_in[3] ,
         \SB2_0_21/Component_Function_3/NAND4_in[1] ,
         \SB2_0_21/Component_Function_3/NAND4_in[0] ,
         \SB2_0_21/Component_Function_4/NAND4_in[3] ,
         \SB2_0_21/Component_Function_4/NAND4_in[1] ,
         \SB2_0_21/Component_Function_4/NAND4_in[0] ,
         \SB2_0_22/Component_Function_2/NAND4_in[3] ,
         \SB2_0_22/Component_Function_2/NAND4_in[2] ,
         \SB2_0_22/Component_Function_2/NAND4_in[1] ,
         \SB2_0_22/Component_Function_2/NAND4_in[0] ,
         \SB2_0_22/Component_Function_3/NAND4_in[3] ,
         \SB2_0_22/Component_Function_3/NAND4_in[1] ,
         \SB2_0_22/Component_Function_4/NAND4_in[3] ,
         \SB2_0_22/Component_Function_4/NAND4_in[1] ,
         \SB2_0_22/Component_Function_4/NAND4_in[0] ,
         \SB2_0_23/Component_Function_2/NAND4_in[3] ,
         \SB2_0_23/Component_Function_2/NAND4_in[2] ,
         \SB2_0_23/Component_Function_2/NAND4_in[1] ,
         \SB2_0_23/Component_Function_3/NAND4_in[2] ,
         \SB2_0_23/Component_Function_3/NAND4_in[1] ,
         \SB2_0_23/Component_Function_3/NAND4_in[0] ,
         \SB2_0_23/Component_Function_4/NAND4_in[3] ,
         \SB2_0_23/Component_Function_4/NAND4_in[1] ,
         \SB2_0_23/Component_Function_4/NAND4_in[0] ,
         \SB2_0_24/Component_Function_2/NAND4_in[3] ,
         \SB2_0_24/Component_Function_2/NAND4_in[2] ,
         \SB2_0_24/Component_Function_2/NAND4_in[0] ,
         \SB2_0_24/Component_Function_3/NAND4_in[3] ,
         \SB2_0_24/Component_Function_3/NAND4_in[2] ,
         \SB2_0_24/Component_Function_3/NAND4_in[0] ,
         \SB2_0_24/Component_Function_4/NAND4_in[3] ,
         \SB2_0_24/Component_Function_4/NAND4_in[2] ,
         \SB2_0_24/Component_Function_4/NAND4_in[1] ,
         \SB2_0_24/Component_Function_4/NAND4_in[0] ,
         \SB2_0_25/Component_Function_2/NAND4_in[3] ,
         \SB2_0_25/Component_Function_2/NAND4_in[2] ,
         \SB2_0_25/Component_Function_2/NAND4_in[1] ,
         \SB2_0_25/Component_Function_2/NAND4_in[0] ,
         \SB2_0_25/Component_Function_3/NAND4_in[3] ,
         \SB2_0_25/Component_Function_3/NAND4_in[2] ,
         \SB2_0_25/Component_Function_3/NAND4_in[1] ,
         \SB2_0_25/Component_Function_3/NAND4_in[0] ,
         \SB2_0_25/Component_Function_4/NAND4_in[3] ,
         \SB2_0_25/Component_Function_4/NAND4_in[2] ,
         \SB2_0_25/Component_Function_4/NAND4_in[0] ,
         \SB2_0_26/Component_Function_2/NAND4_in[3] ,
         \SB2_0_26/Component_Function_2/NAND4_in[2] ,
         \SB2_0_26/Component_Function_2/NAND4_in[1] ,
         \SB2_0_26/Component_Function_2/NAND4_in[0] ,
         \SB2_0_26/Component_Function_3/NAND4_in[3] ,
         \SB2_0_26/Component_Function_3/NAND4_in[2] ,
         \SB2_0_26/Component_Function_3/NAND4_in[1] ,
         \SB2_0_26/Component_Function_3/NAND4_in[0] ,
         \SB2_0_26/Component_Function_4/NAND4_in[3] ,
         \SB2_0_26/Component_Function_4/NAND4_in[2] ,
         \SB2_0_26/Component_Function_4/NAND4_in[1] ,
         \SB2_0_26/Component_Function_4/NAND4_in[0] ,
         \SB2_0_27/Component_Function_2/NAND4_in[2] ,
         \SB2_0_27/Component_Function_2/NAND4_in[1] ,
         \SB2_0_27/Component_Function_2/NAND4_in[0] ,
         \SB2_0_27/Component_Function_3/NAND4_in[3] ,
         \SB2_0_27/Component_Function_3/NAND4_in[2] ,
         \SB2_0_27/Component_Function_3/NAND4_in[1] ,
         \SB2_0_27/Component_Function_3/NAND4_in[0] ,
         \SB2_0_27/Component_Function_4/NAND4_in[3] ,
         \SB2_0_27/Component_Function_4/NAND4_in[2] ,
         \SB2_0_27/Component_Function_4/NAND4_in[1] ,
         \SB2_0_27/Component_Function_4/NAND4_in[0] ,
         \SB2_0_28/Component_Function_2/NAND4_in[3] ,
         \SB2_0_28/Component_Function_2/NAND4_in[2] ,
         \SB2_0_28/Component_Function_2/NAND4_in[1] ,
         \SB2_0_28/Component_Function_2/NAND4_in[0] ,
         \SB2_0_28/Component_Function_3/NAND4_in[3] ,
         \SB2_0_28/Component_Function_3/NAND4_in[1] ,
         \SB2_0_28/Component_Function_3/NAND4_in[0] ,
         \SB2_0_28/Component_Function_4/NAND4_in[3] ,
         \SB2_0_28/Component_Function_4/NAND4_in[1] ,
         \SB2_0_28/Component_Function_4/NAND4_in[0] ,
         \SB2_0_29/Component_Function_2/NAND4_in[3] ,
         \SB2_0_29/Component_Function_2/NAND4_in[1] ,
         \SB2_0_29/Component_Function_2/NAND4_in[0] ,
         \SB2_0_29/Component_Function_3/NAND4_in[3] ,
         \SB2_0_29/Component_Function_3/NAND4_in[2] ,
         \SB2_0_29/Component_Function_3/NAND4_in[1] ,
         \SB2_0_29/Component_Function_4/NAND4_in[3] ,
         \SB2_0_29/Component_Function_4/NAND4_in[2] ,
         \SB2_0_29/Component_Function_4/NAND4_in[1] ,
         \SB2_0_29/Component_Function_4/NAND4_in[0] ,
         \SB2_0_30/Component_Function_2/NAND4_in[3] ,
         \SB2_0_30/Component_Function_2/NAND4_in[1] ,
         \SB2_0_30/Component_Function_2/NAND4_in[0] ,
         \SB2_0_30/Component_Function_3/NAND4_in[3] ,
         \SB2_0_30/Component_Function_3/NAND4_in[2] ,
         \SB2_0_30/Component_Function_3/NAND4_in[1] ,
         \SB2_0_30/Component_Function_3/NAND4_in[0] ,
         \SB2_0_30/Component_Function_4/NAND4_in[3] ,
         \SB2_0_30/Component_Function_4/NAND4_in[1] ,
         \SB2_0_30/Component_Function_4/NAND4_in[0] ,
         \SB2_0_31/Component_Function_2/NAND4_in[3] ,
         \SB2_0_31/Component_Function_2/NAND4_in[2] ,
         \SB2_0_31/Component_Function_2/NAND4_in[1] ,
         \SB2_0_31/Component_Function_2/NAND4_in[0] ,
         \SB2_0_31/Component_Function_3/NAND4_in[2] ,
         \SB2_0_31/Component_Function_3/NAND4_in[1] ,
         \SB2_0_31/Component_Function_3/NAND4_in[0] ,
         \SB2_0_31/Component_Function_4/NAND4_in[2] ,
         \SB2_0_31/Component_Function_4/NAND4_in[1] ,
         \SB2_0_31/Component_Function_4/NAND4_in[0] ,
         \SB1_1_0/Component_Function_2/NAND4_in[3] ,
         \SB1_1_0/Component_Function_2/NAND4_in[1] ,
         \SB1_1_0/Component_Function_3/NAND4_in[1] ,
         \SB1_1_0/Component_Function_3/NAND4_in[0] ,
         \SB1_1_0/Component_Function_4/NAND4_in[3] ,
         \SB1_1_0/Component_Function_4/NAND4_in[2] ,
         \SB1_1_1/Component_Function_2/NAND4_in[3] ,
         \SB1_1_1/Component_Function_2/NAND4_in[2] ,
         \SB1_1_1/Component_Function_2/NAND4_in[0] ,
         \SB1_1_1/Component_Function_3/NAND4_in[2] ,
         \SB1_1_1/Component_Function_3/NAND4_in[1] ,
         \SB1_1_1/Component_Function_4/NAND4_in[3] ,
         \SB1_1_1/Component_Function_4/NAND4_in[1] ,
         \SB1_1_1/Component_Function_4/NAND4_in[0] ,
         \SB1_1_2/Component_Function_2/NAND4_in[3] ,
         \SB1_1_2/Component_Function_2/NAND4_in[2] ,
         \SB1_1_2/Component_Function_2/NAND4_in[1] ,
         \SB1_1_2/Component_Function_2/NAND4_in[0] ,
         \SB1_1_2/Component_Function_3/NAND4_in[3] ,
         \SB1_1_2/Component_Function_3/NAND4_in[1] ,
         \SB1_1_2/Component_Function_3/NAND4_in[0] ,
         \SB1_1_2/Component_Function_4/NAND4_in[2] ,
         \SB1_1_2/Component_Function_4/NAND4_in[1] ,
         \SB1_1_2/Component_Function_4/NAND4_in[0] ,
         \SB1_1_3/Component_Function_2/NAND4_in[1] ,
         \SB1_1_3/Component_Function_2/NAND4_in[0] ,
         \SB1_1_3/Component_Function_3/NAND4_in[1] ,
         \SB1_1_3/Component_Function_3/NAND4_in[0] ,
         \SB1_1_3/Component_Function_4/NAND4_in[2] ,
         \SB1_1_3/Component_Function_4/NAND4_in[1] ,
         \SB1_1_4/Component_Function_2/NAND4_in[2] ,
         \SB1_1_4/Component_Function_2/NAND4_in[1] ,
         \SB1_1_4/Component_Function_3/NAND4_in[1] ,
         \SB1_1_4/Component_Function_3/NAND4_in[0] ,
         \SB1_1_4/Component_Function_4/NAND4_in[2] ,
         \SB1_1_4/Component_Function_4/NAND4_in[1] ,
         \SB1_1_5/Component_Function_2/NAND4_in[3] ,
         \SB1_1_5/Component_Function_2/NAND4_in[2] ,
         \SB1_1_5/Component_Function_2/NAND4_in[1] ,
         \SB1_1_5/Component_Function_3/NAND4_in[2] ,
         \SB1_1_5/Component_Function_3/NAND4_in[1] ,
         \SB1_1_5/Component_Function_3/NAND4_in[0] ,
         \SB1_1_5/Component_Function_4/NAND4_in[3] ,
         \SB1_1_5/Component_Function_4/NAND4_in[2] ,
         \SB1_1_5/Component_Function_4/NAND4_in[1] ,
         \SB1_1_5/Component_Function_4/NAND4_in[0] ,
         \SB1_1_6/Component_Function_2/NAND4_in[1] ,
         \SB1_1_6/Component_Function_3/NAND4_in[2] ,
         \SB1_1_6/Component_Function_3/NAND4_in[0] ,
         \SB1_1_6/Component_Function_4/NAND4_in[3] ,
         \SB1_1_6/Component_Function_4/NAND4_in[1] ,
         \SB1_1_6/Component_Function_4/NAND4_in[0] ,
         \SB1_1_7/Component_Function_2/NAND4_in[2] ,
         \SB1_1_7/Component_Function_2/NAND4_in[1] ,
         \SB1_1_7/Component_Function_2/NAND4_in[0] ,
         \SB1_1_7/Component_Function_3/NAND4_in[3] ,
         \SB1_1_7/Component_Function_3/NAND4_in[2] ,
         \SB1_1_7/Component_Function_3/NAND4_in[1] ,
         \SB1_1_7/Component_Function_4/NAND4_in[3] ,
         \SB1_1_7/Component_Function_4/NAND4_in[1] ,
         \SB1_1_7/Component_Function_4/NAND4_in[0] ,
         \SB1_1_8/Component_Function_2/NAND4_in[2] ,
         \SB1_1_8/Component_Function_2/NAND4_in[1] ,
         \SB1_1_8/Component_Function_2/NAND4_in[0] ,
         \SB1_1_8/Component_Function_3/NAND4_in[1] ,
         \SB1_1_8/Component_Function_3/NAND4_in[0] ,
         \SB1_1_8/Component_Function_4/NAND4_in[3] ,
         \SB1_1_8/Component_Function_4/NAND4_in[1] ,
         \SB1_1_8/Component_Function_4/NAND4_in[0] ,
         \SB1_1_9/Component_Function_2/NAND4_in[2] ,
         \SB1_1_9/Component_Function_2/NAND4_in[1] ,
         \SB1_1_9/Component_Function_3/NAND4_in[2] ,
         \SB1_1_9/Component_Function_3/NAND4_in[1] ,
         \SB1_1_9/Component_Function_3/NAND4_in[0] ,
         \SB1_1_9/Component_Function_4/NAND4_in[2] ,
         \SB1_1_9/Component_Function_4/NAND4_in[1] ,
         \SB1_1_9/Component_Function_4/NAND4_in[0] ,
         \SB1_1_10/Component_Function_2/NAND4_in[1] ,
         \SB1_1_10/Component_Function_2/NAND4_in[0] ,
         \SB1_1_10/Component_Function_3/NAND4_in[2] ,
         \SB1_1_10/Component_Function_3/NAND4_in[1] ,
         \SB1_1_10/Component_Function_4/NAND4_in[3] ,
         \SB1_1_10/Component_Function_4/NAND4_in[2] ,
         \SB1_1_10/Component_Function_4/NAND4_in[1] ,
         \SB1_1_10/Component_Function_4/NAND4_in[0] ,
         \SB1_1_11/Component_Function_2/NAND4_in[1] ,
         \SB1_1_11/Component_Function_2/NAND4_in[0] ,
         \SB1_1_11/Component_Function_3/NAND4_in[2] ,
         \SB1_1_11/Component_Function_3/NAND4_in[1] ,
         \SB1_1_11/Component_Function_3/NAND4_in[0] ,
         \SB1_1_11/Component_Function_4/NAND4_in[3] ,
         \SB1_1_11/Component_Function_4/NAND4_in[2] ,
         \SB1_1_11/Component_Function_4/NAND4_in[1] ,
         \SB1_1_11/Component_Function_4/NAND4_in[0] ,
         \SB1_1_12/Component_Function_2/NAND4_in[3] ,
         \SB1_1_12/Component_Function_2/NAND4_in[2] ,
         \SB1_1_12/Component_Function_2/NAND4_in[0] ,
         \SB1_1_12/Component_Function_3/NAND4_in[2] ,
         \SB1_1_12/Component_Function_3/NAND4_in[1] ,
         \SB1_1_12/Component_Function_3/NAND4_in[0] ,
         \SB1_1_12/Component_Function_4/NAND4_in[3] ,
         \SB1_1_12/Component_Function_4/NAND4_in[2] ,
         \SB1_1_12/Component_Function_4/NAND4_in[1] ,
         \SB1_1_12/Component_Function_4/NAND4_in[0] ,
         \SB1_1_13/Component_Function_2/NAND4_in[3] ,
         \SB1_1_13/Component_Function_2/NAND4_in[2] ,
         \SB1_1_13/Component_Function_2/NAND4_in[1] ,
         \SB1_1_13/Component_Function_2/NAND4_in[0] ,
         \SB1_1_13/Component_Function_3/NAND4_in[3] ,
         \SB1_1_13/Component_Function_3/NAND4_in[1] ,
         \SB1_1_13/Component_Function_3/NAND4_in[0] ,
         \SB1_1_13/Component_Function_4/NAND4_in[3] ,
         \SB1_1_13/Component_Function_4/NAND4_in[1] ,
         \SB1_1_13/Component_Function_4/NAND4_in[0] ,
         \SB1_1_14/Component_Function_2/NAND4_in[3] ,
         \SB1_1_14/Component_Function_2/NAND4_in[2] ,
         \SB1_1_14/Component_Function_2/NAND4_in[1] ,
         \SB1_1_14/Component_Function_2/NAND4_in[0] ,
         \SB1_1_14/Component_Function_3/NAND4_in[2] ,
         \SB1_1_14/Component_Function_3/NAND4_in[1] ,
         \SB1_1_14/Component_Function_3/NAND4_in[0] ,
         \SB1_1_14/Component_Function_4/NAND4_in[3] ,
         \SB1_1_14/Component_Function_4/NAND4_in[1] ,
         \SB1_1_14/Component_Function_4/NAND4_in[0] ,
         \SB1_1_15/Component_Function_2/NAND4_in[2] ,
         \SB1_1_15/Component_Function_2/NAND4_in[1] ,
         \SB1_1_15/Component_Function_2/NAND4_in[0] ,
         \SB1_1_15/Component_Function_3/NAND4_in[2] ,
         \SB1_1_15/Component_Function_3/NAND4_in[1] ,
         \SB1_1_15/Component_Function_4/NAND4_in[3] ,
         \SB1_1_15/Component_Function_4/NAND4_in[2] ,
         \SB1_1_15/Component_Function_4/NAND4_in[1] ,
         \SB1_1_15/Component_Function_4/NAND4_in[0] ,
         \SB1_1_16/Component_Function_2/NAND4_in[2] ,
         \SB1_1_16/Component_Function_2/NAND4_in[1] ,
         \SB1_1_16/Component_Function_2/NAND4_in[0] ,
         \SB1_1_16/Component_Function_3/NAND4_in[2] ,
         \SB1_1_16/Component_Function_3/NAND4_in[1] ,
         \SB1_1_16/Component_Function_4/NAND4_in[3] ,
         \SB1_1_16/Component_Function_4/NAND4_in[1] ,
         \SB1_1_16/Component_Function_4/NAND4_in[0] ,
         \SB1_1_17/Component_Function_2/NAND4_in[3] ,
         \SB1_1_17/Component_Function_2/NAND4_in[1] ,
         \SB1_1_17/Component_Function_3/NAND4_in[2] ,
         \SB1_1_17/Component_Function_3/NAND4_in[1] ,
         \SB1_1_17/Component_Function_4/NAND4_in[1] ,
         \SB1_1_17/Component_Function_4/NAND4_in[0] ,
         \SB1_1_18/Component_Function_2/NAND4_in[2] ,
         \SB1_1_18/Component_Function_2/NAND4_in[1] ,
         \SB1_1_18/Component_Function_2/NAND4_in[0] ,
         \SB1_1_18/Component_Function_3/NAND4_in[3] ,
         \SB1_1_18/Component_Function_3/NAND4_in[1] ,
         \SB1_1_18/Component_Function_4/NAND4_in[3] ,
         \SB1_1_18/Component_Function_4/NAND4_in[2] ,
         \SB1_1_18/Component_Function_4/NAND4_in[1] ,
         \SB1_1_18/Component_Function_4/NAND4_in[0] ,
         \SB1_1_19/Component_Function_2/NAND4_in[3] ,
         \SB1_1_19/Component_Function_2/NAND4_in[2] ,
         \SB1_1_19/Component_Function_2/NAND4_in[1] ,
         \SB1_1_19/Component_Function_2/NAND4_in[0] ,
         \SB1_1_19/Component_Function_3/NAND4_in[2] ,
         \SB1_1_19/Component_Function_3/NAND4_in[1] ,
         \SB1_1_19/Component_Function_3/NAND4_in[0] ,
         \SB1_1_19/Component_Function_4/NAND4_in[3] ,
         \SB1_1_19/Component_Function_4/NAND4_in[2] ,
         \SB1_1_19/Component_Function_4/NAND4_in[1] ,
         \SB1_1_19/Component_Function_4/NAND4_in[0] ,
         \SB1_1_20/Component_Function_2/NAND4_in[2] ,
         \SB1_1_20/Component_Function_2/NAND4_in[1] ,
         \SB1_1_20/Component_Function_3/NAND4_in[3] ,
         \SB1_1_20/Component_Function_3/NAND4_in[2] ,
         \SB1_1_20/Component_Function_3/NAND4_in[1] ,
         \SB1_1_20/Component_Function_3/NAND4_in[0] ,
         \SB1_1_20/Component_Function_4/NAND4_in[3] ,
         \SB1_1_20/Component_Function_4/NAND4_in[0] ,
         \SB1_1_21/Component_Function_2/NAND4_in[2] ,
         \SB1_1_21/Component_Function_2/NAND4_in[1] ,
         \SB1_1_21/Component_Function_2/NAND4_in[0] ,
         \SB1_1_21/Component_Function_3/NAND4_in[3] ,
         \SB1_1_21/Component_Function_3/NAND4_in[2] ,
         \SB1_1_21/Component_Function_3/NAND4_in[1] ,
         \SB1_1_21/Component_Function_3/NAND4_in[0] ,
         \SB1_1_21/Component_Function_4/NAND4_in[1] ,
         \SB1_1_21/Component_Function_4/NAND4_in[0] ,
         \SB1_1_22/Component_Function_2/NAND4_in[3] ,
         \SB1_1_22/Component_Function_2/NAND4_in[2] ,
         \SB1_1_22/Component_Function_3/NAND4_in[2] ,
         \SB1_1_22/Component_Function_3/NAND4_in[0] ,
         \SB1_1_22/Component_Function_4/NAND4_in[3] ,
         \SB1_1_22/Component_Function_4/NAND4_in[1] ,
         \SB1_1_22/Component_Function_4/NAND4_in[0] ,
         \SB1_1_23/Component_Function_2/NAND4_in[3] ,
         \SB1_1_23/Component_Function_2/NAND4_in[0] ,
         \SB1_1_23/Component_Function_3/NAND4_in[1] ,
         \SB1_1_23/Component_Function_3/NAND4_in[0] ,
         \SB1_1_23/Component_Function_4/NAND4_in[3] ,
         \SB1_1_23/Component_Function_4/NAND4_in[2] ,
         \SB1_1_23/Component_Function_4/NAND4_in[1] ,
         \SB1_1_23/Component_Function_4/NAND4_in[0] ,
         \SB1_1_24/Component_Function_2/NAND4_in[1] ,
         \SB1_1_24/Component_Function_3/NAND4_in[3] ,
         \SB1_1_24/Component_Function_3/NAND4_in[0] ,
         \SB1_1_24/Component_Function_4/NAND4_in[1] ,
         \SB1_1_24/Component_Function_4/NAND4_in[0] ,
         \SB1_1_25/Component_Function_2/NAND4_in[2] ,
         \SB1_1_25/Component_Function_2/NAND4_in[1] ,
         \SB1_1_25/Component_Function_2/NAND4_in[0] ,
         \SB1_1_25/Component_Function_3/NAND4_in[2] ,
         \SB1_1_25/Component_Function_3/NAND4_in[1] ,
         \SB1_1_25/Component_Function_3/NAND4_in[0] ,
         \SB1_1_25/Component_Function_4/NAND4_in[3] ,
         \SB1_1_25/Component_Function_4/NAND4_in[2] ,
         \SB1_1_25/Component_Function_4/NAND4_in[1] ,
         \SB1_1_25/Component_Function_4/NAND4_in[0] ,
         \SB1_1_26/Component_Function_2/NAND4_in[2] ,
         \SB1_1_26/Component_Function_3/NAND4_in[3] ,
         \SB1_1_26/Component_Function_3/NAND4_in[1] ,
         \SB1_1_26/Component_Function_3/NAND4_in[0] ,
         \SB1_1_26/Component_Function_4/NAND4_in[3] ,
         \SB1_1_26/Component_Function_4/NAND4_in[2] ,
         \SB1_1_26/Component_Function_4/NAND4_in[1] ,
         \SB1_1_26/Component_Function_4/NAND4_in[0] ,
         \SB1_1_27/Component_Function_2/NAND4_in[2] ,
         \SB1_1_27/Component_Function_2/NAND4_in[0] ,
         \SB1_1_27/Component_Function_3/NAND4_in[3] ,
         \SB1_1_27/Component_Function_3/NAND4_in[1] ,
         \SB1_1_27/Component_Function_3/NAND4_in[0] ,
         \SB1_1_27/Component_Function_4/NAND4_in[2] ,
         \SB1_1_27/Component_Function_4/NAND4_in[1] ,
         \SB1_1_27/Component_Function_4/NAND4_in[0] ,
         \SB1_1_28/Component_Function_2/NAND4_in[3] ,
         \SB1_1_28/Component_Function_2/NAND4_in[2] ,
         \SB1_1_28/Component_Function_2/NAND4_in[1] ,
         \SB1_1_28/Component_Function_3/NAND4_in[1] ,
         \SB1_1_28/Component_Function_3/NAND4_in[0] ,
         \SB1_1_28/Component_Function_4/NAND4_in[3] ,
         \SB1_1_28/Component_Function_4/NAND4_in[2] ,
         \SB1_1_28/Component_Function_4/NAND4_in[1] ,
         \SB1_1_28/Component_Function_4/NAND4_in[0] ,
         \SB1_1_29/Component_Function_2/NAND4_in[3] ,
         \SB1_1_29/Component_Function_2/NAND4_in[2] ,
         \SB1_1_29/Component_Function_2/NAND4_in[1] ,
         \SB1_1_29/Component_Function_2/NAND4_in[0] ,
         \SB1_1_29/Component_Function_3/NAND4_in[1] ,
         \SB1_1_29/Component_Function_3/NAND4_in[0] ,
         \SB1_1_29/Component_Function_4/NAND4_in[1] ,
         \SB1_1_29/Component_Function_4/NAND4_in[0] ,
         \SB1_1_30/Component_Function_2/NAND4_in[2] ,
         \SB1_1_30/Component_Function_2/NAND4_in[0] ,
         \SB1_1_30/Component_Function_3/NAND4_in[1] ,
         \SB1_1_30/Component_Function_3/NAND4_in[0] ,
         \SB1_1_30/Component_Function_4/NAND4_in[1] ,
         \SB1_1_31/Component_Function_2/NAND4_in[1] ,
         \SB1_1_31/Component_Function_2/NAND4_in[0] ,
         \SB1_1_31/Component_Function_3/NAND4_in[3] ,
         \SB1_1_31/Component_Function_3/NAND4_in[1] ,
         \SB1_1_31/Component_Function_3/NAND4_in[0] ,
         \SB1_1_31/Component_Function_4/NAND4_in[2] ,
         \SB1_1_31/Component_Function_4/NAND4_in[1] ,
         \SB1_1_31/Component_Function_4/NAND4_in[0] ,
         \SB2_1_0/Component_Function_2/NAND4_in[3] ,
         \SB2_1_0/Component_Function_2/NAND4_in[2] ,
         \SB2_1_0/Component_Function_3/NAND4_in[3] ,
         \SB2_1_0/Component_Function_4/NAND4_in[3] ,
         \SB2_1_0/Component_Function_4/NAND4_in[2] ,
         \SB2_1_0/Component_Function_4/NAND4_in[1] ,
         \SB2_1_0/Component_Function_4/NAND4_in[0] ,
         \SB2_1_1/Component_Function_2/NAND4_in[3] ,
         \SB2_1_1/Component_Function_3/NAND4_in[3] ,
         \SB2_1_1/Component_Function_3/NAND4_in[0] ,
         \SB2_1_1/Component_Function_4/NAND4_in[2] ,
         \SB2_1_1/Component_Function_4/NAND4_in[1] ,
         \SB2_1_1/Component_Function_4/NAND4_in[0] ,
         \SB2_1_2/Component_Function_2/NAND4_in[3] ,
         \SB2_1_2/Component_Function_2/NAND4_in[2] ,
         \SB2_1_2/Component_Function_3/NAND4_in[2] ,
         \SB2_1_2/Component_Function_3/NAND4_in[1] ,
         \SB2_1_2/Component_Function_3/NAND4_in[0] ,
         \SB2_1_2/Component_Function_4/NAND4_in[3] ,
         \SB2_1_2/Component_Function_4/NAND4_in[1] ,
         \SB2_1_2/Component_Function_4/NAND4_in[0] ,
         \SB2_1_3/Component_Function_2/NAND4_in[3] ,
         \SB2_1_3/Component_Function_2/NAND4_in[2] ,
         \SB2_1_3/Component_Function_2/NAND4_in[1] ,
         \SB2_1_3/Component_Function_2/NAND4_in[0] ,
         \SB2_1_3/Component_Function_3/NAND4_in[2] ,
         \SB2_1_3/Component_Function_4/NAND4_in[3] ,
         \SB2_1_3/Component_Function_4/NAND4_in[1] ,
         \SB2_1_3/Component_Function_4/NAND4_in[0] ,
         \SB2_1_4/Component_Function_2/NAND4_in[2] ,
         \SB2_1_4/Component_Function_2/NAND4_in[0] ,
         \SB2_1_4/Component_Function_3/NAND4_in[3] ,
         \SB2_1_4/Component_Function_3/NAND4_in[1] ,
         \SB2_1_4/Component_Function_4/NAND4_in[2] ,
         \SB2_1_4/Component_Function_4/NAND4_in[1] ,
         \SB2_1_4/Component_Function_4/NAND4_in[0] ,
         \SB2_1_5/Component_Function_2/NAND4_in[3] ,
         \SB2_1_5/Component_Function_2/NAND4_in[0] ,
         \SB2_1_5/Component_Function_3/NAND4_in[3] ,
         \SB2_1_5/Component_Function_3/NAND4_in[2] ,
         \SB2_1_5/Component_Function_3/NAND4_in[1] ,
         \SB2_1_5/Component_Function_3/NAND4_in[0] ,
         \SB2_1_5/Component_Function_4/NAND4_in[3] ,
         \SB2_1_5/Component_Function_4/NAND4_in[2] ,
         \SB2_1_5/Component_Function_4/NAND4_in[1] ,
         \SB2_1_5/Component_Function_4/NAND4_in[0] ,
         \SB2_1_6/Component_Function_2/NAND4_in[2] ,
         \SB2_1_6/Component_Function_2/NAND4_in[1] ,
         \SB2_1_6/Component_Function_2/NAND4_in[0] ,
         \SB2_1_6/Component_Function_3/NAND4_in[2] ,
         \SB2_1_6/Component_Function_3/NAND4_in[0] ,
         \SB2_1_6/Component_Function_4/NAND4_in[3] ,
         \SB2_1_6/Component_Function_4/NAND4_in[2] ,
         \SB2_1_6/Component_Function_4/NAND4_in[1] ,
         \SB2_1_6/Component_Function_4/NAND4_in[0] ,
         \SB2_1_7/Component_Function_2/NAND4_in[3] ,
         \SB2_1_7/Component_Function_2/NAND4_in[2] ,
         \SB2_1_7/Component_Function_2/NAND4_in[0] ,
         \SB2_1_7/Component_Function_4/NAND4_in[3] ,
         \SB2_1_7/Component_Function_4/NAND4_in[2] ,
         \SB2_1_7/Component_Function_4/NAND4_in[1] ,
         \SB2_1_8/Component_Function_2/NAND4_in[3] ,
         \SB2_1_8/Component_Function_2/NAND4_in[2] ,
         \SB2_1_8/Component_Function_2/NAND4_in[1] ,
         \SB2_1_8/Component_Function_2/NAND4_in[0] ,
         \SB2_1_8/Component_Function_3/NAND4_in[2] ,
         \SB2_1_8/Component_Function_3/NAND4_in[1] ,
         \SB2_1_8/Component_Function_3/NAND4_in[0] ,
         \SB2_1_8/Component_Function_4/NAND4_in[3] ,
         \SB2_1_8/Component_Function_4/NAND4_in[2] ,
         \SB2_1_8/Component_Function_4/NAND4_in[1] ,
         \SB2_1_8/Component_Function_4/NAND4_in[0] ,
         \SB2_1_9/Component_Function_2/NAND4_in[3] ,
         \SB2_1_9/Component_Function_2/NAND4_in[2] ,
         \SB2_1_9/Component_Function_2/NAND4_in[0] ,
         \SB2_1_9/Component_Function_3/NAND4_in[3] ,
         \SB2_1_9/Component_Function_3/NAND4_in[2] ,
         \SB2_1_9/Component_Function_3/NAND4_in[1] ,
         \SB2_1_9/Component_Function_3/NAND4_in[0] ,
         \SB2_1_9/Component_Function_4/NAND4_in[3] ,
         \SB2_1_9/Component_Function_4/NAND4_in[2] ,
         \SB2_1_9/Component_Function_4/NAND4_in[1] ,
         \SB2_1_9/Component_Function_4/NAND4_in[0] ,
         \SB2_1_10/Component_Function_2/NAND4_in[2] ,
         \SB2_1_10/Component_Function_2/NAND4_in[1] ,
         \SB2_1_10/Component_Function_2/NAND4_in[0] ,
         \SB2_1_10/Component_Function_3/NAND4_in[3] ,
         \SB2_1_10/Component_Function_4/NAND4_in[3] ,
         \SB2_1_10/Component_Function_4/NAND4_in[1] ,
         \SB2_1_10/Component_Function_4/NAND4_in[0] ,
         \SB2_1_11/Component_Function_2/NAND4_in[3] ,
         \SB2_1_11/Component_Function_2/NAND4_in[1] ,
         \SB2_1_11/Component_Function_2/NAND4_in[0] ,
         \SB2_1_11/Component_Function_3/NAND4_in[3] ,
         \SB2_1_11/Component_Function_3/NAND4_in[2] ,
         \SB2_1_11/Component_Function_3/NAND4_in[1] ,
         \SB2_1_11/Component_Function_3/NAND4_in[0] ,
         \SB2_1_11/Component_Function_4/NAND4_in[3] ,
         \SB2_1_11/Component_Function_4/NAND4_in[2] ,
         \SB2_1_11/Component_Function_4/NAND4_in[1] ,
         \SB2_1_11/Component_Function_4/NAND4_in[0] ,
         \SB2_1_12/Component_Function_2/NAND4_in[2] ,
         \SB2_1_12/Component_Function_2/NAND4_in[1] ,
         \SB2_1_12/Component_Function_2/NAND4_in[0] ,
         \SB2_1_12/Component_Function_3/NAND4_in[3] ,
         \SB2_1_12/Component_Function_3/NAND4_in[0] ,
         \SB2_1_12/Component_Function_4/NAND4_in[3] ,
         \SB2_1_12/Component_Function_4/NAND4_in[0] ,
         \SB2_1_13/Component_Function_2/NAND4_in[2] ,
         \SB2_1_13/Component_Function_2/NAND4_in[0] ,
         \SB2_1_13/Component_Function_3/NAND4_in[3] ,
         \SB2_1_13/Component_Function_3/NAND4_in[1] ,
         \SB2_1_13/Component_Function_4/NAND4_in[3] ,
         \SB2_1_13/Component_Function_4/NAND4_in[1] ,
         \SB2_1_13/Component_Function_4/NAND4_in[0] ,
         \SB2_1_14/Component_Function_2/NAND4_in[2] ,
         \SB2_1_14/Component_Function_2/NAND4_in[1] ,
         \SB2_1_14/Component_Function_2/NAND4_in[0] ,
         \SB2_1_14/Component_Function_3/NAND4_in[3] ,
         \SB2_1_14/Component_Function_3/NAND4_in[2] ,
         \SB2_1_14/Component_Function_3/NAND4_in[1] ,
         \SB2_1_14/Component_Function_3/NAND4_in[0] ,
         \SB2_1_14/Component_Function_4/NAND4_in[3] ,
         \SB2_1_14/Component_Function_4/NAND4_in[1] ,
         \SB2_1_14/Component_Function_4/NAND4_in[0] ,
         \SB2_1_15/Component_Function_2/NAND4_in[3] ,
         \SB2_1_15/Component_Function_2/NAND4_in[1] ,
         \SB2_1_15/Component_Function_2/NAND4_in[0] ,
         \SB2_1_15/Component_Function_3/NAND4_in[3] ,
         \SB2_1_15/Component_Function_3/NAND4_in[2] ,
         \SB2_1_15/Component_Function_3/NAND4_in[1] ,
         \SB2_1_15/Component_Function_4/NAND4_in[3] ,
         \SB2_1_15/Component_Function_4/NAND4_in[1] ,
         \SB2_1_15/Component_Function_4/NAND4_in[0] ,
         \SB2_1_16/Component_Function_2/NAND4_in[2] ,
         \SB2_1_16/Component_Function_2/NAND4_in[0] ,
         \SB2_1_16/Component_Function_3/NAND4_in[0] ,
         \SB2_1_16/Component_Function_4/NAND4_in[3] ,
         \SB2_1_16/Component_Function_4/NAND4_in[1] ,
         \SB2_1_16/Component_Function_4/NAND4_in[0] ,
         \SB2_1_17/Component_Function_2/NAND4_in[3] ,
         \SB2_1_17/Component_Function_2/NAND4_in[1] ,
         \SB2_1_17/Component_Function_2/NAND4_in[0] ,
         \SB2_1_17/Component_Function_3/NAND4_in[2] ,
         \SB2_1_17/Component_Function_3/NAND4_in[1] ,
         \SB2_1_17/Component_Function_3/NAND4_in[0] ,
         \SB2_1_17/Component_Function_4/NAND4_in[3] ,
         \SB2_1_17/Component_Function_4/NAND4_in[1] ,
         \SB2_1_17/Component_Function_4/NAND4_in[0] ,
         \SB2_1_18/Component_Function_2/NAND4_in[3] ,
         \SB2_1_18/Component_Function_2/NAND4_in[1] ,
         \SB2_1_18/Component_Function_2/NAND4_in[0] ,
         \SB2_1_18/Component_Function_3/NAND4_in[3] ,
         \SB2_1_18/Component_Function_3/NAND4_in[1] ,
         \SB2_1_18/Component_Function_3/NAND4_in[0] ,
         \SB2_1_18/Component_Function_4/NAND4_in[3] ,
         \SB2_1_18/Component_Function_4/NAND4_in[2] ,
         \SB2_1_18/Component_Function_4/NAND4_in[1] ,
         \SB2_1_18/Component_Function_4/NAND4_in[0] ,
         \SB2_1_19/Component_Function_2/NAND4_in[1] ,
         \SB2_1_19/Component_Function_2/NAND4_in[0] ,
         \SB2_1_19/Component_Function_3/NAND4_in[3] ,
         \SB2_1_19/Component_Function_3/NAND4_in[2] ,
         \SB2_1_19/Component_Function_3/NAND4_in[1] ,
         \SB2_1_19/Component_Function_3/NAND4_in[0] ,
         \SB2_1_19/Component_Function_4/NAND4_in[3] ,
         \SB2_1_19/Component_Function_4/NAND4_in[1] ,
         \SB2_1_19/Component_Function_4/NAND4_in[0] ,
         \SB2_1_20/Component_Function_2/NAND4_in[3] ,
         \SB2_1_20/Component_Function_2/NAND4_in[2] ,
         \SB2_1_20/Component_Function_2/NAND4_in[1] ,
         \SB2_1_20/Component_Function_2/NAND4_in[0] ,
         \SB2_1_20/Component_Function_4/NAND4_in[3] ,
         \SB2_1_20/Component_Function_4/NAND4_in[1] ,
         \SB2_1_20/Component_Function_4/NAND4_in[0] ,
         \SB2_1_21/Component_Function_2/NAND4_in[2] ,
         \SB2_1_21/Component_Function_2/NAND4_in[1] ,
         \SB2_1_21/Component_Function_3/NAND4_in[3] ,
         \SB2_1_21/Component_Function_3/NAND4_in[2] ,
         \SB2_1_21/Component_Function_3/NAND4_in[1] ,
         \SB2_1_21/Component_Function_3/NAND4_in[0] ,
         \SB2_1_21/Component_Function_4/NAND4_in[3] ,
         \SB2_1_21/Component_Function_4/NAND4_in[2] ,
         \SB2_1_21/Component_Function_4/NAND4_in[1] ,
         \SB2_1_21/Component_Function_4/NAND4_in[0] ,
         \SB2_1_22/Component_Function_2/NAND4_in[3] ,
         \SB2_1_22/Component_Function_2/NAND4_in[2] ,
         \SB2_1_22/Component_Function_2/NAND4_in[1] ,
         \SB2_1_22/Component_Function_2/NAND4_in[0] ,
         \SB2_1_22/Component_Function_3/NAND4_in[2] ,
         \SB2_1_22/Component_Function_3/NAND4_in[0] ,
         \SB2_1_22/Component_Function_4/NAND4_in[3] ,
         \SB2_1_22/Component_Function_4/NAND4_in[1] ,
         \SB2_1_22/Component_Function_4/NAND4_in[0] ,
         \SB2_1_23/Component_Function_2/NAND4_in[2] ,
         \SB2_1_23/Component_Function_2/NAND4_in[1] ,
         \SB2_1_23/Component_Function_2/NAND4_in[0] ,
         \SB2_1_23/Component_Function_3/NAND4_in[3] ,
         \SB2_1_23/Component_Function_3/NAND4_in[2] ,
         \SB2_1_23/Component_Function_3/NAND4_in[1] ,
         \SB2_1_23/Component_Function_3/NAND4_in[0] ,
         \SB2_1_23/Component_Function_4/NAND4_in[3] ,
         \SB2_1_23/Component_Function_4/NAND4_in[1] ,
         \SB2_1_23/Component_Function_4/NAND4_in[0] ,
         \SB2_1_24/Component_Function_2/NAND4_in[2] ,
         \SB2_1_24/Component_Function_2/NAND4_in[1] ,
         \SB2_1_24/Component_Function_2/NAND4_in[0] ,
         \SB2_1_24/Component_Function_3/NAND4_in[3] ,
         \SB2_1_24/Component_Function_3/NAND4_in[2] ,
         \SB2_1_24/Component_Function_3/NAND4_in[0] ,
         \SB2_1_24/Component_Function_4/NAND4_in[3] ,
         \SB2_1_24/Component_Function_4/NAND4_in[2] ,
         \SB2_1_24/Component_Function_4/NAND4_in[1] ,
         \SB2_1_24/Component_Function_4/NAND4_in[0] ,
         \SB2_1_25/Component_Function_2/NAND4_in[1] ,
         \SB2_1_25/Component_Function_2/NAND4_in[0] ,
         \SB2_1_25/Component_Function_3/NAND4_in[2] ,
         \SB2_1_25/Component_Function_3/NAND4_in[1] ,
         \SB2_1_25/Component_Function_3/NAND4_in[0] ,
         \SB2_1_25/Component_Function_4/NAND4_in[2] ,
         \SB2_1_25/Component_Function_4/NAND4_in[1] ,
         \SB2_1_25/Component_Function_4/NAND4_in[0] ,
         \SB2_1_26/Component_Function_2/NAND4_in[2] ,
         \SB2_1_26/Component_Function_2/NAND4_in[1] ,
         \SB2_1_26/Component_Function_2/NAND4_in[0] ,
         \SB2_1_26/Component_Function_3/NAND4_in[3] ,
         \SB2_1_26/Component_Function_3/NAND4_in[2] ,
         \SB2_1_26/Component_Function_3/NAND4_in[1] ,
         \SB2_1_26/Component_Function_3/NAND4_in[0] ,
         \SB2_1_26/Component_Function_4/NAND4_in[3] ,
         \SB2_1_26/Component_Function_4/NAND4_in[1] ,
         \SB2_1_26/Component_Function_4/NAND4_in[0] ,
         \SB2_1_27/Component_Function_2/NAND4_in[3] ,
         \SB2_1_27/Component_Function_2/NAND4_in[2] ,
         \SB2_1_27/Component_Function_2/NAND4_in[1] ,
         \SB2_1_27/Component_Function_2/NAND4_in[0] ,
         \SB2_1_27/Component_Function_3/NAND4_in[3] ,
         \SB2_1_27/Component_Function_3/NAND4_in[2] ,
         \SB2_1_27/Component_Function_3/NAND4_in[0] ,
         \SB2_1_27/Component_Function_4/NAND4_in[3] ,
         \SB2_1_27/Component_Function_4/NAND4_in[2] ,
         \SB2_1_27/Component_Function_4/NAND4_in[1] ,
         \SB2_1_27/Component_Function_4/NAND4_in[0] ,
         \SB2_1_28/Component_Function_2/NAND4_in[1] ,
         \SB2_1_28/Component_Function_2/NAND4_in[0] ,
         \SB2_1_28/Component_Function_3/NAND4_in[1] ,
         \SB2_1_28/Component_Function_3/NAND4_in[0] ,
         \SB2_1_28/Component_Function_4/NAND4_in[3] ,
         \SB2_1_28/Component_Function_4/NAND4_in[2] ,
         \SB2_1_28/Component_Function_4/NAND4_in[1] ,
         \SB2_1_28/Component_Function_4/NAND4_in[0] ,
         \SB2_1_29/Component_Function_2/NAND4_in[2] ,
         \SB2_1_29/Component_Function_2/NAND4_in[1] ,
         \SB2_1_29/Component_Function_2/NAND4_in[0] ,
         \SB2_1_29/Component_Function_3/NAND4_in[3] ,
         \SB2_1_29/Component_Function_3/NAND4_in[2] ,
         \SB2_1_29/Component_Function_3/NAND4_in[1] ,
         \SB2_1_29/Component_Function_3/NAND4_in[0] ,
         \SB2_1_29/Component_Function_4/NAND4_in[2] ,
         \SB2_1_29/Component_Function_4/NAND4_in[1] ,
         \SB2_1_29/Component_Function_4/NAND4_in[0] ,
         \SB2_1_30/Component_Function_2/NAND4_in[2] ,
         \SB2_1_30/Component_Function_2/NAND4_in[1] ,
         \SB2_1_30/Component_Function_2/NAND4_in[0] ,
         \SB2_1_30/Component_Function_3/NAND4_in[2] ,
         \SB2_1_30/Component_Function_3/NAND4_in[0] ,
         \SB2_1_30/Component_Function_4/NAND4_in[2] ,
         \SB2_1_30/Component_Function_4/NAND4_in[1] ,
         \SB2_1_30/Component_Function_4/NAND4_in[0] ,
         \SB2_1_31/Component_Function_2/NAND4_in[3] ,
         \SB2_1_31/Component_Function_2/NAND4_in[2] ,
         \SB2_1_31/Component_Function_2/NAND4_in[1] ,
         \SB2_1_31/Component_Function_2/NAND4_in[0] ,
         \SB2_1_31/Component_Function_3/NAND4_in[3] ,
         \SB2_1_31/Component_Function_3/NAND4_in[2] ,
         \SB2_1_31/Component_Function_4/NAND4_in[3] ,
         \SB2_1_31/Component_Function_4/NAND4_in[1] ,
         \SB2_1_31/Component_Function_4/NAND4_in[0] ,
         \SB1_2_0/Component_Function_2/NAND4_in[3] ,
         \SB1_2_0/Component_Function_2/NAND4_in[2] ,
         \SB1_2_0/Component_Function_2/NAND4_in[1] ,
         \SB1_2_0/Component_Function_2/NAND4_in[0] ,
         \SB1_2_0/Component_Function_3/NAND4_in[3] ,
         \SB1_2_0/Component_Function_3/NAND4_in[2] ,
         \SB1_2_0/Component_Function_3/NAND4_in[1] ,
         \SB1_2_0/Component_Function_3/NAND4_in[0] ,
         \SB1_2_0/Component_Function_4/NAND4_in[2] ,
         \SB1_2_0/Component_Function_4/NAND4_in[1] ,
         \SB1_2_0/Component_Function_4/NAND4_in[0] ,
         \SB1_2_1/Component_Function_2/NAND4_in[2] ,
         \SB1_2_1/Component_Function_2/NAND4_in[1] ,
         \SB1_2_1/Component_Function_3/NAND4_in[0] ,
         \SB1_2_1/Component_Function_4/NAND4_in[3] ,
         \SB1_2_2/Component_Function_2/NAND4_in[3] ,
         \SB1_2_2/Component_Function_2/NAND4_in[2] ,
         \SB1_2_2/Component_Function_2/NAND4_in[1] ,
         \SB1_2_2/Component_Function_2/NAND4_in[0] ,
         \SB1_2_2/Component_Function_3/NAND4_in[2] ,
         \SB1_2_2/Component_Function_3/NAND4_in[1] ,
         \SB1_2_2/Component_Function_4/NAND4_in[3] ,
         \SB1_2_2/Component_Function_4/NAND4_in[1] ,
         \SB1_2_2/Component_Function_4/NAND4_in[0] ,
         \SB1_2_3/Component_Function_2/NAND4_in[1] ,
         \SB1_2_3/Component_Function_2/NAND4_in[0] ,
         \SB1_2_3/Component_Function_3/NAND4_in[3] ,
         \SB1_2_3/Component_Function_3/NAND4_in[2] ,
         \SB1_2_3/Component_Function_3/NAND4_in[1] ,
         \SB1_2_3/Component_Function_3/NAND4_in[0] ,
         \SB1_2_3/Component_Function_4/NAND4_in[3] ,
         \SB1_2_3/Component_Function_4/NAND4_in[2] ,
         \SB1_2_3/Component_Function_4/NAND4_in[1] ,
         \SB1_2_3/Component_Function_4/NAND4_in[0] ,
         \SB1_2_4/Component_Function_2/NAND4_in[3] ,
         \SB1_2_4/Component_Function_2/NAND4_in[2] ,
         \SB1_2_4/Component_Function_2/NAND4_in[1] ,
         \SB1_2_4/Component_Function_2/NAND4_in[0] ,
         \SB1_2_4/Component_Function_3/NAND4_in[1] ,
         \SB1_2_4/Component_Function_3/NAND4_in[0] ,
         \SB1_2_4/Component_Function_4/NAND4_in[3] ,
         \SB1_2_4/Component_Function_4/NAND4_in[1] ,
         \SB1_2_4/Component_Function_4/NAND4_in[0] ,
         \SB1_2_5/Component_Function_2/NAND4_in[2] ,
         \SB1_2_5/Component_Function_2/NAND4_in[1] ,
         \SB1_2_5/Component_Function_2/NAND4_in[0] ,
         \SB1_2_5/Component_Function_3/NAND4_in[3] ,
         \SB1_2_5/Component_Function_3/NAND4_in[1] ,
         \SB1_2_5/Component_Function_4/NAND4_in[3] ,
         \SB1_2_6/Component_Function_2/NAND4_in[2] ,
         \SB1_2_6/Component_Function_2/NAND4_in[1] ,
         \SB1_2_6/Component_Function_2/NAND4_in[0] ,
         \SB1_2_6/Component_Function_3/NAND4_in[3] ,
         \SB1_2_6/Component_Function_3/NAND4_in[1] ,
         \SB1_2_6/Component_Function_3/NAND4_in[0] ,
         \SB1_2_6/Component_Function_4/NAND4_in[2] ,
         \SB1_2_6/Component_Function_4/NAND4_in[1] ,
         \SB1_2_6/Component_Function_4/NAND4_in[0] ,
         \SB1_2_7/Component_Function_2/NAND4_in[3] ,
         \SB1_2_7/Component_Function_2/NAND4_in[1] ,
         \SB1_2_7/Component_Function_2/NAND4_in[0] ,
         \SB1_2_7/Component_Function_3/NAND4_in[2] ,
         \SB1_2_7/Component_Function_3/NAND4_in[1] ,
         \SB1_2_7/Component_Function_3/NAND4_in[0] ,
         \SB1_2_7/Component_Function_4/NAND4_in[3] ,
         \SB1_2_7/Component_Function_4/NAND4_in[2] ,
         \SB1_2_7/Component_Function_4/NAND4_in[1] ,
         \SB1_2_7/Component_Function_4/NAND4_in[0] ,
         \SB1_2_8/Component_Function_2/NAND4_in[3] ,
         \SB1_2_8/Component_Function_2/NAND4_in[2] ,
         \SB1_2_8/Component_Function_3/NAND4_in[3] ,
         \SB1_2_8/Component_Function_3/NAND4_in[2] ,
         \SB1_2_8/Component_Function_3/NAND4_in[1] ,
         \SB1_2_8/Component_Function_3/NAND4_in[0] ,
         \SB1_2_8/Component_Function_4/NAND4_in[3] ,
         \SB1_2_8/Component_Function_4/NAND4_in[2] ,
         \SB1_2_8/Component_Function_4/NAND4_in[1] ,
         \SB1_2_8/Component_Function_4/NAND4_in[0] ,
         \SB1_2_9/Component_Function_2/NAND4_in[3] ,
         \SB1_2_9/Component_Function_2/NAND4_in[1] ,
         \SB1_2_9/Component_Function_3/NAND4_in[1] ,
         \SB1_2_9/Component_Function_3/NAND4_in[0] ,
         \SB1_2_9/Component_Function_4/NAND4_in[3] ,
         \SB1_2_9/Component_Function_4/NAND4_in[1] ,
         \SB1_2_9/Component_Function_4/NAND4_in[0] ,
         \SB1_2_10/Component_Function_2/NAND4_in[1] ,
         \SB1_2_10/Component_Function_3/NAND4_in[1] ,
         \SB1_2_10/Component_Function_3/NAND4_in[0] ,
         \SB1_2_10/Component_Function_4/NAND4_in[2] ,
         \SB1_2_10/Component_Function_4/NAND4_in[1] ,
         \SB1_2_10/Component_Function_4/NAND4_in[0] ,
         \SB1_2_11/Component_Function_2/NAND4_in[0] ,
         \SB1_2_11/Component_Function_3/NAND4_in[1] ,
         \SB1_2_11/Component_Function_3/NAND4_in[0] ,
         \SB1_2_11/Component_Function_4/NAND4_in[2] ,
         \SB1_2_11/Component_Function_4/NAND4_in[1] ,
         \SB1_2_12/Component_Function_2/NAND4_in[2] ,
         \SB1_2_12/Component_Function_2/NAND4_in[0] ,
         \SB1_2_12/Component_Function_3/NAND4_in[3] ,
         \SB1_2_12/Component_Function_3/NAND4_in[1] ,
         \SB1_2_12/Component_Function_4/NAND4_in[3] ,
         \SB1_2_12/Component_Function_4/NAND4_in[1] ,
         \SB1_2_12/Component_Function_4/NAND4_in[0] ,
         \SB1_2_13/Component_Function_2/NAND4_in[2] ,
         \SB1_2_13/Component_Function_2/NAND4_in[1] ,
         \SB1_2_13/Component_Function_2/NAND4_in[0] ,
         \SB1_2_13/Component_Function_3/NAND4_in[3] ,
         \SB1_2_13/Component_Function_3/NAND4_in[1] ,
         \SB1_2_13/Component_Function_3/NAND4_in[0] ,
         \SB1_2_13/Component_Function_4/NAND4_in[2] ,
         \SB1_2_13/Component_Function_4/NAND4_in[1] ,
         \SB1_2_13/Component_Function_4/NAND4_in[0] ,
         \SB1_2_14/Component_Function_2/NAND4_in[0] ,
         \SB1_2_14/Component_Function_3/NAND4_in[1] ,
         \SB1_2_14/Component_Function_4/NAND4_in[3] ,
         \SB1_2_14/Component_Function_4/NAND4_in[2] ,
         \SB1_2_14/Component_Function_4/NAND4_in[1] ,
         \SB1_2_14/Component_Function_4/NAND4_in[0] ,
         \SB1_2_15/Component_Function_2/NAND4_in[3] ,
         \SB1_2_15/Component_Function_2/NAND4_in[1] ,
         \SB1_2_15/Component_Function_2/NAND4_in[0] ,
         \SB1_2_15/Component_Function_3/NAND4_in[2] ,
         \SB1_2_15/Component_Function_3/NAND4_in[0] ,
         \SB1_2_15/Component_Function_4/NAND4_in[0] ,
         \SB1_2_16/Component_Function_2/NAND4_in[3] ,
         \SB1_2_16/Component_Function_2/NAND4_in[2] ,
         \SB1_2_16/Component_Function_2/NAND4_in[1] ,
         \SB1_2_16/Component_Function_2/NAND4_in[0] ,
         \SB1_2_16/Component_Function_3/NAND4_in[1] ,
         \SB1_2_16/Component_Function_3/NAND4_in[0] ,
         \SB1_2_16/Component_Function_4/NAND4_in[3] ,
         \SB1_2_16/Component_Function_4/NAND4_in[1] ,
         \SB1_2_16/Component_Function_4/NAND4_in[0] ,
         \SB1_2_17/Component_Function_2/NAND4_in[2] ,
         \SB1_2_17/Component_Function_2/NAND4_in[1] ,
         \SB1_2_17/Component_Function_3/NAND4_in[3] ,
         \SB1_2_17/Component_Function_3/NAND4_in[2] ,
         \SB1_2_17/Component_Function_3/NAND4_in[0] ,
         \SB1_2_17/Component_Function_4/NAND4_in[2] ,
         \SB1_2_17/Component_Function_4/NAND4_in[1] ,
         \SB1_2_17/Component_Function_4/NAND4_in[0] ,
         \SB1_2_18/Component_Function_2/NAND4_in[2] ,
         \SB1_2_18/Component_Function_3/NAND4_in[1] ,
         \SB1_2_18/Component_Function_3/NAND4_in[0] ,
         \SB1_2_18/Component_Function_4/NAND4_in[3] ,
         \SB1_2_18/Component_Function_4/NAND4_in[1] ,
         \SB1_2_19/Component_Function_2/NAND4_in[2] ,
         \SB1_2_19/Component_Function_2/NAND4_in[1] ,
         \SB1_2_19/Component_Function_3/NAND4_in[1] ,
         \SB1_2_19/Component_Function_3/NAND4_in[0] ,
         \SB1_2_19/Component_Function_4/NAND4_in[3] ,
         \SB1_2_19/Component_Function_4/NAND4_in[1] ,
         \SB1_2_19/Component_Function_4/NAND4_in[0] ,
         \SB1_2_20/Component_Function_2/NAND4_in[3] ,
         \SB1_2_20/Component_Function_2/NAND4_in[2] ,
         \SB1_2_20/Component_Function_2/NAND4_in[1] ,
         \SB1_2_20/Component_Function_2/NAND4_in[0] ,
         \SB1_2_20/Component_Function_3/NAND4_in[1] ,
         \SB1_2_20/Component_Function_3/NAND4_in[0] ,
         \SB1_2_20/Component_Function_4/NAND4_in[3] ,
         \SB1_2_20/Component_Function_4/NAND4_in[2] ,
         \SB1_2_20/Component_Function_4/NAND4_in[1] ,
         \SB1_2_20/Component_Function_4/NAND4_in[0] ,
         \SB1_2_21/Component_Function_2/NAND4_in[3] ,
         \SB1_2_21/Component_Function_2/NAND4_in[1] ,
         \SB1_2_21/Component_Function_3/NAND4_in[3] ,
         \SB1_2_21/Component_Function_3/NAND4_in[2] ,
         \SB1_2_21/Component_Function_3/NAND4_in[0] ,
         \SB1_2_21/Component_Function_4/NAND4_in[3] ,
         \SB1_2_21/Component_Function_4/NAND4_in[1] ,
         \SB1_2_21/Component_Function_4/NAND4_in[0] ,
         \SB1_2_22/Component_Function_2/NAND4_in[1] ,
         \SB1_2_22/Component_Function_4/NAND4_in[2] ,
         \SB1_2_22/Component_Function_4/NAND4_in[1] ,
         \SB1_2_22/Component_Function_4/NAND4_in[0] ,
         \SB1_2_23/Component_Function_2/NAND4_in[2] ,
         \SB1_2_23/Component_Function_2/NAND4_in[1] ,
         \SB1_2_23/Component_Function_2/NAND4_in[0] ,
         \SB1_2_23/Component_Function_3/NAND4_in[2] ,
         \SB1_2_23/Component_Function_3/NAND4_in[1] ,
         \SB1_2_23/Component_Function_3/NAND4_in[0] ,
         \SB1_2_23/Component_Function_4/NAND4_in[3] ,
         \SB1_2_23/Component_Function_4/NAND4_in[2] ,
         \SB1_2_23/Component_Function_4/NAND4_in[1] ,
         \SB1_2_23/Component_Function_4/NAND4_in[0] ,
         \SB1_2_24/Component_Function_3/NAND4_in[1] ,
         \SB1_2_24/Component_Function_3/NAND4_in[0] ,
         \SB1_2_24/Component_Function_4/NAND4_in[3] ,
         \SB1_2_24/Component_Function_4/NAND4_in[2] ,
         \SB1_2_24/Component_Function_4/NAND4_in[1] ,
         \SB1_2_25/Component_Function_2/NAND4_in[2] ,
         \SB1_2_25/Component_Function_2/NAND4_in[0] ,
         \SB1_2_25/Component_Function_3/NAND4_in[1] ,
         \SB1_2_25/Component_Function_3/NAND4_in[0] ,
         \SB1_2_25/Component_Function_4/NAND4_in[2] ,
         \SB1_2_25/Component_Function_4/NAND4_in[1] ,
         \SB1_2_25/Component_Function_4/NAND4_in[0] ,
         \SB1_2_26/Component_Function_2/NAND4_in[3] ,
         \SB1_2_26/Component_Function_2/NAND4_in[2] ,
         \SB1_2_26/Component_Function_2/NAND4_in[1] ,
         \SB1_2_26/Component_Function_2/NAND4_in[0] ,
         \SB1_2_26/Component_Function_3/NAND4_in[1] ,
         \SB1_2_26/Component_Function_3/NAND4_in[0] ,
         \SB1_2_26/Component_Function_4/NAND4_in[3] ,
         \SB1_2_26/Component_Function_4/NAND4_in[1] ,
         \SB1_2_27/Component_Function_2/NAND4_in[1] ,
         \SB1_2_27/Component_Function_3/NAND4_in[2] ,
         \SB1_2_27/Component_Function_3/NAND4_in[1] ,
         \SB1_2_27/Component_Function_3/NAND4_in[0] ,
         \SB1_2_27/Component_Function_4/NAND4_in[3] ,
         \SB1_2_27/Component_Function_4/NAND4_in[1] ,
         \SB1_2_28/Component_Function_2/NAND4_in[2] ,
         \SB1_2_28/Component_Function_2/NAND4_in[1] ,
         \SB1_2_28/Component_Function_2/NAND4_in[0] ,
         \SB1_2_28/Component_Function_3/NAND4_in[1] ,
         \SB1_2_28/Component_Function_3/NAND4_in[0] ,
         \SB1_2_28/Component_Function_4/NAND4_in[2] ,
         \SB1_2_28/Component_Function_4/NAND4_in[1] ,
         \SB1_2_28/Component_Function_4/NAND4_in[0] ,
         \SB1_2_29/Component_Function_2/NAND4_in[3] ,
         \SB1_2_29/Component_Function_2/NAND4_in[2] ,
         \SB1_2_29/Component_Function_2/NAND4_in[0] ,
         \SB1_2_29/Component_Function_3/NAND4_in[2] ,
         \SB1_2_29/Component_Function_3/NAND4_in[1] ,
         \SB1_2_29/Component_Function_4/NAND4_in[2] ,
         \SB1_2_29/Component_Function_4/NAND4_in[1] ,
         \SB1_2_29/Component_Function_4/NAND4_in[0] ,
         \SB1_2_30/Component_Function_3/NAND4_in[3] ,
         \SB1_2_30/Component_Function_3/NAND4_in[1] ,
         \SB1_2_30/Component_Function_3/NAND4_in[0] ,
         \SB1_2_30/Component_Function_4/NAND4_in[3] ,
         \SB1_2_30/Component_Function_4/NAND4_in[1] ,
         \SB1_2_30/Component_Function_4/NAND4_in[0] ,
         \SB1_2_31/Component_Function_2/NAND4_in[1] ,
         \SB1_2_31/Component_Function_2/NAND4_in[0] ,
         \SB1_2_31/Component_Function_3/NAND4_in[1] ,
         \SB1_2_31/Component_Function_3/NAND4_in[0] ,
         \SB1_2_31/Component_Function_4/NAND4_in[3] ,
         \SB1_2_31/Component_Function_4/NAND4_in[1] ,
         \SB1_2_31/Component_Function_4/NAND4_in[0] ,
         \SB2_2_0/Component_Function_2/NAND4_in[2] ,
         \SB2_2_0/Component_Function_2/NAND4_in[1] ,
         \SB2_2_0/Component_Function_2/NAND4_in[0] ,
         \SB2_2_0/Component_Function_3/NAND4_in[3] ,
         \SB2_2_0/Component_Function_3/NAND4_in[2] ,
         \SB2_2_0/Component_Function_3/NAND4_in[1] ,
         \SB2_2_0/Component_Function_3/NAND4_in[0] ,
         \SB2_2_0/Component_Function_4/NAND4_in[3] ,
         \SB2_2_0/Component_Function_4/NAND4_in[1] ,
         \SB2_2_0/Component_Function_4/NAND4_in[0] ,
         \SB2_2_1/Component_Function_2/NAND4_in[2] ,
         \SB2_2_1/Component_Function_2/NAND4_in[1] ,
         \SB2_2_1/Component_Function_2/NAND4_in[0] ,
         \SB2_2_1/Component_Function_3/NAND4_in[0] ,
         \SB2_2_1/Component_Function_4/NAND4_in[3] ,
         \SB2_2_1/Component_Function_4/NAND4_in[1] ,
         \SB2_2_2/Component_Function_2/NAND4_in[2] ,
         \SB2_2_2/Component_Function_2/NAND4_in[0] ,
         \SB2_2_2/Component_Function_3/NAND4_in[2] ,
         \SB2_2_2/Component_Function_3/NAND4_in[1] ,
         \SB2_2_2/Component_Function_3/NAND4_in[0] ,
         \SB2_2_2/Component_Function_4/NAND4_in[3] ,
         \SB2_2_2/Component_Function_4/NAND4_in[1] ,
         \SB2_2_2/Component_Function_4/NAND4_in[0] ,
         \SB2_2_3/Component_Function_2/NAND4_in[2] ,
         \SB2_2_3/Component_Function_2/NAND4_in[1] ,
         \SB2_2_3/Component_Function_3/NAND4_in[3] ,
         \SB2_2_3/Component_Function_3/NAND4_in[1] ,
         \SB2_2_3/Component_Function_3/NAND4_in[0] ,
         \SB2_2_3/Component_Function_4/NAND4_in[3] ,
         \SB2_2_3/Component_Function_4/NAND4_in[1] ,
         \SB2_2_3/Component_Function_4/NAND4_in[0] ,
         \SB2_2_4/Component_Function_2/NAND4_in[2] ,
         \SB2_2_4/Component_Function_2/NAND4_in[1] ,
         \SB2_2_4/Component_Function_2/NAND4_in[0] ,
         \SB2_2_4/Component_Function_3/NAND4_in[3] ,
         \SB2_2_4/Component_Function_3/NAND4_in[2] ,
         \SB2_2_4/Component_Function_4/NAND4_in[2] ,
         \SB2_2_4/Component_Function_4/NAND4_in[1] ,
         \SB2_2_5/Component_Function_2/NAND4_in[3] ,
         \SB2_2_5/Component_Function_2/NAND4_in[2] ,
         \SB2_2_5/Component_Function_2/NAND4_in[1] ,
         \SB2_2_5/Component_Function_3/NAND4_in[2] ,
         \SB2_2_5/Component_Function_3/NAND4_in[1] ,
         \SB2_2_5/Component_Function_3/NAND4_in[0] ,
         \SB2_2_5/Component_Function_4/NAND4_in[3] ,
         \SB2_2_5/Component_Function_4/NAND4_in[1] ,
         \SB2_2_5/Component_Function_4/NAND4_in[0] ,
         \SB2_2_6/Component_Function_2/NAND4_in[3] ,
         \SB2_2_6/Component_Function_2/NAND4_in[1] ,
         \SB2_2_6/Component_Function_2/NAND4_in[0] ,
         \SB2_2_6/Component_Function_3/NAND4_in[3] ,
         \SB2_2_6/Component_Function_3/NAND4_in[1] ,
         \SB2_2_6/Component_Function_3/NAND4_in[0] ,
         \SB2_2_6/Component_Function_4/NAND4_in[1] ,
         \SB2_2_6/Component_Function_4/NAND4_in[0] ,
         \SB2_2_7/Component_Function_2/NAND4_in[0] ,
         \SB2_2_7/Component_Function_3/NAND4_in[3] ,
         \SB2_2_7/Component_Function_3/NAND4_in[0] ,
         \SB2_2_7/Component_Function_4/NAND4_in[3] ,
         \SB2_2_7/Component_Function_4/NAND4_in[2] ,
         \SB2_2_7/Component_Function_4/NAND4_in[0] ,
         \SB2_2_8/Component_Function_2/NAND4_in[0] ,
         \SB2_2_8/Component_Function_4/NAND4_in[3] ,
         \SB2_2_8/Component_Function_4/NAND4_in[0] ,
         \SB2_2_9/Component_Function_3/NAND4_in[3] ,
         \SB2_2_9/Component_Function_3/NAND4_in[2] ,
         \SB2_2_9/Component_Function_3/NAND4_in[1] ,
         \SB2_2_9/Component_Function_3/NAND4_in[0] ,
         \SB2_2_9/Component_Function_4/NAND4_in[3] ,
         \SB2_2_9/Component_Function_4/NAND4_in[2] ,
         \SB2_2_9/Component_Function_4/NAND4_in[1] ,
         \SB2_2_9/Component_Function_4/NAND4_in[0] ,
         \SB2_2_10/Component_Function_2/NAND4_in[2] ,
         \SB2_2_10/Component_Function_2/NAND4_in[1] ,
         \SB2_2_10/Component_Function_3/NAND4_in[3] ,
         \SB2_2_10/Component_Function_3/NAND4_in[1] ,
         \SB2_2_10/Component_Function_4/NAND4_in[1] ,
         \SB2_2_11/Component_Function_2/NAND4_in[2] ,
         \SB2_2_11/Component_Function_2/NAND4_in[1] ,
         \SB2_2_11/Component_Function_2/NAND4_in[0] ,
         \SB2_2_11/Component_Function_3/NAND4_in[3] ,
         \SB2_2_11/Component_Function_3/NAND4_in[2] ,
         \SB2_2_11/Component_Function_4/NAND4_in[2] ,
         \SB2_2_11/Component_Function_4/NAND4_in[1] ,
         \SB2_2_11/Component_Function_4/NAND4_in[0] ,
         \SB2_2_12/Component_Function_2/NAND4_in[2] ,
         \SB2_2_12/Component_Function_2/NAND4_in[1] ,
         \SB2_2_12/Component_Function_2/NAND4_in[0] ,
         \SB2_2_12/Component_Function_3/NAND4_in[3] ,
         \SB2_2_12/Component_Function_3/NAND4_in[2] ,
         \SB2_2_12/Component_Function_4/NAND4_in[2] ,
         \SB2_2_12/Component_Function_4/NAND4_in[1] ,
         \SB2_2_12/Component_Function_4/NAND4_in[0] ,
         \SB2_2_13/Component_Function_2/NAND4_in[3] ,
         \SB2_2_13/Component_Function_2/NAND4_in[1] ,
         \SB2_2_13/Component_Function_2/NAND4_in[0] ,
         \SB2_2_13/Component_Function_3/NAND4_in[2] ,
         \SB2_2_13/Component_Function_3/NAND4_in[1] ,
         \SB2_2_13/Component_Function_3/NAND4_in[0] ,
         \SB2_2_13/Component_Function_4/NAND4_in[3] ,
         \SB2_2_13/Component_Function_4/NAND4_in[2] ,
         \SB2_2_13/Component_Function_4/NAND4_in[1] ,
         \SB2_2_13/Component_Function_4/NAND4_in[0] ,
         \SB2_2_14/Component_Function_2/NAND4_in[2] ,
         \SB2_2_14/Component_Function_2/NAND4_in[1] ,
         \SB2_2_14/Component_Function_3/NAND4_in[3] ,
         \SB2_2_14/Component_Function_3/NAND4_in[1] ,
         \SB2_2_14/Component_Function_3/NAND4_in[0] ,
         \SB2_2_14/Component_Function_4/NAND4_in[2] ,
         \SB2_2_14/Component_Function_4/NAND4_in[1] ,
         \SB2_2_14/Component_Function_4/NAND4_in[0] ,
         \SB2_2_15/Component_Function_2/NAND4_in[3] ,
         \SB2_2_15/Component_Function_2/NAND4_in[2] ,
         \SB2_2_15/Component_Function_2/NAND4_in[1] ,
         \SB2_2_15/Component_Function_2/NAND4_in[0] ,
         \SB2_2_15/Component_Function_3/NAND4_in[3] ,
         \SB2_2_15/Component_Function_3/NAND4_in[1] ,
         \SB2_2_15/Component_Function_4/NAND4_in[3] ,
         \SB2_2_15/Component_Function_4/NAND4_in[1] ,
         \SB2_2_15/Component_Function_4/NAND4_in[0] ,
         \SB2_2_16/Component_Function_2/NAND4_in[3] ,
         \SB2_2_16/Component_Function_2/NAND4_in[2] ,
         \SB2_2_16/Component_Function_3/NAND4_in[3] ,
         \SB2_2_16/Component_Function_3/NAND4_in[2] ,
         \SB2_2_16/Component_Function_3/NAND4_in[0] ,
         \SB2_2_16/Component_Function_4/NAND4_in[1] ,
         \SB2_2_16/Component_Function_4/NAND4_in[0] ,
         \SB2_2_17/Component_Function_2/NAND4_in[3] ,
         \SB2_2_17/Component_Function_2/NAND4_in[1] ,
         \SB2_2_17/Component_Function_2/NAND4_in[0] ,
         \SB2_2_17/Component_Function_3/NAND4_in[2] ,
         \SB2_2_17/Component_Function_3/NAND4_in[1] ,
         \SB2_2_17/Component_Function_3/NAND4_in[0] ,
         \SB2_2_17/Component_Function_4/NAND4_in[3] ,
         \SB2_2_17/Component_Function_4/NAND4_in[0] ,
         \SB2_2_18/Component_Function_2/NAND4_in[3] ,
         \SB2_2_18/Component_Function_2/NAND4_in[2] ,
         \SB2_2_18/Component_Function_2/NAND4_in[0] ,
         \SB2_2_18/Component_Function_3/NAND4_in[3] ,
         \SB2_2_18/Component_Function_3/NAND4_in[2] ,
         \SB2_2_18/Component_Function_3/NAND4_in[1] ,
         \SB2_2_18/Component_Function_4/NAND4_in[3] ,
         \SB2_2_18/Component_Function_4/NAND4_in[1] ,
         \SB2_2_18/Component_Function_4/NAND4_in[0] ,
         \SB2_2_19/Component_Function_2/NAND4_in[3] ,
         \SB2_2_19/Component_Function_2/NAND4_in[1] ,
         \SB2_2_19/Component_Function_2/NAND4_in[0] ,
         \SB2_2_19/Component_Function_3/NAND4_in[3] ,
         \SB2_2_19/Component_Function_3/NAND4_in[1] ,
         \SB2_2_19/Component_Function_3/NAND4_in[0] ,
         \SB2_2_19/Component_Function_4/NAND4_in[3] ,
         \SB2_2_19/Component_Function_4/NAND4_in[2] ,
         \SB2_2_19/Component_Function_4/NAND4_in[1] ,
         \SB2_2_19/Component_Function_4/NAND4_in[0] ,
         \SB2_2_20/Component_Function_2/NAND4_in[2] ,
         \SB2_2_20/Component_Function_3/NAND4_in[2] ,
         \SB2_2_20/Component_Function_3/NAND4_in[1] ,
         \SB2_2_20/Component_Function_3/NAND4_in[0] ,
         \SB2_2_20/Component_Function_4/NAND4_in[3] ,
         \SB2_2_20/Component_Function_4/NAND4_in[1] ,
         \SB2_2_20/Component_Function_4/NAND4_in[0] ,
         \SB2_2_21/Component_Function_2/NAND4_in[0] ,
         \SB2_2_21/Component_Function_3/NAND4_in[3] ,
         \SB2_2_21/Component_Function_3/NAND4_in[1] ,
         \SB2_2_21/Component_Function_3/NAND4_in[0] ,
         \SB2_2_21/Component_Function_4/NAND4_in[3] ,
         \SB2_2_21/Component_Function_4/NAND4_in[1] ,
         \SB2_2_21/Component_Function_4/NAND4_in[0] ,
         \SB2_2_22/Component_Function_2/NAND4_in[3] ,
         \SB2_2_22/Component_Function_2/NAND4_in[0] ,
         \SB2_2_22/Component_Function_3/NAND4_in[3] ,
         \SB2_2_22/Component_Function_3/NAND4_in[2] ,
         \SB2_2_22/Component_Function_3/NAND4_in[1] ,
         \SB2_2_22/Component_Function_3/NAND4_in[0] ,
         \SB2_2_22/Component_Function_4/NAND4_in[3] ,
         \SB2_2_22/Component_Function_4/NAND4_in[1] ,
         \SB2_2_22/Component_Function_4/NAND4_in[0] ,
         \SB2_2_23/Component_Function_2/NAND4_in[2] ,
         \SB2_2_23/Component_Function_2/NAND4_in[0] ,
         \SB2_2_23/Component_Function_3/NAND4_in[3] ,
         \SB2_2_23/Component_Function_3/NAND4_in[1] ,
         \SB2_2_23/Component_Function_3/NAND4_in[0] ,
         \SB2_2_23/Component_Function_4/NAND4_in[2] ,
         \SB2_2_23/Component_Function_4/NAND4_in[1] ,
         \SB2_2_23/Component_Function_4/NAND4_in[0] ,
         \SB2_2_24/Component_Function_2/NAND4_in[3] ,
         \SB2_2_24/Component_Function_2/NAND4_in[2] ,
         \SB2_2_24/Component_Function_2/NAND4_in[1] ,
         \SB2_2_24/Component_Function_2/NAND4_in[0] ,
         \SB2_2_24/Component_Function_3/NAND4_in[3] ,
         \SB2_2_24/Component_Function_3/NAND4_in[1] ,
         \SB2_2_24/Component_Function_4/NAND4_in[3] ,
         \SB2_2_24/Component_Function_4/NAND4_in[1] ,
         \SB2_2_24/Component_Function_4/NAND4_in[0] ,
         \SB2_2_25/Component_Function_2/NAND4_in[2] ,
         \SB2_2_25/Component_Function_2/NAND4_in[1] ,
         \SB2_2_25/Component_Function_2/NAND4_in[0] ,
         \SB2_2_25/Component_Function_3/NAND4_in[3] ,
         \SB2_2_25/Component_Function_3/NAND4_in[0] ,
         \SB2_2_25/Component_Function_4/NAND4_in[3] ,
         \SB2_2_25/Component_Function_4/NAND4_in[2] ,
         \SB2_2_25/Component_Function_4/NAND4_in[1] ,
         \SB2_2_25/Component_Function_4/NAND4_in[0] ,
         \SB2_2_26/Component_Function_2/NAND4_in[2] ,
         \SB2_2_26/Component_Function_2/NAND4_in[1] ,
         \SB2_2_26/Component_Function_2/NAND4_in[0] ,
         \SB2_2_26/Component_Function_3/NAND4_in[2] ,
         \SB2_2_26/Component_Function_3/NAND4_in[0] ,
         \SB2_2_26/Component_Function_4/NAND4_in[2] ,
         \SB2_2_26/Component_Function_4/NAND4_in[1] ,
         \SB2_2_26/Component_Function_4/NAND4_in[0] ,
         \SB2_2_27/Component_Function_2/NAND4_in[3] ,
         \SB2_2_27/Component_Function_3/NAND4_in[2] ,
         \SB2_2_27/Component_Function_3/NAND4_in[1] ,
         \SB2_2_27/Component_Function_3/NAND4_in[0] ,
         \SB2_2_27/Component_Function_4/NAND4_in[3] ,
         \SB2_2_27/Component_Function_4/NAND4_in[2] ,
         \SB2_2_27/Component_Function_4/NAND4_in[1] ,
         \SB2_2_27/Component_Function_4/NAND4_in[0] ,
         \SB2_2_28/Component_Function_2/NAND4_in[2] ,
         \SB2_2_28/Component_Function_2/NAND4_in[1] ,
         \SB2_2_28/Component_Function_2/NAND4_in[0] ,
         \SB2_2_28/Component_Function_3/NAND4_in[3] ,
         \SB2_2_28/Component_Function_3/NAND4_in[0] ,
         \SB2_2_28/Component_Function_4/NAND4_in[3] ,
         \SB2_2_28/Component_Function_4/NAND4_in[0] ,
         \SB2_2_29/Component_Function_2/NAND4_in[0] ,
         \SB2_2_29/Component_Function_3/NAND4_in[2] ,
         \SB2_2_29/Component_Function_3/NAND4_in[1] ,
         \SB2_2_29/Component_Function_3/NAND4_in[0] ,
         \SB2_2_29/Component_Function_4/NAND4_in[3] ,
         \SB2_2_29/Component_Function_4/NAND4_in[0] ,
         \SB2_2_30/Component_Function_2/NAND4_in[2] ,
         \SB2_2_30/Component_Function_2/NAND4_in[1] ,
         \SB2_2_30/Component_Function_2/NAND4_in[0] ,
         \SB2_2_30/Component_Function_3/NAND4_in[3] ,
         \SB2_2_30/Component_Function_3/NAND4_in[1] ,
         \SB2_2_30/Component_Function_3/NAND4_in[0] ,
         \SB2_2_30/Component_Function_4/NAND4_in[3] ,
         \SB2_2_30/Component_Function_4/NAND4_in[1] ,
         \SB2_2_30/Component_Function_4/NAND4_in[0] ,
         \SB2_2_31/Component_Function_2/NAND4_in[1] ,
         \SB2_2_31/Component_Function_2/NAND4_in[0] ,
         \SB2_2_31/Component_Function_3/NAND4_in[2] ,
         \SB2_2_31/Component_Function_3/NAND4_in[1] ,
         \SB2_2_31/Component_Function_4/NAND4_in[2] ,
         \SB2_2_31/Component_Function_4/NAND4_in[1] ,
         \SB2_2_31/Component_Function_4/NAND4_in[0] ,
         \SB1_3_0/Component_Function_2/NAND4_in[0] ,
         \SB1_3_0/Component_Function_3/NAND4_in[2] ,
         \SB1_3_0/Component_Function_3/NAND4_in[0] ,
         \SB1_3_0/Component_Function_4/NAND4_in[3] ,
         \SB1_3_0/Component_Function_4/NAND4_in[2] ,
         \SB1_3_0/Component_Function_4/NAND4_in[1] ,
         \SB1_3_0/Component_Function_4/NAND4_in[0] ,
         \SB1_3_1/Component_Function_2/NAND4_in[1] ,
         \SB1_3_1/Component_Function_2/NAND4_in[0] ,
         \SB1_3_1/Component_Function_3/NAND4_in[3] ,
         \SB1_3_1/Component_Function_3/NAND4_in[2] ,
         \SB1_3_1/Component_Function_3/NAND4_in[1] ,
         \SB1_3_1/Component_Function_3/NAND4_in[0] ,
         \SB1_3_1/Component_Function_4/NAND4_in[3] ,
         \SB1_3_1/Component_Function_4/NAND4_in[1] ,
         \SB1_3_1/Component_Function_4/NAND4_in[0] ,
         \SB1_3_2/Component_Function_2/NAND4_in[2] ,
         \SB1_3_2/Component_Function_2/NAND4_in[1] ,
         \SB1_3_2/Component_Function_2/NAND4_in[0] ,
         \SB1_3_2/Component_Function_3/NAND4_in[0] ,
         \SB1_3_2/Component_Function_4/NAND4_in[3] ,
         \SB1_3_2/Component_Function_4/NAND4_in[1] ,
         \SB1_3_2/Component_Function_4/NAND4_in[0] ,
         \SB1_3_3/Component_Function_2/NAND4_in[3] ,
         \SB1_3_3/Component_Function_2/NAND4_in[2] ,
         \SB1_3_3/Component_Function_3/NAND4_in[3] ,
         \SB1_3_3/Component_Function_3/NAND4_in[2] ,
         \SB1_3_3/Component_Function_3/NAND4_in[1] ,
         \SB1_3_3/Component_Function_3/NAND4_in[0] ,
         \SB1_3_3/Component_Function_4/NAND4_in[2] ,
         \SB1_3_3/Component_Function_4/NAND4_in[1] ,
         \SB1_3_3/Component_Function_4/NAND4_in[0] ,
         \SB1_3_4/Component_Function_2/NAND4_in[1] ,
         \SB1_3_4/Component_Function_2/NAND4_in[0] ,
         \SB1_3_4/Component_Function_3/NAND4_in[3] ,
         \SB1_3_4/Component_Function_3/NAND4_in[0] ,
         \SB1_3_4/Component_Function_4/NAND4_in[1] ,
         \SB1_3_5/Component_Function_2/NAND4_in[3] ,
         \SB1_3_5/Component_Function_2/NAND4_in[2] ,
         \SB1_3_5/Component_Function_2/NAND4_in[1] ,
         \SB1_3_5/Component_Function_2/NAND4_in[0] ,
         \SB1_3_5/Component_Function_3/NAND4_in[2] ,
         \SB1_3_5/Component_Function_3/NAND4_in[1] ,
         \SB1_3_5/Component_Function_3/NAND4_in[0] ,
         \SB1_3_5/Component_Function_4/NAND4_in[3] ,
         \SB1_3_5/Component_Function_4/NAND4_in[2] ,
         \SB1_3_5/Component_Function_4/NAND4_in[1] ,
         \SB1_3_5/Component_Function_4/NAND4_in[0] ,
         \SB1_3_6/Component_Function_2/NAND4_in[1] ,
         \SB1_3_6/Component_Function_3/NAND4_in[1] ,
         \SB1_3_6/Component_Function_3/NAND4_in[0] ,
         \SB1_3_6/Component_Function_4/NAND4_in[3] ,
         \SB1_3_6/Component_Function_4/NAND4_in[1] ,
         \SB1_3_7/Component_Function_2/NAND4_in[2] ,
         \SB1_3_7/Component_Function_2/NAND4_in[1] ,
         \SB1_3_7/Component_Function_2/NAND4_in[0] ,
         \SB1_3_7/Component_Function_3/NAND4_in[1] ,
         \SB1_3_7/Component_Function_3/NAND4_in[0] ,
         \SB1_3_7/Component_Function_4/NAND4_in[2] ,
         \SB1_3_7/Component_Function_4/NAND4_in[1] ,
         \SB1_3_7/Component_Function_4/NAND4_in[0] ,
         \SB1_3_8/Component_Function_2/NAND4_in[2] ,
         \SB1_3_8/Component_Function_2/NAND4_in[1] ,
         \SB1_3_8/Component_Function_2/NAND4_in[0] ,
         \SB1_3_8/Component_Function_3/NAND4_in[3] ,
         \SB1_3_8/Component_Function_3/NAND4_in[1] ,
         \SB1_3_8/Component_Function_3/NAND4_in[0] ,
         \SB1_3_8/Component_Function_4/NAND4_in[3] ,
         \SB1_3_9/Component_Function_2/NAND4_in[3] ,
         \SB1_3_9/Component_Function_2/NAND4_in[2] ,
         \SB1_3_9/Component_Function_2/NAND4_in[1] ,
         \SB1_3_9/Component_Function_2/NAND4_in[0] ,
         \SB1_3_9/Component_Function_3/NAND4_in[3] ,
         \SB1_3_9/Component_Function_3/NAND4_in[2] ,
         \SB1_3_9/Component_Function_3/NAND4_in[1] ,
         \SB1_3_9/Component_Function_3/NAND4_in[0] ,
         \SB1_3_9/Component_Function_4/NAND4_in[3] ,
         \SB1_3_9/Component_Function_4/NAND4_in[1] ,
         \SB1_3_9/Component_Function_4/NAND4_in[0] ,
         \SB1_3_10/Component_Function_2/NAND4_in[3] ,
         \SB1_3_10/Component_Function_2/NAND4_in[1] ,
         \SB1_3_10/Component_Function_2/NAND4_in[0] ,
         \SB1_3_10/Component_Function_3/NAND4_in[1] ,
         \SB1_3_10/Component_Function_3/NAND4_in[0] ,
         \SB1_3_10/Component_Function_4/NAND4_in[3] ,
         \SB1_3_10/Component_Function_4/NAND4_in[1] ,
         \SB1_3_10/Component_Function_4/NAND4_in[0] ,
         \SB1_3_11/Component_Function_2/NAND4_in[3] ,
         \SB1_3_11/Component_Function_2/NAND4_in[1] ,
         \SB1_3_11/Component_Function_3/NAND4_in[1] ,
         \SB1_3_12/Component_Function_2/NAND4_in[3] ,
         \SB1_3_12/Component_Function_2/NAND4_in[1] ,
         \SB1_3_12/Component_Function_2/NAND4_in[0] ,
         \SB1_3_12/Component_Function_3/NAND4_in[3] ,
         \SB1_3_12/Component_Function_3/NAND4_in[1] ,
         \SB1_3_12/Component_Function_3/NAND4_in[0] ,
         \SB1_3_12/Component_Function_4/NAND4_in[3] ,
         \SB1_3_12/Component_Function_4/NAND4_in[1] ,
         \SB1_3_13/Component_Function_2/NAND4_in[2] ,
         \SB1_3_13/Component_Function_2/NAND4_in[1] ,
         \SB1_3_13/Component_Function_3/NAND4_in[1] ,
         \SB1_3_13/Component_Function_3/NAND4_in[0] ,
         \SB1_3_13/Component_Function_4/NAND4_in[3] ,
         \SB1_3_13/Component_Function_4/NAND4_in[2] ,
         \SB1_3_13/Component_Function_4/NAND4_in[1] ,
         \SB1_3_14/Component_Function_2/NAND4_in[3] ,
         \SB1_3_14/Component_Function_2/NAND4_in[0] ,
         \SB1_3_14/Component_Function_3/NAND4_in[3] ,
         \SB1_3_14/Component_Function_3/NAND4_in[1] ,
         \SB1_3_14/Component_Function_4/NAND4_in[3] ,
         \SB1_3_14/Component_Function_4/NAND4_in[1] ,
         \SB1_3_15/Component_Function_2/NAND4_in[3] ,
         \SB1_3_15/Component_Function_2/NAND4_in[2] ,
         \SB1_3_15/Component_Function_2/NAND4_in[1] ,
         \SB1_3_15/Component_Function_2/NAND4_in[0] ,
         \SB1_3_15/Component_Function_3/NAND4_in[2] ,
         \SB1_3_15/Component_Function_3/NAND4_in[1] ,
         \SB1_3_15/Component_Function_4/NAND4_in[2] ,
         \SB1_3_15/Component_Function_4/NAND4_in[1] ,
         \SB1_3_15/Component_Function_4/NAND4_in[0] ,
         \SB1_3_16/Component_Function_2/NAND4_in[1] ,
         \SB1_3_16/Component_Function_3/NAND4_in[1] ,
         \SB1_3_16/Component_Function_4/NAND4_in[3] ,
         \SB1_3_16/Component_Function_4/NAND4_in[2] ,
         \SB1_3_16/Component_Function_4/NAND4_in[1] ,
         \SB1_3_17/Component_Function_2/NAND4_in[2] ,
         \SB1_3_17/Component_Function_2/NAND4_in[1] ,
         \SB1_3_17/Component_Function_3/NAND4_in[3] ,
         \SB1_3_17/Component_Function_3/NAND4_in[2] ,
         \SB1_3_17/Component_Function_4/NAND4_in[2] ,
         \SB1_3_17/Component_Function_4/NAND4_in[1] ,
         \SB1_3_17/Component_Function_4/NAND4_in[0] ,
         \SB1_3_18/Component_Function_2/NAND4_in[2] ,
         \SB1_3_18/Component_Function_2/NAND4_in[1] ,
         \SB1_3_18/Component_Function_2/NAND4_in[0] ,
         \SB1_3_18/Component_Function_3/NAND4_in[1] ,
         \SB1_3_18/Component_Function_3/NAND4_in[0] ,
         \SB1_3_18/Component_Function_4/NAND4_in[2] ,
         \SB1_3_18/Component_Function_4/NAND4_in[1] ,
         \SB1_3_18/Component_Function_4/NAND4_in[0] ,
         \SB1_3_19/Component_Function_2/NAND4_in[3] ,
         \SB1_3_19/Component_Function_2/NAND4_in[0] ,
         \SB1_3_19/Component_Function_3/NAND4_in[2] ,
         \SB1_3_19/Component_Function_3/NAND4_in[1] ,
         \SB1_3_19/Component_Function_3/NAND4_in[0] ,
         \SB1_3_19/Component_Function_4/NAND4_in[3] ,
         \SB1_3_19/Component_Function_4/NAND4_in[2] ,
         \SB1_3_19/Component_Function_4/NAND4_in[1] ,
         \SB1_3_19/Component_Function_4/NAND4_in[0] ,
         \SB1_3_20/Component_Function_2/NAND4_in[3] ,
         \SB1_3_20/Component_Function_2/NAND4_in[1] ,
         \SB1_3_20/Component_Function_2/NAND4_in[0] ,
         \SB1_3_20/Component_Function_3/NAND4_in[3] ,
         \SB1_3_20/Component_Function_3/NAND4_in[2] ,
         \SB1_3_20/Component_Function_3/NAND4_in[0] ,
         \SB1_3_20/Component_Function_4/NAND4_in[3] ,
         \SB1_3_20/Component_Function_4/NAND4_in[2] ,
         \SB1_3_20/Component_Function_4/NAND4_in[0] ,
         \SB1_3_21/Component_Function_2/NAND4_in[2] ,
         \SB1_3_21/Component_Function_2/NAND4_in[1] ,
         \SB1_3_21/Component_Function_2/NAND4_in[0] ,
         \SB1_3_21/Component_Function_3/NAND4_in[3] ,
         \SB1_3_21/Component_Function_3/NAND4_in[2] ,
         \SB1_3_21/Component_Function_3/NAND4_in[0] ,
         \SB1_3_21/Component_Function_4/NAND4_in[3] ,
         \SB1_3_21/Component_Function_4/NAND4_in[1] ,
         \SB1_3_22/Component_Function_2/NAND4_in[3] ,
         \SB1_3_22/Component_Function_2/NAND4_in[1] ,
         \SB1_3_22/Component_Function_3/NAND4_in[2] ,
         \SB1_3_22/Component_Function_3/NAND4_in[0] ,
         \SB1_3_22/Component_Function_4/NAND4_in[2] ,
         \SB1_3_22/Component_Function_4/NAND4_in[1] ,
         \SB1_3_22/Component_Function_4/NAND4_in[0] ,
         \SB1_3_23/Component_Function_2/NAND4_in[3] ,
         \SB1_3_23/Component_Function_2/NAND4_in[2] ,
         \SB1_3_23/Component_Function_2/NAND4_in[1] ,
         \SB1_3_23/Component_Function_3/NAND4_in[1] ,
         \SB1_3_23/Component_Function_3/NAND4_in[0] ,
         \SB1_3_23/Component_Function_4/NAND4_in[3] ,
         \SB1_3_23/Component_Function_4/NAND4_in[1] ,
         \SB1_3_24/Component_Function_2/NAND4_in[1] ,
         \SB1_3_24/Component_Function_2/NAND4_in[0] ,
         \SB1_3_24/Component_Function_3/NAND4_in[3] ,
         \SB1_3_24/Component_Function_3/NAND4_in[2] ,
         \SB1_3_24/Component_Function_3/NAND4_in[1] ,
         \SB1_3_24/Component_Function_3/NAND4_in[0] ,
         \SB1_3_24/Component_Function_4/NAND4_in[3] ,
         \SB1_3_24/Component_Function_4/NAND4_in[1] ,
         \SB1_3_24/Component_Function_4/NAND4_in[0] ,
         \SB1_3_25/Component_Function_2/NAND4_in[2] ,
         \SB1_3_25/Component_Function_2/NAND4_in[1] ,
         \SB1_3_25/Component_Function_2/NAND4_in[0] ,
         \SB1_3_25/Component_Function_3/NAND4_in[2] ,
         \SB1_3_25/Component_Function_3/NAND4_in[1] ,
         \SB1_3_25/Component_Function_3/NAND4_in[0] ,
         \SB1_3_25/Component_Function_4/NAND4_in[3] ,
         \SB1_3_25/Component_Function_4/NAND4_in[2] ,
         \SB1_3_25/Component_Function_4/NAND4_in[1] ,
         \SB1_3_25/Component_Function_4/NAND4_in[0] ,
         \SB1_3_26/Component_Function_2/NAND4_in[3] ,
         \SB1_3_26/Component_Function_2/NAND4_in[1] ,
         \SB1_3_26/Component_Function_2/NAND4_in[0] ,
         \SB1_3_26/Component_Function_3/NAND4_in[2] ,
         \SB1_3_26/Component_Function_3/NAND4_in[0] ,
         \SB1_3_26/Component_Function_4/NAND4_in[3] ,
         \SB1_3_26/Component_Function_4/NAND4_in[1] ,
         \SB1_3_26/Component_Function_4/NAND4_in[0] ,
         \SB1_3_27/Component_Function_2/NAND4_in[1] ,
         \SB1_3_27/Component_Function_2/NAND4_in[0] ,
         \SB1_3_27/Component_Function_3/NAND4_in[0] ,
         \SB1_3_28/Component_Function_2/NAND4_in[2] ,
         \SB1_3_28/Component_Function_2/NAND4_in[0] ,
         \SB1_3_28/Component_Function_3/NAND4_in[2] ,
         \SB1_3_28/Component_Function_3/NAND4_in[1] ,
         \SB1_3_28/Component_Function_3/NAND4_in[0] ,
         \SB1_3_28/Component_Function_4/NAND4_in[3] ,
         \SB1_3_28/Component_Function_4/NAND4_in[2] ,
         \SB1_3_28/Component_Function_4/NAND4_in[1] ,
         \SB1_3_28/Component_Function_4/NAND4_in[0] ,
         \SB1_3_29/Component_Function_2/NAND4_in[2] ,
         \SB1_3_29/Component_Function_2/NAND4_in[1] ,
         \SB1_3_29/Component_Function_2/NAND4_in[0] ,
         \SB1_3_29/Component_Function_3/NAND4_in[1] ,
         \SB1_3_29/Component_Function_3/NAND4_in[0] ,
         \SB1_3_29/Component_Function_4/NAND4_in[2] ,
         \SB1_3_29/Component_Function_4/NAND4_in[1] ,
         \SB1_3_30/Component_Function_2/NAND4_in[3] ,
         \SB1_3_30/Component_Function_2/NAND4_in[2] ,
         \SB1_3_30/Component_Function_2/NAND4_in[1] ,
         \SB1_3_30/Component_Function_3/NAND4_in[3] ,
         \SB1_3_30/Component_Function_3/NAND4_in[1] ,
         \SB1_3_30/Component_Function_3/NAND4_in[0] ,
         \SB1_3_30/Component_Function_4/NAND4_in[1] ,
         \SB1_3_30/Component_Function_4/NAND4_in[0] ,
         \SB1_3_31/Component_Function_2/NAND4_in[3] ,
         \SB1_3_31/Component_Function_2/NAND4_in[2] ,
         \SB1_3_31/Component_Function_3/NAND4_in[3] ,
         \SB1_3_31/Component_Function_3/NAND4_in[2] ,
         \SB1_3_31/Component_Function_3/NAND4_in[1] ,
         \SB1_3_31/Component_Function_3/NAND4_in[0] ,
         \SB1_3_31/Component_Function_4/NAND4_in[0] ,
         \SB2_3_0/Component_Function_2/NAND4_in[2] ,
         \SB2_3_0/Component_Function_2/NAND4_in[1] ,
         \SB2_3_0/Component_Function_3/NAND4_in[3] ,
         \SB2_3_0/Component_Function_3/NAND4_in[2] ,
         \SB2_3_0/Component_Function_3/NAND4_in[1] ,
         \SB2_3_0/Component_Function_3/NAND4_in[0] ,
         \SB2_3_0/Component_Function_4/NAND4_in[3] ,
         \SB2_3_1/Component_Function_2/NAND4_in[2] ,
         \SB2_3_1/Component_Function_2/NAND4_in[0] ,
         \SB2_3_1/Component_Function_3/NAND4_in[3] ,
         \SB2_3_1/Component_Function_3/NAND4_in[2] ,
         \SB2_3_1/Component_Function_3/NAND4_in[0] ,
         \SB2_3_1/Component_Function_4/NAND4_in[2] ,
         \SB2_3_1/Component_Function_4/NAND4_in[1] ,
         \SB2_3_1/Component_Function_4/NAND4_in[0] ,
         \SB2_3_2/Component_Function_2/NAND4_in[0] ,
         \SB2_3_2/Component_Function_3/NAND4_in[2] ,
         \SB2_3_2/Component_Function_3/NAND4_in[1] ,
         \SB2_3_2/Component_Function_3/NAND4_in[0] ,
         \SB2_3_2/Component_Function_4/NAND4_in[3] ,
         \SB2_3_2/Component_Function_4/NAND4_in[1] ,
         \SB2_3_2/Component_Function_4/NAND4_in[0] ,
         \SB2_3_3/Component_Function_2/NAND4_in[1] ,
         \SB2_3_3/Component_Function_2/NAND4_in[0] ,
         \SB2_3_3/Component_Function_3/NAND4_in[2] ,
         \SB2_3_3/Component_Function_3/NAND4_in[1] ,
         \SB2_3_3/Component_Function_3/NAND4_in[0] ,
         \SB2_3_3/Component_Function_4/NAND4_in[3] ,
         \SB2_3_3/Component_Function_4/NAND4_in[2] ,
         \SB2_3_3/Component_Function_4/NAND4_in[1] ,
         \SB2_3_4/Component_Function_2/NAND4_in[2] ,
         \SB2_3_4/Component_Function_2/NAND4_in[1] ,
         \SB2_3_4/Component_Function_2/NAND4_in[0] ,
         \SB2_3_4/Component_Function_3/NAND4_in[3] ,
         \SB2_3_4/Component_Function_3/NAND4_in[2] ,
         \SB2_3_4/Component_Function_3/NAND4_in[0] ,
         \SB2_3_4/Component_Function_4/NAND4_in[3] ,
         \SB2_3_4/Component_Function_4/NAND4_in[1] ,
         \SB2_3_4/Component_Function_4/NAND4_in[0] ,
         \SB2_3_5/Component_Function_2/NAND4_in[2] ,
         \SB2_3_5/Component_Function_2/NAND4_in[0] ,
         \SB2_3_5/Component_Function_3/NAND4_in[3] ,
         \SB2_3_5/Component_Function_3/NAND4_in[2] ,
         \SB2_3_5/Component_Function_3/NAND4_in[1] ,
         \SB2_3_5/Component_Function_3/NAND4_in[0] ,
         \SB2_3_5/Component_Function_4/NAND4_in[1] ,
         \SB2_3_5/Component_Function_4/NAND4_in[0] ,
         \SB2_3_6/Component_Function_2/NAND4_in[2] ,
         \SB2_3_6/Component_Function_2/NAND4_in[1] ,
         \SB2_3_6/Component_Function_2/NAND4_in[0] ,
         \SB2_3_6/Component_Function_3/NAND4_in[3] ,
         \SB2_3_6/Component_Function_3/NAND4_in[1] ,
         \SB2_3_6/Component_Function_3/NAND4_in[0] ,
         \SB2_3_6/Component_Function_4/NAND4_in[3] ,
         \SB2_3_6/Component_Function_4/NAND4_in[1] ,
         \SB2_3_6/Component_Function_4/NAND4_in[0] ,
         \SB2_3_7/Component_Function_2/NAND4_in[2] ,
         \SB2_3_7/Component_Function_2/NAND4_in[0] ,
         \SB2_3_7/Component_Function_3/NAND4_in[3] ,
         \SB2_3_7/Component_Function_3/NAND4_in[2] ,
         \SB2_3_7/Component_Function_3/NAND4_in[0] ,
         \SB2_3_7/Component_Function_4/NAND4_in[3] ,
         \SB2_3_7/Component_Function_4/NAND4_in[1] ,
         \SB2_3_7/Component_Function_4/NAND4_in[0] ,
         \SB2_3_8/Component_Function_2/NAND4_in[2] ,
         \SB2_3_8/Component_Function_2/NAND4_in[0] ,
         \SB2_3_8/Component_Function_3/NAND4_in[2] ,
         \SB2_3_8/Component_Function_3/NAND4_in[1] ,
         \SB2_3_8/Component_Function_3/NAND4_in[0] ,
         \SB2_3_8/Component_Function_4/NAND4_in[3] ,
         \SB2_3_8/Component_Function_4/NAND4_in[2] ,
         \SB2_3_8/Component_Function_4/NAND4_in[1] ,
         \SB2_3_8/Component_Function_4/NAND4_in[0] ,
         \SB2_3_9/Component_Function_2/NAND4_in[2] ,
         \SB2_3_9/Component_Function_2/NAND4_in[1] ,
         \SB2_3_9/Component_Function_2/NAND4_in[0] ,
         \SB2_3_9/Component_Function_3/NAND4_in[3] ,
         \SB2_3_9/Component_Function_3/NAND4_in[1] ,
         \SB2_3_9/Component_Function_3/NAND4_in[0] ,
         \SB2_3_9/Component_Function_4/NAND4_in[3] ,
         \SB2_3_9/Component_Function_4/NAND4_in[1] ,
         \SB2_3_10/Component_Function_2/NAND4_in[2] ,
         \SB2_3_10/Component_Function_2/NAND4_in[0] ,
         \SB2_3_10/Component_Function_3/NAND4_in[3] ,
         \SB2_3_10/Component_Function_3/NAND4_in[0] ,
         \SB2_3_10/Component_Function_4/NAND4_in[3] ,
         \SB2_3_10/Component_Function_4/NAND4_in[0] ,
         \SB2_3_11/Component_Function_2/NAND4_in[2] ,
         \SB2_3_11/Component_Function_3/NAND4_in[3] ,
         \SB2_3_11/Component_Function_4/NAND4_in[1] ,
         \SB2_3_11/Component_Function_4/NAND4_in[0] ,
         \SB2_3_12/Component_Function_2/NAND4_in[3] ,
         \SB2_3_12/Component_Function_2/NAND4_in[1] ,
         \SB2_3_12/Component_Function_2/NAND4_in[0] ,
         \SB2_3_12/Component_Function_3/NAND4_in[3] ,
         \SB2_3_12/Component_Function_3/NAND4_in[2] ,
         \SB2_3_12/Component_Function_3/NAND4_in[1] ,
         \SB2_3_12/Component_Function_3/NAND4_in[0] ,
         \SB2_3_12/Component_Function_4/NAND4_in[3] ,
         \SB2_3_12/Component_Function_4/NAND4_in[2] ,
         \SB2_3_12/Component_Function_4/NAND4_in[1] ,
         \SB2_3_12/Component_Function_4/NAND4_in[0] ,
         \SB2_3_13/Component_Function_2/NAND4_in[2] ,
         \SB2_3_13/Component_Function_2/NAND4_in[0] ,
         \SB2_3_13/Component_Function_3/NAND4_in[3] ,
         \SB2_3_13/Component_Function_3/NAND4_in[2] ,
         \SB2_3_13/Component_Function_4/NAND4_in[3] ,
         \SB2_3_13/Component_Function_4/NAND4_in[2] ,
         \SB2_3_13/Component_Function_4/NAND4_in[1] ,
         \SB2_3_13/Component_Function_4/NAND4_in[0] ,
         \SB2_3_14/Component_Function_2/NAND4_in[2] ,
         \SB2_3_14/Component_Function_2/NAND4_in[0] ,
         \SB2_3_14/Component_Function_3/NAND4_in[3] ,
         \SB2_3_14/Component_Function_3/NAND4_in[1] ,
         \SB2_3_14/Component_Function_3/NAND4_in[0] ,
         \SB2_3_14/Component_Function_4/NAND4_in[3] ,
         \SB2_3_14/Component_Function_4/NAND4_in[2] ,
         \SB2_3_14/Component_Function_4/NAND4_in[1] ,
         \SB2_3_14/Component_Function_4/NAND4_in[0] ,
         \SB2_3_15/Component_Function_2/NAND4_in[2] ,
         \SB2_3_15/Component_Function_2/NAND4_in[0] ,
         \SB2_3_15/Component_Function_3/NAND4_in[3] ,
         \SB2_3_15/Component_Function_3/NAND4_in[0] ,
         \SB2_3_15/Component_Function_4/NAND4_in[3] ,
         \SB2_3_15/Component_Function_4/NAND4_in[1] ,
         \SB2_3_15/Component_Function_4/NAND4_in[0] ,
         \SB2_3_16/Component_Function_2/NAND4_in[2] ,
         \SB2_3_16/Component_Function_2/NAND4_in[1] ,
         \SB2_3_16/Component_Function_2/NAND4_in[0] ,
         \SB2_3_16/Component_Function_3/NAND4_in[3] ,
         \SB2_3_16/Component_Function_3/NAND4_in[2] ,
         \SB2_3_16/Component_Function_3/NAND4_in[0] ,
         \SB2_3_16/Component_Function_4/NAND4_in[3] ,
         \SB2_3_16/Component_Function_4/NAND4_in[2] ,
         \SB2_3_16/Component_Function_4/NAND4_in[1] ,
         \SB2_3_16/Component_Function_4/NAND4_in[0] ,
         \SB2_3_17/Component_Function_2/NAND4_in[2] ,
         \SB2_3_17/Component_Function_2/NAND4_in[1] ,
         \SB2_3_17/Component_Function_2/NAND4_in[0] ,
         \SB2_3_17/Component_Function_3/NAND4_in[0] ,
         \SB2_3_17/Component_Function_4/NAND4_in[3] ,
         \SB2_3_17/Component_Function_4/NAND4_in[1] ,
         \SB2_3_17/Component_Function_4/NAND4_in[0] ,
         \SB2_3_18/Component_Function_2/NAND4_in[0] ,
         \SB2_3_18/Component_Function_3/NAND4_in[3] ,
         \SB2_3_18/Component_Function_3/NAND4_in[1] ,
         \SB2_3_18/Component_Function_3/NAND4_in[0] ,
         \SB2_3_18/Component_Function_4/NAND4_in[3] ,
         \SB2_3_18/Component_Function_4/NAND4_in[2] ,
         \SB2_3_18/Component_Function_4/NAND4_in[1] ,
         \SB2_3_18/Component_Function_4/NAND4_in[0] ,
         \SB2_3_19/Component_Function_2/NAND4_in[2] ,
         \SB2_3_19/Component_Function_2/NAND4_in[0] ,
         \SB2_3_19/Component_Function_3/NAND4_in[3] ,
         \SB2_3_19/Component_Function_3/NAND4_in[0] ,
         \SB2_3_19/Component_Function_4/NAND4_in[2] ,
         \SB2_3_19/Component_Function_4/NAND4_in[1] ,
         \SB2_3_19/Component_Function_4/NAND4_in[0] ,
         \SB2_3_20/Component_Function_2/NAND4_in[2] ,
         \SB2_3_20/Component_Function_2/NAND4_in[1] ,
         \SB2_3_20/Component_Function_2/NAND4_in[0] ,
         \SB2_3_20/Component_Function_3/NAND4_in[3] ,
         \SB2_3_20/Component_Function_3/NAND4_in[0] ,
         \SB2_3_20/Component_Function_4/NAND4_in[1] ,
         \SB2_3_20/Component_Function_4/NAND4_in[0] ,
         \SB2_3_21/Component_Function_2/NAND4_in[2] ,
         \SB2_3_21/Component_Function_2/NAND4_in[0] ,
         \SB2_3_21/Component_Function_3/NAND4_in[3] ,
         \SB2_3_21/Component_Function_3/NAND4_in[1] ,
         \SB2_3_21/Component_Function_3/NAND4_in[0] ,
         \SB2_3_21/Component_Function_4/NAND4_in[2] ,
         \SB2_3_21/Component_Function_4/NAND4_in[1] ,
         \SB2_3_21/Component_Function_4/NAND4_in[0] ,
         \SB2_3_22/Component_Function_2/NAND4_in[2] ,
         \SB2_3_22/Component_Function_2/NAND4_in[1] ,
         \SB2_3_22/Component_Function_2/NAND4_in[0] ,
         \SB2_3_22/Component_Function_3/NAND4_in[3] ,
         \SB2_3_22/Component_Function_3/NAND4_in[2] ,
         \SB2_3_22/Component_Function_3/NAND4_in[1] ,
         \SB2_3_22/Component_Function_3/NAND4_in[0] ,
         \SB2_3_22/Component_Function_4/NAND4_in[3] ,
         \SB2_3_22/Component_Function_4/NAND4_in[2] ,
         \SB2_3_22/Component_Function_4/NAND4_in[1] ,
         \SB2_3_22/Component_Function_4/NAND4_in[0] ,
         \SB2_3_23/Component_Function_2/NAND4_in[2] ,
         \SB2_3_23/Component_Function_2/NAND4_in[0] ,
         \SB2_3_23/Component_Function_3/NAND4_in[3] ,
         \SB2_3_23/Component_Function_4/NAND4_in[3] ,
         \SB2_3_23/Component_Function_4/NAND4_in[0] ,
         \SB2_3_24/Component_Function_2/NAND4_in[2] ,
         \SB2_3_24/Component_Function_2/NAND4_in[1] ,
         \SB2_3_24/Component_Function_2/NAND4_in[0] ,
         \SB2_3_24/Component_Function_3/NAND4_in[1] ,
         \SB2_3_24/Component_Function_3/NAND4_in[0] ,
         \SB2_3_24/Component_Function_4/NAND4_in[3] ,
         \SB2_3_24/Component_Function_4/NAND4_in[2] ,
         \SB2_3_24/Component_Function_4/NAND4_in[1] ,
         \SB2_3_24/Component_Function_4/NAND4_in[0] ,
         \SB2_3_25/Component_Function_2/NAND4_in[3] ,
         \SB2_3_25/Component_Function_2/NAND4_in[1] ,
         \SB2_3_25/Component_Function_2/NAND4_in[0] ,
         \SB2_3_25/Component_Function_3/NAND4_in[3] ,
         \SB2_3_25/Component_Function_3/NAND4_in[1] ,
         \SB2_3_25/Component_Function_3/NAND4_in[0] ,
         \SB2_3_25/Component_Function_4/NAND4_in[3] ,
         \SB2_3_25/Component_Function_4/NAND4_in[2] ,
         \SB2_3_25/Component_Function_4/NAND4_in[1] ,
         \SB2_3_25/Component_Function_4/NAND4_in[0] ,
         \SB2_3_26/Component_Function_2/NAND4_in[2] ,
         \SB2_3_26/Component_Function_2/NAND4_in[1] ,
         \SB2_3_26/Component_Function_2/NAND4_in[0] ,
         \SB2_3_26/Component_Function_3/NAND4_in[3] ,
         \SB2_3_26/Component_Function_3/NAND4_in[2] ,
         \SB2_3_26/Component_Function_3/NAND4_in[1] ,
         \SB2_3_26/Component_Function_3/NAND4_in[0] ,
         \SB2_3_26/Component_Function_4/NAND4_in[3] ,
         \SB2_3_26/Component_Function_4/NAND4_in[1] ,
         \SB2_3_26/Component_Function_4/NAND4_in[0] ,
         \SB2_3_27/Component_Function_2/NAND4_in[3] ,
         \SB2_3_27/Component_Function_2/NAND4_in[1] ,
         \SB2_3_27/Component_Function_2/NAND4_in[0] ,
         \SB2_3_27/Component_Function_3/NAND4_in[3] ,
         \SB2_3_27/Component_Function_3/NAND4_in[1] ,
         \SB2_3_27/Component_Function_4/NAND4_in[3] ,
         \SB2_3_27/Component_Function_4/NAND4_in[1] ,
         \SB2_3_27/Component_Function_4/NAND4_in[0] ,
         \SB2_3_28/Component_Function_2/NAND4_in[3] ,
         \SB2_3_28/Component_Function_2/NAND4_in[0] ,
         \SB2_3_28/Component_Function_3/NAND4_in[2] ,
         \SB2_3_28/Component_Function_3/NAND4_in[0] ,
         \SB2_3_28/Component_Function_4/NAND4_in[0] ,
         \SB2_3_29/Component_Function_2/NAND4_in[2] ,
         \SB2_3_29/Component_Function_2/NAND4_in[1] ,
         \SB2_3_29/Component_Function_2/NAND4_in[0] ,
         \SB2_3_29/Component_Function_3/NAND4_in[3] ,
         \SB2_3_29/Component_Function_4/NAND4_in[3] ,
         \SB2_3_29/Component_Function_4/NAND4_in[0] ,
         \SB2_3_30/Component_Function_2/NAND4_in[2] ,
         \SB2_3_30/Component_Function_2/NAND4_in[1] ,
         \SB2_3_30/Component_Function_2/NAND4_in[0] ,
         \SB2_3_30/Component_Function_3/NAND4_in[3] ,
         \SB2_3_30/Component_Function_3/NAND4_in[0] ,
         \SB2_3_30/Component_Function_4/NAND4_in[3] ,
         \SB2_3_30/Component_Function_4/NAND4_in[1] ,
         \SB2_3_30/Component_Function_4/NAND4_in[0] ,
         \SB2_3_31/Component_Function_2/NAND4_in[3] ,
         \SB2_3_31/Component_Function_2/NAND4_in[2] ,
         \SB2_3_31/Component_Function_2/NAND4_in[1] ,
         \SB2_3_31/Component_Function_2/NAND4_in[0] ,
         \SB2_3_31/Component_Function_3/NAND4_in[3] ,
         \SB2_3_31/Component_Function_3/NAND4_in[2] ,
         \SB2_3_31/Component_Function_3/NAND4_in[1] ,
         \SB2_3_31/Component_Function_3/NAND4_in[0] ,
         \SB2_3_31/Component_Function_4/NAND4_in[3] ,
         \SB2_3_31/Component_Function_4/NAND4_in[2] ,
         \SB2_3_31/Component_Function_4/NAND4_in[1] ,
         \SB2_3_31/Component_Function_4/NAND4_in[0] ,
         \SB1_4_0/Component_Function_2/NAND4_in[1] ,
         \SB1_4_0/Component_Function_2/NAND4_in[0] ,
         \SB1_4_0/Component_Function_3/NAND4_in[3] ,
         \SB1_4_0/Component_Function_4/NAND4_in[2] ,
         \SB1_4_0/Component_Function_4/NAND4_in[1] ,
         \SB1_4_0/Component_Function_4/NAND4_in[0] ,
         \SB1_4_1/Component_Function_2/NAND4_in[3] ,
         \SB1_4_1/Component_Function_2/NAND4_in[1] ,
         \SB1_4_1/Component_Function_2/NAND4_in[0] ,
         \SB1_4_1/Component_Function_3/NAND4_in[2] ,
         \SB1_4_1/Component_Function_3/NAND4_in[1] ,
         \SB1_4_1/Component_Function_3/NAND4_in[0] ,
         \SB1_4_1/Component_Function_4/NAND4_in[1] ,
         \SB1_4_1/Component_Function_4/NAND4_in[0] ,
         \SB1_4_2/Component_Function_2/NAND4_in[3] ,
         \SB1_4_2/Component_Function_2/NAND4_in[1] ,
         \SB1_4_2/Component_Function_2/NAND4_in[0] ,
         \SB1_4_2/Component_Function_3/NAND4_in[2] ,
         \SB1_4_2/Component_Function_3/NAND4_in[1] ,
         \SB1_4_2/Component_Function_3/NAND4_in[0] ,
         \SB1_4_3/Component_Function_2/NAND4_in[3] ,
         \SB1_4_3/Component_Function_2/NAND4_in[1] ,
         \SB1_4_3/Component_Function_3/NAND4_in[1] ,
         \SB1_4_3/Component_Function_4/NAND4_in[2] ,
         \SB1_4_3/Component_Function_4/NAND4_in[1] ,
         \SB1_4_3/Component_Function_4/NAND4_in[0] ,
         \SB1_4_4/Component_Function_2/NAND4_in[2] ,
         \SB1_4_4/Component_Function_2/NAND4_in[0] ,
         \SB1_4_4/Component_Function_3/NAND4_in[1] ,
         \SB1_4_4/Component_Function_3/NAND4_in[0] ,
         \SB1_4_4/Component_Function_4/NAND4_in[3] ,
         \SB1_4_4/Component_Function_4/NAND4_in[2] ,
         \SB1_4_4/Component_Function_4/NAND4_in[1] ,
         \SB1_4_4/Component_Function_4/NAND4_in[0] ,
         \SB1_4_5/Component_Function_2/NAND4_in[3] ,
         \SB1_4_5/Component_Function_2/NAND4_in[2] ,
         \SB1_4_5/Component_Function_2/NAND4_in[0] ,
         \SB1_4_5/Component_Function_3/NAND4_in[3] ,
         \SB1_4_5/Component_Function_3/NAND4_in[1] ,
         \SB1_4_5/Component_Function_3/NAND4_in[0] ,
         \SB1_4_5/Component_Function_4/NAND4_in[3] ,
         \SB1_4_5/Component_Function_4/NAND4_in[1] ,
         \SB1_4_5/Component_Function_4/NAND4_in[0] ,
         \SB1_4_6/Component_Function_3/NAND4_in[1] ,
         \SB1_4_6/Component_Function_3/NAND4_in[0] ,
         \SB1_4_6/Component_Function_4/NAND4_in[3] ,
         \SB1_4_6/Component_Function_4/NAND4_in[0] ,
         \SB1_4_7/Component_Function_2/NAND4_in[2] ,
         \SB1_4_7/Component_Function_2/NAND4_in[1] ,
         \SB1_4_7/Component_Function_3/NAND4_in[1] ,
         \SB1_4_7/Component_Function_4/NAND4_in[2] ,
         \SB1_4_7/Component_Function_4/NAND4_in[1] ,
         \SB1_4_7/Component_Function_4/NAND4_in[0] ,
         \SB1_4_8/Component_Function_2/NAND4_in[3] ,
         \SB1_4_8/Component_Function_2/NAND4_in[1] ,
         \SB1_4_8/Component_Function_3/NAND4_in[2] ,
         \SB1_4_8/Component_Function_3/NAND4_in[1] ,
         \SB1_4_8/Component_Function_4/NAND4_in[3] ,
         \SB1_4_8/Component_Function_4/NAND4_in[2] ,
         \SB1_4_8/Component_Function_4/NAND4_in[1] ,
         \SB1_4_8/Component_Function_4/NAND4_in[0] ,
         \SB1_4_9/Component_Function_2/NAND4_in[2] ,
         \SB1_4_9/Component_Function_2/NAND4_in[0] ,
         \SB1_4_9/Component_Function_3/NAND4_in[2] ,
         \SB1_4_9/Component_Function_3/NAND4_in[1] ,
         \SB1_4_9/Component_Function_4/NAND4_in[2] ,
         \SB1_4_9/Component_Function_4/NAND4_in[0] ,
         \SB1_4_10/Component_Function_2/NAND4_in[2] ,
         \SB1_4_10/Component_Function_2/NAND4_in[1] ,
         \SB1_4_10/Component_Function_2/NAND4_in[0] ,
         \SB1_4_10/Component_Function_3/NAND4_in[2] ,
         \SB1_4_10/Component_Function_3/NAND4_in[1] ,
         \SB1_4_10/Component_Function_3/NAND4_in[0] ,
         \SB1_4_10/Component_Function_4/NAND4_in[3] ,
         \SB1_4_10/Component_Function_4/NAND4_in[0] ,
         \SB1_4_11/Component_Function_2/NAND4_in[2] ,
         \SB1_4_11/Component_Function_2/NAND4_in[1] ,
         \SB1_4_11/Component_Function_2/NAND4_in[0] ,
         \SB1_4_11/Component_Function_3/NAND4_in[2] ,
         \SB1_4_11/Component_Function_3/NAND4_in[1] ,
         \SB1_4_11/Component_Function_3/NAND4_in[0] ,
         \SB1_4_11/Component_Function_4/NAND4_in[2] ,
         \SB1_4_11/Component_Function_4/NAND4_in[1] ,
         \SB1_4_11/Component_Function_4/NAND4_in[0] ,
         \SB1_4_12/Component_Function_2/NAND4_in[1] ,
         \SB1_4_12/Component_Function_2/NAND4_in[0] ,
         \SB1_4_12/Component_Function_3/NAND4_in[3] ,
         \SB1_4_12/Component_Function_3/NAND4_in[1] ,
         \SB1_4_12/Component_Function_3/NAND4_in[0] ,
         \SB1_4_12/Component_Function_4/NAND4_in[1] ,
         \SB1_4_13/Component_Function_2/NAND4_in[3] ,
         \SB1_4_13/Component_Function_2/NAND4_in[1] ,
         \SB1_4_13/Component_Function_3/NAND4_in[3] ,
         \SB1_4_13/Component_Function_3/NAND4_in[1] ,
         \SB1_4_13/Component_Function_3/NAND4_in[0] ,
         \SB1_4_13/Component_Function_4/NAND4_in[3] ,
         \SB1_4_13/Component_Function_4/NAND4_in[1] ,
         \SB1_4_13/Component_Function_4/NAND4_in[0] ,
         \SB1_4_14/Component_Function_2/NAND4_in[2] ,
         \SB1_4_14/Component_Function_2/NAND4_in[0] ,
         \SB1_4_14/Component_Function_3/NAND4_in[0] ,
         \SB1_4_14/Component_Function_4/NAND4_in[1] ,
         \SB1_4_14/Component_Function_4/NAND4_in[0] ,
         \SB1_4_15/Component_Function_2/NAND4_in[1] ,
         \SB1_4_15/Component_Function_3/NAND4_in[2] ,
         \SB1_4_15/Component_Function_3/NAND4_in[1] ,
         \SB1_4_15/Component_Function_4/NAND4_in[2] ,
         \SB1_4_15/Component_Function_4/NAND4_in[1] ,
         \SB1_4_15/Component_Function_4/NAND4_in[0] ,
         \SB1_4_16/Component_Function_2/NAND4_in[1] ,
         \SB1_4_16/Component_Function_2/NAND4_in[0] ,
         \SB1_4_16/Component_Function_3/NAND4_in[1] ,
         \SB1_4_16/Component_Function_4/NAND4_in[2] ,
         \SB1_4_16/Component_Function_4/NAND4_in[1] ,
         \SB1_4_16/Component_Function_4/NAND4_in[0] ,
         \SB1_4_17/Component_Function_2/NAND4_in[1] ,
         \SB1_4_17/Component_Function_2/NAND4_in[0] ,
         \SB1_4_17/Component_Function_3/NAND4_in[1] ,
         \SB1_4_17/Component_Function_4/NAND4_in[3] ,
         \SB1_4_17/Component_Function_4/NAND4_in[2] ,
         \SB1_4_17/Component_Function_4/NAND4_in[1] ,
         \SB1_4_17/Component_Function_4/NAND4_in[0] ,
         \SB1_4_18/Component_Function_2/NAND4_in[1] ,
         \SB1_4_18/Component_Function_2/NAND4_in[0] ,
         \SB1_4_18/Component_Function_3/NAND4_in[1] ,
         \SB1_4_18/Component_Function_4/NAND4_in[3] ,
         \SB1_4_18/Component_Function_4/NAND4_in[1] ,
         \SB1_4_18/Component_Function_4/NAND4_in[0] ,
         \SB1_4_19/Component_Function_2/NAND4_in[1] ,
         \SB1_4_19/Component_Function_3/NAND4_in[0] ,
         \SB1_4_19/Component_Function_4/NAND4_in[3] ,
         \SB1_4_19/Component_Function_4/NAND4_in[2] ,
         \SB1_4_19/Component_Function_4/NAND4_in[0] ,
         \SB1_4_20/Component_Function_2/NAND4_in[2] ,
         \SB1_4_20/Component_Function_3/NAND4_in[3] ,
         \SB1_4_20/Component_Function_3/NAND4_in[1] ,
         \SB1_4_20/Component_Function_3/NAND4_in[0] ,
         \SB1_4_20/Component_Function_4/NAND4_in[3] ,
         \SB1_4_20/Component_Function_4/NAND4_in[2] ,
         \SB1_4_20/Component_Function_4/NAND4_in[1] ,
         \SB1_4_20/Component_Function_4/NAND4_in[0] ,
         \SB1_4_21/Component_Function_2/NAND4_in[1] ,
         \SB1_4_21/Component_Function_3/NAND4_in[2] ,
         \SB1_4_21/Component_Function_3/NAND4_in[1] ,
         \SB1_4_21/Component_Function_3/NAND4_in[0] ,
         \SB1_4_21/Component_Function_4/NAND4_in[3] ,
         \SB1_4_21/Component_Function_4/NAND4_in[1] ,
         \SB1_4_22/Component_Function_2/NAND4_in[3] ,
         \SB1_4_22/Component_Function_2/NAND4_in[2] ,
         \SB1_4_22/Component_Function_2/NAND4_in[1] ,
         \SB1_4_22/Component_Function_2/NAND4_in[0] ,
         \SB1_4_22/Component_Function_3/NAND4_in[2] ,
         \SB1_4_22/Component_Function_3/NAND4_in[0] ,
         \SB1_4_22/Component_Function_4/NAND4_in[3] ,
         \SB1_4_22/Component_Function_4/NAND4_in[1] ,
         \SB1_4_22/Component_Function_4/NAND4_in[0] ,
         \SB1_4_23/Component_Function_2/NAND4_in[3] ,
         \SB1_4_23/Component_Function_2/NAND4_in[1] ,
         \SB1_4_23/Component_Function_2/NAND4_in[0] ,
         \SB1_4_23/Component_Function_3/NAND4_in[1] ,
         \SB1_4_23/Component_Function_3/NAND4_in[0] ,
         \SB1_4_23/Component_Function_4/NAND4_in[3] ,
         \SB1_4_23/Component_Function_4/NAND4_in[2] ,
         \SB1_4_23/Component_Function_4/NAND4_in[1] ,
         \SB1_4_23/Component_Function_4/NAND4_in[0] ,
         \SB1_4_24/Component_Function_2/NAND4_in[3] ,
         \SB1_4_24/Component_Function_2/NAND4_in[2] ,
         \SB1_4_24/Component_Function_2/NAND4_in[0] ,
         \SB1_4_24/Component_Function_3/NAND4_in[1] ,
         \SB1_4_24/Component_Function_3/NAND4_in[0] ,
         \SB1_4_24/Component_Function_4/NAND4_in[2] ,
         \SB1_4_25/Component_Function_2/NAND4_in[1] ,
         \SB1_4_25/Component_Function_3/NAND4_in[3] ,
         \SB1_4_25/Component_Function_3/NAND4_in[1] ,
         \SB1_4_25/Component_Function_4/NAND4_in[2] ,
         \SB1_4_25/Component_Function_4/NAND4_in[1] ,
         \SB1_4_26/Component_Function_2/NAND4_in[0] ,
         \SB1_4_26/Component_Function_3/NAND4_in[3] ,
         \SB1_4_26/Component_Function_3/NAND4_in[1] ,
         \SB1_4_26/Component_Function_3/NAND4_in[0] ,
         \SB1_4_26/Component_Function_4/NAND4_in[3] ,
         \SB1_4_26/Component_Function_4/NAND4_in[2] ,
         \SB1_4_26/Component_Function_4/NAND4_in[1] ,
         \SB1_4_26/Component_Function_4/NAND4_in[0] ,
         \SB1_4_27/Component_Function_2/NAND4_in[2] ,
         \SB1_4_27/Component_Function_2/NAND4_in[1] ,
         \SB1_4_27/Component_Function_2/NAND4_in[0] ,
         \SB1_4_27/Component_Function_3/NAND4_in[2] ,
         \SB1_4_27/Component_Function_3/NAND4_in[1] ,
         \SB1_4_27/Component_Function_3/NAND4_in[0] ,
         \SB1_4_27/Component_Function_4/NAND4_in[2] ,
         \SB1_4_28/Component_Function_2/NAND4_in[2] ,
         \SB1_4_28/Component_Function_2/NAND4_in[1] ,
         \SB1_4_28/Component_Function_3/NAND4_in[2] ,
         \SB1_4_28/Component_Function_3/NAND4_in[0] ,
         \SB1_4_28/Component_Function_4/NAND4_in[2] ,
         \SB1_4_28/Component_Function_4/NAND4_in[1] ,
         \SB1_4_28/Component_Function_4/NAND4_in[0] ,
         \SB1_4_29/Component_Function_2/NAND4_in[3] ,
         \SB1_4_29/Component_Function_2/NAND4_in[1] ,
         \SB1_4_29/Component_Function_2/NAND4_in[0] ,
         \SB1_4_29/Component_Function_3/NAND4_in[3] ,
         \SB1_4_29/Component_Function_3/NAND4_in[1] ,
         \SB1_4_29/Component_Function_3/NAND4_in[0] ,
         \SB1_4_29/Component_Function_4/NAND4_in[0] ,
         \SB1_4_30/Component_Function_2/NAND4_in[0] ,
         \SB1_4_30/Component_Function_3/NAND4_in[3] ,
         \SB1_4_30/Component_Function_3/NAND4_in[1] ,
         \SB1_4_30/Component_Function_3/NAND4_in[0] ,
         \SB1_4_30/Component_Function_4/NAND4_in[3] ,
         \SB1_4_30/Component_Function_4/NAND4_in[1] ,
         \SB1_4_30/Component_Function_4/NAND4_in[0] ,
         \SB1_4_31/Component_Function_2/NAND4_in[2] ,
         \SB1_4_31/Component_Function_2/NAND4_in[1] ,
         \SB1_4_31/Component_Function_2/NAND4_in[0] ,
         \SB1_4_31/Component_Function_3/NAND4_in[3] ,
         \SB1_4_31/Component_Function_3/NAND4_in[2] ,
         \SB1_4_31/Component_Function_3/NAND4_in[1] ,
         \SB1_4_31/Component_Function_3/NAND4_in[0] ,
         \SB1_4_31/Component_Function_4/NAND4_in[1] ,
         \SB2_4_0/Component_Function_2/NAND4_in[2] ,
         \SB2_4_0/Component_Function_2/NAND4_in[1] ,
         \SB2_4_0/Component_Function_2/NAND4_in[0] ,
         \SB2_4_0/Component_Function_3/NAND4_in[3] ,
         \SB2_4_0/Component_Function_3/NAND4_in[0] ,
         \SB2_4_0/Component_Function_4/NAND4_in[3] ,
         \SB2_4_0/Component_Function_4/NAND4_in[1] ,
         \SB2_4_0/Component_Function_4/NAND4_in[0] ,
         \SB2_4_1/Component_Function_2/NAND4_in[3] ,
         \SB2_4_1/Component_Function_2/NAND4_in[2] ,
         \SB2_4_1/Component_Function_2/NAND4_in[0] ,
         \SB2_4_1/Component_Function_3/NAND4_in[3] ,
         \SB2_4_1/Component_Function_3/NAND4_in[1] ,
         \SB2_4_1/Component_Function_3/NAND4_in[0] ,
         \SB2_4_1/Component_Function_4/NAND4_in[1] ,
         \SB2_4_1/Component_Function_4/NAND4_in[0] ,
         \SB2_4_2/Component_Function_2/NAND4_in[3] ,
         \SB2_4_2/Component_Function_2/NAND4_in[1] ,
         \SB2_4_2/Component_Function_2/NAND4_in[0] ,
         \SB2_4_2/Component_Function_3/NAND4_in[3] ,
         \SB2_4_2/Component_Function_3/NAND4_in[2] ,
         \SB2_4_2/Component_Function_3/NAND4_in[1] ,
         \SB2_4_2/Component_Function_3/NAND4_in[0] ,
         \SB2_4_2/Component_Function_4/NAND4_in[3] ,
         \SB2_4_2/Component_Function_4/NAND4_in[1] ,
         \SB2_4_2/Component_Function_4/NAND4_in[0] ,
         \SB2_4_3/Component_Function_2/NAND4_in[3] ,
         \SB2_4_3/Component_Function_2/NAND4_in[2] ,
         \SB2_4_3/Component_Function_2/NAND4_in[0] ,
         \SB2_4_3/Component_Function_3/NAND4_in[3] ,
         \SB2_4_3/Component_Function_3/NAND4_in[1] ,
         \SB2_4_3/Component_Function_3/NAND4_in[0] ,
         \SB2_4_3/Component_Function_4/NAND4_in[3] ,
         \SB2_4_3/Component_Function_4/NAND4_in[2] ,
         \SB2_4_3/Component_Function_4/NAND4_in[1] ,
         \SB2_4_3/Component_Function_4/NAND4_in[0] ,
         \SB2_4_4/Component_Function_2/NAND4_in[2] ,
         \SB2_4_4/Component_Function_2/NAND4_in[1] ,
         \SB2_4_4/Component_Function_2/NAND4_in[0] ,
         \SB2_4_4/Component_Function_3/NAND4_in[2] ,
         \SB2_4_4/Component_Function_3/NAND4_in[0] ,
         \SB2_4_4/Component_Function_4/NAND4_in[3] ,
         \SB2_4_4/Component_Function_4/NAND4_in[1] ,
         \SB2_4_4/Component_Function_4/NAND4_in[0] ,
         \SB2_4_5/Component_Function_2/NAND4_in[3] ,
         \SB2_4_5/Component_Function_2/NAND4_in[2] ,
         \SB2_4_5/Component_Function_2/NAND4_in[1] ,
         \SB2_4_5/Component_Function_2/NAND4_in[0] ,
         \SB2_4_5/Component_Function_3/NAND4_in[2] ,
         \SB2_4_5/Component_Function_4/NAND4_in[2] ,
         \SB2_4_5/Component_Function_4/NAND4_in[1] ,
         \SB2_4_5/Component_Function_4/NAND4_in[0] ,
         \SB2_4_6/Component_Function_2/NAND4_in[3] ,
         \SB2_4_6/Component_Function_2/NAND4_in[2] ,
         \SB2_4_6/Component_Function_2/NAND4_in[1] ,
         \SB2_4_6/Component_Function_2/NAND4_in[0] ,
         \SB2_4_6/Component_Function_3/NAND4_in[3] ,
         \SB2_4_6/Component_Function_3/NAND4_in[2] ,
         \SB2_4_6/Component_Function_3/NAND4_in[0] ,
         \SB2_4_6/Component_Function_4/NAND4_in[2] ,
         \SB2_4_6/Component_Function_4/NAND4_in[1] ,
         \SB2_4_6/Component_Function_4/NAND4_in[0] ,
         \SB2_4_7/Component_Function_2/NAND4_in[0] ,
         \SB2_4_7/Component_Function_3/NAND4_in[2] ,
         \SB2_4_7/Component_Function_3/NAND4_in[0] ,
         \SB2_4_7/Component_Function_4/NAND4_in[3] ,
         \SB2_4_7/Component_Function_4/NAND4_in[1] ,
         \SB2_4_7/Component_Function_4/NAND4_in[0] ,
         \SB2_4_8/Component_Function_2/NAND4_in[2] ,
         \SB2_4_8/Component_Function_2/NAND4_in[1] ,
         \SB2_4_8/Component_Function_2/NAND4_in[0] ,
         \SB2_4_8/Component_Function_3/NAND4_in[3] ,
         \SB2_4_8/Component_Function_3/NAND4_in[2] ,
         \SB2_4_8/Component_Function_3/NAND4_in[0] ,
         \SB2_4_8/Component_Function_4/NAND4_in[3] ,
         \SB2_4_8/Component_Function_4/NAND4_in[0] ,
         \SB2_4_9/Component_Function_2/NAND4_in[2] ,
         \SB2_4_9/Component_Function_3/NAND4_in[0] ,
         \SB2_4_9/Component_Function_4/NAND4_in[2] ,
         \SB2_4_9/Component_Function_4/NAND4_in[1] ,
         \SB2_4_9/Component_Function_4/NAND4_in[0] ,
         \SB2_4_10/Component_Function_2/NAND4_in[3] ,
         \SB2_4_10/Component_Function_3/NAND4_in[2] ,
         \SB2_4_10/Component_Function_3/NAND4_in[1] ,
         \SB2_4_10/Component_Function_3/NAND4_in[0] ,
         \SB2_4_10/Component_Function_4/NAND4_in[3] ,
         \SB2_4_10/Component_Function_4/NAND4_in[2] ,
         \SB2_4_10/Component_Function_4/NAND4_in[1] ,
         \SB2_4_10/Component_Function_4/NAND4_in[0] ,
         \SB2_4_11/Component_Function_2/NAND4_in[2] ,
         \SB2_4_11/Component_Function_2/NAND4_in[1] ,
         \SB2_4_11/Component_Function_2/NAND4_in[0] ,
         \SB2_4_11/Component_Function_3/NAND4_in[3] ,
         \SB2_4_11/Component_Function_3/NAND4_in[0] ,
         \SB2_4_11/Component_Function_4/NAND4_in[3] ,
         \SB2_4_11/Component_Function_4/NAND4_in[2] ,
         \SB2_4_11/Component_Function_4/NAND4_in[1] ,
         \SB2_4_11/Component_Function_4/NAND4_in[0] ,
         \SB2_4_12/Component_Function_2/NAND4_in[2] ,
         \SB2_4_12/Component_Function_2/NAND4_in[0] ,
         \SB2_4_12/Component_Function_3/NAND4_in[2] ,
         \SB2_4_12/Component_Function_3/NAND4_in[1] ,
         \SB2_4_12/Component_Function_3/NAND4_in[0] ,
         \SB2_4_12/Component_Function_4/NAND4_in[3] ,
         \SB2_4_12/Component_Function_4/NAND4_in[2] ,
         \SB2_4_12/Component_Function_4/NAND4_in[1] ,
         \SB2_4_12/Component_Function_4/NAND4_in[0] ,
         \SB2_4_13/Component_Function_2/NAND4_in[2] ,
         \SB2_4_13/Component_Function_2/NAND4_in[0] ,
         \SB2_4_13/Component_Function_3/NAND4_in[3] ,
         \SB2_4_13/Component_Function_3/NAND4_in[1] ,
         \SB2_4_13/Component_Function_3/NAND4_in[0] ,
         \SB2_4_13/Component_Function_4/NAND4_in[1] ,
         \SB2_4_13/Component_Function_4/NAND4_in[0] ,
         \SB2_4_14/Component_Function_2/NAND4_in[3] ,
         \SB2_4_14/Component_Function_2/NAND4_in[2] ,
         \SB2_4_14/Component_Function_2/NAND4_in[0] ,
         \SB2_4_14/Component_Function_3/NAND4_in[3] ,
         \SB2_4_14/Component_Function_3/NAND4_in[2] ,
         \SB2_4_14/Component_Function_3/NAND4_in[1] ,
         \SB2_4_14/Component_Function_3/NAND4_in[0] ,
         \SB2_4_14/Component_Function_4/NAND4_in[1] ,
         \SB2_4_14/Component_Function_4/NAND4_in[0] ,
         \SB2_4_15/Component_Function_3/NAND4_in[3] ,
         \SB2_4_15/Component_Function_3/NAND4_in[2] ,
         \SB2_4_15/Component_Function_3/NAND4_in[0] ,
         \SB2_4_15/Component_Function_4/NAND4_in[3] ,
         \SB2_4_15/Component_Function_4/NAND4_in[1] ,
         \SB2_4_15/Component_Function_4/NAND4_in[0] ,
         \SB2_4_16/Component_Function_2/NAND4_in[2] ,
         \SB2_4_16/Component_Function_2/NAND4_in[0] ,
         \SB2_4_16/Component_Function_3/NAND4_in[3] ,
         \SB2_4_16/Component_Function_3/NAND4_in[0] ,
         \SB2_4_16/Component_Function_4/NAND4_in[3] ,
         \SB2_4_16/Component_Function_4/NAND4_in[0] ,
         \SB2_4_17/Component_Function_2/NAND4_in[3] ,
         \SB2_4_17/Component_Function_2/NAND4_in[2] ,
         \SB2_4_17/Component_Function_2/NAND4_in[1] ,
         \SB2_4_17/Component_Function_2/NAND4_in[0] ,
         \SB2_4_17/Component_Function_3/NAND4_in[3] ,
         \SB2_4_17/Component_Function_3/NAND4_in[0] ,
         \SB2_4_17/Component_Function_4/NAND4_in[3] ,
         \SB2_4_17/Component_Function_4/NAND4_in[1] ,
         \SB2_4_17/Component_Function_4/NAND4_in[0] ,
         \SB2_4_18/Component_Function_2/NAND4_in[2] ,
         \SB2_4_18/Component_Function_2/NAND4_in[0] ,
         \SB2_4_18/Component_Function_3/NAND4_in[3] ,
         \SB2_4_18/Component_Function_3/NAND4_in[1] ,
         \SB2_4_18/Component_Function_3/NAND4_in[0] ,
         \SB2_4_18/Component_Function_4/NAND4_in[3] ,
         \SB2_4_18/Component_Function_4/NAND4_in[1] ,
         \SB2_4_18/Component_Function_4/NAND4_in[0] ,
         \SB2_4_19/Component_Function_2/NAND4_in[3] ,
         \SB2_4_19/Component_Function_2/NAND4_in[1] ,
         \SB2_4_19/Component_Function_2/NAND4_in[0] ,
         \SB2_4_19/Component_Function_3/NAND4_in[3] ,
         \SB2_4_19/Component_Function_3/NAND4_in[1] ,
         \SB2_4_19/Component_Function_3/NAND4_in[0] ,
         \SB2_4_19/Component_Function_4/NAND4_in[2] ,
         \SB2_4_19/Component_Function_4/NAND4_in[1] ,
         \SB2_4_19/Component_Function_4/NAND4_in[0] ,
         \SB2_4_20/Component_Function_2/NAND4_in[3] ,
         \SB2_4_20/Component_Function_2/NAND4_in[2] ,
         \SB2_4_20/Component_Function_2/NAND4_in[1] ,
         \SB2_4_20/Component_Function_2/NAND4_in[0] ,
         \SB2_4_20/Component_Function_3/NAND4_in[2] ,
         \SB2_4_20/Component_Function_3/NAND4_in[0] ,
         \SB2_4_20/Component_Function_4/NAND4_in[3] ,
         \SB2_4_20/Component_Function_4/NAND4_in[1] ,
         \SB2_4_21/Component_Function_2/NAND4_in[2] ,
         \SB2_4_21/Component_Function_2/NAND4_in[0] ,
         \SB2_4_21/Component_Function_3/NAND4_in[3] ,
         \SB2_4_21/Component_Function_3/NAND4_in[2] ,
         \SB2_4_21/Component_Function_3/NAND4_in[1] ,
         \SB2_4_21/Component_Function_3/NAND4_in[0] ,
         \SB2_4_21/Component_Function_4/NAND4_in[3] ,
         \SB2_4_21/Component_Function_4/NAND4_in[1] ,
         \SB2_4_21/Component_Function_4/NAND4_in[0] ,
         \SB2_4_22/Component_Function_2/NAND4_in[0] ,
         \SB2_4_22/Component_Function_3/NAND4_in[3] ,
         \SB2_4_22/Component_Function_3/NAND4_in[1] ,
         \SB2_4_22/Component_Function_3/NAND4_in[0] ,
         \SB2_4_22/Component_Function_4/NAND4_in[3] ,
         \SB2_4_22/Component_Function_4/NAND4_in[1] ,
         \SB2_4_23/Component_Function_2/NAND4_in[3] ,
         \SB2_4_23/Component_Function_2/NAND4_in[2] ,
         \SB2_4_23/Component_Function_2/NAND4_in[1] ,
         \SB2_4_23/Component_Function_2/NAND4_in[0] ,
         \SB2_4_23/Component_Function_3/NAND4_in[3] ,
         \SB2_4_23/Component_Function_3/NAND4_in[2] ,
         \SB2_4_23/Component_Function_3/NAND4_in[1] ,
         \SB2_4_23/Component_Function_3/NAND4_in[0] ,
         \SB2_4_23/Component_Function_4/NAND4_in[3] ,
         \SB2_4_24/Component_Function_2/NAND4_in[3] ,
         \SB2_4_24/Component_Function_2/NAND4_in[1] ,
         \SB2_4_24/Component_Function_3/NAND4_in[3] ,
         \SB2_4_24/Component_Function_3/NAND4_in[1] ,
         \SB2_4_24/Component_Function_3/NAND4_in[0] ,
         \SB2_4_24/Component_Function_4/NAND4_in[3] ,
         \SB2_4_24/Component_Function_4/NAND4_in[1] ,
         \SB2_4_24/Component_Function_4/NAND4_in[0] ,
         \SB2_4_25/Component_Function_2/NAND4_in[0] ,
         \SB2_4_25/Component_Function_3/NAND4_in[2] ,
         \SB2_4_25/Component_Function_3/NAND4_in[1] ,
         \SB2_4_25/Component_Function_3/NAND4_in[0] ,
         \SB2_4_25/Component_Function_4/NAND4_in[1] ,
         \SB2_4_25/Component_Function_4/NAND4_in[0] ,
         \SB2_4_26/Component_Function_2/NAND4_in[1] ,
         \SB2_4_26/Component_Function_2/NAND4_in[0] ,
         \SB2_4_26/Component_Function_3/NAND4_in[3] ,
         \SB2_4_26/Component_Function_3/NAND4_in[1] ,
         \SB2_4_26/Component_Function_3/NAND4_in[0] ,
         \SB2_4_26/Component_Function_4/NAND4_in[3] ,
         \SB2_4_26/Component_Function_4/NAND4_in[2] ,
         \SB2_4_26/Component_Function_4/NAND4_in[1] ,
         \SB2_4_26/Component_Function_4/NAND4_in[0] ,
         \SB2_4_27/Component_Function_2/NAND4_in[3] ,
         \SB2_4_27/Component_Function_2/NAND4_in[2] ,
         \SB2_4_27/Component_Function_2/NAND4_in[1] ,
         \SB2_4_27/Component_Function_3/NAND4_in[2] ,
         \SB2_4_27/Component_Function_3/NAND4_in[0] ,
         \SB2_4_27/Component_Function_4/NAND4_in[3] ,
         \SB2_4_27/Component_Function_4/NAND4_in[1] ,
         \SB2_4_27/Component_Function_4/NAND4_in[0] ,
         \SB2_4_28/Component_Function_2/NAND4_in[2] ,
         \SB2_4_28/Component_Function_2/NAND4_in[1] ,
         \SB2_4_28/Component_Function_2/NAND4_in[0] ,
         \SB2_4_28/Component_Function_3/NAND4_in[3] ,
         \SB2_4_28/Component_Function_3/NAND4_in[2] ,
         \SB2_4_28/Component_Function_3/NAND4_in[1] ,
         \SB2_4_28/Component_Function_3/NAND4_in[0] ,
         \SB2_4_28/Component_Function_4/NAND4_in[3] ,
         \SB2_4_28/Component_Function_4/NAND4_in[2] ,
         \SB2_4_28/Component_Function_4/NAND4_in[1] ,
         \SB2_4_29/Component_Function_2/NAND4_in[2] ,
         \SB2_4_29/Component_Function_2/NAND4_in[1] ,
         \SB2_4_29/Component_Function_2/NAND4_in[0] ,
         \SB2_4_29/Component_Function_3/NAND4_in[1] ,
         \SB2_4_29/Component_Function_3/NAND4_in[0] ,
         \SB2_4_29/Component_Function_4/NAND4_in[3] ,
         \SB2_4_29/Component_Function_4/NAND4_in[0] ,
         \SB2_4_30/Component_Function_2/NAND4_in[2] ,
         \SB2_4_30/Component_Function_2/NAND4_in[0] ,
         \SB2_4_30/Component_Function_3/NAND4_in[3] ,
         \SB2_4_30/Component_Function_3/NAND4_in[0] ,
         \SB2_4_30/Component_Function_4/NAND4_in[3] ,
         \SB2_4_30/Component_Function_4/NAND4_in[2] ,
         \SB2_4_30/Component_Function_4/NAND4_in[1] ,
         \SB2_4_30/Component_Function_4/NAND4_in[0] ,
         \SB2_4_31/Component_Function_2/NAND4_in[3] ,
         \SB2_4_31/Component_Function_2/NAND4_in[2] ,
         \SB2_4_31/Component_Function_2/NAND4_in[1] ,
         \SB2_4_31/Component_Function_2/NAND4_in[0] ,
         \SB2_4_31/Component_Function_3/NAND4_in[3] ,
         \SB2_4_31/Component_Function_3/NAND4_in[2] ,
         \SB2_4_31/Component_Function_3/NAND4_in[1] ,
         \SB2_4_31/Component_Function_3/NAND4_in[0] ,
         \SB2_4_31/Component_Function_4/NAND4_in[1] ,
         \SB2_4_31/Component_Function_4/NAND4_in[0] ,
         \SB3_0/Component_Function_2/NAND4_in[1] ,
         \SB3_0/Component_Function_2/NAND4_in[0] ,
         \SB3_0/Component_Function_3/NAND4_in[1] ,
         \SB3_0/Component_Function_4/NAND4_in[3] ,
         \SB3_0/Component_Function_4/NAND4_in[2] ,
         \SB3_0/Component_Function_4/NAND4_in[1] ,
         \SB3_0/Component_Function_4/NAND4_in[0] ,
         \SB3_1/Component_Function_2/NAND4_in[2] ,
         \SB3_1/Component_Function_2/NAND4_in[1] ,
         \SB3_1/Component_Function_2/NAND4_in[0] ,
         \SB3_1/Component_Function_3/NAND4_in[2] ,
         \SB3_1/Component_Function_3/NAND4_in[1] ,
         \SB3_1/Component_Function_3/NAND4_in[0] ,
         \SB3_1/Component_Function_4/NAND4_in[3] ,
         \SB3_1/Component_Function_4/NAND4_in[2] ,
         \SB3_2/Component_Function_2/NAND4_in[3] ,
         \SB3_2/Component_Function_2/NAND4_in[1] ,
         \SB3_2/Component_Function_3/NAND4_in[0] ,
         \SB3_2/Component_Function_4/NAND4_in[3] ,
         \SB3_2/Component_Function_4/NAND4_in[2] ,
         \SB3_2/Component_Function_4/NAND4_in[1] ,
         \SB3_2/Component_Function_4/NAND4_in[0] ,
         \SB3_3/Component_Function_2/NAND4_in[3] ,
         \SB3_3/Component_Function_2/NAND4_in[2] ,
         \SB3_3/Component_Function_3/NAND4_in[3] ,
         \SB3_3/Component_Function_3/NAND4_in[1] ,
         \SB3_3/Component_Function_3/NAND4_in[0] ,
         \SB3_3/Component_Function_4/NAND4_in[2] ,
         \SB3_3/Component_Function_4/NAND4_in[1] ,
         \SB3_3/Component_Function_4/NAND4_in[0] ,
         \SB3_4/Component_Function_2/NAND4_in[3] ,
         \SB3_4/Component_Function_2/NAND4_in[2] ,
         \SB3_4/Component_Function_2/NAND4_in[0] ,
         \SB3_4/Component_Function_3/NAND4_in[3] ,
         \SB3_4/Component_Function_3/NAND4_in[1] ,
         \SB3_4/Component_Function_3/NAND4_in[0] ,
         \SB3_4/Component_Function_4/NAND4_in[3] ,
         \SB3_4/Component_Function_4/NAND4_in[2] ,
         \SB3_4/Component_Function_4/NAND4_in[1] ,
         \SB3_4/Component_Function_4/NAND4_in[0] ,
         \SB3_5/Component_Function_2/NAND4_in[2] ,
         \SB3_5/Component_Function_2/NAND4_in[1] ,
         \SB3_5/Component_Function_2/NAND4_in[0] ,
         \SB3_5/Component_Function_3/NAND4_in[2] ,
         \SB3_5/Component_Function_3/NAND4_in[1] ,
         \SB3_5/Component_Function_3/NAND4_in[0] ,
         \SB3_5/Component_Function_4/NAND4_in[3] ,
         \SB3_5/Component_Function_4/NAND4_in[2] ,
         \SB3_5/Component_Function_4/NAND4_in[1] ,
         \SB3_5/Component_Function_4/NAND4_in[0] ,
         \SB3_6/Component_Function_2/NAND4_in[2] ,
         \SB3_6/Component_Function_2/NAND4_in[1] ,
         \SB3_6/Component_Function_2/NAND4_in[0] ,
         \SB3_6/Component_Function_3/NAND4_in[3] ,
         \SB3_6/Component_Function_3/NAND4_in[1] ,
         \SB3_6/Component_Function_4/NAND4_in[2] ,
         \SB3_6/Component_Function_4/NAND4_in[1] ,
         \SB3_6/Component_Function_4/NAND4_in[0] ,
         \SB3_7/Component_Function_2/NAND4_in[3] ,
         \SB3_7/Component_Function_2/NAND4_in[2] ,
         \SB3_7/Component_Function_2/NAND4_in[1] ,
         \SB3_7/Component_Function_3/NAND4_in[3] ,
         \SB3_7/Component_Function_3/NAND4_in[1] ,
         \SB3_7/Component_Function_4/NAND4_in[2] ,
         \SB3_7/Component_Function_4/NAND4_in[0] ,
         \SB3_8/Component_Function_2/NAND4_in[2] ,
         \SB3_8/Component_Function_2/NAND4_in[1] ,
         \SB3_8/Component_Function_2/NAND4_in[0] ,
         \SB3_8/Component_Function_3/NAND4_in[3] ,
         \SB3_8/Component_Function_3/NAND4_in[2] ,
         \SB3_8/Component_Function_3/NAND4_in[1] ,
         \SB3_8/Component_Function_3/NAND4_in[0] ,
         \SB3_8/Component_Function_4/NAND4_in[3] ,
         \SB3_8/Component_Function_4/NAND4_in[2] ,
         \SB3_8/Component_Function_4/NAND4_in[1] ,
         \SB3_8/Component_Function_4/NAND4_in[0] ,
         \SB3_9/Component_Function_2/NAND4_in[2] ,
         \SB3_9/Component_Function_3/NAND4_in[3] ,
         \SB3_9/Component_Function_3/NAND4_in[2] ,
         \SB3_9/Component_Function_3/NAND4_in[1] ,
         \SB3_9/Component_Function_3/NAND4_in[0] ,
         \SB3_9/Component_Function_4/NAND4_in[3] ,
         \SB3_9/Component_Function_4/NAND4_in[2] ,
         \SB3_9/Component_Function_4/NAND4_in[1] ,
         \SB3_9/Component_Function_4/NAND4_in[0] ,
         \SB3_10/Component_Function_2/NAND4_in[2] ,
         \SB3_10/Component_Function_2/NAND4_in[1] ,
         \SB3_10/Component_Function_2/NAND4_in[0] ,
         \SB3_10/Component_Function_3/NAND4_in[3] ,
         \SB3_10/Component_Function_3/NAND4_in[2] ,
         \SB3_10/Component_Function_3/NAND4_in[0] ,
         \SB3_10/Component_Function_4/NAND4_in[3] ,
         \SB3_10/Component_Function_4/NAND4_in[1] ,
         \SB3_10/Component_Function_4/NAND4_in[0] ,
         \SB3_11/Component_Function_2/NAND4_in[2] ,
         \SB3_11/Component_Function_2/NAND4_in[1] ,
         \SB3_11/Component_Function_2/NAND4_in[0] ,
         \SB3_11/Component_Function_3/NAND4_in[3] ,
         \SB3_11/Component_Function_3/NAND4_in[2] ,
         \SB3_11/Component_Function_3/NAND4_in[1] ,
         \SB3_11/Component_Function_3/NAND4_in[0] ,
         \SB3_11/Component_Function_4/NAND4_in[2] ,
         \SB3_11/Component_Function_4/NAND4_in[0] ,
         \SB3_12/Component_Function_2/NAND4_in[0] ,
         \SB3_12/Component_Function_3/NAND4_in[3] ,
         \SB3_12/Component_Function_3/NAND4_in[0] ,
         \SB3_12/Component_Function_4/NAND4_in[1] ,
         \SB3_12/Component_Function_4/NAND4_in[0] ,
         \SB3_13/Component_Function_2/NAND4_in[1] ,
         \SB3_13/Component_Function_2/NAND4_in[0] ,
         \SB3_13/Component_Function_3/NAND4_in[0] ,
         \SB3_13/Component_Function_4/NAND4_in[1] ,
         \SB3_13/Component_Function_4/NAND4_in[0] ,
         \SB3_14/Component_Function_2/NAND4_in[3] ,
         \SB3_14/Component_Function_2/NAND4_in[0] ,
         \SB3_14/Component_Function_3/NAND4_in[2] ,
         \SB3_14/Component_Function_3/NAND4_in[1] ,
         \SB3_14/Component_Function_4/NAND4_in[3] ,
         \SB3_14/Component_Function_4/NAND4_in[2] ,
         \SB3_14/Component_Function_4/NAND4_in[0] ,
         \SB3_15/Component_Function_2/NAND4_in[1] ,
         \SB3_15/Component_Function_2/NAND4_in[0] ,
         \SB3_15/Component_Function_3/NAND4_in[3] ,
         \SB3_15/Component_Function_3/NAND4_in[1] ,
         \SB3_15/Component_Function_3/NAND4_in[0] ,
         \SB3_15/Component_Function_4/NAND4_in[3] ,
         \SB3_15/Component_Function_4/NAND4_in[2] ,
         \SB3_15/Component_Function_4/NAND4_in[0] ,
         \SB3_16/Component_Function_2/NAND4_in[2] ,
         \SB3_16/Component_Function_2/NAND4_in[1] ,
         \SB3_16/Component_Function_2/NAND4_in[0] ,
         \SB3_16/Component_Function_3/NAND4_in[1] ,
         \SB3_16/Component_Function_3/NAND4_in[0] ,
         \SB3_16/Component_Function_4/NAND4_in[3] ,
         \SB3_16/Component_Function_4/NAND4_in[1] ,
         \SB3_16/Component_Function_4/NAND4_in[0] ,
         \SB3_17/Component_Function_2/NAND4_in[2] ,
         \SB3_17/Component_Function_2/NAND4_in[1] ,
         \SB3_17/Component_Function_3/NAND4_in[2] ,
         \SB3_17/Component_Function_3/NAND4_in[1] ,
         \SB3_17/Component_Function_3/NAND4_in[0] ,
         \SB3_17/Component_Function_4/NAND4_in[3] ,
         \SB3_17/Component_Function_4/NAND4_in[1] ,
         \SB3_17/Component_Function_4/NAND4_in[0] ,
         \SB3_18/Component_Function_2/NAND4_in[3] ,
         \SB3_18/Component_Function_2/NAND4_in[2] ,
         \SB3_18/Component_Function_2/NAND4_in[0] ,
         \SB3_18/Component_Function_3/NAND4_in[1] ,
         \SB3_18/Component_Function_4/NAND4_in[3] ,
         \SB3_18/Component_Function_4/NAND4_in[2] ,
         \SB3_18/Component_Function_4/NAND4_in[1] ,
         \SB3_18/Component_Function_4/NAND4_in[0] ,
         \SB3_19/Component_Function_2/NAND4_in[3] ,
         \SB3_19/Component_Function_2/NAND4_in[1] ,
         \SB3_19/Component_Function_3/NAND4_in[3] ,
         \SB3_19/Component_Function_3/NAND4_in[2] ,
         \SB3_19/Component_Function_3/NAND4_in[1] ,
         \SB3_19/Component_Function_3/NAND4_in[0] ,
         \SB3_19/Component_Function_4/NAND4_in[3] ,
         \SB3_19/Component_Function_4/NAND4_in[2] ,
         \SB3_19/Component_Function_4/NAND4_in[1] ,
         \SB3_19/Component_Function_4/NAND4_in[0] ,
         \SB3_20/Component_Function_2/NAND4_in[1] ,
         \SB3_20/Component_Function_2/NAND4_in[0] ,
         \SB3_20/Component_Function_3/NAND4_in[2] ,
         \SB3_20/Component_Function_3/NAND4_in[0] ,
         \SB3_20/Component_Function_4/NAND4_in[3] ,
         \SB3_20/Component_Function_4/NAND4_in[1] ,
         \SB3_20/Component_Function_4/NAND4_in[0] ,
         \SB3_21/Component_Function_2/NAND4_in[3] ,
         \SB3_21/Component_Function_2/NAND4_in[2] ,
         \SB3_21/Component_Function_2/NAND4_in[1] ,
         \SB3_21/Component_Function_2/NAND4_in[0] ,
         \SB3_21/Component_Function_3/NAND4_in[1] ,
         \SB3_21/Component_Function_3/NAND4_in[0] ,
         \SB3_21/Component_Function_4/NAND4_in[2] ,
         \SB3_21/Component_Function_4/NAND4_in[1] ,
         \SB3_21/Component_Function_4/NAND4_in[0] ,
         \SB3_22/Component_Function_2/NAND4_in[2] ,
         \SB3_22/Component_Function_2/NAND4_in[1] ,
         \SB3_22/Component_Function_2/NAND4_in[0] ,
         \SB3_22/Component_Function_3/NAND4_in[2] ,
         \SB3_22/Component_Function_3/NAND4_in[1] ,
         \SB3_22/Component_Function_3/NAND4_in[0] ,
         \SB3_22/Component_Function_4/NAND4_in[3] ,
         \SB3_22/Component_Function_4/NAND4_in[2] ,
         \SB3_22/Component_Function_4/NAND4_in[1] ,
         \SB3_22/Component_Function_4/NAND4_in[0] ,
         \SB3_23/Component_Function_2/NAND4_in[3] ,
         \SB3_23/Component_Function_2/NAND4_in[1] ,
         \SB3_23/Component_Function_3/NAND4_in[2] ,
         \SB3_23/Component_Function_3/NAND4_in[1] ,
         \SB3_23/Component_Function_4/NAND4_in[3] ,
         \SB3_23/Component_Function_4/NAND4_in[1] ,
         \SB3_24/Component_Function_2/NAND4_in[3] ,
         \SB3_24/Component_Function_2/NAND4_in[2] ,
         \SB3_24/Component_Function_2/NAND4_in[1] ,
         \SB3_24/Component_Function_2/NAND4_in[0] ,
         \SB3_24/Component_Function_3/NAND4_in[1] ,
         \SB3_24/Component_Function_4/NAND4_in[3] ,
         \SB3_24/Component_Function_4/NAND4_in[1] ,
         \SB3_24/Component_Function_4/NAND4_in[0] ,
         \SB3_25/Component_Function_2/NAND4_in[3] ,
         \SB3_25/Component_Function_2/NAND4_in[2] ,
         \SB3_25/Component_Function_2/NAND4_in[0] ,
         \SB3_25/Component_Function_3/NAND4_in[2] ,
         \SB3_25/Component_Function_3/NAND4_in[1] ,
         \SB3_25/Component_Function_3/NAND4_in[0] ,
         \SB3_25/Component_Function_4/NAND4_in[1] ,
         \SB3_25/Component_Function_4/NAND4_in[0] ,
         \SB3_26/Component_Function_2/NAND4_in[1] ,
         \SB3_26/Component_Function_2/NAND4_in[0] ,
         \SB3_26/Component_Function_3/NAND4_in[3] ,
         \SB3_26/Component_Function_3/NAND4_in[2] ,
         \SB3_26/Component_Function_3/NAND4_in[1] ,
         \SB3_26/Component_Function_3/NAND4_in[0] ,
         \SB3_26/Component_Function_4/NAND4_in[3] ,
         \SB3_26/Component_Function_4/NAND4_in[2] ,
         \SB3_26/Component_Function_4/NAND4_in[1] ,
         \SB3_26/Component_Function_4/NAND4_in[0] ,
         \SB3_27/Component_Function_2/NAND4_in[1] ,
         \SB3_27/Component_Function_2/NAND4_in[0] ,
         \SB3_27/Component_Function_3/NAND4_in[3] ,
         \SB3_27/Component_Function_3/NAND4_in[2] ,
         \SB3_27/Component_Function_3/NAND4_in[0] ,
         \SB3_27/Component_Function_4/NAND4_in[1] ,
         \SB3_27/Component_Function_4/NAND4_in[0] ,
         \SB3_28/Component_Function_2/NAND4_in[3] ,
         \SB3_28/Component_Function_2/NAND4_in[2] ,
         \SB3_28/Component_Function_2/NAND4_in[1] ,
         \SB3_28/Component_Function_2/NAND4_in[0] ,
         \SB3_28/Component_Function_3/NAND4_in[2] ,
         \SB3_28/Component_Function_3/NAND4_in[1] ,
         \SB3_28/Component_Function_3/NAND4_in[0] ,
         \SB3_28/Component_Function_4/NAND4_in[3] ,
         \SB3_28/Component_Function_4/NAND4_in[1] ,
         \SB3_28/Component_Function_4/NAND4_in[0] ,
         \SB3_29/Component_Function_2/NAND4_in[3] ,
         \SB3_29/Component_Function_2/NAND4_in[2] ,
         \SB3_29/Component_Function_2/NAND4_in[1] ,
         \SB3_29/Component_Function_2/NAND4_in[0] ,
         \SB3_29/Component_Function_3/NAND4_in[2] ,
         \SB3_29/Component_Function_3/NAND4_in[1] ,
         \SB3_29/Component_Function_3/NAND4_in[0] ,
         \SB3_29/Component_Function_4/NAND4_in[2] ,
         \SB3_29/Component_Function_4/NAND4_in[1] ,
         \SB3_29/Component_Function_4/NAND4_in[0] ,
         \SB3_30/Component_Function_2/NAND4_in[3] ,
         \SB3_30/Component_Function_2/NAND4_in[2] ,
         \SB3_30/Component_Function_2/NAND4_in[1] ,
         \SB3_30/Component_Function_2/NAND4_in[0] ,
         \SB3_30/Component_Function_3/NAND4_in[1] ,
         \SB3_30/Component_Function_3/NAND4_in[0] ,
         \SB3_30/Component_Function_4/NAND4_in[3] ,
         \SB3_30/Component_Function_4/NAND4_in[1] ,
         \SB3_30/Component_Function_4/NAND4_in[0] ,
         \SB3_31/Component_Function_2/NAND4_in[2] ,
         \SB3_31/Component_Function_2/NAND4_in[1] ,
         \SB3_31/Component_Function_3/NAND4_in[1] ,
         \SB3_31/Component_Function_3/NAND4_in[0] ,
         \SB3_31/Component_Function_4/NAND4_in[3] ,
         \SB3_31/Component_Function_4/NAND4_in[1] ,
         \SB3_31/Component_Function_4/NAND4_in[0] ,
         \SB4_0/Component_Function_2/NAND4_in[2] ,
         \SB4_0/Component_Function_2/NAND4_in[1] ,
         \SB4_0/Component_Function_2/NAND4_in[0] ,
         \SB4_0/Component_Function_3/NAND4_in[3] ,
         \SB4_0/Component_Function_4/NAND4_in[2] ,
         \SB4_0/Component_Function_4/NAND4_in[0] ,
         \SB4_1/Component_Function_2/NAND4_in[0] ,
         \SB4_1/Component_Function_3/NAND4_in[3] ,
         \SB4_1/Component_Function_3/NAND4_in[0] ,
         \SB4_1/Component_Function_4/NAND4_in[3] ,
         \SB4_1/Component_Function_4/NAND4_in[0] ,
         \SB4_2/Component_Function_2/NAND4_in[3] ,
         \SB4_2/Component_Function_2/NAND4_in[1] ,
         \SB4_2/Component_Function_2/NAND4_in[0] ,
         \SB4_2/Component_Function_3/NAND4_in[3] ,
         \SB4_2/Component_Function_3/NAND4_in[2] ,
         \SB4_2/Component_Function_4/NAND4_in[3] ,
         \SB4_2/Component_Function_4/NAND4_in[0] ,
         \SB4_3/Component_Function_2/NAND4_in[2] ,
         \SB4_3/Component_Function_3/NAND4_in[3] ,
         \SB4_3/Component_Function_3/NAND4_in[1] ,
         \SB4_3/Component_Function_4/NAND4_in[0] ,
         \SB4_4/Component_Function_2/NAND4_in[2] ,
         \SB4_4/Component_Function_3/NAND4_in[3] ,
         \SB4_4/Component_Function_3/NAND4_in[1] ,
         \SB4_4/Component_Function_4/NAND4_in[3] ,
         \SB4_4/Component_Function_4/NAND4_in[2] ,
         \SB4_4/Component_Function_4/NAND4_in[1] ,
         \SB4_5/Component_Function_2/NAND4_in[2] ,
         \SB4_5/Component_Function_3/NAND4_in[3] ,
         \SB4_5/Component_Function_3/NAND4_in[1] ,
         \SB4_5/Component_Function_4/NAND4_in[1] ,
         \SB4_5/Component_Function_4/NAND4_in[0] ,
         \SB4_6/Component_Function_2/NAND4_in[3] ,
         \SB4_6/Component_Function_2/NAND4_in[2] ,
         \SB4_6/Component_Function_2/NAND4_in[0] ,
         \SB4_6/Component_Function_3/NAND4_in[3] ,
         \SB4_6/Component_Function_3/NAND4_in[2] ,
         \SB4_6/Component_Function_3/NAND4_in[1] ,
         \SB4_6/Component_Function_4/NAND4_in[3] ,
         \SB4_6/Component_Function_4/NAND4_in[2] ,
         \SB4_6/Component_Function_4/NAND4_in[0] ,
         \SB4_7/Component_Function_2/NAND4_in[2] ,
         \SB4_7/Component_Function_3/NAND4_in[3] ,
         \SB4_7/Component_Function_3/NAND4_in[0] ,
         \SB4_7/Component_Function_4/NAND4_in[1] ,
         \SB4_8/Component_Function_2/NAND4_in[2] ,
         \SB4_8/Component_Function_3/NAND4_in[3] ,
         \SB4_8/Component_Function_3/NAND4_in[1] ,
         \SB4_8/Component_Function_3/NAND4_in[0] ,
         \SB4_8/Component_Function_4/NAND4_in[2] ,
         \SB4_8/Component_Function_4/NAND4_in[1] ,
         \SB4_8/Component_Function_4/NAND4_in[0] ,
         \SB4_9/Component_Function_2/NAND4_in[0] ,
         \SB4_9/Component_Function_4/NAND4_in[3] ,
         \SB4_10/Component_Function_3/NAND4_in[3] ,
         \SB4_10/Component_Function_3/NAND4_in[1] ,
         \SB4_11/Component_Function_2/NAND4_in[2] ,
         \SB4_11/Component_Function_3/NAND4_in[1] ,
         \SB4_11/Component_Function_4/NAND4_in[0] ,
         \SB4_12/Component_Function_2/NAND4_in[2] ,
         \SB4_12/Component_Function_2/NAND4_in[0] ,
         \SB4_12/Component_Function_3/NAND4_in[1] ,
         \SB4_12/Component_Function_3/NAND4_in[0] ,
         \SB4_12/Component_Function_4/NAND4_in[3] ,
         \SB4_12/Component_Function_4/NAND4_in[1] ,
         \SB4_13/Component_Function_2/NAND4_in[2] ,
         \SB4_13/Component_Function_2/NAND4_in[1] ,
         \SB4_13/Component_Function_2/NAND4_in[0] ,
         \SB4_13/Component_Function_3/NAND4_in[3] ,
         \SB4_13/Component_Function_3/NAND4_in[2] ,
         \SB4_13/Component_Function_4/NAND4_in[3] ,
         \SB4_13/Component_Function_4/NAND4_in[2] ,
         \SB4_14/Component_Function_2/NAND4_in[2] ,
         \SB4_14/Component_Function_2/NAND4_in[0] ,
         \SB4_14/Component_Function_3/NAND4_in[3] ,
         \SB4_14/Component_Function_3/NAND4_in[2] ,
         \SB4_14/Component_Function_3/NAND4_in[1] ,
         \SB4_14/Component_Function_3/NAND4_in[0] ,
         \SB4_14/Component_Function_4/NAND4_in[2] ,
         \SB4_15/Component_Function_2/NAND4_in[2] ,
         \SB4_15/Component_Function_2/NAND4_in[1] ,
         \SB4_15/Component_Function_2/NAND4_in[0] ,
         \SB4_15/Component_Function_3/NAND4_in[3] ,
         \SB4_15/Component_Function_3/NAND4_in[1] ,
         \SB4_15/Component_Function_4/NAND4_in[3] ,
         \SB4_15/Component_Function_4/NAND4_in[0] ,
         \SB4_16/Component_Function_2/NAND4_in[2] ,
         \SB4_16/Component_Function_3/NAND4_in[3] ,
         \SB4_16/Component_Function_3/NAND4_in[0] ,
         \SB4_16/Component_Function_4/NAND4_in[1] ,
         \SB4_16/Component_Function_4/NAND4_in[0] ,
         \SB4_17/Component_Function_2/NAND4_in[3] ,
         \SB4_17/Component_Function_2/NAND4_in[1] ,
         \SB4_17/Component_Function_3/NAND4_in[2] ,
         \SB4_17/Component_Function_3/NAND4_in[1] ,
         \SB4_17/Component_Function_3/NAND4_in[0] ,
         \SB4_17/Component_Function_4/NAND4_in[0] ,
         \SB4_18/Component_Function_2/NAND4_in[3] ,
         \SB4_18/Component_Function_2/NAND4_in[2] ,
         \SB4_18/Component_Function_2/NAND4_in[0] ,
         \SB4_18/Component_Function_3/NAND4_in[2] ,
         \SB4_18/Component_Function_3/NAND4_in[1] ,
         \SB4_18/Component_Function_3/NAND4_in[0] ,
         \SB4_18/Component_Function_4/NAND4_in[3] ,
         \SB4_18/Component_Function_4/NAND4_in[1] ,
         \SB4_19/Component_Function_2/NAND4_in[3] ,
         \SB4_19/Component_Function_2/NAND4_in[2] ,
         \SB4_19/Component_Function_3/NAND4_in[3] ,
         \SB4_19/Component_Function_3/NAND4_in[1] ,
         \SB4_19/Component_Function_3/NAND4_in[0] ,
         \SB4_19/Component_Function_4/NAND4_in[3] ,
         \SB4_19/Component_Function_4/NAND4_in[1] ,
         \SB4_20/Component_Function_2/NAND4_in[0] ,
         \SB4_20/Component_Function_3/NAND4_in[3] ,
         \SB4_20/Component_Function_3/NAND4_in[2] ,
         \SB4_20/Component_Function_3/NAND4_in[0] ,
         \SB4_20/Component_Function_4/NAND4_in[2] ,
         \SB4_21/Component_Function_2/NAND4_in[3] ,
         \SB4_21/Component_Function_2/NAND4_in[2] ,
         \SB4_21/Component_Function_2/NAND4_in[1] ,
         \SB4_21/Component_Function_2/NAND4_in[0] ,
         \SB4_21/Component_Function_3/NAND4_in[2] ,
         \SB4_21/Component_Function_3/NAND4_in[1] ,
         \SB4_21/Component_Function_4/NAND4_in[3] ,
         \SB4_21/Component_Function_4/NAND4_in[0] ,
         \SB4_22/Component_Function_2/NAND4_in[2] ,
         \SB4_22/Component_Function_3/NAND4_in[3] ,
         \SB4_22/Component_Function_4/NAND4_in[3] ,
         \SB4_22/Component_Function_4/NAND4_in[2] ,
         \SB4_22/Component_Function_4/NAND4_in[0] ,
         \SB4_23/Component_Function_2/NAND4_in[2] ,
         \SB4_23/Component_Function_2/NAND4_in[0] ,
         \SB4_23/Component_Function_3/NAND4_in[3] ,
         \SB4_23/Component_Function_3/NAND4_in[1] ,
         \SB4_23/Component_Function_4/NAND4_in[3] ,
         \SB4_24/Component_Function_3/NAND4_in[3] ,
         \SB4_24/Component_Function_3/NAND4_in[1] ,
         \SB4_24/Component_Function_4/NAND4_in[0] ,
         \SB4_25/Component_Function_2/NAND4_in[3] ,
         \SB4_25/Component_Function_3/NAND4_in[3] ,
         \SB4_25/Component_Function_3/NAND4_in[1] ,
         \SB4_25/Component_Function_4/NAND4_in[3] ,
         \SB4_25/Component_Function_4/NAND4_in[1] ,
         \SB4_25/Component_Function_4/NAND4_in[0] ,
         \SB4_26/Component_Function_2/NAND4_in[0] ,
         \SB4_26/Component_Function_3/NAND4_in[3] ,
         \SB4_26/Component_Function_4/NAND4_in[1] ,
         \SB4_26/Component_Function_4/NAND4_in[0] ,
         \SB4_27/Component_Function_2/NAND4_in[0] ,
         \SB4_27/Component_Function_3/NAND4_in[3] ,
         \SB4_27/Component_Function_3/NAND4_in[2] ,
         \SB4_27/Component_Function_3/NAND4_in[1] ,
         \SB4_27/Component_Function_4/NAND4_in[1] ,
         \SB4_28/Component_Function_2/NAND4_in[2] ,
         \SB4_28/Component_Function_3/NAND4_in[2] ,
         \SB4_28/Component_Function_4/NAND4_in[2] ,
         \SB4_28/Component_Function_4/NAND4_in[0] ,
         \SB4_29/Component_Function_2/NAND4_in[2] ,
         \SB4_29/Component_Function_2/NAND4_in[0] ,
         \SB4_29/Component_Function_4/NAND4_in[0] ,
         \SB4_30/Component_Function_2/NAND4_in[0] ,
         \SB4_30/Component_Function_3/NAND4_in[3] ,
         \SB4_30/Component_Function_3/NAND4_in[2] ,
         \SB4_30/Component_Function_4/NAND4_in[3] ,
         \SB4_30/Component_Function_4/NAND4_in[1] ,
         \SB4_31/Component_Function_2/NAND4_in[0] ,
         \SB4_31/Component_Function_3/NAND4_in[2] ,
         \SB4_31/Component_Function_4/NAND4_in[3] ,
         \SB1_0_0/Component_Function_0/NAND4_in[3] ,
         \SB1_0_0/Component_Function_0/NAND4_in[1] ,
         \SB1_0_0/Component_Function_0/NAND4_in[0] ,
         \SB1_0_0/Component_Function_1/NAND4_in[3] ,
         \SB1_0_0/Component_Function_1/NAND4_in[2] ,
         \SB1_0_0/Component_Function_1/NAND4_in[1] ,
         \SB1_0_0/Component_Function_5/NAND4_in[2] ,
         \SB1_0_0/Component_Function_5/NAND4_in[1] ,
         \SB1_0_0/Component_Function_5/NAND4_in[0] ,
         \SB1_0_1/Component_Function_0/NAND4_in[3] ,
         \SB1_0_1/Component_Function_0/NAND4_in[2] ,
         \SB1_0_1/Component_Function_0/NAND4_in[1] ,
         \SB1_0_1/Component_Function_0/NAND4_in[0] ,
         \SB1_0_1/Component_Function_1/NAND4_in[3] ,
         \SB1_0_1/Component_Function_1/NAND4_in[2] ,
         \SB1_0_1/Component_Function_1/NAND4_in[1] ,
         \SB1_0_1/Component_Function_1/NAND4_in[0] ,
         \SB1_0_1/Component_Function_5/NAND4_in[3] ,
         \SB1_0_1/Component_Function_5/NAND4_in[1] ,
         \SB1_0_1/Component_Function_5/NAND4_in[0] ,
         \SB1_0_2/Component_Function_0/NAND4_in[3] ,
         \SB1_0_2/Component_Function_0/NAND4_in[2] ,
         \SB1_0_2/Component_Function_0/NAND4_in[1] ,
         \SB1_0_2/Component_Function_0/NAND4_in[0] ,
         \SB1_0_2/Component_Function_1/NAND4_in[2] ,
         \SB1_0_2/Component_Function_1/NAND4_in[1] ,
         \SB1_0_2/Component_Function_1/NAND4_in[0] ,
         \SB1_0_2/Component_Function_5/NAND4_in[3] ,
         \SB1_0_2/Component_Function_5/NAND4_in[2] ,
         \SB1_0_2/Component_Function_5/NAND4_in[1] ,
         \SB1_0_2/Component_Function_5/NAND4_in[0] ,
         \SB1_0_3/Component_Function_0/NAND4_in[3] ,
         \SB1_0_3/Component_Function_0/NAND4_in[2] ,
         \SB1_0_3/Component_Function_0/NAND4_in[1] ,
         \SB1_0_3/Component_Function_0/NAND4_in[0] ,
         \SB1_0_3/Component_Function_1/NAND4_in[2] ,
         \SB1_0_3/Component_Function_1/NAND4_in[1] ,
         \SB1_0_3/Component_Function_1/NAND4_in[0] ,
         \SB1_0_3/Component_Function_5/NAND4_in[3] ,
         \SB1_0_3/Component_Function_5/NAND4_in[2] ,
         \SB1_0_3/Component_Function_5/NAND4_in[1] ,
         \SB1_0_4/Component_Function_0/NAND4_in[3] ,
         \SB1_0_4/Component_Function_0/NAND4_in[2] ,
         \SB1_0_4/Component_Function_0/NAND4_in[1] ,
         \SB1_0_4/Component_Function_0/NAND4_in[0] ,
         \SB1_0_4/Component_Function_1/NAND4_in[3] ,
         \SB1_0_4/Component_Function_1/NAND4_in[2] ,
         \SB1_0_4/Component_Function_1/NAND4_in[1] ,
         \SB1_0_4/Component_Function_1/NAND4_in[0] ,
         \SB1_0_4/Component_Function_5/NAND4_in[2] ,
         \SB1_0_4/Component_Function_5/NAND4_in[1] ,
         \SB1_0_4/Component_Function_5/NAND4_in[0] ,
         \SB1_0_5/Component_Function_0/NAND4_in[3] ,
         \SB1_0_5/Component_Function_0/NAND4_in[1] ,
         \SB1_0_5/Component_Function_0/NAND4_in[0] ,
         \SB1_0_5/Component_Function_1/NAND4_in[3] ,
         \SB1_0_5/Component_Function_1/NAND4_in[1] ,
         \SB1_0_5/Component_Function_1/NAND4_in[0] ,
         \SB1_0_5/Component_Function_5/NAND4_in[3] ,
         \SB1_0_5/Component_Function_5/NAND4_in[2] ,
         \SB1_0_5/Component_Function_5/NAND4_in[1] ,
         \SB1_0_5/Component_Function_5/NAND4_in[0] ,
         \SB1_0_6/Component_Function_0/NAND4_in[3] ,
         \SB1_0_6/Component_Function_0/NAND4_in[1] ,
         \SB1_0_6/Component_Function_0/NAND4_in[0] ,
         \SB1_0_6/Component_Function_1/NAND4_in[2] ,
         \SB1_0_6/Component_Function_1/NAND4_in[1] ,
         \SB1_0_6/Component_Function_1/NAND4_in[0] ,
         \SB1_0_6/Component_Function_5/NAND4_in[2] ,
         \SB1_0_6/Component_Function_5/NAND4_in[1] ,
         \SB1_0_7/Component_Function_0/NAND4_in[3] ,
         \SB1_0_7/Component_Function_0/NAND4_in[2] ,
         \SB1_0_7/Component_Function_0/NAND4_in[1] ,
         \SB1_0_7/Component_Function_0/NAND4_in[0] ,
         \SB1_0_7/Component_Function_1/NAND4_in[3] ,
         \SB1_0_7/Component_Function_1/NAND4_in[2] ,
         \SB1_0_7/Component_Function_1/NAND4_in[1] ,
         \SB1_0_7/Component_Function_1/NAND4_in[0] ,
         \SB1_0_7/Component_Function_5/NAND4_in[2] ,
         \SB1_0_7/Component_Function_5/NAND4_in[1] ,
         \SB1_0_7/Component_Function_5/NAND4_in[0] ,
         \SB1_0_8/Component_Function_0/NAND4_in[2] ,
         \SB1_0_8/Component_Function_0/NAND4_in[1] ,
         \SB1_0_8/Component_Function_0/NAND4_in[0] ,
         \SB1_0_8/Component_Function_1/NAND4_in[3] ,
         \SB1_0_8/Component_Function_1/NAND4_in[2] ,
         \SB1_0_8/Component_Function_1/NAND4_in[1] ,
         \SB1_0_8/Component_Function_1/NAND4_in[0] ,
         \SB1_0_8/Component_Function_5/NAND4_in[1] ,
         \SB1_0_8/Component_Function_5/NAND4_in[0] ,
         \SB1_0_9/Component_Function_0/NAND4_in[2] ,
         \SB1_0_9/Component_Function_0/NAND4_in[1] ,
         \SB1_0_9/Component_Function_0/NAND4_in[0] ,
         \SB1_0_9/Component_Function_1/NAND4_in[3] ,
         \SB1_0_9/Component_Function_1/NAND4_in[2] ,
         \SB1_0_9/Component_Function_1/NAND4_in[1] ,
         \SB1_0_9/Component_Function_1/NAND4_in[0] ,
         \SB1_0_9/Component_Function_5/NAND4_in[3] ,
         \SB1_0_9/Component_Function_5/NAND4_in[2] ,
         \SB1_0_9/Component_Function_5/NAND4_in[1] ,
         \SB1_0_9/Component_Function_5/NAND4_in[0] ,
         \SB1_0_10/Component_Function_0/NAND4_in[3] ,
         \SB1_0_10/Component_Function_0/NAND4_in[2] ,
         \SB1_0_10/Component_Function_0/NAND4_in[1] ,
         \SB1_0_10/Component_Function_0/NAND4_in[0] ,
         \SB1_0_10/Component_Function_1/NAND4_in[3] ,
         \SB1_0_10/Component_Function_1/NAND4_in[2] ,
         \SB1_0_10/Component_Function_1/NAND4_in[1] ,
         \SB1_0_10/Component_Function_1/NAND4_in[0] ,
         \SB1_0_10/Component_Function_5/NAND4_in[1] ,
         \SB1_0_11/Component_Function_0/NAND4_in[3] ,
         \SB1_0_11/Component_Function_0/NAND4_in[2] ,
         \SB1_0_11/Component_Function_0/NAND4_in[1] ,
         \SB1_0_11/Component_Function_1/NAND4_in[3] ,
         \SB1_0_11/Component_Function_1/NAND4_in[2] ,
         \SB1_0_11/Component_Function_1/NAND4_in[1] ,
         \SB1_0_11/Component_Function_1/NAND4_in[0] ,
         \SB1_0_11/Component_Function_5/NAND4_in[3] ,
         \SB1_0_11/Component_Function_5/NAND4_in[2] ,
         \SB1_0_11/Component_Function_5/NAND4_in[0] ,
         \SB1_0_12/Component_Function_0/NAND4_in[3] ,
         \SB1_0_12/Component_Function_0/NAND4_in[2] ,
         \SB1_0_12/Component_Function_0/NAND4_in[1] ,
         \SB1_0_12/Component_Function_0/NAND4_in[0] ,
         \SB1_0_12/Component_Function_1/NAND4_in[3] ,
         \SB1_0_12/Component_Function_1/NAND4_in[2] ,
         \SB1_0_12/Component_Function_1/NAND4_in[1] ,
         \SB1_0_12/Component_Function_1/NAND4_in[0] ,
         \SB1_0_12/Component_Function_5/NAND4_in[1] ,
         \SB1_0_12/Component_Function_5/NAND4_in[0] ,
         \SB1_0_13/Component_Function_0/NAND4_in[3] ,
         \SB1_0_13/Component_Function_0/NAND4_in[2] ,
         \SB1_0_13/Component_Function_0/NAND4_in[1] ,
         \SB1_0_13/Component_Function_0/NAND4_in[0] ,
         \SB1_0_13/Component_Function_1/NAND4_in[3] ,
         \SB1_0_13/Component_Function_1/NAND4_in[2] ,
         \SB1_0_13/Component_Function_1/NAND4_in[1] ,
         \SB1_0_13/Component_Function_1/NAND4_in[0] ,
         \SB1_0_13/Component_Function_5/NAND4_in[3] ,
         \SB1_0_13/Component_Function_5/NAND4_in[2] ,
         \SB1_0_13/Component_Function_5/NAND4_in[1] ,
         \SB1_0_13/Component_Function_5/NAND4_in[0] ,
         \SB1_0_14/Component_Function_0/NAND4_in[3] ,
         \SB1_0_14/Component_Function_0/NAND4_in[1] ,
         \SB1_0_14/Component_Function_1/NAND4_in[3] ,
         \SB1_0_14/Component_Function_1/NAND4_in[2] ,
         \SB1_0_14/Component_Function_1/NAND4_in[1] ,
         \SB1_0_14/Component_Function_1/NAND4_in[0] ,
         \SB1_0_14/Component_Function_5/NAND4_in[2] ,
         \SB1_0_14/Component_Function_5/NAND4_in[1] ,
         \SB1_0_15/Component_Function_0/NAND4_in[3] ,
         \SB1_0_15/Component_Function_0/NAND4_in[2] ,
         \SB1_0_15/Component_Function_0/NAND4_in[1] ,
         \SB1_0_15/Component_Function_0/NAND4_in[0] ,
         \SB1_0_15/Component_Function_1/NAND4_in[3] ,
         \SB1_0_15/Component_Function_1/NAND4_in[2] ,
         \SB1_0_15/Component_Function_1/NAND4_in[1] ,
         \SB1_0_15/Component_Function_5/NAND4_in[1] ,
         \SB1_0_15/Component_Function_5/NAND4_in[0] ,
         \SB1_0_16/Component_Function_0/NAND4_in[3] ,
         \SB1_0_16/Component_Function_0/NAND4_in[2] ,
         \SB1_0_16/Component_Function_0/NAND4_in[1] ,
         \SB1_0_16/Component_Function_0/NAND4_in[0] ,
         \SB1_0_16/Component_Function_1/NAND4_in[3] ,
         \SB1_0_16/Component_Function_1/NAND4_in[2] ,
         \SB1_0_16/Component_Function_1/NAND4_in[1] ,
         \SB1_0_16/Component_Function_1/NAND4_in[0] ,
         \SB1_0_16/Component_Function_5/NAND4_in[2] ,
         \SB1_0_16/Component_Function_5/NAND4_in[1] ,
         \SB1_0_16/Component_Function_5/NAND4_in[0] ,
         \SB1_0_17/Component_Function_0/NAND4_in[3] ,
         \SB1_0_17/Component_Function_0/NAND4_in[2] ,
         \SB1_0_17/Component_Function_0/NAND4_in[1] ,
         \SB1_0_17/Component_Function_0/NAND4_in[0] ,
         \SB1_0_17/Component_Function_1/NAND4_in[3] ,
         \SB1_0_17/Component_Function_1/NAND4_in[2] ,
         \SB1_0_17/Component_Function_1/NAND4_in[1] ,
         \SB1_0_17/Component_Function_1/NAND4_in[0] ,
         \SB1_0_17/Component_Function_5/NAND4_in[3] ,
         \SB1_0_17/Component_Function_5/NAND4_in[2] ,
         \SB1_0_17/Component_Function_5/NAND4_in[1] ,
         \SB1_0_17/Component_Function_5/NAND4_in[0] ,
         \SB1_0_18/Component_Function_0/NAND4_in[3] ,
         \SB1_0_18/Component_Function_0/NAND4_in[2] ,
         \SB1_0_18/Component_Function_0/NAND4_in[1] ,
         \SB1_0_18/Component_Function_0/NAND4_in[0] ,
         \SB1_0_18/Component_Function_1/NAND4_in[3] ,
         \SB1_0_18/Component_Function_1/NAND4_in[0] ,
         \SB1_0_18/Component_Function_5/NAND4_in[2] ,
         \SB1_0_18/Component_Function_5/NAND4_in[1] ,
         \SB1_0_18/Component_Function_5/NAND4_in[0] ,
         \SB1_0_19/Component_Function_0/NAND4_in[2] ,
         \SB1_0_19/Component_Function_0/NAND4_in[1] ,
         \SB1_0_19/Component_Function_0/NAND4_in[0] ,
         \SB1_0_19/Component_Function_1/NAND4_in[3] ,
         \SB1_0_19/Component_Function_1/NAND4_in[2] ,
         \SB1_0_19/Component_Function_1/NAND4_in[1] ,
         \SB1_0_19/Component_Function_5/NAND4_in[3] ,
         \SB1_0_19/Component_Function_5/NAND4_in[1] ,
         \SB1_0_19/Component_Function_5/NAND4_in[0] ,
         \SB1_0_20/Component_Function_0/NAND4_in[3] ,
         \SB1_0_20/Component_Function_0/NAND4_in[2] ,
         \SB1_0_20/Component_Function_0/NAND4_in[1] ,
         \SB1_0_20/Component_Function_0/NAND4_in[0] ,
         \SB1_0_20/Component_Function_1/NAND4_in[2] ,
         \SB1_0_20/Component_Function_1/NAND4_in[1] ,
         \SB1_0_20/Component_Function_1/NAND4_in[0] ,
         \SB1_0_20/Component_Function_5/NAND4_in[3] ,
         \SB1_0_20/Component_Function_5/NAND4_in[2] ,
         \SB1_0_20/Component_Function_5/NAND4_in[1] ,
         \SB1_0_20/Component_Function_5/NAND4_in[0] ,
         \SB1_0_21/Component_Function_0/NAND4_in[3] ,
         \SB1_0_21/Component_Function_0/NAND4_in[2] ,
         \SB1_0_21/Component_Function_0/NAND4_in[1] ,
         \SB1_0_21/Component_Function_0/NAND4_in[0] ,
         \SB1_0_21/Component_Function_1/NAND4_in[3] ,
         \SB1_0_21/Component_Function_1/NAND4_in[2] ,
         \SB1_0_21/Component_Function_1/NAND4_in[1] ,
         \SB1_0_21/Component_Function_1/NAND4_in[0] ,
         \SB1_0_21/Component_Function_5/NAND4_in[3] ,
         \SB1_0_21/Component_Function_5/NAND4_in[2] ,
         \SB1_0_21/Component_Function_5/NAND4_in[1] ,
         \SB1_0_21/Component_Function_5/NAND4_in[0] ,
         \SB1_0_22/Component_Function_0/NAND4_in[2] ,
         \SB1_0_22/Component_Function_0/NAND4_in[1] ,
         \SB1_0_22/Component_Function_0/NAND4_in[0] ,
         \SB1_0_22/Component_Function_1/NAND4_in[3] ,
         \SB1_0_22/Component_Function_1/NAND4_in[2] ,
         \SB1_0_22/Component_Function_1/NAND4_in[1] ,
         \SB1_0_22/Component_Function_1/NAND4_in[0] ,
         \SB1_0_22/Component_Function_5/NAND4_in[1] ,
         \SB1_0_22/Component_Function_5/NAND4_in[0] ,
         \SB1_0_23/Component_Function_0/NAND4_in[3] ,
         \SB1_0_23/Component_Function_0/NAND4_in[2] ,
         \SB1_0_23/Component_Function_0/NAND4_in[1] ,
         \SB1_0_23/Component_Function_0/NAND4_in[0] ,
         \SB1_0_23/Component_Function_1/NAND4_in[1] ,
         \SB1_0_23/Component_Function_1/NAND4_in[0] ,
         \SB1_0_23/Component_Function_5/NAND4_in[3] ,
         \SB1_0_23/Component_Function_5/NAND4_in[2] ,
         \SB1_0_23/Component_Function_5/NAND4_in[1] ,
         \SB1_0_23/Component_Function_5/NAND4_in[0] ,
         \SB1_0_24/Component_Function_0/NAND4_in[3] ,
         \SB1_0_24/Component_Function_0/NAND4_in[2] ,
         \SB1_0_24/Component_Function_0/NAND4_in[1] ,
         \SB1_0_24/Component_Function_1/NAND4_in[2] ,
         \SB1_0_24/Component_Function_1/NAND4_in[1] ,
         \SB1_0_24/Component_Function_1/NAND4_in[0] ,
         \SB1_0_24/Component_Function_5/NAND4_in[3] ,
         \SB1_0_24/Component_Function_5/NAND4_in[2] ,
         \SB1_0_24/Component_Function_5/NAND4_in[1] ,
         \SB1_0_24/Component_Function_5/NAND4_in[0] ,
         \SB1_0_25/Component_Function_0/NAND4_in[1] ,
         \SB1_0_25/Component_Function_0/NAND4_in[0] ,
         \SB1_0_25/Component_Function_1/NAND4_in[3] ,
         \SB1_0_25/Component_Function_1/NAND4_in[1] ,
         \SB1_0_25/Component_Function_1/NAND4_in[0] ,
         \SB1_0_25/Component_Function_5/NAND4_in[3] ,
         \SB1_0_25/Component_Function_5/NAND4_in[2] ,
         \SB1_0_25/Component_Function_5/NAND4_in[0] ,
         \SB1_0_26/Component_Function_0/NAND4_in[3] ,
         \SB1_0_26/Component_Function_0/NAND4_in[2] ,
         \SB1_0_26/Component_Function_0/NAND4_in[1] ,
         \SB1_0_26/Component_Function_0/NAND4_in[0] ,
         \SB1_0_26/Component_Function_1/NAND4_in[3] ,
         \SB1_0_26/Component_Function_1/NAND4_in[1] ,
         \SB1_0_26/Component_Function_1/NAND4_in[0] ,
         \SB1_0_26/Component_Function_5/NAND4_in[2] ,
         \SB1_0_26/Component_Function_5/NAND4_in[1] ,
         \SB1_0_27/Component_Function_0/NAND4_in[3] ,
         \SB1_0_27/Component_Function_0/NAND4_in[2] ,
         \SB1_0_27/Component_Function_0/NAND4_in[1] ,
         \SB1_0_27/Component_Function_0/NAND4_in[0] ,
         \SB1_0_27/Component_Function_1/NAND4_in[2] ,
         \SB1_0_27/Component_Function_1/NAND4_in[1] ,
         \SB1_0_27/Component_Function_1/NAND4_in[0] ,
         \SB1_0_27/Component_Function_5/NAND4_in[3] ,
         \SB1_0_27/Component_Function_5/NAND4_in[2] ,
         \SB1_0_27/Component_Function_5/NAND4_in[0] ,
         \SB1_0_28/Component_Function_0/NAND4_in[2] ,
         \SB1_0_28/Component_Function_0/NAND4_in[1] ,
         \SB1_0_28/Component_Function_0/NAND4_in[0] ,
         \SB1_0_28/Component_Function_1/NAND4_in[3] ,
         \SB1_0_28/Component_Function_1/NAND4_in[2] ,
         \SB1_0_28/Component_Function_1/NAND4_in[1] ,
         \SB1_0_28/Component_Function_1/NAND4_in[0] ,
         \SB1_0_28/Component_Function_5/NAND4_in[2] ,
         \SB1_0_28/Component_Function_5/NAND4_in[1] ,
         \SB1_0_28/Component_Function_5/NAND4_in[0] ,
         \SB1_0_29/Component_Function_0/NAND4_in[3] ,
         \SB1_0_29/Component_Function_0/NAND4_in[2] ,
         \SB1_0_29/Component_Function_0/NAND4_in[1] ,
         \SB1_0_29/Component_Function_0/NAND4_in[0] ,
         \SB1_0_29/Component_Function_1/NAND4_in[3] ,
         \SB1_0_29/Component_Function_1/NAND4_in[2] ,
         \SB1_0_29/Component_Function_1/NAND4_in[1] ,
         \SB1_0_29/Component_Function_1/NAND4_in[0] ,
         \SB1_0_29/Component_Function_5/NAND4_in[2] ,
         \SB1_0_29/Component_Function_5/NAND4_in[1] ,
         \SB1_0_29/Component_Function_5/NAND4_in[0] ,
         \SB1_0_30/Component_Function_0/NAND4_in[3] ,
         \SB1_0_30/Component_Function_0/NAND4_in[2] ,
         \SB1_0_30/Component_Function_0/NAND4_in[1] ,
         \SB1_0_30/Component_Function_0/NAND4_in[0] ,
         \SB1_0_30/Component_Function_1/NAND4_in[3] ,
         \SB1_0_30/Component_Function_1/NAND4_in[2] ,
         \SB1_0_30/Component_Function_1/NAND4_in[1] ,
         \SB1_0_30/Component_Function_1/NAND4_in[0] ,
         \SB1_0_30/Component_Function_5/NAND4_in[2] ,
         \SB1_0_30/Component_Function_5/NAND4_in[1] ,
         \SB1_0_30/Component_Function_5/NAND4_in[0] ,
         \SB1_0_31/Component_Function_0/NAND4_in[2] ,
         \SB1_0_31/Component_Function_0/NAND4_in[1] ,
         \SB1_0_31/Component_Function_0/NAND4_in[0] ,
         \SB1_0_31/Component_Function_1/NAND4_in[3] ,
         \SB1_0_31/Component_Function_1/NAND4_in[2] ,
         \SB1_0_31/Component_Function_1/NAND4_in[1] ,
         \SB1_0_31/Component_Function_1/NAND4_in[0] ,
         \SB1_0_31/Component_Function_5/NAND4_in[2] ,
         \SB1_0_31/Component_Function_5/NAND4_in[0] ,
         \SB2_0_0/Component_Function_0/NAND4_in[1] ,
         \SB2_0_0/Component_Function_0/NAND4_in[0] ,
         \SB2_0_0/Component_Function_1/NAND4_in[3] ,
         \SB2_0_0/Component_Function_1/NAND4_in[1] ,
         \SB2_0_0/Component_Function_1/NAND4_in[0] ,
         \SB2_0_0/Component_Function_5/NAND4_in[1] ,
         \SB2_0_0/Component_Function_5/NAND4_in[0] ,
         \SB2_0_1/Component_Function_0/NAND4_in[3] ,
         \SB2_0_1/Component_Function_0/NAND4_in[1] ,
         \SB2_0_1/Component_Function_0/NAND4_in[0] ,
         \SB2_0_1/Component_Function_1/NAND4_in[2] ,
         \SB2_0_1/Component_Function_1/NAND4_in[1] ,
         \SB2_0_1/Component_Function_1/NAND4_in[0] ,
         \SB2_0_1/Component_Function_5/NAND4_in[2] ,
         \SB2_0_1/Component_Function_5/NAND4_in[0] ,
         \SB2_0_2/Component_Function_0/NAND4_in[3] ,
         \SB2_0_2/Component_Function_0/NAND4_in[2] ,
         \SB2_0_2/Component_Function_0/NAND4_in[1] ,
         \SB2_0_2/Component_Function_0/NAND4_in[0] ,
         \SB2_0_2/Component_Function_1/NAND4_in[3] ,
         \SB2_0_2/Component_Function_1/NAND4_in[2] ,
         \SB2_0_2/Component_Function_1/NAND4_in[1] ,
         \SB2_0_2/Component_Function_1/NAND4_in[0] ,
         \SB2_0_2/Component_Function_5/NAND4_in[3] ,
         \SB2_0_2/Component_Function_5/NAND4_in[2] ,
         \SB2_0_2/Component_Function_5/NAND4_in[0] ,
         \SB2_0_3/Component_Function_0/NAND4_in[3] ,
         \SB2_0_3/Component_Function_0/NAND4_in[2] ,
         \SB2_0_3/Component_Function_0/NAND4_in[1] ,
         \SB2_0_3/Component_Function_0/NAND4_in[0] ,
         \SB2_0_3/Component_Function_1/NAND4_in[3] ,
         \SB2_0_3/Component_Function_1/NAND4_in[1] ,
         \SB2_0_3/Component_Function_1/NAND4_in[0] ,
         \SB2_0_3/Component_Function_5/NAND4_in[3] ,
         \SB2_0_3/Component_Function_5/NAND4_in[2] ,
         \SB2_0_3/Component_Function_5/NAND4_in[1] ,
         \SB2_0_3/Component_Function_5/NAND4_in[0] ,
         \SB2_0_4/Component_Function_0/NAND4_in[2] ,
         \SB2_0_4/Component_Function_0/NAND4_in[1] ,
         \SB2_0_4/Component_Function_0/NAND4_in[0] ,
         \SB2_0_4/Component_Function_1/NAND4_in[3] ,
         \SB2_0_4/Component_Function_1/NAND4_in[2] ,
         \SB2_0_4/Component_Function_1/NAND4_in[1] ,
         \SB2_0_4/Component_Function_1/NAND4_in[0] ,
         \SB2_0_4/Component_Function_5/NAND4_in[2] ,
         \SB2_0_4/Component_Function_5/NAND4_in[1] ,
         \SB2_0_4/Component_Function_5/NAND4_in[0] ,
         \SB2_0_5/Component_Function_0/NAND4_in[2] ,
         \SB2_0_5/Component_Function_0/NAND4_in[1] ,
         \SB2_0_5/Component_Function_0/NAND4_in[0] ,
         \SB2_0_5/Component_Function_1/NAND4_in[3] ,
         \SB2_0_5/Component_Function_1/NAND4_in[2] ,
         \SB2_0_5/Component_Function_1/NAND4_in[1] ,
         \SB2_0_5/Component_Function_1/NAND4_in[0] ,
         \SB2_0_5/Component_Function_5/NAND4_in[3] ,
         \SB2_0_5/Component_Function_5/NAND4_in[1] ,
         \SB2_0_5/Component_Function_5/NAND4_in[0] ,
         \SB2_0_6/Component_Function_0/NAND4_in[1] ,
         \SB2_0_6/Component_Function_1/NAND4_in[3] ,
         \SB2_0_6/Component_Function_1/NAND4_in[2] ,
         \SB2_0_6/Component_Function_1/NAND4_in[1] ,
         \SB2_0_6/Component_Function_1/NAND4_in[0] ,
         \SB2_0_6/Component_Function_5/NAND4_in[2] ,
         \SB2_0_6/Component_Function_5/NAND4_in[0] ,
         \SB2_0_7/Component_Function_0/NAND4_in[2] ,
         \SB2_0_7/Component_Function_0/NAND4_in[1] ,
         \SB2_0_7/Component_Function_0/NAND4_in[0] ,
         \SB2_0_7/Component_Function_1/NAND4_in[3] ,
         \SB2_0_7/Component_Function_1/NAND4_in[2] ,
         \SB2_0_7/Component_Function_1/NAND4_in[1] ,
         \SB2_0_7/Component_Function_1/NAND4_in[0] ,
         \SB2_0_7/Component_Function_5/NAND4_in[0] ,
         \SB2_0_8/Component_Function_0/NAND4_in[3] ,
         \SB2_0_8/Component_Function_0/NAND4_in[2] ,
         \SB2_0_8/Component_Function_0/NAND4_in[1] ,
         \SB2_0_8/Component_Function_0/NAND4_in[0] ,
         \SB2_0_8/Component_Function_1/NAND4_in[3] ,
         \SB2_0_8/Component_Function_1/NAND4_in[2] ,
         \SB2_0_8/Component_Function_1/NAND4_in[1] ,
         \SB2_0_8/Component_Function_1/NAND4_in[0] ,
         \SB2_0_8/Component_Function_5/NAND4_in[1] ,
         \SB2_0_8/Component_Function_5/NAND4_in[0] ,
         \SB2_0_9/Component_Function_0/NAND4_in[2] ,
         \SB2_0_9/Component_Function_0/NAND4_in[1] ,
         \SB2_0_9/Component_Function_0/NAND4_in[0] ,
         \SB2_0_9/Component_Function_1/NAND4_in[3] ,
         \SB2_0_9/Component_Function_1/NAND4_in[2] ,
         \SB2_0_9/Component_Function_1/NAND4_in[1] ,
         \SB2_0_9/Component_Function_1/NAND4_in[0] ,
         \SB2_0_9/Component_Function_5/NAND4_in[2] ,
         \SB2_0_9/Component_Function_5/NAND4_in[0] ,
         \SB2_0_10/Component_Function_0/NAND4_in[2] ,
         \SB2_0_10/Component_Function_0/NAND4_in[1] ,
         \SB2_0_10/Component_Function_0/NAND4_in[0] ,
         \SB2_0_10/Component_Function_1/NAND4_in[3] ,
         \SB2_0_10/Component_Function_1/NAND4_in[2] ,
         \SB2_0_10/Component_Function_1/NAND4_in[1] ,
         \SB2_0_10/Component_Function_1/NAND4_in[0] ,
         \SB2_0_10/Component_Function_5/NAND4_in[3] ,
         \SB2_0_10/Component_Function_5/NAND4_in[1] ,
         \SB2_0_10/Component_Function_5/NAND4_in[0] ,
         \SB2_0_11/Component_Function_0/NAND4_in[2] ,
         \SB2_0_11/Component_Function_0/NAND4_in[1] ,
         \SB2_0_11/Component_Function_0/NAND4_in[0] ,
         \SB2_0_11/Component_Function_1/NAND4_in[3] ,
         \SB2_0_11/Component_Function_1/NAND4_in[2] ,
         \SB2_0_11/Component_Function_1/NAND4_in[1] ,
         \SB2_0_11/Component_Function_1/NAND4_in[0] ,
         \SB2_0_11/Component_Function_5/NAND4_in[2] ,
         \SB2_0_11/Component_Function_5/NAND4_in[0] ,
         \SB2_0_12/Component_Function_0/NAND4_in[3] ,
         \SB2_0_12/Component_Function_0/NAND4_in[2] ,
         \SB2_0_12/Component_Function_0/NAND4_in[0] ,
         \SB2_0_12/Component_Function_1/NAND4_in[3] ,
         \SB2_0_12/Component_Function_1/NAND4_in[2] ,
         \SB2_0_12/Component_Function_1/NAND4_in[1] ,
         \SB2_0_12/Component_Function_1/NAND4_in[0] ,
         \SB2_0_12/Component_Function_5/NAND4_in[2] ,
         \SB2_0_12/Component_Function_5/NAND4_in[1] ,
         \SB2_0_12/Component_Function_5/NAND4_in[0] ,
         \SB2_0_13/Component_Function_0/NAND4_in[2] ,
         \SB2_0_13/Component_Function_0/NAND4_in[1] ,
         \SB2_0_13/Component_Function_0/NAND4_in[0] ,
         \SB2_0_13/Component_Function_1/NAND4_in[3] ,
         \SB2_0_13/Component_Function_1/NAND4_in[2] ,
         \SB2_0_13/Component_Function_1/NAND4_in[1] ,
         \SB2_0_13/Component_Function_1/NAND4_in[0] ,
         \SB2_0_13/Component_Function_5/NAND4_in[1] ,
         \SB2_0_13/Component_Function_5/NAND4_in[0] ,
         \SB2_0_14/Component_Function_0/NAND4_in[3] ,
         \SB2_0_14/Component_Function_0/NAND4_in[2] ,
         \SB2_0_14/Component_Function_0/NAND4_in[1] ,
         \SB2_0_14/Component_Function_0/NAND4_in[0] ,
         \SB2_0_14/Component_Function_1/NAND4_in[3] ,
         \SB2_0_14/Component_Function_1/NAND4_in[2] ,
         \SB2_0_14/Component_Function_1/NAND4_in[1] ,
         \SB2_0_14/Component_Function_1/NAND4_in[0] ,
         \SB2_0_14/Component_Function_5/NAND4_in[3] ,
         \SB2_0_14/Component_Function_5/NAND4_in[2] ,
         \SB2_0_14/Component_Function_5/NAND4_in[1] ,
         \SB2_0_14/Component_Function_5/NAND4_in[0] ,
         \SB2_0_15/Component_Function_0/NAND4_in[3] ,
         \SB2_0_15/Component_Function_0/NAND4_in[2] ,
         \SB2_0_15/Component_Function_0/NAND4_in[1] ,
         \SB2_0_15/Component_Function_0/NAND4_in[0] ,
         \SB2_0_15/Component_Function_1/NAND4_in[3] ,
         \SB2_0_15/Component_Function_5/NAND4_in[0] ,
         \SB2_0_16/Component_Function_0/NAND4_in[3] ,
         \SB2_0_16/Component_Function_0/NAND4_in[2] ,
         \SB2_0_16/Component_Function_0/NAND4_in[1] ,
         \SB2_0_16/Component_Function_0/NAND4_in[0] ,
         \SB2_0_16/Component_Function_1/NAND4_in[3] ,
         \SB2_0_16/Component_Function_1/NAND4_in[2] ,
         \SB2_0_16/Component_Function_1/NAND4_in[1] ,
         \SB2_0_16/Component_Function_1/NAND4_in[0] ,
         \SB2_0_16/Component_Function_5/NAND4_in[2] ,
         \SB2_0_16/Component_Function_5/NAND4_in[1] ,
         \SB2_0_16/Component_Function_5/NAND4_in[0] ,
         \SB2_0_17/Component_Function_0/NAND4_in[3] ,
         \SB2_0_17/Component_Function_0/NAND4_in[2] ,
         \SB2_0_17/Component_Function_0/NAND4_in[1] ,
         \SB2_0_17/Component_Function_0/NAND4_in[0] ,
         \SB2_0_17/Component_Function_1/NAND4_in[3] ,
         \SB2_0_17/Component_Function_1/NAND4_in[1] ,
         \SB2_0_17/Component_Function_1/NAND4_in[0] ,
         \SB2_0_17/Component_Function_5/NAND4_in[3] ,
         \SB2_0_17/Component_Function_5/NAND4_in[2] ,
         \SB2_0_17/Component_Function_5/NAND4_in[1] ,
         \SB2_0_17/Component_Function_5/NAND4_in[0] ,
         \SB2_0_18/Component_Function_0/NAND4_in[2] ,
         \SB2_0_18/Component_Function_0/NAND4_in[1] ,
         \SB2_0_18/Component_Function_0/NAND4_in[0] ,
         \SB2_0_18/Component_Function_1/NAND4_in[2] ,
         \SB2_0_18/Component_Function_1/NAND4_in[1] ,
         \SB2_0_18/Component_Function_1/NAND4_in[0] ,
         \SB2_0_18/Component_Function_5/NAND4_in[3] ,
         \SB2_0_18/Component_Function_5/NAND4_in[1] ,
         \SB2_0_18/Component_Function_5/NAND4_in[0] ,
         \SB2_0_19/Component_Function_0/NAND4_in[1] ,
         \SB2_0_19/Component_Function_0/NAND4_in[0] ,
         \SB2_0_19/Component_Function_1/NAND4_in[2] ,
         \SB2_0_19/Component_Function_1/NAND4_in[1] ,
         \SB2_0_19/Component_Function_1/NAND4_in[0] ,
         \SB2_0_19/Component_Function_5/NAND4_in[3] ,
         \SB2_0_19/Component_Function_5/NAND4_in[2] ,
         \SB2_0_19/Component_Function_5/NAND4_in[1] ,
         \SB2_0_19/Component_Function_5/NAND4_in[0] ,
         \SB2_0_20/Component_Function_0/NAND4_in[3] ,
         \SB2_0_20/Component_Function_0/NAND4_in[2] ,
         \SB2_0_20/Component_Function_0/NAND4_in[1] ,
         \SB2_0_20/Component_Function_0/NAND4_in[0] ,
         \SB2_0_20/Component_Function_1/NAND4_in[3] ,
         \SB2_0_20/Component_Function_1/NAND4_in[2] ,
         \SB2_0_20/Component_Function_1/NAND4_in[1] ,
         \SB2_0_20/Component_Function_1/NAND4_in[0] ,
         \SB2_0_20/Component_Function_5/NAND4_in[1] ,
         \SB2_0_20/Component_Function_5/NAND4_in[0] ,
         \SB2_0_21/Component_Function_0/NAND4_in[2] ,
         \SB2_0_21/Component_Function_0/NAND4_in[1] ,
         \SB2_0_21/Component_Function_0/NAND4_in[0] ,
         \SB2_0_21/Component_Function_1/NAND4_in[3] ,
         \SB2_0_21/Component_Function_1/NAND4_in[2] ,
         \SB2_0_21/Component_Function_1/NAND4_in[1] ,
         \SB2_0_21/Component_Function_1/NAND4_in[0] ,
         \SB2_0_21/Component_Function_5/NAND4_in[3] ,
         \SB2_0_21/Component_Function_5/NAND4_in[2] ,
         \SB2_0_21/Component_Function_5/NAND4_in[0] ,
         \SB2_0_22/Component_Function_0/NAND4_in[2] ,
         \SB2_0_22/Component_Function_0/NAND4_in[0] ,
         \SB2_0_22/Component_Function_1/NAND4_in[3] ,
         \SB2_0_22/Component_Function_1/NAND4_in[2] ,
         \SB2_0_22/Component_Function_1/NAND4_in[1] ,
         \SB2_0_22/Component_Function_5/NAND4_in[3] ,
         \SB2_0_22/Component_Function_5/NAND4_in[2] ,
         \SB2_0_22/Component_Function_5/NAND4_in[1] ,
         \SB2_0_22/Component_Function_5/NAND4_in[0] ,
         \SB2_0_23/Component_Function_0/NAND4_in[3] ,
         \SB2_0_23/Component_Function_0/NAND4_in[2] ,
         \SB2_0_23/Component_Function_0/NAND4_in[0] ,
         \SB2_0_23/Component_Function_1/NAND4_in[3] ,
         \SB2_0_23/Component_Function_1/NAND4_in[2] ,
         \SB2_0_23/Component_Function_1/NAND4_in[1] ,
         \SB2_0_23/Component_Function_5/NAND4_in[3] ,
         \SB2_0_23/Component_Function_5/NAND4_in[0] ,
         \SB2_0_24/Component_Function_0/NAND4_in[3] ,
         \SB2_0_24/Component_Function_0/NAND4_in[2] ,
         \SB2_0_24/Component_Function_0/NAND4_in[1] ,
         \SB2_0_24/Component_Function_0/NAND4_in[0] ,
         \SB2_0_24/Component_Function_1/NAND4_in[3] ,
         \SB2_0_24/Component_Function_1/NAND4_in[2] ,
         \SB2_0_24/Component_Function_1/NAND4_in[1] ,
         \SB2_0_24/Component_Function_1/NAND4_in[0] ,
         \SB2_0_24/Component_Function_5/NAND4_in[3] ,
         \SB2_0_25/Component_Function_0/NAND4_in[1] ,
         \SB2_0_25/Component_Function_0/NAND4_in[0] ,
         \SB2_0_25/Component_Function_1/NAND4_in[3] ,
         \SB2_0_25/Component_Function_1/NAND4_in[2] ,
         \SB2_0_25/Component_Function_1/NAND4_in[1] ,
         \SB2_0_25/Component_Function_1/NAND4_in[0] ,
         \SB2_0_25/Component_Function_5/NAND4_in[3] ,
         \SB2_0_25/Component_Function_5/NAND4_in[1] ,
         \SB2_0_25/Component_Function_5/NAND4_in[0] ,
         \SB2_0_26/Component_Function_0/NAND4_in[3] ,
         \SB2_0_26/Component_Function_0/NAND4_in[2] ,
         \SB2_0_26/Component_Function_0/NAND4_in[1] ,
         \SB2_0_26/Component_Function_0/NAND4_in[0] ,
         \SB2_0_26/Component_Function_1/NAND4_in[2] ,
         \SB2_0_26/Component_Function_1/NAND4_in[1] ,
         \SB2_0_26/Component_Function_1/NAND4_in[0] ,
         \SB2_0_26/Component_Function_5/NAND4_in[3] ,
         \SB2_0_26/Component_Function_5/NAND4_in[2] ,
         \SB2_0_26/Component_Function_5/NAND4_in[1] ,
         \SB2_0_26/Component_Function_5/NAND4_in[0] ,
         \SB2_0_27/Component_Function_0/NAND4_in[3] ,
         \SB2_0_27/Component_Function_0/NAND4_in[2] ,
         \SB2_0_27/Component_Function_0/NAND4_in[0] ,
         \SB2_0_27/Component_Function_1/NAND4_in[2] ,
         \SB2_0_27/Component_Function_1/NAND4_in[1] ,
         \SB2_0_27/Component_Function_1/NAND4_in[0] ,
         \SB2_0_27/Component_Function_5/NAND4_in[2] ,
         \SB2_0_28/Component_Function_0/NAND4_in[3] ,
         \SB2_0_28/Component_Function_0/NAND4_in[2] ,
         \SB2_0_28/Component_Function_0/NAND4_in[1] ,
         \SB2_0_28/Component_Function_0/NAND4_in[0] ,
         \SB2_0_28/Component_Function_1/NAND4_in[3] ,
         \SB2_0_28/Component_Function_1/NAND4_in[2] ,
         \SB2_0_28/Component_Function_1/NAND4_in[1] ,
         \SB2_0_28/Component_Function_1/NAND4_in[0] ,
         \SB2_0_28/Component_Function_5/NAND4_in[3] ,
         \SB2_0_28/Component_Function_5/NAND4_in[1] ,
         \SB2_0_28/Component_Function_5/NAND4_in[0] ,
         \SB2_0_29/Component_Function_0/NAND4_in[3] ,
         \SB2_0_29/Component_Function_0/NAND4_in[1] ,
         \SB2_0_29/Component_Function_0/NAND4_in[0] ,
         \SB2_0_29/Component_Function_1/NAND4_in[3] ,
         \SB2_0_29/Component_Function_1/NAND4_in[2] ,
         \SB2_0_29/Component_Function_1/NAND4_in[1] ,
         \SB2_0_29/Component_Function_1/NAND4_in[0] ,
         \SB2_0_29/Component_Function_5/NAND4_in[3] ,
         \SB2_0_29/Component_Function_5/NAND4_in[2] ,
         \SB2_0_29/Component_Function_5/NAND4_in[1] ,
         \SB2_0_29/Component_Function_5/NAND4_in[0] ,
         \SB2_0_30/Component_Function_0/NAND4_in[1] ,
         \SB2_0_30/Component_Function_0/NAND4_in[0] ,
         \SB2_0_30/Component_Function_1/NAND4_in[3] ,
         \SB2_0_30/Component_Function_1/NAND4_in[2] ,
         \SB2_0_30/Component_Function_1/NAND4_in[1] ,
         \SB2_0_30/Component_Function_1/NAND4_in[0] ,
         \SB2_0_30/Component_Function_5/NAND4_in[3] ,
         \SB2_0_30/Component_Function_5/NAND4_in[1] ,
         \SB2_0_30/Component_Function_5/NAND4_in[0] ,
         \SB2_0_31/Component_Function_0/NAND4_in[3] ,
         \SB2_0_31/Component_Function_0/NAND4_in[2] ,
         \SB2_0_31/Component_Function_0/NAND4_in[0] ,
         \SB2_0_31/Component_Function_1/NAND4_in[3] ,
         \SB2_0_31/Component_Function_1/NAND4_in[2] ,
         \SB2_0_31/Component_Function_1/NAND4_in[1] ,
         \SB2_0_31/Component_Function_1/NAND4_in[0] ,
         \SB2_0_31/Component_Function_5/NAND4_in[2] ,
         \SB2_0_31/Component_Function_5/NAND4_in[0] ,
         \SB1_1_0/Component_Function_0/NAND4_in[3] ,
         \SB1_1_0/Component_Function_0/NAND4_in[2] ,
         \SB1_1_0/Component_Function_0/NAND4_in[1] ,
         \SB1_1_0/Component_Function_0/NAND4_in[0] ,
         \SB1_1_0/Component_Function_1/NAND4_in[3] ,
         \SB1_1_0/Component_Function_1/NAND4_in[2] ,
         \SB1_1_0/Component_Function_1/NAND4_in[1] ,
         \SB1_1_0/Component_Function_1/NAND4_in[0] ,
         \SB1_1_0/Component_Function_5/NAND4_in[3] ,
         \SB1_1_0/Component_Function_5/NAND4_in[0] ,
         \SB1_1_1/Component_Function_0/NAND4_in[3] ,
         \SB1_1_1/Component_Function_0/NAND4_in[2] ,
         \SB1_1_1/Component_Function_0/NAND4_in[1] ,
         \SB1_1_1/Component_Function_0/NAND4_in[0] ,
         \SB1_1_1/Component_Function_1/NAND4_in[3] ,
         \SB1_1_1/Component_Function_1/NAND4_in[2] ,
         \SB1_1_1/Component_Function_1/NAND4_in[1] ,
         \SB1_1_1/Component_Function_1/NAND4_in[0] ,
         \SB1_1_1/Component_Function_5/NAND4_in[3] ,
         \SB1_1_1/Component_Function_5/NAND4_in[2] ,
         \SB1_1_2/Component_Function_0/NAND4_in[2] ,
         \SB1_1_2/Component_Function_0/NAND4_in[1] ,
         \SB1_1_2/Component_Function_0/NAND4_in[0] ,
         \SB1_1_2/Component_Function_1/NAND4_in[3] ,
         \SB1_1_2/Component_Function_1/NAND4_in[1] ,
         \SB1_1_2/Component_Function_5/NAND4_in[2] ,
         \SB1_1_2/Component_Function_5/NAND4_in[0] ,
         \SB1_1_3/Component_Function_0/NAND4_in[3] ,
         \SB1_1_3/Component_Function_0/NAND4_in[2] ,
         \SB1_1_3/Component_Function_0/NAND4_in[1] ,
         \SB1_1_3/Component_Function_0/NAND4_in[0] ,
         \SB1_1_3/Component_Function_1/NAND4_in[0] ,
         \SB1_1_3/Component_Function_5/NAND4_in[1] ,
         \SB1_1_3/Component_Function_5/NAND4_in[0] ,
         \SB1_1_4/Component_Function_0/NAND4_in[3] ,
         \SB1_1_4/Component_Function_0/NAND4_in[2] ,
         \SB1_1_4/Component_Function_0/NAND4_in[1] ,
         \SB1_1_4/Component_Function_0/NAND4_in[0] ,
         \SB1_1_4/Component_Function_1/NAND4_in[2] ,
         \SB1_1_4/Component_Function_1/NAND4_in[1] ,
         \SB1_1_4/Component_Function_1/NAND4_in[0] ,
         \SB1_1_4/Component_Function_5/NAND4_in[0] ,
         \SB1_1_5/Component_Function_0/NAND4_in[3] ,
         \SB1_1_5/Component_Function_0/NAND4_in[2] ,
         \SB1_1_5/Component_Function_0/NAND4_in[1] ,
         \SB1_1_5/Component_Function_0/NAND4_in[0] ,
         \SB1_1_5/Component_Function_1/NAND4_in[3] ,
         \SB1_1_5/Component_Function_1/NAND4_in[2] ,
         \SB1_1_5/Component_Function_1/NAND4_in[1] ,
         \SB1_1_5/Component_Function_1/NAND4_in[0] ,
         \SB1_1_5/Component_Function_5/NAND4_in[1] ,
         \SB1_1_5/Component_Function_5/NAND4_in[0] ,
         \SB1_1_6/Component_Function_0/NAND4_in[1] ,
         \SB1_1_6/Component_Function_0/NAND4_in[0] ,
         \SB1_1_6/Component_Function_1/NAND4_in[2] ,
         \SB1_1_6/Component_Function_1/NAND4_in[1] ,
         \SB1_1_6/Component_Function_1/NAND4_in[0] ,
         \SB1_1_6/Component_Function_5/NAND4_in[3] ,
         \SB1_1_6/Component_Function_5/NAND4_in[2] ,
         \SB1_1_7/Component_Function_0/NAND4_in[2] ,
         \SB1_1_7/Component_Function_0/NAND4_in[1] ,
         \SB1_1_7/Component_Function_0/NAND4_in[0] ,
         \SB1_1_7/Component_Function_1/NAND4_in[3] ,
         \SB1_1_7/Component_Function_1/NAND4_in[2] ,
         \SB1_1_7/Component_Function_1/NAND4_in[1] ,
         \SB1_1_7/Component_Function_1/NAND4_in[0] ,
         \SB1_1_7/Component_Function_5/NAND4_in[2] ,
         \SB1_1_7/Component_Function_5/NAND4_in[1] ,
         \SB1_1_7/Component_Function_5/NAND4_in[0] ,
         \SB1_1_8/Component_Function_0/NAND4_in[3] ,
         \SB1_1_8/Component_Function_0/NAND4_in[1] ,
         \SB1_1_8/Component_Function_0/NAND4_in[0] ,
         \SB1_1_8/Component_Function_1/NAND4_in[3] ,
         \SB1_1_8/Component_Function_1/NAND4_in[2] ,
         \SB1_1_8/Component_Function_1/NAND4_in[1] ,
         \SB1_1_8/Component_Function_1/NAND4_in[0] ,
         \SB1_1_8/Component_Function_5/NAND4_in[1] ,
         \SB1_1_8/Component_Function_5/NAND4_in[0] ,
         \SB1_1_9/Component_Function_0/NAND4_in[3] ,
         \SB1_1_9/Component_Function_0/NAND4_in[1] ,
         \SB1_1_9/Component_Function_0/NAND4_in[0] ,
         \SB1_1_9/Component_Function_1/NAND4_in[3] ,
         \SB1_1_9/Component_Function_1/NAND4_in[2] ,
         \SB1_1_9/Component_Function_1/NAND4_in[1] ,
         \SB1_1_9/Component_Function_1/NAND4_in[0] ,
         \SB1_1_9/Component_Function_5/NAND4_in[2] ,
         \SB1_1_9/Component_Function_5/NAND4_in[0] ,
         \SB1_1_10/Component_Function_0/NAND4_in[3] ,
         \SB1_1_10/Component_Function_0/NAND4_in[2] ,
         \SB1_1_10/Component_Function_0/NAND4_in[1] ,
         \SB1_1_10/Component_Function_0/NAND4_in[0] ,
         \SB1_1_10/Component_Function_1/NAND4_in[3] ,
         \SB1_1_10/Component_Function_1/NAND4_in[2] ,
         \SB1_1_10/Component_Function_1/NAND4_in[1] ,
         \SB1_1_10/Component_Function_1/NAND4_in[0] ,
         \SB1_1_10/Component_Function_5/NAND4_in[1] ,
         \SB1_1_10/Component_Function_5/NAND4_in[0] ,
         \SB1_1_11/Component_Function_0/NAND4_in[3] ,
         \SB1_1_11/Component_Function_0/NAND4_in[1] ,
         \SB1_1_11/Component_Function_0/NAND4_in[0] ,
         \SB1_1_11/Component_Function_1/NAND4_in[2] ,
         \SB1_1_11/Component_Function_1/NAND4_in[1] ,
         \SB1_1_11/Component_Function_1/NAND4_in[0] ,
         \SB1_1_11/Component_Function_5/NAND4_in[3] ,
         \SB1_1_11/Component_Function_5/NAND4_in[1] ,
         \SB1_1_11/Component_Function_5/NAND4_in[0] ,
         \SB1_1_12/Component_Function_0/NAND4_in[3] ,
         \SB1_1_12/Component_Function_0/NAND4_in[2] ,
         \SB1_1_12/Component_Function_0/NAND4_in[1] ,
         \SB1_1_12/Component_Function_0/NAND4_in[0] ,
         \SB1_1_12/Component_Function_1/NAND4_in[2] ,
         \SB1_1_12/Component_Function_1/NAND4_in[1] ,
         \SB1_1_12/Component_Function_1/NAND4_in[0] ,
         \SB1_1_12/Component_Function_5/NAND4_in[2] ,
         \SB1_1_12/Component_Function_5/NAND4_in[1] ,
         \SB1_1_12/Component_Function_5/NAND4_in[0] ,
         \SB1_1_13/Component_Function_0/NAND4_in[3] ,
         \SB1_1_13/Component_Function_0/NAND4_in[2] ,
         \SB1_1_13/Component_Function_0/NAND4_in[1] ,
         \SB1_1_13/Component_Function_0/NAND4_in[0] ,
         \SB1_1_13/Component_Function_1/NAND4_in[3] ,
         \SB1_1_13/Component_Function_1/NAND4_in[2] ,
         \SB1_1_13/Component_Function_1/NAND4_in[1] ,
         \SB1_1_13/Component_Function_1/NAND4_in[0] ,
         \SB1_1_13/Component_Function_5/NAND4_in[2] ,
         \SB1_1_13/Component_Function_5/NAND4_in[1] ,
         \SB1_1_13/Component_Function_5/NAND4_in[0] ,
         \SB1_1_14/Component_Function_0/NAND4_in[3] ,
         \SB1_1_14/Component_Function_0/NAND4_in[2] ,
         \SB1_1_14/Component_Function_0/NAND4_in[1] ,
         \SB1_1_14/Component_Function_0/NAND4_in[0] ,
         \SB1_1_14/Component_Function_1/NAND4_in[2] ,
         \SB1_1_14/Component_Function_1/NAND4_in[1] ,
         \SB1_1_14/Component_Function_5/NAND4_in[2] ,
         \SB1_1_14/Component_Function_5/NAND4_in[0] ,
         \SB1_1_15/Component_Function_0/NAND4_in[3] ,
         \SB1_1_15/Component_Function_0/NAND4_in[1] ,
         \SB1_1_15/Component_Function_0/NAND4_in[0] ,
         \SB1_1_15/Component_Function_1/NAND4_in[3] ,
         \SB1_1_15/Component_Function_1/NAND4_in[2] ,
         \SB1_1_15/Component_Function_1/NAND4_in[1] ,
         \SB1_1_15/Component_Function_1/NAND4_in[0] ,
         \SB1_1_15/Component_Function_5/NAND4_in[1] ,
         \SB1_1_15/Component_Function_5/NAND4_in[0] ,
         \SB1_1_16/Component_Function_0/NAND4_in[3] ,
         \SB1_1_16/Component_Function_0/NAND4_in[2] ,
         \SB1_1_16/Component_Function_0/NAND4_in[1] ,
         \SB1_1_16/Component_Function_0/NAND4_in[0] ,
         \SB1_1_16/Component_Function_1/NAND4_in[2] ,
         \SB1_1_16/Component_Function_1/NAND4_in[1] ,
         \SB1_1_16/Component_Function_1/NAND4_in[0] ,
         \SB1_1_16/Component_Function_5/NAND4_in[2] ,
         \SB1_1_16/Component_Function_5/NAND4_in[0] ,
         \SB1_1_17/Component_Function_0/NAND4_in[3] ,
         \SB1_1_17/Component_Function_0/NAND4_in[2] ,
         \SB1_1_17/Component_Function_0/NAND4_in[1] ,
         \SB1_1_17/Component_Function_0/NAND4_in[0] ,
         \SB1_1_17/Component_Function_1/NAND4_in[3] ,
         \SB1_1_17/Component_Function_1/NAND4_in[1] ,
         \SB1_1_17/Component_Function_1/NAND4_in[0] ,
         \SB1_1_17/Component_Function_5/NAND4_in[3] ,
         \SB1_1_17/Component_Function_5/NAND4_in[1] ,
         \SB1_1_17/Component_Function_5/NAND4_in[0] ,
         \SB1_1_18/Component_Function_0/NAND4_in[3] ,
         \SB1_1_18/Component_Function_0/NAND4_in[2] ,
         \SB1_1_18/Component_Function_0/NAND4_in[1] ,
         \SB1_1_18/Component_Function_0/NAND4_in[0] ,
         \SB1_1_18/Component_Function_1/NAND4_in[3] ,
         \SB1_1_18/Component_Function_1/NAND4_in[2] ,
         \SB1_1_18/Component_Function_1/NAND4_in[1] ,
         \SB1_1_18/Component_Function_1/NAND4_in[0] ,
         \SB1_1_18/Component_Function_5/NAND4_in[1] ,
         \SB1_1_18/Component_Function_5/NAND4_in[0] ,
         \SB1_1_19/Component_Function_0/NAND4_in[3] ,
         \SB1_1_19/Component_Function_0/NAND4_in[2] ,
         \SB1_1_19/Component_Function_0/NAND4_in[1] ,
         \SB1_1_19/Component_Function_0/NAND4_in[0] ,
         \SB1_1_19/Component_Function_1/NAND4_in[3] ,
         \SB1_1_19/Component_Function_1/NAND4_in[2] ,
         \SB1_1_19/Component_Function_1/NAND4_in[1] ,
         \SB1_1_19/Component_Function_1/NAND4_in[0] ,
         \SB1_1_19/Component_Function_5/NAND4_in[1] ,
         \SB1_1_19/Component_Function_5/NAND4_in[0] ,
         \SB1_1_20/Component_Function_0/NAND4_in[3] ,
         \SB1_1_20/Component_Function_0/NAND4_in[2] ,
         \SB1_1_20/Component_Function_0/NAND4_in[1] ,
         \SB1_1_20/Component_Function_0/NAND4_in[0] ,
         \SB1_1_20/Component_Function_1/NAND4_in[2] ,
         \SB1_1_20/Component_Function_1/NAND4_in[1] ,
         \SB1_1_20/Component_Function_1/NAND4_in[0] ,
         \SB1_1_20/Component_Function_5/NAND4_in[2] ,
         \SB1_1_20/Component_Function_5/NAND4_in[1] ,
         \SB1_1_20/Component_Function_5/NAND4_in[0] ,
         \SB1_1_21/Component_Function_0/NAND4_in[3] ,
         \SB1_1_21/Component_Function_0/NAND4_in[2] ,
         \SB1_1_21/Component_Function_0/NAND4_in[1] ,
         \SB1_1_21/Component_Function_0/NAND4_in[0] ,
         \SB1_1_21/Component_Function_1/NAND4_in[2] ,
         \SB1_1_21/Component_Function_1/NAND4_in[1] ,
         \SB1_1_21/Component_Function_1/NAND4_in[0] ,
         \SB1_1_22/Component_Function_0/NAND4_in[2] ,
         \SB1_1_22/Component_Function_0/NAND4_in[1] ,
         \SB1_1_22/Component_Function_0/NAND4_in[0] ,
         \SB1_1_22/Component_Function_1/NAND4_in[3] ,
         \SB1_1_22/Component_Function_1/NAND4_in[2] ,
         \SB1_1_22/Component_Function_1/NAND4_in[1] ,
         \SB1_1_22/Component_Function_1/NAND4_in[0] ,
         \SB1_1_22/Component_Function_5/NAND4_in[2] ,
         \SB1_1_22/Component_Function_5/NAND4_in[0] ,
         \SB1_1_23/Component_Function_0/NAND4_in[3] ,
         \SB1_1_23/Component_Function_0/NAND4_in[2] ,
         \SB1_1_23/Component_Function_0/NAND4_in[1] ,
         \SB1_1_23/Component_Function_0/NAND4_in[0] ,
         \SB1_1_23/Component_Function_1/NAND4_in[2] ,
         \SB1_1_23/Component_Function_1/NAND4_in[1] ,
         \SB1_1_23/Component_Function_1/NAND4_in[0] ,
         \SB1_1_23/Component_Function_5/NAND4_in[2] ,
         \SB1_1_24/Component_Function_0/NAND4_in[2] ,
         \SB1_1_24/Component_Function_0/NAND4_in[1] ,
         \SB1_1_24/Component_Function_0/NAND4_in[0] ,
         \SB1_1_24/Component_Function_1/NAND4_in[2] ,
         \SB1_1_24/Component_Function_1/NAND4_in[1] ,
         \SB1_1_24/Component_Function_1/NAND4_in[0] ,
         \SB1_1_24/Component_Function_5/NAND4_in[0] ,
         \SB1_1_25/Component_Function_0/NAND4_in[2] ,
         \SB1_1_25/Component_Function_0/NAND4_in[1] ,
         \SB1_1_25/Component_Function_0/NAND4_in[0] ,
         \SB1_1_25/Component_Function_1/NAND4_in[3] ,
         \SB1_1_25/Component_Function_1/NAND4_in[2] ,
         \SB1_1_25/Component_Function_1/NAND4_in[1] ,
         \SB1_1_25/Component_Function_1/NAND4_in[0] ,
         \SB1_1_25/Component_Function_5/NAND4_in[2] ,
         \SB1_1_25/Component_Function_5/NAND4_in[1] ,
         \SB1_1_26/Component_Function_0/NAND4_in[3] ,
         \SB1_1_26/Component_Function_0/NAND4_in[2] ,
         \SB1_1_26/Component_Function_0/NAND4_in[1] ,
         \SB1_1_26/Component_Function_0/NAND4_in[0] ,
         \SB1_1_26/Component_Function_1/NAND4_in[2] ,
         \SB1_1_26/Component_Function_1/NAND4_in[1] ,
         \SB1_1_26/Component_Function_1/NAND4_in[0] ,
         \SB1_1_26/Component_Function_5/NAND4_in[2] ,
         \SB1_1_26/Component_Function_5/NAND4_in[1] ,
         \SB1_1_26/Component_Function_5/NAND4_in[0] ,
         \SB1_1_27/Component_Function_0/NAND4_in[3] ,
         \SB1_1_27/Component_Function_0/NAND4_in[1] ,
         \SB1_1_27/Component_Function_0/NAND4_in[0] ,
         \SB1_1_27/Component_Function_1/NAND4_in[2] ,
         \SB1_1_27/Component_Function_1/NAND4_in[1] ,
         \SB1_1_27/Component_Function_1/NAND4_in[0] ,
         \SB1_1_27/Component_Function_5/NAND4_in[1] ,
         \SB1_1_28/Component_Function_0/NAND4_in[2] ,
         \SB1_1_28/Component_Function_0/NAND4_in[0] ,
         \SB1_1_28/Component_Function_1/NAND4_in[3] ,
         \SB1_1_28/Component_Function_1/NAND4_in[2] ,
         \SB1_1_28/Component_Function_1/NAND4_in[1] ,
         \SB1_1_28/Component_Function_1/NAND4_in[0] ,
         \SB1_1_28/Component_Function_5/NAND4_in[1] ,
         \SB1_1_28/Component_Function_5/NAND4_in[0] ,
         \SB1_1_29/Component_Function_0/NAND4_in[2] ,
         \SB1_1_29/Component_Function_0/NAND4_in[1] ,
         \SB1_1_29/Component_Function_0/NAND4_in[0] ,
         \SB1_1_29/Component_Function_1/NAND4_in[3] ,
         \SB1_1_29/Component_Function_1/NAND4_in[2] ,
         \SB1_1_29/Component_Function_1/NAND4_in[1] ,
         \SB1_1_29/Component_Function_1/NAND4_in[0] ,
         \SB1_1_29/Component_Function_5/NAND4_in[2] ,
         \SB1_1_29/Component_Function_5/NAND4_in[1] ,
         \SB1_1_29/Component_Function_5/NAND4_in[0] ,
         \SB1_1_30/Component_Function_0/NAND4_in[3] ,
         \SB1_1_30/Component_Function_0/NAND4_in[2] ,
         \SB1_1_30/Component_Function_0/NAND4_in[1] ,
         \SB1_1_30/Component_Function_0/NAND4_in[0] ,
         \SB1_1_30/Component_Function_1/NAND4_in[2] ,
         \SB1_1_30/Component_Function_1/NAND4_in[1] ,
         \SB1_1_30/Component_Function_1/NAND4_in[0] ,
         \SB1_1_30/Component_Function_5/NAND4_in[2] ,
         \SB1_1_30/Component_Function_5/NAND4_in[1] ,
         \SB1_1_30/Component_Function_5/NAND4_in[0] ,
         \SB1_1_31/Component_Function_0/NAND4_in[3] ,
         \SB1_1_31/Component_Function_0/NAND4_in[2] ,
         \SB1_1_31/Component_Function_0/NAND4_in[1] ,
         \SB1_1_31/Component_Function_0/NAND4_in[0] ,
         \SB1_1_31/Component_Function_1/NAND4_in[2] ,
         \SB1_1_31/Component_Function_1/NAND4_in[1] ,
         \SB1_1_31/Component_Function_1/NAND4_in[0] ,
         \SB1_1_31/Component_Function_5/NAND4_in[3] ,
         \SB1_1_31/Component_Function_5/NAND4_in[2] ,
         \SB1_1_31/Component_Function_5/NAND4_in[1] ,
         \SB1_1_31/Component_Function_5/NAND4_in[0] ,
         \SB2_1_0/Component_Function_0/NAND4_in[3] ,
         \SB2_1_0/Component_Function_0/NAND4_in[2] ,
         \SB2_1_0/Component_Function_0/NAND4_in[0] ,
         \SB2_1_0/Component_Function_1/NAND4_in[2] ,
         \SB2_1_0/Component_Function_1/NAND4_in[1] ,
         \SB2_1_0/Component_Function_1/NAND4_in[0] ,
         \SB2_1_0/Component_Function_5/NAND4_in[2] ,
         \SB2_1_0/Component_Function_5/NAND4_in[1] ,
         \SB2_1_0/Component_Function_5/NAND4_in[0] ,
         \SB2_1_1/Component_Function_0/NAND4_in[3] ,
         \SB2_1_1/Component_Function_0/NAND4_in[2] ,
         \SB2_1_1/Component_Function_0/NAND4_in[1] ,
         \SB2_1_1/Component_Function_0/NAND4_in[0] ,
         \SB2_1_1/Component_Function_1/NAND4_in[3] ,
         \SB2_1_1/Component_Function_1/NAND4_in[2] ,
         \SB2_1_1/Component_Function_5/NAND4_in[0] ,
         \SB2_1_2/Component_Function_0/NAND4_in[2] ,
         \SB2_1_2/Component_Function_0/NAND4_in[1] ,
         \SB2_1_2/Component_Function_0/NAND4_in[0] ,
         \SB2_1_2/Component_Function_1/NAND4_in[2] ,
         \SB2_1_2/Component_Function_1/NAND4_in[1] ,
         \SB2_1_2/Component_Function_1/NAND4_in[0] ,
         \SB2_1_2/Component_Function_5/NAND4_in[2] ,
         \SB2_1_2/Component_Function_5/NAND4_in[0] ,
         \SB2_1_3/Component_Function_0/NAND4_in[3] ,
         \SB2_1_3/Component_Function_0/NAND4_in[2] ,
         \SB2_1_3/Component_Function_0/NAND4_in[1] ,
         \SB2_1_3/Component_Function_1/NAND4_in[2] ,
         \SB2_1_3/Component_Function_1/NAND4_in[1] ,
         \SB2_1_3/Component_Function_1/NAND4_in[0] ,
         \SB2_1_3/Component_Function_5/NAND4_in[0] ,
         \SB2_1_4/Component_Function_0/NAND4_in[2] ,
         \SB2_1_4/Component_Function_0/NAND4_in[1] ,
         \SB2_1_4/Component_Function_0/NAND4_in[0] ,
         \SB2_1_4/Component_Function_1/NAND4_in[3] ,
         \SB2_1_4/Component_Function_1/NAND4_in[2] ,
         \SB2_1_4/Component_Function_1/NAND4_in[1] ,
         \SB2_1_4/Component_Function_1/NAND4_in[0] ,
         \SB2_1_4/Component_Function_5/NAND4_in[3] ,
         \SB2_1_4/Component_Function_5/NAND4_in[2] ,
         \SB2_1_5/Component_Function_0/NAND4_in[1] ,
         \SB2_1_5/Component_Function_0/NAND4_in[0] ,
         \SB2_1_5/Component_Function_1/NAND4_in[3] ,
         \SB2_1_5/Component_Function_1/NAND4_in[1] ,
         \SB2_1_5/Component_Function_1/NAND4_in[0] ,
         \SB2_1_5/Component_Function_5/NAND4_in[2] ,
         \SB2_1_5/Component_Function_5/NAND4_in[0] ,
         \SB2_1_6/Component_Function_0/NAND4_in[3] ,
         \SB2_1_6/Component_Function_0/NAND4_in[1] ,
         \SB2_1_6/Component_Function_0/NAND4_in[0] ,
         \SB2_1_6/Component_Function_1/NAND4_in[3] ,
         \SB2_1_6/Component_Function_1/NAND4_in[2] ,
         \SB2_1_6/Component_Function_1/NAND4_in[1] ,
         \SB2_1_6/Component_Function_1/NAND4_in[0] ,
         \SB2_1_6/Component_Function_5/NAND4_in[3] ,
         \SB2_1_6/Component_Function_5/NAND4_in[1] ,
         \SB2_1_6/Component_Function_5/NAND4_in[0] ,
         \SB2_1_7/Component_Function_0/NAND4_in[3] ,
         \SB2_1_7/Component_Function_0/NAND4_in[2] ,
         \SB2_1_7/Component_Function_0/NAND4_in[1] ,
         \SB2_1_7/Component_Function_0/NAND4_in[0] ,
         \SB2_1_7/Component_Function_1/NAND4_in[3] ,
         \SB2_1_7/Component_Function_1/NAND4_in[2] ,
         \SB2_1_7/Component_Function_1/NAND4_in[1] ,
         \SB2_1_7/Component_Function_1/NAND4_in[0] ,
         \SB2_1_7/Component_Function_5/NAND4_in[2] ,
         \SB2_1_7/Component_Function_5/NAND4_in[1] ,
         \SB2_1_7/Component_Function_5/NAND4_in[0] ,
         \SB2_1_8/Component_Function_0/NAND4_in[3] ,
         \SB2_1_8/Component_Function_0/NAND4_in[2] ,
         \SB2_1_8/Component_Function_0/NAND4_in[0] ,
         \SB2_1_8/Component_Function_1/NAND4_in[2] ,
         \SB2_1_8/Component_Function_1/NAND4_in[1] ,
         \SB2_1_8/Component_Function_1/NAND4_in[0] ,
         \SB2_1_8/Component_Function_5/NAND4_in[3] ,
         \SB2_1_8/Component_Function_5/NAND4_in[1] ,
         \SB2_1_8/Component_Function_5/NAND4_in[0] ,
         \SB2_1_9/Component_Function_0/NAND4_in[1] ,
         \SB2_1_9/Component_Function_0/NAND4_in[0] ,
         \SB2_1_9/Component_Function_1/NAND4_in[3] ,
         \SB2_1_9/Component_Function_1/NAND4_in[2] ,
         \SB2_1_9/Component_Function_1/NAND4_in[0] ,
         \SB2_1_9/Component_Function_5/NAND4_in[1] ,
         \SB2_1_9/Component_Function_5/NAND4_in[0] ,
         \SB2_1_10/Component_Function_0/NAND4_in[3] ,
         \SB2_1_10/Component_Function_0/NAND4_in[1] ,
         \SB2_1_10/Component_Function_0/NAND4_in[0] ,
         \SB2_1_10/Component_Function_1/NAND4_in[3] ,
         \SB2_1_10/Component_Function_1/NAND4_in[2] ,
         \SB2_1_10/Component_Function_1/NAND4_in[0] ,
         \SB2_1_10/Component_Function_5/NAND4_in[1] ,
         \SB2_1_10/Component_Function_5/NAND4_in[0] ,
         \SB2_1_11/Component_Function_0/NAND4_in[2] ,
         \SB2_1_11/Component_Function_0/NAND4_in[1] ,
         \SB2_1_11/Component_Function_0/NAND4_in[0] ,
         \SB2_1_11/Component_Function_1/NAND4_in[3] ,
         \SB2_1_11/Component_Function_1/NAND4_in[1] ,
         \SB2_1_11/Component_Function_1/NAND4_in[0] ,
         \SB2_1_11/Component_Function_5/NAND4_in[2] ,
         \SB2_1_11/Component_Function_5/NAND4_in[1] ,
         \SB2_1_11/Component_Function_5/NAND4_in[0] ,
         \SB2_1_12/Component_Function_0/NAND4_in[3] ,
         \SB2_1_12/Component_Function_0/NAND4_in[1] ,
         \SB2_1_12/Component_Function_0/NAND4_in[0] ,
         \SB2_1_12/Component_Function_1/NAND4_in[3] ,
         \SB2_1_12/Component_Function_1/NAND4_in[2] ,
         \SB2_1_12/Component_Function_1/NAND4_in[1] ,
         \SB2_1_12/Component_Function_1/NAND4_in[0] ,
         \SB2_1_12/Component_Function_5/NAND4_in[2] ,
         \SB2_1_13/Component_Function_0/NAND4_in[3] ,
         \SB2_1_13/Component_Function_0/NAND4_in[2] ,
         \SB2_1_13/Component_Function_0/NAND4_in[0] ,
         \SB2_1_13/Component_Function_1/NAND4_in[3] ,
         \SB2_1_13/Component_Function_1/NAND4_in[2] ,
         \SB2_1_13/Component_Function_1/NAND4_in[0] ,
         \SB2_1_13/Component_Function_5/NAND4_in[0] ,
         \SB2_1_14/Component_Function_0/NAND4_in[3] ,
         \SB2_1_14/Component_Function_0/NAND4_in[1] ,
         \SB2_1_14/Component_Function_0/NAND4_in[0] ,
         \SB2_1_14/Component_Function_1/NAND4_in[3] ,
         \SB2_1_14/Component_Function_1/NAND4_in[2] ,
         \SB2_1_14/Component_Function_1/NAND4_in[1] ,
         \SB2_1_14/Component_Function_1/NAND4_in[0] ,
         \SB2_1_14/Component_Function_5/NAND4_in[2] ,
         \SB2_1_14/Component_Function_5/NAND4_in[1] ,
         \SB2_1_15/Component_Function_0/NAND4_in[2] ,
         \SB2_1_15/Component_Function_0/NAND4_in[1] ,
         \SB2_1_15/Component_Function_0/NAND4_in[0] ,
         \SB2_1_15/Component_Function_1/NAND4_in[2] ,
         \SB2_1_15/Component_Function_1/NAND4_in[1] ,
         \SB2_1_15/Component_Function_1/NAND4_in[0] ,
         \SB2_1_15/Component_Function_5/NAND4_in[3] ,
         \SB2_1_15/Component_Function_5/NAND4_in[2] ,
         \SB2_1_15/Component_Function_5/NAND4_in[0] ,
         \SB2_1_16/Component_Function_0/NAND4_in[3] ,
         \SB2_1_16/Component_Function_0/NAND4_in[1] ,
         \SB2_1_16/Component_Function_1/NAND4_in[2] ,
         \SB2_1_16/Component_Function_1/NAND4_in[1] ,
         \SB2_1_16/Component_Function_1/NAND4_in[0] ,
         \SB2_1_16/Component_Function_5/NAND4_in[0] ,
         \SB2_1_17/Component_Function_0/NAND4_in[3] ,
         \SB2_1_17/Component_Function_0/NAND4_in[1] ,
         \SB2_1_17/Component_Function_0/NAND4_in[0] ,
         \SB2_1_17/Component_Function_1/NAND4_in[3] ,
         \SB2_1_17/Component_Function_1/NAND4_in[2] ,
         \SB2_1_17/Component_Function_1/NAND4_in[1] ,
         \SB2_1_17/Component_Function_1/NAND4_in[0] ,
         \SB2_1_17/Component_Function_5/NAND4_in[2] ,
         \SB2_1_17/Component_Function_5/NAND4_in[0] ,
         \SB2_1_18/Component_Function_0/NAND4_in[1] ,
         \SB2_1_18/Component_Function_0/NAND4_in[0] ,
         \SB2_1_18/Component_Function_1/NAND4_in[3] ,
         \SB2_1_18/Component_Function_1/NAND4_in[2] ,
         \SB2_1_18/Component_Function_1/NAND4_in[1] ,
         \SB2_1_18/Component_Function_1/NAND4_in[0] ,
         \SB2_1_19/Component_Function_0/NAND4_in[2] ,
         \SB2_1_19/Component_Function_0/NAND4_in[1] ,
         \SB2_1_19/Component_Function_1/NAND4_in[2] ,
         \SB2_1_19/Component_Function_1/NAND4_in[1] ,
         \SB2_1_19/Component_Function_1/NAND4_in[0] ,
         \SB2_1_19/Component_Function_5/NAND4_in[3] ,
         \SB2_1_19/Component_Function_5/NAND4_in[0] ,
         \SB2_1_20/Component_Function_0/NAND4_in[1] ,
         \SB2_1_20/Component_Function_0/NAND4_in[0] ,
         \SB2_1_20/Component_Function_1/NAND4_in[2] ,
         \SB2_1_20/Component_Function_1/NAND4_in[1] ,
         \SB2_1_20/Component_Function_1/NAND4_in[0] ,
         \SB2_1_20/Component_Function_5/NAND4_in[1] ,
         \SB2_1_20/Component_Function_5/NAND4_in[0] ,
         \SB2_1_21/Component_Function_0/NAND4_in[2] ,
         \SB2_1_21/Component_Function_0/NAND4_in[1] ,
         \SB2_1_21/Component_Function_0/NAND4_in[0] ,
         \SB2_1_21/Component_Function_1/NAND4_in[3] ,
         \SB2_1_21/Component_Function_1/NAND4_in[2] ,
         \SB2_1_21/Component_Function_1/NAND4_in[1] ,
         \SB2_1_21/Component_Function_1/NAND4_in[0] ,
         \SB2_1_21/Component_Function_5/NAND4_in[3] ,
         \SB2_1_21/Component_Function_5/NAND4_in[0] ,
         \SB2_1_22/Component_Function_0/NAND4_in[2] ,
         \SB2_1_22/Component_Function_0/NAND4_in[1] ,
         \SB2_1_22/Component_Function_0/NAND4_in[0] ,
         \SB2_1_22/Component_Function_1/NAND4_in[3] ,
         \SB2_1_22/Component_Function_1/NAND4_in[1] ,
         \SB2_1_22/Component_Function_1/NAND4_in[0] ,
         \SB2_1_22/Component_Function_5/NAND4_in[3] ,
         \SB2_1_22/Component_Function_5/NAND4_in[2] ,
         \SB2_1_22/Component_Function_5/NAND4_in[1] ,
         \SB2_1_22/Component_Function_5/NAND4_in[0] ,
         \SB2_1_23/Component_Function_0/NAND4_in[3] ,
         \SB2_1_23/Component_Function_0/NAND4_in[1] ,
         \SB2_1_23/Component_Function_0/NAND4_in[0] ,
         \SB2_1_23/Component_Function_1/NAND4_in[3] ,
         \SB2_1_23/Component_Function_1/NAND4_in[2] ,
         \SB2_1_23/Component_Function_1/NAND4_in[1] ,
         \SB2_1_23/Component_Function_1/NAND4_in[0] ,
         \SB2_1_23/Component_Function_5/NAND4_in[1] ,
         \SB2_1_23/Component_Function_5/NAND4_in[0] ,
         \SB2_1_24/Component_Function_0/NAND4_in[3] ,
         \SB2_1_24/Component_Function_0/NAND4_in[1] ,
         \SB2_1_24/Component_Function_1/NAND4_in[2] ,
         \SB2_1_24/Component_Function_1/NAND4_in[1] ,
         \SB2_1_24/Component_Function_1/NAND4_in[0] ,
         \SB2_1_24/Component_Function_5/NAND4_in[3] ,
         \SB2_1_24/Component_Function_5/NAND4_in[1] ,
         \SB2_1_24/Component_Function_5/NAND4_in[0] ,
         \SB2_1_25/Component_Function_0/NAND4_in[3] ,
         \SB2_1_25/Component_Function_0/NAND4_in[1] ,
         \SB2_1_25/Component_Function_0/NAND4_in[0] ,
         \SB2_1_25/Component_Function_1/NAND4_in[3] ,
         \SB2_1_25/Component_Function_1/NAND4_in[2] ,
         \SB2_1_25/Component_Function_1/NAND4_in[1] ,
         \SB2_1_25/Component_Function_1/NAND4_in[0] ,
         \SB2_1_25/Component_Function_5/NAND4_in[3] ,
         \SB2_1_25/Component_Function_5/NAND4_in[0] ,
         \SB2_1_26/Component_Function_0/NAND4_in[1] ,
         \SB2_1_26/Component_Function_1/NAND4_in[2] ,
         \SB2_1_26/Component_Function_1/NAND4_in[1] ,
         \SB2_1_26/Component_Function_1/NAND4_in[0] ,
         \SB2_1_26/Component_Function_5/NAND4_in[2] ,
         \SB2_1_26/Component_Function_5/NAND4_in[1] ,
         \SB2_1_26/Component_Function_5/NAND4_in[0] ,
         \SB2_1_27/Component_Function_0/NAND4_in[2] ,
         \SB2_1_27/Component_Function_0/NAND4_in[1] ,
         \SB2_1_27/Component_Function_0/NAND4_in[0] ,
         \SB2_1_27/Component_Function_1/NAND4_in[3] ,
         \SB2_1_27/Component_Function_1/NAND4_in[1] ,
         \SB2_1_27/Component_Function_1/NAND4_in[0] ,
         \SB2_1_27/Component_Function_5/NAND4_in[2] ,
         \SB2_1_27/Component_Function_5/NAND4_in[1] ,
         \SB2_1_27/Component_Function_5/NAND4_in[0] ,
         \SB2_1_28/Component_Function_0/NAND4_in[2] ,
         \SB2_1_28/Component_Function_0/NAND4_in[1] ,
         \SB2_1_28/Component_Function_0/NAND4_in[0] ,
         \SB2_1_28/Component_Function_1/NAND4_in[2] ,
         \SB2_1_28/Component_Function_1/NAND4_in[1] ,
         \SB2_1_28/Component_Function_1/NAND4_in[0] ,
         \SB2_1_28/Component_Function_5/NAND4_in[2] ,
         \SB2_1_28/Component_Function_5/NAND4_in[1] ,
         \SB2_1_28/Component_Function_5/NAND4_in[0] ,
         \SB2_1_29/Component_Function_0/NAND4_in[3] ,
         \SB2_1_29/Component_Function_0/NAND4_in[2] ,
         \SB2_1_29/Component_Function_0/NAND4_in[1] ,
         \SB2_1_29/Component_Function_0/NAND4_in[0] ,
         \SB2_1_29/Component_Function_1/NAND4_in[3] ,
         \SB2_1_29/Component_Function_1/NAND4_in[2] ,
         \SB2_1_29/Component_Function_1/NAND4_in[1] ,
         \SB2_1_29/Component_Function_1/NAND4_in[0] ,
         \SB2_1_29/Component_Function_5/NAND4_in[2] ,
         \SB2_1_29/Component_Function_5/NAND4_in[0] ,
         \SB2_1_30/Component_Function_0/NAND4_in[2] ,
         \SB2_1_30/Component_Function_0/NAND4_in[1] ,
         \SB2_1_30/Component_Function_0/NAND4_in[0] ,
         \SB2_1_30/Component_Function_1/NAND4_in[3] ,
         \SB2_1_30/Component_Function_1/NAND4_in[1] ,
         \SB2_1_30/Component_Function_1/NAND4_in[0] ,
         \SB2_1_30/Component_Function_5/NAND4_in[0] ,
         \SB2_1_31/Component_Function_0/NAND4_in[3] ,
         \SB2_1_31/Component_Function_0/NAND4_in[2] ,
         \SB2_1_31/Component_Function_0/NAND4_in[1] ,
         \SB2_1_31/Component_Function_0/NAND4_in[0] ,
         \SB2_1_31/Component_Function_1/NAND4_in[3] ,
         \SB2_1_31/Component_Function_1/NAND4_in[2] ,
         \SB2_1_31/Component_Function_1/NAND4_in[1] ,
         \SB2_1_31/Component_Function_1/NAND4_in[0] ,
         \SB2_1_31/Component_Function_5/NAND4_in[0] ,
         \SB1_2_0/Component_Function_0/NAND4_in[3] ,
         \SB1_2_0/Component_Function_0/NAND4_in[2] ,
         \SB1_2_0/Component_Function_0/NAND4_in[1] ,
         \SB1_2_0/Component_Function_0/NAND4_in[0] ,
         \SB1_2_0/Component_Function_1/NAND4_in[3] ,
         \SB1_2_0/Component_Function_1/NAND4_in[2] ,
         \SB1_2_0/Component_Function_1/NAND4_in[1] ,
         \SB1_2_0/Component_Function_1/NAND4_in[0] ,
         \SB1_2_0/Component_Function_5/NAND4_in[2] ,
         \SB1_2_0/Component_Function_5/NAND4_in[1] ,
         \SB1_2_0/Component_Function_5/NAND4_in[0] ,
         \SB1_2_1/Component_Function_0/NAND4_in[2] ,
         \SB1_2_1/Component_Function_0/NAND4_in[1] ,
         \SB1_2_1/Component_Function_0/NAND4_in[0] ,
         \SB1_2_1/Component_Function_1/NAND4_in[2] ,
         \SB1_2_1/Component_Function_1/NAND4_in[1] ,
         \SB1_2_1/Component_Function_1/NAND4_in[0] ,
         \SB1_2_1/Component_Function_5/NAND4_in[1] ,
         \SB1_2_1/Component_Function_5/NAND4_in[0] ,
         \SB1_2_2/Component_Function_0/NAND4_in[2] ,
         \SB1_2_2/Component_Function_0/NAND4_in[1] ,
         \SB1_2_2/Component_Function_0/NAND4_in[0] ,
         \SB1_2_2/Component_Function_1/NAND4_in[3] ,
         \SB1_2_2/Component_Function_1/NAND4_in[2] ,
         \SB1_2_2/Component_Function_1/NAND4_in[1] ,
         \SB1_2_2/Component_Function_1/NAND4_in[0] ,
         \SB1_2_2/Component_Function_5/NAND4_in[3] ,
         \SB1_2_2/Component_Function_5/NAND4_in[2] ,
         \SB1_2_2/Component_Function_5/NAND4_in[1] ,
         \SB1_2_2/Component_Function_5/NAND4_in[0] ,
         \SB1_2_3/Component_Function_0/NAND4_in[3] ,
         \SB1_2_3/Component_Function_0/NAND4_in[1] ,
         \SB1_2_3/Component_Function_0/NAND4_in[0] ,
         \SB1_2_3/Component_Function_1/NAND4_in[3] ,
         \SB1_2_3/Component_Function_1/NAND4_in[2] ,
         \SB1_2_3/Component_Function_1/NAND4_in[1] ,
         \SB1_2_3/Component_Function_1/NAND4_in[0] ,
         \SB1_2_3/Component_Function_5/NAND4_in[2] ,
         \SB1_2_3/Component_Function_5/NAND4_in[0] ,
         \SB1_2_4/Component_Function_0/NAND4_in[2] ,
         \SB1_2_4/Component_Function_0/NAND4_in[1] ,
         \SB1_2_4/Component_Function_0/NAND4_in[0] ,
         \SB1_2_4/Component_Function_1/NAND4_in[3] ,
         \SB1_2_4/Component_Function_1/NAND4_in[2] ,
         \SB1_2_4/Component_Function_1/NAND4_in[1] ,
         \SB1_2_4/Component_Function_1/NAND4_in[0] ,
         \SB1_2_4/Component_Function_5/NAND4_in[2] ,
         \SB1_2_4/Component_Function_5/NAND4_in[0] ,
         \SB1_2_5/Component_Function_0/NAND4_in[2] ,
         \SB1_2_5/Component_Function_0/NAND4_in[1] ,
         \SB1_2_5/Component_Function_0/NAND4_in[0] ,
         \SB1_2_5/Component_Function_1/NAND4_in[3] ,
         \SB1_2_5/Component_Function_1/NAND4_in[1] ,
         \SB1_2_5/Component_Function_1/NAND4_in[0] ,
         \SB1_2_5/Component_Function_5/NAND4_in[2] ,
         \SB1_2_5/Component_Function_5/NAND4_in[1] ,
         \SB1_2_6/Component_Function_0/NAND4_in[2] ,
         \SB1_2_6/Component_Function_0/NAND4_in[1] ,
         \SB1_2_6/Component_Function_0/NAND4_in[0] ,
         \SB1_2_6/Component_Function_1/NAND4_in[2] ,
         \SB1_2_6/Component_Function_1/NAND4_in[1] ,
         \SB1_2_6/Component_Function_1/NAND4_in[0] ,
         \SB1_2_6/Component_Function_5/NAND4_in[3] ,
         \SB1_2_6/Component_Function_5/NAND4_in[0] ,
         \SB1_2_7/Component_Function_0/NAND4_in[1] ,
         \SB1_2_7/Component_Function_0/NAND4_in[0] ,
         \SB1_2_7/Component_Function_1/NAND4_in[3] ,
         \SB1_2_7/Component_Function_1/NAND4_in[1] ,
         \SB1_2_7/Component_Function_1/NAND4_in[0] ,
         \SB1_2_7/Component_Function_5/NAND4_in[1] ,
         \SB1_2_7/Component_Function_5/NAND4_in[0] ,
         \SB1_2_8/Component_Function_0/NAND4_in[3] ,
         \SB1_2_8/Component_Function_0/NAND4_in[1] ,
         \SB1_2_8/Component_Function_0/NAND4_in[0] ,
         \SB1_2_8/Component_Function_1/NAND4_in[3] ,
         \SB1_2_8/Component_Function_1/NAND4_in[2] ,
         \SB1_2_8/Component_Function_1/NAND4_in[1] ,
         \SB1_2_8/Component_Function_1/NAND4_in[0] ,
         \SB1_2_8/Component_Function_5/NAND4_in[2] ,
         \SB1_2_8/Component_Function_5/NAND4_in[1] ,
         \SB1_2_8/Component_Function_5/NAND4_in[0] ,
         \SB1_2_9/Component_Function_0/NAND4_in[3] ,
         \SB1_2_9/Component_Function_0/NAND4_in[2] ,
         \SB1_2_9/Component_Function_0/NAND4_in[1] ,
         \SB1_2_9/Component_Function_0/NAND4_in[0] ,
         \SB1_2_9/Component_Function_1/NAND4_in[1] ,
         \SB1_2_9/Component_Function_1/NAND4_in[0] ,
         \SB1_2_9/Component_Function_5/NAND4_in[2] ,
         \SB1_2_10/Component_Function_0/NAND4_in[2] ,
         \SB1_2_10/Component_Function_0/NAND4_in[1] ,
         \SB1_2_10/Component_Function_0/NAND4_in[0] ,
         \SB1_2_10/Component_Function_1/NAND4_in[0] ,
         \SB1_2_10/Component_Function_5/NAND4_in[3] ,
         \SB1_2_10/Component_Function_5/NAND4_in[2] ,
         \SB1_2_10/Component_Function_5/NAND4_in[1] ,
         \SB1_2_10/Component_Function_5/NAND4_in[0] ,
         \SB1_2_11/Component_Function_0/NAND4_in[2] ,
         \SB1_2_11/Component_Function_0/NAND4_in[1] ,
         \SB1_2_11/Component_Function_0/NAND4_in[0] ,
         \SB1_2_11/Component_Function_1/NAND4_in[2] ,
         \SB1_2_11/Component_Function_1/NAND4_in[1] ,
         \SB1_2_11/Component_Function_1/NAND4_in[0] ,
         \SB1_2_11/Component_Function_5/NAND4_in[1] ,
         \SB1_2_11/Component_Function_5/NAND4_in[0] ,
         \SB1_2_12/Component_Function_0/NAND4_in[3] ,
         \SB1_2_12/Component_Function_0/NAND4_in[2] ,
         \SB1_2_12/Component_Function_0/NAND4_in[1] ,
         \SB1_2_12/Component_Function_0/NAND4_in[0] ,
         \SB1_2_12/Component_Function_1/NAND4_in[3] ,
         \SB1_2_12/Component_Function_1/NAND4_in[1] ,
         \SB1_2_12/Component_Function_5/NAND4_in[3] ,
         \SB1_2_12/Component_Function_5/NAND4_in[2] ,
         \SB1_2_12/Component_Function_5/NAND4_in[1] ,
         \SB1_2_12/Component_Function_5/NAND4_in[0] ,
         \SB1_2_13/Component_Function_0/NAND4_in[3] ,
         \SB1_2_13/Component_Function_0/NAND4_in[2] ,
         \SB1_2_13/Component_Function_0/NAND4_in[1] ,
         \SB1_2_13/Component_Function_0/NAND4_in[0] ,
         \SB1_2_13/Component_Function_1/NAND4_in[3] ,
         \SB1_2_13/Component_Function_1/NAND4_in[2] ,
         \SB1_2_13/Component_Function_1/NAND4_in[1] ,
         \SB1_2_13/Component_Function_1/NAND4_in[0] ,
         \SB1_2_13/Component_Function_5/NAND4_in[2] ,
         \SB1_2_13/Component_Function_5/NAND4_in[1] ,
         \SB1_2_13/Component_Function_5/NAND4_in[0] ,
         \SB1_2_14/Component_Function_0/NAND4_in[3] ,
         \SB1_2_14/Component_Function_0/NAND4_in[2] ,
         \SB1_2_14/Component_Function_0/NAND4_in[1] ,
         \SB1_2_14/Component_Function_0/NAND4_in[0] ,
         \SB1_2_14/Component_Function_1/NAND4_in[2] ,
         \SB1_2_14/Component_Function_1/NAND4_in[1] ,
         \SB1_2_14/Component_Function_5/NAND4_in[1] ,
         \SB1_2_14/Component_Function_5/NAND4_in[0] ,
         \SB1_2_15/Component_Function_0/NAND4_in[2] ,
         \SB1_2_15/Component_Function_0/NAND4_in[1] ,
         \SB1_2_15/Component_Function_0/NAND4_in[0] ,
         \SB1_2_15/Component_Function_1/NAND4_in[3] ,
         \SB1_2_15/Component_Function_1/NAND4_in[2] ,
         \SB1_2_15/Component_Function_1/NAND4_in[1] ,
         \SB1_2_15/Component_Function_5/NAND4_in[3] ,
         \SB1_2_15/Component_Function_5/NAND4_in[0] ,
         \SB1_2_16/Component_Function_0/NAND4_in[2] ,
         \SB1_2_16/Component_Function_0/NAND4_in[1] ,
         \SB1_2_16/Component_Function_0/NAND4_in[0] ,
         \SB1_2_16/Component_Function_1/NAND4_in[2] ,
         \SB1_2_16/Component_Function_1/NAND4_in[1] ,
         \SB1_2_16/Component_Function_1/NAND4_in[0] ,
         \SB1_2_16/Component_Function_5/NAND4_in[2] ,
         \SB1_2_16/Component_Function_5/NAND4_in[1] ,
         \SB1_2_16/Component_Function_5/NAND4_in[0] ,
         \SB1_2_17/Component_Function_0/NAND4_in[3] ,
         \SB1_2_17/Component_Function_0/NAND4_in[0] ,
         \SB1_2_17/Component_Function_1/NAND4_in[2] ,
         \SB1_2_17/Component_Function_1/NAND4_in[1] ,
         \SB1_2_17/Component_Function_1/NAND4_in[0] ,
         \SB1_2_17/Component_Function_5/NAND4_in[3] ,
         \SB1_2_17/Component_Function_5/NAND4_in[0] ,
         \SB1_2_18/Component_Function_0/NAND4_in[2] ,
         \SB1_2_18/Component_Function_0/NAND4_in[1] ,
         \SB1_2_18/Component_Function_0/NAND4_in[0] ,
         \SB1_2_18/Component_Function_1/NAND4_in[3] ,
         \SB1_2_18/Component_Function_1/NAND4_in[2] ,
         \SB1_2_18/Component_Function_1/NAND4_in[1] ,
         \SB1_2_18/Component_Function_1/NAND4_in[0] ,
         \SB1_2_18/Component_Function_5/NAND4_in[2] ,
         \SB1_2_18/Component_Function_5/NAND4_in[1] ,
         \SB1_2_18/Component_Function_5/NAND4_in[0] ,
         \SB1_2_19/Component_Function_0/NAND4_in[3] ,
         \SB1_2_19/Component_Function_0/NAND4_in[2] ,
         \SB1_2_19/Component_Function_0/NAND4_in[1] ,
         \SB1_2_19/Component_Function_0/NAND4_in[0] ,
         \SB1_2_19/Component_Function_1/NAND4_in[3] ,
         \SB1_2_19/Component_Function_1/NAND4_in[2] ,
         \SB1_2_19/Component_Function_1/NAND4_in[0] ,
         \SB1_2_19/Component_Function_5/NAND4_in[2] ,
         \SB1_2_19/Component_Function_5/NAND4_in[1] ,
         \SB1_2_19/Component_Function_5/NAND4_in[0] ,
         \SB1_2_20/Component_Function_0/NAND4_in[3] ,
         \SB1_2_20/Component_Function_0/NAND4_in[2] ,
         \SB1_2_20/Component_Function_0/NAND4_in[1] ,
         \SB1_2_20/Component_Function_0/NAND4_in[0] ,
         \SB1_2_20/Component_Function_1/NAND4_in[3] ,
         \SB1_2_20/Component_Function_1/NAND4_in[2] ,
         \SB1_2_20/Component_Function_1/NAND4_in[1] ,
         \SB1_2_20/Component_Function_1/NAND4_in[0] ,
         \SB1_2_20/Component_Function_5/NAND4_in[2] ,
         \SB1_2_20/Component_Function_5/NAND4_in[1] ,
         \SB1_2_20/Component_Function_5/NAND4_in[0] ,
         \SB1_2_21/Component_Function_0/NAND4_in[3] ,
         \SB1_2_21/Component_Function_0/NAND4_in[2] ,
         \SB1_2_21/Component_Function_0/NAND4_in[1] ,
         \SB1_2_21/Component_Function_0/NAND4_in[0] ,
         \SB1_2_21/Component_Function_1/NAND4_in[3] ,
         \SB1_2_21/Component_Function_1/NAND4_in[2] ,
         \SB1_2_21/Component_Function_1/NAND4_in[1] ,
         \SB1_2_21/Component_Function_1/NAND4_in[0] ,
         \SB1_2_21/Component_Function_5/NAND4_in[0] ,
         \SB1_2_22/Component_Function_0/NAND4_in[2] ,
         \SB1_2_22/Component_Function_0/NAND4_in[1] ,
         \SB1_2_22/Component_Function_1/NAND4_in[1] ,
         \SB1_2_22/Component_Function_1/NAND4_in[0] ,
         \SB1_2_22/Component_Function_5/NAND4_in[3] ,
         \SB1_2_22/Component_Function_5/NAND4_in[2] ,
         \SB1_2_22/Component_Function_5/NAND4_in[1] ,
         \SB1_2_22/Component_Function_5/NAND4_in[0] ,
         \SB1_2_23/Component_Function_0/NAND4_in[2] ,
         \SB1_2_23/Component_Function_0/NAND4_in[1] ,
         \SB1_2_23/Component_Function_0/NAND4_in[0] ,
         \SB1_2_23/Component_Function_1/NAND4_in[2] ,
         \SB1_2_23/Component_Function_1/NAND4_in[1] ,
         \SB1_2_23/Component_Function_1/NAND4_in[0] ,
         \SB1_2_23/Component_Function_5/NAND4_in[3] ,
         \SB1_2_23/Component_Function_5/NAND4_in[0] ,
         \SB1_2_24/Component_Function_0/NAND4_in[3] ,
         \SB1_2_24/Component_Function_0/NAND4_in[2] ,
         \SB1_2_24/Component_Function_0/NAND4_in[1] ,
         \SB1_2_24/Component_Function_1/NAND4_in[3] ,
         \SB1_2_24/Component_Function_1/NAND4_in[2] ,
         \SB1_2_24/Component_Function_1/NAND4_in[1] ,
         \SB1_2_24/Component_Function_1/NAND4_in[0] ,
         \SB1_2_24/Component_Function_5/NAND4_in[0] ,
         \SB1_2_25/Component_Function_0/NAND4_in[3] ,
         \SB1_2_25/Component_Function_0/NAND4_in[2] ,
         \SB1_2_25/Component_Function_0/NAND4_in[1] ,
         \SB1_2_25/Component_Function_0/NAND4_in[0] ,
         \SB1_2_25/Component_Function_1/NAND4_in[3] ,
         \SB1_2_25/Component_Function_1/NAND4_in[2] ,
         \SB1_2_25/Component_Function_1/NAND4_in[1] ,
         \SB1_2_25/Component_Function_1/NAND4_in[0] ,
         \SB1_2_25/Component_Function_5/NAND4_in[2] ,
         \SB1_2_25/Component_Function_5/NAND4_in[1] ,
         \SB1_2_25/Component_Function_5/NAND4_in[0] ,
         \SB1_2_26/Component_Function_0/NAND4_in[2] ,
         \SB1_2_26/Component_Function_0/NAND4_in[1] ,
         \SB1_2_26/Component_Function_0/NAND4_in[0] ,
         \SB1_2_26/Component_Function_1/NAND4_in[3] ,
         \SB1_2_26/Component_Function_1/NAND4_in[1] ,
         \SB1_2_26/Component_Function_1/NAND4_in[0] ,
         \SB1_2_26/Component_Function_5/NAND4_in[2] ,
         \SB1_2_26/Component_Function_5/NAND4_in[0] ,
         \SB1_2_27/Component_Function_0/NAND4_in[2] ,
         \SB1_2_27/Component_Function_0/NAND4_in[1] ,
         \SB1_2_27/Component_Function_1/NAND4_in[3] ,
         \SB1_2_27/Component_Function_1/NAND4_in[1] ,
         \SB1_2_27/Component_Function_1/NAND4_in[0] ,
         \SB1_2_27/Component_Function_5/NAND4_in[0] ,
         \SB1_2_28/Component_Function_0/NAND4_in[3] ,
         \SB1_2_28/Component_Function_0/NAND4_in[2] ,
         \SB1_2_28/Component_Function_0/NAND4_in[1] ,
         \SB1_2_28/Component_Function_0/NAND4_in[0] ,
         \SB1_2_28/Component_Function_1/NAND4_in[2] ,
         \SB1_2_28/Component_Function_1/NAND4_in[1] ,
         \SB1_2_28/Component_Function_1/NAND4_in[0] ,
         \SB1_2_28/Component_Function_5/NAND4_in[1] ,
         \SB1_2_28/Component_Function_5/NAND4_in[0] ,
         \SB1_2_29/Component_Function_0/NAND4_in[2] ,
         \SB1_2_29/Component_Function_0/NAND4_in[1] ,
         \SB1_2_29/Component_Function_0/NAND4_in[0] ,
         \SB1_2_29/Component_Function_1/NAND4_in[2] ,
         \SB1_2_29/Component_Function_1/NAND4_in[1] ,
         \SB1_2_29/Component_Function_1/NAND4_in[0] ,
         \SB1_2_29/Component_Function_5/NAND4_in[1] ,
         \SB1_2_29/Component_Function_5/NAND4_in[0] ,
         \SB1_2_30/Component_Function_0/NAND4_in[2] ,
         \SB1_2_30/Component_Function_0/NAND4_in[1] ,
         \SB1_2_30/Component_Function_0/NAND4_in[0] ,
         \SB1_2_30/Component_Function_1/NAND4_in[3] ,
         \SB1_2_30/Component_Function_1/NAND4_in[2] ,
         \SB1_2_30/Component_Function_1/NAND4_in[1] ,
         \SB1_2_30/Component_Function_1/NAND4_in[0] ,
         \SB1_2_30/Component_Function_5/NAND4_in[2] ,
         \SB1_2_30/Component_Function_5/NAND4_in[1] ,
         \SB1_2_30/Component_Function_5/NAND4_in[0] ,
         \SB1_2_31/Component_Function_0/NAND4_in[1] ,
         \SB1_2_31/Component_Function_0/NAND4_in[0] ,
         \SB1_2_31/Component_Function_1/NAND4_in[3] ,
         \SB1_2_31/Component_Function_1/NAND4_in[2] ,
         \SB1_2_31/Component_Function_1/NAND4_in[1] ,
         \SB1_2_31/Component_Function_1/NAND4_in[0] ,
         \SB1_2_31/Component_Function_5/NAND4_in[3] ,
         \SB1_2_31/Component_Function_5/NAND4_in[1] ,
         \SB1_2_31/Component_Function_5/NAND4_in[0] ,
         \SB2_2_0/Component_Function_0/NAND4_in[3] ,
         \SB2_2_0/Component_Function_0/NAND4_in[0] ,
         \SB2_2_0/Component_Function_1/NAND4_in[3] ,
         \SB2_2_0/Component_Function_1/NAND4_in[2] ,
         \SB2_2_0/Component_Function_1/NAND4_in[0] ,
         \SB2_2_0/Component_Function_5/NAND4_in[2] ,
         \SB2_2_1/Component_Function_0/NAND4_in[3] ,
         \SB2_2_1/Component_Function_0/NAND4_in[2] ,
         \SB2_2_1/Component_Function_0/NAND4_in[1] ,
         \SB2_2_1/Component_Function_0/NAND4_in[0] ,
         \SB2_2_1/Component_Function_1/NAND4_in[3] ,
         \SB2_2_1/Component_Function_1/NAND4_in[2] ,
         \SB2_2_1/Component_Function_1/NAND4_in[1] ,
         \SB2_2_1/Component_Function_1/NAND4_in[0] ,
         \SB2_2_1/Component_Function_5/NAND4_in[2] ,
         \SB2_2_1/Component_Function_5/NAND4_in[1] ,
         \SB2_2_1/Component_Function_5/NAND4_in[0] ,
         \SB2_2_2/Component_Function_0/NAND4_in[3] ,
         \SB2_2_2/Component_Function_0/NAND4_in[1] ,
         \SB2_2_2/Component_Function_0/NAND4_in[0] ,
         \SB2_2_2/Component_Function_1/NAND4_in[2] ,
         \SB2_2_2/Component_Function_1/NAND4_in[1] ,
         \SB2_2_2/Component_Function_1/NAND4_in[0] ,
         \SB2_2_2/Component_Function_5/NAND4_in[0] ,
         \SB2_2_3/Component_Function_0/NAND4_in[1] ,
         \SB2_2_3/Component_Function_0/NAND4_in[0] ,
         \SB2_2_3/Component_Function_1/NAND4_in[3] ,
         \SB2_2_3/Component_Function_1/NAND4_in[2] ,
         \SB2_2_3/Component_Function_1/NAND4_in[1] ,
         \SB2_2_3/Component_Function_1/NAND4_in[0] ,
         \SB2_2_3/Component_Function_5/NAND4_in[2] ,
         \SB2_2_3/Component_Function_5/NAND4_in[1] ,
         \SB2_2_3/Component_Function_5/NAND4_in[0] ,
         \SB2_2_4/Component_Function_0/NAND4_in[2] ,
         \SB2_2_4/Component_Function_0/NAND4_in[1] ,
         \SB2_2_4/Component_Function_0/NAND4_in[0] ,
         \SB2_2_4/Component_Function_1/NAND4_in[3] ,
         \SB2_2_4/Component_Function_1/NAND4_in[2] ,
         \SB2_2_4/Component_Function_1/NAND4_in[1] ,
         \SB2_2_4/Component_Function_5/NAND4_in[2] ,
         \SB2_2_4/Component_Function_5/NAND4_in[1] ,
         \SB2_2_5/Component_Function_0/NAND4_in[3] ,
         \SB2_2_5/Component_Function_0/NAND4_in[2] ,
         \SB2_2_5/Component_Function_0/NAND4_in[1] ,
         \SB2_2_5/Component_Function_0/NAND4_in[0] ,
         \SB2_2_5/Component_Function_1/NAND4_in[3] ,
         \SB2_2_5/Component_Function_1/NAND4_in[1] ,
         \SB2_2_5/Component_Function_1/NAND4_in[0] ,
         \SB2_2_5/Component_Function_5/NAND4_in[1] ,
         \SB2_2_5/Component_Function_5/NAND4_in[0] ,
         \SB2_2_6/Component_Function_0/NAND4_in[3] ,
         \SB2_2_6/Component_Function_0/NAND4_in[1] ,
         \SB2_2_6/Component_Function_0/NAND4_in[0] ,
         \SB2_2_6/Component_Function_1/NAND4_in[3] ,
         \SB2_2_6/Component_Function_1/NAND4_in[2] ,
         \SB2_2_6/Component_Function_1/NAND4_in[1] ,
         \SB2_2_6/Component_Function_1/NAND4_in[0] ,
         \SB2_2_6/Component_Function_5/NAND4_in[2] ,
         \SB2_2_6/Component_Function_5/NAND4_in[0] ,
         \SB2_2_7/Component_Function_0/NAND4_in[2] ,
         \SB2_2_7/Component_Function_0/NAND4_in[1] ,
         \SB2_2_7/Component_Function_0/NAND4_in[0] ,
         \SB2_2_7/Component_Function_1/NAND4_in[2] ,
         \SB2_2_7/Component_Function_1/NAND4_in[1] ,
         \SB2_2_7/Component_Function_1/NAND4_in[0] ,
         \SB2_2_7/Component_Function_5/NAND4_in[1] ,
         \SB2_2_7/Component_Function_5/NAND4_in[0] ,
         \SB2_2_8/Component_Function_0/NAND4_in[2] ,
         \SB2_2_8/Component_Function_0/NAND4_in[1] ,
         \SB2_2_8/Component_Function_0/NAND4_in[0] ,
         \SB2_2_8/Component_Function_1/NAND4_in[2] ,
         \SB2_2_8/Component_Function_1/NAND4_in[1] ,
         \SB2_2_8/Component_Function_1/NAND4_in[0] ,
         \SB2_2_8/Component_Function_5/NAND4_in[2] ,
         \SB2_2_8/Component_Function_5/NAND4_in[1] ,
         \SB2_2_8/Component_Function_5/NAND4_in[0] ,
         \SB2_2_9/Component_Function_0/NAND4_in[2] ,
         \SB2_2_9/Component_Function_0/NAND4_in[1] ,
         \SB2_2_9/Component_Function_0/NAND4_in[0] ,
         \SB2_2_9/Component_Function_1/NAND4_in[2] ,
         \SB2_2_9/Component_Function_5/NAND4_in[3] ,
         \SB2_2_9/Component_Function_5/NAND4_in[0] ,
         \SB2_2_10/Component_Function_0/NAND4_in[3] ,
         \SB2_2_10/Component_Function_0/NAND4_in[2] ,
         \SB2_2_10/Component_Function_0/NAND4_in[1] ,
         \SB2_2_10/Component_Function_0/NAND4_in[0] ,
         \SB2_2_10/Component_Function_1/NAND4_in[2] ,
         \SB2_2_10/Component_Function_1/NAND4_in[1] ,
         \SB2_2_10/Component_Function_1/NAND4_in[0] ,
         \SB2_2_10/Component_Function_5/NAND4_in[2] ,
         \SB2_2_10/Component_Function_5/NAND4_in[1] ,
         \SB2_2_11/Component_Function_0/NAND4_in[3] ,
         \SB2_2_11/Component_Function_0/NAND4_in[1] ,
         \SB2_2_11/Component_Function_0/NAND4_in[0] ,
         \SB2_2_11/Component_Function_1/NAND4_in[2] ,
         \SB2_2_11/Component_Function_1/NAND4_in[1] ,
         \SB2_2_11/Component_Function_1/NAND4_in[0] ,
         \SB2_2_11/Component_Function_5/NAND4_in[3] ,
         \SB2_2_12/Component_Function_0/NAND4_in[1] ,
         \SB2_2_12/Component_Function_0/NAND4_in[0] ,
         \SB2_2_12/Component_Function_1/NAND4_in[2] ,
         \SB2_2_12/Component_Function_1/NAND4_in[1] ,
         \SB2_2_12/Component_Function_1/NAND4_in[0] ,
         \SB2_2_12/Component_Function_5/NAND4_in[2] ,
         \SB2_2_12/Component_Function_5/NAND4_in[1] ,
         \SB2_2_12/Component_Function_5/NAND4_in[0] ,
         \SB2_2_13/Component_Function_0/NAND4_in[2] ,
         \SB2_2_13/Component_Function_0/NAND4_in[1] ,
         \SB2_2_13/Component_Function_0/NAND4_in[0] ,
         \SB2_2_13/Component_Function_1/NAND4_in[3] ,
         \SB2_2_13/Component_Function_1/NAND4_in[2] ,
         \SB2_2_13/Component_Function_1/NAND4_in[1] ,
         \SB2_2_13/Component_Function_1/NAND4_in[0] ,
         \SB2_2_13/Component_Function_5/NAND4_in[3] ,
         \SB2_2_13/Component_Function_5/NAND4_in[2] ,
         \SB2_2_13/Component_Function_5/NAND4_in[1] ,
         \SB2_2_13/Component_Function_5/NAND4_in[0] ,
         \SB2_2_14/Component_Function_0/NAND4_in[3] ,
         \SB2_2_14/Component_Function_0/NAND4_in[2] ,
         \SB2_2_14/Component_Function_0/NAND4_in[1] ,
         \SB2_2_14/Component_Function_0/NAND4_in[0] ,
         \SB2_2_14/Component_Function_1/NAND4_in[3] ,
         \SB2_2_14/Component_Function_1/NAND4_in[2] ,
         \SB2_2_14/Component_Function_1/NAND4_in[1] ,
         \SB2_2_14/Component_Function_1/NAND4_in[0] ,
         \SB2_2_14/Component_Function_5/NAND4_in[1] ,
         \SB2_2_14/Component_Function_5/NAND4_in[0] ,
         \SB2_2_15/Component_Function_0/NAND4_in[3] ,
         \SB2_2_15/Component_Function_0/NAND4_in[2] ,
         \SB2_2_15/Component_Function_0/NAND4_in[1] ,
         \SB2_2_15/Component_Function_0/NAND4_in[0] ,
         \SB2_2_15/Component_Function_1/NAND4_in[3] ,
         \SB2_2_15/Component_Function_1/NAND4_in[1] ,
         \SB2_2_15/Component_Function_1/NAND4_in[0] ,
         \SB2_2_15/Component_Function_5/NAND4_in[3] ,
         \SB2_2_15/Component_Function_5/NAND4_in[1] ,
         \SB2_2_15/Component_Function_5/NAND4_in[0] ,
         \SB2_2_16/Component_Function_0/NAND4_in[1] ,
         \SB2_2_16/Component_Function_0/NAND4_in[0] ,
         \SB2_2_16/Component_Function_1/NAND4_in[3] ,
         \SB2_2_16/Component_Function_1/NAND4_in[2] ,
         \SB2_2_16/Component_Function_1/NAND4_in[0] ,
         \SB2_2_16/Component_Function_5/NAND4_in[3] ,
         \SB2_2_16/Component_Function_5/NAND4_in[1] ,
         \SB2_2_16/Component_Function_5/NAND4_in[0] ,
         \SB2_2_17/Component_Function_0/NAND4_in[1] ,
         \SB2_2_17/Component_Function_0/NAND4_in[0] ,
         \SB2_2_17/Component_Function_1/NAND4_in[3] ,
         \SB2_2_17/Component_Function_1/NAND4_in[2] ,
         \SB2_2_17/Component_Function_1/NAND4_in[1] ,
         \SB2_2_17/Component_Function_5/NAND4_in[2] ,
         \SB2_2_17/Component_Function_5/NAND4_in[1] ,
         \SB2_2_17/Component_Function_5/NAND4_in[0] ,
         \SB2_2_18/Component_Function_0/NAND4_in[3] ,
         \SB2_2_18/Component_Function_0/NAND4_in[2] ,
         \SB2_2_18/Component_Function_0/NAND4_in[0] ,
         \SB2_2_18/Component_Function_1/NAND4_in[3] ,
         \SB2_2_18/Component_Function_1/NAND4_in[2] ,
         \SB2_2_18/Component_Function_1/NAND4_in[1] ,
         \SB2_2_18/Component_Function_1/NAND4_in[0] ,
         \SB2_2_18/Component_Function_5/NAND4_in[3] ,
         \SB2_2_18/Component_Function_5/NAND4_in[2] ,
         \SB2_2_18/Component_Function_5/NAND4_in[1] ,
         \SB2_2_18/Component_Function_5/NAND4_in[0] ,
         \SB2_2_19/Component_Function_0/NAND4_in[2] ,
         \SB2_2_19/Component_Function_0/NAND4_in[1] ,
         \SB2_2_19/Component_Function_0/NAND4_in[0] ,
         \SB2_2_19/Component_Function_1/NAND4_in[3] ,
         \SB2_2_19/Component_Function_1/NAND4_in[2] ,
         \SB2_2_19/Component_Function_1/NAND4_in[1] ,
         \SB2_2_19/Component_Function_1/NAND4_in[0] ,
         \SB2_2_19/Component_Function_5/NAND4_in[3] ,
         \SB2_2_19/Component_Function_5/NAND4_in[1] ,
         \SB2_2_19/Component_Function_5/NAND4_in[0] ,
         \SB2_2_20/Component_Function_0/NAND4_in[3] ,
         \SB2_2_20/Component_Function_0/NAND4_in[1] ,
         \SB2_2_20/Component_Function_0/NAND4_in[0] ,
         \SB2_2_20/Component_Function_1/NAND4_in[3] ,
         \SB2_2_20/Component_Function_1/NAND4_in[2] ,
         \SB2_2_20/Component_Function_1/NAND4_in[1] ,
         \SB2_2_20/Component_Function_1/NAND4_in[0] ,
         \SB2_2_20/Component_Function_5/NAND4_in[3] ,
         \SB2_2_20/Component_Function_5/NAND4_in[2] ,
         \SB2_2_20/Component_Function_5/NAND4_in[1] ,
         \SB2_2_20/Component_Function_5/NAND4_in[0] ,
         \SB2_2_21/Component_Function_0/NAND4_in[1] ,
         \SB2_2_21/Component_Function_0/NAND4_in[0] ,
         \SB2_2_21/Component_Function_1/NAND4_in[3] ,
         \SB2_2_21/Component_Function_1/NAND4_in[2] ,
         \SB2_2_21/Component_Function_1/NAND4_in[1] ,
         \SB2_2_21/Component_Function_1/NAND4_in[0] ,
         \SB2_2_21/Component_Function_5/NAND4_in[2] ,
         \SB2_2_21/Component_Function_5/NAND4_in[1] ,
         \SB2_2_21/Component_Function_5/NAND4_in[0] ,
         \SB2_2_22/Component_Function_0/NAND4_in[1] ,
         \SB2_2_22/Component_Function_0/NAND4_in[0] ,
         \SB2_2_22/Component_Function_1/NAND4_in[3] ,
         \SB2_2_22/Component_Function_1/NAND4_in[1] ,
         \SB2_2_22/Component_Function_1/NAND4_in[0] ,
         \SB2_2_22/Component_Function_5/NAND4_in[2] ,
         \SB2_2_22/Component_Function_5/NAND4_in[1] ,
         \SB2_2_23/Component_Function_0/NAND4_in[3] ,
         \SB2_2_23/Component_Function_0/NAND4_in[2] ,
         \SB2_2_23/Component_Function_0/NAND4_in[1] ,
         \SB2_2_23/Component_Function_0/NAND4_in[0] ,
         \SB2_2_23/Component_Function_1/NAND4_in[3] ,
         \SB2_2_23/Component_Function_1/NAND4_in[1] ,
         \SB2_2_23/Component_Function_1/NAND4_in[0] ,
         \SB2_2_23/Component_Function_5/NAND4_in[3] ,
         \SB2_2_23/Component_Function_5/NAND4_in[2] ,
         \SB2_2_23/Component_Function_5/NAND4_in[0] ,
         \SB2_2_24/Component_Function_0/NAND4_in[2] ,
         \SB2_2_24/Component_Function_0/NAND4_in[1] ,
         \SB2_2_24/Component_Function_0/NAND4_in[0] ,
         \SB2_2_24/Component_Function_1/NAND4_in[3] ,
         \SB2_2_24/Component_Function_1/NAND4_in[2] ,
         \SB2_2_24/Component_Function_1/NAND4_in[1] ,
         \SB2_2_24/Component_Function_1/NAND4_in[0] ,
         \SB2_2_24/Component_Function_5/NAND4_in[2] ,
         \SB2_2_24/Component_Function_5/NAND4_in[0] ,
         \SB2_2_25/Component_Function_0/NAND4_in[0] ,
         \SB2_2_25/Component_Function_1/NAND4_in[2] ,
         \SB2_2_25/Component_Function_1/NAND4_in[1] ,
         \SB2_2_25/Component_Function_1/NAND4_in[0] ,
         \SB2_2_25/Component_Function_5/NAND4_in[2] ,
         \SB2_2_25/Component_Function_5/NAND4_in[1] ,
         \SB2_2_25/Component_Function_5/NAND4_in[0] ,
         \SB2_2_26/Component_Function_0/NAND4_in[1] ,
         \SB2_2_26/Component_Function_0/NAND4_in[0] ,
         \SB2_2_26/Component_Function_1/NAND4_in[2] ,
         \SB2_2_26/Component_Function_1/NAND4_in[1] ,
         \SB2_2_26/Component_Function_1/NAND4_in[0] ,
         \SB2_2_26/Component_Function_5/NAND4_in[2] ,
         \SB2_2_26/Component_Function_5/NAND4_in[0] ,
         \SB2_2_27/Component_Function_0/NAND4_in[3] ,
         \SB2_2_27/Component_Function_0/NAND4_in[1] ,
         \SB2_2_27/Component_Function_0/NAND4_in[0] ,
         \SB2_2_27/Component_Function_1/NAND4_in[2] ,
         \SB2_2_27/Component_Function_1/NAND4_in[1] ,
         \SB2_2_27/Component_Function_1/NAND4_in[0] ,
         \SB2_2_27/Component_Function_5/NAND4_in[0] ,
         \SB2_2_28/Component_Function_0/NAND4_in[1] ,
         \SB2_2_28/Component_Function_0/NAND4_in[0] ,
         \SB2_2_28/Component_Function_1/NAND4_in[2] ,
         \SB2_2_28/Component_Function_1/NAND4_in[1] ,
         \SB2_2_28/Component_Function_1/NAND4_in[0] ,
         \SB2_2_28/Component_Function_5/NAND4_in[2] ,
         \SB2_2_28/Component_Function_5/NAND4_in[1] ,
         \SB2_2_28/Component_Function_5/NAND4_in[0] ,
         \SB2_2_29/Component_Function_0/NAND4_in[3] ,
         \SB2_2_29/Component_Function_0/NAND4_in[2] ,
         \SB2_2_29/Component_Function_0/NAND4_in[1] ,
         \SB2_2_29/Component_Function_0/NAND4_in[0] ,
         \SB2_2_29/Component_Function_1/NAND4_in[3] ,
         \SB2_2_29/Component_Function_1/NAND4_in[2] ,
         \SB2_2_29/Component_Function_1/NAND4_in[1] ,
         \SB2_2_29/Component_Function_1/NAND4_in[0] ,
         \SB2_2_29/Component_Function_5/NAND4_in[2] ,
         \SB2_2_29/Component_Function_5/NAND4_in[1] ,
         \SB2_2_29/Component_Function_5/NAND4_in[0] ,
         \SB2_2_30/Component_Function_0/NAND4_in[1] ,
         \SB2_2_30/Component_Function_0/NAND4_in[0] ,
         \SB2_2_30/Component_Function_1/NAND4_in[3] ,
         \SB2_2_30/Component_Function_1/NAND4_in[2] ,
         \SB2_2_30/Component_Function_1/NAND4_in[1] ,
         \SB2_2_30/Component_Function_1/NAND4_in[0] ,
         \SB2_2_30/Component_Function_5/NAND4_in[3] ,
         \SB2_2_30/Component_Function_5/NAND4_in[0] ,
         \SB2_2_31/Component_Function_0/NAND4_in[1] ,
         \SB2_2_31/Component_Function_1/NAND4_in[1] ,
         \SB2_2_31/Component_Function_1/NAND4_in[0] ,
         \SB2_2_31/Component_Function_5/NAND4_in[0] ,
         \SB1_3_0/Component_Function_0/NAND4_in[1] ,
         \SB1_3_0/Component_Function_0/NAND4_in[0] ,
         \SB1_3_0/Component_Function_1/NAND4_in[3] ,
         \SB1_3_0/Component_Function_1/NAND4_in[1] ,
         \SB1_3_0/Component_Function_1/NAND4_in[0] ,
         \SB1_3_0/Component_Function_5/NAND4_in[2] ,
         \SB1_3_0/Component_Function_5/NAND4_in[1] ,
         \SB1_3_0/Component_Function_5/NAND4_in[0] ,
         \SB1_3_1/Component_Function_0/NAND4_in[2] ,
         \SB1_3_1/Component_Function_0/NAND4_in[1] ,
         \SB1_3_1/Component_Function_0/NAND4_in[0] ,
         \SB1_3_1/Component_Function_1/NAND4_in[3] ,
         \SB1_3_1/Component_Function_1/NAND4_in[2] ,
         \SB1_3_1/Component_Function_1/NAND4_in[1] ,
         \SB1_3_1/Component_Function_1/NAND4_in[0] ,
         \SB1_3_1/Component_Function_5/NAND4_in[2] ,
         \SB1_3_1/Component_Function_5/NAND4_in[0] ,
         \SB1_3_2/Component_Function_0/NAND4_in[2] ,
         \SB1_3_2/Component_Function_0/NAND4_in[1] ,
         \SB1_3_2/Component_Function_0/NAND4_in[0] ,
         \SB1_3_2/Component_Function_1/NAND4_in[2] ,
         \SB1_3_2/Component_Function_1/NAND4_in[1] ,
         \SB1_3_2/Component_Function_1/NAND4_in[0] ,
         \SB1_3_2/Component_Function_5/NAND4_in[1] ,
         \SB1_3_2/Component_Function_5/NAND4_in[0] ,
         \SB1_3_3/Component_Function_0/NAND4_in[3] ,
         \SB1_3_3/Component_Function_0/NAND4_in[2] ,
         \SB1_3_3/Component_Function_0/NAND4_in[0] ,
         \SB1_3_3/Component_Function_1/NAND4_in[3] ,
         \SB1_3_3/Component_Function_1/NAND4_in[1] ,
         \SB1_3_3/Component_Function_1/NAND4_in[0] ,
         \SB1_3_3/Component_Function_5/NAND4_in[2] ,
         \SB1_3_3/Component_Function_5/NAND4_in[1] ,
         \SB1_3_3/Component_Function_5/NAND4_in[0] ,
         \SB1_3_4/Component_Function_0/NAND4_in[3] ,
         \SB1_3_4/Component_Function_0/NAND4_in[2] ,
         \SB1_3_4/Component_Function_0/NAND4_in[1] ,
         \SB1_3_4/Component_Function_0/NAND4_in[0] ,
         \SB1_3_4/Component_Function_1/NAND4_in[3] ,
         \SB1_3_4/Component_Function_1/NAND4_in[2] ,
         \SB1_3_4/Component_Function_1/NAND4_in[0] ,
         \SB1_3_4/Component_Function_5/NAND4_in[1] ,
         \SB1_3_4/Component_Function_5/NAND4_in[0] ,
         \SB1_3_5/Component_Function_0/NAND4_in[2] ,
         \SB1_3_5/Component_Function_0/NAND4_in[1] ,
         \SB1_3_5/Component_Function_0/NAND4_in[0] ,
         \SB1_3_5/Component_Function_1/NAND4_in[3] ,
         \SB1_3_5/Component_Function_1/NAND4_in[2] ,
         \SB1_3_5/Component_Function_1/NAND4_in[1] ,
         \SB1_3_5/Component_Function_1/NAND4_in[0] ,
         \SB1_3_5/Component_Function_5/NAND4_in[0] ,
         \SB1_3_6/Component_Function_0/NAND4_in[3] ,
         \SB1_3_6/Component_Function_0/NAND4_in[1] ,
         \SB1_3_6/Component_Function_0/NAND4_in[0] ,
         \SB1_3_6/Component_Function_1/NAND4_in[2] ,
         \SB1_3_6/Component_Function_1/NAND4_in[1] ,
         \SB1_3_6/Component_Function_1/NAND4_in[0] ,
         \SB1_3_6/Component_Function_5/NAND4_in[1] ,
         \SB1_3_6/Component_Function_5/NAND4_in[0] ,
         \SB1_3_7/Component_Function_0/NAND4_in[2] ,
         \SB1_3_7/Component_Function_0/NAND4_in[1] ,
         \SB1_3_7/Component_Function_0/NAND4_in[0] ,
         \SB1_3_7/Component_Function_1/NAND4_in[3] ,
         \SB1_3_7/Component_Function_1/NAND4_in[2] ,
         \SB1_3_7/Component_Function_1/NAND4_in[1] ,
         \SB1_3_7/Component_Function_1/NAND4_in[0] ,
         \SB1_3_7/Component_Function_5/NAND4_in[2] ,
         \SB1_3_7/Component_Function_5/NAND4_in[1] ,
         \SB1_3_8/Component_Function_0/NAND4_in[3] ,
         \SB1_3_8/Component_Function_0/NAND4_in[2] ,
         \SB1_3_8/Component_Function_0/NAND4_in[1] ,
         \SB1_3_8/Component_Function_1/NAND4_in[3] ,
         \SB1_3_8/Component_Function_1/NAND4_in[2] ,
         \SB1_3_8/Component_Function_1/NAND4_in[1] ,
         \SB1_3_8/Component_Function_1/NAND4_in[0] ,
         \SB1_3_8/Component_Function_5/NAND4_in[1] ,
         \SB1_3_9/Component_Function_0/NAND4_in[3] ,
         \SB1_3_9/Component_Function_0/NAND4_in[2] ,
         \SB1_3_9/Component_Function_0/NAND4_in[1] ,
         \SB1_3_9/Component_Function_0/NAND4_in[0] ,
         \SB1_3_9/Component_Function_1/NAND4_in[3] ,
         \SB1_3_9/Component_Function_1/NAND4_in[2] ,
         \SB1_3_9/Component_Function_1/NAND4_in[1] ,
         \SB1_3_9/Component_Function_1/NAND4_in[0] ,
         \SB1_3_9/Component_Function_5/NAND4_in[2] ,
         \SB1_3_10/Component_Function_0/NAND4_in[2] ,
         \SB1_3_10/Component_Function_0/NAND4_in[1] ,
         \SB1_3_10/Component_Function_0/NAND4_in[0] ,
         \SB1_3_10/Component_Function_1/NAND4_in[3] ,
         \SB1_3_10/Component_Function_1/NAND4_in[1] ,
         \SB1_3_10/Component_Function_1/NAND4_in[0] ,
         \SB1_3_10/Component_Function_5/NAND4_in[3] ,
         \SB1_3_10/Component_Function_5/NAND4_in[1] ,
         \SB1_3_10/Component_Function_5/NAND4_in[0] ,
         \SB1_3_11/Component_Function_0/NAND4_in[3] ,
         \SB1_3_11/Component_Function_0/NAND4_in[2] ,
         \SB1_3_11/Component_Function_0/NAND4_in[1] ,
         \SB1_3_11/Component_Function_0/NAND4_in[0] ,
         \SB1_3_11/Component_Function_1/NAND4_in[3] ,
         \SB1_3_11/Component_Function_1/NAND4_in[1] ,
         \SB1_3_11/Component_Function_1/NAND4_in[0] ,
         \SB1_3_11/Component_Function_5/NAND4_in[3] ,
         \SB1_3_11/Component_Function_5/NAND4_in[2] ,
         \SB1_3_11/Component_Function_5/NAND4_in[1] ,
         \SB1_3_11/Component_Function_5/NAND4_in[0] ,
         \SB1_3_12/Component_Function_0/NAND4_in[3] ,
         \SB1_3_12/Component_Function_0/NAND4_in[2] ,
         \SB1_3_12/Component_Function_0/NAND4_in[1] ,
         \SB1_3_12/Component_Function_0/NAND4_in[0] ,
         \SB1_3_12/Component_Function_1/NAND4_in[3] ,
         \SB1_3_12/Component_Function_1/NAND4_in[1] ,
         \SB1_3_12/Component_Function_1/NAND4_in[0] ,
         \SB1_3_12/Component_Function_5/NAND4_in[1] ,
         \SB1_3_12/Component_Function_5/NAND4_in[0] ,
         \SB1_3_13/Component_Function_0/NAND4_in[3] ,
         \SB1_3_13/Component_Function_0/NAND4_in[2] ,
         \SB1_3_13/Component_Function_0/NAND4_in[1] ,
         \SB1_3_13/Component_Function_0/NAND4_in[0] ,
         \SB1_3_13/Component_Function_1/NAND4_in[3] ,
         \SB1_3_13/Component_Function_1/NAND4_in[2] ,
         \SB1_3_13/Component_Function_1/NAND4_in[1] ,
         \SB1_3_13/Component_Function_1/NAND4_in[0] ,
         \SB1_3_13/Component_Function_5/NAND4_in[2] ,
         \SB1_3_13/Component_Function_5/NAND4_in[1] ,
         \SB1_3_13/Component_Function_5/NAND4_in[0] ,
         \SB1_3_14/Component_Function_0/NAND4_in[3] ,
         \SB1_3_14/Component_Function_0/NAND4_in[2] ,
         \SB1_3_14/Component_Function_0/NAND4_in[1] ,
         \SB1_3_14/Component_Function_0/NAND4_in[0] ,
         \SB1_3_14/Component_Function_1/NAND4_in[3] ,
         \SB1_3_14/Component_Function_1/NAND4_in[2] ,
         \SB1_3_14/Component_Function_1/NAND4_in[1] ,
         \SB1_3_14/Component_Function_1/NAND4_in[0] ,
         \SB1_3_14/Component_Function_5/NAND4_in[3] ,
         \SB1_3_14/Component_Function_5/NAND4_in[2] ,
         \SB1_3_14/Component_Function_5/NAND4_in[1] ,
         \SB1_3_15/Component_Function_0/NAND4_in[3] ,
         \SB1_3_15/Component_Function_0/NAND4_in[2] ,
         \SB1_3_15/Component_Function_0/NAND4_in[1] ,
         \SB1_3_15/Component_Function_0/NAND4_in[0] ,
         \SB1_3_15/Component_Function_1/NAND4_in[3] ,
         \SB1_3_15/Component_Function_1/NAND4_in[2] ,
         \SB1_3_15/Component_Function_1/NAND4_in[1] ,
         \SB1_3_15/Component_Function_1/NAND4_in[0] ,
         \SB1_3_15/Component_Function_5/NAND4_in[2] ,
         \SB1_3_15/Component_Function_5/NAND4_in[0] ,
         \SB1_3_16/Component_Function_0/NAND4_in[3] ,
         \SB1_3_16/Component_Function_0/NAND4_in[2] ,
         \SB1_3_16/Component_Function_0/NAND4_in[1] ,
         \SB1_3_16/Component_Function_0/NAND4_in[0] ,
         \SB1_3_16/Component_Function_1/NAND4_in[2] ,
         \SB1_3_16/Component_Function_1/NAND4_in[1] ,
         \SB1_3_16/Component_Function_1/NAND4_in[0] ,
         \SB1_3_16/Component_Function_5/NAND4_in[2] ,
         \SB1_3_16/Component_Function_5/NAND4_in[1] ,
         \SB1_3_16/Component_Function_5/NAND4_in[0] ,
         \SB1_3_17/Component_Function_0/NAND4_in[3] ,
         \SB1_3_17/Component_Function_0/NAND4_in[2] ,
         \SB1_3_17/Component_Function_0/NAND4_in[1] ,
         \SB1_3_17/Component_Function_0/NAND4_in[0] ,
         \SB1_3_17/Component_Function_1/NAND4_in[3] ,
         \SB1_3_17/Component_Function_5/NAND4_in[3] ,
         \SB1_3_17/Component_Function_5/NAND4_in[1] ,
         \SB1_3_17/Component_Function_5/NAND4_in[0] ,
         \SB1_3_18/Component_Function_0/NAND4_in[3] ,
         \SB1_3_18/Component_Function_0/NAND4_in[2] ,
         \SB1_3_18/Component_Function_0/NAND4_in[1] ,
         \SB1_3_18/Component_Function_0/NAND4_in[0] ,
         \SB1_3_18/Component_Function_1/NAND4_in[3] ,
         \SB1_3_18/Component_Function_1/NAND4_in[2] ,
         \SB1_3_18/Component_Function_1/NAND4_in[1] ,
         \SB1_3_18/Component_Function_1/NAND4_in[0] ,
         \SB1_3_18/Component_Function_5/NAND4_in[1] ,
         \SB1_3_18/Component_Function_5/NAND4_in[0] ,
         \SB1_3_19/Component_Function_0/NAND4_in[2] ,
         \SB1_3_19/Component_Function_0/NAND4_in[1] ,
         \SB1_3_19/Component_Function_0/NAND4_in[0] ,
         \SB1_3_19/Component_Function_1/NAND4_in[2] ,
         \SB1_3_19/Component_Function_1/NAND4_in[1] ,
         \SB1_3_19/Component_Function_1/NAND4_in[0] ,
         \SB1_3_19/Component_Function_5/NAND4_in[3] ,
         \SB1_3_19/Component_Function_5/NAND4_in[0] ,
         \SB1_3_20/Component_Function_0/NAND4_in[3] ,
         \SB1_3_20/Component_Function_0/NAND4_in[2] ,
         \SB1_3_20/Component_Function_0/NAND4_in[1] ,
         \SB1_3_20/Component_Function_0/NAND4_in[0] ,
         \SB1_3_20/Component_Function_1/NAND4_in[2] ,
         \SB1_3_20/Component_Function_1/NAND4_in[1] ,
         \SB1_3_20/Component_Function_1/NAND4_in[0] ,
         \SB1_3_20/Component_Function_5/NAND4_in[0] ,
         \SB1_3_21/Component_Function_0/NAND4_in[2] ,
         \SB1_3_21/Component_Function_0/NAND4_in[1] ,
         \SB1_3_21/Component_Function_0/NAND4_in[0] ,
         \SB1_3_21/Component_Function_1/NAND4_in[2] ,
         \SB1_3_21/Component_Function_1/NAND4_in[1] ,
         \SB1_3_21/Component_Function_1/NAND4_in[0] ,
         \SB1_3_21/Component_Function_5/NAND4_in[2] ,
         \SB1_3_21/Component_Function_5/NAND4_in[1] ,
         \SB1_3_22/Component_Function_0/NAND4_in[3] ,
         \SB1_3_22/Component_Function_0/NAND4_in[2] ,
         \SB1_3_22/Component_Function_0/NAND4_in[1] ,
         \SB1_3_22/Component_Function_0/NAND4_in[0] ,
         \SB1_3_22/Component_Function_1/NAND4_in[2] ,
         \SB1_3_22/Component_Function_1/NAND4_in[1] ,
         \SB1_3_22/Component_Function_1/NAND4_in[0] ,
         \SB1_3_22/Component_Function_5/NAND4_in[3] ,
         \SB1_3_23/Component_Function_0/NAND4_in[2] ,
         \SB1_3_23/Component_Function_0/NAND4_in[1] ,
         \SB1_3_23/Component_Function_0/NAND4_in[0] ,
         \SB1_3_23/Component_Function_1/NAND4_in[2] ,
         \SB1_3_23/Component_Function_1/NAND4_in[1] ,
         \SB1_3_23/Component_Function_1/NAND4_in[0] ,
         \SB1_3_23/Component_Function_5/NAND4_in[2] ,
         \SB1_3_23/Component_Function_5/NAND4_in[1] ,
         \SB1_3_23/Component_Function_5/NAND4_in[0] ,
         \SB1_3_24/Component_Function_0/NAND4_in[3] ,
         \SB1_3_24/Component_Function_0/NAND4_in[2] ,
         \SB1_3_24/Component_Function_0/NAND4_in[1] ,
         \SB1_3_24/Component_Function_0/NAND4_in[0] ,
         \SB1_3_24/Component_Function_1/NAND4_in[3] ,
         \SB1_3_24/Component_Function_1/NAND4_in[2] ,
         \SB1_3_24/Component_Function_1/NAND4_in[1] ,
         \SB1_3_24/Component_Function_1/NAND4_in[0] ,
         \SB1_3_24/Component_Function_5/NAND4_in[2] ,
         \SB1_3_24/Component_Function_5/NAND4_in[1] ,
         \SB1_3_24/Component_Function_5/NAND4_in[0] ,
         \SB1_3_25/Component_Function_0/NAND4_in[2] ,
         \SB1_3_25/Component_Function_0/NAND4_in[1] ,
         \SB1_3_25/Component_Function_1/NAND4_in[3] ,
         \SB1_3_25/Component_Function_1/NAND4_in[2] ,
         \SB1_3_25/Component_Function_1/NAND4_in[1] ,
         \SB1_3_25/Component_Function_1/NAND4_in[0] ,
         \SB1_3_25/Component_Function_5/NAND4_in[3] ,
         \SB1_3_25/Component_Function_5/NAND4_in[0] ,
         \SB1_3_26/Component_Function_0/NAND4_in[2] ,
         \SB1_3_26/Component_Function_0/NAND4_in[1] ,
         \SB1_3_26/Component_Function_0/NAND4_in[0] ,
         \SB1_3_26/Component_Function_1/NAND4_in[3] ,
         \SB1_3_26/Component_Function_1/NAND4_in[1] ,
         \SB1_3_26/Component_Function_1/NAND4_in[0] ,
         \SB1_3_26/Component_Function_5/NAND4_in[3] ,
         \SB1_3_26/Component_Function_5/NAND4_in[2] ,
         \SB1_3_26/Component_Function_5/NAND4_in[0] ,
         \SB1_3_27/Component_Function_0/NAND4_in[3] ,
         \SB1_3_27/Component_Function_0/NAND4_in[2] ,
         \SB1_3_27/Component_Function_0/NAND4_in[0] ,
         \SB1_3_27/Component_Function_1/NAND4_in[3] ,
         \SB1_3_27/Component_Function_1/NAND4_in[1] ,
         \SB1_3_27/Component_Function_1/NAND4_in[0] ,
         \SB1_3_27/Component_Function_5/NAND4_in[1] ,
         \SB1_3_27/Component_Function_5/NAND4_in[0] ,
         \SB1_3_28/Component_Function_0/NAND4_in[3] ,
         \SB1_3_28/Component_Function_0/NAND4_in[2] ,
         \SB1_3_28/Component_Function_0/NAND4_in[1] ,
         \SB1_3_28/Component_Function_1/NAND4_in[3] ,
         \SB1_3_28/Component_Function_1/NAND4_in[2] ,
         \SB1_3_28/Component_Function_1/NAND4_in[1] ,
         \SB1_3_28/Component_Function_1/NAND4_in[0] ,
         \SB1_3_28/Component_Function_5/NAND4_in[2] ,
         \SB1_3_28/Component_Function_5/NAND4_in[1] ,
         \SB1_3_28/Component_Function_5/NAND4_in[0] ,
         \SB1_3_29/Component_Function_0/NAND4_in[2] ,
         \SB1_3_29/Component_Function_0/NAND4_in[1] ,
         \SB1_3_29/Component_Function_0/NAND4_in[0] ,
         \SB1_3_29/Component_Function_1/NAND4_in[3] ,
         \SB1_3_29/Component_Function_1/NAND4_in[2] ,
         \SB1_3_29/Component_Function_1/NAND4_in[1] ,
         \SB1_3_29/Component_Function_1/NAND4_in[0] ,
         \SB1_3_29/Component_Function_5/NAND4_in[2] ,
         \SB1_3_29/Component_Function_5/NAND4_in[0] ,
         \SB1_3_30/Component_Function_0/NAND4_in[3] ,
         \SB1_3_30/Component_Function_0/NAND4_in[1] ,
         \SB1_3_30/Component_Function_1/NAND4_in[2] ,
         \SB1_3_30/Component_Function_1/NAND4_in[1] ,
         \SB1_3_30/Component_Function_1/NAND4_in[0] ,
         \SB1_3_30/Component_Function_5/NAND4_in[2] ,
         \SB1_3_30/Component_Function_5/NAND4_in[1] ,
         \SB1_3_30/Component_Function_5/NAND4_in[0] ,
         \SB1_3_31/Component_Function_0/NAND4_in[2] ,
         \SB1_3_31/Component_Function_0/NAND4_in[1] ,
         \SB1_3_31/Component_Function_1/NAND4_in[3] ,
         \SB1_3_31/Component_Function_1/NAND4_in[0] ,
         \SB1_3_31/Component_Function_5/NAND4_in[2] ,
         \SB1_3_31/Component_Function_5/NAND4_in[1] ,
         \SB1_3_31/Component_Function_5/NAND4_in[0] ,
         \SB2_3_0/Component_Function_0/NAND4_in[2] ,
         \SB2_3_0/Component_Function_0/NAND4_in[1] ,
         \SB2_3_0/Component_Function_0/NAND4_in[0] ,
         \SB2_3_0/Component_Function_1/NAND4_in[3] ,
         \SB2_3_0/Component_Function_1/NAND4_in[2] ,
         \SB2_3_0/Component_Function_1/NAND4_in[1] ,
         \SB2_3_0/Component_Function_1/NAND4_in[0] ,
         \SB2_3_0/Component_Function_5/NAND4_in[3] ,
         \SB2_3_0/Component_Function_5/NAND4_in[0] ,
         \SB2_3_1/Component_Function_0/NAND4_in[2] ,
         \SB2_3_1/Component_Function_0/NAND4_in[1] ,
         \SB2_3_1/Component_Function_1/NAND4_in[1] ,
         \SB2_3_1/Component_Function_1/NAND4_in[0] ,
         \SB2_3_1/Component_Function_5/NAND4_in[0] ,
         \SB2_3_2/Component_Function_0/NAND4_in[2] ,
         \SB2_3_2/Component_Function_0/NAND4_in[1] ,
         \SB2_3_2/Component_Function_1/NAND4_in[3] ,
         \SB2_3_2/Component_Function_1/NAND4_in[2] ,
         \SB2_3_2/Component_Function_1/NAND4_in[0] ,
         \SB2_3_2/Component_Function_5/NAND4_in[3] ,
         \SB2_3_2/Component_Function_5/NAND4_in[0] ,
         \SB2_3_3/Component_Function_0/NAND4_in[2] ,
         \SB2_3_3/Component_Function_0/NAND4_in[1] ,
         \SB2_3_3/Component_Function_0/NAND4_in[0] ,
         \SB2_3_3/Component_Function_1/NAND4_in[3] ,
         \SB2_3_3/Component_Function_1/NAND4_in[2] ,
         \SB2_3_3/Component_Function_1/NAND4_in[1] ,
         \SB2_3_3/Component_Function_1/NAND4_in[0] ,
         \SB2_3_3/Component_Function_5/NAND4_in[1] ,
         \SB2_3_3/Component_Function_5/NAND4_in[0] ,
         \SB2_3_4/Component_Function_0/NAND4_in[1] ,
         \SB2_3_4/Component_Function_0/NAND4_in[0] ,
         \SB2_3_4/Component_Function_1/NAND4_in[3] ,
         \SB2_3_4/Component_Function_1/NAND4_in[2] ,
         \SB2_3_4/Component_Function_1/NAND4_in[1] ,
         \SB2_3_4/Component_Function_1/NAND4_in[0] ,
         \SB2_3_5/Component_Function_0/NAND4_in[3] ,
         \SB2_3_5/Component_Function_0/NAND4_in[2] ,
         \SB2_3_5/Component_Function_0/NAND4_in[1] ,
         \SB2_3_5/Component_Function_0/NAND4_in[0] ,
         \SB2_3_5/Component_Function_1/NAND4_in[3] ,
         \SB2_3_5/Component_Function_1/NAND4_in[2] ,
         \SB2_3_5/Component_Function_1/NAND4_in[1] ,
         \SB2_3_5/Component_Function_1/NAND4_in[0] ,
         \SB2_3_5/Component_Function_5/NAND4_in[2] ,
         \SB2_3_5/Component_Function_5/NAND4_in[0] ,
         \SB2_3_6/Component_Function_0/NAND4_in[3] ,
         \SB2_3_6/Component_Function_0/NAND4_in[1] ,
         \SB2_3_6/Component_Function_0/NAND4_in[0] ,
         \SB2_3_6/Component_Function_1/NAND4_in[3] ,
         \SB2_3_6/Component_Function_1/NAND4_in[2] ,
         \SB2_3_6/Component_Function_1/NAND4_in[1] ,
         \SB2_3_6/Component_Function_1/NAND4_in[0] ,
         \SB2_3_6/Component_Function_5/NAND4_in[2] ,
         \SB2_3_6/Component_Function_5/NAND4_in[0] ,
         \SB2_3_7/Component_Function_0/NAND4_in[3] ,
         \SB2_3_7/Component_Function_0/NAND4_in[2] ,
         \SB2_3_7/Component_Function_0/NAND4_in[0] ,
         \SB2_3_7/Component_Function_1/NAND4_in[3] ,
         \SB2_3_7/Component_Function_1/NAND4_in[1] ,
         \SB2_3_7/Component_Function_1/NAND4_in[0] ,
         \SB2_3_7/Component_Function_5/NAND4_in[2] ,
         \SB2_3_7/Component_Function_5/NAND4_in[1] ,
         \SB2_3_7/Component_Function_5/NAND4_in[0] ,
         \SB2_3_8/Component_Function_0/NAND4_in[3] ,
         \SB2_3_8/Component_Function_0/NAND4_in[2] ,
         \SB2_3_8/Component_Function_0/NAND4_in[0] ,
         \SB2_3_8/Component_Function_1/NAND4_in[3] ,
         \SB2_3_8/Component_Function_1/NAND4_in[1] ,
         \SB2_3_8/Component_Function_1/NAND4_in[0] ,
         \SB2_3_8/Component_Function_5/NAND4_in[2] ,
         \SB2_3_8/Component_Function_5/NAND4_in[1] ,
         \SB2_3_8/Component_Function_5/NAND4_in[0] ,
         \SB2_3_9/Component_Function_0/NAND4_in[3] ,
         \SB2_3_9/Component_Function_0/NAND4_in[1] ,
         \SB2_3_9/Component_Function_0/NAND4_in[0] ,
         \SB2_3_9/Component_Function_1/NAND4_in[3] ,
         \SB2_3_9/Component_Function_1/NAND4_in[2] ,
         \SB2_3_9/Component_Function_1/NAND4_in[1] ,
         \SB2_3_9/Component_Function_1/NAND4_in[0] ,
         \SB2_3_9/Component_Function_5/NAND4_in[3] ,
         \SB2_3_9/Component_Function_5/NAND4_in[2] ,
         \SB2_3_9/Component_Function_5/NAND4_in[0] ,
         \SB2_3_10/Component_Function_0/NAND4_in[2] ,
         \SB2_3_10/Component_Function_0/NAND4_in[1] ,
         \SB2_3_10/Component_Function_0/NAND4_in[0] ,
         \SB2_3_10/Component_Function_1/NAND4_in[2] ,
         \SB2_3_10/Component_Function_1/NAND4_in[1] ,
         \SB2_3_10/Component_Function_1/NAND4_in[0] ,
         \SB2_3_10/Component_Function_5/NAND4_in[2] ,
         \SB2_3_10/Component_Function_5/NAND4_in[0] ,
         \SB2_3_11/Component_Function_0/NAND4_in[3] ,
         \SB2_3_11/Component_Function_0/NAND4_in[1] ,
         \SB2_3_11/Component_Function_0/NAND4_in[0] ,
         \SB2_3_11/Component_Function_1/NAND4_in[3] ,
         \SB2_3_11/Component_Function_1/NAND4_in[2] ,
         \SB2_3_11/Component_Function_1/NAND4_in[0] ,
         \SB2_3_11/Component_Function_5/NAND4_in[3] ,
         \SB2_3_11/Component_Function_5/NAND4_in[0] ,
         \SB2_3_12/Component_Function_0/NAND4_in[3] ,
         \SB2_3_12/Component_Function_0/NAND4_in[2] ,
         \SB2_3_12/Component_Function_0/NAND4_in[0] ,
         \SB2_3_12/Component_Function_1/NAND4_in[2] ,
         \SB2_3_12/Component_Function_1/NAND4_in[1] ,
         \SB2_3_12/Component_Function_1/NAND4_in[0] ,
         \SB2_3_12/Component_Function_5/NAND4_in[2] ,
         \SB2_3_12/Component_Function_5/NAND4_in[0] ,
         \SB2_3_13/Component_Function_0/NAND4_in[3] ,
         \SB2_3_13/Component_Function_0/NAND4_in[2] ,
         \SB2_3_13/Component_Function_0/NAND4_in[1] ,
         \SB2_3_13/Component_Function_0/NAND4_in[0] ,
         \SB2_3_13/Component_Function_1/NAND4_in[2] ,
         \SB2_3_13/Component_Function_1/NAND4_in[1] ,
         \SB2_3_13/Component_Function_1/NAND4_in[0] ,
         \SB2_3_13/Component_Function_5/NAND4_in[2] ,
         \SB2_3_13/Component_Function_5/NAND4_in[1] ,
         \SB2_3_13/Component_Function_5/NAND4_in[0] ,
         \SB2_3_14/Component_Function_0/NAND4_in[2] ,
         \SB2_3_14/Component_Function_0/NAND4_in[1] ,
         \SB2_3_14/Component_Function_0/NAND4_in[0] ,
         \SB2_3_14/Component_Function_1/NAND4_in[3] ,
         \SB2_3_14/Component_Function_1/NAND4_in[2] ,
         \SB2_3_14/Component_Function_1/NAND4_in[1] ,
         \SB2_3_14/Component_Function_1/NAND4_in[0] ,
         \SB2_3_14/Component_Function_5/NAND4_in[3] ,
         \SB2_3_14/Component_Function_5/NAND4_in[2] ,
         \SB2_3_14/Component_Function_5/NAND4_in[0] ,
         \SB2_3_15/Component_Function_0/NAND4_in[3] ,
         \SB2_3_15/Component_Function_0/NAND4_in[1] ,
         \SB2_3_15/Component_Function_0/NAND4_in[0] ,
         \SB2_3_15/Component_Function_1/NAND4_in[3] ,
         \SB2_3_15/Component_Function_1/NAND4_in[1] ,
         \SB2_3_15/Component_Function_1/NAND4_in[0] ,
         \SB2_3_15/Component_Function_5/NAND4_in[0] ,
         \SB2_3_16/Component_Function_0/NAND4_in[1] ,
         \SB2_3_16/Component_Function_0/NAND4_in[0] ,
         \SB2_3_16/Component_Function_1/NAND4_in[3] ,
         \SB2_3_16/Component_Function_1/NAND4_in[2] ,
         \SB2_3_16/Component_Function_1/NAND4_in[1] ,
         \SB2_3_16/Component_Function_1/NAND4_in[0] ,
         \SB2_3_16/Component_Function_5/NAND4_in[2] ,
         \SB2_3_17/Component_Function_0/NAND4_in[3] ,
         \SB2_3_17/Component_Function_0/NAND4_in[1] ,
         \SB2_3_17/Component_Function_0/NAND4_in[0] ,
         \SB2_3_17/Component_Function_1/NAND4_in[2] ,
         \SB2_3_17/Component_Function_1/NAND4_in[1] ,
         \SB2_3_17/Component_Function_1/NAND4_in[0] ,
         \SB2_3_17/Component_Function_5/NAND4_in[1] ,
         \SB2_3_17/Component_Function_5/NAND4_in[0] ,
         \SB2_3_18/Component_Function_0/NAND4_in[2] ,
         \SB2_3_18/Component_Function_0/NAND4_in[1] ,
         \SB2_3_18/Component_Function_0/NAND4_in[0] ,
         \SB2_3_18/Component_Function_1/NAND4_in[3] ,
         \SB2_3_18/Component_Function_1/NAND4_in[2] ,
         \SB2_3_18/Component_Function_1/NAND4_in[1] ,
         \SB2_3_18/Component_Function_1/NAND4_in[0] ,
         \SB2_3_18/Component_Function_5/NAND4_in[2] ,
         \SB2_3_18/Component_Function_5/NAND4_in[0] ,
         \SB2_3_19/Component_Function_0/NAND4_in[2] ,
         \SB2_3_19/Component_Function_0/NAND4_in[1] ,
         \SB2_3_19/Component_Function_0/NAND4_in[0] ,
         \SB2_3_19/Component_Function_1/NAND4_in[1] ,
         \SB2_3_19/Component_Function_1/NAND4_in[0] ,
         \SB2_3_19/Component_Function_5/NAND4_in[3] ,
         \SB2_3_19/Component_Function_5/NAND4_in[2] ,
         \SB2_3_19/Component_Function_5/NAND4_in[0] ,
         \SB2_3_20/Component_Function_0/NAND4_in[3] ,
         \SB2_3_20/Component_Function_0/NAND4_in[1] ,
         \SB2_3_20/Component_Function_0/NAND4_in[0] ,
         \SB2_3_20/Component_Function_1/NAND4_in[3] ,
         \SB2_3_20/Component_Function_1/NAND4_in[2] ,
         \SB2_3_20/Component_Function_1/NAND4_in[1] ,
         \SB2_3_20/Component_Function_1/NAND4_in[0] ,
         \SB2_3_20/Component_Function_5/NAND4_in[2] ,
         \SB2_3_20/Component_Function_5/NAND4_in[0] ,
         \SB2_3_21/Component_Function_0/NAND4_in[3] ,
         \SB2_3_21/Component_Function_0/NAND4_in[1] ,
         \SB2_3_21/Component_Function_0/NAND4_in[0] ,
         \SB2_3_21/Component_Function_1/NAND4_in[3] ,
         \SB2_3_21/Component_Function_1/NAND4_in[2] ,
         \SB2_3_21/Component_Function_1/NAND4_in[1] ,
         \SB2_3_21/Component_Function_1/NAND4_in[0] ,
         \SB2_3_21/Component_Function_5/NAND4_in[2] ,
         \SB2_3_21/Component_Function_5/NAND4_in[1] ,
         \SB2_3_22/Component_Function_0/NAND4_in[3] ,
         \SB2_3_22/Component_Function_0/NAND4_in[1] ,
         \SB2_3_22/Component_Function_0/NAND4_in[0] ,
         \SB2_3_22/Component_Function_1/NAND4_in[3] ,
         \SB2_3_22/Component_Function_1/NAND4_in[2] ,
         \SB2_3_22/Component_Function_1/NAND4_in[1] ,
         \SB2_3_22/Component_Function_1/NAND4_in[0] ,
         \SB2_3_22/Component_Function_5/NAND4_in[2] ,
         \SB2_3_22/Component_Function_5/NAND4_in[0] ,
         \SB2_3_23/Component_Function_0/NAND4_in[1] ,
         \SB2_3_23/Component_Function_0/NAND4_in[0] ,
         \SB2_3_23/Component_Function_1/NAND4_in[3] ,
         \SB2_3_23/Component_Function_1/NAND4_in[2] ,
         \SB2_3_23/Component_Function_1/NAND4_in[1] ,
         \SB2_3_23/Component_Function_5/NAND4_in[2] ,
         \SB2_3_23/Component_Function_5/NAND4_in[0] ,
         \SB2_3_24/Component_Function_0/NAND4_in[3] ,
         \SB2_3_24/Component_Function_0/NAND4_in[1] ,
         \SB2_3_24/Component_Function_0/NAND4_in[0] ,
         \SB2_3_24/Component_Function_1/NAND4_in[2] ,
         \SB2_3_24/Component_Function_1/NAND4_in[1] ,
         \SB2_3_24/Component_Function_1/NAND4_in[0] ,
         \SB2_3_24/Component_Function_5/NAND4_in[3] ,
         \SB2_3_24/Component_Function_5/NAND4_in[0] ,
         \SB2_3_25/Component_Function_0/NAND4_in[2] ,
         \SB2_3_25/Component_Function_0/NAND4_in[1] ,
         \SB2_3_25/Component_Function_1/NAND4_in[3] ,
         \SB2_3_25/Component_Function_1/NAND4_in[2] ,
         \SB2_3_25/Component_Function_1/NAND4_in[1] ,
         \SB2_3_25/Component_Function_1/NAND4_in[0] ,
         \SB2_3_25/Component_Function_5/NAND4_in[2] ,
         \SB2_3_25/Component_Function_5/NAND4_in[1] ,
         \SB2_3_25/Component_Function_5/NAND4_in[0] ,
         \SB2_3_26/Component_Function_0/NAND4_in[2] ,
         \SB2_3_26/Component_Function_0/NAND4_in[1] ,
         \SB2_3_26/Component_Function_0/NAND4_in[0] ,
         \SB2_3_26/Component_Function_1/NAND4_in[3] ,
         \SB2_3_26/Component_Function_1/NAND4_in[2] ,
         \SB2_3_26/Component_Function_1/NAND4_in[1] ,
         \SB2_3_26/Component_Function_1/NAND4_in[0] ,
         \SB2_3_26/Component_Function_5/NAND4_in[3] ,
         \SB2_3_26/Component_Function_5/NAND4_in[2] ,
         \SB2_3_27/Component_Function_0/NAND4_in[2] ,
         \SB2_3_27/Component_Function_0/NAND4_in[1] ,
         \SB2_3_27/Component_Function_0/NAND4_in[0] ,
         \SB2_3_27/Component_Function_1/NAND4_in[3] ,
         \SB2_3_27/Component_Function_1/NAND4_in[2] ,
         \SB2_3_27/Component_Function_1/NAND4_in[1] ,
         \SB2_3_27/Component_Function_5/NAND4_in[1] ,
         \SB2_3_27/Component_Function_5/NAND4_in[0] ,
         \SB2_3_28/Component_Function_0/NAND4_in[3] ,
         \SB2_3_28/Component_Function_0/NAND4_in[1] ,
         \SB2_3_28/Component_Function_0/NAND4_in[0] ,
         \SB2_3_28/Component_Function_1/NAND4_in[1] ,
         \SB2_3_28/Component_Function_1/NAND4_in[0] ,
         \SB2_3_28/Component_Function_5/NAND4_in[3] ,
         \SB2_3_28/Component_Function_5/NAND4_in[1] ,
         \SB2_3_29/Component_Function_0/NAND4_in[3] ,
         \SB2_3_29/Component_Function_0/NAND4_in[2] ,
         \SB2_3_29/Component_Function_0/NAND4_in[1] ,
         \SB2_3_29/Component_Function_0/NAND4_in[0] ,
         \SB2_3_29/Component_Function_1/NAND4_in[3] ,
         \SB2_3_29/Component_Function_1/NAND4_in[1] ,
         \SB2_3_29/Component_Function_1/NAND4_in[0] ,
         \SB2_3_29/Component_Function_5/NAND4_in[2] ,
         \SB2_3_29/Component_Function_5/NAND4_in[0] ,
         \SB2_3_30/Component_Function_0/NAND4_in[2] ,
         \SB2_3_30/Component_Function_0/NAND4_in[1] ,
         \SB2_3_30/Component_Function_0/NAND4_in[0] ,
         \SB2_3_30/Component_Function_1/NAND4_in[3] ,
         \SB2_3_30/Component_Function_1/NAND4_in[1] ,
         \SB2_3_30/Component_Function_1/NAND4_in[0] ,
         \SB2_3_30/Component_Function_5/NAND4_in[0] ,
         \SB2_3_31/Component_Function_0/NAND4_in[2] ,
         \SB2_3_31/Component_Function_0/NAND4_in[1] ,
         \SB2_3_31/Component_Function_0/NAND4_in[0] ,
         \SB2_3_31/Component_Function_1/NAND4_in[3] ,
         \SB2_3_31/Component_Function_1/NAND4_in[2] ,
         \SB2_3_31/Component_Function_1/NAND4_in[1] ,
         \SB2_3_31/Component_Function_1/NAND4_in[0] ,
         \SB2_3_31/Component_Function_5/NAND4_in[0] ,
         \SB1_4_0/Component_Function_0/NAND4_in[2] ,
         \SB1_4_0/Component_Function_0/NAND4_in[1] ,
         \SB1_4_0/Component_Function_0/NAND4_in[0] ,
         \SB1_4_0/Component_Function_1/NAND4_in[3] ,
         \SB1_4_0/Component_Function_1/NAND4_in[2] ,
         \SB1_4_0/Component_Function_1/NAND4_in[1] ,
         \SB1_4_0/Component_Function_1/NAND4_in[0] ,
         \SB1_4_0/Component_Function_5/NAND4_in[3] ,
         \SB1_4_0/Component_Function_5/NAND4_in[2] ,
         \SB1_4_1/Component_Function_0/NAND4_in[2] ,
         \SB1_4_1/Component_Function_0/NAND4_in[1] ,
         \SB1_4_1/Component_Function_0/NAND4_in[0] ,
         \SB1_4_1/Component_Function_1/NAND4_in[3] ,
         \SB1_4_1/Component_Function_1/NAND4_in[2] ,
         \SB1_4_1/Component_Function_1/NAND4_in[1] ,
         \SB1_4_1/Component_Function_1/NAND4_in[0] ,
         \SB1_4_1/Component_Function_5/NAND4_in[2] ,
         \SB1_4_1/Component_Function_5/NAND4_in[1] ,
         \SB1_4_1/Component_Function_5/NAND4_in[0] ,
         \SB1_4_2/Component_Function_0/NAND4_in[3] ,
         \SB1_4_2/Component_Function_0/NAND4_in[2] ,
         \SB1_4_2/Component_Function_0/NAND4_in[1] ,
         \SB1_4_2/Component_Function_0/NAND4_in[0] ,
         \SB1_4_2/Component_Function_1/NAND4_in[2] ,
         \SB1_4_2/Component_Function_1/NAND4_in[1] ,
         \SB1_4_2/Component_Function_1/NAND4_in[0] ,
         \SB1_4_2/Component_Function_5/NAND4_in[2] ,
         \SB1_4_2/Component_Function_5/NAND4_in[0] ,
         \SB1_4_3/Component_Function_0/NAND4_in[3] ,
         \SB1_4_3/Component_Function_0/NAND4_in[2] ,
         \SB1_4_3/Component_Function_0/NAND4_in[1] ,
         \SB1_4_3/Component_Function_0/NAND4_in[0] ,
         \SB1_4_3/Component_Function_1/NAND4_in[3] ,
         \SB1_4_3/Component_Function_1/NAND4_in[1] ,
         \SB1_4_3/Component_Function_1/NAND4_in[0] ,
         \SB1_4_3/Component_Function_5/NAND4_in[1] ,
         \SB1_4_3/Component_Function_5/NAND4_in[0] ,
         \SB1_4_4/Component_Function_0/NAND4_in[3] ,
         \SB1_4_4/Component_Function_0/NAND4_in[1] ,
         \SB1_4_4/Component_Function_0/NAND4_in[0] ,
         \SB1_4_4/Component_Function_1/NAND4_in[3] ,
         \SB1_4_4/Component_Function_1/NAND4_in[0] ,
         \SB1_4_4/Component_Function_5/NAND4_in[1] ,
         \SB1_4_4/Component_Function_5/NAND4_in[0] ,
         \SB1_4_5/Component_Function_0/NAND4_in[3] ,
         \SB1_4_5/Component_Function_0/NAND4_in[2] ,
         \SB1_4_5/Component_Function_0/NAND4_in[1] ,
         \SB1_4_5/Component_Function_0/NAND4_in[0] ,
         \SB1_4_5/Component_Function_1/NAND4_in[3] ,
         \SB1_4_5/Component_Function_1/NAND4_in[2] ,
         \SB1_4_5/Component_Function_1/NAND4_in[1] ,
         \SB1_4_5/Component_Function_1/NAND4_in[0] ,
         \SB1_4_5/Component_Function_5/NAND4_in[1] ,
         \SB1_4_5/Component_Function_5/NAND4_in[0] ,
         \SB1_4_6/Component_Function_0/NAND4_in[1] ,
         \SB1_4_6/Component_Function_0/NAND4_in[0] ,
         \SB1_4_6/Component_Function_1/NAND4_in[1] ,
         \SB1_4_6/Component_Function_5/NAND4_in[3] ,
         \SB1_4_6/Component_Function_5/NAND4_in[1] ,
         \SB1_4_6/Component_Function_5/NAND4_in[0] ,
         \SB1_4_7/Component_Function_0/NAND4_in[2] ,
         \SB1_4_7/Component_Function_0/NAND4_in[1] ,
         \SB1_4_7/Component_Function_0/NAND4_in[0] ,
         \SB1_4_7/Component_Function_1/NAND4_in[3] ,
         \SB1_4_7/Component_Function_1/NAND4_in[2] ,
         \SB1_4_7/Component_Function_1/NAND4_in[1] ,
         \SB1_4_7/Component_Function_1/NAND4_in[0] ,
         \SB1_4_7/Component_Function_5/NAND4_in[3] ,
         \SB1_4_8/Component_Function_0/NAND4_in[2] ,
         \SB1_4_8/Component_Function_0/NAND4_in[1] ,
         \SB1_4_8/Component_Function_0/NAND4_in[0] ,
         \SB1_4_8/Component_Function_1/NAND4_in[3] ,
         \SB1_4_8/Component_Function_1/NAND4_in[2] ,
         \SB1_4_8/Component_Function_1/NAND4_in[1] ,
         \SB1_4_8/Component_Function_1/NAND4_in[0] ,
         \SB1_4_8/Component_Function_5/NAND4_in[3] ,
         \SB1_4_8/Component_Function_5/NAND4_in[1] ,
         \SB1_4_9/Component_Function_0/NAND4_in[2] ,
         \SB1_4_9/Component_Function_0/NAND4_in[1] ,
         \SB1_4_9/Component_Function_0/NAND4_in[0] ,
         \SB1_4_9/Component_Function_1/NAND4_in[3] ,
         \SB1_4_9/Component_Function_1/NAND4_in[2] ,
         \SB1_4_9/Component_Function_1/NAND4_in[1] ,
         \SB1_4_9/Component_Function_1/NAND4_in[0] ,
         \SB1_4_9/Component_Function_5/NAND4_in[1] ,
         \SB1_4_9/Component_Function_5/NAND4_in[0] ,
         \SB1_4_10/Component_Function_0/NAND4_in[1] ,
         \SB1_4_10/Component_Function_0/NAND4_in[0] ,
         \SB1_4_10/Component_Function_1/NAND4_in[3] ,
         \SB1_4_10/Component_Function_1/NAND4_in[2] ,
         \SB1_4_10/Component_Function_1/NAND4_in[1] ,
         \SB1_4_10/Component_Function_1/NAND4_in[0] ,
         \SB1_4_10/Component_Function_5/NAND4_in[3] ,
         \SB1_4_10/Component_Function_5/NAND4_in[2] ,
         \SB1_4_10/Component_Function_5/NAND4_in[1] ,
         \SB1_4_10/Component_Function_5/NAND4_in[0] ,
         \SB1_4_11/Component_Function_0/NAND4_in[3] ,
         \SB1_4_11/Component_Function_0/NAND4_in[2] ,
         \SB1_4_11/Component_Function_0/NAND4_in[1] ,
         \SB1_4_11/Component_Function_0/NAND4_in[0] ,
         \SB1_4_11/Component_Function_1/NAND4_in[3] ,
         \SB1_4_11/Component_Function_1/NAND4_in[1] ,
         \SB1_4_11/Component_Function_1/NAND4_in[0] ,
         \SB1_4_11/Component_Function_5/NAND4_in[1] ,
         \SB1_4_11/Component_Function_5/NAND4_in[0] ,
         \SB1_4_12/Component_Function_0/NAND4_in[3] ,
         \SB1_4_12/Component_Function_0/NAND4_in[2] ,
         \SB1_4_12/Component_Function_0/NAND4_in[1] ,
         \SB1_4_12/Component_Function_0/NAND4_in[0] ,
         \SB1_4_12/Component_Function_1/NAND4_in[3] ,
         \SB1_4_12/Component_Function_1/NAND4_in[1] ,
         \SB1_4_12/Component_Function_1/NAND4_in[0] ,
         \SB1_4_12/Component_Function_5/NAND4_in[2] ,
         \SB1_4_12/Component_Function_5/NAND4_in[1] ,
         \SB1_4_12/Component_Function_5/NAND4_in[0] ,
         \SB1_4_13/Component_Function_0/NAND4_in[3] ,
         \SB1_4_13/Component_Function_0/NAND4_in[2] ,
         \SB1_4_13/Component_Function_0/NAND4_in[1] ,
         \SB1_4_13/Component_Function_0/NAND4_in[0] ,
         \SB1_4_13/Component_Function_1/NAND4_in[2] ,
         \SB1_4_13/Component_Function_1/NAND4_in[1] ,
         \SB1_4_13/Component_Function_1/NAND4_in[0] ,
         \SB1_4_13/Component_Function_5/NAND4_in[1] ,
         \SB1_4_13/Component_Function_5/NAND4_in[0] ,
         \SB1_4_14/Component_Function_0/NAND4_in[3] ,
         \SB1_4_14/Component_Function_0/NAND4_in[2] ,
         \SB1_4_14/Component_Function_0/NAND4_in[1] ,
         \SB1_4_14/Component_Function_0/NAND4_in[0] ,
         \SB1_4_14/Component_Function_1/NAND4_in[3] ,
         \SB1_4_14/Component_Function_1/NAND4_in[1] ,
         \SB1_4_14/Component_Function_5/NAND4_in[3] ,
         \SB1_4_14/Component_Function_5/NAND4_in[2] ,
         \SB1_4_15/Component_Function_0/NAND4_in[3] ,
         \SB1_4_15/Component_Function_0/NAND4_in[2] ,
         \SB1_4_15/Component_Function_0/NAND4_in[1] ,
         \SB1_4_15/Component_Function_0/NAND4_in[0] ,
         \SB1_4_15/Component_Function_1/NAND4_in[2] ,
         \SB1_4_15/Component_Function_1/NAND4_in[1] ,
         \SB1_4_15/Component_Function_1/NAND4_in[0] ,
         \SB1_4_15/Component_Function_5/NAND4_in[1] ,
         \SB1_4_15/Component_Function_5/NAND4_in[0] ,
         \SB1_4_16/Component_Function_0/NAND4_in[2] ,
         \SB1_4_16/Component_Function_0/NAND4_in[1] ,
         \SB1_4_16/Component_Function_0/NAND4_in[0] ,
         \SB1_4_16/Component_Function_1/NAND4_in[3] ,
         \SB1_4_16/Component_Function_1/NAND4_in[1] ,
         \SB1_4_16/Component_Function_1/NAND4_in[0] ,
         \SB1_4_16/Component_Function_5/NAND4_in[1] ,
         \SB1_4_17/Component_Function_0/NAND4_in[3] ,
         \SB1_4_17/Component_Function_0/NAND4_in[2] ,
         \SB1_4_17/Component_Function_0/NAND4_in[1] ,
         \SB1_4_17/Component_Function_0/NAND4_in[0] ,
         \SB1_4_17/Component_Function_1/NAND4_in[2] ,
         \SB1_4_17/Component_Function_1/NAND4_in[1] ,
         \SB1_4_17/Component_Function_1/NAND4_in[0] ,
         \SB1_4_17/Component_Function_5/NAND4_in[1] ,
         \SB1_4_18/Component_Function_0/NAND4_in[3] ,
         \SB1_4_18/Component_Function_0/NAND4_in[2] ,
         \SB1_4_18/Component_Function_0/NAND4_in[1] ,
         \SB1_4_18/Component_Function_0/NAND4_in[0] ,
         \SB1_4_18/Component_Function_1/NAND4_in[3] ,
         \SB1_4_18/Component_Function_1/NAND4_in[2] ,
         \SB1_4_18/Component_Function_1/NAND4_in[1] ,
         \SB1_4_18/Component_Function_1/NAND4_in[0] ,
         \SB1_4_18/Component_Function_5/NAND4_in[2] ,
         \SB1_4_18/Component_Function_5/NAND4_in[0] ,
         \SB1_4_19/Component_Function_0/NAND4_in[3] ,
         \SB1_4_19/Component_Function_0/NAND4_in[2] ,
         \SB1_4_19/Component_Function_0/NAND4_in[1] ,
         \SB1_4_19/Component_Function_0/NAND4_in[0] ,
         \SB1_4_19/Component_Function_1/NAND4_in[3] ,
         \SB1_4_19/Component_Function_1/NAND4_in[2] ,
         \SB1_4_19/Component_Function_1/NAND4_in[1] ,
         \SB1_4_19/Component_Function_1/NAND4_in[0] ,
         \SB1_4_19/Component_Function_5/NAND4_in[1] ,
         \SB1_4_20/Component_Function_0/NAND4_in[3] ,
         \SB1_4_20/Component_Function_0/NAND4_in[2] ,
         \SB1_4_20/Component_Function_0/NAND4_in[1] ,
         \SB1_4_20/Component_Function_0/NAND4_in[0] ,
         \SB1_4_20/Component_Function_1/NAND4_in[2] ,
         \SB1_4_20/Component_Function_1/NAND4_in[1] ,
         \SB1_4_20/Component_Function_1/NAND4_in[0] ,
         \SB1_4_20/Component_Function_5/NAND4_in[1] ,
         \SB1_4_21/Component_Function_0/NAND4_in[3] ,
         \SB1_4_21/Component_Function_0/NAND4_in[2] ,
         \SB1_4_21/Component_Function_0/NAND4_in[1] ,
         \SB1_4_21/Component_Function_0/NAND4_in[0] ,
         \SB1_4_21/Component_Function_1/NAND4_in[3] ,
         \SB1_4_21/Component_Function_1/NAND4_in[1] ,
         \SB1_4_21/Component_Function_1/NAND4_in[0] ,
         \SB1_4_21/Component_Function_5/NAND4_in[1] ,
         \SB1_4_22/Component_Function_0/NAND4_in[2] ,
         \SB1_4_22/Component_Function_0/NAND4_in[1] ,
         \SB1_4_22/Component_Function_0/NAND4_in[0] ,
         \SB1_4_22/Component_Function_1/NAND4_in[3] ,
         \SB1_4_22/Component_Function_1/NAND4_in[2] ,
         \SB1_4_22/Component_Function_1/NAND4_in[1] ,
         \SB1_4_22/Component_Function_1/NAND4_in[0] ,
         \SB1_4_22/Component_Function_5/NAND4_in[3] ,
         \SB1_4_22/Component_Function_5/NAND4_in[1] ,
         \SB1_4_23/Component_Function_0/NAND4_in[2] ,
         \SB1_4_23/Component_Function_0/NAND4_in[1] ,
         \SB1_4_23/Component_Function_0/NAND4_in[0] ,
         \SB1_4_23/Component_Function_1/NAND4_in[1] ,
         \SB1_4_23/Component_Function_1/NAND4_in[0] ,
         \SB1_4_23/Component_Function_5/NAND4_in[2] ,
         \SB1_4_23/Component_Function_5/NAND4_in[1] ,
         \SB1_4_23/Component_Function_5/NAND4_in[0] ,
         \SB1_4_24/Component_Function_0/NAND4_in[2] ,
         \SB1_4_24/Component_Function_0/NAND4_in[1] ,
         \SB1_4_24/Component_Function_0/NAND4_in[0] ,
         \SB1_4_24/Component_Function_1/NAND4_in[3] ,
         \SB1_4_24/Component_Function_1/NAND4_in[2] ,
         \SB1_4_24/Component_Function_1/NAND4_in[1] ,
         \SB1_4_24/Component_Function_1/NAND4_in[0] ,
         \SB1_4_24/Component_Function_5/NAND4_in[1] ,
         \SB1_4_24/Component_Function_5/NAND4_in[0] ,
         \SB1_4_25/Component_Function_0/NAND4_in[2] ,
         \SB1_4_25/Component_Function_0/NAND4_in[0] ,
         \SB1_4_25/Component_Function_1/NAND4_in[3] ,
         \SB1_4_25/Component_Function_1/NAND4_in[1] ,
         \SB1_4_25/Component_Function_1/NAND4_in[0] ,
         \SB1_4_25/Component_Function_5/NAND4_in[3] ,
         \SB1_4_25/Component_Function_5/NAND4_in[1] ,
         \SB1_4_25/Component_Function_5/NAND4_in[0] ,
         \SB1_4_26/Component_Function_0/NAND4_in[3] ,
         \SB1_4_26/Component_Function_0/NAND4_in[2] ,
         \SB1_4_26/Component_Function_0/NAND4_in[1] ,
         \SB1_4_26/Component_Function_0/NAND4_in[0] ,
         \SB1_4_26/Component_Function_1/NAND4_in[3] ,
         \SB1_4_26/Component_Function_1/NAND4_in[2] ,
         \SB1_4_26/Component_Function_1/NAND4_in[1] ,
         \SB1_4_26/Component_Function_1/NAND4_in[0] ,
         \SB1_4_26/Component_Function_5/NAND4_in[2] ,
         \SB1_4_26/Component_Function_5/NAND4_in[0] ,
         \SB1_4_27/Component_Function_0/NAND4_in[3] ,
         \SB1_4_27/Component_Function_0/NAND4_in[2] ,
         \SB1_4_27/Component_Function_0/NAND4_in[1] ,
         \SB1_4_27/Component_Function_1/NAND4_in[3] ,
         \SB1_4_27/Component_Function_1/NAND4_in[2] ,
         \SB1_4_27/Component_Function_1/NAND4_in[1] ,
         \SB1_4_27/Component_Function_1/NAND4_in[0] ,
         \SB1_4_27/Component_Function_5/NAND4_in[3] ,
         \SB1_4_27/Component_Function_5/NAND4_in[2] ,
         \SB1_4_27/Component_Function_5/NAND4_in[1] ,
         \SB1_4_28/Component_Function_0/NAND4_in[2] ,
         \SB1_4_28/Component_Function_0/NAND4_in[0] ,
         \SB1_4_28/Component_Function_1/NAND4_in[3] ,
         \SB1_4_28/Component_Function_1/NAND4_in[1] ,
         \SB1_4_28/Component_Function_1/NAND4_in[0] ,
         \SB1_4_28/Component_Function_5/NAND4_in[2] ,
         \SB1_4_28/Component_Function_5/NAND4_in[1] ,
         \SB1_4_29/Component_Function_0/NAND4_in[2] ,
         \SB1_4_29/Component_Function_0/NAND4_in[1] ,
         \SB1_4_29/Component_Function_0/NAND4_in[0] ,
         \SB1_4_29/Component_Function_1/NAND4_in[3] ,
         \SB1_4_29/Component_Function_1/NAND4_in[2] ,
         \SB1_4_29/Component_Function_1/NAND4_in[0] ,
         \SB1_4_29/Component_Function_5/NAND4_in[0] ,
         \SB1_4_30/Component_Function_0/NAND4_in[2] ,
         \SB1_4_30/Component_Function_0/NAND4_in[1] ,
         \SB1_4_30/Component_Function_0/NAND4_in[0] ,
         \SB1_4_30/Component_Function_1/NAND4_in[3] ,
         \SB1_4_30/Component_Function_1/NAND4_in[2] ,
         \SB1_4_30/Component_Function_1/NAND4_in[1] ,
         \SB1_4_30/Component_Function_1/NAND4_in[0] ,
         \SB1_4_30/Component_Function_5/NAND4_in[3] ,
         \SB1_4_30/Component_Function_5/NAND4_in[2] ,
         \SB1_4_30/Component_Function_5/NAND4_in[1] ,
         \SB1_4_31/Component_Function_0/NAND4_in[2] ,
         \SB1_4_31/Component_Function_0/NAND4_in[1] ,
         \SB1_4_31/Component_Function_0/NAND4_in[0] ,
         \SB1_4_31/Component_Function_1/NAND4_in[3] ,
         \SB1_4_31/Component_Function_1/NAND4_in[1] ,
         \SB1_4_31/Component_Function_1/NAND4_in[0] ,
         \SB1_4_31/Component_Function_5/NAND4_in[3] ,
         \SB1_4_31/Component_Function_5/NAND4_in[2] ,
         \SB1_4_31/Component_Function_5/NAND4_in[1] ,
         \SB1_4_31/Component_Function_5/NAND4_in[0] ,
         \SB2_4_0/Component_Function_0/NAND4_in[3] ,
         \SB2_4_0/Component_Function_0/NAND4_in[2] ,
         \SB2_4_0/Component_Function_0/NAND4_in[1] ,
         \SB2_4_0/Component_Function_0/NAND4_in[0] ,
         \SB2_4_0/Component_Function_1/NAND4_in[3] ,
         \SB2_4_0/Component_Function_1/NAND4_in[2] ,
         \SB2_4_0/Component_Function_1/NAND4_in[1] ,
         \SB2_4_0/Component_Function_1/NAND4_in[0] ,
         \SB2_4_0/Component_Function_5/NAND4_in[2] ,
         \SB2_4_1/Component_Function_0/NAND4_in[3] ,
         \SB2_4_1/Component_Function_0/NAND4_in[2] ,
         \SB2_4_1/Component_Function_0/NAND4_in[0] ,
         \SB2_4_1/Component_Function_1/NAND4_in[2] ,
         \SB2_4_1/Component_Function_1/NAND4_in[1] ,
         \SB2_4_1/Component_Function_1/NAND4_in[0] ,
         \SB2_4_1/Component_Function_5/NAND4_in[3] ,
         \SB2_4_1/Component_Function_5/NAND4_in[2] ,
         \SB2_4_1/Component_Function_5/NAND4_in[1] ,
         \SB2_4_1/Component_Function_5/NAND4_in[0] ,
         \SB2_4_2/Component_Function_0/NAND4_in[3] ,
         \SB2_4_2/Component_Function_0/NAND4_in[2] ,
         \SB2_4_2/Component_Function_0/NAND4_in[1] ,
         \SB2_4_2/Component_Function_0/NAND4_in[0] ,
         \SB2_4_2/Component_Function_1/NAND4_in[3] ,
         \SB2_4_2/Component_Function_1/NAND4_in[1] ,
         \SB2_4_2/Component_Function_1/NAND4_in[0] ,
         \SB2_4_2/Component_Function_5/NAND4_in[1] ,
         \SB2_4_2/Component_Function_5/NAND4_in[0] ,
         \SB2_4_3/Component_Function_0/NAND4_in[2] ,
         \SB2_4_3/Component_Function_0/NAND4_in[1] ,
         \SB2_4_3/Component_Function_0/NAND4_in[0] ,
         \SB2_4_3/Component_Function_1/NAND4_in[3] ,
         \SB2_4_3/Component_Function_1/NAND4_in[2] ,
         \SB2_4_3/Component_Function_1/NAND4_in[1] ,
         \SB2_4_3/Component_Function_1/NAND4_in[0] ,
         \SB2_4_3/Component_Function_5/NAND4_in[3] ,
         \SB2_4_3/Component_Function_5/NAND4_in[1] ,
         \SB2_4_3/Component_Function_5/NAND4_in[0] ,
         \SB2_4_4/Component_Function_0/NAND4_in[3] ,
         \SB2_4_4/Component_Function_0/NAND4_in[1] ,
         \SB2_4_4/Component_Function_0/NAND4_in[0] ,
         \SB2_4_4/Component_Function_1/NAND4_in[3] ,
         \SB2_4_4/Component_Function_1/NAND4_in[2] ,
         \SB2_4_4/Component_Function_1/NAND4_in[1] ,
         \SB2_4_4/Component_Function_1/NAND4_in[0] ,
         \SB2_4_4/Component_Function_5/NAND4_in[1] ,
         \SB2_4_4/Component_Function_5/NAND4_in[0] ,
         \SB2_4_5/Component_Function_0/NAND4_in[2] ,
         \SB2_4_5/Component_Function_0/NAND4_in[1] ,
         \SB2_4_5/Component_Function_0/NAND4_in[0] ,
         \SB2_4_5/Component_Function_1/NAND4_in[3] ,
         \SB2_4_5/Component_Function_1/NAND4_in[2] ,
         \SB2_4_5/Component_Function_1/NAND4_in[1] ,
         \SB2_4_5/Component_Function_1/NAND4_in[0] ,
         \SB2_4_5/Component_Function_5/NAND4_in[2] ,
         \SB2_4_5/Component_Function_5/NAND4_in[0] ,
         \SB2_4_6/Component_Function_0/NAND4_in[2] ,
         \SB2_4_6/Component_Function_0/NAND4_in[1] ,
         \SB2_4_6/Component_Function_0/NAND4_in[0] ,
         \SB2_4_6/Component_Function_1/NAND4_in[3] ,
         \SB2_4_6/Component_Function_1/NAND4_in[2] ,
         \SB2_4_6/Component_Function_1/NAND4_in[1] ,
         \SB2_4_6/Component_Function_1/NAND4_in[0] ,
         \SB2_4_6/Component_Function_5/NAND4_in[0] ,
         \SB2_4_7/Component_Function_0/NAND4_in[2] ,
         \SB2_4_7/Component_Function_0/NAND4_in[0] ,
         \SB2_4_7/Component_Function_1/NAND4_in[3] ,
         \SB2_4_7/Component_Function_1/NAND4_in[2] ,
         \SB2_4_7/Component_Function_1/NAND4_in[1] ,
         \SB2_4_7/Component_Function_1/NAND4_in[0] ,
         \SB2_4_7/Component_Function_5/NAND4_in[0] ,
         \SB2_4_8/Component_Function_0/NAND4_in[3] ,
         \SB2_4_8/Component_Function_0/NAND4_in[2] ,
         \SB2_4_8/Component_Function_0/NAND4_in[0] ,
         \SB2_4_8/Component_Function_1/NAND4_in[3] ,
         \SB2_4_8/Component_Function_1/NAND4_in[2] ,
         \SB2_4_8/Component_Function_1/NAND4_in[1] ,
         \SB2_4_8/Component_Function_1/NAND4_in[0] ,
         \SB2_4_8/Component_Function_5/NAND4_in[2] ,
         \SB2_4_9/Component_Function_0/NAND4_in[2] ,
         \SB2_4_9/Component_Function_0/NAND4_in[1] ,
         \SB2_4_9/Component_Function_0/NAND4_in[0] ,
         \SB2_4_9/Component_Function_1/NAND4_in[3] ,
         \SB2_4_9/Component_Function_1/NAND4_in[1] ,
         \SB2_4_9/Component_Function_1/NAND4_in[0] ,
         \SB2_4_9/Component_Function_5/NAND4_in[1] ,
         \SB2_4_10/Component_Function_0/NAND4_in[3] ,
         \SB2_4_10/Component_Function_0/NAND4_in[2] ,
         \SB2_4_10/Component_Function_0/NAND4_in[1] ,
         \SB2_4_10/Component_Function_0/NAND4_in[0] ,
         \SB2_4_10/Component_Function_1/NAND4_in[3] ,
         \SB2_4_10/Component_Function_1/NAND4_in[2] ,
         \SB2_4_10/Component_Function_1/NAND4_in[1] ,
         \SB2_4_10/Component_Function_1/NAND4_in[0] ,
         \SB2_4_10/Component_Function_5/NAND4_in[2] ,
         \SB2_4_11/Component_Function_0/NAND4_in[2] ,
         \SB2_4_11/Component_Function_0/NAND4_in[1] ,
         \SB2_4_11/Component_Function_0/NAND4_in[0] ,
         \SB2_4_11/Component_Function_1/NAND4_in[1] ,
         \SB2_4_11/Component_Function_1/NAND4_in[0] ,
         \SB2_4_12/Component_Function_0/NAND4_in[3] ,
         \SB2_4_12/Component_Function_0/NAND4_in[2] ,
         \SB2_4_12/Component_Function_0/NAND4_in[0] ,
         \SB2_4_12/Component_Function_1/NAND4_in[3] ,
         \SB2_4_12/Component_Function_1/NAND4_in[2] ,
         \SB2_4_12/Component_Function_1/NAND4_in[1] ,
         \SB2_4_12/Component_Function_1/NAND4_in[0] ,
         \SB2_4_13/Component_Function_0/NAND4_in[3] ,
         \SB2_4_13/Component_Function_0/NAND4_in[1] ,
         \SB2_4_13/Component_Function_0/NAND4_in[0] ,
         \SB2_4_13/Component_Function_1/NAND4_in[2] ,
         \SB2_4_13/Component_Function_1/NAND4_in[1] ,
         \SB2_4_13/Component_Function_1/NAND4_in[0] ,
         \SB2_4_13/Component_Function_5/NAND4_in[0] ,
         \SB2_4_14/Component_Function_0/NAND4_in[2] ,
         \SB2_4_14/Component_Function_0/NAND4_in[1] ,
         \SB2_4_14/Component_Function_1/NAND4_in[3] ,
         \SB2_4_14/Component_Function_1/NAND4_in[2] ,
         \SB2_4_14/Component_Function_1/NAND4_in[1] ,
         \SB2_4_14/Component_Function_5/NAND4_in[0] ,
         \SB2_4_15/Component_Function_0/NAND4_in[2] ,
         \SB2_4_15/Component_Function_0/NAND4_in[1] ,
         \SB2_4_15/Component_Function_0/NAND4_in[0] ,
         \SB2_4_15/Component_Function_1/NAND4_in[3] ,
         \SB2_4_15/Component_Function_1/NAND4_in[2] ,
         \SB2_4_15/Component_Function_1/NAND4_in[1] ,
         \SB2_4_15/Component_Function_1/NAND4_in[0] ,
         \SB2_4_15/Component_Function_5/NAND4_in[3] ,
         \SB2_4_16/Component_Function_0/NAND4_in[2] ,
         \SB2_4_16/Component_Function_0/NAND4_in[1] ,
         \SB2_4_16/Component_Function_0/NAND4_in[0] ,
         \SB2_4_16/Component_Function_1/NAND4_in[3] ,
         \SB2_4_16/Component_Function_1/NAND4_in[2] ,
         \SB2_4_16/Component_Function_1/NAND4_in[1] ,
         \SB2_4_16/Component_Function_1/NAND4_in[0] ,
         \SB2_4_17/Component_Function_0/NAND4_in[3] ,
         \SB2_4_17/Component_Function_0/NAND4_in[2] ,
         \SB2_4_17/Component_Function_0/NAND4_in[1] ,
         \SB2_4_17/Component_Function_0/NAND4_in[0] ,
         \SB2_4_17/Component_Function_1/NAND4_in[3] ,
         \SB2_4_17/Component_Function_1/NAND4_in[2] ,
         \SB2_4_17/Component_Function_1/NAND4_in[1] ,
         \SB2_4_17/Component_Function_1/NAND4_in[0] ,
         \SB2_4_17/Component_Function_5/NAND4_in[2] ,
         \SB2_4_18/Component_Function_0/NAND4_in[3] ,
         \SB2_4_18/Component_Function_0/NAND4_in[1] ,
         \SB2_4_18/Component_Function_0/NAND4_in[0] ,
         \SB2_4_18/Component_Function_1/NAND4_in[2] ,
         \SB2_4_18/Component_Function_1/NAND4_in[1] ,
         \SB2_4_18/Component_Function_5/NAND4_in[0] ,
         \SB2_4_19/Component_Function_0/NAND4_in[2] ,
         \SB2_4_19/Component_Function_0/NAND4_in[1] ,
         \SB2_4_19/Component_Function_0/NAND4_in[0] ,
         \SB2_4_19/Component_Function_1/NAND4_in[3] ,
         \SB2_4_19/Component_Function_1/NAND4_in[2] ,
         \SB2_4_19/Component_Function_1/NAND4_in[1] ,
         \SB2_4_19/Component_Function_1/NAND4_in[0] ,
         \SB2_4_19/Component_Function_5/NAND4_in[2] ,
         \SB2_4_19/Component_Function_5/NAND4_in[1] ,
         \SB2_4_19/Component_Function_5/NAND4_in[0] ,
         \SB2_4_20/Component_Function_0/NAND4_in[3] ,
         \SB2_4_20/Component_Function_0/NAND4_in[1] ,
         \SB2_4_20/Component_Function_0/NAND4_in[0] ,
         \SB2_4_20/Component_Function_1/NAND4_in[3] ,
         \SB2_4_20/Component_Function_1/NAND4_in[2] ,
         \SB2_4_20/Component_Function_1/NAND4_in[1] ,
         \SB2_4_20/Component_Function_1/NAND4_in[0] ,
         \SB2_4_20/Component_Function_5/NAND4_in[1] ,
         \SB2_4_20/Component_Function_5/NAND4_in[0] ,
         \SB2_4_21/Component_Function_0/NAND4_in[2] ,
         \SB2_4_21/Component_Function_0/NAND4_in[1] ,
         \SB2_4_21/Component_Function_0/NAND4_in[0] ,
         \SB2_4_21/Component_Function_1/NAND4_in[3] ,
         \SB2_4_21/Component_Function_1/NAND4_in[1] ,
         \SB2_4_21/Component_Function_1/NAND4_in[0] ,
         \SB2_4_21/Component_Function_5/NAND4_in[2] ,
         \SB2_4_21/Component_Function_5/NAND4_in[1] ,
         \SB2_4_21/Component_Function_5/NAND4_in[0] ,
         \SB2_4_22/Component_Function_0/NAND4_in[3] ,
         \SB2_4_22/Component_Function_0/NAND4_in[1] ,
         \SB2_4_22/Component_Function_0/NAND4_in[0] ,
         \SB2_4_22/Component_Function_1/NAND4_in[3] ,
         \SB2_4_22/Component_Function_1/NAND4_in[1] ,
         \SB2_4_22/Component_Function_1/NAND4_in[0] ,
         \SB2_4_22/Component_Function_5/NAND4_in[3] ,
         \SB2_4_22/Component_Function_5/NAND4_in[2] ,
         \SB2_4_22/Component_Function_5/NAND4_in[1] ,
         \SB2_4_22/Component_Function_5/NAND4_in[0] ,
         \SB2_4_23/Component_Function_0/NAND4_in[2] ,
         \SB2_4_23/Component_Function_0/NAND4_in[1] ,
         \SB2_4_23/Component_Function_0/NAND4_in[0] ,
         \SB2_4_23/Component_Function_1/NAND4_in[2] ,
         \SB2_4_23/Component_Function_1/NAND4_in[1] ,
         \SB2_4_23/Component_Function_1/NAND4_in[0] ,
         \SB2_4_23/Component_Function_5/NAND4_in[1] ,
         \SB2_4_23/Component_Function_5/NAND4_in[0] ,
         \SB2_4_24/Component_Function_0/NAND4_in[3] ,
         \SB2_4_24/Component_Function_0/NAND4_in[1] ,
         \SB2_4_24/Component_Function_0/NAND4_in[0] ,
         \SB2_4_24/Component_Function_1/NAND4_in[3] ,
         \SB2_4_24/Component_Function_1/NAND4_in[2] ,
         \SB2_4_24/Component_Function_1/NAND4_in[1] ,
         \SB2_4_24/Component_Function_1/NAND4_in[0] ,
         \SB2_4_24/Component_Function_5/NAND4_in[2] ,
         \SB2_4_24/Component_Function_5/NAND4_in[0] ,
         \SB2_4_25/Component_Function_0/NAND4_in[1] ,
         \SB2_4_25/Component_Function_0/NAND4_in[0] ,
         \SB2_4_25/Component_Function_1/NAND4_in[2] ,
         \SB2_4_25/Component_Function_1/NAND4_in[1] ,
         \SB2_4_25/Component_Function_1/NAND4_in[0] ,
         \SB2_4_26/Component_Function_0/NAND4_in[2] ,
         \SB2_4_26/Component_Function_0/NAND4_in[1] ,
         \SB2_4_26/Component_Function_0/NAND4_in[0] ,
         \SB2_4_26/Component_Function_1/NAND4_in[2] ,
         \SB2_4_26/Component_Function_1/NAND4_in[1] ,
         \SB2_4_26/Component_Function_1/NAND4_in[0] ,
         \SB2_4_26/Component_Function_5/NAND4_in[1] ,
         \SB2_4_26/Component_Function_5/NAND4_in[0] ,
         \SB2_4_27/Component_Function_0/NAND4_in[2] ,
         \SB2_4_27/Component_Function_0/NAND4_in[1] ,
         \SB2_4_27/Component_Function_0/NAND4_in[0] ,
         \SB2_4_27/Component_Function_1/NAND4_in[2] ,
         \SB2_4_27/Component_Function_1/NAND4_in[1] ,
         \SB2_4_27/Component_Function_1/NAND4_in[0] ,
         \SB2_4_27/Component_Function_5/NAND4_in[0] ,
         \SB2_4_28/Component_Function_0/NAND4_in[3] ,
         \SB2_4_28/Component_Function_0/NAND4_in[1] ,
         \SB2_4_28/Component_Function_0/NAND4_in[0] ,
         \SB2_4_28/Component_Function_1/NAND4_in[3] ,
         \SB2_4_28/Component_Function_1/NAND4_in[2] ,
         \SB2_4_28/Component_Function_1/NAND4_in[1] ,
         \SB2_4_28/Component_Function_1/NAND4_in[0] ,
         \SB2_4_28/Component_Function_5/NAND4_in[0] ,
         \SB2_4_29/Component_Function_0/NAND4_in[2] ,
         \SB2_4_29/Component_Function_0/NAND4_in[1] ,
         \SB2_4_29/Component_Function_0/NAND4_in[0] ,
         \SB2_4_29/Component_Function_1/NAND4_in[2] ,
         \SB2_4_29/Component_Function_1/NAND4_in[1] ,
         \SB2_4_29/Component_Function_1/NAND4_in[0] ,
         \SB2_4_29/Component_Function_5/NAND4_in[3] ,
         \SB2_4_29/Component_Function_5/NAND4_in[0] ,
         \SB2_4_30/Component_Function_0/NAND4_in[3] ,
         \SB2_4_30/Component_Function_0/NAND4_in[2] ,
         \SB2_4_30/Component_Function_0/NAND4_in[1] ,
         \SB2_4_30/Component_Function_0/NAND4_in[0] ,
         \SB2_4_30/Component_Function_1/NAND4_in[2] ,
         \SB2_4_30/Component_Function_1/NAND4_in[1] ,
         \SB2_4_30/Component_Function_1/NAND4_in[0] ,
         \SB2_4_30/Component_Function_5/NAND4_in[2] ,
         \SB2_4_30/Component_Function_5/NAND4_in[1] ,
         \SB2_4_30/Component_Function_5/NAND4_in[0] ,
         \SB2_4_31/Component_Function_0/NAND4_in[2] ,
         \SB2_4_31/Component_Function_0/NAND4_in[1] ,
         \SB2_4_31/Component_Function_0/NAND4_in[0] ,
         \SB2_4_31/Component_Function_1/NAND4_in[3] ,
         \SB2_4_31/Component_Function_1/NAND4_in[2] ,
         \SB2_4_31/Component_Function_1/NAND4_in[1] ,
         \SB2_4_31/Component_Function_1/NAND4_in[0] ,
         \SB2_4_31/Component_Function_5/NAND4_in[1] ,
         \SB2_4_31/Component_Function_5/NAND4_in[0] ,
         \SB3_0/Component_Function_0/NAND4_in[3] ,
         \SB3_0/Component_Function_0/NAND4_in[2] ,
         \SB3_0/Component_Function_0/NAND4_in[1] ,
         \SB3_0/Component_Function_0/NAND4_in[0] ,
         \SB3_0/Component_Function_1/NAND4_in[2] ,
         \SB3_0/Component_Function_1/NAND4_in[1] ,
         \SB3_0/Component_Function_5/NAND4_in[1] ,
         \SB3_0/Component_Function_5/NAND4_in[0] ,
         \SB3_1/Component_Function_0/NAND4_in[1] ,
         \SB3_1/Component_Function_0/NAND4_in[0] ,
         \SB3_1/Component_Function_1/NAND4_in[2] ,
         \SB3_1/Component_Function_1/NAND4_in[1] ,
         \SB3_1/Component_Function_1/NAND4_in[0] ,
         \SB3_1/Component_Function_5/NAND4_in[2] ,
         \SB3_1/Component_Function_5/NAND4_in[1] ,
         \SB3_1/Component_Function_5/NAND4_in[0] ,
         \SB3_2/Component_Function_0/NAND4_in[2] ,
         \SB3_2/Component_Function_0/NAND4_in[1] ,
         \SB3_2/Component_Function_0/NAND4_in[0] ,
         \SB3_2/Component_Function_1/NAND4_in[3] ,
         \SB3_2/Component_Function_1/NAND4_in[1] ,
         \SB3_2/Component_Function_5/NAND4_in[1] ,
         \SB3_2/Component_Function_5/NAND4_in[0] ,
         \SB3_3/Component_Function_0/NAND4_in[2] ,
         \SB3_3/Component_Function_0/NAND4_in[1] ,
         \SB3_3/Component_Function_0/NAND4_in[0] ,
         \SB3_3/Component_Function_1/NAND4_in[3] ,
         \SB3_3/Component_Function_1/NAND4_in[2] ,
         \SB3_3/Component_Function_1/NAND4_in[1] ,
         \SB3_3/Component_Function_1/NAND4_in[0] ,
         \SB3_3/Component_Function_5/NAND4_in[3] ,
         \SB3_3/Component_Function_5/NAND4_in[1] ,
         \SB3_3/Component_Function_5/NAND4_in[0] ,
         \SB3_4/Component_Function_0/NAND4_in[3] ,
         \SB3_4/Component_Function_0/NAND4_in[2] ,
         \SB3_4/Component_Function_0/NAND4_in[1] ,
         \SB3_4/Component_Function_0/NAND4_in[0] ,
         \SB3_4/Component_Function_1/NAND4_in[3] ,
         \SB3_4/Component_Function_1/NAND4_in[2] ,
         \SB3_4/Component_Function_1/NAND4_in[1] ,
         \SB3_4/Component_Function_1/NAND4_in[0] ,
         \SB3_4/Component_Function_5/NAND4_in[3] ,
         \SB3_4/Component_Function_5/NAND4_in[1] ,
         \SB3_4/Component_Function_5/NAND4_in[0] ,
         \SB3_5/Component_Function_0/NAND4_in[2] ,
         \SB3_5/Component_Function_0/NAND4_in[1] ,
         \SB3_5/Component_Function_0/NAND4_in[0] ,
         \SB3_5/Component_Function_1/NAND4_in[3] ,
         \SB3_5/Component_Function_1/NAND4_in[2] ,
         \SB3_5/Component_Function_1/NAND4_in[1] ,
         \SB3_5/Component_Function_1/NAND4_in[0] ,
         \SB3_5/Component_Function_5/NAND4_in[3] ,
         \SB3_5/Component_Function_5/NAND4_in[2] ,
         \SB3_5/Component_Function_5/NAND4_in[1] ,
         \SB3_5/Component_Function_5/NAND4_in[0] ,
         \SB3_6/Component_Function_0/NAND4_in[3] ,
         \SB3_6/Component_Function_0/NAND4_in[2] ,
         \SB3_6/Component_Function_0/NAND4_in[1] ,
         \SB3_6/Component_Function_0/NAND4_in[0] ,
         \SB3_6/Component_Function_1/NAND4_in[3] ,
         \SB3_6/Component_Function_1/NAND4_in[2] ,
         \SB3_6/Component_Function_1/NAND4_in[1] ,
         \SB3_6/Component_Function_1/NAND4_in[0] ,
         \SB3_6/Component_Function_5/NAND4_in[2] ,
         \SB3_6/Component_Function_5/NAND4_in[1] ,
         \SB3_6/Component_Function_5/NAND4_in[0] ,
         \SB3_7/Component_Function_0/NAND4_in[3] ,
         \SB3_7/Component_Function_0/NAND4_in[2] ,
         \SB3_7/Component_Function_0/NAND4_in[0] ,
         \SB3_7/Component_Function_1/NAND4_in[3] ,
         \SB3_7/Component_Function_1/NAND4_in[2] ,
         \SB3_7/Component_Function_1/NAND4_in[1] ,
         \SB3_7/Component_Function_1/NAND4_in[0] ,
         \SB3_7/Component_Function_5/NAND4_in[3] ,
         \SB3_7/Component_Function_5/NAND4_in[2] ,
         \SB3_7/Component_Function_5/NAND4_in[0] ,
         \SB3_8/Component_Function_0/NAND4_in[3] ,
         \SB3_8/Component_Function_0/NAND4_in[2] ,
         \SB3_8/Component_Function_0/NAND4_in[1] ,
         \SB3_8/Component_Function_0/NAND4_in[0] ,
         \SB3_8/Component_Function_1/NAND4_in[3] ,
         \SB3_8/Component_Function_1/NAND4_in[2] ,
         \SB3_8/Component_Function_1/NAND4_in[1] ,
         \SB3_8/Component_Function_1/NAND4_in[0] ,
         \SB3_8/Component_Function_5/NAND4_in[2] ,
         \SB3_8/Component_Function_5/NAND4_in[1] ,
         \SB3_9/Component_Function_0/NAND4_in[3] ,
         \SB3_9/Component_Function_0/NAND4_in[2] ,
         \SB3_9/Component_Function_0/NAND4_in[1] ,
         \SB3_9/Component_Function_0/NAND4_in[0] ,
         \SB3_9/Component_Function_1/NAND4_in[2] ,
         \SB3_9/Component_Function_1/NAND4_in[1] ,
         \SB3_9/Component_Function_1/NAND4_in[0] ,
         \SB3_9/Component_Function_5/NAND4_in[1] ,
         \SB3_9/Component_Function_5/NAND4_in[0] ,
         \SB3_10/Component_Function_0/NAND4_in[3] ,
         \SB3_10/Component_Function_0/NAND4_in[2] ,
         \SB3_10/Component_Function_0/NAND4_in[1] ,
         \SB3_10/Component_Function_0/NAND4_in[0] ,
         \SB3_10/Component_Function_1/NAND4_in[3] ,
         \SB3_10/Component_Function_1/NAND4_in[2] ,
         \SB3_10/Component_Function_1/NAND4_in[1] ,
         \SB3_10/Component_Function_1/NAND4_in[0] ,
         \SB3_10/Component_Function_5/NAND4_in[1] ,
         \SB3_10/Component_Function_5/NAND4_in[0] ,
         \SB3_11/Component_Function_0/NAND4_in[2] ,
         \SB3_11/Component_Function_0/NAND4_in[1] ,
         \SB3_11/Component_Function_0/NAND4_in[0] ,
         \SB3_11/Component_Function_1/NAND4_in[3] ,
         \SB3_11/Component_Function_1/NAND4_in[2] ,
         \SB3_11/Component_Function_1/NAND4_in[1] ,
         \SB3_11/Component_Function_1/NAND4_in[0] ,
         \SB3_11/Component_Function_5/NAND4_in[2] ,
         \SB3_11/Component_Function_5/NAND4_in[1] ,
         \SB3_11/Component_Function_5/NAND4_in[0] ,
         \SB3_12/Component_Function_0/NAND4_in[1] ,
         \SB3_12/Component_Function_0/NAND4_in[0] ,
         \SB3_12/Component_Function_1/NAND4_in[3] ,
         \SB3_12/Component_Function_1/NAND4_in[2] ,
         \SB3_12/Component_Function_1/NAND4_in[1] ,
         \SB3_12/Component_Function_1/NAND4_in[0] ,
         \SB3_12/Component_Function_5/NAND4_in[2] ,
         \SB3_12/Component_Function_5/NAND4_in[1] ,
         \SB3_12/Component_Function_5/NAND4_in[0] ,
         \SB3_13/Component_Function_0/NAND4_in[2] ,
         \SB3_13/Component_Function_0/NAND4_in[1] ,
         \SB3_13/Component_Function_0/NAND4_in[0] ,
         \SB3_13/Component_Function_1/NAND4_in[2] ,
         \SB3_13/Component_Function_1/NAND4_in[1] ,
         \SB3_13/Component_Function_5/NAND4_in[2] ,
         \SB3_13/Component_Function_5/NAND4_in[1] ,
         \SB3_13/Component_Function_5/NAND4_in[0] ,
         \SB3_14/Component_Function_0/NAND4_in[2] ,
         \SB3_14/Component_Function_0/NAND4_in[1] ,
         \SB3_14/Component_Function_0/NAND4_in[0] ,
         \SB3_14/Component_Function_1/NAND4_in[2] ,
         \SB3_14/Component_Function_1/NAND4_in[1] ,
         \SB3_14/Component_Function_1/NAND4_in[0] ,
         \SB3_14/Component_Function_5/NAND4_in[2] ,
         \SB3_14/Component_Function_5/NAND4_in[1] ,
         \SB3_14/Component_Function_5/NAND4_in[0] ,
         \SB3_15/Component_Function_0/NAND4_in[2] ,
         \SB3_15/Component_Function_0/NAND4_in[1] ,
         \SB3_15/Component_Function_0/NAND4_in[0] ,
         \SB3_15/Component_Function_1/NAND4_in[2] ,
         \SB3_15/Component_Function_1/NAND4_in[1] ,
         \SB3_15/Component_Function_1/NAND4_in[0] ,
         \SB3_15/Component_Function_5/NAND4_in[2] ,
         \SB3_16/Component_Function_0/NAND4_in[3] ,
         \SB3_16/Component_Function_0/NAND4_in[1] ,
         \SB3_16/Component_Function_0/NAND4_in[0] ,
         \SB3_16/Component_Function_1/NAND4_in[3] ,
         \SB3_16/Component_Function_1/NAND4_in[2] ,
         \SB3_16/Component_Function_1/NAND4_in[1] ,
         \SB3_16/Component_Function_1/NAND4_in[0] ,
         \SB3_16/Component_Function_5/NAND4_in[3] ,
         \SB3_16/Component_Function_5/NAND4_in[1] ,
         \SB3_16/Component_Function_5/NAND4_in[0] ,
         \SB3_17/Component_Function_0/NAND4_in[2] ,
         \SB3_17/Component_Function_0/NAND4_in[1] ,
         \SB3_17/Component_Function_0/NAND4_in[0] ,
         \SB3_17/Component_Function_1/NAND4_in[2] ,
         \SB3_17/Component_Function_1/NAND4_in[1] ,
         \SB3_17/Component_Function_1/NAND4_in[0] ,
         \SB3_17/Component_Function_5/NAND4_in[1] ,
         \SB3_17/Component_Function_5/NAND4_in[0] ,
         \SB3_18/Component_Function_0/NAND4_in[3] ,
         \SB3_18/Component_Function_0/NAND4_in[2] ,
         \SB3_18/Component_Function_0/NAND4_in[1] ,
         \SB3_18/Component_Function_0/NAND4_in[0] ,
         \SB3_18/Component_Function_1/NAND4_in[3] ,
         \SB3_18/Component_Function_1/NAND4_in[2] ,
         \SB3_18/Component_Function_1/NAND4_in[1] ,
         \SB3_18/Component_Function_1/NAND4_in[0] ,
         \SB3_18/Component_Function_5/NAND4_in[3] ,
         \SB3_18/Component_Function_5/NAND4_in[2] ,
         \SB3_18/Component_Function_5/NAND4_in[1] ,
         \SB3_18/Component_Function_5/NAND4_in[0] ,
         \SB3_19/Component_Function_0/NAND4_in[2] ,
         \SB3_19/Component_Function_0/NAND4_in[1] ,
         \SB3_19/Component_Function_0/NAND4_in[0] ,
         \SB3_19/Component_Function_1/NAND4_in[2] ,
         \SB3_19/Component_Function_1/NAND4_in[1] ,
         \SB3_19/Component_Function_1/NAND4_in[0] ,
         \SB3_19/Component_Function_5/NAND4_in[1] ,
         \SB3_19/Component_Function_5/NAND4_in[0] ,
         \SB3_20/Component_Function_0/NAND4_in[3] ,
         \SB3_20/Component_Function_0/NAND4_in[2] ,
         \SB3_20/Component_Function_0/NAND4_in[1] ,
         \SB3_20/Component_Function_0/NAND4_in[0] ,
         \SB3_20/Component_Function_1/NAND4_in[1] ,
         \SB3_20/Component_Function_1/NAND4_in[0] ,
         \SB3_20/Component_Function_5/NAND4_in[1] ,
         \SB3_21/Component_Function_0/NAND4_in[2] ,
         \SB3_21/Component_Function_0/NAND4_in[1] ,
         \SB3_21/Component_Function_0/NAND4_in[0] ,
         \SB3_21/Component_Function_1/NAND4_in[2] ,
         \SB3_21/Component_Function_1/NAND4_in[1] ,
         \SB3_21/Component_Function_1/NAND4_in[0] ,
         \SB3_21/Component_Function_5/NAND4_in[1] ,
         \SB3_21/Component_Function_5/NAND4_in[0] ,
         \SB3_22/Component_Function_0/NAND4_in[3] ,
         \SB3_22/Component_Function_0/NAND4_in[2] ,
         \SB3_22/Component_Function_0/NAND4_in[1] ,
         \SB3_22/Component_Function_0/NAND4_in[0] ,
         \SB3_22/Component_Function_1/NAND4_in[3] ,
         \SB3_22/Component_Function_1/NAND4_in[2] ,
         \SB3_22/Component_Function_1/NAND4_in[1] ,
         \SB3_22/Component_Function_1/NAND4_in[0] ,
         \SB3_22/Component_Function_5/NAND4_in[2] ,
         \SB3_22/Component_Function_5/NAND4_in[1] ,
         \SB3_22/Component_Function_5/NAND4_in[0] ,
         \SB3_23/Component_Function_0/NAND4_in[3] ,
         \SB3_23/Component_Function_0/NAND4_in[2] ,
         \SB3_23/Component_Function_0/NAND4_in[0] ,
         \SB3_23/Component_Function_1/NAND4_in[3] ,
         \SB3_23/Component_Function_1/NAND4_in[2] ,
         \SB3_23/Component_Function_1/NAND4_in[1] ,
         \SB3_23/Component_Function_1/NAND4_in[0] ,
         \SB3_23/Component_Function_5/NAND4_in[3] ,
         \SB3_23/Component_Function_5/NAND4_in[2] ,
         \SB3_23/Component_Function_5/NAND4_in[1] ,
         \SB3_23/Component_Function_5/NAND4_in[0] ,
         \SB3_24/Component_Function_0/NAND4_in[3] ,
         \SB3_24/Component_Function_0/NAND4_in[2] ,
         \SB3_24/Component_Function_0/NAND4_in[1] ,
         \SB3_24/Component_Function_0/NAND4_in[0] ,
         \SB3_24/Component_Function_1/NAND4_in[2] ,
         \SB3_24/Component_Function_1/NAND4_in[1] ,
         \SB3_24/Component_Function_1/NAND4_in[0] ,
         \SB3_24/Component_Function_5/NAND4_in[3] ,
         \SB3_24/Component_Function_5/NAND4_in[1] ,
         \SB3_24/Component_Function_5/NAND4_in[0] ,
         \SB3_25/Component_Function_0/NAND4_in[2] ,
         \SB3_25/Component_Function_0/NAND4_in[1] ,
         \SB3_25/Component_Function_0/NAND4_in[0] ,
         \SB3_25/Component_Function_1/NAND4_in[3] ,
         \SB3_25/Component_Function_1/NAND4_in[2] ,
         \SB3_25/Component_Function_1/NAND4_in[1] ,
         \SB3_25/Component_Function_1/NAND4_in[0] ,
         \SB3_25/Component_Function_5/NAND4_in[2] ,
         \SB3_25/Component_Function_5/NAND4_in[1] ,
         \SB3_25/Component_Function_5/NAND4_in[0] ,
         \SB3_26/Component_Function_0/NAND4_in[1] ,
         \SB3_26/Component_Function_0/NAND4_in[0] ,
         \SB3_26/Component_Function_1/NAND4_in[3] ,
         \SB3_26/Component_Function_1/NAND4_in[2] ,
         \SB3_26/Component_Function_1/NAND4_in[1] ,
         \SB3_26/Component_Function_1/NAND4_in[0] ,
         \SB3_26/Component_Function_5/NAND4_in[1] ,
         \SB3_27/Component_Function_0/NAND4_in[3] ,
         \SB3_27/Component_Function_0/NAND4_in[2] ,
         \SB3_27/Component_Function_0/NAND4_in[1] ,
         \SB3_27/Component_Function_0/NAND4_in[0] ,
         \SB3_27/Component_Function_1/NAND4_in[3] ,
         \SB3_27/Component_Function_1/NAND4_in[1] ,
         \SB3_27/Component_Function_1/NAND4_in[0] ,
         \SB3_27/Component_Function_5/NAND4_in[3] ,
         \SB3_27/Component_Function_5/NAND4_in[1] ,
         \SB3_27/Component_Function_5/NAND4_in[0] ,
         \SB3_28/Component_Function_0/NAND4_in[3] ,
         \SB3_28/Component_Function_0/NAND4_in[2] ,
         \SB3_28/Component_Function_0/NAND4_in[1] ,
         \SB3_28/Component_Function_0/NAND4_in[0] ,
         \SB3_28/Component_Function_1/NAND4_in[3] ,
         \SB3_28/Component_Function_1/NAND4_in[1] ,
         \SB3_28/Component_Function_1/NAND4_in[0] ,
         \SB3_28/Component_Function_5/NAND4_in[1] ,
         \SB3_28/Component_Function_5/NAND4_in[0] ,
         \SB3_29/Component_Function_0/NAND4_in[3] ,
         \SB3_29/Component_Function_0/NAND4_in[2] ,
         \SB3_29/Component_Function_0/NAND4_in[1] ,
         \SB3_29/Component_Function_0/NAND4_in[0] ,
         \SB3_29/Component_Function_1/NAND4_in[3] ,
         \SB3_29/Component_Function_1/NAND4_in[2] ,
         \SB3_29/Component_Function_1/NAND4_in[1] ,
         \SB3_29/Component_Function_1/NAND4_in[0] ,
         \SB3_29/Component_Function_5/NAND4_in[3] ,
         \SB3_29/Component_Function_5/NAND4_in[2] ,
         \SB3_29/Component_Function_5/NAND4_in[1] ,
         \SB3_29/Component_Function_5/NAND4_in[0] ,
         \SB3_30/Component_Function_0/NAND4_in[3] ,
         \SB3_30/Component_Function_0/NAND4_in[1] ,
         \SB3_30/Component_Function_0/NAND4_in[0] ,
         \SB3_30/Component_Function_1/NAND4_in[3] ,
         \SB3_30/Component_Function_1/NAND4_in[1] ,
         \SB3_30/Component_Function_1/NAND4_in[0] ,
         \SB3_30/Component_Function_5/NAND4_in[1] ,
         \SB3_30/Component_Function_5/NAND4_in[0] ,
         \SB3_31/Component_Function_0/NAND4_in[3] ,
         \SB3_31/Component_Function_0/NAND4_in[2] ,
         \SB3_31/Component_Function_0/NAND4_in[1] ,
         \SB3_31/Component_Function_0/NAND4_in[0] ,
         \SB3_31/Component_Function_1/NAND4_in[3] ,
         \SB3_31/Component_Function_1/NAND4_in[2] ,
         \SB3_31/Component_Function_1/NAND4_in[1] ,
         \SB3_31/Component_Function_1/NAND4_in[0] ,
         \SB3_31/Component_Function_5/NAND4_in[2] ,
         \SB3_31/Component_Function_5/NAND4_in[0] ,
         \SB4_0/Component_Function_0/NAND4_in[2] ,
         \SB4_0/Component_Function_0/NAND4_in[1] ,
         \SB4_0/Component_Function_1/NAND4_in[1] ,
         \SB4_0/Component_Function_1/NAND4_in[0] ,
         \SB4_0/Component_Function_5/NAND4_in[3] ,
         \SB4_0/Component_Function_5/NAND4_in[2] ,
         \SB4_0/Component_Function_5/NAND4_in[0] ,
         \SB4_1/Component_Function_0/NAND4_in[3] ,
         \SB4_1/Component_Function_0/NAND4_in[2] ,
         \SB4_1/Component_Function_0/NAND4_in[1] ,
         \SB4_1/Component_Function_0/NAND4_in[0] ,
         \SB4_1/Component_Function_1/NAND4_in[2] ,
         \SB4_1/Component_Function_1/NAND4_in[1] ,
         \SB4_1/Component_Function_1/NAND4_in[0] ,
         \SB4_1/Component_Function_5/NAND4_in[3] ,
         \SB4_1/Component_Function_5/NAND4_in[1] ,
         \SB4_1/Component_Function_5/NAND4_in[0] ,
         \SB4_2/Component_Function_0/NAND4_in[3] ,
         \SB4_2/Component_Function_0/NAND4_in[1] ,
         \SB4_2/Component_Function_0/NAND4_in[0] ,
         \SB4_2/Component_Function_1/NAND4_in[3] ,
         \SB4_2/Component_Function_1/NAND4_in[2] ,
         \SB4_2/Component_Function_1/NAND4_in[1] ,
         \SB4_2/Component_Function_1/NAND4_in[0] ,
         \SB4_2/Component_Function_5/NAND4_in[3] ,
         \SB4_2/Component_Function_5/NAND4_in[2] ,
         \SB4_2/Component_Function_5/NAND4_in[0] ,
         \SB4_3/Component_Function_0/NAND4_in[3] ,
         \SB4_3/Component_Function_0/NAND4_in[2] ,
         \SB4_3/Component_Function_0/NAND4_in[1] ,
         \SB4_3/Component_Function_0/NAND4_in[0] ,
         \SB4_3/Component_Function_1/NAND4_in[3] ,
         \SB4_3/Component_Function_1/NAND4_in[2] ,
         \SB4_3/Component_Function_1/NAND4_in[1] ,
         \SB4_3/Component_Function_1/NAND4_in[0] ,
         \SB4_3/Component_Function_5/NAND4_in[3] ,
         \SB4_3/Component_Function_5/NAND4_in[2] ,
         \SB4_4/Component_Function_0/NAND4_in[2] ,
         \SB4_4/Component_Function_0/NAND4_in[1] ,
         \SB4_4/Component_Function_1/NAND4_in[3] ,
         \SB4_4/Component_Function_1/NAND4_in[2] ,
         \SB4_4/Component_Function_1/NAND4_in[1] ,
         \SB4_4/Component_Function_1/NAND4_in[0] ,
         \SB4_4/Component_Function_5/NAND4_in[2] ,
         \SB4_4/Component_Function_5/NAND4_in[1] ,
         \SB4_4/Component_Function_5/NAND4_in[0] ,
         \SB4_5/Component_Function_0/NAND4_in[3] ,
         \SB4_5/Component_Function_0/NAND4_in[2] ,
         \SB4_5/Component_Function_0/NAND4_in[1] ,
         \SB4_5/Component_Function_0/NAND4_in[0] ,
         \SB4_5/Component_Function_1/NAND4_in[3] ,
         \SB4_5/Component_Function_1/NAND4_in[2] ,
         \SB4_5/Component_Function_1/NAND4_in[1] ,
         \SB4_5/Component_Function_1/NAND4_in[0] ,
         \SB4_5/Component_Function_5/NAND4_in[2] ,
         \SB4_5/Component_Function_5/NAND4_in[1] ,
         \SB4_5/Component_Function_5/NAND4_in[0] ,
         \SB4_6/Component_Function_0/NAND4_in[3] ,
         \SB4_6/Component_Function_0/NAND4_in[2] ,
         \SB4_6/Component_Function_0/NAND4_in[1] ,
         \SB4_6/Component_Function_0/NAND4_in[0] ,
         \SB4_6/Component_Function_1/NAND4_in[3] ,
         \SB4_6/Component_Function_1/NAND4_in[2] ,
         \SB4_6/Component_Function_1/NAND4_in[1] ,
         \SB4_6/Component_Function_1/NAND4_in[0] ,
         \SB4_6/Component_Function_5/NAND4_in[3] ,
         \SB4_6/Component_Function_5/NAND4_in[0] ,
         \SB4_7/Component_Function_0/NAND4_in[3] ,
         \SB4_7/Component_Function_0/NAND4_in[2] ,
         \SB4_7/Component_Function_0/NAND4_in[1] ,
         \SB4_7/Component_Function_0/NAND4_in[0] ,
         \SB4_7/Component_Function_1/NAND4_in[3] ,
         \SB4_7/Component_Function_1/NAND4_in[1] ,
         \SB4_7/Component_Function_1/NAND4_in[0] ,
         \SB4_7/Component_Function_5/NAND4_in[3] ,
         \SB4_7/Component_Function_5/NAND4_in[2] ,
         \SB4_7/Component_Function_5/NAND4_in[1] ,
         \SB4_7/Component_Function_5/NAND4_in[0] ,
         \SB4_8/Component_Function_0/NAND4_in[1] ,
         \SB4_8/Component_Function_1/NAND4_in[3] ,
         \SB4_8/Component_Function_1/NAND4_in[2] ,
         \SB4_8/Component_Function_1/NAND4_in[1] ,
         \SB4_8/Component_Function_1/NAND4_in[0] ,
         \SB4_8/Component_Function_5/NAND4_in[3] ,
         \SB4_8/Component_Function_5/NAND4_in[0] ,
         \SB4_9/Component_Function_0/NAND4_in[3] ,
         \SB4_9/Component_Function_0/NAND4_in[2] ,
         \SB4_9/Component_Function_0/NAND4_in[1] ,
         \SB4_9/Component_Function_1/NAND4_in[3] ,
         \SB4_9/Component_Function_1/NAND4_in[2] ,
         \SB4_9/Component_Function_1/NAND4_in[1] ,
         \SB4_9/Component_Function_1/NAND4_in[0] ,
         \SB4_9/Component_Function_5/NAND4_in[3] ,
         \SB4_9/Component_Function_5/NAND4_in[1] ,
         \SB4_9/Component_Function_5/NAND4_in[0] ,
         \SB4_10/Component_Function_0/NAND4_in[0] ,
         \SB4_10/Component_Function_1/NAND4_in[3] ,
         \SB4_10/Component_Function_1/NAND4_in[0] ,
         \SB4_10/Component_Function_5/NAND4_in[2] ,
         \SB4_10/Component_Function_5/NAND4_in[1] ,
         \SB4_11/Component_Function_0/NAND4_in[2] ,
         \SB4_11/Component_Function_0/NAND4_in[1] ,
         \SB4_11/Component_Function_0/NAND4_in[0] ,
         \SB4_11/Component_Function_1/NAND4_in[3] ,
         \SB4_11/Component_Function_1/NAND4_in[2] ,
         \SB4_11/Component_Function_1/NAND4_in[1] ,
         \SB4_11/Component_Function_1/NAND4_in[0] ,
         \SB4_11/Component_Function_5/NAND4_in[3] ,
         \SB4_11/Component_Function_5/NAND4_in[2] ,
         \SB4_11/Component_Function_5/NAND4_in[1] ,
         \SB4_11/Component_Function_5/NAND4_in[0] ,
         \SB4_12/Component_Function_0/NAND4_in[3] ,
         \SB4_12/Component_Function_0/NAND4_in[2] ,
         \SB4_12/Component_Function_0/NAND4_in[1] ,
         \SB4_12/Component_Function_1/NAND4_in[2] ,
         \SB4_12/Component_Function_1/NAND4_in[1] ,
         \SB4_12/Component_Function_1/NAND4_in[0] ,
         \SB4_12/Component_Function_5/NAND4_in[3] ,
         \SB4_12/Component_Function_5/NAND4_in[2] ,
         \SB4_13/Component_Function_0/NAND4_in[1] ,
         \SB4_13/Component_Function_0/NAND4_in[0] ,
         \SB4_13/Component_Function_1/NAND4_in[2] ,
         \SB4_13/Component_Function_1/NAND4_in[1] ,
         \SB4_13/Component_Function_1/NAND4_in[0] ,
         \SB4_13/Component_Function_5/NAND4_in[2] ,
         \SB4_13/Component_Function_5/NAND4_in[1] ,
         \SB4_13/Component_Function_5/NAND4_in[0] ,
         \SB4_14/Component_Function_0/NAND4_in[3] ,
         \SB4_14/Component_Function_0/NAND4_in[2] ,
         \SB4_14/Component_Function_0/NAND4_in[0] ,
         \SB4_14/Component_Function_1/NAND4_in[3] ,
         \SB4_14/Component_Function_1/NAND4_in[2] ,
         \SB4_14/Component_Function_1/NAND4_in[1] ,
         \SB4_14/Component_Function_1/NAND4_in[0] ,
         \SB4_14/Component_Function_5/NAND4_in[3] ,
         \SB4_14/Component_Function_5/NAND4_in[2] ,
         \SB4_14/Component_Function_5/NAND4_in[1] ,
         \SB4_14/Component_Function_5/NAND4_in[0] ,
         \SB4_15/Component_Function_0/NAND4_in[3] ,
         \SB4_15/Component_Function_0/NAND4_in[2] ,
         \SB4_15/Component_Function_0/NAND4_in[1] ,
         \SB4_15/Component_Function_0/NAND4_in[0] ,
         \SB4_15/Component_Function_1/NAND4_in[2] ,
         \SB4_15/Component_Function_1/NAND4_in[1] ,
         \SB4_15/Component_Function_5/NAND4_in[3] ,
         \SB4_15/Component_Function_5/NAND4_in[1] ,
         \SB4_15/Component_Function_5/NAND4_in[0] ,
         \SB4_16/Component_Function_0/NAND4_in[2] ,
         \SB4_16/Component_Function_0/NAND4_in[1] ,
         \SB4_16/Component_Function_0/NAND4_in[0] ,
         \SB4_16/Component_Function_1/NAND4_in[3] ,
         \SB4_16/Component_Function_1/NAND4_in[1] ,
         \SB4_16/Component_Function_1/NAND4_in[0] ,
         \SB4_16/Component_Function_5/NAND4_in[3] ,
         \SB4_16/Component_Function_5/NAND4_in[2] ,
         \SB4_17/Component_Function_0/NAND4_in[3] ,
         \SB4_17/Component_Function_0/NAND4_in[1] ,
         \SB4_17/Component_Function_1/NAND4_in[3] ,
         \SB4_17/Component_Function_1/NAND4_in[2] ,
         \SB4_17/Component_Function_1/NAND4_in[1] ,
         \SB4_17/Component_Function_1/NAND4_in[0] ,
         \SB4_17/Component_Function_5/NAND4_in[3] ,
         \SB4_17/Component_Function_5/NAND4_in[2] ,
         \SB4_17/Component_Function_5/NAND4_in[1] ,
         \SB4_17/Component_Function_5/NAND4_in[0] ,
         \SB4_18/Component_Function_0/NAND4_in[3] ,
         \SB4_18/Component_Function_0/NAND4_in[2] ,
         \SB4_18/Component_Function_0/NAND4_in[1] ,
         \SB4_18/Component_Function_0/NAND4_in[0] ,
         \SB4_18/Component_Function_1/NAND4_in[3] ,
         \SB4_18/Component_Function_1/NAND4_in[2] ,
         \SB4_18/Component_Function_1/NAND4_in[1] ,
         \SB4_18/Component_Function_1/NAND4_in[0] ,
         \SB4_18/Component_Function_5/NAND4_in[3] ,
         \SB4_18/Component_Function_5/NAND4_in[2] ,
         \SB4_18/Component_Function_5/NAND4_in[1] ,
         \SB4_18/Component_Function_5/NAND4_in[0] ,
         \SB4_19/Component_Function_0/NAND4_in[3] ,
         \SB4_19/Component_Function_0/NAND4_in[2] ,
         \SB4_19/Component_Function_1/NAND4_in[3] ,
         \SB4_19/Component_Function_1/NAND4_in[2] ,
         \SB4_19/Component_Function_5/NAND4_in[1] ,
         \SB4_19/Component_Function_5/NAND4_in[0] ,
         \SB4_20/Component_Function_0/NAND4_in[0] ,
         \SB4_20/Component_Function_1/NAND4_in[3] ,
         \SB4_20/Component_Function_1/NAND4_in[2] ,
         \SB4_20/Component_Function_1/NAND4_in[1] ,
         \SB4_20/Component_Function_1/NAND4_in[0] ,
         \SB4_20/Component_Function_5/NAND4_in[3] ,
         \SB4_20/Component_Function_5/NAND4_in[2] ,
         \SB4_20/Component_Function_5/NAND4_in[0] ,
         \SB4_21/Component_Function_0/NAND4_in[3] ,
         \SB4_21/Component_Function_0/NAND4_in[2] ,
         \SB4_21/Component_Function_0/NAND4_in[0] ,
         \SB4_21/Component_Function_1/NAND4_in[3] ,
         \SB4_21/Component_Function_1/NAND4_in[1] ,
         \SB4_21/Component_Function_5/NAND4_in[3] ,
         \SB4_21/Component_Function_5/NAND4_in[1] ,
         \SB4_21/Component_Function_5/NAND4_in[0] ,
         \SB4_22/Component_Function_0/NAND4_in[2] ,
         \SB4_22/Component_Function_0/NAND4_in[1] ,
         \SB4_22/Component_Function_0/NAND4_in[0] ,
         \SB4_22/Component_Function_1/NAND4_in[3] ,
         \SB4_22/Component_Function_1/NAND4_in[2] ,
         \SB4_22/Component_Function_1/NAND4_in[1] ,
         \SB4_22/Component_Function_1/NAND4_in[0] ,
         \SB4_22/Component_Function_5/NAND4_in[2] ,
         \SB4_22/Component_Function_5/NAND4_in[1] ,
         \SB4_22/Component_Function_5/NAND4_in[0] ,
         \SB4_23/Component_Function_0/NAND4_in[3] ,
         \SB4_23/Component_Function_0/NAND4_in[2] ,
         \SB4_23/Component_Function_0/NAND4_in[1] ,
         \SB4_23/Component_Function_0/NAND4_in[0] ,
         \SB4_23/Component_Function_1/NAND4_in[3] ,
         \SB4_23/Component_Function_1/NAND4_in[2] ,
         \SB4_23/Component_Function_1/NAND4_in[1] ,
         \SB4_23/Component_Function_1/NAND4_in[0] ,
         \SB4_23/Component_Function_5/NAND4_in[2] ,
         \SB4_23/Component_Function_5/NAND4_in[1] ,
         \SB4_23/Component_Function_5/NAND4_in[0] ,
         \SB4_24/Component_Function_0/NAND4_in[3] ,
         \SB4_24/Component_Function_0/NAND4_in[2] ,
         \SB4_24/Component_Function_0/NAND4_in[0] ,
         \SB4_24/Component_Function_1/NAND4_in[3] ,
         \SB4_24/Component_Function_1/NAND4_in[2] ,
         \SB4_24/Component_Function_1/NAND4_in[1] ,
         \SB4_24/Component_Function_1/NAND4_in[0] ,
         \SB4_24/Component_Function_5/NAND4_in[2] ,
         \SB4_24/Component_Function_5/NAND4_in[1] ,
         \SB4_24/Component_Function_5/NAND4_in[0] ,
         \SB4_25/Component_Function_0/NAND4_in[3] ,
         \SB4_25/Component_Function_0/NAND4_in[2] ,
         \SB4_25/Component_Function_0/NAND4_in[1] ,
         \SB4_25/Component_Function_0/NAND4_in[0] ,
         \SB4_25/Component_Function_1/NAND4_in[3] ,
         \SB4_25/Component_Function_1/NAND4_in[2] ,
         \SB4_25/Component_Function_1/NAND4_in[1] ,
         \SB4_25/Component_Function_5/NAND4_in[2] ,
         \SB4_25/Component_Function_5/NAND4_in[1] ,
         \SB4_25/Component_Function_5/NAND4_in[0] ,
         \SB4_26/Component_Function_0/NAND4_in[2] ,
         \SB4_26/Component_Function_0/NAND4_in[1] ,
         \SB4_26/Component_Function_1/NAND4_in[3] ,
         \SB4_26/Component_Function_1/NAND4_in[2] ,
         \SB4_26/Component_Function_1/NAND4_in[1] ,
         \SB4_26/Component_Function_1/NAND4_in[0] ,
         \SB4_26/Component_Function_5/NAND4_in[3] ,
         \SB4_26/Component_Function_5/NAND4_in[2] ,
         \SB4_26/Component_Function_5/NAND4_in[0] ,
         \SB4_27/Component_Function_0/NAND4_in[2] ,
         \SB4_27/Component_Function_0/NAND4_in[0] ,
         \SB4_27/Component_Function_1/NAND4_in[3] ,
         \SB4_27/Component_Function_1/NAND4_in[2] ,
         \SB4_27/Component_Function_1/NAND4_in[1] ,
         \SB4_27/Component_Function_1/NAND4_in[0] ,
         \SB4_27/Component_Function_5/NAND4_in[3] ,
         \SB4_27/Component_Function_5/NAND4_in[2] ,
         \SB4_27/Component_Function_5/NAND4_in[1] ,
         \SB4_27/Component_Function_5/NAND4_in[0] ,
         \SB4_28/Component_Function_0/NAND4_in[2] ,
         \SB4_28/Component_Function_0/NAND4_in[1] ,
         \SB4_28/Component_Function_1/NAND4_in[3] ,
         \SB4_28/Component_Function_1/NAND4_in[1] ,
         \SB4_28/Component_Function_5/NAND4_in[1] ,
         \SB4_28/Component_Function_5/NAND4_in[0] ,
         \SB4_29/Component_Function_0/NAND4_in[1] ,
         \SB4_29/Component_Function_0/NAND4_in[0] ,
         \SB4_29/Component_Function_1/NAND4_in[3] ,
         \SB4_29/Component_Function_1/NAND4_in[2] ,
         \SB4_29/Component_Function_1/NAND4_in[1] ,
         \SB4_29/Component_Function_1/NAND4_in[0] ,
         \SB4_29/Component_Function_5/NAND4_in[2] ,
         \SB4_29/Component_Function_5/NAND4_in[1] ,
         \SB4_29/Component_Function_5/NAND4_in[0] ,
         \SB4_30/Component_Function_0/NAND4_in[3] ,
         \SB4_30/Component_Function_0/NAND4_in[1] ,
         \SB4_30/Component_Function_0/NAND4_in[0] ,
         \SB4_30/Component_Function_1/NAND4_in[3] ,
         \SB4_30/Component_Function_1/NAND4_in[2] ,
         \SB4_30/Component_Function_1/NAND4_in[1] ,
         \SB4_30/Component_Function_1/NAND4_in[0] ,
         \SB4_30/Component_Function_5/NAND4_in[2] ,
         \SB4_30/Component_Function_5/NAND4_in[1] ,
         \SB4_30/Component_Function_5/NAND4_in[0] ,
         \SB4_31/Component_Function_0/NAND4_in[2] ,
         \SB4_31/Component_Function_0/NAND4_in[1] ,
         \SB4_31/Component_Function_0/NAND4_in[0] ,
         \SB4_31/Component_Function_1/NAND4_in[3] ,
         \SB4_31/Component_Function_1/NAND4_in[2] ,
         \SB4_31/Component_Function_1/NAND4_in[1] ,
         \SB4_31/Component_Function_1/NAND4_in[0] ,
         \SB4_31/Component_Function_5/NAND4_in[3] ,
         \SB4_31/Component_Function_5/NAND4_in[1] ,
         \SB4_31/Component_Function_5/NAND4_in[0] , n8, n9, n13, n20, n33, n44,
         n45, n50, n51, n64, n84, n87, n89, n90, n94, n99, n102, n113, n115,
         n127, n145, n148, n153, n158, n164, n167, n171, n1, n2, n3, n4, n5,
         n6, n7, n10, n11, n12, n14, n15, n16, n17, n18, n19, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n46, n47, n48, n49, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n85, n86,
         n88, n91, n92, n95, n96, n97, n98, n100, n101, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n114, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n146, n147, n149, n150, n151, n152, n154, n155, n156,
         n157, n159, n160, n161, n162, n163, n165, n166, n168, n169, n170,
         n172, n173, n174, n175, n176, n177, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n571, n572, n573, n575, n578, n583, n588, n589, n590, n592,
         n593, n594, n595, n597, n598, n599, n600, n601, n602, n603, n604,
         n606, n610, n611, n614, n615, n617, n621, n626, n630, n633, n634,
         n635, n639, n641, n642, n643, n646, n647, n648, n649, n650, n655,
         n656, n660, n665, n666, n669, n671, n673, n674, n675, n681, n683,
         n684, n685, n686, n687, n690, n694, n702, n706, n709, n710, n714,
         n715, n716, n724, n727, n729, n733, n736, n739, n741, n742, n744,
         n745, n746, n748, n750, n753, n756, n757, n758, n759, n761, n763,
         n766, n774, n775, n784, n788, n790, n792, n795, n796, n797, n798,
         n801, n802, n804, n806, n807, n809, n813, n816, n817, n818, n821,
         n823, n826, n829, n830, n833, n835, n836, n840, n845, n849, n851,
         n852, n853, n854, n855, n857, n859, n861, n862, n863, n864, n865,
         n869, n871, n874, n877, n878, n879, n880, n881, n882, n883, n885,
         n886, n887, n890, n893, n895, n897, n898, n901, n903, n904, n905,
         n906, n907, n910, n911, n912, n913, n914, n916, n917, n919, n920,
         n922, n924, n929, n931, n932, n933, n934, n935, n936, n939, n940,
         n942, n944, n945, n946, n954, n955, n958, n959, n960, n961, n964,
         n965, n966, n967, n969, n971, n973, n974, n976, n979, n980, n982,
         n986, n988, n993, n994, n996, n997, n998, n1000, n1002, n1003, n1004,
         n1005, n1010, n1012, n1014, n1016, n1018, n1019, n1020, n1025, n1026,
         n1027, n1029, n1030, n1032, n1034, n1035, n1037, n1043, n1045, n1046,
         n1047, n1048, n1049, n1052, n1054, n1061, n1062, n1066, n1067, n1068,
         n1069, n1071, n1073, n1075, n1076, n1077, n1078, n1079, n1080, n1082,
         n1083, n1087, n1089, n1090, n1091, n1092, n1095, n1096, n1097, n1101,
         n1102, n1103, n1104, n1105, n1106, n1109, n1111, n1112, n1115, n1116,
         n1117, n1120, n1121, n1122, n1123, n1125, n1126, n1128, n1131, n1133,
         n1137, n1142, n1143, n1144, n1146, n1148, n1154, n1155, n1156, n1157,
         n1158, n1161, n1163, n1165, n1166, n1167, n1169, n1170, n1171, n1176,
         n1179, n1182, n1183, n1184, n1187, n1188, n1189, n1191, n1192, n1195,
         n1196, n1197, n1199, n1200, n1203, n1205, n1208, n1209, n1210, n1211,
         n1212, n1214, n1216, n1222, n1223, n1224, n1228, n1230, n1233, n1234,
         n1235, n1236, n1237, n1239, n1242, n1243, n1244, n1246, n1247, n1248,
         n1251, n1253, n1254, n1255, n1256, n1259, n1260, n1261, n1262, n1263,
         n1266, n1268, n1270, n1271, n1274, n1277, n1282, n1283, n1284, n1287,
         n1291, n1294, n1295, n1296, n1303, n1304, n1305, n1311, n1312, n1313,
         n1315, n1317, n1318, n1319, n1321, n1324, n1327, n1333, n1335, n1337,
         n1339, n1341, n1344, n1348, n1351, n1353, n1355, n1356, n1359, n1360,
         n1361, n1363, n1364, n1366, n1369, n1371, n1372, n1375, n1376, n1379,
         n1381, n1383, n1384, n1387, n1389, n1390, n1391, n1392, n1393, n1394,
         n1398, n1399, n1400, n1401, n1403, n1407, n1411, n1412, n1414, n1415,
         n1417, n1420, n1422, n1423, n1424, n1426, n1427, n1428, n1429, n1431,
         n1432, n1433, n1436, n1447, n1448, n1449, n1450, n1453, n1454, n1457,
         n1460, n1461, n1465, n1466, n1467, n1468, n1469, n1470, n1475, n1479,
         n1480, n1481, n1482, n1483, n1485, n1487, n1488, n1490, n1491, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1504, n1506,
         n1507, n1508, n1509, n1510, n1512, n1518, n1519, n1520, n1523, n1526,
         n1529, n1532, n1534, n1535, n1536, n1537, n1538, n1541, n1543, n1544,
         n1545, n1546, n1547, n1548, n1550, n1551, n1552, n1557, n1558, n1560,
         n1562, n1564, n1566, n1568, n1569, n1571, n1573, n1574, n1575, n1576,
         n1577, n1579, n1580, n1582, n1584, n1587, n1589, n1590, n1591, n1592,
         n1593, n1594, n1596, n1599, n1600, n1604, n1608, n1609, n1610, n1612,
         n1613, n1614, n1615, n1617, n1618, n1622, n1623, n1624, n1625, n1628,
         n1630, n1631, n1634, n1636, n1637, n1638, n1640, n1641, n1642, n1643,
         n1645, n1647, n1650, n1651, n1653, n1654, n1655, n1656, n1659, n1660,
         n1662, n1663, n1666, n1669, n1670, n1671, n1672, n1677, n1678, n1680,
         n1682, n1683, n1685, n1689, n1693, n1694, n1695, n1696, n1698, n1699,
         n1700, n1702, n1704, n1705, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1723, n1725,
         n1726, n1728, n1729, n1732, n1733, n1734, n1736, n1739, n1742, n1743,
         n1744, n1745, n1746, n1749, n1752, n1753, n1759, n1763, n1764, n1765,
         n1766, n1767, n1769, n1770, n1771, n1772, n1773, n1775, n1776, n1777,
         n1778, n1780, n1781, n1782, n1786, n1787, n1788, n1789, n1790, n1793,
         n1794, n1795, n1796, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1813, n1814, n1815, n1817,
         n1818, n1819, n1821, n1823, n1825, n1826, n1827, n1828, n1832, n1833,
         n1835, n1836, n1838, n1839, n1841, n1844, n1845, n1846, n1848, n1849,
         n1850, n1851, n1853, n1854, n1855, n1856, n1861, n1862, n1863, n1866,
         n1868, n1870, n1871, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1882, n1883, n1884, n1890, n1892, n1893, n1896, n1898, n1902, n1903,
         n1904, n1905, n1908, n1910, n1911, n1912, n1913, n1915, n1916, n1918,
         n1919, n1920, n1922, n1923, n1925, n1927, n1928, n1930, n1931, n1932,
         n1933, n1935, n1936, n1937, n1938, n1940, n1942, n1946, n1947, n1949,
         n1950, n1952, n1953, n1956, n1957, n1958, n1959, n1962, n1963, n1965,
         n1967, n1968, n1970, n1972, n1973, n1974, n1975, n1980, n1982, n1983,
         n1984, n1985, n1986, n1991, n1993, n1994, n1995, n1997, n1999, n2001,
         n2003, n2004, n2005, n2006, n2009, n2011, n2012, n2013, n2014, n2015,
         n2017, n2018, n2021, n2022, n2024, n2025, n2026, n2027, n2030, n2031,
         n2032, n2033, n2034, n2037, n2039, n2041, n2042, n2043, n2045, n2046,
         n2047, n2048, n2049, n2053, n2054, n2055, n2056, n2059, n2060, n2061,
         n2062, n2063, n2064, n2066, n2067, n2069, n2070, n2071, n2073, n2074,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2085, n2086,
         n2088, n2089, n2091, n2092, n2093, n2094, n2096, n2097, n2098, n2100,
         n2101, n2103, n2104, n2105, n2107, n2109, n2110, n2111, n2115, n2116,
         n2117, n2119, n2120, n2121, n2124, n2126, n2128, n2129, n2132, n2134,
         n2135, n2136, n2137, n2140, n2141, n2142, n2145, n2147, n2149, n2150,
         n2151, n2152, n2153, n2156, n2157, n2159, n2160, n2161, n2163, n2164,
         n2165, n2167, n2168, n2170, n2172, n2174, n2175, n2177, n2178, n2179,
         n2180, n2181, n2183, n2185, n2186, n2188, n2189, n2190, n2191, n2192,
         n2193, n2195, n2196, n2197, n2199, n2200, n2202, n2203, n2204, n2206,
         n2207, n2209, n2210, n2211, n2212, n2213, n2215, n2216, n2217, n2221,
         n2222, n2223, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2245, n2246, n2248, n2251, n2253, n2254, n2255, n2256, n2258, n2261,
         n2262, n2263, n2265, n2266, n2268, n2270, n2273, n2274, n2278, n2279,
         n2280, n2281, n2283, n2284, n2285, n2286, n2287, n2291, n2292, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2304, n2305, n2306, n2308,
         n2309, n2310, n2311, n2312, n2313, n2315, n2316, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2326, n2328, n2330, n2332, n2333, n2334,
         n2335, n2337, n2340, n2343, n2344, n2346, n2347, n2348, n2349, n2350,
         n2351, n2353, n2355, n2359, n2360, n2361, n2364, n2365, n2366, n2367,
         n2369, n2371, n2372, n2374, n2375, n2377, n2378, n2379, n2380, n2381,
         n2382, n2384, n2387, n2388, n2389, n2390, n2392, n2393, n2394, n2395,
         n2396, n2398, n2399, n2400, n2401, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2416, n2417, n2418,
         n2421, n2422, n2423, n2424, n2425, n2427, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2444, n2445, n2446, n2447, n2450, n2452, n2453, n2454, n2455, n2457,
         n2458, n2459, n2460, n2462, n2463, n2467, n2469, n2474, n2476, n2479,
         n2480, n2482, n2483, n2485, n2486, n2487, n2490, n2495, n2496, n2497,
         n2498, n2500, n2501, n2502, n2503, n2506, n2507, n2508, n2509, n2511,
         n2514, n2515, n2516, n2518, n2519, n2520, n2521, n2522, n2525, n2528,
         n2530, n2531, n2532, n2533, n2534, n2535, n2537, n2538, n2540, n2544,
         n2546, n2547, n2552, n2553, n2554, n2555, n2556, n2558, n2561, n2562,
         n2563, n2564, n2565, n2566, n2569, n2570, n2572, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2588, n2589, n2590, n2592,
         n2593, n2594, n2595, n2597, n2599, n2600, n2601, n2602, n2604, n2605,
         n2606, n2609, n2610, n2611, n2612, n2613, n2614, n2616, n2618, n2619,
         n2620, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2632, n2633, n2634, n2635, n2636, n2641, n2642, n2643, n2645, n2648,
         n2649, n2651, n2652, n2653, n2655, n2656, n2657, n2660, n2661, n2662,
         n2663, n2664, n2665, n2667, n2668, n2669, n2670, n2672, n2673, n2674,
         n2675, n2676, n2680, n2682, n2683, n2684, n2685, n2687, n2693, n2694,
         n2695, n2697, n2698, n2700, n2702, n2703, n2707, n2708, n2712, n2713,
         n2717, n2718, n2721, n2723, n2724, n2725, n2728, n2730, n2731, n2733,
         n2735, n2736, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2753, n2755, n2756, n2759, n2760, n2761,
         n2762, n2763, n2764, n2767, n2768, n2769, n2771, n2772, n2775, n2776,
         n2778, n2779, n2780, n2781, n2783, n2786, n2787, n2788, n2789, n2791,
         n2792, n2795, n2797, n2801, n2802, n2803, n2804, n2805, n2806, n2810,
         n2811, n2814, n2815, n2816, n2819, n2821, n2822, n2823, n2824, n2826,
         n2827, n2828, n2829, n2831, n2832, n2833, n2834, n2835, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2852, n2854, n2855, n2856, n2857, n2858, n2860, n2861, n2862, n2864,
         n2869, n2870, n2872, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2890, n2891, n2893, n2894, n2897, n2898,
         n2901, n2902, n2903, n2905, n2907, n2909, n2910, n2911, n2912, n2914,
         n2915, n2916, n2917, n2918, n2921, n2922, n2923, n2924, n2925, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2936, n2938, n2939, n2941,
         n2943, n2945, n2946, n2948, n2950, n2951, n2952, n2955, n2957, n2960,
         n2961, n2962, n2963, n2965, n2966, n2967, n2968, n2969, n2971, n2972,
         n2973, n2976, n2977, n2978, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2991, n2993, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3009,
         n3011, n3012, n3013, n3016, n3018, n3020, n3023, n3025, n3027, n3029,
         n3030, n3031, n3033, n3034, n3037, n3038, n3039, n3041, n3044, n3046,
         n3049, n3051, n3053, n3055, n3056, n3060, n3061, n3063, n3064, n3065,
         n3067, n3068, n3069, n3070, n3073, n3075, n3076, n3078, n3079, n3080,
         n3082, n3083, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3096, n3097, n3098, n3100, n3101, n3102, n3103, n3104,
         n3106, n3107, n3109, n3110, n3113, n3114, n3115, n3116, n3117, n3118,
         n3122, n3123, n3125, n3127, n3131, n3133, n3134, n3135, n3136, n3137,
         n3139, n3140, n3141, n3145, n3147, n3148, n3149, n3150, n3152, n3153,
         n3154, n3157, n3158, n3159, n3161, n3162, n3165, n3166, n3167, n3168,
         n3169, n3171, n3173, n3175, n3177, n3178, n3179, n3180, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3190, n3191, n3193, n3194, n3195,
         n3196, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3212, n3213, n3214, n3215, n3216, n3218, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3229, n3231, n3233, n3234,
         n3236, n3242, n3246, n3248, n3249, n3252, n3253, n3254, n3255, n3256,
         n3257, n3262, n3263, n3265, n3266, n3270, n3271, n3272, n3274, n3276,
         n3279, n3280, n3284, n3286, n3287, n3288, n3289, n3290, n3292, n3293,
         n3295, n3298, n3299, n3301, n3302, n3303, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3316, n3317, n3318, n3319, n3322, n3325,
         n3326, n3327, n3329, n3330, n3331, n3334, n3335, n3337, n3338, n3343,
         n3344, n3349, n3350, n3352, n3354, n3355, n3357, n3358, n3359, n3361,
         n3362, n3363, n3364, n3365, n3367, n3368, n3370, n3373, n3374, n3375,
         n3376, n3377, n3378, n3380, n3381, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3402,
         n3403, n3404, n3408, n3411, n3412, n3413, n3416, n3417, n3421, n3422,
         n3423, n3424, n3425, n3428, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3439, n3440, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3454, n3455, n3456, n3457, n3458, n3460, n3464, n3465,
         n3466, n3467, n3468, n3471, n3472, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3484, n3485, n3486, n3487, n3489, n3490, n3491, n3494,
         n3495, n3496, n3497, n3499, n3500, n3501, n3503, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3515, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3530,
         n3532, n3534, n3535, n3537, n3539, n3540, n3541, n3542, n3543, n3544,
         n3546, n3548, n3551, n3552, n3553, n3554, n3556, n3557, n3561, n3562,
         n3563, n3568, n3570, n3573, n3574, n3575, n3576, n3579, n3580, n3581,
         n3583, n3584, n3585, n3586, n3588, n3590, n3591, n3596, n3597, n3598,
         n3602, n3605, n3607, n3608, n3609, n3611, n3613, n3617, n3620, n3621,
         n3622, n3623, n3625, n3626, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3639, n3640, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3651, n3652, n3654, n3660, n3661, n3662, n3664,
         n3666, n3668, n3672, n3674, n3676, n3678, n3680, n3681, n3683, n3684,
         n3685, n3688, n3689, n3690, n3691, n3697, n3698, n3699, n3700, n3701,
         n3703, n3704, n3707, n3708, n3710, n3711, n3712, n3714, n3716, n3717,
         n3718, n3721, n3722, n3723, n3724, n3725, n3726, n3728, n3729, n3730,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3740, n3742, n3743,
         n3744, n3745, n3746, n3747, n3749, n3750, n3751, n3752, n3753, n3754,
         n3756, n3757, n3758, n3762, n3763, n3765, n3766, n3769, n3770, n3773,
         n3774, n3775, n3776, n3777, n3780, n3781, n3782, n3783, n3785, n3787,
         n3788, n3789, n3790, n3792, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3802, n3804, n3805, n3806, n3807, n3808, n3810, n3811, n3812,
         n3813, n3814, n3815, n3817, n3819, n3820, n3822, n3824, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3836, n3838, n3839, n3840, n3842,
         n3843, n3844, n3846, n3847, n3848, n3851, n3852, n3854, n3855, n3857,
         n3858, n3860, n3862, n3863, n3864, n3865, n3866, n3868, n3870, n3872,
         n3874, n3875, n3877, n3878, n3879, n3880, n3882, n3883, n3884, n3885,
         n3886, n3887, n3891, n3892, n3898, n3900, n3902, n3904, n3905, n3907,
         n3909, n3912, n3914, n3916, n3919, n3920, n3921, n3922, n3923, n3924,
         n3927, n3928, n3930, n3931, n3932, n3933, n3935, n3936, n3937, n3938,
         n3939, n3940, n3942, n3943, n3946, n3948, n3949, n3950, n3951, n3953,
         n3954, n3956, n3957, n3960, n3961, n3963, n3965, n3966, n3967, n3968,
         n3970, n3971, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4009, n4010, n4012, n4015,
         n4016, n4017, n4018, n4020, n4022, n4023, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4036, n4037, n4038, n4043, n4044,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4055, n4056,
         n4058, n4060, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4073, n4074, n4075, n4077, n4079, n4081, n4082, n4083, n4084,
         n4086, n4087, n4088, n4089, n4090, n4093, n4096, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4107, n4108, n4109, n4111, n4112,
         n4113, n4114, n4115, n4117, n4118, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4129, n4130, n4132, n4133, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4159, n4160, n4161,
         n4162, n4165, n4167, n4169, n4170, n4171, n4172, n4174, n4175, n4176,
         n4177, n4178, n4180, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4207, n4213, n4214, n4219, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4231, n4232,
         n4233, n4235, n4236, n4238, n4239, n4240, n4245, n4246, n4248, n4249,
         n4250, n4252, n4255, n4257, n4258, n4259, n4261, n4263, n4264, n4266,
         n4267, n4268, n4269, n4270, n4272, n4274, n4275, n4276, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4291, n4292,
         n4293, n4295, n4297, n4298, n4299, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4309, n4310, n4314, n4315, n4316, n4317, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4339, n4340, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4350, n4351, n4352, n4355, n4357, n4359,
         n4360, n4361, n4362, n4365, n4366, n4367, n4370, n4371, n4372, n4373,
         n4375, n4376, n4377, n4378, n4380, n4381, n4382, n4383, n4385, n4387,
         n4388, n4390, n4391, n4392, n4393, n4394, n4395, n4398, n4399, n4401,
         n4402, n4403, n4404, n4405, n4406, n4408, n4409, n4411, n4412, n4414,
         n4417, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4427, n4429,
         n4430, n4431, n4432, n4433, n4434, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4469, n4470, n4471, n4473, n4474, n4476,
         n4477, n4478, n4479, n4480, n4483, n4485, n4486, n4487, n4488, n4490,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4516, n4517, n4518, n4519, n4524, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4565, n4568, n4569, n4570, n4571, n4574, n4575, n4576, n4577,
         n4579, n4581, n4582, n4584, n4585, n4586, n4587, n4588, n4589, n4591,
         n4592, n4595, n4596, n4597, n4598, n4599, n4601, n4602, n4603, n4604,
         n4606, n4607, n4608, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4620, n4621, n4622, n4623, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4634, n4635, n4636, n4637, n4639, n4640,
         n4641, n4642, n4643, n4645, n4647, n4649, n4650, n4651, n4652, n4654,
         n4657, n4658, n4659, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4692, n4693, n4694, n4695, n4696, n4698, n4699, n4700,
         n4702, n4704, n4705, n4708, n4710, n4711, n4712, n4713, n4714, n4715,
         n4717, n4718, n4719, n4722, n4724, n4727, n4729, n4730, n4732, n4734,
         n4735, n4737, n4738, n4739, n4740, n4741, n4743, n4744, n4745, n4746,
         n4747, n4748, n4750, n4751, n4752, n4754, n4755, n4756, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4777, n4778, n4780, n4781, n4782,
         n4784, n4785, n4786, n4787, n4790, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4803, n4804, n4805, n4806, n4808,
         n4809, n4812, n4813, n4814, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4827, n4828, n4829, n4830, n4832, n4834,
         n4835, n4837, n4838, n4839, n4840, n4842, n4845, n4846, n4847, n4848,
         n4849, n4850, n4852, n4853, n4855, n4856, n4857, n4858, n4859, n4861,
         n4862, n4863, n4865, n4868, n4869, n4872, n4873, n4875, n4876, n4878,
         n4879, n4881, n4882, n4883, n4885, n4886, n4889, n4891, n4892, n4893,
         n4894, n4898, n4899, n4900, n4901, n4902, n4903, n4906, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4921,
         n4922, n4924, n4926, n4929, n4930, n4931, n4933, n4936, n4937, n4938,
         n4940, n4942, n4943, n4944, n4946, n4947, n4948, n4949, n4950, n4951,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4966, n4967, n4969, n4970, n4972, n4974, n4975, n4976,
         n4977, n4978, n4979, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4992, n4996, n4997, n4998, n5000, n5001, n5003,
         n5004, n5005, n5006, n5007, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5031, n5032, n5033, n5034, n5035,
         n5037, n5038, n5039, n5040, n5042, n5043, n5046, n5047, n5049, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5059, n5060, n5062, n5064,
         n5065, n5066, n5067, n5068, n5069, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5100, n5101, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5117, n5118, n5119, n5120,
         n5122, n5123, n5124, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5138, n5140, n5142, n5143, n5144, n5145, n5147, n5148,
         n5149, n5151, n5153, n5155, n5156, n5157, n5158, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5193, n5197, n5198,
         n5200, n5201, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5214, n5215, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5226, n5228, n5229, n5231, n5232, n5233, n5235, n5237, n5238,
         n5239, n5242, n5243, n5244, n5245, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5257, n5258, n5259, n5260, n5261, n5262,
         n5264, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5275, n5276,
         n5277, n5278, n5279, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5293, n5294, n5295, n5296, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5309, n5311,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5323,
         n5324, n5325, n5326, n5327, n5328, n5330, n5331, n5332, n5335, n5336,
         n5338, n5339, n5340, n5342, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5352, n5353, n5355, n5356, n5357, n5358, n5362, n5363, n5364,
         n5365, n5366, n5367, n5369, n5370, n5372, n5373, n5374, n5375, n5379,
         n5380, n5381, n5383, n5385, n5387, n5388, n5389, n5390, n5392, n5393,
         n5394, n5395, n5396, n5397, n5400, n5401, n5402, n5403, n5405, n5406,
         n5408, n5410, n5411, n5412, n5413, n5414, n5418, n5419, n5421, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590;

  XOR2_X1 \MC_ARK_ARC_1_0/X7_31_5  ( .A1(\MC_ARK_ARC_1_0/temp5[0] ), .A2(
        \MC_ARK_ARC_1_0/temp6[0] ), .Z(\MC_ARK_ARC_1_0/buf_output[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_31_5  ( .A1(\MC_ARK_ARC_1_0/temp3[0] ), .A2(
        \MC_ARK_ARC_1_0/temp4[0] ), .Z(\MC_ARK_ARC_1_0/temp6[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_5  ( .A1(\RI5[0][36] ), .A2(n41), .Z(
        \MC_ARK_ARC_1_0/temp4[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_31_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .A2(\RI5[0][66] ), .Z(\MC_ARK_ARC_1_0/temp3[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_31_5  ( .A1(\RI5[0][138] ), .A2(\RI5[0][162] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_4  ( .A1(\RI5[0][37] ), .A2(n95), .Z(
        \MC_ARK_ARC_1_0/temp4[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_31_4  ( .A1(\RI5[0][103] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[67] ), .Z(\MC_ARK_ARC_1_0/temp3[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_31_4  ( .A1(\RI5[0][163] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[139] ), .Z(\MC_ARK_ARC_1_0/temp2[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_31_4  ( .A1(\RI5[0][1] ), .A2(\RI5[0][187] ), .Z(
        \MC_ARK_ARC_1_0/temp1[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_31_3  ( .A1(\MC_ARK_ARC_1_0/temp6[2] ), .A2(
        \MC_ARK_ARC_1_0/temp5[2] ), .Z(\MC_ARK_ARC_1_0/buf_output[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_31_3  ( .A1(\MC_ARK_ARC_1_0/temp4[2] ), .A2(
        \MC_ARK_ARC_1_0/temp3[2] ), .Z(\MC_ARK_ARC_1_0/temp6[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_3  ( .A1(\RI5[0][38] ), .A2(n215), .Z(
        \MC_ARK_ARC_1_0/temp4[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_2  ( .A1(\RI5[0][39] ), .A2(n155), .Z(
        \MC_ARK_ARC_1_0/temp4[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_1  ( .A1(\RI5[0][40] ), .A2(n153), .Z(
        \MC_ARK_ARC_1_0/temp4[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_31_1  ( .A1(\RI5[0][142] ), .A2(\RI5[0][166] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_31_1  ( .A1(\RI5[0][4] ), .A2(\RI5[0][190] ), .Z(
        \MC_ARK_ARC_1_0/temp1[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_31_0  ( .A1(\MC_ARK_ARC_1_0/temp3[5] ), .A2(
        \MC_ARK_ARC_1_0/temp4[5] ), .Z(\MC_ARK_ARC_1_0/temp6[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[41] ), 
        .A2(n143), .Z(\MC_ARK_ARC_1_0/temp4[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_31_0  ( .A1(\RI5[0][107] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[71] ), .Z(\MC_ARK_ARC_1_0/temp3[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_31_0  ( .A1(\RI5[0][143] ), .A2(\RI5[0][167] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_31_0  ( .A1(\RI5[0][5] ), .A2(\RI5[0][191] ), .Z(
        \MC_ARK_ARC_1_0/temp1[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_30_5  ( .A1(\MC_ARK_ARC_1_0/temp4[6] ), .A2(
        \MC_ARK_ARC_1_0/temp3[6] ), .Z(\MC_ARK_ARC_1_0/temp6[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_5  ( .A1(\RI5[0][42] ), .A2(n532), .Z(
        \MC_ARK_ARC_1_0/temp4[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_30_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[108] ), 
        .A2(\RI5[0][72] ), .Z(\MC_ARK_ARC_1_0/temp3[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_30_5  ( .A1(\RI5[0][0] ), .A2(\RI5[0][6] ), .Z(
        \MC_ARK_ARC_1_0/temp1[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_30_4  ( .A1(\MC_ARK_ARC_1_0/temp6[7] ), .A2(
        \MC_ARK_ARC_1_0/temp5[7] ), .Z(\MC_ARK_ARC_1_0/buf_output[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_30_4  ( .A1(\MC_ARK_ARC_1_0/temp1[7] ), .A2(
        \MC_ARK_ARC_1_0/temp2[7] ), .Z(\MC_ARK_ARC_1_0/temp5[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .A2(n525), .Z(\MC_ARK_ARC_1_0/temp4[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_30_4  ( .A1(\RI5[0][169] ), .A2(\RI5[0][145] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_30_4  ( .A1(\RI5[0][7] ), .A2(\RI5[0][1] ), .Z(
        \MC_ARK_ARC_1_0/temp1[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_30_3  ( .A1(\MC_ARK_ARC_1_0/temp3[8] ), .A2(
        \MC_ARK_ARC_1_0/temp4[8] ), .Z(\MC_ARK_ARC_1_0/temp6[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_3  ( .A1(\RI5[0][44] ), .A2(n519), .Z(
        \MC_ARK_ARC_1_0/temp4[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_30_3  ( .A1(\RI5[0][2] ), .A2(\RI5[0][8] ), .Z(
        \MC_ARK_ARC_1_0/temp1[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_2  ( .A1(\RI5[0][45] ), .A2(n138), .Z(
        \MC_ARK_ARC_1_0/temp4[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_30_2  ( .A1(\RI5[0][147] ), .A2(\RI5[0][171] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_1  ( .A1(\RI5[0][46] ), .A2(n141), .Z(
        \MC_ARK_ARC_1_0/temp4[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_30_1  ( .A1(\RI5[0][112] ), .A2(\RI5[0][76] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_30_1  ( .A1(\RI5[0][148] ), .A2(\RI5[0][172] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_0  ( .A1(\SB2_0_24/buf_output[5] ), .A2(n132), 
        .Z(\MC_ARK_ARC_1_0/temp4[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_29_5  ( .A1(\MC_ARK_ARC_1_0/temp5[12] ), .A2(
        \MC_ARK_ARC_1_0/temp6[12] ), .Z(\MC_ARK_ARC_1_0/buf_output[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_29_5  ( .A1(\MC_ARK_ARC_1_0/temp3[12] ), .A2(
        \MC_ARK_ARC_1_0/temp4[12] ), .Z(\MC_ARK_ARC_1_0/temp6[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_5  ( .A1(\RI5[0][48] ), .A2(n496), .Z(
        \MC_ARK_ARC_1_0/temp4[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_29_5  ( .A1(\RI5[0][78] ), .A2(\RI5[0][114] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_29_5  ( .A1(\RI5[0][12] ), .A2(\RI5[0][6] ), .Z(
        \MC_ARK_ARC_1_0/temp1[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_29_4  ( .A1(\MC_ARK_ARC_1_0/temp3[13] ), .A2(
        \MC_ARK_ARC_1_0/temp4[13] ), .Z(\MC_ARK_ARC_1_0/temp6[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_29_4  ( .A1(\MC_ARK_ARC_1_0/temp1[13] ), .A2(
        \MC_ARK_ARC_1_0/temp2[13] ), .Z(\MC_ARK_ARC_1_0/temp5[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_4  ( .A1(\RI5[0][49] ), .A2(n94), .Z(
        \MC_ARK_ARC_1_0/temp4[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_29_4  ( .A1(\RI5[0][115] ), .A2(\RI5[0][79] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_29_4  ( .A1(\RI5[0][175] ), .A2(\RI5[0][151] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_29_4  ( .A1(\RI5[0][13] ), .A2(\RI5[0][7] ), .Z(
        \MC_ARK_ARC_1_0/temp1[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_3  ( .A1(\RI5[0][50] ), .A2(
        \MC_ARK_ARC_1_1/buf_keyinput[111] ), .Z(\MC_ARK_ARC_1_0/temp4[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_29_3  ( .A1(\RI5[0][176] ), .A2(\RI5[0][152] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_29_3  ( .A1(\RI5[0][8] ), .A2(\RI5[0][14] ), .Z(
        \MC_ARK_ARC_1_0/temp1[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_29_2  ( .A1(\MC_ARK_ARC_1_0/temp1[15] ), .A2(
        \MC_ARK_ARC_1_0/temp2[15] ), .Z(\MC_ARK_ARC_1_0/temp5[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_2  ( .A1(\RI5[0][51] ), .A2(n149), .Z(
        \MC_ARK_ARC_1_0/temp4[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_29_2  ( .A1(\RI5[0][153] ), .A2(\RI5[0][177] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_29_2  ( .A1(\RI5[0][9] ), .A2(\RI5[0][15] ), .Z(
        \MC_ARK_ARC_1_0/temp1[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_29_1  ( .A1(\MC_ARK_ARC_1_0/temp5[16] ), .A2(
        \MC_ARK_ARC_1_0/temp6[16] ), .Z(\MC_ARK_ARC_1_0/buf_output[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_29_1  ( .A1(\MC_ARK_ARC_1_0/temp3[16] ), .A2(
        \MC_ARK_ARC_1_0/temp4[16] ), .Z(\MC_ARK_ARC_1_0/temp6[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_29_1  ( .A1(\MC_ARK_ARC_1_0/temp1[16] ), .A2(
        \MC_ARK_ARC_1_0/temp2[16] ), .Z(\MC_ARK_ARC_1_0/temp5[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_1  ( .A1(\RI5[0][52] ), .A2(n475), .Z(
        \MC_ARK_ARC_1_0/temp4[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_29_1  ( .A1(\RI5[0][178] ), .A2(\RI5[0][154] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_29_0  ( .A1(\RI5[0][83] ), .A2(\RI5[0][119] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_28_5  ( .A1(\MC_ARK_ARC_1_0/temp1[18] ), .A2(
        \MC_ARK_ARC_1_0/temp2[18] ), .Z(\MC_ARK_ARC_1_0/temp5[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_5  ( .A1(\RI5[0][54] ), .A2(n463), .Z(
        \MC_ARK_ARC_1_0/temp4[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_28_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[84] ), 
        .A2(\RI5[0][120] ), .Z(\MC_ARK_ARC_1_0/temp3[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_28_5  ( .A1(\RI5[0][180] ), .A2(\RI5[0][156] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_28_5  ( .A1(\RI5[0][12] ), .A2(\RI5[0][18] ), .Z(
        \MC_ARK_ARC_1_0/temp1[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_28_4  ( .A1(\MC_ARK_ARC_1_0/temp4[19] ), .A2(
        \MC_ARK_ARC_1_0/temp3[19] ), .Z(\MC_ARK_ARC_1_0/temp6[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_4  ( .A1(\RI5[0][55] ), .A2(n457), .Z(
        \MC_ARK_ARC_1_0/temp4[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_28_4  ( .A1(\RI5[0][181] ), .A2(\RI5[0][157] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_28_4  ( .A1(\RI5[0][19] ), .A2(\RI5[0][13] ), .Z(
        \MC_ARK_ARC_1_0/temp1[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_28_2  ( .A1(\MC_ARK_ARC_1_0/temp3[21] ), .A2(
        \MC_ARK_ARC_1_0/temp4[21] ), .Z(\MC_ARK_ARC_1_0/temp6[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_2  ( .A1(\RI5[0][57] ), .A2(n114), .Z(
        \MC_ARK_ARC_1_0/temp4[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_28_2  ( .A1(\RI5[0][87] ), .A2(\RI5[0][123] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_28_2  ( .A1(\RI5[0][15] ), .A2(\RI5[0][21] ), .Z(
        \MC_ARK_ARC_1_0/temp1[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_1  ( .A1(\RI5[0][58] ), .A2(n172), .Z(
        \MC_ARK_ARC_1_0/temp4[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_28_1  ( .A1(\RI5[0][88] ), .A2(\RI5[0][124] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_28_1  ( .A1(\RI5[0][184] ), .A2(\RI5[0][160] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_28_1  ( .A1(\RI5[0][16] ), .A2(\RI5[0][22] ), .Z(
        \MC_ARK_ARC_1_0/temp1[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_0  ( .A1(\RI5[0][59] ), .A2(n434), .Z(
        \MC_ARK_ARC_1_0/temp4[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_28_0  ( .A1(\RI5[0][125] ), .A2(\RI5[0][89] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_28_0  ( .A1(\RI5[0][23] ), .A2(\RI5[0][17] ), .Z(
        \MC_ARK_ARC_1_0/temp1[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_27_5  ( .A1(\MC_ARK_ARC_1_0/temp3[24] ), .A2(
        \MC_ARK_ARC_1_0/temp4[24] ), .Z(\MC_ARK_ARC_1_0/temp6[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_5  ( .A1(\RI5[0][60] ), .A2(n428), .Z(
        \MC_ARK_ARC_1_0/temp4[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_27_5  ( .A1(\RI5[0][186] ), .A2(\RI5[0][162] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_27_5  ( .A1(\RI5[0][18] ), .A2(\RI5[0][24] ), .Z(
        \MC_ARK_ARC_1_0/temp1[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_27_4  ( .A1(\MC_ARK_ARC_1_0/temp6[25] ), .A2(
        \MC_ARK_ARC_1_0/temp5[25] ), .Z(\MC_ARK_ARC_1_0/buf_output[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_27_4  ( .A1(\MC_ARK_ARC_1_0/temp3[25] ), .A2(
        \MC_ARK_ARC_1_0/temp4[25] ), .Z(\MC_ARK_ARC_1_0/temp6[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_4  ( .A1(\RI5[0][61] ), .A2(n111), .Z(
        \MC_ARK_ARC_1_0/temp4[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_27_4  ( .A1(\RI5[0][127] ), .A2(\RI5[0][91] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_2  ( .A1(\RI5[0][63] ), .A2(n567), .Z(
        \MC_ARK_ARC_1_0/temp4[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_27_2  ( .A1(\RI5[0][93] ), .A2(\RI5[0][129] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .A2(n133), .Z(\MC_ARK_ARC_1_0/temp4[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_26_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[67] ), 
        .A2(n30), .Z(\MC_ARK_ARC_1_0/temp4[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_26_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[97] ), 
        .A2(\RI5[0][133] ), .Z(\MC_ARK_ARC_1_0/temp3[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_26_4  ( .A1(\RI5[0][1] ), .A2(\RI5[0][169] ), .Z(
        \MC_ARK_ARC_1_0/temp2[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_26_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .A2(\RI5[0][25] ), .Z(\MC_ARK_ARC_1_0/temp1[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_26_3  ( .A1(\RI5[0][170] ), .A2(\RI5[0][2] ), .Z(
        \MC_ARK_ARC_1_0/temp2[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_26_2  ( .A1(\MC_ARK_ARC_1_0/temp6[33] ), .A2(
        \MC_ARK_ARC_1_0/temp5[33] ), .Z(\MC_ARK_ARC_1_0/buf_output[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_26_2  ( .A1(\MC_ARK_ARC_1_0/temp1[33] ), .A2(
        \MC_ARK_ARC_1_0/temp2[33] ), .Z(\MC_ARK_ARC_1_0/temp5[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_26_2  ( .A1(\RI5[0][69] ), .A2(n535), .Z(
        \MC_ARK_ARC_1_0/temp4[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_26_2  ( .A1(\RI5[0][3] ), .A2(\RI5[0][171] ), .Z(
        \MC_ARK_ARC_1_0/temp2[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_26_2  ( .A1(\RI5[0][33] ), .A2(\RI5[0][27] ), .Z(
        \MC_ARK_ARC_1_0/temp1[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_26_0  ( .A1(\MC_ARK_ARC_1_0/temp4[35] ), .A2(
        \MC_ARK_ARC_1_0/temp3[35] ), .Z(\MC_ARK_ARC_1_0/temp6[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_26_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[71] ), 
        .A2(n199), .Z(\MC_ARK_ARC_1_0/temp4[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_26_0  ( .A1(\RI5[0][101] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[137] ), .Z(\MC_ARK_ARC_1_0/temp3[35] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_25_5  ( .A1(\MC_ARK_ARC_1_0/temp3[36] ), .A2(
        \MC_ARK_ARC_1_0/temp4[36] ), .Z(\MC_ARK_ARC_1_0/temp6[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_5  ( .A1(\RI5[0][72] ), .A2(n194), .Z(
        \MC_ARK_ARC_1_0/temp4[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_25_5  ( .A1(\RI5[0][6] ), .A2(\RI5[0][174] ), .Z(
        \MC_ARK_ARC_1_0/temp2[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_25_5  ( .A1(\RI5[0][36] ), .A2(\RI5[0][30] ), .Z(
        \MC_ARK_ARC_1_0/temp1[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_25_4  ( .A1(\MC_ARK_ARC_1_0/temp3[37] ), .A2(
        \MC_ARK_ARC_1_0/temp4[37] ), .Z(\MC_ARK_ARC_1_0/temp6[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_25_4  ( .A1(\MC_ARK_ARC_1_0/temp1[37] ), .A2(
        \MC_ARK_ARC_1_0/temp2[37] ), .Z(\MC_ARK_ARC_1_0/temp5[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_4  ( .A1(\RI5[0][73] ), .A2(n509), .Z(
        \MC_ARK_ARC_1_0/temp4[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_25_4  ( .A1(\RI5[0][7] ), .A2(\RI5[0][175] ), .Z(
        \MC_ARK_ARC_1_0/temp2[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_25_4  ( .A1(\RI5[0][37] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[31] ), .Z(\MC_ARK_ARC_1_0/temp1[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_25_2  ( .A1(\MC_ARK_ARC_1_0/temp5[39] ), .A2(
        \MC_ARK_ARC_1_0/temp6[39] ), .Z(\MC_ARK_ARC_1_0/buf_output[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_25_2  ( .A1(\MC_ARK_ARC_1_0/temp4[39] ), .A2(
        \MC_ARK_ARC_1_0/temp3[39] ), .Z(\MC_ARK_ARC_1_0/temp6[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[75] ), 
        .A2(n196), .Z(\MC_ARK_ARC_1_0/temp4[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_25_2  ( .A1(\RI5[0][105] ), .A2(\RI5[0][141] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_25_2  ( .A1(\RI5[0][9] ), .A2(\RI5[0][177] ), .Z(
        \MC_ARK_ARC_1_0/temp2[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_25_1  ( .A1(\MC_ARK_ARC_1_0/temp3[40] ), .A2(
        \MC_ARK_ARC_1_0/temp4[40] ), .Z(\MC_ARK_ARC_1_0/temp6[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_1  ( .A1(\RI5[0][76] ), .A2(n73), .Z(
        \MC_ARK_ARC_1_0/temp4[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_25_1  ( .A1(\RI5[0][10] ), .A2(\RI5[0][178] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[77] ), 
        .A2(n213), .Z(\MC_ARK_ARC_1_0/temp4[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_25_0  ( .A1(\RI5[0][143] ), .A2(\RI5[0][107] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_25_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[35] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[41] ), .Z(\MC_ARK_ARC_1_0/temp1[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_5  ( .A1(\RI5[0][78] ), .A2(n65), .Z(
        \MC_ARK_ARC_1_0/temp4[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_24_5  ( .A1(\RI5[0][144] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[108] ), .Z(\MC_ARK_ARC_1_0/temp3[42] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_24_5  ( .A1(\RI5[0][12] ), .A2(\RI5[0][180] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_24_5  ( .A1(\RI5[0][36] ), .A2(\RI5[0][42] ), .Z(
        \MC_ARK_ARC_1_0/temp1[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_24_4  ( .A1(\MC_ARK_ARC_1_0/temp5[43] ), .A2(
        \MC_ARK_ARC_1_0/temp6[43] ), .Z(\MC_ARK_ARC_1_0/buf_output[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_4  ( .A1(\RI5[0][79] ), .A2(n478), .Z(
        \MC_ARK_ARC_1_0/temp4[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_3  ( .A1(\RI5[0][80] ), .A2(n471), .Z(
        \MC_ARK_ARC_1_0/temp4[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_24_2  ( .A1(\MC_ARK_ARC_1_0/temp3[45] ), .A2(
        \MC_ARK_ARC_1_0/temp4[45] ), .Z(\MC_ARK_ARC_1_0/temp6[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_2  ( .A1(\RI5[0][81] ), .A2(n465), .Z(
        \MC_ARK_ARC_1_0/temp4[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_1  ( .A1(\RI5[0][82] ), .A2(n129), .Z(
        \MC_ARK_ARC_1_0/temp4[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_24_1  ( .A1(\RI5[0][148] ), .A2(\RI5[0][112] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_24_1  ( .A1(\RI5[0][46] ), .A2(\RI5[0][40] ), .Z(
        \MC_ARK_ARC_1_0/temp1[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_23_5  ( .A1(\MC_ARK_ARC_1_0/temp5[48] ), .A2(
        \MC_ARK_ARC_1_0/temp6[48] ), .Z(\MC_ARK_ARC_1_0/buf_output[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_23_5  ( .A1(\MC_ARK_ARC_1_0/temp3[48] ), .A2(
        \MC_ARK_ARC_1_0/temp4[48] ), .Z(\MC_ARK_ARC_1_0/temp6[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_5  ( .A1(\SB2_0_22/buf_output[0] ), .A2(n450), 
        .Z(\MC_ARK_ARC_1_0/temp4[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_23_5  ( .A1(\RI5[0][114] ), .A2(\RI5[0][150] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_23_5  ( .A1(\RI5[0][18] ), .A2(\RI5[0][186] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_23_5  ( .A1(\RI5[0][48] ), .A2(\RI5[0][42] ), .Z(
        \MC_ARK_ARC_1_0/temp1[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_23_4  ( .A1(\MC_ARK_ARC_1_0/temp3[49] ), .A2(
        \MC_ARK_ARC_1_0/temp4[49] ), .Z(\MC_ARK_ARC_1_0/temp6[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_4  ( .A1(\RI5[0][85] ), .A2(n82), .Z(
        \MC_ARK_ARC_1_0/temp4[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_23_4  ( .A1(\RI5[0][19] ), .A2(\RI5[0][187] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_23_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .A2(\RI5[0][49] ), .Z(\MC_ARK_ARC_1_0/temp1[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_3  ( .A1(\RI5[0][86] ), .A2(n96), .Z(
        \MC_ARK_ARC_1_0/temp4[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_2  ( .A1(\RI5[0][87] ), .A2(n430), .Z(
        \MC_ARK_ARC_1_0/temp4[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_1  ( .A1(\RI5[0][88] ), .A2(n180), .Z(
        \MC_ARK_ARC_1_0/temp4[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_23_1  ( .A1(\RI5[0][154] ), .A2(\RI5[0][118] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_23_1  ( .A1(\RI5[0][190] ), .A2(\RI5[0][22] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_0  ( .A1(\RI5[0][89] ), .A2(n195), .Z(
        \MC_ARK_ARC_1_0/temp4[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_23_0  ( .A1(\RI5[0][119] ), .A2(\RI5[0][155] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_23_0  ( .A1(\RI5[0][47] ), .A2(\RI5[0][53] ), .Z(
        \MC_ARK_ARC_1_0/temp1[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_22_5  ( .A1(\MC_ARK_ARC_1_0/temp2[54] ), .A2(
        \MC_ARK_ARC_1_0/temp1[54] ), .Z(\MC_ARK_ARC_1_0/temp5[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_5  ( .A1(\RI5[0][90] ), .A2(n174), .Z(
        \MC_ARK_ARC_1_0/temp4[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_22_5  ( .A1(\RI5[0][54] ), .A2(\RI5[0][48] ), .Z(
        \MC_ARK_ARC_1_0/temp1[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_4  ( .A1(\RI5[0][91] ), .A2(n46), .Z(
        \MC_ARK_ARC_1_0/temp4[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_22_4  ( .A1(\RI5[0][55] ), .A2(\RI5[0][49] ), .Z(
        \MC_ARK_ARC_1_0/temp1[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_2  ( .A1(\SB2_0_18/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_0/buf_keyinput[57] ), .Z(\MC_ARK_ARC_1_0/temp4[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_22_1  ( .A1(\MC_ARK_ARC_1_0/temp5[58] ), .A2(
        \MC_ARK_ARC_1_0/temp6[58] ), .Z(\MC_ARK_ARC_1_0/buf_output[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_22_1  ( .A1(\MC_ARK_ARC_1_0/temp3[58] ), .A2(
        \MC_ARK_ARC_1_0/temp4[58] ), .Z(\MC_ARK_ARC_1_0/temp6[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_22_1  ( .A1(\MC_ARK_ARC_1_0/temp2[58] ), .A2(
        \MC_ARK_ARC_1_0/temp1[58] ), .Z(\MC_ARK_ARC_1_0/temp5[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_1  ( .A1(\RI5[0][94] ), .A2(n546), .Z(
        \MC_ARK_ARC_1_0/temp4[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_22_1  ( .A1(\RI5[0][160] ), .A2(\RI5[0][124] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_22_1  ( .A1(\RI5[0][4] ), .A2(\RI5[0][28] ), .Z(
        \MC_ARK_ARC_1_0/temp2[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_22_1  ( .A1(\RI5[0][58] ), .A2(\RI5[0][52] ), .Z(
        \MC_ARK_ARC_1_0/temp1[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_21_5  ( .A1(\MC_ARK_ARC_1_0/temp4[60] ), .A2(
        \MC_ARK_ARC_1_0/temp3[60] ), .Z(\MC_ARK_ARC_1_0/temp6[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_21_5  ( .A1(\RI5[0][96] ), .A2(n77), .Z(
        \MC_ARK_ARC_1_0/temp4[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_21_5  ( .A1(\RI5[0][6] ), .A2(\RI5[0][30] ), .Z(
        \MC_ARK_ARC_1_0/temp2[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_21_5  ( .A1(\RI5[0][60] ), .A2(\RI5[0][54] ), .Z(
        \MC_ARK_ARC_1_0/temp1[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_21_4  ( .A1(\MC_ARK_ARC_1_0/temp6[61] ), .A2(
        \MC_ARK_ARC_1_0/temp5[61] ), .Z(\MC_ARK_ARC_1_0/buf_output[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_21_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[97] ), 
        .A2(n531), .Z(\MC_ARK_ARC_1_0/temp4[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_21_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .A2(\RI5[0][7] ), .Z(\MC_ARK_ARC_1_0/temp2[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_21_3  ( .A1(\MC_ARK_ARC_1_0/temp4[62] ), .A2(
        \MC_ARK_ARC_1_0/temp3[62] ), .Z(\MC_ARK_ARC_1_0/temp6[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_21_3  ( .A1(\MC_ARK_ARC_1_0/temp1[62] ), .A2(
        \MC_ARK_ARC_1_0/temp2[62] ), .Z(\MC_ARK_ARC_1_0/temp5[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_21_3  ( .A1(\RI5[0][98] ), .A2(n197), .Z(
        \MC_ARK_ARC_1_0/temp4[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_21_3  ( .A1(\RI5[0][128] ), .A2(\RI5[0][164] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_21_3  ( .A1(\RI5[0][32] ), .A2(\RI5[0][8] ), .Z(
        \MC_ARK_ARC_1_0/temp2[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_21_3  ( .A1(\RI5[0][56] ), .A2(\RI5[0][62] ), .Z(
        \MC_ARK_ARC_1_0/temp1[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_21_2  ( .A1(\SB2_0_17/buf_output[3] ), .A2(n127), 
        .Z(\MC_ARK_ARC_1_0/temp4[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_21_1  ( .A1(\RI5[0][100] ), .A2(n151), .Z(
        \MC_ARK_ARC_1_0/temp4[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_21_1  ( .A1(\RI5[0][166] ), .A2(\RI5[0][130] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .A2(n501), .Z(\MC_ARK_ARC_1_0/temp4[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_20_5  ( .A1(\RI5[0][168] ), .A2(\RI5[0][132] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_4  ( .A1(\RI5[0][103] ), .A2(n25), .Z(
        \MC_ARK_ARC_1_0/temp4[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_20_4  ( .A1(\RI5[0][133] ), .A2(\RI5[0][169] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_20_4  ( .A1(\RI5[0][37] ), .A2(\RI5[0][13] ), .Z(
        \MC_ARK_ARC_1_0/temp2[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_20_4  ( .A1(\RI5[0][61] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[67] ), .Z(\MC_ARK_ARC_1_0/temp1[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_3  ( .A1(\SB2_0_17/buf_output[2] ), .A2(n168), 
        .Z(\MC_ARK_ARC_1_0/temp4[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_20_3  ( .A1(\RI5[0][134] ), .A2(\RI5[0][170] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_20_2  ( .A1(\MC_ARK_ARC_1_0/temp1[69] ), .A2(
        \MC_ARK_ARC_1_0/temp2[69] ), .Z(\MC_ARK_ARC_1_0/temp5[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_2  ( .A1(\RI5[0][105] ), .A2(n175), .Z(
        \MC_ARK_ARC_1_0/temp4[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_20_2  ( .A1(\RI5[0][135] ), .A2(\RI5[0][171] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_20_2  ( .A1(\RI5[0][15] ), .A2(\RI5[0][39] ), .Z(
        \MC_ARK_ARC_1_0/temp2[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_20_2  ( .A1(\RI5[0][69] ), .A2(\RI5[0][63] ), .Z(
        \MC_ARK_ARC_1_0/temp1[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_20_1  ( .A1(\MC_ARK_ARC_1_0/temp6[70] ), .A2(
        \MC_ARK_ARC_1_0/temp5[70] ), .Z(\MC_ARK_ARC_1_0/buf_output[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_20_1  ( .A1(\MC_ARK_ARC_1_0/temp3[70] ), .A2(
        \MC_ARK_ARC_1_0/temp4[70] ), .Z(\MC_ARK_ARC_1_0/temp6[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_20_1  ( .A1(\MC_ARK_ARC_1_0/temp1[70] ), .A2(
        \MC_ARK_ARC_1_0/temp2[70] ), .Z(\MC_ARK_ARC_1_0/temp5[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_1  ( .A1(\RI5[0][106] ), .A2(n481), .Z(
        \MC_ARK_ARC_1_0/temp4[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_20_1  ( .A1(\RI5[0][172] ), .A2(\RI5[0][136] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_20_1  ( .A1(\RI5[0][16] ), .A2(\RI5[0][40] ), .Z(
        \MC_ARK_ARC_1_0/temp2[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_20_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[70] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[64] ), .Z(\MC_ARK_ARC_1_0/temp1[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_20_0  ( .A1(\MC_ARK_ARC_1_0/temp1[71] ), .A2(
        \MC_ARK_ARC_1_0/temp2[71] ), .Z(\MC_ARK_ARC_1_0/temp5[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_0  ( .A1(\RI5[0][107] ), .A2(
        \MC_ARK_ARC_1_0/buf_keyinput[71] ), .Z(\MC_ARK_ARC_1_0/temp4[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_20_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[41] ), 
        .A2(\RI5[0][17] ), .Z(\MC_ARK_ARC_1_0/temp2[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_19_5  ( .A1(\MC_ARK_ARC_1_0/temp6[72] ), .A2(
        \MC_ARK_ARC_1_0/temp5[72] ), .Z(\MC_ARK_ARC_1_0/buf_output[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_19_5  ( .A1(\MC_ARK_ARC_1_0/temp3[72] ), .A2(
        \MC_ARK_ARC_1_0/temp4[72] ), .Z(\MC_ARK_ARC_1_0/temp6[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[108] ), 
        .A2(n467), .Z(\MC_ARK_ARC_1_0/temp4[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_19_5  ( .A1(\RI5[0][174] ), .A2(\RI5[0][138] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_19_5  ( .A1(\RI5[0][42] ), .A2(\RI5[0][18] ), .Z(
        \MC_ARK_ARC_1_0/temp2[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_19_5  ( .A1(\RI5[0][72] ), .A2(\RI5[0][66] ), .Z(
        \MC_ARK_ARC_1_0/temp1[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_19_4  ( .A1(\MC_ARK_ARC_1_0/temp2[73] ), .A2(
        \MC_ARK_ARC_1_0/temp1[73] ), .Z(\MC_ARK_ARC_1_0/temp5[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_4  ( .A1(\RI5[0][109] ), .A2(n462), .Z(
        \MC_ARK_ARC_1_0/temp4[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_19_4  ( .A1(\RI5[0][175] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[139] ), .Z(\MC_ARK_ARC_1_0/temp3[73] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_19_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .A2(\RI5[0][19] ), .Z(\MC_ARK_ARC_1_0/temp2[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_19_4  ( .A1(\RI5[0][73] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[67] ), .Z(\MC_ARK_ARC_1_0/temp1[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_3  ( .A1(\RI5[0][110] ), .A2(n100), .Z(
        \MC_ARK_ARC_1_0/temp4[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_19_3  ( .A1(\RI5[0][74] ), .A2(\RI5[0][68] ), .Z(
        \MC_ARK_ARC_1_0/temp1[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_2  ( .A1(\RI5[0][111] ), .A2(n137), .Z(
        \MC_ARK_ARC_1_0/temp4[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_19_1  ( .A1(\MC_ARK_ARC_1_0/temp6[76] ), .A2(
        \MC_ARK_ARC_1_0/temp5[76] ), .Z(\MC_ARK_ARC_1_0/buf_output[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_19_1  ( .A1(\MC_ARK_ARC_1_0/temp3[76] ), .A2(
        \MC_ARK_ARC_1_0/temp4[76] ), .Z(\MC_ARK_ARC_1_0/temp6[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_19_1  ( .A1(\MC_ARK_ARC_1_0/temp2[76] ), .A2(
        \MC_ARK_ARC_1_0/temp1[76] ), .Z(\MC_ARK_ARC_1_0/temp5[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_1  ( .A1(\RI5[0][112] ), .A2(n446), .Z(
        \MC_ARK_ARC_1_0/temp4[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_19_1  ( .A1(\RI5[0][46] ), .A2(\RI5[0][22] ), .Z(
        \MC_ARK_ARC_1_0/temp2[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_19_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[70] ), 
        .A2(\RI5[0][76] ), .Z(\MC_ARK_ARC_1_0/temp1[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_19_0  ( .A1(\MC_ARK_ARC_1_0/temp3[77] ), .A2(
        \MC_ARK_ARC_1_0/temp4[77] ), .Z(\MC_ARK_ARC_1_0/temp6[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_19_0  ( .A1(\MC_ARK_ARC_1_0/temp1[77] ), .A2(
        \MC_ARK_ARC_1_0/temp2[77] ), .Z(\MC_ARK_ARC_1_0/temp5[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[113] ), 
        .A2(n440), .Z(\MC_ARK_ARC_1_0/temp4[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_19_0  ( .A1(\RI5[0][143] ), .A2(\RI5[0][179] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_19_0  ( .A1(\RI5[0][47] ), .A2(\RI5[0][23] ), .Z(
        \MC_ARK_ARC_1_0/temp2[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_18_5  ( .A1(\MC_ARK_ARC_1_0/temp3[78] ), .A2(
        \MC_ARK_ARC_1_0/temp4[78] ), .Z(\MC_ARK_ARC_1_0/temp6[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_5  ( .A1(\RI5[0][114] ), .A2(n433), .Z(
        \MC_ARK_ARC_1_0/temp4[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_18_5  ( .A1(\RI5[0][144] ), .A2(\RI5[0][180] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_18_5  ( .A1(\RI5[0][78] ), .A2(\RI5[0][72] ), .Z(
        \MC_ARK_ARC_1_0/temp1[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_4  ( .A1(\RI5[0][115] ), .A2(n39), .Z(
        \MC_ARK_ARC_1_0/temp4[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_18_4  ( .A1(\RI5[0][49] ), .A2(\RI5[0][25] ), .Z(
        \MC_ARK_ARC_1_0/temp2[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_18_4  ( .A1(\RI5[0][73] ), .A2(\RI5[0][79] ), .Z(
        \MC_ARK_ARC_1_0/temp1[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_3  ( .A1(\SB2_0_15/buf_output[2] ), .A2(n118), 
        .Z(\MC_ARK_ARC_1_0/temp4[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_18_3  ( .A1(\RI5[0][146] ), .A2(\RI5[0][182] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_2  ( .A1(\SB2_0_14/buf_output[3] ), .A2(n166), 
        .Z(\MC_ARK_ARC_1_0/temp4[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_18_2  ( .A1(\RI5[0][147] ), .A2(\RI5[0][183] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_18_2  ( .A1(\RI5[0][51] ), .A2(\RI5[0][27] ), .Z(
        \MC_ARK_ARC_1_0/temp2[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_18_1  ( .A1(\MC_ARK_ARC_1_0/temp3[82] ), .A2(
        \MC_ARK_ARC_1_0/temp4[82] ), .Z(\MC_ARK_ARC_1_0/temp6[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_1  ( .A1(\RI5[0][118] ), .A2(n169), .Z(
        \MC_ARK_ARC_1_0/temp4[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_18_1  ( .A1(\RI5[0][148] ), .A2(\RI5[0][184] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_18_1  ( .A1(\RI5[0][52] ), .A2(\RI5[0][28] ), .Z(
        \MC_ARK_ARC_1_0/temp2[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_18_1  ( .A1(\RI5[0][76] ), .A2(\RI5[0][82] ), .Z(
        \MC_ARK_ARC_1_0/temp1[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_18_0  ( .A1(\MC_ARK_ARC_1_0/temp5[83] ), .A2(
        \MC_ARK_ARC_1_0/temp6[83] ), .Z(\MC_ARK_ARC_1_0/buf_output[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_18_0  ( .A1(\MC_ARK_ARC_1_0/temp3[83] ), .A2(
        \MC_ARK_ARC_1_0/temp4[83] ), .Z(\MC_ARK_ARC_1_0/temp6[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_18_0  ( .A1(\MC_ARK_ARC_1_0/temp1[83] ), .A2(
        \MC_ARK_ARC_1_0/temp2[83] ), .Z(\MC_ARK_ARC_1_0/temp5[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_0  ( .A1(\RI5[0][119] ), .A2(n103), .Z(
        \MC_ARK_ARC_1_0/temp4[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_18_0  ( .A1(\RI5[0][185] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[149] ), .Z(\MC_ARK_ARC_1_0/temp3[83] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_18_0  ( .A1(\RI5[0][29] ), .A2(\RI5[0][53] ), .Z(
        \MC_ARK_ARC_1_0/temp2[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_17_5  ( .A1(\MC_ARK_ARC_1_0/temp6[84] ), .A2(
        \MC_ARK_ARC_1_0/temp5[84] ), .Z(\MC_ARK_ARC_1_0/buf_output[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_17_5  ( .A1(\MC_ARK_ARC_1_0/temp3[84] ), .A2(
        \MC_ARK_ARC_1_0/temp4[84] ), .Z(\MC_ARK_ARC_1_0/temp6[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_5  ( .A1(\RI5[0][120] ), .A2(n554), .Z(
        \MC_ARK_ARC_1_0/temp4[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_17_5  ( .A1(\RI5[0][186] ), .A2(\RI5[0][150] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_17_5  ( .A1(\RI5[0][54] ), .A2(\RI5[0][30] ), .Z(
        \MC_ARK_ARC_1_0/temp2[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_17_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[84] ), 
        .A2(\RI5[0][78] ), .Z(\MC_ARK_ARC_1_0/temp1[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_17_4  ( .A1(\MC_ARK_ARC_1_0/temp2[85] ), .A2(
        \MC_ARK_ARC_1_0/temp1[85] ), .Z(\MC_ARK_ARC_1_0/temp5[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_4  ( .A1(n7134), .A2(n549), .Z(
        \MC_ARK_ARC_1_0/temp4[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_17_4  ( .A1(\RI5[0][187] ), .A2(\RI5[0][151] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_17_4  ( .A1(\RI5[0][79] ), .A2(\RI5[0][85] ), .Z(
        \MC_ARK_ARC_1_0/temp1[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_3  ( .A1(\RI5[0][122] ), .A2(n543), .Z(
        \MC_ARK_ARC_1_0/temp4[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_17_3  ( .A1(\RI5[0][188] ), .A2(\RI5[0][152] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_17_2  ( .A1(\RI5[0][33] ), .A2(\RI5[0][57] ), .Z(
        \MC_ARK_ARC_1_0/temp2[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_1  ( .A1(\RI5[0][124] ), .A2(n534), .Z(
        \MC_ARK_ARC_1_0/temp4[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_17_1  ( .A1(\RI5[0][88] ), .A2(\RI5[0][82] ), .Z(
        \MC_ARK_ARC_1_0/temp1[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_5  ( .A1(\RI5[0][126] ), .A2(n144), .Z(
        \MC_ARK_ARC_1_0/temp4[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_16_5  ( .A1(\RI5[0][0] ), .A2(\RI5[0][156] ), .Z(
        \MC_ARK_ARC_1_0/temp3[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_16_5  ( .A1(\RI5[0][60] ), .A2(\RI5[0][36] ), .Z(
        \MC_ARK_ARC_1_0/temp2[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_16_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[84] ), 
        .A2(\RI5[0][90] ), .Z(\MC_ARK_ARC_1_0/temp1[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_16_4  ( .A1(\MC_ARK_ARC_1_0/temp6[91] ), .A2(
        \MC_ARK_ARC_1_0/temp5[91] ), .Z(\MC_ARK_ARC_1_0/buf_output[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_16_4  ( .A1(\MC_ARK_ARC_1_0/temp3[91] ), .A2(
        \MC_ARK_ARC_1_0/temp4[91] ), .Z(\MC_ARK_ARC_1_0/temp6[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_16_4  ( .A1(\MC_ARK_ARC_1_0/temp2[91] ), .A2(
        \MC_ARK_ARC_1_0/temp1[91] ), .Z(\MC_ARK_ARC_1_0/temp5[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_4  ( .A1(\RI5[0][127] ), .A2(n121), .Z(
        \MC_ARK_ARC_1_0/temp4[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_16_4  ( .A1(\RI5[0][1] ), .A2(\RI5[0][157] ), .Z(
        \MC_ARK_ARC_1_0/temp3[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_16_4  ( .A1(\RI5[0][37] ), .A2(\RI5[0][61] ), .Z(
        \MC_ARK_ARC_1_0/temp2[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_16_4  ( .A1(\RI5[0][91] ), .A2(\RI5[0][85] ), .Z(
        \MC_ARK_ARC_1_0/temp1[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_3  ( .A1(\RI5[0][128] ), .A2(
        \MC_ARK_ARC_1_0/buf_keyinput[92] ), .Z(\MC_ARK_ARC_1_0/temp4[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_2  ( .A1(\RI5[0][129] ), .A2(n207), .Z(
        \MC_ARK_ARC_1_0/temp4[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_16_2  ( .A1(\RI5[0][39] ), .A2(\RI5[0][63] ), .Z(
        \MC_ARK_ARC_1_0/temp2[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_1  ( .A1(\RI5[0][130] ), .A2(n75), .Z(
        \MC_ARK_ARC_1_0/temp4[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_16_1  ( .A1(\RI5[0][4] ), .A2(\RI5[0][160] ), .Z(
        \MC_ARK_ARC_1_0/temp3[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_16_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .A2(\RI5[0][40] ), .Z(\MC_ARK_ARC_1_0/temp2[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_16_1  ( .A1(\RI5[0][88] ), .A2(\RI5[0][94] ), .Z(
        \MC_ARK_ARC_1_0/temp1[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_0  ( .A1(\RI5[0][131] ), .A2(n21), .Z(
        \MC_ARK_ARC_1_0/temp4[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_15_5  ( .A1(\MC_ARK_ARC_1_0/temp1[96] ), .A2(
        \MC_ARK_ARC_1_0/temp2[96] ), .Z(\MC_ARK_ARC_1_0/temp5[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_5  ( .A1(\RI5[0][132] ), .A2(n212), .Z(
        \MC_ARK_ARC_1_0/temp4[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_15_5  ( .A1(\RI5[0][6] ), .A2(\RI5[0][162] ), .Z(
        \MC_ARK_ARC_1_0/temp3[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_15_5  ( .A1(\RI5[0][66] ), .A2(\RI5[0][42] ), .Z(
        \MC_ARK_ARC_1_0/temp2[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_15_5  ( .A1(\RI5[0][96] ), .A2(\RI5[0][90] ), .Z(
        \MC_ARK_ARC_1_0/temp1[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_15_4  ( .A1(\MC_ARK_ARC_1_0/temp2[97] ), .A2(
        \MC_ARK_ARC_1_0/temp1[97] ), .Z(\MC_ARK_ARC_1_0/temp5[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_4  ( .A1(\RI5[0][133] ), .A2(n484), .Z(
        \MC_ARK_ARC_1_0/temp4[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_15_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[67] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[43] ), .Z(\MC_ARK_ARC_1_0/temp2[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_3  ( .A1(\RI5[0][134] ), .A2(n477), .Z(
        \MC_ARK_ARC_1_0/temp4[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_2  ( .A1(\RI5[0][135] ), .A2(n470), .Z(
        \MC_ARK_ARC_1_0/temp4[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_15_1  ( .A1(\MC_ARK_ARC_1_0/temp3[100] ), .A2(
        \MC_ARK_ARC_1_0/temp4[100] ), .Z(\MC_ARK_ARC_1_0/temp6[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_1  ( .A1(\RI5[0][136] ), .A2(n63), .Z(
        \MC_ARK_ARC_1_0/temp4[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_15_1  ( .A1(\RI5[0][10] ), .A2(\RI5[0][166] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_15_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[70] ), 
        .A2(\RI5[0][46] ), .Z(\MC_ARK_ARC_1_0/temp2[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_15_1  ( .A1(\RI5[0][100] ), .A2(\RI5[0][94] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_15_0  ( .A1(\MC_ARK_ARC_1_0/temp5[101] ), .A2(
        \MC_ARK_ARC_1_0/temp6[101] ), .Z(\MC_ARK_ARC_1_0/buf_output[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_15_0  ( .A1(\MC_ARK_ARC_1_0/temp3[101] ), .A2(
        \MC_ARK_ARC_1_0/temp4[101] ), .Z(\MC_ARK_ARC_1_0/temp6[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_15_0  ( .A1(\MC_ARK_ARC_1_0/temp1[101] ), .A2(
        \MC_ARK_ARC_1_0/temp2[101] ), .Z(\MC_ARK_ARC_1_0/temp5[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[137] ), 
        .A2(n458), .Z(\MC_ARK_ARC_1_0/temp4[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_15_0  ( .A1(\RI5[0][95] ), .A2(\RI5[0][101] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_5  ( .A1(\SB2_0_13/buf_output[0] ), .A2(n209), 
        .Z(\MC_ARK_ARC_1_0/temp4[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_14_4  ( .A1(\MC_ARK_ARC_1_0/temp1[103] ), .A2(
        \MC_ARK_ARC_1_0/temp2[103] ), .Z(\MC_ARK_ARC_1_0/temp5[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[139] ), 
        .A2(n88), .Z(\MC_ARK_ARC_1_0/temp4[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_14_4  ( .A1(\RI5[0][13] ), .A2(\RI5[0][169] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_14_4  ( .A1(\RI5[0][73] ), .A2(\RI5[0][49] ), .Z(
        \MC_ARK_ARC_1_0/temp2[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_3  ( .A1(\RI5[0][140] ), .A2(n49), .Z(
        \MC_ARK_ARC_1_0/temp4[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_2  ( .A1(\RI5[0][141] ), .A2(n436), .Z(
        \MC_ARK_ARC_1_0/temp4[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_14_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[75] ), 
        .A2(\RI5[0][51] ), .Z(\MC_ARK_ARC_1_0/temp2[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_14_1  ( .A1(\MC_ARK_ARC_1_0/temp6[106] ), .A2(
        \MC_ARK_ARC_1_0/temp5[106] ), .Z(\MC_ARK_ARC_1_0/buf_output[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_14_1  ( .A1(\MC_ARK_ARC_1_0/temp3[106] ), .A2(
        \MC_ARK_ARC_1_0/temp4[106] ), .Z(\MC_ARK_ARC_1_0/temp6[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_14_1  ( .A1(\MC_ARK_ARC_1_0/temp1[106] ), .A2(
        \MC_ARK_ARC_1_0/temp2[106] ), .Z(\MC_ARK_ARC_1_0/temp5[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_1  ( .A1(\RI5[0][142] ), .A2(n58), .Z(
        \MC_ARK_ARC_1_0/temp4[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_14_1  ( .A1(\RI5[0][16] ), .A2(\RI5[0][172] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_14_1  ( .A1(\RI5[0][76] ), .A2(\RI5[0][52] ), .Z(
        \MC_ARK_ARC_1_0/temp2[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_0  ( .A1(\RI5[0][143] ), .A2(n423), .Z(
        \MC_ARK_ARC_1_0/temp4[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_13_5  ( .A1(\MC_ARK_ARC_1_0/temp3[108] ), .A2(
        \MC_ARK_ARC_1_0/temp4[108] ), .Z(\MC_ARK_ARC_1_0/temp6[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_5  ( .A1(\RI5[0][144] ), .A2(n187), .Z(
        \MC_ARK_ARC_1_0/temp4[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_13_5  ( .A1(\RI5[0][18] ), .A2(\RI5[0][174] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_13_5  ( .A1(\RI5[0][78] ), .A2(\RI5[0][54] ), .Z(
        \MC_ARK_ARC_1_0/temp2[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_13_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[108] ), .Z(
        \MC_ARK_ARC_1_0/temp1[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_4  ( .A1(\RI5[0][145] ), .A2(n37), .Z(
        \MC_ARK_ARC_1_0/temp4[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_13_4  ( .A1(\SB2_0_18/buf_output[1] ), .A2(
        \RI5[0][109] ), .Z(\MC_ARK_ARC_1_0/temp1[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_3  ( .A1(\RI5[0][146] ), .A2(n193), .Z(
        \MC_ARK_ARC_1_0/temp4[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_13_2  ( .A1(\MC_ARK_ARC_1_0/temp4[111] ), .A2(
        \MC_ARK_ARC_1_0/temp3[111] ), .Z(\MC_ARK_ARC_1_0/temp6[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_13_2  ( .A1(\MC_ARK_ARC_1_0/temp1[111] ), .A2(
        \MC_ARK_ARC_1_0/temp2[111] ), .Z(\MC_ARK_ARC_1_0/temp5[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_2  ( .A1(\RI5[0][147] ), .A2(n556), .Z(
        \MC_ARK_ARC_1_0/temp4[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_13_2  ( .A1(\RI5[0][21] ), .A2(\RI5[0][177] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_13_2  ( .A1(\RI5[0][81] ), .A2(\RI5[0][57] ), .Z(
        \MC_ARK_ARC_1_0/temp2[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_13_1  ( .A1(\MC_ARK_ARC_1_0/temp1[112] ), .A2(
        \MC_ARK_ARC_1_0/temp2[112] ), .Z(\MC_ARK_ARC_1_0/temp5[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_1  ( .A1(\RI5[0][148] ), .A2(n551), .Z(
        \MC_ARK_ARC_1_0/temp4[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_13_1  ( .A1(\SB2_0_23/buf_output[4] ), .A2(
        \RI5[0][82] ), .Z(\MC_ARK_ARC_1_0/temp2[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_13_1  ( .A1(\RI5[0][112] ), .A2(\RI5[0][106] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_13_0  ( .A1(\MC_ARK_ARC_1_0/temp3[113] ), .A2(
        \MC_ARK_ARC_1_0/temp4[113] ), .Z(\MC_ARK_ARC_1_0/temp6[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[149] ), 
        .A2(n220), .Z(\MC_ARK_ARC_1_0/temp4[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_12_5  ( .A1(\MC_ARK_ARC_1_0/temp5[114] ), .A2(
        \MC_ARK_ARC_1_0/temp6[114] ), .Z(\MC_ARK_ARC_1_0/buf_output[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_12_5  ( .A1(\MC_ARK_ARC_1_0/temp3[114] ), .A2(
        \MC_ARK_ARC_1_0/temp4[114] ), .Z(\MC_ARK_ARC_1_0/temp6[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_12_5  ( .A1(\MC_ARK_ARC_1_0/temp2[114] ), .A2(
        \MC_ARK_ARC_1_0/temp1[114] ), .Z(\MC_ARK_ARC_1_0/temp5[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_5  ( .A1(\RI5[0][150] ), .A2(n123), .Z(
        \MC_ARK_ARC_1_0/temp4[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_12_5  ( .A1(\RI5[0][24] ), .A2(\RI5[0][180] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_12_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[84] ), 
        .A2(\RI5[0][60] ), .Z(\MC_ARK_ARC_1_0/temp2[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_12_4  ( .A1(\MC_ARK_ARC_1_0/temp3[115] ), .A2(
        \MC_ARK_ARC_1_0/temp4[115] ), .Z(\MC_ARK_ARC_1_0/temp6[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_12_4  ( .A1(\MC_ARK_ARC_1_0/temp1[115] ), .A2(
        \MC_ARK_ARC_1_0/temp2[115] ), .Z(\MC_ARK_ARC_1_0/temp5[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_4  ( .A1(\RI5[0][151] ), .A2(n536), .Z(
        \MC_ARK_ARC_1_0/temp4[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_12_4  ( .A1(\RI5[0][25] ), .A2(\RI5[0][181] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_12_4  ( .A1(\RI5[0][85] ), .A2(\RI5[0][61] ), .Z(
        \MC_ARK_ARC_1_0/temp2[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_12_4  ( .A1(\RI5[0][115] ), .A2(\RI5[0][109] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_12_3  ( .A1(\MC_ARK_ARC_1_0/temp1[116] ), .A2(
        \MC_ARK_ARC_1_0/temp2[116] ), .Z(\MC_ARK_ARC_1_0/temp5[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_3  ( .A1(\RI5[0][152] ), .A2(n530), .Z(
        \MC_ARK_ARC_1_0/temp4[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_12_3  ( .A1(\RI5[0][62] ), .A2(\RI5[0][86] ), .Z(
        \MC_ARK_ARC_1_0/temp2[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_2  ( .A1(\RI5[0][153] ), .A2(n154), .Z(
        \MC_ARK_ARC_1_0/temp4[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_12_1  ( .A1(\MC_ARK_ARC_1_0/temp5[118] ), .A2(
        \MC_ARK_ARC_1_0/temp6[118] ), .Z(\MC_ARK_ARC_1_0/buf_output[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_12_1  ( .A1(\MC_ARK_ARC_1_0/temp3[118] ), .A2(
        \MC_ARK_ARC_1_0/temp4[118] ), .Z(\MC_ARK_ARC_1_0/temp6[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_12_1  ( .A1(\MC_ARK_ARC_1_0/temp2[118] ), .A2(
        \MC_ARK_ARC_1_0/temp1[118] ), .Z(\MC_ARK_ARC_1_0/temp5[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_1  ( .A1(\SB2_0_7/buf_output[4] ), .A2(n110), 
        .Z(\MC_ARK_ARC_1_0/temp4[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_12_1  ( .A1(\RI5[0][28] ), .A2(\RI5[0][184] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_12_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .A2(\RI5[0][88] ), .Z(\MC_ARK_ARC_1_0/temp2[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_12_1  ( .A1(\RI5[0][118] ), .A2(\RI5[0][112] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_12_0  ( .A1(\MC_ARK_ARC_1_0/temp3[119] ), .A2(
        \MC_ARK_ARC_1_0/temp4[119] ), .Z(\MC_ARK_ARC_1_0/temp6[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_12_0  ( .A1(\MC_ARK_ARC_1_0/temp2[119] ), .A2(
        \MC_ARK_ARC_1_0/temp1[119] ), .Z(\MC_ARK_ARC_1_0/temp5[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_0  ( .A1(\RI5[0][155] ), .A2(n106), .Z(
        \MC_ARK_ARC_1_0/temp4[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_12_0  ( .A1(\RI5[0][89] ), .A2(\RI5[0][65] ), .Z(
        \MC_ARK_ARC_1_0/temp2[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_12_0  ( .A1(\RI5[0][119] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[113] ), .Z(\MC_ARK_ARC_1_0/temp1[119] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_11_5  ( .A1(\MC_ARK_ARC_1_0/temp5[120] ), .A2(
        \MC_ARK_ARC_1_0/temp6[120] ), .Z(\MC_ARK_ARC_1_0/buf_output[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_11_5  ( .A1(\MC_ARK_ARC_1_0/temp1[120] ), .A2(
        \MC_ARK_ARC_1_0/temp2[120] ), .Z(\MC_ARK_ARC_1_0/temp5[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_5  ( .A1(\RI5[0][156] ), .A2(n506), .Z(
        \MC_ARK_ARC_1_0/temp4[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_11_5  ( .A1(\RI5[0][30] ), .A2(\RI5[0][186] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_11_5  ( .A1(\RI5[0][90] ), .A2(\RI5[0][66] ), .Z(
        \MC_ARK_ARC_1_0/temp2[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_11_5  ( .A1(\RI5[0][120] ), .A2(\RI5[0][114] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_11_4  ( .A1(\MC_ARK_ARC_1_0/temp5[121] ), .A2(
        \MC_ARK_ARC_1_0/temp6[121] ), .Z(\MC_ARK_ARC_1_0/buf_output[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_11_4  ( .A1(\MC_ARK_ARC_1_0/temp3[121] ), .A2(
        \MC_ARK_ARC_1_0/temp4[121] ), .Z(\MC_ARK_ARC_1_0/temp6[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_11_4  ( .A1(\MC_ARK_ARC_1_0/temp1[121] ), .A2(
        \MC_ARK_ARC_1_0/temp2[121] ), .Z(\MC_ARK_ARC_1_0/temp5[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_4  ( .A1(\RI5[0][157] ), .A2(n500), .Z(
        \MC_ARK_ARC_1_0/temp4[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_11_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .A2(\RI5[0][187] ), .Z(\MC_ARK_ARC_1_0/temp3[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_11_4  ( .A1(\RI5[0][91] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[67] ), .Z(\MC_ARK_ARC_1_0/temp2[121] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_11_4  ( .A1(n7134), .A2(\RI5[0][115] ), .Z(
        \MC_ARK_ARC_1_0/temp1[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_3  ( .A1(\RI5[0][158] ), .A2(n192), .Z(
        \MC_ARK_ARC_1_0/temp4[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_11_3  ( .A1(\RI5[0][68] ), .A2(\RI5[0][92] ), .Z(
        \MC_ARK_ARC_1_0/temp2[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_2  ( .A1(\RI5[0][159] ), .A2(n4), .Z(
        \MC_ARK_ARC_1_0/temp4[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_11_2  ( .A1(\RI5[0][33] ), .A2(\RI5[0][189] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_11_1  ( .A1(\MC_ARK_ARC_1_0/temp6[124] ), .A2(
        \MC_ARK_ARC_1_0/temp5[124] ), .Z(\MC_ARK_ARC_1_0/buf_output[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_11_1  ( .A1(\MC_ARK_ARC_1_0/temp3[124] ), .A2(
        \MC_ARK_ARC_1_0/temp4[124] ), .Z(\MC_ARK_ARC_1_0/temp6[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_1  ( .A1(\RI5[0][160] ), .A2(n486), .Z(
        \MC_ARK_ARC_1_0/temp4[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_11_1  ( .A1(\RI5[0][34] ), .A2(\RI5[0][190] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_11_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[70] ), 
        .A2(\RI5[0][94] ), .Z(\MC_ARK_ARC_1_0/temp2[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_0  ( .A1(\RI5[0][161] ), .A2(n69), .Z(
        \MC_ARK_ARC_1_0/temp4[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_11_0  ( .A1(\RI5[0][125] ), .A2(\RI5[0][119] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_10_5  ( .A1(\MC_ARK_ARC_1_0/temp3[126] ), .A2(
        \MC_ARK_ARC_1_0/temp4[126] ), .Z(\MC_ARK_ARC_1_0/temp6[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_5  ( .A1(\RI5[0][162] ), .A2(n159), .Z(
        \MC_ARK_ARC_1_0/temp4[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_10_5  ( .A1(\RI5[0][0] ), .A2(\RI5[0][36] ), .Z(
        \MC_ARK_ARC_1_0/temp3[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_10_5  ( .A1(\RI5[0][96] ), .A2(\RI5[0][72] ), .Z(
        \MC_ARK_ARC_1_0/temp2[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_4  ( .A1(\RI5[0][163] ), .A2(n139), .Z(
        \MC_ARK_ARC_1_0/temp4[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_10_4  ( .A1(\RI5[0][37] ), .A2(\RI5[0][1] ), .Z(
        \MC_ARK_ARC_1_0/temp3[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_10_4  ( .A1(n7134), .A2(\RI5[0][127] ), .Z(
        \MC_ARK_ARC_1_0/temp1[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_3  ( .A1(\RI5[0][164] ), .A2(n461), .Z(
        \MC_ARK_ARC_1_0/temp4[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_10_3  ( .A1(\RI5[0][38] ), .A2(\RI5[0][2] ), .Z(
        \MC_ARK_ARC_1_0/temp3[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_10_3  ( .A1(\RI5[0][122] ), .A2(\RI5[0][128] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_10_2  ( .A1(\MC_ARK_ARC_1_0/temp5[129] ), .A2(
        \MC_ARK_ARC_1_0/temp6[129] ), .Z(\MC_ARK_ARC_1_0/buf_output[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_10_2  ( .A1(\MC_ARK_ARC_1_0/temp3[129] ), .A2(
        \MC_ARK_ARC_1_0/temp4[129] ), .Z(\MC_ARK_ARC_1_0/temp6[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_2  ( .A1(\RI5[0][165] ), .A2(n455), .Z(
        \MC_ARK_ARC_1_0/temp4[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_10_2  ( .A1(\RI5[0][39] ), .A2(\RI5[0][3] ), .Z(
        \MC_ARK_ARC_1_0/temp3[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_10_2  ( .A1(\RI5[0][123] ), .A2(\RI5[0][129] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_10_1  ( .A1(\MC_ARK_ARC_1_0/temp5[130] ), .A2(
        \MC_ARK_ARC_1_0/temp6[130] ), .Z(\MC_ARK_ARC_1_0/buf_output[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_10_1  ( .A1(\MC_ARK_ARC_1_0/temp2[130] ), .A2(
        \MC_ARK_ARC_1_0/temp1[130] ), .Z(\MC_ARK_ARC_1_0/temp5[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_1  ( .A1(\RI5[0][166] ), .A2(n206), .Z(
        \MC_ARK_ARC_1_0/temp4[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_10_1  ( .A1(\RI5[0][4] ), .A2(\RI5[0][40] ), .Z(
        \MC_ARK_ARC_1_0/temp3[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_10_1  ( .A1(\RI5[0][130] ), .A2(\RI5[0][124] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_0  ( .A1(\RI5[0][167] ), .A2(n211), .Z(
        \MC_ARK_ARC_1_0/temp4[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_10_0  ( .A1(\RI5[0][125] ), .A2(\RI5[0][131] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_5  ( .A1(\RI5[0][168] ), .A2(n439), .Z(
        \MC_ARK_ARC_1_0/temp4[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_9_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .A2(\RI5[0][78] ), .Z(\MC_ARK_ARC_1_0/temp2[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_9_4  ( .A1(\MC_ARK_ARC_1_0/temp5[133] ), .A2(
        \MC_ARK_ARC_1_0/temp6[133] ), .Z(\MC_ARK_ARC_1_0/buf_output[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_9_4  ( .A1(\MC_ARK_ARC_1_0/temp3[133] ), .A2(
        \MC_ARK_ARC_1_0/temp4[133] ), .Z(\MC_ARK_ARC_1_0/temp6[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_4  ( .A1(\RI5[0][169] ), .A2(n119), .Z(
        \MC_ARK_ARC_1_0/temp4[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_9_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .A2(\RI5[0][7] ), .Z(\MC_ARK_ARC_1_0/temp3[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_9_4  ( .A1(\RI5[0][133] ), .A2(\RI5[0][127] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_9_2  ( .A1(\MC_ARK_ARC_1_0/temp3[135] ), .A2(
        \MC_ARK_ARC_1_0/temp4[135] ), .Z(\MC_ARK_ARC_1_0/temp6[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_2  ( .A1(\RI5[0][171] ), .A2(n420), .Z(
        \MC_ARK_ARC_1_0/temp4[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_1  ( .A1(\RI5[0][172] ), .A2(n47), .Z(
        \MC_ARK_ARC_1_0/temp4[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_9_1  ( .A1(\RI5[0][10] ), .A2(\RI5[0][46] ), .Z(
        \MC_ARK_ARC_1_0/temp3[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_9_1  ( .A1(\RI5[0][106] ), .A2(\RI5[0][82] ), .Z(
        \MC_ARK_ARC_1_0/temp2[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_9_1  ( .A1(\RI5[0][136] ), .A2(\RI5[0][130] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_9_0  ( .A1(\MC_ARK_ARC_1_0/temp3[137] ), .A2(
        \MC_ARK_ARC_1_0/temp4[137] ), .Z(\MC_ARK_ARC_1_0/temp6[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[173] ), 
        .A2(n173), .Z(\MC_ARK_ARC_1_0/temp4[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_9_0  ( .A1(\RI5[0][83] ), .A2(\RI5[0][107] ), .Z(
        \MC_ARK_ARC_1_0/temp2[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_5  ( .A1(\RI5[0][174] ), .A2(n163), .Z(
        \MC_ARK_ARC_1_0/temp4[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_8_5  ( .A1(\RI5[0][12] ), .A2(\RI5[0][48] ), .Z(
        \MC_ARK_ARC_1_0/temp3[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_8_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[84] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[108] ), .Z(
        \MC_ARK_ARC_1_0/temp2[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_8_5  ( .A1(\RI5[0][138] ), .A2(\RI5[0][132] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_8_4  ( .A1(\MC_ARK_ARC_1_0/temp3[139] ), .A2(
        \MC_ARK_ARC_1_0/temp4[139] ), .Z(\MC_ARK_ARC_1_0/temp6[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_4  ( .A1(\RI5[0][175] ), .A2(n553), .Z(
        \MC_ARK_ARC_1_0/temp4[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_8_4  ( .A1(\RI5[0][49] ), .A2(\RI5[0][13] ), .Z(
        \MC_ARK_ARC_1_0/temp3[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_8_4  ( .A1(\RI5[0][109] ), .A2(\RI5[0][85] ), .Z(
        \MC_ARK_ARC_1_0/temp2[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_3  ( .A1(\SB2_0_5/buf_output[2] ), .A2(n146), 
        .Z(\MC_ARK_ARC_1_0/temp4[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_2  ( .A1(\RI5[0][177] ), .A2(n130), .Z(
        \MC_ARK_ARC_1_0/temp4[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_8_1  ( .A1(\MC_ARK_ARC_1_0/temp5[142] ), .A2(
        \MC_ARK_ARC_1_0/temp6[142] ), .Z(\MC_ARK_ARC_1_0/buf_output[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_1  ( .A1(\SB2_0_3/buf_output[4] ), .A2(n210), 
        .Z(\MC_ARK_ARC_1_0/temp4[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_0  ( .A1(\RI5[0][179] ), .A2(n181), .Z(
        \MC_ARK_ARC_1_0/temp4[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_8_0  ( .A1(\RI5[0][143] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[137] ), .Z(\MC_ARK_ARC_1_0/temp1[143] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_7_5  ( .A1(\MC_ARK_ARC_1_0/temp5[144] ), .A2(
        \MC_ARK_ARC_1_0/temp6[144] ), .Z(\MC_ARK_ARC_1_0/buf_output[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_7_5  ( .A1(\MC_ARK_ARC_1_0/temp3[144] ), .A2(
        \MC_ARK_ARC_1_0/temp4[144] ), .Z(\MC_ARK_ARC_1_0/temp6[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_7_5  ( .A1(\MC_ARK_ARC_1_0/temp1[144] ), .A2(
        \MC_ARK_ARC_1_0/temp2[144] ), .Z(\MC_ARK_ARC_1_0/temp5[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_5  ( .A1(\RI5[0][180] ), .A2(n526), .Z(
        \MC_ARK_ARC_1_0/temp4[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_7_5  ( .A1(\RI5[0][54] ), .A2(\RI5[0][18] ), .Z(
        \MC_ARK_ARC_1_0/temp3[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_7_5  ( .A1(\RI5[0][138] ), .A2(\RI5[0][144] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_7_4  ( .A1(\MC_ARK_ARC_1_0/temp6[145] ), .A2(
        \MC_ARK_ARC_1_0/temp5[145] ), .Z(\MC_ARK_ARC_1_0/buf_output[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_7_4  ( .A1(\MC_ARK_ARC_1_0/temp3[145] ), .A2(
        \MC_ARK_ARC_1_0/temp4[145] ), .Z(\MC_ARK_ARC_1_0/temp6[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_4  ( .A1(\RI5[0][181] ), .A2(n520), .Z(
        \MC_ARK_ARC_1_0/temp4[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_7_4  ( .A1(\RI5[0][55] ), .A2(\RI5[0][19] ), .Z(
        \MC_ARK_ARC_1_0/temp3[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_7_4  ( .A1(\RI5[0][91] ), .A2(\RI5[0][115] ), .Z(
        \MC_ARK_ARC_1_0/temp2[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_7_4  ( .A1(\RI5[0][145] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[139] ), .Z(\MC_ARK_ARC_1_0/temp1[145] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_3  ( .A1(\RI5[0][182] ), .A2(n135), .Z(
        \MC_ARK_ARC_1_0/temp4[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_7_3  ( .A1(\RI5[0][140] ), .A2(\RI5[0][146] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_2  ( .A1(\RI5[0][183] ), .A2(n202), .Z(
        \MC_ARK_ARC_1_0/temp4[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_7_2  ( .A1(\RI5[0][93] ), .A2(\RI5[0][117] ), .Z(
        \MC_ARK_ARC_1_0/temp2[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_7_1  ( .A1(\MC_ARK_ARC_1_0/temp1[148] ), .A2(
        \MC_ARK_ARC_1_0/temp2[148] ), .Z(\MC_ARK_ARC_1_0/temp5[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_1  ( .A1(\RI5[0][184] ), .A2(n85), .Z(
        \MC_ARK_ARC_1_0/temp4[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_7_1  ( .A1(\RI5[0][58] ), .A2(\RI5[0][22] ), .Z(
        \MC_ARK_ARC_1_0/temp3[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_7_1  ( .A1(\RI5[0][118] ), .A2(\RI5[0][94] ), .Z(
        \MC_ARK_ARC_1_0/temp2[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_7_0  ( .A1(\RI5[0][59] ), .A2(\RI5[0][23] ), .Z(
        \MC_ARK_ARC_1_0/temp3[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_6_5  ( .A1(\MC_ARK_ARC_1_0/temp3[150] ), .A2(
        \MC_ARK_ARC_1_0/temp4[150] ), .Z(\MC_ARK_ARC_1_0/temp6[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_5  ( .A1(\RI5[0][186] ), .A2(n160), .Z(
        \MC_ARK_ARC_1_0/temp4[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_6_5  ( .A1(\RI5[0][60] ), .A2(\RI5[0][24] ), .Z(
        \MC_ARK_ARC_1_0/temp3[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_6_5  ( .A1(\RI5[0][120] ), .A2(\RI5[0][96] ), .Z(
        \MC_ARK_ARC_1_0/temp2[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_6_4  ( .A1(\MC_ARK_ARC_1_0/temp5[151] ), .A2(
        \MC_ARK_ARC_1_0/temp6[151] ), .Z(\MC_ARK_ARC_1_0/buf_output[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_6_4  ( .A1(\MC_ARK_ARC_1_0/temp3[151] ), .A2(
        \MC_ARK_ARC_1_0/temp4[151] ), .Z(\MC_ARK_ARC_1_0/temp6[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_4  ( .A1(\RI5[0][187] ), .A2(n488), .Z(
        \MC_ARK_ARC_1_0/temp4[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_6_4  ( .A1(\RI5[0][61] ), .A2(\RI5[0][25] ), .Z(
        \MC_ARK_ARC_1_0/temp3[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_6_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[97] ), 
        .A2(n7134), .Z(\MC_ARK_ARC_1_0/temp2[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_6_4  ( .A1(\RI5[0][151] ), .A2(\RI5[0][145] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_3  ( .A1(\RI5[0][188] ), .A2(n483), .Z(
        \MC_ARK_ARC_1_0/temp4[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_2  ( .A1(\RI5[0][189] ), .A2(n205), .Z(
        \MC_ARK_ARC_1_0/temp4[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_6_1  ( .A1(\MC_ARK_ARC_1_0/temp5[154] ), .A2(
        \MC_ARK_ARC_1_0/temp6[154] ), .Z(\MC_ARK_ARC_1_0/buf_output[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_6_1  ( .A1(\MC_ARK_ARC_1_0/temp3[154] ), .A2(
        \MC_ARK_ARC_1_0/temp4[154] ), .Z(\MC_ARK_ARC_1_0/temp6[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_6_1  ( .A1(\MC_ARK_ARC_1_0/temp2[154] ), .A2(
        \MC_ARK_ARC_1_0/temp1[154] ), .Z(\MC_ARK_ARC_1_0/temp5[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_1  ( .A1(\RI5[0][190] ), .A2(n469), .Z(
        \MC_ARK_ARC_1_0/temp4[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_6_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .A2(\RI5[0][28] ), .Z(\MC_ARK_ARC_1_0/temp3[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_6_1  ( .A1(\RI5[0][154] ), .A2(\RI5[0][148] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_5  ( .A1(\SB2_0_4/buf_output[0] ), .A2(n131), 
        .Z(\MC_ARK_ARC_1_0/temp4[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_5_5  ( .A1(\RI5[0][66] ), .A2(\RI5[0][30] ), .Z(
        \MC_ARK_ARC_1_0/temp3[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_5_5  ( .A1(\RI5[0][156] ), .A2(\RI5[0][150] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_5_4  ( .A1(\MC_ARK_ARC_1_0/temp5[157] ), .A2(
        \MC_ARK_ARC_1_0/temp6[157] ), .Z(\MC_ARK_ARC_1_0/buf_output[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_5_4  ( .A1(\MC_ARK_ARC_1_0/temp3[157] ), .A2(
        \MC_ARK_ARC_1_0/temp4[157] ), .Z(\MC_ARK_ARC_1_0/temp6[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_5_4  ( .A1(\MC_ARK_ARC_1_0/temp2[157] ), .A2(
        \MC_ARK_ARC_1_0/temp1[157] ), .Z(\MC_ARK_ARC_1_0/temp5[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_4  ( .A1(\RI5[0][1] ), .A2(n53), .Z(
        \MC_ARK_ARC_1_0/temp4[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_5_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[67] ), .Z(
        \MC_ARK_ARC_1_0/temp3[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_5_4  ( .A1(\RI5[0][157] ), .A2(\RI5[0][151] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_3  ( .A1(\RI5[0][2] ), .A2(n5), .Z(
        \MC_ARK_ARC_1_0/temp4[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_5_3  ( .A1(\RI5[0][32] ), .A2(\RI5[0][68] ), .Z(
        \MC_ARK_ARC_1_0/temp3[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_5_3  ( .A1(\RI5[0][104] ), .A2(\RI5[0][128] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_5_3  ( .A1(\RI5[0][158] ), .A2(\RI5[0][152] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_2  ( .A1(\RI5[0][3] ), .A2(n441), .Z(
        \MC_ARK_ARC_1_0/temp4[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_5_2  ( .A1(\RI5[0][33] ), .A2(\RI5[0][69] ), .Z(
        \MC_ARK_ARC_1_0/temp3[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_5_2  ( .A1(\RI5[0][105] ), .A2(\RI5[0][129] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_5_1  ( .A1(\MC_ARK_ARC_1_0/temp3[160] ), .A2(
        \MC_ARK_ARC_1_0/temp4[160] ), .Z(\MC_ARK_ARC_1_0/temp6[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_1  ( .A1(\RI5[0][4] ), .A2(n109), .Z(
        \MC_ARK_ARC_1_0/temp4[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_5_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[70] ), 
        .A2(\RI5[0][34] ), .Z(\MC_ARK_ARC_1_0/temp3[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_5_1  ( .A1(\RI5[0][154] ), .A2(\RI5[0][160] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_5_0  ( .A1(\MC_ARK_ARC_1_0/temp6[161] ), .A2(
        \MC_ARK_ARC_1_0/temp5[161] ), .Z(\MC_ARK_ARC_1_0/buf_output[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_5_0  ( .A1(\MC_ARK_ARC_1_0/temp4[161] ), .A2(
        \MC_ARK_ARC_1_0/temp3[161] ), .Z(\MC_ARK_ARC_1_0/temp6[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_0  ( .A1(\RI5[0][5] ), .A2(n184), .Z(
        \MC_ARK_ARC_1_0/temp4[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_4_5  ( .A1(\MC_ARK_ARC_1_0/temp6[162] ), .A2(
        \MC_ARK_ARC_1_0/temp5[162] ), .Z(\MC_ARK_ARC_1_0/buf_output[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_4_5  ( .A1(\MC_ARK_ARC_1_0/temp1[162] ), .A2(
        \MC_ARK_ARC_1_0/temp2[162] ), .Z(\MC_ARK_ARC_1_0/temp5[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_4_5  ( .A1(\RI5[0][6] ), .A2(n216), .Z(
        \MC_ARK_ARC_1_0/temp4[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_4_5  ( .A1(\RI5[0][72] ), .A2(\RI5[0][36] ), .Z(
        \MC_ARK_ARC_1_0/temp3[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_4_5  ( .A1(\RI5[0][132] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[108] ), .Z(\MC_ARK_ARC_1_0/temp2[162] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_4_5  ( .A1(\RI5[0][162] ), .A2(\RI5[0][156] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_4_4  ( .A1(\MC_ARK_ARC_1_0/temp3[163] ), .A2(
        \MC_ARK_ARC_1_0/temp4[163] ), .Z(\MC_ARK_ARC_1_0/temp6[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_4_4  ( .A1(\RI5[0][7] ), .A2(n418), .Z(
        \MC_ARK_ARC_1_0/temp4[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_4_4  ( .A1(\RI5[0][73] ), .A2(\RI5[0][37] ), .Z(
        \MC_ARK_ARC_1_0/temp3[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_4_4  ( .A1(\SB2_0_13/buf_output[1] ), .A2(
        \RI5[0][109] ), .Z(\MC_ARK_ARC_1_0/temp2[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_4_4  ( .A1(\RI5[0][157] ), .A2(\RI5[0][163] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_4_2  ( .A1(\RI5[0][9] ), .A2(n157), .Z(
        \MC_ARK_ARC_1_0/temp4[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_4_2  ( .A1(\RI5[0][135] ), .A2(\RI5[0][111] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_4_1  ( .A1(\MC_ARK_ARC_1_0/temp1[166] ), .A2(
        \MC_ARK_ARC_1_0/temp2[166] ), .Z(\MC_ARK_ARC_1_0/temp5[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_4_1  ( .A1(\RI5[0][136] ), .A2(\RI5[0][112] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_4_0  ( .A1(\RI5[0][11] ), .A2(n164), .Z(
        \MC_ARK_ARC_1_0/temp4[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_4_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[77] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[41] ), .Z(
        \MC_ARK_ARC_1_0/temp3[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_5  ( .A1(\RI5[0][12] ), .A2(n108), .Z(
        \MC_ARK_ARC_1_0/temp4[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_3_5  ( .A1(\RI5[0][78] ), .A2(\RI5[0][42] ), .Z(
        \MC_ARK_ARC_1_0/temp3[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_3_5  ( .A1(\RI5[0][168] ), .A2(\RI5[0][162] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_3_4  ( .A1(\MC_ARK_ARC_1_0/temp6[169] ), .A2(
        \MC_ARK_ARC_1_0/temp5[169] ), .Z(\MC_ARK_ARC_1_0/buf_output[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_3_4  ( .A1(\MC_ARK_ARC_1_0/temp3[169] ), .A2(
        \MC_ARK_ARC_1_0/temp4[169] ), .Z(\MC_ARK_ARC_1_0/temp6[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_4  ( .A1(\RI5[0][13] ), .A2(n540), .Z(
        \MC_ARK_ARC_1_0/temp4[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_3_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .A2(\RI5[0][79] ), .Z(\MC_ARK_ARC_1_0/temp3[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_3_4  ( .A1(\RI5[0][163] ), .A2(\RI5[0][169] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_3  ( .A1(\RI5[0][14] ), .A2(n214), .Z(
        \MC_ARK_ARC_1_0/temp4[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_3_3  ( .A1(\RI5[0][170] ), .A2(\RI5[0][164] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_3_2  ( .A1(\MC_ARK_ARC_1_0/temp4[171] ), .A2(
        \MC_ARK_ARC_1_0/temp3[171] ), .Z(\MC_ARK_ARC_1_0/temp6[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_2  ( .A1(\RI5[0][15] ), .A2(n529), .Z(
        \MC_ARK_ARC_1_0/temp4[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_1  ( .A1(\RI5[0][16] ), .A2(n72), .Z(
        \MC_ARK_ARC_1_0/temp4[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_3_1  ( .A1(\RI5[0][46] ), .A2(\RI5[0][82] ), .Z(
        \MC_ARK_ARC_1_0/temp3[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_3_1  ( .A1(\RI5[0][172] ), .A2(\RI5[0][166] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_0  ( .A1(\RI5[0][17] ), .A2(n517), .Z(
        \MC_ARK_ARC_1_0/temp4[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_2_5  ( .A1(\MC_ARK_ARC_1_0/temp5[174] ), .A2(
        \MC_ARK_ARC_1_0/temp6[174] ), .Z(\MC_ARK_ARC_1_0/buf_output[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_2_5  ( .A1(\MC_ARK_ARC_1_0/temp3[174] ), .A2(
        \MC_ARK_ARC_1_0/temp4[174] ), .Z(\MC_ARK_ARC_1_0/temp6[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_2_5  ( .A1(\MC_ARK_ARC_1_0/temp2[174] ), .A2(
        \MC_ARK_ARC_1_0/temp1[174] ), .Z(\MC_ARK_ARC_1_0/temp5[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_5  ( .A1(\RI5[0][18] ), .A2(n510), .Z(
        \MC_ARK_ARC_1_0/temp4[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_2_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[84] ), 
        .A2(\RI5[0][48] ), .Z(\MC_ARK_ARC_1_0/temp3[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_2_5  ( .A1(\RI5[0][174] ), .A2(\RI5[0][168] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_2_4  ( .A1(\MC_ARK_ARC_1_0/temp5[175] ), .A2(
        \MC_ARK_ARC_1_0/temp6[175] ), .Z(\MC_ARK_ARC_1_0/buf_output[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_4  ( .A1(\RI5[0][19] ), .A2(n71), .Z(
        \MC_ARK_ARC_1_0/temp4[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_2_4  ( .A1(\RI5[0][145] ), .A2(n7134), .Z(
        \MC_ARK_ARC_1_0/temp2[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_2_4  ( .A1(\RI5[0][175] ), .A2(\RI5[0][169] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_2_2  ( .A1(\MC_ARK_ARC_1_0/temp3[177] ), .A2(
        \MC_ARK_ARC_1_0/temp4[177] ), .Z(\MC_ARK_ARC_1_0/temp6[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_2  ( .A1(\RI5[0][21] ), .A2(n494), .Z(
        \MC_ARK_ARC_1_0/temp4[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_2_2  ( .A1(\RI5[0][177] ), .A2(\RI5[0][171] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_2_1  ( .A1(\MC_ARK_ARC_1_0/temp5[178] ), .A2(
        \MC_ARK_ARC_1_0/temp6[178] ), .Z(\MC_ARK_ARC_1_0/buf_output[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_2_1  ( .A1(\MC_ARK_ARC_1_0/temp4[178] ), .A2(
        \MC_ARK_ARC_1_0/temp3[178] ), .Z(\MC_ARK_ARC_1_0/temp6[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_1  ( .A1(\RI5[0][22] ), .A2(n489), .Z(
        \MC_ARK_ARC_1_0/temp4[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_2_1  ( .A1(\RI5[0][88] ), .A2(\RI5[0][52] ), .Z(
        \MC_ARK_ARC_1_0/temp3[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_2_1  ( .A1(\RI5[0][148] ), .A2(\RI5[0][124] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_2_1  ( .A1(\RI5[0][178] ), .A2(\RI5[0][172] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_0  ( .A1(\RI5[0][23] ), .A2(n84), .Z(
        \MC_ARK_ARC_1_0/temp4[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_1_5  ( .A1(\MC_ARK_ARC_1_0/temp6[180] ), .A2(
        \MC_ARK_ARC_1_0/temp5[180] ), .Z(\MC_ARK_ARC_1_0/buf_output[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_1_5  ( .A1(\MC_ARK_ARC_1_0/temp3[180] ), .A2(
        \MC_ARK_ARC_1_0/temp4[180] ), .Z(\MC_ARK_ARC_1_0/temp6[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_1_5  ( .A1(\MC_ARK_ARC_1_0/temp2[180] ), .A2(
        \MC_ARK_ARC_1_0/temp1[180] ), .Z(\MC_ARK_ARC_1_0/temp5[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_5  ( .A1(\RI5[0][24] ), .A2(n479), .Z(
        \MC_ARK_ARC_1_0/temp4[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_1_5  ( .A1(\RI5[0][90] ), .A2(\RI5[0][54] ), .Z(
        \MC_ARK_ARC_1_0/temp3[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_1_5  ( .A1(\RI5[0][150] ), .A2(\RI5[0][126] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_1_5  ( .A1(\RI5[0][180] ), .A2(\RI5[0][174] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_4  ( .A1(\RI5[0][25] ), .A2(n472), .Z(
        \MC_ARK_ARC_1_0/temp4[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_1_4  ( .A1(\RI5[0][55] ), .A2(\RI5[0][91] ), .Z(
        \MC_ARK_ARC_1_0/temp3[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_1_4  ( .A1(\RI5[0][151] ), .A2(\RI5[0][127] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_1_4  ( .A1(\RI5[0][181] ), .A2(\RI5[0][175] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_1_3  ( .A1(\MC_ARK_ARC_1_0/temp6[182] ), .A2(
        \MC_ARK_ARC_1_0/temp5[182] ), .Z(\MC_ARK_ARC_1_0/buf_output[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_1_3  ( .A1(\MC_ARK_ARC_1_0/temp3[182] ), .A2(
        \MC_ARK_ARC_1_0/temp4[182] ), .Z(\MC_ARK_ARC_1_0/temp6[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_3  ( .A1(\RI5[0][26] ), .A2(n18), .Z(
        \MC_ARK_ARC_1_0/temp4[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_1_3  ( .A1(\RI5[0][92] ), .A2(\RI5[0][56] ), .Z(
        \MC_ARK_ARC_1_0/temp3[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_1_3  ( .A1(\RI5[0][176] ), .A2(\RI5[0][182] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_1_2  ( .A1(\MC_ARK_ARC_1_0/temp3[183] ), .A2(
        \MC_ARK_ARC_1_0/temp4[183] ), .Z(\MC_ARK_ARC_1_0/temp6[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_2  ( .A1(\RI5[0][27] ), .A2(n112), .Z(
        \MC_ARK_ARC_1_0/temp4[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_1_1  ( .A1(\MC_ARK_ARC_1_0/temp3[184] ), .A2(
        \MC_ARK_ARC_1_0/temp4[184] ), .Z(\MC_ARK_ARC_1_0/temp6[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_1_1  ( .A1(\MC_ARK_ARC_1_0/temp2[184] ), .A2(
        \MC_ARK_ARC_1_0/temp1[184] ), .Z(\MC_ARK_ARC_1_0/temp5[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_1  ( .A1(\RI5[0][28] ), .A2(n203), .Z(
        \MC_ARK_ARC_1_0/temp4[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_1_1  ( .A1(\RI5[0][58] ), .A2(\RI5[0][94] ), .Z(
        \MC_ARK_ARC_1_0/temp3[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_1_1  ( .A1(\RI5[0][154] ), .A2(\RI5[0][130] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_1_1  ( .A1(\RI5[0][178] ), .A2(\RI5[0][184] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_1_0  ( .A1(\MC_ARK_ARC_1_0/temp6[185] ), .A2(
        \MC_ARK_ARC_1_0/temp5[185] ), .Z(\MC_ARK_ARC_1_0/buf_output[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_1_0  ( .A1(\MC_ARK_ARC_1_0/temp3[185] ), .A2(
        \MC_ARK_ARC_1_0/temp4[185] ), .Z(\MC_ARK_ARC_1_0/temp6[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_0  ( .A1(\RI5[0][29] ), .A2(n219), .Z(
        \MC_ARK_ARC_1_0/temp4[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_1_0  ( .A1(\RI5[0][59] ), .A2(\RI5[0][95] ), .Z(
        \MC_ARK_ARC_1_0/temp3[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_1_0  ( .A1(\RI5[0][185] ), .A2(\RI5[0][179] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_0_5  ( .A1(\MC_ARK_ARC_1_0/temp3[186] ), .A2(
        \MC_ARK_ARC_1_0/temp4[186] ), .Z(\MC_ARK_ARC_1_0/temp6[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_5  ( .A1(\RI5[0][30] ), .A2(n444), .Z(
        \MC_ARK_ARC_1_0/temp4[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_0_5  ( .A1(\RI5[0][156] ), .A2(\RI5[0][132] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_0_4  ( .A1(\MC_ARK_ARC_1_0/temp5[187] ), .A2(
        \MC_ARK_ARC_1_0/temp6[187] ), .Z(\MC_ARK_ARC_1_0/buf_output[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_0_4  ( .A1(\MC_ARK_ARC_1_0/temp1[187] ), .A2(
        \MC_ARK_ARC_1_0/temp2[187] ), .Z(\MC_ARK_ARC_1_0/temp5[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .A2(n43), .Z(\MC_ARK_ARC_1_0/temp4[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_0_4  ( .A1(\SB2_0_19/buf_output[1] ), .A2(
        \RI5[0][61] ), .Z(\MC_ARK_ARC_1_0/temp3[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_0_4  ( .A1(\RI5[0][157] ), .A2(\RI5[0][133] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_0_4  ( .A1(\RI5[0][181] ), .A2(\RI5[0][187] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_3  ( .A1(\RI5[0][32] ), .A2(n101), .Z(
        \MC_ARK_ARC_1_0/temp4[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_0_2  ( .A1(\MC_ARK_ARC_1_0/temp3[189] ), .A2(
        \MC_ARK_ARC_1_0/temp4[189] ), .Z(\MC_ARK_ARC_1_0/temp6[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_2  ( .A1(\RI5[0][33] ), .A2(n425), .Z(
        \MC_ARK_ARC_1_0/temp4[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_0_1  ( .A1(\MC_ARK_ARC_1_0/temp6[190] ), .A2(
        \MC_ARK_ARC_1_0/temp5[190] ), .Z(\MC_ARK_ARC_1_0/buf_output[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_0_1  ( .A1(\MC_ARK_ARC_1_0/temp4[190] ), .A2(
        \MC_ARK_ARC_1_0/temp3[190] ), .Z(\MC_ARK_ARC_1_0/temp6[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_1  ( .A1(\RI5[0][34] ), .A2(n208), .Z(
        \MC_ARK_ARC_1_0/temp4[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_0_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .A2(\RI5[0][100] ), .Z(\MC_ARK_ARC_1_0/temp3[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_0_1  ( .A1(\RI5[0][160] ), .A2(\RI5[0][136] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[35] ), 
        .A2(n122), .Z(\MC_ARK_ARC_1_0/temp4[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_0_0  ( .A1(\RI5[0][101] ), .A2(\RI5[0][65] ), .Z(
        \MC_ARK_ARC_1_0/temp3[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_0_0  ( .A1(\SB2_0_5/buf_output[5] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[137] ), .Z(\MC_ARK_ARC_1_0/temp2[191] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_31_5  ( .A1(\MC_ARK_ARC_1_1/temp5[0] ), .A2(
        \MC_ARK_ARC_1_1/temp6[0] ), .Z(\MC_ARK_ARC_1_1/buf_output[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_31_5  ( .A1(\MC_ARK_ARC_1_1/temp3[0] ), .A2(
        \MC_ARK_ARC_1_1/temp4[0] ), .Z(\MC_ARK_ARC_1_1/temp6[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[36] ), 
        .A2(n143), .Z(\MC_ARK_ARC_1_1/temp4[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_31_5  ( .A1(\RI5[1][102] ), .A2(\RI5[1][66] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_31_4  ( .A1(\MC_ARK_ARC_1_1/temp3[1] ), .A2(
        \MC_ARK_ARC_1_1/temp4[1] ), .Z(\MC_ARK_ARC_1_1/temp6[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_31_4  ( .A1(\MC_ARK_ARC_1_1/temp1[1] ), .A2(
        \MC_ARK_ARC_1_1/temp2[1] ), .Z(\MC_ARK_ARC_1_1/temp5[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[37] ), 
        .A2(n98), .Z(\MC_ARK_ARC_1_1/temp4[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_31_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[103] ), 
        .A2(\RI5[1][67] ), .Z(\MC_ARK_ARC_1_1/temp3[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_31_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .A2(\RI5[1][139] ), .Z(\MC_ARK_ARC_1_1/temp2[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_31_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[187] ), .Z(\MC_ARK_ARC_1_1/temp1[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_31_3  ( .A1(\MC_ARK_ARC_1_1/temp1[2] ), .A2(
        \MC_ARK_ARC_1_1/temp2[2] ), .Z(\MC_ARK_ARC_1_1/temp5[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[38] ), 
        .A2(n457), .Z(\MC_ARK_ARC_1_1/temp4[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_31_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[164] ), 
        .A2(\RI5[1][140] ), .Z(\MC_ARK_ARC_1_1/temp2[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_31_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .A2(\RI5[1][2] ), .Z(\MC_ARK_ARC_1_1/temp1[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_2  ( .A1(\RI5[1][39] ), .A2(n417), .Z(
        \MC_ARK_ARC_1_1/temp4[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_31_2  ( .A1(\RI5[1][165] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_1/temp2[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_31_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[189] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[3] ), .Z(\MC_ARK_ARC_1_1/temp1[3] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_1  ( .A1(\RI5[1][40] ), .A2(n177), .Z(
        \MC_ARK_ARC_1_1/temp4[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_31_1  ( .A1(\RI5[1][70] ), .A2(\RI5[1][106] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_31_1  ( .A1(\RI5[1][142] ), .A2(\RI5[1][166] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_31_0  ( .A1(\MC_ARK_ARC_1_1/temp1[5] ), .A2(
        \MC_ARK_ARC_1_1/temp2[5] ), .Z(\MC_ARK_ARC_1_1/temp5[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_0  ( .A1(\RI5[1][41] ), .A2(n493), .Z(
        \MC_ARK_ARC_1_1/temp4[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_31_0  ( .A1(\RI5[1][143] ), .A2(\RI5[1][167] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_30_5  ( .A1(\MC_ARK_ARC_1_1/temp2[6] ), .A2(
        \MC_ARK_ARC_1_1/temp1[6] ), .Z(\MC_ARK_ARC_1_1/temp5[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_5  ( .A1(\RI5[1][42] ), .A2(n50), .Z(
        \MC_ARK_ARC_1_1/temp4[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_30_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[108] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[72] ), .Z(\MC_ARK_ARC_1_1/temp3[6] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_30_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[168] ), 
        .A2(\RI5[1][144] ), .Z(\MC_ARK_ARC_1_1/temp2[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_30_5  ( .A1(\RI5[1][6] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[0] ), .Z(\MC_ARK_ARC_1_1/temp1[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_4  ( .A1(\RI5[1][43] ), .A2(n174), .Z(
        \MC_ARK_ARC_1_1/temp4[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[44] ), 
        .A2(n67), .Z(\MC_ARK_ARC_1_1/temp4[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_30_3  ( .A1(\SB2_1_22/buf_output[2] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[110] ), .Z(\MC_ARK_ARC_1_1/temp3[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_30_3  ( .A1(n3168), .A2(\RI5[1][2] ), .Z(
        \MC_ARK_ARC_1_1/temp1[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_30_2  ( .A1(\MC_ARK_ARC_1_1/temp3[9] ), .A2(
        \MC_ARK_ARC_1_1/temp4[9] ), .Z(\MC_ARK_ARC_1_1/temp6[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[45] ), 
        .A2(n168), .Z(\MC_ARK_ARC_1_1/temp4[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_30_2  ( .A1(\RI5[1][75] ), .A2(\RI5[1][111] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_30_2  ( .A1(\RI5[1][147] ), .A2(\RI5[1][171] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_1  ( .A1(\RI5[1][46] ), .A2(n451), .Z(
        \MC_ARK_ARC_1_1/temp4[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_30_1  ( .A1(\RI5[1][112] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_1/temp3[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_30_1  ( .A1(\RI5[1][10] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[4] ), .Z(\MC_ARK_ARC_1_1/temp1[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_30_0  ( .A1(\MC_ARK_ARC_1_1/temp3[11] ), .A2(
        \MC_ARK_ARC_1_1/temp4[11] ), .Z(\MC_ARK_ARC_1_1/temp6[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_0  ( .A1(\RI5[1][47] ), .A2(n566), .Z(
        \MC_ARK_ARC_1_1/temp4[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_30_0  ( .A1(\RI5[1][113] ), .A2(\RI5[1][77] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_30_0  ( .A1(\RI5[1][173] ), .A2(\RI5[1][149] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_30_0  ( .A1(\RI5[1][5] ), .A2(\RI5[1][11] ), .Z(
        \MC_ARK_ARC_1_1/temp1[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_29_5  ( .A1(\MC_ARK_ARC_1_1/temp5[12] ), .A2(
        \MC_ARK_ARC_1_1/temp6[12] ), .Z(\MC_ARK_ARC_1_1/buf_output[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_29_5  ( .A1(\MC_ARK_ARC_1_1/temp2[12] ), .A2(
        \MC_ARK_ARC_1_1/temp1[12] ), .Z(\MC_ARK_ARC_1_1/temp5[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[48] ), 
        .A2(n142), .Z(\MC_ARK_ARC_1_1/temp4[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_29_5  ( .A1(\RI5[1][174] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[150] ), .Z(\MC_ARK_ARC_1_1/temp2[12] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_29_5  ( .A1(\RI5[1][12] ), .A2(\RI5[1][6] ), .Z(
        \MC_ARK_ARC_1_1/temp1[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_29_4  ( .A1(\MC_ARK_ARC_1_1/temp4[13] ), .A2(
        \MC_ARK_ARC_1_1/temp3[13] ), .Z(\MC_ARK_ARC_1_1/temp6[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_4  ( .A1(\RI5[1][49] ), .A2(n212), .Z(
        \MC_ARK_ARC_1_1/temp4[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_29_4  ( .A1(\RI5[1][115] ), .A2(\RI5[1][79] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_2  ( .A1(\SB2_1_25/buf_output[3] ), .A2(n193), 
        .Z(\MC_ARK_ARC_1_1/temp4[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_29_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[177] ), 
        .A2(\RI5[1][153] ), .Z(\MC_ARK_ARC_1_1/temp2[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_29_1  ( .A1(\MC_ARK_ARC_1_1/temp6[16] ), .A2(
        \MC_ARK_ARC_1_1/temp5[16] ), .Z(\MC_ARK_ARC_1_1/buf_output[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_29_1  ( .A1(\MC_ARK_ARC_1_1/temp1[16] ), .A2(
        \MC_ARK_ARC_1_1/temp2[16] ), .Z(\MC_ARK_ARC_1_1/temp5[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_1  ( .A1(\RI5[1][52] ), .A2(n523), .Z(
        \MC_ARK_ARC_1_1/temp4[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_29_1  ( .A1(\RI5[1][118] ), .A2(\RI5[1][82] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_29_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[178] ), 
        .A2(\RI5[1][154] ), .Z(\MC_ARK_ARC_1_1/temp2[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_29_1  ( .A1(\RI5[1][16] ), .A2(\RI5[1][10] ), .Z(
        \MC_ARK_ARC_1_1/temp1[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_0  ( .A1(\RI5[1][53] ), .A2(n120), .Z(
        \MC_ARK_ARC_1_1/temp4[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_29_0  ( .A1(\RI5[1][17] ), .A2(\RI5[1][11] ), .Z(
        \MC_ARK_ARC_1_1/temp1[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_28_5  ( .A1(\MC_ARK_ARC_1_1/temp3[18] ), .A2(
        \MC_ARK_ARC_1_1/temp4[18] ), .Z(\MC_ARK_ARC_1_1/temp6[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_5  ( .A1(\RI5[1][54] ), .A2(n211), .Z(
        \MC_ARK_ARC_1_1/temp4[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_28_5  ( .A1(\RI5[1][120] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[84] ), .Z(\MC_ARK_ARC_1_1/temp3[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_28_5  ( .A1(\RI5[1][180] ), .A2(\RI5[1][156] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_28_4  ( .A1(\MC_ARK_ARC_1_1/temp5[19] ), .A2(
        \MC_ARK_ARC_1_1/temp6[19] ), .Z(\MC_ARK_ARC_1_1/buf_output[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_28_4  ( .A1(\MC_ARK_ARC_1_1/temp3[19] ), .A2(
        \MC_ARK_ARC_1_1/temp4[19] ), .Z(\MC_ARK_ARC_1_1/temp6[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_28_4  ( .A1(\MC_ARK_ARC_1_1/temp1[19] ), .A2(
        \MC_ARK_ARC_1_1/temp2[19] ), .Z(\MC_ARK_ARC_1_1/temp5[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_4  ( .A1(\RI5[1][55] ), .A2(n559), .Z(
        \MC_ARK_ARC_1_1/temp4[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_28_4  ( .A1(\RI5[1][181] ), .A2(\RI5[1][157] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_28_4  ( .A1(\RI5[1][19] ), .A2(\RI5[1][13] ), .Z(
        \MC_ARK_ARC_1_1/temp1[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_28_3  ( .A1(\MC_ARK_ARC_1_1/temp3[20] ), .A2(
        \MC_ARK_ARC_1_1/temp4[20] ), .Z(\MC_ARK_ARC_1_1/temp6[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_3  ( .A1(\RI5[1][56] ), .A2(n79), .Z(
        \MC_ARK_ARC_1_1/temp4[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_28_2  ( .A1(\MC_ARK_ARC_1_1/temp3[21] ), .A2(
        \MC_ARK_ARC_1_1/temp4[21] ), .Z(\MC_ARK_ARC_1_1/temp6[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_2  ( .A1(\RI5[1][57] ), .A2(n483), .Z(
        \MC_ARK_ARC_1_1/temp4[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_28_1  ( .A1(\MC_ARK_ARC_1_1/temp5[22] ), .A2(
        \MC_ARK_ARC_1_1/temp6[22] ), .Z(\MC_ARK_ARC_1_1/buf_output[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_28_1  ( .A1(\MC_ARK_ARC_1_1/temp3[22] ), .A2(
        \MC_ARK_ARC_1_1/temp4[22] ), .Z(\MC_ARK_ARC_1_1/temp6[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_28_1  ( .A1(\MC_ARK_ARC_1_1/temp1[22] ), .A2(
        \MC_ARK_ARC_1_1/temp2[22] ), .Z(\MC_ARK_ARC_1_1/temp5[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .A2(n441), .Z(\MC_ARK_ARC_1_1/temp4[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_28_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[124] ), 
        .A2(\RI5[1][88] ), .Z(\MC_ARK_ARC_1_1/temp3[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_28_1  ( .A1(\RI5[1][184] ), .A2(\RI5[1][160] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_28_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .A2(\RI5[1][16] ), .Z(\MC_ARK_ARC_1_1/temp1[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_0  ( .A1(\RI5[1][59] ), .A2(n171), .Z(
        \MC_ARK_ARC_1_1/temp4[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_27_5  ( .A1(\MC_ARK_ARC_1_1/temp2[24] ), .A2(
        \MC_ARK_ARC_1_1/temp1[24] ), .Z(\MC_ARK_ARC_1_1/temp5[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_5  ( .A1(\RI5[1][60] ), .A2(n40), .Z(
        \MC_ARK_ARC_1_1/temp4[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_27_5  ( .A1(\RI5[1][90] ), .A2(\RI5[1][126] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_27_5  ( .A1(\RI5[1][186] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[162] ), .Z(\MC_ARK_ARC_1_1/temp2[24] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_27_5  ( .A1(\RI5[1][24] ), .A2(\RI5[1][18] ), .Z(
        \MC_ARK_ARC_1_1/temp1[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_27_4  ( .A1(\MC_ARK_ARC_1_1/temp3[25] ), .A2(
        \MC_ARK_ARC_1_1/temp4[25] ), .Z(\MC_ARK_ARC_1_1/temp6[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_4  ( .A1(\RI5[1][61] ), .A2(n176), .Z(
        \MC_ARK_ARC_1_1/temp4[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_27_4  ( .A1(\RI5[1][127] ), .A2(\RI5[1][91] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_27_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[163] ), .Z(
        \MC_ARK_ARC_1_1/temp2[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .A2(n438), .Z(\MC_ARK_ARC_1_1/temp4[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_2  ( .A1(\RI5[1][63] ), .A2(n215), .Z(
        \MC_ARK_ARC_1_1/temp4[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_27_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[21] ), 
        .A2(\RI5[1][27] ), .Z(\MC_ARK_ARC_1_1/temp1[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_27_1  ( .A1(\MC_ARK_ARC_1_1/temp6[28] ), .A2(
        \MC_ARK_ARC_1_1/temp5[28] ), .Z(\MC_ARK_ARC_1_1/buf_output[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_27_1  ( .A1(\MC_ARK_ARC_1_1/temp3[28] ), .A2(
        \MC_ARK_ARC_1_1/temp4[28] ), .Z(\MC_ARK_ARC_1_1/temp6[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_1  ( .A1(\RI5[1][64] ), .A2(n513), .Z(
        \MC_ARK_ARC_1_1/temp4[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_27_1  ( .A1(\RI5[1][130] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[94] ), .Z(\MC_ARK_ARC_1_1/temp3[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_27_1  ( .A1(\RI5[1][28] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_1/temp1[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_0  ( .A1(\RI5[1][65] ), .A2(n475), .Z(
        \MC_ARK_ARC_1_1/temp4[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_26_5  ( .A1(\MC_ARK_ARC_1_1/temp3[30] ), .A2(
        \MC_ARK_ARC_1_1/temp4[30] ), .Z(\MC_ARK_ARC_1_1/temp6[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_26_5  ( .A1(\MC_ARK_ARC_1_1/temp1[30] ), .A2(
        \MC_ARK_ARC_1_1/temp2[30] ), .Z(\MC_ARK_ARC_1_1/temp5[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_5  ( .A1(\RI5[1][66] ), .A2(n34), .Z(
        \MC_ARK_ARC_1_1/temp4[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_26_5  ( .A1(\RI5[1][132] ), .A2(\RI5[1][96] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_26_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[168] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[0] ), .Z(\MC_ARK_ARC_1_1/temp2[30] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_26_5  ( .A1(\RI5[1][30] ), .A2(\RI5[1][24] ), .Z(
        \MC_ARK_ARC_1_1/temp1[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_4  ( .A1(\RI5[1][67] ), .A2(n91), .Z(
        \MC_ARK_ARC_1_1/temp4[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_26_4  ( .A1(\RI5[1][31] ), .A2(\RI5[1][25] ), .Z(
        \MC_ARK_ARC_1_1/temp1[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_2  ( .A1(\SB2_1_22/buf_output[3] ), .A2(n471), 
        .Z(\MC_ARK_ARC_1_1/temp4[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_26_2  ( .A1(\RI5[1][171] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[3] ), .Z(\MC_ARK_ARC_1_1/temp2[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_26_1  ( .A1(\MC_ARK_ARC_1_1/temp5[34] ), .A2(
        \MC_ARK_ARC_1_1/temp6[34] ), .Z(\MC_ARK_ARC_1_1/buf_output[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_26_1  ( .A1(\MC_ARK_ARC_1_1/temp3[34] ), .A2(
        \MC_ARK_ARC_1_1/temp4[34] ), .Z(\MC_ARK_ARC_1_1/temp6[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_26_1  ( .A1(\MC_ARK_ARC_1_1/temp2[34] ), .A2(
        \MC_ARK_ARC_1_1/temp1[34] ), .Z(\MC_ARK_ARC_1_1/temp5[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_1  ( .A1(\RI5[1][70] ), .A2(n430), .Z(
        \MC_ARK_ARC_1_1/temp4[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_26_1  ( .A1(\RI5[1][136] ), .A2(\RI5[1][100] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_26_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[34] ), 
        .A2(\RI5[1][28] ), .Z(\MC_ARK_ARC_1_1/temp1[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_25_5  ( .A1(\MC_ARK_ARC_1_1/temp5[36] ), .A2(
        \MC_ARK_ARC_1_1/temp6[36] ), .Z(\MC_ARK_ARC_1_1/buf_output[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_25_5  ( .A1(\MC_ARK_ARC_1_1/temp3[36] ), .A2(
        \MC_ARK_ARC_1_1/temp4[36] ), .Z(\MC_ARK_ARC_1_1/temp6[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_25_5  ( .A1(\MC_ARK_ARC_1_1/temp1[36] ), .A2(
        \MC_ARK_ARC_1_1/temp2[36] ), .Z(\MC_ARK_ARC_1_1/temp5[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_25_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[72] ), 
        .A2(n200), .Z(\MC_ARK_ARC_1_1/temp4[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_25_5  ( .A1(\RI5[1][138] ), .A2(\RI5[1][102] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_25_5  ( .A1(\RI5[1][6] ), .A2(\RI5[1][174] ), .Z(
        \MC_ARK_ARC_1_1/temp2[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_25_5  ( .A1(\RI5[1][30] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[36] ), .Z(\MC_ARK_ARC_1_1/temp1[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_25_4  ( .A1(\MC_ARK_ARC_1_1/temp3[37] ), .A2(
        \MC_ARK_ARC_1_1/temp4[37] ), .Z(\MC_ARK_ARC_1_1/temp6[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_25_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[73] ), 
        .A2(n170), .Z(\MC_ARK_ARC_1_1/temp4[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_25_4  ( .A1(\RI5[1][139] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[103] ), .Z(\MC_ARK_ARC_1_1/temp3[37] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_25_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[7] ), 
        .A2(\RI5[1][175] ), .Z(\MC_ARK_ARC_1_1/temp2[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_25_3  ( .A1(n3167), .A2(\RI5[1][176] ), .Z(
        \MC_ARK_ARC_1_1/temp2[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_25_2  ( .A1(\MC_ARK_ARC_1_1/temp6[39] ), .A2(
        \MC_ARK_ARC_1_1/temp5[39] ), .Z(\MC_ARK_ARC_1_1/buf_output[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_25_2  ( .A1(\MC_ARK_ARC_1_1/temp4[39] ), .A2(
        \MC_ARK_ARC_1_1/temp3[39] ), .Z(\MC_ARK_ARC_1_1/temp6[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_25_2  ( .A1(\RI5[1][75] ), .A2(n543), .Z(
        \MC_ARK_ARC_1_1/temp4[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_25_2  ( .A1(\RI5[1][105] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_1/temp3[39] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_25_2  ( .A1(\RI5[1][9] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[177] ), .Z(\MC_ARK_ARC_1_1/temp2[39] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_25_1  ( .A1(\MC_ARK_ARC_1_1/temp6[40] ), .A2(
        \MC_ARK_ARC_1_1/temp5[40] ), .Z(\MC_ARK_ARC_1_1/buf_output[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_25_1  ( .A1(\MC_ARK_ARC_1_1/temp3[40] ), .A2(
        \MC_ARK_ARC_1_1/temp4[40] ), .Z(\MC_ARK_ARC_1_1/temp6[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_25_1  ( .A1(\MC_ARK_ARC_1_1/temp1[40] ), .A2(
        \MC_ARK_ARC_1_1/temp2[40] ), .Z(\MC_ARK_ARC_1_1/temp5[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_25_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[76] ), 
        .A2(n207), .Z(\MC_ARK_ARC_1_1/temp4[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_25_1  ( .A1(\RI5[1][142] ), .A2(\RI5[1][106] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_25_1  ( .A1(\RI5[1][10] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[178] ), .Z(\MC_ARK_ARC_1_1/temp2[40] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_25_1  ( .A1(\RI5[1][40] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[34] ), .Z(\MC_ARK_ARC_1_1/temp1[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_25_0  ( .A1(\RI5[1][11] ), .A2(\RI5[1][179] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_24_5  ( .A1(\RI5[1][78] ), .A2(n423), .Z(
        \MC_ARK_ARC_1_1/temp4[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_24_5  ( .A1(\RI5[1][144] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[108] ), .Z(\MC_ARK_ARC_1_1/temp3[42] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_24_5  ( .A1(\RI5[1][42] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[36] ), .Z(\MC_ARK_ARC_1_1/temp1[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_24_4  ( .A1(\SB2_1_22/buf_output[1] ), .A2(n123), 
        .Z(\MC_ARK_ARC_1_1/temp4[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_24_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[145] ), 
        .A2(\RI5[1][109] ), .Z(\MC_ARK_ARC_1_1/temp3[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_24_4  ( .A1(\RI5[1][43] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[37] ), .Z(\MC_ARK_ARC_1_1/temp1[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_24_3  ( .A1(\SB2_1_27/buf_output[2] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[38] ), .Z(\MC_ARK_ARC_1_1/temp1[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_24_2  ( .A1(\RI5[1][81] ), .A2(n461), .Z(
        \MC_ARK_ARC_1_1/temp4[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_24_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[15] ), 
        .A2(\RI5[1][183] ), .Z(\MC_ARK_ARC_1_1/temp2[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_24_1  ( .A1(\MC_ARK_ARC_1_1/temp3[46] ), .A2(
        \MC_ARK_ARC_1_1/temp4[46] ), .Z(\MC_ARK_ARC_1_1/temp6[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_24_1  ( .A1(\MC_ARK_ARC_1_1/temp1[46] ), .A2(
        \MC_ARK_ARC_1_1/temp2[46] ), .Z(\MC_ARK_ARC_1_1/temp5[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_24_1  ( .A1(\RI5[1][82] ), .A2(n420), .Z(
        \MC_ARK_ARC_1_1/temp4[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_24_1  ( .A1(\RI5[1][148] ), .A2(\RI5[1][112] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_24_1  ( .A1(\RI5[1][16] ), .A2(\RI5[1][184] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_24_1  ( .A1(\RI5[1][46] ), .A2(\RI5[1][40] ), .Z(
        \MC_ARK_ARC_1_1/temp1[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_23_5  ( .A1(\MC_ARK_ARC_1_1/temp5[48] ), .A2(
        \MC_ARK_ARC_1_1/temp6[48] ), .Z(\MC_ARK_ARC_1_1/buf_output[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_23_5  ( .A1(\MC_ARK_ARC_1_1/temp3[48] ), .A2(
        \MC_ARK_ARC_1_1/temp4[48] ), .Z(\MC_ARK_ARC_1_1/temp6[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_23_5  ( .A1(\MC_ARK_ARC_1_1/temp2[48] ), .A2(
        \MC_ARK_ARC_1_1/temp1[48] ), .Z(\MC_ARK_ARC_1_1/temp5[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .A2(n218), .Z(\MC_ARK_ARC_1_1/temp4[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_23_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[150] ), 
        .A2(\RI5[1][114] ), .Z(\MC_ARK_ARC_1_1/temp3[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_23_5  ( .A1(\RI5[1][186] ), .A2(\RI5[1][18] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_23_5  ( .A1(\RI5[1][42] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[48] ), .Z(\MC_ARK_ARC_1_1/temp1[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_4  ( .A1(\RI5[1][85] ), .A2(n131), .Z(
        \MC_ARK_ARC_1_1/temp4[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_23_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[151] ), 
        .A2(\RI5[1][115] ), .Z(\MC_ARK_ARC_1_1/temp3[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_23_4  ( .A1(\RI5[1][43] ), .A2(\RI5[1][49] ), .Z(
        \MC_ARK_ARC_1_1/temp1[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_3  ( .A1(\RI5[1][86] ), .A2(n418), .Z(
        \MC_ARK_ARC_1_1/temp4[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_23_3  ( .A1(\RI5[1][116] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[152] ), .Z(\MC_ARK_ARC_1_1/temp3[50] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_2  ( .A1(\RI5[1][87] ), .A2(n214), .Z(
        \MC_ARK_ARC_1_1/temp4[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_23_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[189] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[21] ), .Z(\MC_ARK_ARC_1_1/temp2[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_23_2  ( .A1(\RI5[1][51] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[45] ), .Z(\MC_ARK_ARC_1_1/temp1[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_23_1  ( .A1(\MC_ARK_ARC_1_1/temp5[52] ), .A2(
        \MC_ARK_ARC_1_1/temp6[52] ), .Z(\MC_ARK_ARC_1_1/buf_output[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_23_1  ( .A1(\MC_ARK_ARC_1_1/temp4[52] ), .A2(
        \MC_ARK_ARC_1_1/temp3[52] ), .Z(\MC_ARK_ARC_1_1/temp6[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_23_1  ( .A1(\MC_ARK_ARC_1_1/temp2[52] ), .A2(
        \MC_ARK_ARC_1_1/temp1[52] ), .Z(\MC_ARK_ARC_1_1/temp5[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_1  ( .A1(\RI5[1][88] ), .A2(n494), .Z(
        \MC_ARK_ARC_1_1/temp4[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_23_1  ( .A1(\RI5[1][154] ), .A2(\RI5[1][118] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_23_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .A2(\RI5[1][190] ), .Z(\MC_ARK_ARC_1_1/temp2[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_23_1  ( .A1(\RI5[1][52] ), .A2(\RI5[1][46] ), .Z(
        \MC_ARK_ARC_1_1/temp1[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_23_0  ( .A1(\MC_ARK_ARC_1_1/temp5[53] ), .A2(
        \MC_ARK_ARC_1_1/temp6[53] ), .Z(\MC_ARK_ARC_1_1/buf_output[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_0  ( .A1(\RI5[1][89] ), .A2(n203), .Z(
        \MC_ARK_ARC_1_1/temp4[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_23_0  ( .A1(\RI5[1][119] ), .A2(\RI5[1][155] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_23_0  ( .A1(\RI5[1][191] ), .A2(\RI5[1][23] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_5  ( .A1(\RI5[1][90] ), .A2(n414), .Z(
        \MC_ARK_ARC_1_1/temp4[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_22_5  ( .A1(\RI5[1][54] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[48] ), .Z(\MC_ARK_ARC_1_1/temp1[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_4  ( .A1(\RI5[1][91] ), .A2(n185), .Z(
        \MC_ARK_ARC_1_1/temp4[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_22_4  ( .A1(\RI5[1][157] ), .A2(\RI5[1][121] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_22_4  ( .A1(\RI5[1][55] ), .A2(\RI5[1][49] ), .Z(
        \MC_ARK_ARC_1_1/temp1[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_2  ( .A1(\SB2_1_18/buf_output[3] ), .A2(n452), 
        .Z(\MC_ARK_ARC_1_1/temp4[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_22_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[3] ), 
        .A2(\RI5[1][27] ), .Z(\MC_ARK_ARC_1_1/temp2[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_22_1  ( .A1(\MC_ARK_ARC_1_1/temp3[58] ), .A2(
        \MC_ARK_ARC_1_1/temp4[58] ), .Z(\MC_ARK_ARC_1_1/temp6[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[94] ), 
        .A2(n567), .Z(\MC_ARK_ARC_1_1/temp4[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_22_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[124] ), 
        .A2(\RI5[1][160] ), .Z(\MC_ARK_ARC_1_1/temp3[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_22_1  ( .A1(\RI5[1][28] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[4] ), .Z(\MC_ARK_ARC_1_1/temp2[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_0  ( .A1(\RI5[1][95] ), .A2(n528), .Z(
        \MC_ARK_ARC_1_1/temp4[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_5  ( .A1(\RI5[1][96] ), .A2(n90), .Z(
        \MC_ARK_ARC_1_1/temp4[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_21_4  ( .A1(\MC_ARK_ARC_1_1/temp5[61] ), .A2(
        \MC_ARK_ARC_1_1/temp6[61] ), .Z(\MC_ARK_ARC_1_1/buf_output[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_21_4  ( .A1(\MC_ARK_ARC_1_1/temp3[61] ), .A2(
        \MC_ARK_ARC_1_1/temp4[61] ), .Z(\MC_ARK_ARC_1_1/temp6[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_4  ( .A1(\RI5[1][97] ), .A2(n450), .Z(
        \MC_ARK_ARC_1_1/temp4[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_21_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .A2(\RI5[1][127] ), .Z(\MC_ARK_ARC_1_1/temp3[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_21_4  ( .A1(\RI5[1][31] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[7] ), .Z(\MC_ARK_ARC_1_1/temp2[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_21_4  ( .A1(\RI5[1][61] ), .A2(\RI5[1][55] ), .Z(
        \MC_ARK_ARC_1_1/temp1[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_3  ( .A1(\RI5[1][98] ), .A2(n46), .Z(
        \MC_ARK_ARC_1_1/temp4[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_21_3  ( .A1(\RI5[1][128] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[164] ), .Z(\MC_ARK_ARC_1_1/temp3[62] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_2  ( .A1(\RI5[1][99] ), .A2(n524), .Z(
        \MC_ARK_ARC_1_1/temp4[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_21_2  ( .A1(\RI5[1][9] ), .A2(\RI5[1][33] ), .Z(
        \MC_ARK_ARC_1_1/temp2[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_1  ( .A1(\RI5[1][100] ), .A2(n487), .Z(
        \MC_ARK_ARC_1_1/temp4[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_21_1  ( .A1(\RI5[1][166] ), .A2(\RI5[1][130] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_21_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[34] ), 
        .A2(\RI5[1][10] ), .Z(\MC_ARK_ARC_1_1/temp2[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_21_0  ( .A1(\MC_ARK_ARC_1_1/temp3[65] ), .A2(
        \MC_ARK_ARC_1_1/temp4[65] ), .Z(\MC_ARK_ARC_1_1/temp6[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_0  ( .A1(\RI5[1][101] ), .A2(n446), .Z(
        \MC_ARK_ARC_1_1/temp4[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_21_0  ( .A1(\RI5[1][131] ), .A2(\RI5[1][167] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_20_5  ( .A1(\MC_ARK_ARC_1_1/temp5[66] ), .A2(
        \MC_ARK_ARC_1_1/temp6[66] ), .Z(\MC_ARK_ARC_1_1/buf_output[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_20_5  ( .A1(\MC_ARK_ARC_1_1/temp2[66] ), .A2(
        \MC_ARK_ARC_1_1/temp1[66] ), .Z(\MC_ARK_ARC_1_1/temp5[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_20_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[36] ), 
        .A2(\RI5[1][12] ), .Z(\MC_ARK_ARC_1_1/temp2[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_20_5  ( .A1(\RI5[1][66] ), .A2(\RI5[1][60] ), .Z(
        \MC_ARK_ARC_1_1/temp1[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_20_4  ( .A1(\MC_ARK_ARC_1_1/temp5[67] ), .A2(
        \MC_ARK_ARC_1_1/temp6[67] ), .Z(\MC_ARK_ARC_1_1/buf_output[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_20_4  ( .A1(\MC_ARK_ARC_1_1/temp3[67] ), .A2(
        \MC_ARK_ARC_1_1/temp4[67] ), .Z(\MC_ARK_ARC_1_1/temp6[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[103] ), 
        .A2(n144), .Z(\MC_ARK_ARC_1_1/temp4[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_20_4  ( .A1(\RI5[1][169] ), .A2(\RI5[1][133] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_20_4  ( .A1(\RI5[1][13] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[37] ), .Z(\MC_ARK_ARC_1_1/temp2[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_20_4  ( .A1(\RI5[1][67] ), .A2(\RI5[1][61] ), .Z(
        \MC_ARK_ARC_1_1/temp1[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_20_3  ( .A1(\MC_ARK_ARC_1_1/temp3[68] ), .A2(
        \MC_ARK_ARC_1_1/temp4[68] ), .Z(\MC_ARK_ARC_1_1/temp6[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_3  ( .A1(\RI5[1][104] ), .A2(n484), .Z(
        \MC_ARK_ARC_1_1/temp4[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_20_3  ( .A1(\RI5[1][134] ), .A2(\RI5[1][170] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_20_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[38] ), 
        .A2(\RI5[1][14] ), .Z(\MC_ARK_ARC_1_1/temp2[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_2  ( .A1(\RI5[1][105] ), .A2(n442), .Z(
        \MC_ARK_ARC_1_1/temp4[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_20_2  ( .A1(\RI5[1][135] ), .A2(\RI5[1][171] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_20_1  ( .A1(\MC_ARK_ARC_1_1/temp3[70] ), .A2(
        \MC_ARK_ARC_1_1/temp4[70] ), .Z(\MC_ARK_ARC_1_1/temp6[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_20_1  ( .A1(\MC_ARK_ARC_1_1/temp1[70] ), .A2(
        \MC_ARK_ARC_1_1/temp2[70] ), .Z(\MC_ARK_ARC_1_1/temp5[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_1  ( .A1(\RI5[1][106] ), .A2(n556), .Z(
        \MC_ARK_ARC_1_1/temp4[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_20_1  ( .A1(n578), .A2(\RI5[1][136] ), .Z(
        \MC_ARK_ARC_1_1/temp3[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_20_1  ( .A1(\RI5[1][40] ), .A2(\RI5[1][16] ), .Z(
        \MC_ARK_ARC_1_1/temp2[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_20_1  ( .A1(\RI5[1][64] ), .A2(\RI5[1][70] ), .Z(
        \MC_ARK_ARC_1_1/temp1[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_0  ( .A1(\RI5[1][107] ), .A2(n110), .Z(
        \MC_ARK_ARC_1_1/temp4[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_20_0  ( .A1(\RI5[1][65] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[71] ), .Z(\MC_ARK_ARC_1_1/temp1[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_19_5  ( .A1(\MC_ARK_ARC_1_1/temp3[72] ), .A2(
        \MC_ARK_ARC_1_1/temp4[72] ), .Z(\MC_ARK_ARC_1_1/temp6[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_19_5  ( .A1(\MC_ARK_ARC_1_1/temp2[72] ), .A2(
        \MC_ARK_ARC_1_1/temp1[72] ), .Z(\MC_ARK_ARC_1_1/temp5[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[108] ), 
        .A2(n480), .Z(\MC_ARK_ARC_1_1/temp4[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_19_5  ( .A1(\RI5[1][138] ), .A2(\RI5[1][174] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_19_5  ( .A1(\RI5[1][18] ), .A2(\RI5[1][42] ), .Z(
        \MC_ARK_ARC_1_1/temp2[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_19_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[72] ), 
        .A2(\RI5[1][66] ), .Z(\MC_ARK_ARC_1_1/temp1[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_19_4  ( .A1(\MC_ARK_ARC_1_1/temp2[73] ), .A2(
        \MC_ARK_ARC_1_1/temp1[73] ), .Z(\MC_ARK_ARC_1_1/temp5[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_4  ( .A1(\RI5[1][109] ), .A2(n439), .Z(
        \MC_ARK_ARC_1_1/temp4[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_19_4  ( .A1(\RI5[1][43] ), .A2(\RI5[1][19] ), .Z(
        \MC_ARK_ARC_1_1/temp2[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_19_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[73] ), 
        .A2(\RI5[1][67] ), .Z(\MC_ARK_ARC_1_1/temp1[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .A2(n56), .Z(\MC_ARK_ARC_1_1/temp4[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_2  ( .A1(\RI5[1][111] ), .A2(n135), .Z(
        \MC_ARK_ARC_1_1/temp4[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_19_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[141] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[177] ), .Z(
        \MC_ARK_ARC_1_1/temp3[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_19_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[21] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[45] ), .Z(\MC_ARK_ARC_1_1/temp2[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_19_2  ( .A1(\RI5[1][75] ), .A2(\RI5[1][69] ), .Z(
        \MC_ARK_ARC_1_1/temp1[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_19_1  ( .A1(\MC_ARK_ARC_1_1/temp3[76] ), .A2(
        \MC_ARK_ARC_1_1/temp4[76] ), .Z(\MC_ARK_ARC_1_1/temp6[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_19_1  ( .A1(\MC_ARK_ARC_1_1/temp2[76] ), .A2(
        \MC_ARK_ARC_1_1/temp1[76] ), .Z(\MC_ARK_ARC_1_1/temp5[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_1  ( .A1(\RI5[1][112] ), .A2(n476), .Z(
        \MC_ARK_ARC_1_1/temp4[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_19_1  ( .A1(\RI5[1][142] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[178] ), .Z(\MC_ARK_ARC_1_1/temp3[76] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_19_1  ( .A1(\RI5[1][46] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_1/temp2[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_19_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[76] ), 
        .A2(\RI5[1][70] ), .Z(\MC_ARK_ARC_1_1/temp1[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_0  ( .A1(\RI5[1][113] ), .A2(n109), .Z(
        \MC_ARK_ARC_1_1/temp4[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_19_0  ( .A1(\RI5[1][143] ), .A2(\RI5[1][179] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_19_0  ( .A1(\RI5[1][77] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[71] ), .Z(\MC_ARK_ARC_1_1/temp1[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_18_5  ( .A1(\RI5[1][114] ), .A2(n188), .Z(
        \MC_ARK_ARC_1_1/temp4[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_18_5  ( .A1(\RI5[1][180] ), .A2(\RI5[1][144] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_18_5  ( .A1(\RI5[1][24] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[48] ), .Z(\MC_ARK_ARC_1_1/temp2[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_18_4  ( .A1(\MC_ARK_ARC_1_1/temp5[79] ), .A2(
        \MC_ARK_ARC_1_1/temp6[79] ), .Z(\MC_ARK_ARC_1_1/buf_output[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_18_4  ( .A1(\RI5[1][115] ), .A2(n150), .Z(
        \MC_ARK_ARC_1_1/temp4[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_18_4  ( .A1(\RI5[1][25] ), .A2(\RI5[1][49] ), .Z(
        \MC_ARK_ARC_1_1/temp2[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_18_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[117] ), 
        .A2(n101), .Z(\MC_ARK_ARC_1_1/temp4[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_18_2  ( .A1(\RI5[1][147] ), .A2(\RI5[1][183] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_18_2  ( .A1(\RI5[1][51] ), .A2(\RI5[1][27] ), .Z(
        \MC_ARK_ARC_1_1/temp2[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_18_1  ( .A1(\RI5[1][118] ), .A2(n155), .Z(
        \MC_ARK_ARC_1_1/temp4[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_17_5  ( .A1(\MC_ARK_ARC_1_1/temp2[84] ), .A2(
        \MC_ARK_ARC_1_1/temp1[84] ), .Z(\MC_ARK_ARC_1_1/temp5[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_5  ( .A1(\RI5[1][120] ), .A2(n468), .Z(
        \MC_ARK_ARC_1_1/temp4[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_17_5  ( .A1(\RI5[1][186] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[150] ), .Z(\MC_ARK_ARC_1_1/temp3[84] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_17_5  ( .A1(\RI5[1][30] ), .A2(\RI5[1][54] ), .Z(
        \MC_ARK_ARC_1_1/temp2[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_17_5  ( .A1(\RI5[1][78] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[84] ), .Z(\MC_ARK_ARC_1_1/temp1[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_17_4  ( .A1(\MC_ARK_ARC_1_1/temp6[85] ), .A2(
        \MC_ARK_ARC_1_1/temp5[85] ), .Z(\MC_ARK_ARC_1_1/buf_output[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_17_4  ( .A1(\MC_ARK_ARC_1_1/temp1[85] ), .A2(
        \MC_ARK_ARC_1_1/temp2[85] ), .Z(\MC_ARK_ARC_1_1/temp5[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_4  ( .A1(\RI5[1][121] ), .A2(n165), .Z(
        \MC_ARK_ARC_1_1/temp4[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_17_4  ( .A1(\SB2_1_30/buf_output[1] ), .A2(
        \RI5[1][55] ), .Z(\MC_ARK_ARC_1_1/temp2[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_17_4  ( .A1(\RI5[1][85] ), .A2(\RI5[1][79] ), .Z(
        \MC_ARK_ARC_1_1/temp1[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_17_3  ( .A1(\MC_ARK_ARC_1_1/temp4[86] ), .A2(
        \MC_ARK_ARC_1_1/temp3[86] ), .Z(\MC_ARK_ARC_1_1/temp6[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[122] ), 
        .A2(n544), .Z(\MC_ARK_ARC_1_1/temp4[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_17_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[152] ), .Z(
        \MC_ARK_ARC_1_1/temp3[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_17_3  ( .A1(\RI5[1][86] ), .A2(\RI5[1][80] ), .Z(
        \MC_ARK_ARC_1_1/temp1[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_17_2  ( .A1(\MC_ARK_ARC_1_1/temp5[87] ), .A2(
        \MC_ARK_ARC_1_1/temp6[87] ), .Z(\MC_ARK_ARC_1_1/buf_output[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_2  ( .A1(\RI5[1][123] ), .A2(n504), .Z(
        \MC_ARK_ARC_1_1/temp4[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_17_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[189] ), 
        .A2(\RI5[1][153] ), .Z(\MC_ARK_ARC_1_1/temp3[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[124] ), 
        .A2(n62), .Z(\MC_ARK_ARC_1_1/temp4[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_17_0  ( .A1(\MC_ARK_ARC_1_1/temp5[89] ), .A2(
        \MC_ARK_ARC_1_1/temp6[89] ), .Z(\MC_ARK_ARC_1_1/buf_output[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_17_0  ( .A1(\MC_ARK_ARC_1_1/temp3[89] ), .A2(
        \MC_ARK_ARC_1_1/temp4[89] ), .Z(\MC_ARK_ARC_1_1/temp6[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[125] ), 
        .A2(n180), .Z(\MC_ARK_ARC_1_1/temp4[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_17_0  ( .A1(\RI5[1][191] ), .A2(\RI5[1][155] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_16_5  ( .A1(\MC_ARK_ARC_1_1/temp2[90] ), .A2(
        \MC_ARK_ARC_1_1/temp1[90] ), .Z(\MC_ARK_ARC_1_1/temp5[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_5  ( .A1(\RI5[1][126] ), .A2(n189), .Z(
        \MC_ARK_ARC_1_1/temp4[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_16_5  ( .A1(\RI5[1][90] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[84] ), .Z(\MC_ARK_ARC_1_1/temp1[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_4  ( .A1(\RI5[1][127] ), .A2(n501), .Z(
        \MC_ARK_ARC_1_1/temp4[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_16_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .A2(\RI5[1][157] ), .Z(\MC_ARK_ARC_1_1/temp3[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_16_4  ( .A1(\RI5[1][61] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[37] ), .Z(\MC_ARK_ARC_1_1/temp2[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_16_4  ( .A1(\RI5[1][91] ), .A2(\RI5[1][85] ), .Z(
        \MC_ARK_ARC_1_1/temp1[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_16_3  ( .A1(\MC_ARK_ARC_1_1/temp4[92] ), .A2(
        \MC_ARK_ARC_1_1/temp3[92] ), .Z(\MC_ARK_ARC_1_1/temp6[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_3  ( .A1(\RI5[1][128] ), .A2(n462), .Z(
        \MC_ARK_ARC_1_1/temp4[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_16_3  ( .A1(\RI5[1][86] ), .A2(\RI5[1][92] ), .Z(
        \MC_ARK_ARC_1_1/temp1[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_2  ( .A1(\RI5[1][129] ), .A2(n421), .Z(
        \MC_ARK_ARC_1_1/temp4[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_16_1  ( .A1(\MC_ARK_ARC_1_1/temp3[94] ), .A2(
        \MC_ARK_ARC_1_1/temp4[94] ), .Z(\MC_ARK_ARC_1_1/temp6[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_16_1  ( .A1(\MC_ARK_ARC_1_1/temp2[94] ), .A2(
        \MC_ARK_ARC_1_1/temp1[94] ), .Z(\MC_ARK_ARC_1_1/temp5[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_1  ( .A1(\RI5[1][130] ), .A2(n152), .Z(
        \MC_ARK_ARC_1_1/temp4[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_16_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[4] ), 
        .A2(\RI5[1][160] ), .Z(\MC_ARK_ARC_1_1/temp3[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_16_1  ( .A1(\RI5[1][64] ), .A2(\RI5[1][40] ), .Z(
        \MC_ARK_ARC_1_1/temp2[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_16_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[94] ), 
        .A2(\RI5[1][88] ), .Z(\MC_ARK_ARC_1_1/temp1[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_0  ( .A1(\RI5[1][131] ), .A2(n75), .Z(
        \MC_ARK_ARC_1_1/temp4[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_15_5  ( .A1(\MC_ARK_ARC_1_1/temp2[96] ), .A2(
        \MC_ARK_ARC_1_1/temp1[96] ), .Z(\MC_ARK_ARC_1_1/temp5[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_5  ( .A1(\RI5[1][132] ), .A2(n61), .Z(
        \MC_ARK_ARC_1_1/temp4[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_15_5  ( .A1(\RI5[1][6] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[162] ), .Z(\MC_ARK_ARC_1_1/temp3[96] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_15_5  ( .A1(\RI5[1][90] ), .A2(\RI5[1][96] ), .Z(
        \MC_ARK_ARC_1_1/temp1[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_15_4  ( .A1(\MC_ARK_ARC_1_1/temp5[97] ), .A2(
        \MC_ARK_ARC_1_1/temp6[97] ), .Z(\MC_ARK_ARC_1_1/buf_output[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_15_4  ( .A1(\MC_ARK_ARC_1_1/temp3[97] ), .A2(
        \MC_ARK_ARC_1_1/temp4[97] ), .Z(\MC_ARK_ARC_1_1/temp6[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_4  ( .A1(\RI5[1][133] ), .A2(n419), .Z(
        \MC_ARK_ARC_1_1/temp4[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_15_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[7] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[163] ), .Z(
        \MC_ARK_ARC_1_1/temp3[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_15_4  ( .A1(\RI5[1][97] ), .A2(\RI5[1][91] ), .Z(
        \MC_ARK_ARC_1_1/temp1[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_2  ( .A1(\RI5[1][135] ), .A2(n192), .Z(
        \MC_ARK_ARC_1_1/temp4[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_15_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[45] ), 
        .A2(\RI5[1][69] ), .Z(\MC_ARK_ARC_1_1/temp2[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_15_2  ( .A1(\RI5[1][93] ), .A2(\RI5[1][99] ), .Z(
        \MC_ARK_ARC_1_1/temp1[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_15_1  ( .A1(\MC_ARK_ARC_1_1/temp3[100] ), .A2(
        \MC_ARK_ARC_1_1/temp4[100] ), .Z(\MC_ARK_ARC_1_1/temp6[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_15_1  ( .A1(\MC_ARK_ARC_1_1/temp1[100] ), .A2(
        \MC_ARK_ARC_1_1/temp2[100] ), .Z(\MC_ARK_ARC_1_1/temp5[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_1  ( .A1(\RI5[1][136] ), .A2(n140), .Z(
        \MC_ARK_ARC_1_1/temp4[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_15_1  ( .A1(\RI5[1][10] ), .A2(\RI5[1][166] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_15_1  ( .A1(\RI5[1][46] ), .A2(\RI5[1][70] ), .Z(
        \MC_ARK_ARC_1_1/temp2[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_15_1  ( .A1(\RI5[1][100] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[94] ), .Z(\MC_ARK_ARC_1_1/temp1[100] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_0  ( .A1(\RI5[1][137] ), .A2(n415), .Z(
        \MC_ARK_ARC_1_1/temp4[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_14_5  ( .A1(\MC_ARK_ARC_1_1/temp6[102] ), .A2(
        \MC_ARK_ARC_1_1/temp5[102] ), .Z(\MC_ARK_ARC_1_1/buf_output[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_14_5  ( .A1(\MC_ARK_ARC_1_1/temp1[102] ), .A2(
        \MC_ARK_ARC_1_1/temp2[102] ), .Z(\MC_ARK_ARC_1_1/temp5[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_14_4  ( .A1(\RI5[1][139] ), .A2(n491), .Z(
        \MC_ARK_ARC_1_1/temp4[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_14_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[73] ), 
        .A2(\RI5[1][49] ), .Z(\MC_ARK_ARC_1_1/temp2[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_14_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[103] ), 
        .A2(\RI5[1][97] ), .Z(\MC_ARK_ARC_1_1/temp1[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_14_3  ( .A1(\RI5[1][140] ), .A2(n453), .Z(
        \MC_ARK_ARC_1_1/temp4[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_14_3  ( .A1(\RI5[1][98] ), .A2(\RI5[1][104] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_14_2  ( .A1(\MC_ARK_ARC_1_1/temp6[105] ), .A2(
        \MC_ARK_ARC_1_1/temp5[105] ), .Z(\MC_ARK_ARC_1_1/buf_output[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_14_2  ( .A1(\MC_ARK_ARC_1_1/temp3[105] ), .A2(
        \MC_ARK_ARC_1_1/temp4[105] ), .Z(\MC_ARK_ARC_1_1/temp6[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_14_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[141] ), 
        .A2(n78), .Z(\MC_ARK_ARC_1_1/temp4[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_14_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[15] ), 
        .A2(\RI5[1][171] ), .Z(\MC_ARK_ARC_1_1/temp3[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_14_2  ( .A1(\RI5[1][105] ), .A2(\RI5[1][99] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_14_1  ( .A1(\MC_ARK_ARC_1_1/temp3[106] ), .A2(
        \MC_ARK_ARC_1_1/temp4[106] ), .Z(\MC_ARK_ARC_1_1/temp6[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_14_1  ( .A1(\SB2_1_9/buf_output[4] ), .A2(n36), 
        .Z(\MC_ARK_ARC_1_1/temp4[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_14_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[76] ), 
        .A2(\RI5[1][52] ), .Z(\MC_ARK_ARC_1_1/temp2[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_13_5  ( .A1(\MC_ARK_ARC_1_1/temp6[108] ), .A2(
        \MC_ARK_ARC_1_1/temp5[108] ), .Z(\MC_ARK_ARC_1_1/buf_output[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_13_5  ( .A1(\MC_ARK_ARC_1_1/temp3[108] ), .A2(
        \MC_ARK_ARC_1_1/temp4[108] ), .Z(\MC_ARK_ARC_1_1/temp6[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_13_5  ( .A1(\MC_ARK_ARC_1_1/temp1[108] ), .A2(
        \MC_ARK_ARC_1_1/temp2[108] ), .Z(\MC_ARK_ARC_1_1/temp5[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_5  ( .A1(\RI5[1][144] ), .A2(n219), .Z(
        \MC_ARK_ARC_1_1/temp4[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_13_5  ( .A1(\RI5[1][18] ), .A2(\RI5[1][174] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_13_5  ( .A1(\RI5[1][54] ), .A2(\RI5[1][78] ), .Z(
        \MC_ARK_ARC_1_1/temp2[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_13_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[108] ), 
        .A2(\RI5[1][102] ), .Z(\MC_ARK_ARC_1_1/temp1[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[145] ), 
        .A2(n564), .Z(\MC_ARK_ARC_1_1/temp4[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_13_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[103] ), 
        .A2(\RI5[1][109] ), .Z(\MC_ARK_ARC_1_1/temp1[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_13_3  ( .A1(\MC_ARK_ARC_1_1/temp3[110] ), .A2(
        \MC_ARK_ARC_1_1/temp4[110] ), .Z(\MC_ARK_ARC_1_1/temp6[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[146] ), 
        .A2(n38), .Z(\MC_ARK_ARC_1_1/temp4[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_13_3  ( .A1(\RI5[1][176] ), .A2(\RI5[1][20] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_13_3  ( .A1(\RI5[1][56] ), .A2(\RI5[1][80] ), .Z(
        \MC_ARK_ARC_1_1/temp2[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_13_2  ( .A1(\MC_ARK_ARC_1_1/temp5[111] ), .A2(
        \MC_ARK_ARC_1_1/temp6[111] ), .Z(\MC_ARK_ARC_1_1/buf_output[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_13_2  ( .A1(\MC_ARK_ARC_1_1/temp3[111] ), .A2(
        \MC_ARK_ARC_1_1/temp4[111] ), .Z(\MC_ARK_ARC_1_1/temp6[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_2  ( .A1(\SB2_1_9/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_1/buf_keyinput[111] ), .Z(\MC_ARK_ARC_1_1/temp4[111] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_13_2  ( .A1(\RI5[1][111] ), .A2(\RI5[1][105] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_1  ( .A1(\RI5[1][148] ), .A2(n114), .Z(
        \MC_ARK_ARC_1_1/temp4[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_0  ( .A1(\RI5[1][149] ), .A2(n133), .Z(
        \MC_ARK_ARC_1_1/temp4[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_12_5  ( .A1(\MC_ARK_ARC_1_1/temp5[114] ), .A2(
        \MC_ARK_ARC_1_1/temp6[114] ), .Z(\MC_ARK_ARC_1_1/buf_output[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_12_5  ( .A1(\MC_ARK_ARC_1_1/temp4[114] ), .A2(
        \MC_ARK_ARC_1_1/temp3[114] ), .Z(\MC_ARK_ARC_1_1/temp6[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_12_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[150] ), 
        .A2(n199), .Z(\MC_ARK_ARC_1_1/temp4[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_12_5  ( .A1(\RI5[1][24] ), .A2(\RI5[1][180] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_12_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[151] ), 
        .A2(n485), .Z(\MC_ARK_ARC_1_1/temp4[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_12_4  ( .A1(\RI5[1][115] ), .A2(\RI5[1][109] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_12_2  ( .A1(\RI5[1][153] ), .A2(n557), .Z(
        \MC_ARK_ARC_1_1/temp4[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_12_2  ( .A1(\SB2_1_19/buf_output[3] ), .A2(
        \RI5[1][63] ), .Z(\MC_ARK_ARC_1_1/temp2[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_12_1  ( .A1(\MC_ARK_ARC_1_1/temp3[118] ), .A2(
        \MC_ARK_ARC_1_1/temp4[118] ), .Z(\MC_ARK_ARC_1_1/temp6[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_12_1  ( .A1(\MC_ARK_ARC_1_1/temp2[118] ), .A2(
        \MC_ARK_ARC_1_1/temp1[118] ), .Z(\MC_ARK_ARC_1_1/temp5[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_12_1  ( .A1(\RI5[1][154] ), .A2(n182), .Z(
        \MC_ARK_ARC_1_1/temp4[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_12_1  ( .A1(\RI5[1][28] ), .A2(\RI5[1][184] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_12_1  ( .A1(\RI5[1][88] ), .A2(\RI5[1][64] ), .Z(
        \MC_ARK_ARC_1_1/temp2[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_12_1  ( .A1(\RI5[1][118] ), .A2(\RI5[1][112] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_12_0  ( .A1(\MC_ARK_ARC_1_1/temp5[119] ), .A2(
        \MC_ARK_ARC_1_1/temp6[119] ), .Z(\MC_ARK_ARC_1_1/buf_output[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_12_0  ( .A1(\RI5[1][155] ), .A2(
        \MC_ARK_ARC_1_1/buf_keyinput[119] ), .Z(\MC_ARK_ARC_1_1/temp4[119] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_5  ( .A1(\RI5[1][156] ), .A2(n440), .Z(
        \MC_ARK_ARC_1_1/temp4[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_4  ( .A1(\RI5[1][157] ), .A2(n92), .Z(
        \MC_ARK_ARC_1_1/temp4[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_3  ( .A1(\RI5[1][158] ), .A2(n515), .Z(
        \MC_ARK_ARC_1_1/temp4[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_2  ( .A1(\RI5[1][159] ), .A2(n81), .Z(
        \MC_ARK_ARC_1_1/temp4[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_11_2  ( .A1(\RI5[1][33] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[189] ), .Z(\MC_ARK_ARC_1_1/temp3[123] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_11_1  ( .A1(\MC_ARK_ARC_1_1/temp3[124] ), .A2(
        \MC_ARK_ARC_1_1/temp4[124] ), .Z(\MC_ARK_ARC_1_1/temp6[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_1  ( .A1(\RI5[1][160] ), .A2(n183), .Z(
        \MC_ARK_ARC_1_1/temp4[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_11_1  ( .A1(\RI5[1][118] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[124] ), .Z(\MC_ARK_ARC_1_1/temp1[124] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_11_0  ( .A1(\MC_ARK_ARC_1_1/temp3[125] ), .A2(
        \MC_ARK_ARC_1_1/temp4[125] ), .Z(\MC_ARK_ARC_1_1/temp6[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_0  ( .A1(\RI5[1][161] ), .A2(n104), .Z(
        \MC_ARK_ARC_1_1/temp4[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_11_0  ( .A1(\RI5[1][191] ), .A2(\RI5[1][35] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_10_5  ( .A1(\MC_ARK_ARC_1_1/temp3[126] ), .A2(
        \MC_ARK_ARC_1_1/temp4[126] ), .Z(\MC_ARK_ARC_1_1/temp6[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_10_5  ( .A1(\MC_ARK_ARC_1_1/temp1[126] ), .A2(
        \MC_ARK_ARC_1_1/temp2[126] ), .Z(\MC_ARK_ARC_1_1/temp5[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[162] ), 
        .A2(n511), .Z(\MC_ARK_ARC_1_1/temp4[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_10_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[0] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[36] ), .Z(
        \MC_ARK_ARC_1_1/temp3[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_10_5  ( .A1(\RI5[1][96] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[72] ), .Z(\MC_ARK_ARC_1_1/temp2[126] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_10_5  ( .A1(\RI5[1][120] ), .A2(\RI5[1][126] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .A2(n159), .Z(\MC_ARK_ARC_1_1/temp4[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_10_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[37] ), .Z(
        \MC_ARK_ARC_1_1/temp3[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_10_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[73] ), 
        .A2(\RI5[1][97] ), .Z(\MC_ARK_ARC_1_1/temp2[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_10_4  ( .A1(\RI5[1][127] ), .A2(\RI5[1][121] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[164] ), 
        .A2(n432), .Z(\MC_ARK_ARC_1_1/temp4[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_10_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[38] ), 
        .A2(\RI5[1][2] ), .Z(\MC_ARK_ARC_1_1/temp3[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_10_3  ( .A1(\SB2_1_22/buf_output[2] ), .A2(
        \RI5[1][98] ), .Z(\MC_ARK_ARC_1_1/temp2[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_10_2  ( .A1(\MC_ARK_ARC_1_1/temp4[129] ), .A2(
        \MC_ARK_ARC_1_1/temp3[129] ), .Z(\MC_ARK_ARC_1_1/temp6[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_2  ( .A1(\RI5[1][165] ), .A2(n146), .Z(
        \MC_ARK_ARC_1_1/temp4[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_10_2  ( .A1(\RI5[1][39] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[3] ), .Z(\MC_ARK_ARC_1_1/temp3[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_10_1  ( .A1(\MC_ARK_ARC_1_1/temp1[130] ), .A2(
        \MC_ARK_ARC_1_1/temp2[130] ), .Z(\MC_ARK_ARC_1_1/temp5[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_1  ( .A1(\RI5[1][166] ), .A2(n202), .Z(
        \MC_ARK_ARC_1_1/temp4[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_10_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[4] ), 
        .A2(\RI5[1][40] ), .Z(\MC_ARK_ARC_1_1/temp3[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_10_1  ( .A1(\RI5[1][100] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_1/temp2[130] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_10_1  ( .A1(\RI5[1][130] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[124] ), .Z(\MC_ARK_ARC_1_1/temp1[130] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_0  ( .A1(\RI5[1][167] ), .A2(n469), .Z(
        \MC_ARK_ARC_1_1/temp4[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_10_0  ( .A1(\RI5[1][41] ), .A2(\RI5[1][5] ), .Z(
        \MC_ARK_ARC_1_1/temp3[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_9_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[168] ), 
        .A2(n184), .Z(\MC_ARK_ARC_1_1/temp4[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_9_5  ( .A1(\RI5[1][102] ), .A2(\RI5[1][78] ), .Z(
        \MC_ARK_ARC_1_1/temp2[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_9_5  ( .A1(\RI5[1][132] ), .A2(\RI5[1][126] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_9_4  ( .A1(\MC_ARK_ARC_1_1/temp1[133] ), .A2(
        \MC_ARK_ARC_1_1/temp2[133] ), .Z(\MC_ARK_ARC_1_1/temp5[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_9_4  ( .A1(\RI5[1][169] ), .A2(n108), .Z(
        \MC_ARK_ARC_1_1/temp4[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_9_4  ( .A1(\RI5[1][79] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[103] ), .Z(\MC_ARK_ARC_1_1/temp2[133] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_9_1  ( .A1(\MC_ARK_ARC_1_1/temp1[136] ), .A2(
        \MC_ARK_ARC_1_1/temp2[136] ), .Z(\MC_ARK_ARC_1_1/temp5[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_9_1  ( .A1(n578), .A2(n19), .Z(
        \MC_ARK_ARC_1_1/temp4[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_9_1  ( .A1(\RI5[1][46] ), .A2(\RI5[1][10] ), .Z(
        \MC_ARK_ARC_1_1/temp3[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_9_1  ( .A1(\RI5[1][82] ), .A2(\RI5[1][106] ), .Z(
        \MC_ARK_ARC_1_1/temp2[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_9_1  ( .A1(\RI5[1][136] ), .A2(\RI5[1][130] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_9_0  ( .A1(\RI5[1][173] ), .A2(n201), .Z(
        \MC_ARK_ARC_1_1/temp4[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_8_5  ( .A1(\MC_ARK_ARC_1_1/temp3[138] ), .A2(
        \MC_ARK_ARC_1_1/temp4[138] ), .Z(\MC_ARK_ARC_1_1/temp6[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_5  ( .A1(\RI5[1][174] ), .A2(n502), .Z(
        \MC_ARK_ARC_1_1/temp4[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_8_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[48] ), 
        .A2(\RI5[1][12] ), .Z(\MC_ARK_ARC_1_1/temp3[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_8_5  ( .A1(\RI5[1][138] ), .A2(\RI5[1][132] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_8_4  ( .A1(\MC_ARK_ARC_1_1/temp3[139] ), .A2(
        \MC_ARK_ARC_1_1/temp4[139] ), .Z(\MC_ARK_ARC_1_1/temp6[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_4  ( .A1(\RI5[1][175] ), .A2(n463), .Z(
        \MC_ARK_ARC_1_1/temp4[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_8_4  ( .A1(\RI5[1][85] ), .A2(\RI5[1][109] ), .Z(
        \MC_ARK_ARC_1_1/temp2[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_8_4  ( .A1(\RI5[1][139] ), .A2(\RI5[1][133] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_8_3  ( .A1(\MC_ARK_ARC_1_1/temp3[140] ), .A2(
        \MC_ARK_ARC_1_1/temp4[140] ), .Z(\MC_ARK_ARC_1_1/temp6[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_3  ( .A1(\RI5[1][176] ), .A2(n111), .Z(
        \MC_ARK_ARC_1_1/temp4[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_8_3  ( .A1(\RI5[1][86] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[110] ), .Z(\MC_ARK_ARC_1_1/temp2[140] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[177] ), 
        .A2(n539), .Z(\MC_ARK_ARC_1_1/temp4[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_8_2  ( .A1(\RI5[1][111] ), .A2(\RI5[1][87] ), .Z(
        \MC_ARK_ARC_1_1/temp2[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_8_1  ( .A1(\MC_ARK_ARC_1_1/temp5[142] ), .A2(
        \MC_ARK_ARC_1_1/temp6[142] ), .Z(\MC_ARK_ARC_1_1/buf_output[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_8_1  ( .A1(\MC_ARK_ARC_1_1/temp3[142] ), .A2(
        \MC_ARK_ARC_1_1/temp4[142] ), .Z(\MC_ARK_ARC_1_1/temp6[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_8_1  ( .A1(\MC_ARK_ARC_1_1/temp1[142] ), .A2(
        \MC_ARK_ARC_1_1/temp2[142] ), .Z(\MC_ARK_ARC_1_1/temp5[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[178] ), 
        .A2(n498), .Z(\MC_ARK_ARC_1_1/temp4[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_8_1  ( .A1(\RI5[1][52] ), .A2(\RI5[1][16] ), .Z(
        \MC_ARK_ARC_1_1/temp3[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_8_1  ( .A1(\RI5[1][112] ), .A2(\RI5[1][88] ), .Z(
        \MC_ARK_ARC_1_1/temp2[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_8_1  ( .A1(\RI5[1][136] ), .A2(\RI5[1][142] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_8_0  ( .A1(\MC_ARK_ARC_1_1/temp3[143] ), .A2(
        \MC_ARK_ARC_1_1/temp4[143] ), .Z(\MC_ARK_ARC_1_1/temp6[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_0  ( .A1(\RI5[1][179] ), .A2(n129), .Z(
        \MC_ARK_ARC_1_1/temp4[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_8_0  ( .A1(\RI5[1][17] ), .A2(\RI5[1][53] ), .Z(
        \MC_ARK_ARC_1_1/temp3[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_5  ( .A1(\RI5[1][180] ), .A2(n195), .Z(
        \MC_ARK_ARC_1_1/temp4[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_7_5  ( .A1(\RI5[1][90] ), .A2(\RI5[1][114] ), .Z(
        \MC_ARK_ARC_1_1/temp2[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_7_4  ( .A1(\MC_ARK_ARC_1_1/temp3[145] ), .A2(
        \MC_ARK_ARC_1_1/temp4[145] ), .Z(\MC_ARK_ARC_1_1/temp6[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_4  ( .A1(\RI5[1][181] ), .A2(n537), .Z(
        \MC_ARK_ARC_1_1/temp4[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_7_4  ( .A1(\RI5[1][115] ), .A2(\RI5[1][91] ), .Z(
        \MC_ARK_ARC_1_1/temp2[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_7_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[145] ), 
        .A2(\RI5[1][139] ), .Z(\MC_ARK_ARC_1_1/temp1[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[182] ), 
        .A2(n495), .Z(\MC_ARK_ARC_1_1/temp4[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_7_1  ( .A1(\MC_ARK_ARC_1_1/temp3[148] ), .A2(
        \MC_ARK_ARC_1_1/temp4[148] ), .Z(\MC_ARK_ARC_1_1/temp6[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_1  ( .A1(\RI5[1][184] ), .A2(
        \MC_ARK_ARC_1_1/buf_keyinput[148] ), .Z(\MC_ARK_ARC_1_1/temp4[148] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_7_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[22] ), .Z(
        \MC_ARK_ARC_1_1/temp3[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_7_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[94] ), 
        .A2(\RI5[1][118] ), .Z(\MC_ARK_ARC_1_1/temp2[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_0  ( .A1(\RI5[1][185] ), .A2(n198), .Z(
        \MC_ARK_ARC_1_1/temp4[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_6_5  ( .A1(\MC_ARK_ARC_1_1/temp3[150] ), .A2(
        \MC_ARK_ARC_1_1/temp4[150] ), .Z(\MC_ARK_ARC_1_1/temp6[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_5  ( .A1(\RI5[1][186] ), .A2(n492), .Z(
        \MC_ARK_ARC_1_1/temp4[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_6_5  ( .A1(\RI5[1][24] ), .A2(\RI5[1][60] ), .Z(
        \MC_ARK_ARC_1_1/temp3[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_6_5  ( .A1(\RI5[1][120] ), .A2(\RI5[1][96] ), .Z(
        \MC_ARK_ARC_1_1/temp2[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_6_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[150] ), 
        .A2(\RI5[1][144] ), .Z(\MC_ARK_ARC_1_1/temp1[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_6_4  ( .A1(\MC_ARK_ARC_1_1/temp3[151] ), .A2(
        \MC_ARK_ARC_1_1/temp4[151] ), .Z(\MC_ARK_ARC_1_1/temp6[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_6_4  ( .A1(\MC_ARK_ARC_1_1/temp2[151] ), .A2(
        \MC_ARK_ARC_1_1/temp1[151] ), .Z(\MC_ARK_ARC_1_1/temp5[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .A2(n209), .Z(\MC_ARK_ARC_1_1/temp4[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_6_4  ( .A1(\RI5[1][25] ), .A2(\RI5[1][61] ), .Z(
        \MC_ARK_ARC_1_1/temp3[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_6_4  ( .A1(\RI5[1][97] ), .A2(\RI5[1][121] ), .Z(
        \MC_ARK_ARC_1_1/temp2[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_6_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[151] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[145] ), .Z(
        \MC_ARK_ARC_1_1/temp1[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_6_3  ( .A1(\MC_ARK_ARC_1_1/temp5[152] ), .A2(
        \MC_ARK_ARC_1_1/temp6[152] ), .Z(\MC_ARK_ARC_1_1/buf_output[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .A2(n37), .Z(\MC_ARK_ARC_1_1/temp4[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_6_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[146] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[152] ), .Z(
        \MC_ARK_ARC_1_1/temp1[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_6_2  ( .A1(\MC_ARK_ARC_1_1/temp3[153] ), .A2(
        \MC_ARK_ARC_1_1/temp4[153] ), .Z(\MC_ARK_ARC_1_1/temp6[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[189] ), 
        .A2(n105), .Z(\MC_ARK_ARC_1_1/temp4[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_6_2  ( .A1(\RI5[1][27] ), .A2(\RI5[1][63] ), .Z(
        \MC_ARK_ARC_1_1/temp3[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_6_2  ( .A1(\RI5[1][123] ), .A2(\RI5[1][99] ), .Z(
        \MC_ARK_ARC_1_1/temp2[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_6_2  ( .A1(\RI5[1][147] ), .A2(\RI5[1][153] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_6_1  ( .A1(\MC_ARK_ARC_1_1/temp3[154] ), .A2(
        \MC_ARK_ARC_1_1/temp4[154] ), .Z(\MC_ARK_ARC_1_1/temp6[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_1  ( .A1(\RI5[1][190] ), .A2(n490), .Z(
        \MC_ARK_ARC_1_1/temp4[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_6_1  ( .A1(\RI5[1][64] ), .A2(\RI5[1][28] ), .Z(
        \MC_ARK_ARC_1_1/temp3[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_6_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[124] ), 
        .A2(\RI5[1][100] ), .Z(\MC_ARK_ARC_1_1/temp2[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_6_0  ( .A1(\MC_ARK_ARC_1_1/temp3[155] ), .A2(
        \MC_ARK_ARC_1_1/temp4[155] ), .Z(\MC_ARK_ARC_1_1/temp6[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_0  ( .A1(\RI5[1][191] ), .A2(n45), .Z(
        \MC_ARK_ARC_1_1/temp4[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_6_0  ( .A1(\RI5[1][155] ), .A2(\RI5[1][149] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[0] ), 
        .A2(n173), .Z(\MC_ARK_ARC_1_1/temp4[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_5_5  ( .A1(\RI5[1][30] ), .A2(\RI5[1][66] ), .Z(
        \MC_ARK_ARC_1_1/temp3[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_5_5  ( .A1(\RI5[1][102] ), .A2(\RI5[1][126] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_5_4  ( .A1(\MC_ARK_ARC_1_1/temp3[157] ), .A2(
        \MC_ARK_ARC_1_1/temp4[157] ), .Z(\MC_ARK_ARC_1_1/temp6[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .A2(n526), .Z(\MC_ARK_ARC_1_1/temp4[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_5_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[151] ), 
        .A2(\RI5[1][157] ), .Z(\MC_ARK_ARC_1_1/temp1[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_3  ( .A1(\RI5[1][2] ), .A2(n488), .Z(
        \MC_ARK_ARC_1_1/temp4[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[3] ), 
        .A2(n448), .Z(\MC_ARK_ARC_1_1/temp4[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_5_2  ( .A1(\RI5[1][159] ), .A2(\RI5[1][153] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_5_1  ( .A1(\MC_ARK_ARC_1_1/temp4[160] ), .A2(
        \MC_ARK_ARC_1_1/temp3[160] ), .Z(\MC_ARK_ARC_1_1/temp6[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[4] ), 
        .A2(n157), .Z(\MC_ARK_ARC_1_1/temp4[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_5_1  ( .A1(\RI5[1][130] ), .A2(\RI5[1][106] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_5_1  ( .A1(\RI5[1][154] ), .A2(\RI5[1][160] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_0  ( .A1(\RI5[1][5] ), .A2(n72), .Z(
        \MC_ARK_ARC_1_1/temp4[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_5_0  ( .A1(\RI5[1][131] ), .A2(\RI5[1][107] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_4_5  ( .A1(\MC_ARK_ARC_1_1/temp6[162] ), .A2(
        \MC_ARK_ARC_1_1/temp5[162] ), .Z(\MC_ARK_ARC_1_1/buf_output[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_4_5  ( .A1(\MC_ARK_ARC_1_1/temp1[162] ), .A2(
        \MC_ARK_ARC_1_1/temp2[162] ), .Z(\MC_ARK_ARC_1_1/temp5[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_4_5  ( .A1(\RI5[1][6] ), .A2(n191), .Z(
        \MC_ARK_ARC_1_1/temp4[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_4_5  ( .A1(\RI5[1][132] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[108] ), .Z(\MC_ARK_ARC_1_1/temp2[162] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_4_5  ( .A1(\RI5[1][156] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[162] ), .Z(\MC_ARK_ARC_1_1/temp1[162] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_4_4  ( .A1(\MC_ARK_ARC_1_1/temp3[163] ), .A2(
        \MC_ARK_ARC_1_1/temp4[163] ), .Z(\MC_ARK_ARC_1_1/temp6[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_4_4  ( .A1(\MC_ARK_ARC_1_1/temp2[163] ), .A2(
        \MC_ARK_ARC_1_1/temp1[163] ), .Z(\MC_ARK_ARC_1_1/temp5[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_4_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[7] ), 
        .A2(n444), .Z(\MC_ARK_ARC_1_1/temp4[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_4_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[73] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[37] ), .Z(
        \MC_ARK_ARC_1_1/temp3[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_4_4  ( .A1(\RI5[1][133] ), .A2(\RI5[1][109] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_4_4  ( .A1(\RI5[1][157] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[163] ), .Z(\MC_ARK_ARC_1_1/temp1[163] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_4_3  ( .A1(n3167), .A2(n558), .Z(
        \MC_ARK_ARC_1_1/temp4[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_4_3  ( .A1(\SB2_1_22/buf_output[2] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[38] ), .Z(\MC_ARK_ARC_1_1/temp3[164] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_4_2  ( .A1(\RI5[1][111] ), .A2(\RI5[1][135] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_4_1  ( .A1(\RI5[1][10] ), .A2(n149), .Z(
        \MC_ARK_ARC_1_1/temp4[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_4_1  ( .A1(\RI5[1][40] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_1/temp3[166] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_4_1  ( .A1(\RI5[1][136] ), .A2(\RI5[1][112] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_5  ( .A1(\RI5[1][12] ), .A2(n126), .Z(
        \MC_ARK_ARC_1_1/temp4[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_3_5  ( .A1(\RI5[1][42] ), .A2(\RI5[1][78] ), .Z(
        \MC_ARK_ARC_1_1/temp3[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_3_5  ( .A1(\RI5[1][138] ), .A2(\RI5[1][114] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_3_4  ( .A1(\MC_ARK_ARC_1_1/temp6[169] ), .A2(
        \MC_ARK_ARC_1_1/temp5[169] ), .Z(\MC_ARK_ARC_1_1/buf_output[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_3_4  ( .A1(\MC_ARK_ARC_1_1/temp3[169] ), .A2(
        \MC_ARK_ARC_1_1/temp4[169] ), .Z(\MC_ARK_ARC_1_1/temp6[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_3_4  ( .A1(\MC_ARK_ARC_1_1/temp2[169] ), .A2(
        \MC_ARK_ARC_1_1/temp1[169] ), .Z(\MC_ARK_ARC_1_1/temp5[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_4  ( .A1(\RI5[1][13] ), .A2(n516), .Z(
        \MC_ARK_ARC_1_1/temp4[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_3_4  ( .A1(\RI5[1][43] ), .A2(\RI5[1][79] ), .Z(
        \MC_ARK_ARC_1_1/temp3[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_3_4  ( .A1(\RI5[1][115] ), .A2(\RI5[1][139] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_3_4  ( .A1(\RI5[1][169] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[163] ), .Z(\MC_ARK_ARC_1_1/temp1[169] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_3  ( .A1(\RI5[1][14] ), .A2(n83), .Z(
        \MC_ARK_ARC_1_1/temp4[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_3_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[44] ), 
        .A2(\RI5[1][80] ), .Z(\MC_ARK_ARC_1_1/temp3[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_2  ( .A1(\SB2_1_31/buf_output[3] ), .A2(n437), 
        .Z(\MC_ARK_ARC_1_1/temp4[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_1  ( .A1(\RI5[1][16] ), .A2(n552), .Z(
        \MC_ARK_ARC_1_1/temp4[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_0  ( .A1(\SB2_1_29/buf_output[5] ), .A2(n512), 
        .Z(\MC_ARK_ARC_1_1/temp4[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_2_5  ( .A1(\MC_ARK_ARC_1_1/temp5[174] ), .A2(
        \MC_ARK_ARC_1_1/temp6[174] ), .Z(\MC_ARK_ARC_1_1/buf_output[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_2_5  ( .A1(\MC_ARK_ARC_1_1/temp3[174] ), .A2(
        \MC_ARK_ARC_1_1/temp4[174] ), .Z(\MC_ARK_ARC_1_1/temp6[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_5  ( .A1(\RI5[1][18] ), .A2(n474), .Z(
        \MC_ARK_ARC_1_1/temp4[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_2_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[48] ), .Z(
        \MC_ARK_ARC_1_1/temp3[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_2_5  ( .A1(\RI5[1][120] ), .A2(\RI5[1][144] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_2_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[168] ), 
        .A2(\RI5[1][174] ), .Z(\MC_ARK_ARC_1_1/temp1[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_4  ( .A1(\RI5[1][19] ), .A2(n433), .Z(
        \MC_ARK_ARC_1_1/temp4[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_2_4  ( .A1(\RI5[1][85] ), .A2(\RI5[1][49] ), .Z(
        \MC_ARK_ARC_1_1/temp3[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_3  ( .A1(\RI5[1][20] ), .A2(n186), .Z(
        \MC_ARK_ARC_1_1/temp4[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_2_2  ( .A1(\MC_ARK_ARC_1_1/temp6[177] ), .A2(
        \MC_ARK_ARC_1_1/temp5[177] ), .Z(\MC_ARK_ARC_1_1/buf_output[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_2_2  ( .A1(\MC_ARK_ARC_1_1/temp3[177] ), .A2(
        \MC_ARK_ARC_1_1/temp4[177] ), .Z(\MC_ARK_ARC_1_1/temp6[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[21] ), 
        .A2(n508), .Z(\MC_ARK_ARC_1_1/temp4[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_2_2  ( .A1(\RI5[1][87] ), .A2(\RI5[1][51] ), .Z(
        \MC_ARK_ARC_1_1/temp3[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_2_2  ( .A1(\RI5[1][147] ), .A2(\RI5[1][123] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_2_1  ( .A1(\MC_ARK_ARC_1_1/temp5[178] ), .A2(
        \MC_ARK_ARC_1_1/temp6[178] ), .Z(\MC_ARK_ARC_1_1/buf_output[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_2_1  ( .A1(\MC_ARK_ARC_1_1/temp3[178] ), .A2(
        \MC_ARK_ARC_1_1/temp4[178] ), .Z(\MC_ARK_ARC_1_1/temp6[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .A2(n470), .Z(\MC_ARK_ARC_1_1/temp4[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_2_1  ( .A1(\RI5[1][88] ), .A2(\RI5[1][52] ), .Z(
        \MC_ARK_ARC_1_1/temp3[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_2_1  ( .A1(\RI5[1][148] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[124] ), .Z(\MC_ARK_ARC_1_1/temp2[178] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_0  ( .A1(\RI5[1][23] ), .A2(n429), .Z(
        \MC_ARK_ARC_1_1/temp4[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_2_0  ( .A1(\RI5[1][173] ), .A2(\RI5[1][179] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_1_5  ( .A1(\MC_ARK_ARC_1_1/temp4[180] ), .A2(
        \MC_ARK_ARC_1_1/temp3[180] ), .Z(\MC_ARK_ARC_1_1/temp6[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_5  ( .A1(\RI5[1][24] ), .A2(n220), .Z(
        \MC_ARK_ARC_1_1/temp4[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_1_5  ( .A1(\RI5[1][90] ), .A2(\RI5[1][54] ), .Z(
        \MC_ARK_ARC_1_1/temp3[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_1_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[150] ), 
        .A2(\RI5[1][126] ), .Z(\MC_ARK_ARC_1_1/temp2[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_1_4  ( .A1(\MC_ARK_ARC_1_1/temp2[181] ), .A2(
        \MC_ARK_ARC_1_1/temp1[181] ), .Z(\MC_ARK_ARC_1_1/temp5[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_4  ( .A1(\RI5[1][25] ), .A2(n506), .Z(
        \MC_ARK_ARC_1_1/temp4[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_1_4  ( .A1(\RI5[1][55] ), .A2(\RI5[1][91] ), .Z(
        \MC_ARK_ARC_1_1/temp3[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_1_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[151] ), 
        .A2(\RI5[1][127] ), .Z(\MC_ARK_ARC_1_1/temp2[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_1_4  ( .A1(\RI5[1][175] ), .A2(\RI5[1][181] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_3  ( .A1(\RI5[1][26] ), .A2(n139), .Z(
        \MC_ARK_ARC_1_1/temp4[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_2  ( .A1(\RI5[1][27] ), .A2(n57), .Z(
        \MC_ARK_ARC_1_1/temp4[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_1_2  ( .A1(\RI5[1][57] ), .A2(\RI5[1][93] ), .Z(
        \MC_ARK_ARC_1_1/temp3[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_1_1  ( .A1(\MC_ARK_ARC_1_1/temp2[184] ), .A2(
        \MC_ARK_ARC_1_1/temp1[184] ), .Z(\MC_ARK_ARC_1_1/temp5[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_1  ( .A1(\RI5[1][28] ), .A2(n130), .Z(
        \MC_ARK_ARC_1_1/temp4[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_1_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[94] ), .Z(
        \MC_ARK_ARC_1_1/temp3[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_1_1  ( .A1(\RI5[1][154] ), .A2(\RI5[1][130] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_1_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[178] ), 
        .A2(\RI5[1][184] ), .Z(\MC_ARK_ARC_1_1/temp1[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_1_0  ( .A1(\MC_ARK_ARC_1_1/temp3[185] ), .A2(
        \MC_ARK_ARC_1_1/temp4[185] ), .Z(\MC_ARK_ARC_1_1/temp6[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_0  ( .A1(\RI5[1][29] ), .A2(n85), .Z(
        \MC_ARK_ARC_1_1/temp4[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_1_0  ( .A1(\RI5[1][131] ), .A2(\RI5[1][155] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_5  ( .A1(\RI5[1][30] ), .A2(n134), .Z(
        \MC_ARK_ARC_1_1/temp4[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_0_5  ( .A1(\RI5[1][96] ), .A2(\RI5[1][60] ), .Z(
        \MC_ARK_ARC_1_1/temp3[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_0_5  ( .A1(\RI5[1][156] ), .A2(\RI5[1][132] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_0_5  ( .A1(\RI5[1][186] ), .A2(\RI5[1][180] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_4  ( .A1(\RI5[1][31] ), .A2(n13), .Z(
        \MC_ARK_ARC_1_1/temp4[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_0_4  ( .A1(\RI5[1][157] ), .A2(\RI5[1][133] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[32] ), 
        .A2(n7), .Z(\MC_ARK_ARC_1_1/temp4[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_0_2  ( .A1(\MC_ARK_ARC_1_1/temp2[189] ), .A2(
        \MC_ARK_ARC_1_1/temp1[189] ), .Z(\MC_ARK_ARC_1_1/temp5[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_2  ( .A1(\RI5[1][33] ), .A2(n116), .Z(
        \MC_ARK_ARC_1_1/temp4[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_0_2  ( .A1(\RI5[1][99] ), .A2(\RI5[1][63] ), .Z(
        \MC_ARK_ARC_1_1/temp3[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_0_2  ( .A1(\RI5[1][135] ), .A2(\RI5[1][159] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_0_1  ( .A1(\MC_ARK_ARC_1_1/temp1[190] ), .A2(
        \MC_ARK_ARC_1_1/temp2[190] ), .Z(\MC_ARK_ARC_1_1/temp5[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[34] ), 
        .A2(n112), .Z(\MC_ARK_ARC_1_1/temp4[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_0_1  ( .A1(\RI5[1][190] ), .A2(\RI5[1][184] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_0  ( .A1(\RI5[1][35] ), .A2(n208), .Z(
        \MC_ARK_ARC_1_1/temp4[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_5  ( .A1(\RI5[2][36] ), .A2(n493), .Z(
        \MC_ARK_ARC_1_2/temp4[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_31_5  ( .A1(\RI5[2][102] ), .A2(\RI5[2][66] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_31_5  ( .A1(\RI5[2][0] ), .A2(\RI5[2][186] ), .Z(
        \MC_ARK_ARC_1_2/temp1[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_4  ( .A1(\RI5[2][37] ), .A2(n527), .Z(
        \MC_ARK_ARC_1_2/temp4[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_31_4  ( .A1(\RI5[2][163] ), .A2(\RI5[2][139] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_3  ( .A1(\RI5[2][38] ), .A2(n163), .Z(
        \MC_ARK_ARC_1_2/temp4[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_2  ( .A1(\RI5[2][39] ), .A2(n438), .Z(
        \MC_ARK_ARC_1_2/temp4[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_31_1  ( .A1(\MC_ARK_ARC_1_2/temp6[4] ), .A2(
        \MC_ARK_ARC_1_2/temp5[4] ), .Z(\MC_ARK_ARC_1_2/buf_output[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_31_1  ( .A1(\MC_ARK_ARC_1_2/temp4[4] ), .A2(
        \MC_ARK_ARC_1_2/temp3[4] ), .Z(\MC_ARK_ARC_1_2/temp6[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_31_1  ( .A1(\MC_ARK_ARC_1_2/temp1[4] ), .A2(
        \MC_ARK_ARC_1_2/temp2[4] ), .Z(\MC_ARK_ARC_1_2/temp5[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[40] ), 
        .A2(n471), .Z(\MC_ARK_ARC_1_2/temp4[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_31_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[70] ), .Z(\MC_ARK_ARC_1_2/temp3[4] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_31_1  ( .A1(\RI5[2][166] ), .A2(\RI5[2][142] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_31_1  ( .A1(\RI5[2][4] ), .A2(\RI5[2][190] ), .Z(
        \MC_ARK_ARC_1_2/temp1[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_31_0  ( .A1(\MC_ARK_ARC_1_2/temp3[5] ), .A2(
        \MC_ARK_ARC_1_2/temp4[5] ), .Z(\MC_ARK_ARC_1_2/temp6[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_0  ( .A1(\SB2_2_25/buf_output[5] ), .A2(n207), 
        .Z(\MC_ARK_ARC_1_2/temp4[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_30_5  ( .A1(\MC_ARK_ARC_1_2/temp1[6] ), .A2(
        \MC_ARK_ARC_1_2/temp2[6] ), .Z(\MC_ARK_ARC_1_2/temp5[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_5  ( .A1(\RI5[2][42] ), .A2(n210), .Z(
        \MC_ARK_ARC_1_2/temp4[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_30_5  ( .A1(\RI5[2][108] ), .A2(\RI5[2][72] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_30_5  ( .A1(\RI5[2][168] ), .A2(\RI5[2][144] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_30_5  ( .A1(\RI5[2][6] ), .A2(\RI5[2][0] ), .Z(
        \MC_ARK_ARC_1_2/temp1[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_4  ( .A1(\RI5[2][43] ), .A2(n122), .Z(
        \MC_ARK_ARC_1_2/temp4[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_30_4  ( .A1(\RI5[2][73] ), .A2(\RI5[2][109] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_30_4  ( .A1(\RI5[2][145] ), .A2(\RI5[2][169] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_3  ( .A1(\RI5[2][44] ), .A2(n450), .Z(
        \MC_ARK_ARC_1_2/temp4[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .A2(n484), .Z(\MC_ARK_ARC_1_2/temp4[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_1  ( .A1(\RI5[2][46] ), .A2(n135), .Z(
        \MC_ARK_ARC_1_2/temp4[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_30_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[172] ), 
        .A2(\RI5[2][148] ), .Z(\MC_ARK_ARC_1_2/temp2[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_0  ( .A1(\RI5[2][47] ), .A2(n547), .Z(
        \MC_ARK_ARC_1_2/temp4[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_30_0  ( .A1(\RI5[2][149] ), .A2(\RI5[2][173] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_29_5  ( .A1(\MC_ARK_ARC_1_2/temp1[12] ), .A2(
        \MC_ARK_ARC_1_2/temp2[12] ), .Z(\MC_ARK_ARC_1_2/temp5[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_5  ( .A1(\RI5[2][48] ), .A2(n424), .Z(
        \MC_ARK_ARC_1_2/temp4[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_29_5  ( .A1(\RI5[2][114] ), .A2(\RI5[2][78] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_29_5  ( .A1(\RI5[2][174] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[150] ), .Z(\MC_ARK_ARC_1_2/temp2[12] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_29_4  ( .A1(\MC_ARK_ARC_1_2/temp3[13] ), .A2(
        \MC_ARK_ARC_1_2/temp4[13] ), .Z(\MC_ARK_ARC_1_2/temp6[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .A2(n458), .Z(\MC_ARK_ARC_1_2/temp4[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_29_4  ( .A1(\RI5[2][175] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[151] ), .Z(\MC_ARK_ARC_1_2/temp2[13] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_3  ( .A1(\RI5[2][50] ), .A2(n491), .Z(
        \MC_ARK_ARC_1_2/temp4[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_2  ( .A1(\RI5[2][51] ), .A2(n525), .Z(
        \MC_ARK_ARC_1_2/temp4[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_29_2  ( .A1(\RI5[2][9] ), .A2(\RI5[2][15] ), .Z(
        \MC_ARK_ARC_1_2/temp1[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_29_1  ( .A1(\MC_ARK_ARC_1_2/temp1[16] ), .A2(
        \MC_ARK_ARC_1_2/temp2[16] ), .Z(\MC_ARK_ARC_1_2/temp5[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .A2(n557), .Z(\MC_ARK_ARC_1_2/temp4[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_29_1  ( .A1(\RI5[2][118] ), .A2(\RI5[2][82] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_29_1  ( .A1(\RI5[2][178] ), .A2(\RI5[2][154] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_29_1  ( .A1(\RI5[2][16] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[10] ), .Z(\MC_ARK_ARC_1_2/temp1[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_29_0  ( .A1(\RI5[2][17] ), .A2(\RI5[2][11] ), .Z(
        \MC_ARK_ARC_1_2/temp1[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_28_5  ( .A1(\MC_ARK_ARC_1_2/temp4[18] ), .A2(
        \MC_ARK_ARC_1_2/temp3[18] ), .Z(\MC_ARK_ARC_1_2/temp6[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_28_5  ( .A1(\RI5[2][54] ), .A2(n161), .Z(
        \MC_ARK_ARC_1_2/temp4[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_28_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[84] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[120] ), .Z(
        \MC_ARK_ARC_1_2/temp3[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_28_5  ( .A1(\RI5[2][18] ), .A2(\RI5[2][12] ), .Z(
        \MC_ARK_ARC_1_2/temp1[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_28_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[55] ), 
        .A2(n502), .Z(\MC_ARK_ARC_1_2/temp4[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_28_3  ( .A1(\RI5[2][158] ), .A2(\RI5[2][182] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_28_2  ( .A1(\RI5[2][57] ), .A2(n569), .Z(
        \MC_ARK_ARC_1_2/temp4[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_28_2  ( .A1(\RI5[2][159] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[183] ), .Z(\MC_ARK_ARC_1_2/temp2[21] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_28_2  ( .A1(\RI5[2][15] ), .A2(\RI5[2][21] ), .Z(
        \MC_ARK_ARC_1_2/temp1[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_28_1  ( .A1(\RI5[2][58] ), .A2(n448), .Z(
        \MC_ARK_ARC_1_2/temp4[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_28_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[22] ), 
        .A2(\RI5[2][16] ), .Z(\MC_ARK_ARC_1_2/temp1[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_28_0  ( .A1(\RI5[2][185] ), .A2(\RI5[2][161] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[60] ), 
        .A2(n512), .Z(\MC_ARK_ARC_1_2/temp4[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_27_5  ( .A1(\RI5[2][90] ), .A2(\RI5[2][126] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_27_5  ( .A1(\RI5[2][186] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[162] ), .Z(\MC_ARK_ARC_1_2/temp2[24] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_27_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[24] ), 
        .A2(\RI5[2][18] ), .Z(\MC_ARK_ARC_1_2/temp1[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_27_4  ( .A1(\MC_ARK_ARC_1_2/temp5[25] ), .A2(
        \MC_ARK_ARC_1_2/temp6[25] ), .Z(\MC_ARK_ARC_1_2/buf_output[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_27_4  ( .A1(\MC_ARK_ARC_1_2/temp1[25] ), .A2(
        \MC_ARK_ARC_1_2/temp2[25] ), .Z(\MC_ARK_ARC_1_2/temp5[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .A2(n220), .Z(\MC_ARK_ARC_1_2/temp4[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_27_4  ( .A1(\RI5[2][187] ), .A2(\RI5[2][163] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_27_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[25] ), 
        .A2(\RI5[2][19] ), .Z(\MC_ARK_ARC_1_2/temp1[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_3  ( .A1(\RI5[2][62] ), .A2(n216), .Z(
        \MC_ARK_ARC_1_2/temp4[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_27_3  ( .A1(\RI5[2][128] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[92] ), .Z(\MC_ARK_ARC_1_2/temp3[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_27_2  ( .A1(\MC_ARK_ARC_1_2/temp3[27] ), .A2(
        \MC_ARK_ARC_1_2/temp4[27] ), .Z(\MC_ARK_ARC_1_2/temp6[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_27_2  ( .A1(\MC_ARK_ARC_1_2/temp2[27] ), .A2(
        \MC_ARK_ARC_1_2/temp1[27] ), .Z(\MC_ARK_ARC_1_2/temp5[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[63] ), 
        .A2(n457), .Z(\MC_ARK_ARC_1_2/temp4[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_27_2  ( .A1(\RI5[2][189] ), .A2(\RI5[2][165] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_27_2  ( .A1(\RI5[2][27] ), .A2(\RI5[2][21] ), .Z(
        \MC_ARK_ARC_1_2/temp1[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_1  ( .A1(\SB2_2_22/buf_output[4] ), .A2(n168), 
        .Z(\MC_ARK_ARC_1_2/temp4[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .A2(n154), .Z(\MC_ARK_ARC_1_2/temp4[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_27_0  ( .A1(\RI5[2][95] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[131] ), .Z(\MC_ARK_ARC_1_2/temp3[29] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_27_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[23] ), .Z(\MC_ARK_ARC_1_2/temp1[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_26_5  ( .A1(\MC_ARK_ARC_1_2/temp6[30] ), .A2(
        \MC_ARK_ARC_1_2/temp5[30] ), .Z(\MC_ARK_ARC_1_2/buf_output[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_26_5  ( .A1(\MC_ARK_ARC_1_2/temp3[30] ), .A2(
        \MC_ARK_ARC_1_2/temp4[30] ), .Z(\MC_ARK_ARC_1_2/temp6[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_5  ( .A1(\RI5[2][66] ), .A2(n204), .Z(
        \MC_ARK_ARC_1_2/temp4[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_26_5  ( .A1(\RI5[2][132] ), .A2(\RI5[2][96] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_26_5  ( .A1(\RI5[2][0] ), .A2(\RI5[2][168] ), .Z(
        \MC_ARK_ARC_1_2/temp2[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_26_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[24] ), 
        .A2(\RI5[2][30] ), .Z(\MC_ARK_ARC_1_2/temp1[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_26_4  ( .A1(\MC_ARK_ARC_1_2/temp3[31] ), .A2(
        \MC_ARK_ARC_1_2/temp4[31] ), .Z(\MC_ARK_ARC_1_2/temp6[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_26_4  ( .A1(\MC_ARK_ARC_1_2/temp1[31] ), .A2(
        \MC_ARK_ARC_1_2/temp2[31] ), .Z(\MC_ARK_ARC_1_2/temp5[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_4  ( .A1(\RI5[2][67] ), .A2(n434), .Z(
        \MC_ARK_ARC_1_2/temp4[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_26_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[133] ), 
        .A2(\RI5[2][97] ), .Z(\MC_ARK_ARC_1_2/temp3[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_26_4  ( .A1(\RI5[2][1] ), .A2(\RI5[2][169] ), .Z(
        \MC_ARK_ARC_1_2/temp2[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_26_4  ( .A1(\RI5[2][31] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[25] ), .Z(\MC_ARK_ARC_1_2/temp1[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), 
        .A2(n467), .Z(\MC_ARK_ARC_1_2/temp4[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_26_3  ( .A1(\RI5[2][170] ), .A2(\RI5[2][2] ), .Z(
        \MC_ARK_ARC_1_2/temp2[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_26_1  ( .A1(\MC_ARK_ARC_1_2/temp4[34] ), .A2(
        \MC_ARK_ARC_1_2/temp3[34] ), .Z(\MC_ARK_ARC_1_2/temp6[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[70] ), 
        .A2(n214), .Z(\MC_ARK_ARC_1_2/temp4[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_0  ( .A1(\RI5[2][71] ), .A2(n567), .Z(
        \MC_ARK_ARC_1_2/temp4[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_25_5  ( .A1(\MC_ARK_ARC_1_2/temp1[36] ), .A2(
        \MC_ARK_ARC_1_2/temp2[36] ), .Z(\MC_ARK_ARC_1_2/temp5[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_5  ( .A1(\RI5[2][72] ), .A2(n446), .Z(
        \MC_ARK_ARC_1_2/temp4[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_25_5  ( .A1(\SB2_2_13/buf_output[0] ), .A2(
        \RI5[2][102] ), .Z(\MC_ARK_ARC_1_2/temp3[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_25_5  ( .A1(\RI5[2][6] ), .A2(\RI5[2][174] ), .Z(
        \MC_ARK_ARC_1_2/temp2[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_25_5  ( .A1(\RI5[2][30] ), .A2(\RI5[2][36] ), .Z(
        \MC_ARK_ARC_1_2/temp1[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_25_4  ( .A1(\MC_ARK_ARC_1_2/temp3[37] ), .A2(
        \MC_ARK_ARC_1_2/temp4[37] ), .Z(\MC_ARK_ARC_1_2/temp6[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_25_4  ( .A1(\MC_ARK_ARC_1_2/temp1[37] ), .A2(
        \MC_ARK_ARC_1_2/temp2[37] ), .Z(\MC_ARK_ARC_1_2/temp5[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_4  ( .A1(\RI5[2][73] ), .A2(n69), .Z(
        \MC_ARK_ARC_1_2/temp4[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_25_4  ( .A1(\RI5[2][139] ), .A2(\RI5[2][103] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_25_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .A2(\RI5[2][175] ), .Z(\MC_ARK_ARC_1_2/temp2[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_25_4  ( .A1(\RI5[2][37] ), .A2(\RI5[2][31] ), .Z(
        \MC_ARK_ARC_1_2/temp1[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[74] ), 
        .A2(n510), .Z(\MC_ARK_ARC_1_2/temp4[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_25_3  ( .A1(\RI5[2][104] ), .A2(\RI5[2][140] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_2  ( .A1(\RI5[2][75] ), .A2(n544), .Z(
        \MC_ARK_ARC_1_2/temp4[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_25_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[141] ), 
        .A2(\RI5[2][105] ), .Z(\MC_ARK_ARC_1_2/temp3[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_1  ( .A1(\RI5[2][76] ), .A2(n421), .Z(
        \MC_ARK_ARC_1_2/temp4[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_25_1  ( .A1(\RI5[2][142] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[106] ), .Z(\MC_ARK_ARC_1_2/temp3[40] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_25_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[10] ), 
        .A2(\RI5[2][178] ), .Z(\MC_ARK_ARC_1_2/temp2[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_25_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[40] ), 
        .A2(\RI5[2][34] ), .Z(\MC_ARK_ARC_1_2/temp1[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_24_5  ( .A1(\MC_ARK_ARC_1_2/temp6[42] ), .A2(
        \MC_ARK_ARC_1_2/temp5[42] ), .Z(\MC_ARK_ARC_1_2/buf_output[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_24_5  ( .A1(\MC_ARK_ARC_1_2/temp1[42] ), .A2(
        \MC_ARK_ARC_1_2/temp2[42] ), .Z(\MC_ARK_ARC_1_2/temp5[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_5  ( .A1(\RI5[2][78] ), .A2(n489), .Z(
        \MC_ARK_ARC_1_2/temp4[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_24_5  ( .A1(\RI5[2][12] ), .A2(\RI5[2][180] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_24_5  ( .A1(\RI5[2][42] ), .A2(\RI5[2][36] ), .Z(
        \MC_ARK_ARC_1_2/temp1[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[79] ), 
        .A2(n199), .Z(\MC_ARK_ARC_1_2/temp4[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_24_4  ( .A1(\RI5[2][109] ), .A2(\RI5[2][145] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_24_4  ( .A1(\RI5[2][43] ), .A2(\RI5[2][37] ), .Z(
        \MC_ARK_ARC_1_2/temp1[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_24_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[14] ), 
        .A2(\RI5[2][182] ), .Z(\MC_ARK_ARC_1_2/temp2[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_24_2  ( .A1(\MC_ARK_ARC_1_2/temp2[45] ), .A2(
        \MC_ARK_ARC_1_2/temp1[45] ), .Z(\MC_ARK_ARC_1_2/temp5[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_2  ( .A1(\RI5[2][81] ), .A2(n119), .Z(
        \MC_ARK_ARC_1_2/temp4[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_24_2  ( .A1(\RI5[2][15] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[183] ), .Z(\MC_ARK_ARC_1_2/temp2[45] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_24_1  ( .A1(\MC_ARK_ARC_1_2/temp3[46] ), .A2(
        \MC_ARK_ARC_1_2/temp4[46] ), .Z(\MC_ARK_ARC_1_2/temp6[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_1  ( .A1(\RI5[2][82] ), .A2(n466), .Z(
        \MC_ARK_ARC_1_2/temp4[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_24_1  ( .A1(\RI5[2][148] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[112] ), .Z(\MC_ARK_ARC_1_2/temp3[46] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_24_1  ( .A1(\RI5[2][16] ), .A2(\RI5[2][184] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_24_1  ( .A1(\RI5[2][46] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[40] ), .Z(\MC_ARK_ARC_1_2/temp1[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_0  ( .A1(\RI5[2][83] ), .A2(n498), .Z(
        \MC_ARK_ARC_1_2/temp4[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_24_0  ( .A1(\RI5[2][17] ), .A2(\RI5[2][185] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_24_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[41] ), 
        .A2(\RI5[2][47] ), .Z(\MC_ARK_ARC_1_2/temp1[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_23_5  ( .A1(\MC_ARK_ARC_1_2/temp5[48] ), .A2(
        \MC_ARK_ARC_1_2/temp6[48] ), .Z(\MC_ARK_ARC_1_2/buf_output[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_5  ( .A1(\SB2_2_22/buf_output[0] ), .A2(n198), 
        .Z(\MC_ARK_ARC_1_2/temp4[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_23_5  ( .A1(\RI5[2][18] ), .A2(\RI5[2][186] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_4  ( .A1(\RI5[2][85] ), .A2(n565), .Z(
        \MC_ARK_ARC_1_2/temp4[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_23_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[115] ), .Z(
        \MC_ARK_ARC_1_2/temp3[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_23_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .A2(\RI5[2][43] ), .Z(\MC_ARK_ARC_1_2/temp1[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_3  ( .A1(\RI5[2][86] ), .A2(n444), .Z(
        \MC_ARK_ARC_1_2/temp4[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_23_2  ( .A1(\MC_ARK_ARC_1_2/temp3[51] ), .A2(
        \MC_ARK_ARC_1_2/temp4[51] ), .Z(\MC_ARK_ARC_1_2/temp6[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_2  ( .A1(\SB2_2_19/buf_output[3] ), .A2(n83), 
        .Z(\MC_ARK_ARC_1_2/temp4[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_23_1  ( .A1(\MC_ARK_ARC_1_2/temp3[52] ), .A2(
        \MC_ARK_ARC_1_2/temp4[52] ), .Z(\MC_ARK_ARC_1_2/temp6[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_23_1  ( .A1(\MC_ARK_ARC_1_2/temp2[52] ), .A2(
        \MC_ARK_ARC_1_2/temp1[52] ), .Z(\MC_ARK_ARC_1_2/temp5[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_1  ( .A1(\RI5[2][88] ), .A2(n508), .Z(
        \MC_ARK_ARC_1_2/temp4[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_23_1  ( .A1(\RI5[2][154] ), .A2(\RI5[2][118] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_23_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[22] ), 
        .A2(\RI5[2][190] ), .Z(\MC_ARK_ARC_1_2/temp2[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_23_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .A2(\RI5[2][46] ), .Z(\MC_ARK_ARC_1_2/temp1[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[89] ), 
        .A2(n130), .Z(\MC_ARK_ARC_1_2/temp4[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_5  ( .A1(\RI5[2][90] ), .A2(n208), .Z(
        \MC_ARK_ARC_1_2/temp4[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_22_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[24] ), 
        .A2(\RI5[2][0] ), .Z(\MC_ARK_ARC_1_2/temp2[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_4  ( .A1(\RI5[2][91] ), .A2(n217), .Z(
        \MC_ARK_ARC_1_2/temp4[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_22_4  ( .A1(\RI5[2][1] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[25] ), .Z(\MC_ARK_ARC_1_2/temp2[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_22_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[55] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[49] ), .Z(\MC_ARK_ARC_1_2/temp1[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[92] ), 
        .A2(n212), .Z(\MC_ARK_ARC_1_2/temp4[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_22_3  ( .A1(\RI5[2][2] ), .A2(\RI5[2][26] ), .Z(
        \MC_ARK_ARC_1_2/temp2[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_22_3  ( .A1(\RI5[2][50] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[56] ), .Z(\MC_ARK_ARC_1_2/temp1[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_1  ( .A1(\RI5[2][94] ), .A2(n215), .Z(
        \MC_ARK_ARC_1_2/temp4[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_22_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[28] ), 
        .A2(\RI5[2][4] ), .Z(\MC_ARK_ARC_1_2/temp2[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_22_0  ( .A1(\RI5[2][59] ), .A2(\RI5[2][53] ), .Z(
        \MC_ARK_ARC_1_2/temp1[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_5  ( .A1(\RI5[2][96] ), .A2(n464), .Z(
        \MC_ARK_ARC_1_2/temp4[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_21_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .A2(\RI5[2][126] ), .Z(\MC_ARK_ARC_1_2/temp3[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_21_5  ( .A1(\RI5[2][30] ), .A2(\RI5[2][6] ), .Z(
        \MC_ARK_ARC_1_2/temp2[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_21_4  ( .A1(\MC_ARK_ARC_1_2/temp3[61] ), .A2(
        \MC_ARK_ARC_1_2/temp4[61] ), .Z(\MC_ARK_ARC_1_2/temp6[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_4  ( .A1(\RI5[2][97] ), .A2(n218), .Z(
        \MC_ARK_ARC_1_2/temp4[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_21_4  ( .A1(\RI5[2][31] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[7] ), .Z(\MC_ARK_ARC_1_2/temp2[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_21_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[55] ), .Z(\MC_ARK_ARC_1_2/temp1[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_21_3  ( .A1(\MC_ARK_ARC_1_2/temp3[62] ), .A2(
        \MC_ARK_ARC_1_2/temp4[62] ), .Z(\MC_ARK_ARC_1_2/temp6[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[98] ), 
        .A2(n185), .Z(\MC_ARK_ARC_1_2/temp4[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_21_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[164] ), 
        .A2(\RI5[2][128] ), .Z(\MC_ARK_ARC_1_2/temp3[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_21_3  ( .A1(\RI5[2][8] ), .A2(\RI5[2][32] ), .Z(
        \MC_ARK_ARC_1_2/temp2[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_21_3  ( .A1(\RI5[2][62] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[56] ), .Z(\MC_ARK_ARC_1_2/temp1[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_21_2  ( .A1(\MC_ARK_ARC_1_2/temp3[63] ), .A2(
        \MC_ARK_ARC_1_2/temp4[63] ), .Z(\MC_ARK_ARC_1_2/temp6[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), 
        .A2(n563), .Z(\MC_ARK_ARC_1_2/temp4[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_21_1  ( .A1(\MC_ARK_ARC_1_2/temp1[64] ), .A2(
        \MC_ARK_ARC_1_2/temp2[64] ), .Z(\MC_ARK_ARC_1_2/temp5[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[100] ), 
        .A2(n442), .Z(\MC_ARK_ARC_1_2/temp4[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_21_1  ( .A1(\RI5[2][166] ), .A2(\RI5[2][130] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_21_1  ( .A1(\RI5[2][34] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[10] ), .Z(\MC_ARK_ARC_1_2/temp2[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_21_1  ( .A1(\RI5[2][64] ), .A2(\RI5[2][58] ), .Z(
        \MC_ARK_ARC_1_2/temp1[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_5  ( .A1(\RI5[2][102] ), .A2(n507), .Z(
        \MC_ARK_ARC_1_2/temp4[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_20_5  ( .A1(\RI5[2][168] ), .A2(\RI5[2][132] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_20_5  ( .A1(\RI5[2][36] ), .A2(\RI5[2][12] ), .Z(
        \MC_ARK_ARC_1_2/temp2[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_20_4  ( .A1(\MC_ARK_ARC_1_2/temp2[67] ), .A2(
        \MC_ARK_ARC_1_2/temp1[67] ), .Z(\MC_ARK_ARC_1_2/temp5[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_4  ( .A1(\RI5[2][103] ), .A2(n189), .Z(
        \MC_ARK_ARC_1_2/temp4[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_20_4  ( .A1(\RI5[2][13] ), .A2(\RI5[2][37] ), .Z(
        \MC_ARK_ARC_1_2/temp2[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_3  ( .A1(\RI5[2][104] ), .A2(n419), .Z(
        \MC_ARK_ARC_1_2/temp4[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_2  ( .A1(\RI5[2][105] ), .A2(n53), .Z(
        \MC_ARK_ARC_1_2/temp4[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_20_1  ( .A1(\MC_ARK_ARC_1_2/temp4[70] ), .A2(
        \MC_ARK_ARC_1_2/temp3[70] ), .Z(\MC_ARK_ARC_1_2/temp6[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .A2(\MC_ARK_ARC_1_1/buf_keyinput[111] ), .Z(\MC_ARK_ARC_1_2/temp4[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_20_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[172] ), 
        .A2(\RI5[2][136] ), .Z(\MC_ARK_ARC_1_2/temp3[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_20_1  ( .A1(\RI5[2][64] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[70] ), .Z(\MC_ARK_ARC_1_2/temp1[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_0  ( .A1(\RI5[2][107] ), .A2(n182), .Z(
        \MC_ARK_ARC_1_2/temp4[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_20_0  ( .A1(\RI5[2][173] ), .A2(\RI5[2][137] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_19_5  ( .A1(\MC_ARK_ARC_1_2/temp6[72] ), .A2(
        \MC_ARK_ARC_1_2/temp5[72] ), .Z(\MC_ARK_ARC_1_2/buf_output[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_19_5  ( .A1(\MC_ARK_ARC_1_2/temp3[72] ), .A2(
        \MC_ARK_ARC_1_2/temp4[72] ), .Z(\MC_ARK_ARC_1_2/temp6[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_19_5  ( .A1(\MC_ARK_ARC_1_2/temp2[72] ), .A2(
        \MC_ARK_ARC_1_2/temp1[72] ), .Z(\MC_ARK_ARC_1_2/temp5[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_5  ( .A1(\RI5[2][108] ), .A2(n551), .Z(
        \MC_ARK_ARC_1_2/temp4[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_19_5  ( .A1(\RI5[2][138] ), .A2(\RI5[2][174] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_19_5  ( .A1(\RI5[2][18] ), .A2(\RI5[2][42] ), .Z(
        \MC_ARK_ARC_1_2/temp2[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_19_5  ( .A1(\RI5[2][72] ), .A2(\RI5[2][66] ), .Z(
        \MC_ARK_ARC_1_2/temp1[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_19_4  ( .A1(\MC_ARK_ARC_1_2/temp2[73] ), .A2(
        \MC_ARK_ARC_1_2/temp1[73] ), .Z(\MC_ARK_ARC_1_2/temp5[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_4  ( .A1(\RI5[2][109] ), .A2(n184), .Z(
        \MC_ARK_ARC_1_2/temp4[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_19_4  ( .A1(\RI5[2][139] ), .A2(\RI5[2][175] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_19_4  ( .A1(\RI5[2][43] ), .A2(\RI5[2][19] ), .Z(
        \MC_ARK_ARC_1_2/temp2[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_19_4  ( .A1(\RI5[2][73] ), .A2(\RI5[2][67] ), .Z(
        \MC_ARK_ARC_1_2/temp1[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_2  ( .A1(\RI5[2][111] ), .A2(n495), .Z(
        \MC_ARK_ARC_1_2/temp4[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_19_1  ( .A1(\MC_ARK_ARC_1_2/temp6[76] ), .A2(
        \MC_ARK_ARC_1_2/temp5[76] ), .Z(\MC_ARK_ARC_1_2/buf_output[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_19_1  ( .A1(\MC_ARK_ARC_1_2/temp3[76] ), .A2(
        \MC_ARK_ARC_1_2/temp4[76] ), .Z(\MC_ARK_ARC_1_2/temp6[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_19_1  ( .A1(\MC_ARK_ARC_1_2/temp1[76] ), .A2(
        \MC_ARK_ARC_1_2/temp2[76] ), .Z(\MC_ARK_ARC_1_2/temp5[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[112] ), 
        .A2(n105), .Z(\MC_ARK_ARC_1_2/temp4[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_19_1  ( .A1(\RI5[2][178] ), .A2(\RI5[2][142] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_19_1  ( .A1(\RI5[2][46] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_2/temp2[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_19_1  ( .A1(\RI5[2][76] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[70] ), .Z(\MC_ARK_ARC_1_2/temp1[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_0  ( .A1(\RI5[2][113] ), .A2(n157), .Z(
        \MC_ARK_ARC_1_2/temp4[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_19_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[143] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[179] ), .Z(
        \MC_ARK_ARC_1_2/temp3[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_19_0  ( .A1(\RI5[2][77] ), .A2(\RI5[2][71] ), .Z(
        \MC_ARK_ARC_1_2/temp1[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_5  ( .A1(\RI5[2][114] ), .A2(n172), .Z(
        \MC_ARK_ARC_1_2/temp4[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_18_5  ( .A1(\RI5[2][180] ), .A2(\RI5[2][144] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_18_5  ( .A1(\RI5[2][72] ), .A2(\RI5[2][78] ), .Z(
        \MC_ARK_ARC_1_2/temp1[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_18_4  ( .A1(\MC_ARK_ARC_1_2/temp5[79] ), .A2(
        \MC_ARK_ARC_1_2/temp6[79] ), .Z(\MC_ARK_ARC_1_2/buf_output[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_18_4  ( .A1(\MC_ARK_ARC_1_2/temp3[79] ), .A2(
        \MC_ARK_ARC_1_2/temp4[79] ), .Z(\MC_ARK_ARC_1_2/temp6[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_18_4  ( .A1(\MC_ARK_ARC_1_2/temp2[79] ), .A2(
        \MC_ARK_ARC_1_2/temp1[79] ), .Z(\MC_ARK_ARC_1_2/temp5[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .A2(\MC_ARK_ARC_1_2/buf_keyinput[79] ), .Z(\MC_ARK_ARC_1_2/temp4[79] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_18_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[181] ), 
        .A2(\RI5[2][145] ), .Z(\MC_ARK_ARC_1_2/temp3[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_18_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[25] ), .Z(\MC_ARK_ARC_1_2/temp2[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_18_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[79] ), 
        .A2(\RI5[2][73] ), .Z(\MC_ARK_ARC_1_2/temp1[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_18_3  ( .A1(\MC_ARK_ARC_1_2/temp5[80] ), .A2(
        \MC_ARK_ARC_1_2/temp6[80] ), .Z(\MC_ARK_ARC_1_2/buf_output[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_3  ( .A1(\SB2_2_15/buf_output[2] ), .A2(n506), 
        .Z(\MC_ARK_ARC_1_2/temp4[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_18_3  ( .A1(\RI5[2][50] ), .A2(\RI5[2][26] ), .Z(
        \MC_ARK_ARC_1_2/temp2[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_18_2  ( .A1(\RI5[2][51] ), .A2(\RI5[2][27] ), .Z(
        \MC_ARK_ARC_1_2/temp2[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_18_2  ( .A1(\RI5[2][75] ), .A2(\RI5[2][81] ), .Z(
        \MC_ARK_ARC_1_2/temp1[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_18_1  ( .A1(\MC_ARK_ARC_1_2/temp6[82] ), .A2(
        \MC_ARK_ARC_1_2/temp5[82] ), .Z(\MC_ARK_ARC_1_2/buf_output[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_18_1  ( .A1(\MC_ARK_ARC_1_2/temp3[82] ), .A2(
        \MC_ARK_ARC_1_2/temp4[82] ), .Z(\MC_ARK_ARC_1_2/temp6[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_18_1  ( .A1(\MC_ARK_ARC_1_2/temp1[82] ), .A2(
        \MC_ARK_ARC_1_2/temp2[82] ), .Z(\MC_ARK_ARC_1_2/temp5[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_1  ( .A1(\RI5[2][118] ), .A2(n417), .Z(
        \MC_ARK_ARC_1_2/temp4[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_18_1  ( .A1(\RI5[2][148] ), .A2(\RI5[2][184] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_18_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[28] ), .Z(\MC_ARK_ARC_1_2/temp2[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_18_1  ( .A1(\RI5[2][82] ), .A2(\RI5[2][76] ), .Z(
        \MC_ARK_ARC_1_2/temp1[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_18_0  ( .A1(\MC_ARK_ARC_1_2/temp3[83] ), .A2(
        \MC_ARK_ARC_1_2/temp4[83] ), .Z(\MC_ARK_ARC_1_2/temp6[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_18_0  ( .A1(\MC_ARK_ARC_1_2/temp1[83] ), .A2(
        \MC_ARK_ARC_1_2/temp2[83] ), .Z(\MC_ARK_ARC_1_2/temp5[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_0  ( .A1(\RI5[2][119] ), .A2(n137), .Z(
        \MC_ARK_ARC_1_2/temp4[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_18_0  ( .A1(\RI5[2][149] ), .A2(\RI5[2][185] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_18_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .A2(\RI5[2][53] ), .Z(\MC_ARK_ARC_1_2/temp2[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_18_0  ( .A1(\RI5[2][77] ), .A2(\RI5[2][83] ), .Z(
        \MC_ARK_ARC_1_2/temp1[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_17_5  ( .A1(\MC_ARK_ARC_1_2/temp5[84] ), .A2(
        \MC_ARK_ARC_1_2/temp6[84] ), .Z(\MC_ARK_ARC_1_2/buf_output[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_17_5  ( .A1(\MC_ARK_ARC_1_2/temp3[84] ), .A2(
        \MC_ARK_ARC_1_2/temp4[84] ), .Z(\MC_ARK_ARC_1_2/temp6[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[120] ), 
        .A2(n120), .Z(\MC_ARK_ARC_1_2/temp4[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_17_5  ( .A1(\RI5[2][186] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[150] ), .Z(\MC_ARK_ARC_1_2/temp3[84] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_17_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[84] ), 
        .A2(\RI5[2][78] ), .Z(\MC_ARK_ARC_1_2/temp1[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[121] ), 
        .A2(n40), .Z(\MC_ARK_ARC_1_2/temp4[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_17_4  ( .A1(\RI5[2][187] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[151] ), .Z(\MC_ARK_ARC_1_2/temp3[85] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_17_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[55] ), 
        .A2(\RI5[2][31] ), .Z(\MC_ARK_ARC_1_2/temp2[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[122] ), 
        .A2(n550), .Z(\MC_ARK_ARC_1_2/temp4[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_17_3  ( .A1(\RI5[2][86] ), .A2(\RI5[2][80] ), .Z(
        \MC_ARK_ARC_1_2/temp1[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_2  ( .A1(\RI5[2][123] ), .A2(n39), .Z(
        \MC_ARK_ARC_1_2/temp4[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .A2(n461), .Z(\MC_ARK_ARC_1_2/temp4[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_17_1  ( .A1(\RI5[2][154] ), .A2(\RI5[2][190] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_17_1  ( .A1(\RI5[2][58] ), .A2(\RI5[2][34] ), .Z(
        \MC_ARK_ARC_1_2/temp2[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_17_1  ( .A1(\RI5[2][88] ), .A2(\RI5[2][82] ), .Z(
        \MC_ARK_ARC_1_2/temp1[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_0  ( .A1(\RI5[2][125] ), .A2(n22), .Z(
        \MC_ARK_ARC_1_2/temp4[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_17_0  ( .A1(\RI5[2][191] ), .A2(\RI5[2][155] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_5  ( .A1(\RI5[2][126] ), .A2(n528), .Z(
        \MC_ARK_ARC_1_2/temp4[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_16_5  ( .A1(\RI5[2][0] ), .A2(\RI5[2][156] ), .Z(
        \MC_ARK_ARC_1_2/temp3[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_16_4  ( .A1(\MC_ARK_ARC_1_2/temp5[91] ), .A2(
        \MC_ARK_ARC_1_2/temp6[91] ), .Z(\MC_ARK_ARC_1_2/buf_output[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_16_4  ( .A1(\MC_ARK_ARC_1_2/temp3[91] ), .A2(
        \MC_ARK_ARC_1_2/temp4[91] ), .Z(\MC_ARK_ARC_1_2/temp6[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_4  ( .A1(\RI5[2][127] ), .A2(n103), .Z(
        \MC_ARK_ARC_1_2/temp4[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_16_4  ( .A1(\RI5[2][157] ), .A2(\RI5[2][1] ), .Z(
        \MC_ARK_ARC_1_2/temp3[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_16_4  ( .A1(\RI5[2][37] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[61] ), .Z(\MC_ARK_ARC_1_2/temp2[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_16_4  ( .A1(\RI5[2][85] ), .A2(\RI5[2][91] ), .Z(
        \MC_ARK_ARC_1_2/temp1[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_16_3  ( .A1(\RI5[2][62] ), .A2(\RI5[2][38] ), .Z(
        \MC_ARK_ARC_1_2/temp2[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_2  ( .A1(\RI5[2][129] ), .A2(n472), .Z(
        \MC_ARK_ARC_1_2/temp4[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_16_2  ( .A1(\RI5[2][93] ), .A2(\RI5[2][87] ), .Z(
        \MC_ARK_ARC_1_2/temp1[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_16_1  ( .A1(\MC_ARK_ARC_1_2/temp3[94] ), .A2(
        \MC_ARK_ARC_1_2/temp4[94] ), .Z(\MC_ARK_ARC_1_2/temp6[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_1  ( .A1(\RI5[2][130] ), .A2(n190), .Z(
        \MC_ARK_ARC_1_2/temp4[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_16_1  ( .A1(\RI5[2][4] ), .A2(\RI5[2][160] ), .Z(
        \MC_ARK_ARC_1_2/temp3[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_16_1  ( .A1(\RI5[2][64] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[40] ), .Z(\MC_ARK_ARC_1_2/temp2[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_16_1  ( .A1(\RI5[2][94] ), .A2(\RI5[2][88] ), .Z(
        \MC_ARK_ARC_1_2/temp1[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_16_0  ( .A1(\MC_ARK_ARC_1_2/temp5[95] ), .A2(
        \MC_ARK_ARC_1_2/temp6[95] ), .Z(\MC_ARK_ARC_1_2/buf_output[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_16_0  ( .A1(\MC_ARK_ARC_1_2/temp4[95] ), .A2(
        \MC_ARK_ARC_1_2/temp3[95] ), .Z(\MC_ARK_ARC_1_2/temp6[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .A2(n538), .Z(\MC_ARK_ARC_1_2/temp4[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_16_0  ( .A1(\RI5[2][5] ), .A2(\RI5[2][161] ), .Z(
        \MC_ARK_ARC_1_2/temp3[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_16_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[41] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[65] ), .Z(\MC_ARK_ARC_1_2/temp2[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_15_5  ( .A1(\RI5[2][132] ), .A2(n415), .Z(
        \MC_ARK_ARC_1_2/temp4[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_15_5  ( .A1(\RI5[2][6] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[162] ), .Z(\MC_ARK_ARC_1_2/temp3[96] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_15_5  ( .A1(\RI5[2][90] ), .A2(\RI5[2][96] ), .Z(
        \MC_ARK_ARC_1_2/temp1[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_15_4  ( .A1(\MC_ARK_ARC_1_2/temp2[97] ), .A2(
        \MC_ARK_ARC_1_2/temp1[97] ), .Z(\MC_ARK_ARC_1_2/temp5[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_15_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[133] ), 
        .A2(n219), .Z(\MC_ARK_ARC_1_2/temp4[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_15_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .A2(\RI5[2][163] ), .Z(\MC_ARK_ARC_1_2/temp3[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_15_4  ( .A1(\RI5[2][67] ), .A2(\RI5[2][43] ), .Z(
        \MC_ARK_ARC_1_2/temp2[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_15_4  ( .A1(\RI5[2][97] ), .A2(\RI5[2][91] ), .Z(
        \MC_ARK_ARC_1_2/temp1[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_15_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), 
        .A2(\RI5[2][44] ), .Z(\MC_ARK_ARC_1_2/temp2[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_15_2  ( .A1(\RI5[2][135] ), .A2(n121), .Z(
        \MC_ARK_ARC_1_2/temp4[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_15_1  ( .A1(\MC_ARK_ARC_1_2/temp1[100] ), .A2(
        \MC_ARK_ARC_1_2/temp2[100] ), .Z(\MC_ARK_ARC_1_2/temp5[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_15_1  ( .A1(\RI5[2][136] ), .A2(n548), .Z(
        \MC_ARK_ARC_1_2/temp4[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_15_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[70] ), 
        .A2(\RI5[2][46] ), .Z(\MC_ARK_ARC_1_2/temp2[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_15_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[100] ), 
        .A2(\RI5[2][94] ), .Z(\MC_ARK_ARC_1_2/temp1[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_15_0  ( .A1(\RI5[2][137] ), .A2(n425), .Z(
        \MC_ARK_ARC_1_2/temp4[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_15_0  ( .A1(\RI5[2][95] ), .A2(\RI5[2][101] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_14_5  ( .A1(\MC_ARK_ARC_1_2/temp1[102] ), .A2(
        \MC_ARK_ARC_1_2/temp2[102] ), .Z(\MC_ARK_ARC_1_2/temp5[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_5  ( .A1(\RI5[2][138] ), .A2(n129), .Z(
        \MC_ARK_ARC_1_2/temp4[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_14_5  ( .A1(\RI5[2][12] ), .A2(\RI5[2][168] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_14_5  ( .A1(\RI5[2][72] ), .A2(\RI5[2][48] ), .Z(
        \MC_ARK_ARC_1_2/temp2[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_14_5  ( .A1(\RI5[2][96] ), .A2(\RI5[2][102] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_4  ( .A1(\RI5[2][139] ), .A2(n492), .Z(
        \MC_ARK_ARC_1_2/temp4[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_14_4  ( .A1(\RI5[2][73] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[49] ), .Z(\MC_ARK_ARC_1_2/temp2[103] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_14_4  ( .A1(\RI5[2][103] ), .A2(\RI5[2][97] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_3  ( .A1(\RI5[2][140] ), .A2(n526), .Z(
        \MC_ARK_ARC_1_2/temp4[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[141] ), 
        .A2(n95), .Z(\MC_ARK_ARC_1_2/temp4[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_14_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[171] ), 
        .A2(\RI5[2][15] ), .Z(\MC_ARK_ARC_1_2/temp3[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_14_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), 
        .A2(\RI5[2][105] ), .Z(\MC_ARK_ARC_1_2/temp1[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_14_1  ( .A1(\MC_ARK_ARC_1_2/temp3[106] ), .A2(
        \MC_ARK_ARC_1_2/temp4[106] ), .Z(\MC_ARK_ARC_1_2/temp6[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_1  ( .A1(\RI5[2][142] ), .A2(n437), .Z(
        \MC_ARK_ARC_1_2/temp4[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_14_1  ( .A1(\RI5[2][16] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[172] ), .Z(\MC_ARK_ARC_1_2/temp3[106] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_14_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .A2(\RI5[2][76] ), .Z(\MC_ARK_ARC_1_2/temp2[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_14_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[100] ), .Z(
        \MC_ARK_ARC_1_2/temp1[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[143] ), 
        .A2(n147), .Z(\MC_ARK_ARC_1_2/temp4[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_14_0  ( .A1(\RI5[2][77] ), .A2(\RI5[2][53] ), .Z(
        \MC_ARK_ARC_1_2/temp2[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_5  ( .A1(\RI5[2][144] ), .A2(n503), .Z(
        \MC_ARK_ARC_1_2/temp4[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_13_5  ( .A1(\RI5[2][18] ), .A2(\RI5[2][174] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_13_5  ( .A1(\RI5[2][108] ), .A2(\RI5[2][102] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_4  ( .A1(\RI5[2][145] ), .A2(n143), .Z(
        \MC_ARK_ARC_1_2/temp4[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_13_4  ( .A1(\RI5[2][175] ), .A2(\RI5[2][19] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_13_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[79] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[55] ), .Z(
        \MC_ARK_ARC_1_2/temp2[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_13_4  ( .A1(\RI5[2][109] ), .A2(\RI5[2][103] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[147] ), 
        .A2(n449), .Z(\MC_ARK_ARC_1_2/temp4[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_13_2  ( .A1(\RI5[2][57] ), .A2(\RI5[2][81] ), .Z(
        \MC_ARK_ARC_1_2/temp2[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_13_1  ( .A1(\MC_ARK_ARC_1_2/temp6[112] ), .A2(
        \MC_ARK_ARC_1_2/temp5[112] ), .Z(\MC_ARK_ARC_1_2/buf_output[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_13_1  ( .A1(\MC_ARK_ARC_1_2/temp3[112] ), .A2(
        \MC_ARK_ARC_1_2/temp4[112] ), .Z(\MC_ARK_ARC_1_2/temp6[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_13_1  ( .A1(\MC_ARK_ARC_1_2/temp2[112] ), .A2(
        \MC_ARK_ARC_1_2/temp1[112] ), .Z(\MC_ARK_ARC_1_2/temp5[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_1  ( .A1(\RI5[2][148] ), .A2(n60), .Z(
        \MC_ARK_ARC_1_2/temp4[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_13_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[22] ), 
        .A2(\RI5[2][178] ), .Z(\MC_ARK_ARC_1_2/temp3[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_13_1  ( .A1(\RI5[2][82] ), .A2(\RI5[2][58] ), .Z(
        \MC_ARK_ARC_1_2/temp2[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_13_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[112] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[106] ), .Z(
        \MC_ARK_ARC_1_2/temp1[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_0  ( .A1(\RI5[2][149] ), .A2(n138), .Z(
        \MC_ARK_ARC_1_2/temp4[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_12_5  ( .A1(\MC_ARK_ARC_1_2/temp3[114] ), .A2(
        \MC_ARK_ARC_1_2/temp4[114] ), .Z(\MC_ARK_ARC_1_2/temp6[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[150] ), 
        .A2(n546), .Z(\MC_ARK_ARC_1_2/temp4[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_12_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[24] ), 
        .A2(\RI5[2][180] ), .Z(\MC_ARK_ARC_1_2/temp3[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .A2(n124), .Z(\MC_ARK_ARC_1_2/temp4[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_12_4  ( .A1(\RI5[2][85] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[61] ), .Z(\MC_ARK_ARC_1_2/temp2[115] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_3  ( .A1(\RI5[2][152] ), .A2(n131), .Z(
        \MC_ARK_ARC_1_2/temp4[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_2  ( .A1(\RI5[2][153] ), .A2(n156), .Z(
        \MC_ARK_ARC_1_2/temp4[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_12_2  ( .A1(\RI5[2][27] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[183] ), .Z(\MC_ARK_ARC_1_2/temp3[117] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_12_1  ( .A1(\MC_ARK_ARC_1_2/temp2[118] ), .A2(
        \MC_ARK_ARC_1_2/temp1[118] ), .Z(\MC_ARK_ARC_1_2/temp5[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_1  ( .A1(\RI5[2][154] ), .A2(n197), .Z(
        \MC_ARK_ARC_1_2/temp4[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_12_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[112] ), 
        .A2(\RI5[2][118] ), .Z(\MC_ARK_ARC_1_2/temp1[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_0  ( .A1(\RI5[2][155] ), .A2(n556), .Z(
        \MC_ARK_ARC_1_2/temp4[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_11_5  ( .A1(\MC_ARK_ARC_1_2/temp5[120] ), .A2(
        \MC_ARK_ARC_1_2/temp6[120] ), .Z(\MC_ARK_ARC_1_2/buf_output[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_11_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[120] ), 
        .A2(\RI5[2][114] ), .Z(\MC_ARK_ARC_1_2/temp1[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_11_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[121] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[115] ), .Z(
        \MC_ARK_ARC_1_2/temp1[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_11_3  ( .A1(\MC_ARK_ARC_1_2/temp3[122] ), .A2(
        \MC_ARK_ARC_1_2/temp4[122] ), .Z(\MC_ARK_ARC_1_2/temp6[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_11_3  ( .A1(\RI5[2][158] ), .A2(n501), .Z(
        \MC_ARK_ARC_1_2/temp4[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_11_2  ( .A1(\RI5[2][159] ), .A2(n536), .Z(
        \MC_ARK_ARC_1_2/temp4[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_11_1  ( .A1(\RI5[2][160] ), .A2(n568), .Z(
        \MC_ARK_ARC_1_2/temp4[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_11_1  ( .A1(\RI5[2][34] ), .A2(\RI5[2][190] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_11_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[70] ), 
        .A2(\RI5[2][94] ), .Z(\MC_ARK_ARC_1_2/temp2[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_11_0  ( .A1(\MC_ARK_ARC_1_2/temp3[125] ), .A2(
        \MC_ARK_ARC_1_2/temp4[125] ), .Z(\MC_ARK_ARC_1_2/temp6[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_11_0  ( .A1(\RI5[2][161] ), .A2(n447), .Z(
        \MC_ARK_ARC_1_2/temp4[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_11_0  ( .A1(\RI5[2][191] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[35] ), .Z(\MC_ARK_ARC_1_2/temp3[125] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_10_5  ( .A1(\MC_ARK_ARC_1_2/temp3[126] ), .A2(
        \MC_ARK_ARC_1_2/temp4[126] ), .Z(\MC_ARK_ARC_1_2/temp6[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .A2(\MC_ARK_ARC_1_1/buf_keyinput[119] ), .Z(
        \MC_ARK_ARC_1_2/temp4[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_10_5  ( .A1(\RI5[2][0] ), .A2(\RI5[2][36] ), .Z(
        \MC_ARK_ARC_1_2/temp3[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_10_5  ( .A1(\RI5[2][96] ), .A2(\RI5[2][72] ), .Z(
        \MC_ARK_ARC_1_2/temp2[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_4  ( .A1(\RI5[2][163] ), .A2(n106), .Z(
        \MC_ARK_ARC_1_2/temp4[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_10_4  ( .A1(\RI5[2][97] ), .A2(\RI5[2][73] ), .Z(
        \MC_ARK_ARC_1_2/temp2[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_10_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[121] ), 
        .A2(\RI5[2][127] ), .Z(\MC_ARK_ARC_1_2/temp1[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_10_3  ( .A1(\MC_ARK_ARC_1_2/temp3[128] ), .A2(
        \MC_ARK_ARC_1_2/temp4[128] ), .Z(\MC_ARK_ARC_1_2/temp6[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[164] ), 
        .A2(n545), .Z(\MC_ARK_ARC_1_2/temp4[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_10_3  ( .A1(\RI5[2][2] ), .A2(\RI5[2][38] ), .Z(
        \MC_ARK_ARC_1_2/temp3[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_2  ( .A1(\RI5[2][165] ), .A2(n111), .Z(
        \MC_ARK_ARC_1_2/temp4[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_10_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), 
        .A2(\RI5[2][75] ), .Z(\MC_ARK_ARC_1_2/temp2[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_10_1  ( .A1(\MC_ARK_ARC_1_2/temp5[130] ), .A2(
        \MC_ARK_ARC_1_2/temp6[130] ), .Z(\MC_ARK_ARC_1_2/buf_output[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_10_1  ( .A1(\MC_ARK_ARC_1_2/temp3[130] ), .A2(
        \MC_ARK_ARC_1_2/temp4[130] ), .Z(\MC_ARK_ARC_1_2/temp6[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_10_1  ( .A1(\MC_ARK_ARC_1_2/temp2[130] ), .A2(
        \MC_ARK_ARC_1_2/temp1[130] ), .Z(\MC_ARK_ARC_1_2/temp5[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_1  ( .A1(\RI5[2][166] ), .A2(n456), .Z(
        \MC_ARK_ARC_1_2/temp4[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_10_1  ( .A1(\RI5[2][4] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[40] ), .Z(\MC_ARK_ARC_1_2/temp3[130] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_10_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[100] ), 
        .A2(\RI5[2][76] ), .Z(\MC_ARK_ARC_1_2/temp2[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_10_1  ( .A1(\RI5[2][130] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[124] ), .Z(\MC_ARK_ARC_1_2/temp1[130] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_0  ( .A1(\RI5[2][167] ), .A2(n490), .Z(
        \MC_ARK_ARC_1_2/temp4[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_10_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[41] ), 
        .A2(\RI5[2][5] ), .Z(\MC_ARK_ARC_1_2/temp3[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_10_0  ( .A1(\RI5[2][101] ), .A2(\RI5[2][77] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_9_5  ( .A1(\MC_ARK_ARC_1_2/temp3[132] ), .A2(
        \MC_ARK_ARC_1_2/temp4[132] ), .Z(\MC_ARK_ARC_1_2/temp6[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_5  ( .A1(\RI5[2][168] ), .A2(n522), .Z(
        \MC_ARK_ARC_1_2/temp4[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_9_5  ( .A1(\RI5[2][132] ), .A2(\RI5[2][126] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_9_4  ( .A1(\MC_ARK_ARC_1_2/temp3[133] ), .A2(
        \MC_ARK_ARC_1_2/temp4[133] ), .Z(\MC_ARK_ARC_1_2/temp6[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_4  ( .A1(\RI5[2][169] ), .A2(n126), .Z(
        \MC_ARK_ARC_1_2/temp4[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_9_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .A2(\RI5[2][43] ), .Z(\MC_ARK_ARC_1_2/temp3[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_9_4  ( .A1(\RI5[2][127] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[133] ), .Z(\MC_ARK_ARC_1_2/temp1[133] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_3  ( .A1(\RI5[2][170] ), .A2(n433), .Z(
        \MC_ARK_ARC_1_2/temp4[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_9_2  ( .A1(\MC_ARK_ARC_1_2/temp1[135] ), .A2(
        \MC_ARK_ARC_1_2/temp2[135] ), .Z(\MC_ARK_ARC_1_2/temp5[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[171] ), 
        .A2(n64), .Z(\MC_ARK_ARC_1_2/temp4[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_9_2  ( .A1(\RI5[2][9] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[45] ), .Z(\MC_ARK_ARC_1_2/temp3[135] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_9_2  ( .A1(\RI5[2][105] ), .A2(\RI5[2][81] ), .Z(
        \MC_ARK_ARC_1_2/temp2[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[172] ), 
        .A2(n116), .Z(\MC_ARK_ARC_1_2/temp4[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_9_1  ( .A1(\RI5[2][46] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[10] ), .Z(\MC_ARK_ARC_1_2/temp3[136] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_9_1  ( .A1(\RI5[2][82] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[106] ), .Z(\MC_ARK_ARC_1_2/temp2[136] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_9_1  ( .A1(\RI5[2][136] ), .A2(\RI5[2][130] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_0  ( .A1(\RI5[2][173] ), .A2(n177), .Z(
        \MC_ARK_ARC_1_2/temp4[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_9_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .A2(\RI5[2][137] ), .Z(\MC_ARK_ARC_1_2/temp1[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_8_5  ( .A1(\MC_ARK_ARC_1_2/temp5[138] ), .A2(
        \MC_ARK_ARC_1_2/temp6[138] ), .Z(\MC_ARK_ARC_1_2/buf_output[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_8_5  ( .A1(\MC_ARK_ARC_1_2/temp4[138] ), .A2(
        \MC_ARK_ARC_1_2/temp3[138] ), .Z(\MC_ARK_ARC_1_2/temp6[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_5  ( .A1(\RI5[2][174] ), .A2(n169), .Z(
        \MC_ARK_ARC_1_2/temp4[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_8_5  ( .A1(\RI5[2][12] ), .A2(\RI5[2][48] ), .Z(
        \MC_ARK_ARC_1_2/temp3[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_8_4  ( .A1(\MC_ARK_ARC_1_2/temp5[139] ), .A2(
        \MC_ARK_ARC_1_2/temp6[139] ), .Z(\MC_ARK_ARC_1_2/buf_output[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_8_4  ( .A1(\RI5[2][139] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[133] ), .Z(\MC_ARK_ARC_1_2/temp1[139] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_3  ( .A1(\RI5[2][176] ), .A2(n479), .Z(
        \MC_ARK_ARC_1_2/temp4[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_8_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[110] ), 
        .A2(\RI5[2][86] ), .Z(\MC_ARK_ARC_1_2/temp2[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_8_2  ( .A1(\MC_ARK_ARC_1_2/temp3[141] ), .A2(
        \MC_ARK_ARC_1_2/temp4[141] ), .Z(\MC_ARK_ARC_1_2/temp6[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_2  ( .A1(\RI5[2][177] ), .A2(n16), .Z(
        \MC_ARK_ARC_1_2/temp4[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_8_2  ( .A1(\RI5[2][87] ), .A2(\RI5[2][111] ), .Z(
        \MC_ARK_ARC_1_2/temp2[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_8_2  ( .A1(\RI5[2][135] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_2/temp1[141] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_8_1  ( .A1(\MC_ARK_ARC_1_2/temp2[142] ), .A2(
        \MC_ARK_ARC_1_2/temp1[142] ), .Z(\MC_ARK_ARC_1_2/temp5[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_1  ( .A1(\RI5[2][178] ), .A2(n543), .Z(
        \MC_ARK_ARC_1_2/temp4[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_8_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[52] ), 
        .A2(\RI5[2][16] ), .Z(\MC_ARK_ARC_1_2/temp3[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_8_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[112] ), 
        .A2(\RI5[2][88] ), .Z(\MC_ARK_ARC_1_2/temp2[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_8_1  ( .A1(\RI5[2][142] ), .A2(\RI5[2][136] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_8_0  ( .A1(\MC_ARK_ARC_1_2/temp5[143] ), .A2(
        \MC_ARK_ARC_1_2/temp6[143] ), .Z(\MC_ARK_ARC_1_2/buf_output[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_8_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[143] ), 
        .A2(\RI5[2][137] ), .Z(\MC_ARK_ARC_1_2/temp1[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_7_5  ( .A1(\MC_ARK_ARC_1_2/temp3[144] ), .A2(
        \MC_ARK_ARC_1_2/temp4[144] ), .Z(\MC_ARK_ARC_1_2/temp6[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_5  ( .A1(\RI5[2][180] ), .A2(n203), .Z(
        \MC_ARK_ARC_1_2/temp4[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_7_5  ( .A1(\RI5[2][54] ), .A2(\RI5[2][18] ), .Z(
        \MC_ARK_ARC_1_2/temp3[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[181] ), 
        .A2(n213), .Z(\MC_ARK_ARC_1_2/temp4[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_7_4  ( .A1(\RI5[2][19] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[55] ), .Z(\MC_ARK_ARC_1_2/temp3[145] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_7_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .A2(\RI5[2][91] ), .Z(\MC_ARK_ARC_1_2/temp2[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_7_4  ( .A1(\RI5[2][139] ), .A2(\RI5[2][145] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_3  ( .A1(\RI5[2][182] ), .A2(n521), .Z(
        \MC_ARK_ARC_1_2/temp4[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_7_3  ( .A1(\RI5[2][116] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[92] ), .Z(\MC_ARK_ARC_1_2/temp2[146] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_7_2  ( .A1(\MC_ARK_ARC_1_2/temp5[147] ), .A2(
        \MC_ARK_ARC_1_2/temp6[147] ), .Z(\MC_ARK_ARC_1_2/buf_output[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_7_2  ( .A1(\MC_ARK_ARC_1_2/temp3[147] ), .A2(
        \MC_ARK_ARC_1_2/temp4[147] ), .Z(\MC_ARK_ARC_1_2/temp6[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_2  ( .A1(\SB2_2_3/buf_output[3] ), .A2(n553), 
        .Z(\MC_ARK_ARC_1_2/temp4[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_7_2  ( .A1(\RI5[2][57] ), .A2(\RI5[2][21] ), .Z(
        \MC_ARK_ARC_1_2/temp3[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_7_1  ( .A1(\MC_ARK_ARC_1_2/temp5[148] ), .A2(
        \MC_ARK_ARC_1_2/temp6[148] ), .Z(\MC_ARK_ARC_1_2/buf_output[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_7_1  ( .A1(\MC_ARK_ARC_1_2/temp4[148] ), .A2(
        \MC_ARK_ARC_1_2/temp3[148] ), .Z(\MC_ARK_ARC_1_2/temp6[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_7_1  ( .A1(\MC_ARK_ARC_1_2/temp2[148] ), .A2(
        \MC_ARK_ARC_1_2/temp1[148] ), .Z(\MC_ARK_ARC_1_2/temp5[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_1  ( .A1(\RI5[2][184] ), .A2(n431), .Z(
        \MC_ARK_ARC_1_2/temp4[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_7_1  ( .A1(\RI5[2][58] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_2/temp3[148] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_7_1  ( .A1(\RI5[2][118] ), .A2(\RI5[2][94] ), .Z(
        \MC_ARK_ARC_1_2/temp2[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_7_1  ( .A1(\RI5[2][148] ), .A2(\RI5[2][142] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_7_0  ( .A1(\MC_ARK_ARC_1_2/temp1[149] ), .A2(
        \MC_ARK_ARC_1_2/temp2[149] ), .Z(\MC_ARK_ARC_1_2/temp5[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_0  ( .A1(\RI5[2][185] ), .A2(n465), .Z(
        \MC_ARK_ARC_1_2/temp4[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_7_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[23] ), 
        .A2(\RI5[2][59] ), .Z(\MC_ARK_ARC_1_2/temp3[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_7_0  ( .A1(\RI5[2][119] ), .A2(\RI5[2][95] ), .Z(
        \MC_ARK_ARC_1_2/temp2[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_7_0  ( .A1(\RI5[2][149] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[143] ), .Z(\MC_ARK_ARC_1_2/temp1[149] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_6_5  ( .A1(\MC_ARK_ARC_1_2/temp6[150] ), .A2(
        \MC_ARK_ARC_1_2/temp5[150] ), .Z(\MC_ARK_ARC_1_2/buf_output[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_6_5  ( .A1(\MC_ARK_ARC_1_2/temp3[150] ), .A2(
        \MC_ARK_ARC_1_2/temp4[150] ), .Z(\MC_ARK_ARC_1_2/temp6[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_6_5  ( .A1(\MC_ARK_ARC_1_2/temp2[150] ), .A2(
        \MC_ARK_ARC_1_2/temp1[150] ), .Z(\MC_ARK_ARC_1_2/temp5[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_5  ( .A1(\RI5[2][186] ), .A2(n497), .Z(
        \MC_ARK_ARC_1_2/temp4[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_6_5  ( .A1(\RI5[2][96] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[120] ), .Z(\MC_ARK_ARC_1_2/temp2[150] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_6_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[150] ), 
        .A2(\RI5[2][144] ), .Z(\MC_ARK_ARC_1_2/temp1[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_6_4  ( .A1(\MC_ARK_ARC_1_2/temp6[151] ), .A2(
        \MC_ARK_ARC_1_2/temp5[151] ), .Z(\MC_ARK_ARC_1_2/buf_output[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_4  ( .A1(\RI5[2][187] ), .A2(n181), .Z(
        \MC_ARK_ARC_1_2/temp4[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_6_4  ( .A1(\SB2_2_15/buf_output[1] ), .A2(
        \RI5[2][97] ), .Z(\MC_ARK_ARC_1_2/temp2[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_6_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .A2(\RI5[2][145] ), .Z(\MC_ARK_ARC_1_2/temp1[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_3  ( .A1(\RI5[2][188] ), .A2(n564), .Z(
        \MC_ARK_ARC_1_2/temp4[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_6_2  ( .A1(\RI5[2][123] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[99] ), .Z(\MC_ARK_ARC_1_2/temp2[153] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_1  ( .A1(\RI5[2][190] ), .A2(n81), .Z(
        \MC_ARK_ARC_1_2/temp4[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_5_5  ( .A1(\MC_ARK_ARC_1_2/temp3[156] ), .A2(
        \MC_ARK_ARC_1_2/temp4[156] ), .Z(\MC_ARK_ARC_1_2/temp6[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_5_5  ( .A1(\MC_ARK_ARC_1_2/temp1[156] ), .A2(
        \MC_ARK_ARC_1_2/temp2[156] ), .Z(\MC_ARK_ARC_1_2/temp5[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_5  ( .A1(\RI5[2][0] ), .A2(n201), .Z(
        \MC_ARK_ARC_1_2/temp4[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_5_5  ( .A1(\RI5[2][66] ), .A2(\RI5[2][30] ), .Z(
        \MC_ARK_ARC_1_2/temp3[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_5_5  ( .A1(\RI5[2][102] ), .A2(\RI5[2][126] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_5_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[150] ), 
        .A2(\RI5[2][156] ), .Z(\MC_ARK_ARC_1_2/temp1[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_5_4  ( .A1(\MC_ARK_ARC_1_2/temp1[157] ), .A2(
        \MC_ARK_ARC_1_2/temp2[157] ), .Z(\MC_ARK_ARC_1_2/temp5[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_4  ( .A1(\RI5[2][1] ), .A2(n195), .Z(
        \MC_ARK_ARC_1_2/temp4[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_5_4  ( .A1(\RI5[2][67] ), .A2(\RI5[2][31] ), .Z(
        \MC_ARK_ARC_1_2/temp3[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_5_4  ( .A1(\SB2_2_14/buf_output[1] ), .A2(
        \RI5[2][103] ), .Z(\MC_ARK_ARC_1_2/temp2[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_5_4  ( .A1(\RI5[2][157] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[151] ), .Z(\MC_ARK_ARC_1_2/temp1[157] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_3  ( .A1(\RI5[2][2] ), .A2(n454), .Z(
        \MC_ARK_ARC_1_2/temp4[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_5_2  ( .A1(\MC_ARK_ARC_1_2/temp3[159] ), .A2(
        \MC_ARK_ARC_1_2/temp4[159] ), .Z(\MC_ARK_ARC_1_2/temp6[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[3] ), 
        .A2(n488), .Z(\MC_ARK_ARC_1_2/temp4[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_5_2  ( .A1(\RI5[2][129] ), .A2(\RI5[2][105] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_5_1  ( .A1(\MC_ARK_ARC_1_2/temp5[160] ), .A2(
        \MC_ARK_ARC_1_2/temp6[160] ), .Z(\MC_ARK_ARC_1_2/buf_output[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_1  ( .A1(\RI5[2][4] ), .A2(n519), .Z(
        \MC_ARK_ARC_1_2/temp4[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_5_1  ( .A1(\RI5[2][34] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[70] ), .Z(\MC_ARK_ARC_1_2/temp3[160] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_5_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .A2(\RI5[2][130] ), .Z(\MC_ARK_ARC_1_2/temp2[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_0  ( .A1(\RI5[2][5] ), .A2(n552), .Z(
        \MC_ARK_ARC_1_2/temp4[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_5  ( .A1(\SB2_2_3/buf_output[0] ), .A2(n429), 
        .Z(\MC_ARK_ARC_1_2/temp4[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .A2(n134), .Z(\MC_ARK_ARC_1_2/temp4[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_4_4  ( .A1(\RI5[2][73] ), .A2(\RI5[2][37] ), .Z(
        \MC_ARK_ARC_1_2/temp3[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_4_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[133] ), 
        .A2(\RI5[2][109] ), .Z(\MC_ARK_ARC_1_2/temp2[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_4_4  ( .A1(\RI5[2][157] ), .A2(\RI5[2][163] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_3  ( .A1(\RI5[2][8] ), .A2(n496), .Z(
        \MC_ARK_ARC_1_2/temp4[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_4_2  ( .A1(\MC_ARK_ARC_1_2/temp4[165] ), .A2(
        \MC_ARK_ARC_1_2/temp3[165] ), .Z(\MC_ARK_ARC_1_2/temp6[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_2  ( .A1(\RI5[2][9] ), .A2(n531), .Z(
        \MC_ARK_ARC_1_2/temp4[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_4_2  ( .A1(\RI5[2][39] ), .A2(\RI5[2][75] ), .Z(
        \MC_ARK_ARC_1_2/temp3[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_4_2  ( .A1(\RI5[2][111] ), .A2(\RI5[2][135] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_4_2  ( .A1(\RI5[2][159] ), .A2(\RI5[2][165] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_4_1  ( .A1(\MC_ARK_ARC_1_2/temp3[166] ), .A2(
        \MC_ARK_ARC_1_2/temp4[166] ), .Z(\MC_ARK_ARC_1_2/temp6[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[10] ), 
        .A2(n193), .Z(\MC_ARK_ARC_1_2/temp4[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_4_1  ( .A1(\RI5[2][76] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[40] ), .Z(\MC_ARK_ARC_1_2/temp3[166] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_4_1  ( .A1(\RI5[2][166] ), .A2(\RI5[2][160] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_4_0  ( .A1(\MC_ARK_ARC_1_2/temp3[167] ), .A2(
        \MC_ARK_ARC_1_2/temp4[167] ), .Z(\MC_ARK_ARC_1_2/temp6[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_0  ( .A1(\RI5[2][11] ), .A2(n441), .Z(
        \MC_ARK_ARC_1_2/temp4[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_4_0  ( .A1(\RI5[2][167] ), .A2(\RI5[2][161] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_3_5  ( .A1(\MC_ARK_ARC_1_2/temp4[168] ), .A2(
        \MC_ARK_ARC_1_2/temp3[168] ), .Z(\MC_ARK_ARC_1_2/temp6[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_5  ( .A1(\RI5[2][12] ), .A2(n475), .Z(
        \MC_ARK_ARC_1_2/temp4[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_3_5  ( .A1(\RI5[2][78] ), .A2(\RI5[2][42] ), .Z(
        \MC_ARK_ARC_1_2/temp3[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_3_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .A2(\RI5[2][168] ), .Z(\MC_ARK_ARC_1_2/temp1[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_3_4  ( .A1(\MC_ARK_ARC_1_2/temp3[169] ), .A2(
        \MC_ARK_ARC_1_2/temp4[169] ), .Z(\MC_ARK_ARC_1_2/temp6[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_4  ( .A1(\RI5[2][13] ), .A2(n200), .Z(
        \MC_ARK_ARC_1_2/temp4[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_3_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .A2(\RI5[2][139] ), .Z(\MC_ARK_ARC_1_2/temp2[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_3_3  ( .A1(\MC_ARK_ARC_1_2/temp6[170] ), .A2(
        \MC_ARK_ARC_1_2/temp5[170] ), .Z(\MC_ARK_ARC_1_2/buf_output[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_3_2  ( .A1(\MC_ARK_ARC_1_2/temp5[171] ), .A2(
        \MC_ARK_ARC_1_2/temp6[171] ), .Z(\MC_ARK_ARC_1_2/buf_output[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_2  ( .A1(\RI5[2][15] ), .A2(n418), .Z(
        \MC_ARK_ARC_1_2/temp4[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_3_2  ( .A1(\RI5[2][117] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_2/temp2[171] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_3_1  ( .A1(\MC_ARK_ARC_1_2/temp4[172] ), .A2(
        \MC_ARK_ARC_1_2/temp3[172] ), .Z(\MC_ARK_ARC_1_2/temp6[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_1  ( .A1(\RI5[2][16] ), .A2(n1), .Z(
        \MC_ARK_ARC_1_2/temp4[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_3_1  ( .A1(\RI5[2][82] ), .A2(\RI5[2][46] ), .Z(
        \MC_ARK_ARC_1_2/temp3[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_0  ( .A1(\RI5[2][17] ), .A2(n487), .Z(
        \MC_ARK_ARC_1_2/temp4[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_3_0  ( .A1(\RI5[2][167] ), .A2(\RI5[2][173] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_2_5  ( .A1(\MC_ARK_ARC_1_2/temp3[174] ), .A2(
        \MC_ARK_ARC_1_2/temp4[174] ), .Z(\MC_ARK_ARC_1_2/temp6[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_5  ( .A1(\RI5[2][18] ), .A2(n110), .Z(
        \MC_ARK_ARC_1_2/temp4[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_2_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[84] ), 
        .A2(\RI5[2][48] ), .Z(\MC_ARK_ARC_1_2/temp3[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_2_5  ( .A1(\RI5[2][174] ), .A2(\RI5[2][168] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_4  ( .A1(\RI5[2][19] ), .A2(n188), .Z(
        \MC_ARK_ARC_1_2/temp4[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_2_4  ( .A1(\RI5[2][175] ), .A2(\RI5[2][169] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_2_3  ( .A1(\MC_ARK_ARC_1_2/temp1[176] ), .A2(
        \MC_ARK_ARC_1_2/temp2[176] ), .Z(\MC_ARK_ARC_1_2/temp5[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_2_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[122] ), .Z(
        \MC_ARK_ARC_1_2/temp2[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_2  ( .A1(\RI5[2][21] ), .A2(n55), .Z(
        \MC_ARK_ARC_1_2/temp4[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_2_2  ( .A1(\SB2_2_13/buf_output[3] ), .A2(
        \SB2_2_9/buf_output[3] ), .Z(\MC_ARK_ARC_1_2/temp2[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[22] ), 
        .A2(n99), .Z(\MC_ARK_ARC_1_2/temp4[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_2_1  ( .A1(\RI5[2][148] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[124] ), .Z(\MC_ARK_ARC_1_2/temp2[178] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_2_1  ( .A1(\RI5[2][178] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[172] ), .Z(\MC_ARK_ARC_1_2/temp1[178] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[24] ), 
        .A2(n133), .Z(\MC_ARK_ARC_1_2/temp4[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_1_5  ( .A1(\RI5[2][126] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[150] ), .Z(\MC_ARK_ARC_1_2/temp2[180] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_1_5  ( .A1(\RI5[2][180] ), .A2(\RI5[2][174] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_1_4  ( .A1(\MC_ARK_ARC_1_2/temp2[181] ), .A2(
        \MC_ARK_ARC_1_2/temp1[181] ), .Z(\MC_ARK_ARC_1_2/temp5[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_4  ( .A1(\SB2_2_31/buf_output[1] ), .A2(n440), 
        .Z(\MC_ARK_ARC_1_2/temp4[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_1_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[181] ), 
        .A2(\RI5[2][175] ), .Z(\MC_ARK_ARC_1_2/temp1[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_3  ( .A1(\RI5[2][26] ), .A2(n159), .Z(
        \MC_ARK_ARC_1_2/temp4[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_1_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[92] ), .Z(
        \MC_ARK_ARC_1_2/temp3[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_1_3  ( .A1(\RI5[2][176] ), .A2(\RI5[2][182] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_2  ( .A1(\RI5[2][27] ), .A2(n505), .Z(
        \MC_ARK_ARC_1_2/temp4[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_1_1  ( .A1(\MC_ARK_ARC_1_2/temp5[184] ), .A2(
        \MC_ARK_ARC_1_2/temp6[184] ), .Z(\MC_ARK_ARC_1_2/buf_output[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_1_1  ( .A1(\MC_ARK_ARC_1_2/temp3[184] ), .A2(
        \MC_ARK_ARC_1_2/temp4[184] ), .Z(\MC_ARK_ARC_1_2/temp6[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[28] ), 
        .A2(n107), .Z(\MC_ARK_ARC_1_2/temp4[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_1_1  ( .A1(\RI5[2][94] ), .A2(\RI5[2][58] ), .Z(
        \MC_ARK_ARC_1_2/temp3[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_1_0  ( .A1(\MC_ARK_ARC_1_2/temp4[185] ), .A2(
        \MC_ARK_ARC_1_2/temp3[185] ), .Z(\MC_ARK_ARC_1_2/temp6[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .A2(\MC_ARK_ARC_1_1/buf_keyinput[148] ), .Z(
        \MC_ARK_ARC_1_2/temp4[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_1_0  ( .A1(\RI5[2][95] ), .A2(\RI5[2][59] ), .Z(
        \MC_ARK_ARC_1_2/temp3[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_1_0  ( .A1(\RI5[2][155] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[131] ), .Z(\MC_ARK_ARC_1_2/temp2[185] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_1_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[179] ), 
        .A2(\RI5[2][185] ), .Z(\MC_ARK_ARC_1_2/temp1[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_5  ( .A1(\RI5[2][30] ), .A2(n206), .Z(
        \MC_ARK_ARC_1_2/temp4[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_0_5  ( .A1(\SB2_2_26/buf_output[0] ), .A2(
        \RI5[2][96] ), .Z(\MC_ARK_ARC_1_2/temp3[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_4  ( .A1(\RI5[2][31] ), .A2(n191), .Z(
        \MC_ARK_ARC_1_2/temp4[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_0_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .A2(\RI5[2][97] ), .Z(\MC_ARK_ARC_1_2/temp3[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_0_3  ( .A1(\MC_ARK_ARC_1_2/temp3[188] ), .A2(
        \MC_ARK_ARC_1_2/temp4[188] ), .Z(\MC_ARK_ARC_1_2/temp6[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_0_3  ( .A1(\MC_ARK_ARC_1_2/temp1[188] ), .A2(
        \MC_ARK_ARC_1_2/temp2[188] ), .Z(\MC_ARK_ARC_1_2/temp5[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_3  ( .A1(\RI5[2][32] ), .A2(n194), .Z(
        \MC_ARK_ARC_1_2/temp4[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_0_3  ( .A1(\RI5[2][158] ), .A2(\RI5[2][134] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_0_3  ( .A1(\RI5[2][188] ), .A2(\RI5[2][182] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_2  ( .A1(\RI5[2][33] ), .A2(n186), .Z(
        \MC_ARK_ARC_1_2/temp4[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_0_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[63] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[99] ), .Z(
        \MC_ARK_ARC_1_2/temp3[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_0_2  ( .A1(\RI5[2][189] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[183] ), .Z(\MC_ARK_ARC_1_2/temp1[189] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_0_1  ( .A1(\MC_ARK_ARC_1_2/temp1[190] ), .A2(
        \MC_ARK_ARC_1_2/temp2[190] ), .Z(\MC_ARK_ARC_1_2/temp5[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_1  ( .A1(\RI5[2][34] ), .A2(n426), .Z(
        \MC_ARK_ARC_1_2/temp4[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_0_1  ( .A1(\RI5[2][64] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[100] ), .Z(\MC_ARK_ARC_1_2/temp3[190] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_0_1  ( .A1(\RI5[2][160] ), .A2(\RI5[2][136] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_0_0  ( .A1(\MC_ARK_ARC_1_2/temp1[191] ), .A2(
        \MC_ARK_ARC_1_2/temp2[191] ), .Z(\MC_ARK_ARC_1_2/temp5[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[35] ), 
        .A2(n460), .Z(\MC_ARK_ARC_1_2/temp4[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_0_0  ( .A1(\RI5[2][161] ), .A2(\RI5[2][137] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_31_5  ( .A1(\MC_ARK_ARC_1_3/temp2[0] ), .A2(
        \MC_ARK_ARC_1_3/temp1[0] ), .Z(\MC_ARK_ARC_1_3/temp5[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_5  ( .A1(\RI5[3][36] ), .A2(n207), .Z(
        \MC_ARK_ARC_1_3/temp4[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_31_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[102] ), 
        .A2(\RI5[3][66] ), .Z(\MC_ARK_ARC_1_3/temp3[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_31_4  ( .A1(\MC_ARK_ARC_1_3/temp3[1] ), .A2(
        \MC_ARK_ARC_1_3/temp4[1] ), .Z(\MC_ARK_ARC_1_3/temp6[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[37] ), 
        .A2(n424), .Z(\MC_ARK_ARC_1_3/temp4[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_31_4  ( .A1(\RI5[3][67] ), .A2(\RI5[3][103] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_31_4  ( .A1(\RI5[3][139] ), .A2(\RI5[3][163] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_31_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[1] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[187] ), .Z(\MC_ARK_ARC_1_3/temp1[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_31_3  ( .A1(\MC_ARK_ARC_1_3/temp6[2] ), .A2(
        \MC_ARK_ARC_1_3/temp5[2] ), .Z(\MC_ARK_ARC_1_3/buf_output[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_31_3  ( .A1(\MC_ARK_ARC_1_3/temp1[2] ), .A2(
        \MC_ARK_ARC_1_3/temp2[2] ), .Z(\MC_ARK_ARC_1_3/temp5[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_3  ( .A1(\RI5[3][38] ), .A2(n502), .Z(
        \MC_ARK_ARC_1_3/temp4[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_31_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[164] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[140] ), .Z(\MC_ARK_ARC_1_3/temp2[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_31_3  ( .A1(n1506), .A2(\RI5[3][2] ), .Z(
        \MC_ARK_ARC_1_3/temp1[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[39] ), 
        .A2(n216), .Z(\MC_ARK_ARC_1_3/temp4[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_31_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[105] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[69] ), .Z(\MC_ARK_ARC_1_3/temp3[3] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_31_2  ( .A1(\RI5[3][189] ), .A2(\RI5[3][3] ), .Z(
        \MC_ARK_ARC_1_3/temp1[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_31_1  ( .A1(\MC_ARK_ARC_1_3/temp5[4] ), .A2(
        \MC_ARK_ARC_1_3/temp6[4] ), .Z(\MC_ARK_ARC_1_3/buf_output[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_31_1  ( .A1(\MC_ARK_ARC_1_3/temp3[4] ), .A2(
        \MC_ARK_ARC_1_3/temp4[4] ), .Z(\MC_ARK_ARC_1_3/temp6[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_31_1  ( .A1(\MC_ARK_ARC_1_3/temp2[4] ), .A2(
        \MC_ARK_ARC_1_3/temp1[4] ), .Z(\MC_ARK_ARC_1_3/temp5[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_1  ( .A1(\RI5[3][40] ), .A2(n500), .Z(
        \MC_ARK_ARC_1_3/temp4[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_31_1  ( .A1(\RI5[3][106] ), .A2(\RI5[3][70] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_31_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .A2(\RI5[3][166] ), .Z(\MC_ARK_ARC_1_3/temp2[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_31_0  ( .A1(\RI5[3][167] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[143] ), .Z(\MC_ARK_ARC_1_3/temp2[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_30_5  ( .A1(\MC_ARK_ARC_1_3/temp6[6] ), .A2(
        \MC_ARK_ARC_1_3/temp5[6] ), .Z(\MC_ARK_ARC_1_3/buf_output[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_30_5  ( .A1(\MC_ARK_ARC_1_3/temp1[6] ), .A2(
        \MC_ARK_ARC_1_3/temp2[6] ), .Z(\MC_ARK_ARC_1_3/temp5[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_5  ( .A1(\RI5[3][42] ), .A2(n196), .Z(
        \MC_ARK_ARC_1_3/temp4[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_30_5  ( .A1(\RI5[3][108] ), .A2(\RI5[3][72] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_30_5  ( .A1(\RI5[3][168] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[144] ), .Z(\MC_ARK_ARC_1_3/temp2[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_30_5  ( .A1(\RI5[3][6] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[0] ), .Z(\MC_ARK_ARC_1_3/temp1[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[43] ), 
        .A2(n9), .Z(\MC_ARK_ARC_1_3/temp4[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_30_3  ( .A1(\MC_ARK_ARC_1_3/temp2[8] ), .A2(
        \MC_ARK_ARC_1_3/temp1[8] ), .Z(\MC_ARK_ARC_1_3/temp5[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_3  ( .A1(\RI5[3][44] ), .A2(n218), .Z(
        \MC_ARK_ARC_1_3/temp4[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_30_3  ( .A1(\RI5[3][146] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[170] ), .Z(\MC_ARK_ARC_1_3/temp2[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_30_3  ( .A1(\RI5[3][8] ), .A2(\RI5[3][2] ), .Z(
        \MC_ARK_ARC_1_3/temp1[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_30_2  ( .A1(\MC_ARK_ARC_1_3/temp6[9] ), .A2(
        \MC_ARK_ARC_1_3/temp5[9] ), .Z(\MC_ARK_ARC_1_3/buf_output[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_30_2  ( .A1(\MC_ARK_ARC_1_3/temp3[9] ), .A2(
        \MC_ARK_ARC_1_3/temp4[9] ), .Z(\MC_ARK_ARC_1_3/temp6[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_2  ( .A1(\RI5[3][45] ), .A2(n419), .Z(
        \MC_ARK_ARC_1_3/temp4[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_30_2  ( .A1(\RI5[3][75] ), .A2(\RI5[3][111] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[46] ), 
        .A2(n495), .Z(\MC_ARK_ARC_1_3/temp4[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_30_1  ( .A1(\RI5[3][172] ), .A2(\RI5[3][148] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_30_1  ( .A1(\RI5[3][10] ), .A2(\RI5[3][4] ), .Z(
        \MC_ARK_ARC_1_3/temp1[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_30_0  ( .A1(\MC_ARK_ARC_1_3/temp3[11] ), .A2(
        \MC_ARK_ARC_1_3/temp4[11] ), .Z(\MC_ARK_ARC_1_3/temp6[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_0  ( .A1(\RI5[3][47] ), .A2(n417), .Z(
        \MC_ARK_ARC_1_3/temp4[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_29_5  ( .A1(\MC_ARK_ARC_1_3/temp1[12] ), .A2(
        \MC_ARK_ARC_1_3/temp2[12] ), .Z(\MC_ARK_ARC_1_3/temp5[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_5  ( .A1(\RI5[3][48] ), .A2(n494), .Z(
        \MC_ARK_ARC_1_3/temp4[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_29_5  ( .A1(\RI5[3][174] ), .A2(\RI5[3][150] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), 
        .A2(n415), .Z(\MC_ARK_ARC_1_3/temp4[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_29_4  ( .A1(\RI5[3][175] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[151] ), .Z(\MC_ARK_ARC_1_3/temp2[13] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_3  ( .A1(\RI5[3][50] ), .A2(n492), .Z(
        \MC_ARK_ARC_1_3/temp4[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_29_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[176] ), 
        .A2(\RI5[3][152] ), .Z(\MC_ARK_ARC_1_3/temp2[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_29_3  ( .A1(\RI5[3][8] ), .A2(\RI5[3][14] ), .Z(
        \MC_ARK_ARC_1_3/temp1[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_29_1  ( .A1(\MC_ARK_ARC_1_3/temp1[16] ), .A2(
        \MC_ARK_ARC_1_3/temp2[16] ), .Z(\MC_ARK_ARC_1_3/temp5[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_1  ( .A1(\RI5[3][52] ), .A2(n156), .Z(
        \MC_ARK_ARC_1_3/temp4[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_29_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[118] ), 
        .A2(\RI5[3][82] ), .Z(\MC_ARK_ARC_1_3/temp3[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_29_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .A2(\RI5[3][154] ), .Z(\MC_ARK_ARC_1_3/temp2[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_29_1  ( .A1(\RI5[3][10] ), .A2(\RI5[3][16] ), .Z(
        \MC_ARK_ARC_1_3/temp1[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .A2(n568), .Z(\MC_ARK_ARC_1_3/temp4[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_29_0  ( .A1(\RI5[3][179] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[155] ), .Z(\MC_ARK_ARC_1_3/temp2[17] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_5  ( .A1(\RI5[3][54] ), .A2(n490), .Z(
        \MC_ARK_ARC_1_3/temp4[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_4  ( .A1(\RI5[3][55] ), .A2(n169), .Z(
        \MC_ARK_ARC_1_3/temp4[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_3  ( .A1(\RI5[3][56] ), .A2(n213), .Z(
        \MC_ARK_ARC_1_3/temp4[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_2  ( .A1(\RI5[3][57] ), .A2(n564), .Z(
        \MC_ARK_ARC_1_3/temp4[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_28_2  ( .A1(n575), .A2(\RI5[3][87] ), .Z(
        \MC_ARK_ARC_1_3/temp3[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_28_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[15] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[21] ), .Z(\MC_ARK_ARC_1_3/temp1[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_28_1  ( .A1(\MC_ARK_ARC_1_3/temp3[22] ), .A2(
        \MC_ARK_ARC_1_3/temp4[22] ), .Z(\MC_ARK_ARC_1_3/temp6[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_1  ( .A1(\RI5[3][58] ), .A2(n54), .Z(
        \MC_ARK_ARC_1_3/temp4[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_28_1  ( .A1(\RI5[3][124] ), .A2(\RI5[3][88] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_5  ( .A1(\SB2_3_26/buf_output[0] ), .A2(n175), 
        .Z(\MC_ARK_ARC_1_3/temp4[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_27_5  ( .A1(\SB2_3_0/buf_output[0] ), .A2(
        \RI5[3][18] ), .Z(\MC_ARK_ARC_1_3/temp1[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_27_4  ( .A1(\MC_ARK_ARC_1_3/temp3[25] ), .A2(
        \MC_ARK_ARC_1_3/temp4[25] ), .Z(\MC_ARK_ARC_1_3/temp6[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_4  ( .A1(\RI5[3][61] ), .A2(n561), .Z(
        \MC_ARK_ARC_1_3/temp4[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_27_4  ( .A1(\RI5[3][91] ), .A2(\RI5[3][127] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[62] ), 
        .A2(n191), .Z(\MC_ARK_ARC_1_3/temp4[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_2  ( .A1(\RI5[3][63] ), .A2(n559), .Z(
        \MC_ARK_ARC_1_3/temp4[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_27_2  ( .A1(\RI5[3][93] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[129] ), .Z(\MC_ARK_ARC_1_3/temp3[27] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_1  ( .A1(\SB2_3_22/buf_output[4] ), .A2(n52), 
        .Z(\MC_ARK_ARC_1_3/temp4[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_27_1  ( .A1(\RI5[3][130] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[94] ), .Z(\MC_ARK_ARC_1_3/temp3[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_27_1  ( .A1(\RI5[3][28] ), .A2(\RI5[3][22] ), .Z(
        \MC_ARK_ARC_1_3/temp1[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_0  ( .A1(\RI5[3][65] ), .A2(n557), .Z(
        \MC_ARK_ARC_1_3/temp4[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_26_5  ( .A1(\MC_ARK_ARC_1_3/temp3[30] ), .A2(
        \MC_ARK_ARC_1_3/temp4[30] ), .Z(\MC_ARK_ARC_1_3/temp6[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_26_5  ( .A1(\MC_ARK_ARC_1_3/temp1[30] ), .A2(
        \MC_ARK_ARC_1_3/temp2[30] ), .Z(\MC_ARK_ARC_1_3/temp5[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_5  ( .A1(\RI5[3][66] ), .A2(n482), .Z(
        \MC_ARK_ARC_1_3/temp4[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_26_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[96] ), 
        .A2(\RI5[3][132] ), .Z(\MC_ARK_ARC_1_3/temp3[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_26_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[0] ), 
        .A2(\RI5[3][168] ), .Z(\MC_ARK_ARC_1_3/temp2[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_4  ( .A1(\SB2_3_24/buf_output[1] ), .A2(n204), 
        .Z(\MC_ARK_ARC_1_3/temp4[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_4  ( .A1(\RI5[3][25] ), .A2(\RI5[3][31] ), .Z(
        \MC_ARK_ARC_1_3/temp1[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_3  ( .A1(\RI5[3][68] ), .A2(n480), .Z(
        \MC_ARK_ARC_1_3/temp4[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_26_3  ( .A1(\RI5[3][2] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[170] ), .Z(\MC_ARK_ARC_1_3/temp2[32] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_3  ( .A1(\RI5[3][26] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[32] ), .Z(\MC_ARK_ARC_1_3/temp1[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[69] ), 
        .A2(n92), .Z(\MC_ARK_ARC_1_3/temp4[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_26_2  ( .A1(\RI5[3][171] ), .A2(\RI5[3][3] ), .Z(
        \MC_ARK_ARC_1_3/temp2[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_26_1  ( .A1(\MC_ARK_ARC_1_3/temp5[34] ), .A2(
        \MC_ARK_ARC_1_3/temp6[34] ), .Z(\MC_ARK_ARC_1_3/buf_output[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_26_1  ( .A1(\MC_ARK_ARC_1_3/temp3[34] ), .A2(
        \MC_ARK_ARC_1_3/temp4[34] ), .Z(\MC_ARK_ARC_1_3/temp6[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_26_1  ( .A1(\MC_ARK_ARC_1_3/temp1[34] ), .A2(
        \MC_ARK_ARC_1_3/temp2[34] ), .Z(\MC_ARK_ARC_1_3/temp5[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_1  ( .A1(\RI5[3][70] ), .A2(n478), .Z(
        \MC_ARK_ARC_1_3/temp4[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_26_1  ( .A1(\RI5[3][136] ), .A2(\RI5[3][100] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_26_1  ( .A1(\RI5[3][4] ), .A2(\RI5[3][172] ), .Z(
        \MC_ARK_ARC_1_3/temp2[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_1  ( .A1(\RI5[3][34] ), .A2(\RI5[3][28] ), .Z(
        \MC_ARK_ARC_1_3/temp1[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[29] ), 
        .A2(\RI5[3][35] ), .Z(\MC_ARK_ARC_1_3/temp1[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_5  ( .A1(\RI5[3][72] ), .A2(n205), .Z(
        \MC_ARK_ARC_1_3/temp4[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_4  ( .A1(\RI5[3][73] ), .A2(n551), .Z(
        \MC_ARK_ARC_1_3/temp4[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_25_4  ( .A1(\SB2_3_12/buf_output[1] ), .A2(
        \RI5[3][103] ), .Z(\MC_ARK_ARC_1_3/temp3[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_25_3  ( .A1(\RI5[3][8] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[176] ), .Z(\MC_ARK_ARC_1_3/temp2[38] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_2  ( .A1(\SB2_3_21/buf_output[3] ), .A2(n550), 
        .Z(\MC_ARK_ARC_1_3/temp4[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_25_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[141] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[105] ), .Z(
        \MC_ARK_ARC_1_3/temp3[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_25_1  ( .A1(\MC_ARK_ARC_1_3/temp5[40] ), .A2(
        \MC_ARK_ARC_1_3/temp6[40] ), .Z(\MC_ARK_ARC_1_3/buf_output[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_25_1  ( .A1(\MC_ARK_ARC_1_3/temp3[40] ), .A2(
        \MC_ARK_ARC_1_3/temp4[40] ), .Z(\MC_ARK_ARC_1_3/temp6[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_1  ( .A1(\RI5[3][76] ), .A2(n472), .Z(
        \MC_ARK_ARC_1_3/temp4[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_25_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .A2(\RI5[3][106] ), .Z(\MC_ARK_ARC_1_3/temp3[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_25_1  ( .A1(\RI5[3][10] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[178] ), .Z(\MC_ARK_ARC_1_3/temp2[40] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_25_1  ( .A1(\RI5[3][40] ), .A2(\RI5[3][34] ), .Z(
        \MC_ARK_ARC_1_3/temp1[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_0  ( .A1(\RI5[3][77] ), .A2(n548), .Z(
        \MC_ARK_ARC_1_3/temp4[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_5  ( .A1(\RI5[3][78] ), .A2(n470), .Z(
        \MC_ARK_ARC_1_3/temp4[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_24_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[144] ), 
        .A2(\RI5[3][108] ), .Z(\MC_ARK_ARC_1_3/temp3[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_4  ( .A1(\SB2_3_22/buf_output[1] ), .A2(n546), 
        .Z(\MC_ARK_ARC_1_3/temp4[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_24_4  ( .A1(\RI5[3][181] ), .A2(\RI5[3][13] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[80] ), 
        .A2(n12), .Z(\MC_ARK_ARC_1_3/temp4[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_2  ( .A1(\RI5[3][81] ), .A2(n545), .Z(
        \MC_ARK_ARC_1_3/temp4[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_24_1  ( .A1(\MC_ARK_ARC_1_3/temp3[46] ), .A2(
        \MC_ARK_ARC_1_3/temp4[46] ), .Z(\MC_ARK_ARC_1_3/temp6[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_24_1  ( .A1(\MC_ARK_ARC_1_3/temp1[46] ), .A2(
        \MC_ARK_ARC_1_3/temp2[46] ), .Z(\MC_ARK_ARC_1_3/temp5[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_1  ( .A1(\RI5[3][82] ), .A2(n139), .Z(
        \MC_ARK_ARC_1_3/temp4[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_24_1  ( .A1(\RI5[3][148] ), .A2(\RI5[3][112] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_24_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[46] ), 
        .A2(\RI5[3][40] ), .Z(\MC_ARK_ARC_1_3/temp1[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_23_5  ( .A1(\MC_ARK_ARC_1_3/temp5[48] ), .A2(
        \MC_ARK_ARC_1_3/temp6[48] ), .Z(\MC_ARK_ARC_1_3/buf_output[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_23_5  ( .A1(\MC_ARK_ARC_1_3/temp4[48] ), .A2(
        \MC_ARK_ARC_1_3/temp3[48] ), .Z(\MC_ARK_ARC_1_3/temp6[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_23_5  ( .A1(\MC_ARK_ARC_1_3/temp1[48] ), .A2(
        \MC_ARK_ARC_1_3/temp2[48] ), .Z(\MC_ARK_ARC_1_3/temp5[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_5  ( .A1(\RI5[3][84] ), .A2(n465), .Z(
        \MC_ARK_ARC_1_3/temp4[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_23_5  ( .A1(\RI5[3][150] ), .A2(\RI5[3][114] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_23_5  ( .A1(\RI5[3][186] ), .A2(\RI5[3][18] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_23_5  ( .A1(\RI5[3][42] ), .A2(\RI5[3][48] ), .Z(
        \MC_ARK_ARC_1_3/temp1[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_23_4  ( .A1(\MC_ARK_ARC_1_3/temp4[49] ), .A2(
        \MC_ARK_ARC_1_3/temp3[49] ), .Z(\MC_ARK_ARC_1_3/temp6[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_23_4  ( .A1(\MC_ARK_ARC_1_3/temp1[49] ), .A2(
        \MC_ARK_ARC_1_3/temp2[49] ), .Z(\MC_ARK_ARC_1_3/temp5[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_4  ( .A1(\RI5[3][85] ), .A2(n201), .Z(
        \MC_ARK_ARC_1_3/temp4[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_23_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[151] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[115] ), .Z(
        \MC_ARK_ARC_1_3/temp3[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_23_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[19] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[187] ), .Z(
        \MC_ARK_ARC_1_3/temp2[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_23_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[43] ), .Z(\MC_ARK_ARC_1_3/temp1[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_23_3  ( .A1(\MC_ARK_ARC_1_3/temp5[50] ), .A2(
        \MC_ARK_ARC_1_3/temp6[50] ), .Z(\MC_ARK_ARC_1_3/buf_output[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_3  ( .A1(\RI5[3][86] ), .A2(n134), .Z(
        \MC_ARK_ARC_1_3/temp4[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_23_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[20] ), 
        .A2(n1506), .Z(\MC_ARK_ARC_1_3/temp2[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_2  ( .A1(\RI5[3][87] ), .A2(n123), .Z(
        \MC_ARK_ARC_1_3/temp4[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_23_2  ( .A1(\RI5[3][153] ), .A2(\RI5[3][117] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_23_1  ( .A1(\MC_ARK_ARC_1_3/temp4[52] ), .A2(
        \MC_ARK_ARC_1_3/temp3[52] ), .Z(\MC_ARK_ARC_1_3/temp6[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_1  ( .A1(\RI5[3][88] ), .A2(n55), .Z(
        \MC_ARK_ARC_1_3/temp4[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_23_1  ( .A1(\RI5[3][154] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[118] ), .Z(\MC_ARK_ARC_1_3/temp3[52] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_23_1  ( .A1(\RI5[3][22] ), .A2(\RI5[3][190] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_23_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[46] ), 
        .A2(\RI5[3][52] ), .Z(\MC_ARK_ARC_1_3/temp1[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_23_0  ( .A1(\MC_ARK_ARC_1_3/temp2[53] ), .A2(
        \MC_ARK_ARC_1_3/temp1[53] ), .Z(\MC_ARK_ARC_1_3/temp5[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_0  ( .A1(\RI5[3][89] ), .A2(n539), .Z(
        \MC_ARK_ARC_1_3/temp4[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_23_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), 
        .A2(\RI5[3][119] ), .Z(\MC_ARK_ARC_1_3/temp3[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_23_0  ( .A1(\RI5[3][191] ), .A2(\RI5[3][23] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_22_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[24] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[0] ), .Z(\MC_ARK_ARC_1_3/temp2[54] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_22_5  ( .A1(\RI5[3][48] ), .A2(\RI5[3][54] ), .Z(
        \MC_ARK_ARC_1_3/temp1[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_4  ( .A1(\RI5[3][91] ), .A2(n148), .Z(
        \MC_ARK_ARC_1_3/temp4[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_22_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[157] ), 
        .A2(\RI5[3][121] ), .Z(\MC_ARK_ARC_1_3/temp3[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_22_4  ( .A1(\RI5[3][25] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[1] ), .Z(\MC_ARK_ARC_1_3/temp2[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_22_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), 
        .A2(\RI5[3][55] ), .Z(\MC_ARK_ARC_1_3/temp1[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_22_3  ( .A1(\RI5[3][2] ), .A2(\RI5[3][26] ), .Z(
        \MC_ARK_ARC_1_3/temp2[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_2  ( .A1(\RI5[3][93] ), .A2(n77), .Z(
        \MC_ARK_ARC_1_3/temp4[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_22_2  ( .A1(n575), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[159] ), .Z(\MC_ARK_ARC_1_3/temp3[57] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_22_2  ( .A1(\RI5[3][27] ), .A2(\RI5[3][3] ), .Z(
        \MC_ARK_ARC_1_3/temp2[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[94] ), 
        .A2(n28), .Z(\MC_ARK_ARC_1_3/temp4[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_22_1  ( .A1(\RI5[3][160] ), .A2(\RI5[3][124] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_22_1  ( .A1(\RI5[3][28] ), .A2(\RI5[3][4] ), .Z(
        \MC_ARK_ARC_1_3/temp2[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_22_1  ( .A1(\RI5[3][58] ), .A2(\RI5[3][52] ), .Z(
        \MC_ARK_ARC_1_3/temp1[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_0  ( .A1(\RI5[3][95] ), .A2(n145), .Z(
        \MC_ARK_ARC_1_3/temp4[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[96] ), 
        .A2(n455), .Z(\MC_ARK_ARC_1_3/temp4[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_21_5  ( .A1(\RI5[3][162] ), .A2(\RI5[3][126] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_21_4  ( .A1(\MC_ARK_ARC_1_3/temp6[61] ), .A2(
        \MC_ARK_ARC_1_3/temp5[61] ), .Z(\MC_ARK_ARC_1_3/buf_output[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_4  ( .A1(\RI5[3][97] ), .A2(n534), .Z(
        \MC_ARK_ARC_1_3/temp4[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_21_4  ( .A1(\RI5[3][163] ), .A2(\RI5[3][127] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_21_4  ( .A1(\RI5[3][31] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[7] ), .Z(\MC_ARK_ARC_1_3/temp2[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_21_4  ( .A1(\RI5[3][55] ), .A2(\RI5[3][61] ), .Z(
        \MC_ARK_ARC_1_3/temp1[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_3  ( .A1(\RI5[3][98] ), .A2(n217), .Z(
        \MC_ARK_ARC_1_3/temp4[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_21_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[32] ), 
        .A2(\RI5[3][8] ), .Z(\MC_ARK_ARC_1_3/temp2[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_21_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[62] ), 
        .A2(\RI5[3][56] ), .Z(\MC_ARK_ARC_1_3/temp1[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[99] ), 
        .A2(n532), .Z(\MC_ARK_ARC_1_3/temp4[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_21_1  ( .A1(\MC_ARK_ARC_1_3/temp2[64] ), .A2(
        \MC_ARK_ARC_1_3/temp1[64] ), .Z(\MC_ARK_ARC_1_3/temp5[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_1  ( .A1(\RI5[3][100] ), .A2(n453), .Z(
        \MC_ARK_ARC_1_3/temp4[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_21_1  ( .A1(\RI5[3][166] ), .A2(\RI5[3][130] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_21_1  ( .A1(\RI5[3][10] ), .A2(\RI5[3][34] ), .Z(
        \MC_ARK_ARC_1_3/temp2[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_21_1  ( .A1(\RI5[3][64] ), .A2(\RI5[3][58] ), .Z(
        \MC_ARK_ARC_1_3/temp1[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_21_0  ( .A1(\MC_ARK_ARC_1_3/temp3[65] ), .A2(
        \MC_ARK_ARC_1_3/temp4[65] ), .Z(\MC_ARK_ARC_1_3/temp6[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_0  ( .A1(\RI5[3][101] ), .A2(n530), .Z(
        \MC_ARK_ARC_1_3/temp4[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_21_0  ( .A1(\RI5[3][11] ), .A2(\RI5[3][35] ), .Z(
        \MC_ARK_ARC_1_3/temp2[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_20_5  ( .A1(\MC_ARK_ARC_1_3/temp4[66] ), .A2(
        \MC_ARK_ARC_1_3/temp3[66] ), .Z(\MC_ARK_ARC_1_3/temp6[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_20_5  ( .A1(\MC_ARK_ARC_1_3/temp1[66] ), .A2(
        \MC_ARK_ARC_1_3/temp2[66] ), .Z(\MC_ARK_ARC_1_3/temp5[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[102] ), 
        .A2(n451), .Z(\MC_ARK_ARC_1_3/temp4[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_20_5  ( .A1(\RI5[3][168] ), .A2(\RI5[3][132] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_20_5  ( .A1(\RI5[3][36] ), .A2(\RI5[3][12] ), .Z(
        \MC_ARK_ARC_1_3/temp2[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_4  ( .A1(\RI5[3][103] ), .A2(n117), .Z(
        \MC_ARK_ARC_1_3/temp4[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_20_4  ( .A1(\RI5[3][169] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[133] ), .Z(\MC_ARK_ARC_1_3/temp3[67] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_20_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[37] ), 
        .A2(\RI5[3][13] ), .Z(\MC_ARK_ARC_1_3/temp2[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_20_4  ( .A1(\RI5[3][67] ), .A2(\RI5[3][61] ), .Z(
        \MC_ARK_ARC_1_3/temp1[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_20_3  ( .A1(\MC_ARK_ARC_1_3/temp5[68] ), .A2(
        \MC_ARK_ARC_1_3/temp6[68] ), .Z(\MC_ARK_ARC_1_3/buf_output[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_20_3  ( .A1(\MC_ARK_ARC_1_3/temp2[68] ), .A2(
        \MC_ARK_ARC_1_3/temp1[68] ), .Z(\MC_ARK_ARC_1_3/temp5[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_3  ( .A1(\RI5[3][104] ), .A2(n44), .Z(
        \MC_ARK_ARC_1_3/temp4[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_20_3  ( .A1(\RI5[3][38] ), .A2(\RI5[3][14] ), .Z(
        \MC_ARK_ARC_1_3/temp2[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_20_3  ( .A1(\RI5[3][68] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[62] ), .Z(\MC_ARK_ARC_1_3/temp1[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[105] ), 
        .A2(n526), .Z(\MC_ARK_ARC_1_3/temp4[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_20_1  ( .A1(\MC_ARK_ARC_1_3/temp6[70] ), .A2(
        \MC_ARK_ARC_1_3/temp5[70] ), .Z(\MC_ARK_ARC_1_3/buf_output[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_1  ( .A1(\RI5[3][106] ), .A2(n88), .Z(
        \MC_ARK_ARC_1_3/temp4[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_20_1  ( .A1(\RI5[3][40] ), .A2(\RI5[3][16] ), .Z(
        \MC_ARK_ARC_1_3/temp2[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_0  ( .A1(\RI5[3][107] ), .A2(n524), .Z(
        \MC_ARK_ARC_1_3/temp4[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_19_5  ( .A1(\MC_ARK_ARC_1_3/temp3[72] ), .A2(
        \MC_ARK_ARC_1_3/temp4[72] ), .Z(\MC_ARK_ARC_1_3/temp6[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_5  ( .A1(\RI5[3][108] ), .A2(n447), .Z(
        \MC_ARK_ARC_1_3/temp4[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_19_5  ( .A1(\RI5[3][42] ), .A2(\RI5[3][18] ), .Z(
        \MC_ARK_ARC_1_3/temp2[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_19_5  ( .A1(\RI5[3][72] ), .A2(\RI5[3][66] ), .Z(
        \MC_ARK_ARC_1_3/temp1[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_4  ( .A1(\SB2_3_17/buf_output[1] ), .A2(n522), 
        .Z(\MC_ARK_ARC_1_3/temp4[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_3  ( .A1(\RI5[3][110] ), .A2(n445), .Z(
        \MC_ARK_ARC_1_3/temp4[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_19_3  ( .A1(\RI5[3][74] ), .A2(\RI5[3][68] ), .Z(
        \MC_ARK_ARC_1_3/temp1[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_2  ( .A1(\RI5[3][111] ), .A2(n521), .Z(
        \MC_ARK_ARC_1_3/temp4[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_19_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[177] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[141] ), .Z(
        \MC_ARK_ARC_1_3/temp3[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_19_2  ( .A1(\RI5[3][75] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[69] ), .Z(\MC_ARK_ARC_1_3/temp1[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_1  ( .A1(\RI5[3][112] ), .A2(n443), .Z(
        \MC_ARK_ARC_1_3/temp4[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_19_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[178] ), .Z(
        \MC_ARK_ARC_1_3/temp3[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_0  ( .A1(\RI5[3][113] ), .A2(n48), .Z(
        \MC_ARK_ARC_1_3/temp4[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_19_0  ( .A1(\RI5[3][77] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[71] ), .Z(\MC_ARK_ARC_1_3/temp1[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_18_5  ( .A1(\MC_ARK_ARC_1_3/temp3[78] ), .A2(
        \MC_ARK_ARC_1_3/temp4[78] ), .Z(\MC_ARK_ARC_1_3/temp6[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_5  ( .A1(\RI5[3][114] ), .A2(n441), .Z(
        \MC_ARK_ARC_1_3/temp4[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_18_5  ( .A1(\RI5[3][78] ), .A2(\RI5[3][72] ), .Z(
        \MC_ARK_ARC_1_3/temp1[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[115] ), 
        .A2(n518), .Z(\MC_ARK_ARC_1_3/temp4[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_18_4  ( .A1(\RI5[3][181] ), .A2(\RI5[3][145] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), 
        .A2(n23), .Z(\MC_ARK_ARC_1_3/temp4[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_18_3  ( .A1(\RI5[3][146] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[182] ), .Z(\MC_ARK_ARC_1_3/temp3[80] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_18_1  ( .A1(\MC_ARK_ARC_1_3/temp5[82] ), .A2(
        \MC_ARK_ARC_1_3/temp6[82] ), .Z(\MC_ARK_ARC_1_3/buf_output[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_18_1  ( .A1(\MC_ARK_ARC_1_3/temp4[82] ), .A2(
        \MC_ARK_ARC_1_3/temp3[82] ), .Z(\MC_ARK_ARC_1_3/temp6[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_18_1  ( .A1(\MC_ARK_ARC_1_3/temp2[82] ), .A2(
        \MC_ARK_ARC_1_3/temp1[82] ), .Z(\MC_ARK_ARC_1_3/temp5[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[118] ), 
        .A2(n43), .Z(\MC_ARK_ARC_1_3/temp4[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_18_1  ( .A1(\RI5[3][148] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[184] ), .Z(\MC_ARK_ARC_1_3/temp3[82] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_18_1  ( .A1(\RI5[3][82] ), .A2(\RI5[3][76] ), .Z(
        \MC_ARK_ARC_1_3/temp1[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_18_0  ( .A1(\MC_ARK_ARC_1_3/temp1[83] ), .A2(
        \MC_ARK_ARC_1_3/temp2[83] ), .Z(\MC_ARK_ARC_1_3/temp5[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_18_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[29] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[53] ), .Z(\MC_ARK_ARC_1_3/temp2[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_18_0  ( .A1(\RI5[3][83] ), .A2(\RI5[3][77] ), .Z(
        \MC_ARK_ARC_1_3/temp1[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_17_5  ( .A1(\MC_ARK_ARC_1_3/temp3[84] ), .A2(
        \MC_ARK_ARC_1_3/temp4[84] ), .Z(\MC_ARK_ARC_1_3/temp6[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_17_5  ( .A1(\MC_ARK_ARC_1_3/temp1[84] ), .A2(
        \MC_ARK_ARC_1_3/temp2[84] ), .Z(\MC_ARK_ARC_1_3/temp5[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_5  ( .A1(\RI5[3][120] ), .A2(n436), .Z(
        \MC_ARK_ARC_1_3/temp4[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_17_5  ( .A1(\RI5[3][186] ), .A2(\RI5[3][150] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_17_5  ( .A1(\RI5[3][30] ), .A2(\RI5[3][54] ), .Z(
        \MC_ARK_ARC_1_3/temp2[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_17_4  ( .A1(\MC_ARK_ARC_1_3/temp3[85] ), .A2(
        \MC_ARK_ARC_1_3/temp4[85] ), .Z(\MC_ARK_ARC_1_3/temp6[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_4  ( .A1(\RI5[3][121] ), .A2(n151), .Z(
        \MC_ARK_ARC_1_3/temp4[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_17_4  ( .A1(\RI5[3][85] ), .A2(\RI5[3][79] ), .Z(
        \MC_ARK_ARC_1_3/temp1[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_3  ( .A1(\RI5[3][122] ), .A2(n34), .Z(
        \MC_ARK_ARC_1_3/temp4[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_17_3  ( .A1(n1506), .A2(\RI5[3][152] ), .Z(
        \MC_ARK_ARC_1_3/temp3[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_2  ( .A1(n575), .A2(n150), .Z(
        \MC_ARK_ARC_1_3/temp4[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_17_2  ( .A1(\RI5[3][189] ), .A2(\RI5[3][153] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_17_2  ( .A1(\RI5[3][33] ), .A2(\RI5[3][57] ), .Z(
        \MC_ARK_ARC_1_3/temp2[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_17_2  ( .A1(\RI5[3][81] ), .A2(\RI5[3][87] ), .Z(
        \MC_ARK_ARC_1_3/temp1[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_17_1  ( .A1(\MC_ARK_ARC_1_3/temp4[88] ), .A2(
        \MC_ARK_ARC_1_3/temp3[88] ), .Z(\MC_ARK_ARC_1_3/temp6[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_17_1  ( .A1(\MC_ARK_ARC_1_3/temp1[88] ), .A2(
        \MC_ARK_ARC_1_3/temp2[88] ), .Z(\MC_ARK_ARC_1_3/temp5[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_1  ( .A1(\RI5[3][124] ), .A2(n119), .Z(
        \MC_ARK_ARC_1_3/temp4[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_17_1  ( .A1(\RI5[3][190] ), .A2(\RI5[3][154] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_17_1  ( .A1(\RI5[3][58] ), .A2(\RI5[3][34] ), .Z(
        \MC_ARK_ARC_1_3/temp2[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_17_1  ( .A1(\RI5[3][88] ), .A2(\RI5[3][82] ), .Z(
        \MC_ARK_ARC_1_3/temp1[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_0  ( .A1(\RI5[3][125] ), .A2(n68), .Z(
        \MC_ARK_ARC_1_3/temp4[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_17_0  ( .A1(\RI5[3][83] ), .A2(\RI5[3][89] ), .Z(
        \MC_ARK_ARC_1_3/temp1[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_5  ( .A1(\RI5[3][126] ), .A2(n136), .Z(
        \MC_ARK_ARC_1_3/temp4[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_16_5  ( .A1(\RI5[3][60] ), .A2(\RI5[3][36] ), .Z(
        \MC_ARK_ARC_1_3/temp2[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_16_5  ( .A1(\RI5[3][84] ), .A2(\RI5[3][90] ), .Z(
        \MC_ARK_ARC_1_3/temp1[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_4  ( .A1(\RI5[3][127] ), .A2(n141), .Z(
        \MC_ARK_ARC_1_3/temp4[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_16_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[1] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[157] ), .Z(
        \MC_ARK_ARC_1_3/temp3[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[128] ), 
        .A2(n20), .Z(\MC_ARK_ARC_1_3/temp4[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_16_3  ( .A1(\RI5[3][92] ), .A2(\RI5[3][86] ), .Z(
        \MC_ARK_ARC_1_3/temp1[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[129] ), 
        .A2(n80), .Z(\MC_ARK_ARC_1_3/temp4[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_16_1  ( .A1(\MC_ARK_ARC_1_3/temp4[94] ), .A2(
        \MC_ARK_ARC_1_3/temp3[94] ), .Z(\MC_ARK_ARC_1_3/temp6[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_1  ( .A1(\RI5[3][130] ), .A2(n427), .Z(
        \MC_ARK_ARC_1_3/temp4[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_16_1  ( .A1(\RI5[3][40] ), .A2(\RI5[3][64] ), .Z(
        \MC_ARK_ARC_1_3/temp2[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_0  ( .A1(\RI5[3][131] ), .A2(n504), .Z(
        \MC_ARK_ARC_1_3/temp4[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_15_5  ( .A1(\MC_ARK_ARC_1_3/temp5[96] ), .A2(
        \MC_ARK_ARC_1_3/temp6[96] ), .Z(\MC_ARK_ARC_1_3/buf_output[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_15_5  ( .A1(\MC_ARK_ARC_1_3/temp3[96] ), .A2(
        \MC_ARK_ARC_1_3/temp4[96] ), .Z(\MC_ARK_ARC_1_3/temp6[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_5  ( .A1(\RI5[3][132] ), .A2(n425), .Z(
        \MC_ARK_ARC_1_3/temp4[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_15_5  ( .A1(\RI5[3][6] ), .A2(\RI5[3][162] ), .Z(
        \MC_ARK_ARC_1_3/temp3[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_15_5  ( .A1(\RI5[3][42] ), .A2(\RI5[3][66] ), .Z(
        \MC_ARK_ARC_1_3/temp2[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_15_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[96] ), 
        .A2(\RI5[3][90] ), .Z(\MC_ARK_ARC_1_3/temp1[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_15_4  ( .A1(\MC_ARK_ARC_1_3/temp4[97] ), .A2(
        \MC_ARK_ARC_1_3/temp3[97] ), .Z(\MC_ARK_ARC_1_3/temp6[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[133] ), 
        .A2(n503), .Z(\MC_ARK_ARC_1_3/temp4[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_15_4  ( .A1(\RI5[3][163] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[7] ), .Z(\MC_ARK_ARC_1_3/temp3[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_3  ( .A1(\RI5[3][134] ), .A2(n124), .Z(
        \MC_ARK_ARC_1_3/temp4[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_15_3  ( .A1(\RI5[3][68] ), .A2(\RI5[3][44] ), .Z(
        \MC_ARK_ARC_1_3/temp2[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_2  ( .A1(\RI5[3][135] ), .A2(n501), .Z(
        \MC_ARK_ARC_1_3/temp4[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_15_2  ( .A1(\RI5[3][45] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[69] ), .Z(\MC_ARK_ARC_1_3/temp2[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_1  ( .A1(\RI5[3][136] ), .A2(n422), .Z(
        \MC_ARK_ARC_1_3/temp4[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_15_0  ( .A1(\MC_ARK_ARC_1_3/temp3[101] ), .A2(
        \MC_ARK_ARC_1_3/temp4[101] ), .Z(\MC_ARK_ARC_1_3/temp6[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_0  ( .A1(\RI5[3][137] ), .A2(n116), .Z(
        \MC_ARK_ARC_1_3/temp4[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_15_0  ( .A1(\RI5[3][167] ), .A2(\RI5[3][11] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_15_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .A2(\RI5[3][47] ), .Z(\MC_ARK_ARC_1_3/temp2[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_15_0  ( .A1(\RI5[3][101] ), .A2(\RI5[3][95] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_14_5  ( .A1(\RI5[3][138] ), .A2(n420), .Z(
        \MC_ARK_ARC_1_3/temp4[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_14_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[102] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[96] ), .Z(
        \MC_ARK_ARC_1_3/temp1[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_14_4  ( .A1(\RI5[3][139] ), .A2(n497), .Z(
        \MC_ARK_ARC_1_3/temp4[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_14_4  ( .A1(\SB2_3_27/buf_output[1] ), .A2(
        \RI5[3][73] ), .Z(\MC_ARK_ARC_1_3/temp2[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_14_4  ( .A1(\SB2_3_19/buf_output[1] ), .A2(
        \RI5[3][103] ), .Z(\MC_ARK_ARC_1_3/temp1[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_14_2  ( .A1(\MC_ARK_ARC_1_3/temp3[105] ), .A2(
        \MC_ARK_ARC_1_3/temp4[105] ), .Z(\MC_ARK_ARC_1_3/temp6[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_14_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[141] ), 
        .A2(n496), .Z(\MC_ARK_ARC_1_3/temp4[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_14_2  ( .A1(\RI5[3][75] ), .A2(\RI5[3][51] ), .Z(
        \MC_ARK_ARC_1_3/temp2[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_14_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .A2(n2), .Z(\MC_ARK_ARC_1_3/temp4[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_14_1  ( .A1(\RI5[3][76] ), .A2(\RI5[3][52] ), .Z(
        \MC_ARK_ARC_1_3/temp2[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_14_1  ( .A1(\RI5[3][106] ), .A2(\RI5[3][100] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_14_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[143] ), 
        .A2(n192), .Z(\MC_ARK_ARC_1_3/temp4[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_13_5  ( .A1(\MC_ARK_ARC_1_3/temp3[108] ), .A2(
        \MC_ARK_ARC_1_3/temp4[108] ), .Z(\MC_ARK_ARC_1_3/temp6[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[144] ), 
        .A2(n416), .Z(\MC_ARK_ARC_1_3/temp4[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_13_5  ( .A1(\RI5[3][174] ), .A2(\RI5[3][18] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_13_5  ( .A1(\RI5[3][54] ), .A2(\RI5[3][78] ), .Z(
        \MC_ARK_ARC_1_3/temp2[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_4  ( .A1(\RI5[3][145] ), .A2(n493), .Z(
        \MC_ARK_ARC_1_3/temp4[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_13_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[19] ), 
        .A2(\RI5[3][175] ), .Z(\MC_ARK_ARC_1_3/temp3[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_13_4  ( .A1(\RI5[3][79] ), .A2(\RI5[3][55] ), .Z(
        \MC_ARK_ARC_1_3/temp2[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_13_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[109] ), 
        .A2(\RI5[3][103] ), .Z(\MC_ARK_ARC_1_3/temp1[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_3  ( .A1(\RI5[3][146] ), .A2(n414), .Z(
        \MC_ARK_ARC_1_3/temp4[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_13_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[20] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[176] ), .Z(
        \MC_ARK_ARC_1_3/temp3[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_13_2  ( .A1(\MC_ARK_ARC_1_3/temp5[111] ), .A2(
        \MC_ARK_ARC_1_3/temp6[111] ), .Z(\MC_ARK_ARC_1_3/buf_output[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_13_2  ( .A1(\MC_ARK_ARC_1_3/temp3[111] ), .A2(
        \MC_ARK_ARC_1_3/temp4[111] ), .Z(\MC_ARK_ARC_1_3/temp6[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_13_2  ( .A1(\MC_ARK_ARC_1_3/temp2[111] ), .A2(
        \MC_ARK_ARC_1_3/temp1[111] ), .Z(\MC_ARK_ARC_1_3/temp5[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[147] ), 
        .A2(n160), .Z(\MC_ARK_ARC_1_3/temp4[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_13_2  ( .A1(\RI5[3][57] ), .A2(\RI5[3][81] ), .Z(
        \MC_ARK_ARC_1_3/temp2[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_13_2  ( .A1(\RI5[3][111] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[105] ), .Z(\MC_ARK_ARC_1_3/temp1[111] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_13_1  ( .A1(\MC_ARK_ARC_1_3/temp5[112] ), .A2(
        \MC_ARK_ARC_1_3/temp6[112] ), .Z(\MC_ARK_ARC_1_3/buf_output[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_13_1  ( .A1(\MC_ARK_ARC_1_3/temp4[112] ), .A2(
        \MC_ARK_ARC_1_3/temp3[112] ), .Z(\MC_ARK_ARC_1_3/temp6[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_1  ( .A1(\RI5[3][148] ), .A2(n569), .Z(
        \MC_ARK_ARC_1_3/temp4[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_13_1  ( .A1(\RI5[3][22] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[178] ), .Z(\MC_ARK_ARC_1_3/temp3[112] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_13_1  ( .A1(\RI5[3][82] ), .A2(\RI5[3][58] ), .Z(
        \MC_ARK_ARC_1_3/temp2[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_13_0  ( .A1(\MC_ARK_ARC_1_3/temp3[113] ), .A2(
        \MC_ARK_ARC_1_3/temp4[113] ), .Z(\MC_ARK_ARC_1_3/temp6[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_0  ( .A1(\RI5[3][149] ), .A2(n168), .Z(
        \MC_ARK_ARC_1_3/temp4[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_13_0  ( .A1(\RI5[3][83] ), .A2(\RI5[3][59] ), .Z(
        \MC_ARK_ARC_1_3/temp2[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_13_0  ( .A1(\RI5[3][107] ), .A2(\RI5[3][113] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_4  ( .A1(\SB2_3_10/buf_output[1] ), .A2(n489), 
        .Z(\MC_ARK_ARC_1_3/temp4[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_12_4  ( .A1(\RI5[3][181] ), .A2(\RI5[3][25] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_12_3  ( .A1(\MC_ARK_ARC_1_3/temp3[116] ), .A2(
        \MC_ARK_ARC_1_3/temp4[116] ), .Z(\MC_ARK_ARC_1_3/temp6[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_3  ( .A1(\RI5[3][152] ), .A2(n565), .Z(
        \MC_ARK_ARC_1_3/temp4[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_12_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[62] ), 
        .A2(\RI5[3][86] ), .Z(\MC_ARK_ARC_1_3/temp2[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_12_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), 
        .A2(\RI5[3][110] ), .Z(\MC_ARK_ARC_1_3/temp1[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_2  ( .A1(\RI5[3][153] ), .A2(n89), .Z(
        \MC_ARK_ARC_1_3/temp4[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_12_2  ( .A1(\RI5[3][111] ), .A2(\RI5[3][117] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_1  ( .A1(\RI5[3][154] ), .A2(n563), .Z(
        \MC_ARK_ARC_1_3/temp4[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_12_1  ( .A1(\RI5[3][28] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[184] ), .Z(\MC_ARK_ARC_1_3/temp3[118] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_12_1  ( .A1(\RI5[3][112] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[118] ), .Z(\MC_ARK_ARC_1_3/temp1[118] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_11_5  ( .A1(\MC_ARK_ARC_1_3/temp6[120] ), .A2(
        \MC_ARK_ARC_1_3/temp5[120] ), .Z(\MC_ARK_ARC_1_3/buf_output[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[156] ), 
        .A2(n562), .Z(\MC_ARK_ARC_1_3/temp4[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_11_5  ( .A1(\RI5[3][186] ), .A2(\RI5[3][30] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_11_4  ( .A1(\MC_ARK_ARC_1_3/temp5[121] ), .A2(
        \MC_ARK_ARC_1_3/temp6[121] ), .Z(\MC_ARK_ARC_1_3/buf_output[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_11_4  ( .A1(\MC_ARK_ARC_1_3/temp3[121] ), .A2(
        \MC_ARK_ARC_1_3/temp4[121] ), .Z(\MC_ARK_ARC_1_3/temp6[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_11_4  ( .A1(\MC_ARK_ARC_1_3/temp2[121] ), .A2(
        \MC_ARK_ARC_1_3/temp1[121] ), .Z(\MC_ARK_ARC_1_3/temp5[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[157] ), 
        .A2(n486), .Z(\MC_ARK_ARC_1_3/temp4[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_11_4  ( .A1(\RI5[3][31] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[187] ), .Z(\MC_ARK_ARC_1_3/temp3[121] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_11_4  ( .A1(\RI5[3][121] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_3/temp1[121] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[158] ), 
        .A2(n560), .Z(\MC_ARK_ARC_1_3/temp4[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_11_3  ( .A1(\RI5[3][92] ), .A2(\RI5[3][68] ), .Z(
        \MC_ARK_ARC_1_3/temp2[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[159] ), 
        .A2(n485), .Z(\MC_ARK_ARC_1_3/temp4[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_11_2  ( .A1(\RI5[3][33] ), .A2(\RI5[3][189] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_11_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[69] ), 
        .A2(\RI5[3][93] ), .Z(\MC_ARK_ARC_1_3/temp2[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_11_2  ( .A1(\RI5[3][117] ), .A2(n575), .Z(
        \MC_ARK_ARC_1_3/temp1[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_1  ( .A1(\RI5[3][160] ), .A2(n95), .Z(
        \MC_ARK_ARC_1_3/temp4[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_11_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[94] ), 
        .A2(\RI5[3][70] ), .Z(\MC_ARK_ARC_1_3/temp2[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_11_1  ( .A1(\RI5[3][124] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[118] ), .Z(\MC_ARK_ARC_1_3/temp1[124] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_0  ( .A1(\RI5[3][161] ), .A2(n483), .Z(
        \MC_ARK_ARC_1_3/temp4[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_11_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .A2(\RI5[3][95] ), .Z(\MC_ARK_ARC_1_3/temp2[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_11_0  ( .A1(\RI5[3][119] ), .A2(\RI5[3][125] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_10_5  ( .A1(\MC_ARK_ARC_1_3/temp3[126] ), .A2(
        \MC_ARK_ARC_1_3/temp4[126] ), .Z(\MC_ARK_ARC_1_3/temp6[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_5  ( .A1(\RI5[3][162] ), .A2(n31), .Z(
        \MC_ARK_ARC_1_3/temp4[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_10_5  ( .A1(\RI5[3][36] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[0] ), .Z(\MC_ARK_ARC_1_3/temp3[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_10_5  ( .A1(\RI5[3][72] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[96] ), .Z(\MC_ARK_ARC_1_3/temp2[126] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_10_5  ( .A1(\RI5[3][126] ), .A2(\RI5[3][120] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_10_4  ( .A1(\MC_ARK_ARC_1_3/temp2[127] ), .A2(
        \MC_ARK_ARC_1_3/temp1[127] ), .Z(\MC_ARK_ARC_1_3/temp5[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_4  ( .A1(\RI5[3][163] ), .A2(
        \MC_ARK_ARC_1_1/buf_keyinput[119] ), .Z(\MC_ARK_ARC_1_3/temp4[127] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_10_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[37] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[1] ), .Z(\MC_ARK_ARC_1_3/temp3[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_10_4  ( .A1(\RI5[3][97] ), .A2(\RI5[3][73] ), .Z(
        \MC_ARK_ARC_1_3/temp2[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_10_4  ( .A1(\RI5[3][127] ), .A2(\RI5[3][121] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_10_3  ( .A1(\MC_ARK_ARC_1_3/temp3[128] ), .A2(
        \MC_ARK_ARC_1_3/temp4[128] ), .Z(\MC_ARK_ARC_1_3/temp6[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_10_3  ( .A1(\MC_ARK_ARC_1_3/temp2[128] ), .A2(
        \MC_ARK_ARC_1_3/temp1[128] ), .Z(\MC_ARK_ARC_1_3/temp5[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[164] ), 
        .A2(n126), .Z(\MC_ARK_ARC_1_3/temp4[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_10_3  ( .A1(\RI5[3][74] ), .A2(\RI5[3][98] ), .Z(
        \MC_ARK_ARC_1_3/temp2[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_10_3  ( .A1(\RI5[3][122] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[128] ), .Z(\MC_ARK_ARC_1_3/temp1[128] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_2  ( .A1(\RI5[3][165] ), .A2(n176), .Z(
        \MC_ARK_ARC_1_3/temp4[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_10_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[39] ), 
        .A2(\RI5[3][3] ), .Z(\MC_ARK_ARC_1_3/temp3[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_10_1  ( .A1(\MC_ARK_ARC_1_3/temp3[130] ), .A2(
        \MC_ARK_ARC_1_3/temp4[130] ), .Z(\MC_ARK_ARC_1_3/temp6[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_1  ( .A1(\RI5[3][166] ), .A2(n553), .Z(
        \MC_ARK_ARC_1_3/temp4[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_10_1  ( .A1(\RI5[3][40] ), .A2(\RI5[3][4] ), .Z(
        \MC_ARK_ARC_1_3/temp3[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_10_1  ( .A1(\RI5[3][100] ), .A2(\RI5[3][76] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_10_1  ( .A1(\RI5[3][130] ), .A2(\RI5[3][124] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_0  ( .A1(\SB2_3_4/buf_output[5] ), .A2(n477), 
        .Z(\MC_ARK_ARC_1_3/temp4[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_5  ( .A1(\RI5[3][168] ), .A2(
        \MC_ARK_ARC_1_3/buf_keyinput[132] ), .Z(\MC_ARK_ARC_1_3/temp4[132] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_9_5  ( .A1(\RI5[3][78] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[102] ), .Z(\MC_ARK_ARC_1_3/temp2[132] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_4  ( .A1(\RI5[3][169] ), .A2(n475), .Z(
        \MC_ARK_ARC_1_3/temp4[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_9_4  ( .A1(\RI5[3][79] ), .A2(\RI5[3][103] ), .Z(
        \MC_ARK_ARC_1_3/temp2[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[133] ), 
        .A2(\RI5[3][127] ), .Z(\MC_ARK_ARC_1_3/temp1[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[170] ), 
        .A2(n188), .Z(\MC_ARK_ARC_1_3/temp4[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_3  ( .A1(\RI5[3][134] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[128] ), .Z(\MC_ARK_ARC_1_3/temp1[134] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_2  ( .A1(\RI5[3][171] ), .A2(n473), .Z(
        \MC_ARK_ARC_1_3/temp4[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_9_2  ( .A1(\RI5[3][81] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[105] ), .Z(\MC_ARK_ARC_1_3/temp2[135] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_2  ( .A1(\RI5[3][135] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[129] ), .Z(\MC_ARK_ARC_1_3/temp1[135] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_1  ( .A1(\RI5[3][172] ), .A2(n549), .Z(
        \MC_ARK_ARC_1_3/temp4[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_9_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[46] ), 
        .A2(\RI5[3][10] ), .Z(\MC_ARK_ARC_1_3/temp3[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_1  ( .A1(\RI5[3][136] ), .A2(\RI5[3][130] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_8_5  ( .A1(\MC_ARK_ARC_1_3/temp4[138] ), .A2(
        \MC_ARK_ARC_1_3/temp3[138] ), .Z(\MC_ARK_ARC_1_3/temp6[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_5  ( .A1(\RI5[3][174] ), .A2(n547), .Z(
        \MC_ARK_ARC_1_3/temp4[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_8_5  ( .A1(\RI5[3][48] ), .A2(\RI5[3][12] ), .Z(
        \MC_ARK_ARC_1_3/temp3[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_8_4  ( .A1(\MC_ARK_ARC_1_3/temp5[139] ), .A2(
        \MC_ARK_ARC_1_3/temp6[139] ), .Z(\MC_ARK_ARC_1_3/buf_output[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_8_4  ( .A1(\MC_ARK_ARC_1_3/temp3[139] ), .A2(
        \MC_ARK_ARC_1_3/temp4[139] ), .Z(\MC_ARK_ARC_1_3/temp6[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_8_4  ( .A1(\MC_ARK_ARC_1_3/temp2[139] ), .A2(
        \MC_ARK_ARC_1_3/temp1[139] ), .Z(\MC_ARK_ARC_1_3/temp5[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_4  ( .A1(\RI5[3][175] ), .A2(n161), .Z(
        \MC_ARK_ARC_1_3/temp4[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_8_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), 
        .A2(\RI5[3][13] ), .Z(\MC_ARK_ARC_1_3/temp3[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_8_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[109] ), 
        .A2(\RI5[3][85] ), .Z(\MC_ARK_ARC_1_3/temp2[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_8_4  ( .A1(\RI5[3][139] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[133] ), .Z(\MC_ARK_ARC_1_3/temp1[139] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_8_3  ( .A1(\MC_ARK_ARC_1_3/temp1[140] ), .A2(
        \MC_ARK_ARC_1_3/temp2[140] ), .Z(\MC_ARK_ARC_1_3/temp5[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[176] ), 
        .A2(n158), .Z(\MC_ARK_ARC_1_3/temp4[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_8_3  ( .A1(\RI5[3][50] ), .A2(\RI5[3][14] ), .Z(
        \MC_ARK_ARC_1_3/temp3[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[177] ), 
        .A2(n467), .Z(\MC_ARK_ARC_1_3/temp4[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_8_1  ( .A1(\MC_ARK_ARC_1_3/temp5[142] ), .A2(
        \MC_ARK_ARC_1_3/temp6[142] ), .Z(\MC_ARK_ARC_1_3/buf_output[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_8_1  ( .A1(\MC_ARK_ARC_1_3/temp4[142] ), .A2(
        \MC_ARK_ARC_1_3/temp3[142] ), .Z(\MC_ARK_ARC_1_3/temp6[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_8_1  ( .A1(\MC_ARK_ARC_1_3/temp1[142] ), .A2(
        \MC_ARK_ARC_1_3/temp2[142] ), .Z(\MC_ARK_ARC_1_3/temp5[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .A2(n30), .Z(\MC_ARK_ARC_1_3/temp4[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_8_1  ( .A1(\RI5[3][52] ), .A2(\RI5[3][16] ), .Z(
        \MC_ARK_ARC_1_3/temp3[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_8_1  ( .A1(\RI5[3][112] ), .A2(\RI5[3][88] ), .Z(
        \MC_ARK_ARC_1_3/temp2[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_8_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .A2(\RI5[3][136] ), .Z(\MC_ARK_ARC_1_3/temp1[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_0  ( .A1(\RI5[3][179] ), .A2(n466), .Z(
        \MC_ARK_ARC_1_3/temp4[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_8_0  ( .A1(\RI5[3][17] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[53] ), .Z(\MC_ARK_ARC_1_3/temp3[143] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_7_5  ( .A1(\MC_ARK_ARC_1_3/temp5[144] ), .A2(
        \MC_ARK_ARC_1_3/temp6[144] ), .Z(\MC_ARK_ARC_1_3/buf_output[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_7_5  ( .A1(\MC_ARK_ARC_1_3/temp3[144] ), .A2(
        \MC_ARK_ARC_1_3/temp4[144] ), .Z(\MC_ARK_ARC_1_3/temp6[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_5  ( .A1(\RI5[3][180] ), .A2(n542), .Z(
        \MC_ARK_ARC_1_3/temp4[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_7_5  ( .A1(\RI5[3][54] ), .A2(\RI5[3][18] ), .Z(
        \MC_ARK_ARC_1_3/temp3[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_7_5  ( .A1(\RI5[3][90] ), .A2(\RI5[3][114] ), .Z(
        \MC_ARK_ARC_1_3/temp2[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_7_5  ( .A1(\RI5[3][138] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[144] ), .Z(\MC_ARK_ARC_1_3/temp1[144] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_7_4  ( .A1(\MC_ARK_ARC_1_3/temp3[145] ), .A2(
        \MC_ARK_ARC_1_3/temp4[145] ), .Z(\MC_ARK_ARC_1_3/temp6[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_4  ( .A1(\RI5[3][181] ), .A2(n464), .Z(
        \MC_ARK_ARC_1_3/temp4[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_7_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[19] ), 
        .A2(\RI5[3][55] ), .Z(\MC_ARK_ARC_1_3/temp3[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_7_4  ( .A1(\RI5[3][139] ), .A2(\RI5[3][145] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_7_3  ( .A1(\MC_ARK_ARC_1_3/temp5[146] ), .A2(
        \MC_ARK_ARC_1_3/temp6[146] ), .Z(\MC_ARK_ARC_1_3/buf_output[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_7_3  ( .A1(\MC_ARK_ARC_1_3/temp3[146] ), .A2(
        \MC_ARK_ARC_1_3/temp4[146] ), .Z(\MC_ARK_ARC_1_3/temp6[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[182] ), 
        .A2(n541), .Z(\MC_ARK_ARC_1_3/temp4[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[183] ), 
        .A2(n463), .Z(\MC_ARK_ARC_1_3/temp4[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_7_2  ( .A1(\RI5[3][57] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[21] ), .Z(\MC_ARK_ARC_1_3/temp3[147] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_7_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[94] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[118] ), .Z(
        \MC_ARK_ARC_1_3/temp2[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_7_0  ( .A1(\MC_ARK_ARC_1_3/temp3[149] ), .A2(
        \MC_ARK_ARC_1_3/temp4[149] ), .Z(\MC_ARK_ARC_1_3/temp6[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_0  ( .A1(\RI5[3][185] ), .A2(n32), .Z(
        \MC_ARK_ARC_1_3/temp4[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_7_0  ( .A1(\RI5[3][23] ), .A2(\RI5[3][59] ), .Z(
        \MC_ARK_ARC_1_3/temp3[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_7_0  ( .A1(\RI5[3][119] ), .A2(\RI5[3][95] ), .Z(
        \MC_ARK_ARC_1_3/temp2[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_5  ( .A1(\RI5[3][186] ), .A2(n538), .Z(
        \MC_ARK_ARC_1_3/temp4[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_6_4  ( .A1(\MC_ARK_ARC_1_3/temp3[151] ), .A2(
        \MC_ARK_ARC_1_3/temp4[151] ), .Z(\MC_ARK_ARC_1_3/temp6[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[187] ), 
        .A2(n459), .Z(\MC_ARK_ARC_1_3/temp4[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_6_4  ( .A1(\RI5[3][61] ), .A2(\RI5[3][25] ), .Z(
        \MC_ARK_ARC_1_3/temp3[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_6_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[151] ), 
        .A2(\RI5[3][145] ), .Z(\MC_ARK_ARC_1_3/temp1[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_3  ( .A1(n1506), .A2(n143), .Z(
        \MC_ARK_ARC_1_3/temp4[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_2  ( .A1(\RI5[3][189] ), .A2(n131), .Z(
        \MC_ARK_ARC_1_3/temp4[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_1  ( .A1(\RI5[3][190] ), .A2(n10), .Z(
        \MC_ARK_ARC_1_3/temp4[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_6_1  ( .A1(\RI5[3][28] ), .A2(\RI5[3][64] ), .Z(
        \MC_ARK_ARC_1_3/temp3[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_6_1  ( .A1(\RI5[3][124] ), .A2(\RI5[3][100] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_6_0  ( .A1(\RI5[3][101] ), .A2(\RI5[3][125] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_5_5  ( .A1(\MC_ARK_ARC_1_3/temp5[156] ), .A2(
        \MC_ARK_ARC_1_3/temp6[156] ), .Z(\MC_ARK_ARC_1_3/buf_output[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_5_5  ( .A1(\MC_ARK_ARC_1_3/temp3[156] ), .A2(
        \MC_ARK_ARC_1_3/temp4[156] ), .Z(\MC_ARK_ARC_1_3/temp6[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_5_5  ( .A1(\MC_ARK_ARC_1_3/temp2[156] ), .A2(
        \MC_ARK_ARC_1_3/temp1[156] ), .Z(\MC_ARK_ARC_1_3/temp5[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[0] ), 
        .A2(n535), .Z(\MC_ARK_ARC_1_3/temp4[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_5_5  ( .A1(\RI5[3][66] ), .A2(\RI5[3][30] ), .Z(
        \MC_ARK_ARC_1_3/temp3[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_5_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[102] ), 
        .A2(\RI5[3][126] ), .Z(\MC_ARK_ARC_1_3/temp2[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_5_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[156] ), 
        .A2(\RI5[3][150] ), .Z(\MC_ARK_ARC_1_3/temp1[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_5_4  ( .A1(\MC_ARK_ARC_1_3/temp4[157] ), .A2(
        \MC_ARK_ARC_1_3/temp3[157] ), .Z(\MC_ARK_ARC_1_3/temp6[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[1] ), 
        .A2(n203), .Z(\MC_ARK_ARC_1_3/temp4[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_5_4  ( .A1(\RI5[3][67] ), .A2(\RI5[3][31] ), .Z(
        \MC_ARK_ARC_1_3/temp3[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_5_4  ( .A1(\RI5[3][127] ), .A2(\RI5[3][103] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_3  ( .A1(\RI5[3][2] ), .A2(n181), .Z(
        \MC_ARK_ARC_1_3/temp4[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_5_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[32] ), 
        .A2(\RI5[3][68] ), .Z(\MC_ARK_ARC_1_3/temp3[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_5_3  ( .A1(\RI5[3][152] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[158] ), .Z(\MC_ARK_ARC_1_3/temp1[158] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_5_2  ( .A1(\MC_ARK_ARC_1_3/temp2[159] ), .A2(
        \MC_ARK_ARC_1_3/temp1[159] ), .Z(\MC_ARK_ARC_1_3/temp5[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_2  ( .A1(\RI5[3][3] ), .A2(n454), .Z(
        \MC_ARK_ARC_1_3/temp4[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_5_2  ( .A1(\RI5[3][33] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[69] ), .Z(\MC_ARK_ARC_1_3/temp3[159] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_5_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[129] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[105] ), .Z(
        \MC_ARK_ARC_1_3/temp2[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_5_2  ( .A1(\RI5[3][153] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[159] ), .Z(\MC_ARK_ARC_1_3/temp1[159] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_5_1  ( .A1(\MC_ARK_ARC_1_3/temp5[160] ), .A2(
        \MC_ARK_ARC_1_3/temp6[160] ), .Z(\MC_ARK_ARC_1_3/buf_output[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_5_1  ( .A1(\MC_ARK_ARC_1_3/temp4[160] ), .A2(
        \MC_ARK_ARC_1_3/temp3[160] ), .Z(\MC_ARK_ARC_1_3/temp6[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_1  ( .A1(\RI5[3][4] ), .A2(n67), .Z(
        \MC_ARK_ARC_1_3/temp4[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_5_1  ( .A1(\RI5[3][70] ), .A2(\RI5[3][34] ), .Z(
        \MC_ARK_ARC_1_3/temp3[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_5_1  ( .A1(\RI5[3][130] ), .A2(\RI5[3][106] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_5_1  ( .A1(\RI5[3][160] ), .A2(\RI5[3][154] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_5_0  ( .A1(\MC_ARK_ARC_1_3/temp5[161] ), .A2(
        \MC_ARK_ARC_1_3/temp6[161] ), .Z(\MC_ARK_ARC_1_3/buf_output[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_5_0  ( .A1(\MC_ARK_ARC_1_3/temp4[161] ), .A2(
        \MC_ARK_ARC_1_3/temp3[161] ), .Z(\MC_ARK_ARC_1_3/temp6[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_5_0  ( .A1(\MC_ARK_ARC_1_3/temp2[161] ), .A2(
        \MC_ARK_ARC_1_3/temp1[161] ), .Z(\MC_ARK_ARC_1_3/temp5[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[5] ), 
        .A2(n452), .Z(\MC_ARK_ARC_1_3/temp4[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_5_0  ( .A1(\RI5[3][35] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[71] ), .Z(\MC_ARK_ARC_1_3/temp3[161] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_5_0  ( .A1(\RI5[3][107] ), .A2(\RI5[3][131] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_5_0  ( .A1(\RI5[3][161] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[155] ), .Z(\MC_ARK_ARC_1_3/temp1[161] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_4_5  ( .A1(\RI5[3][6] ), .A2(n529), .Z(
        \MC_ARK_ARC_1_3/temp4[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_4_5  ( .A1(\RI5[3][72] ), .A2(\RI5[3][36] ), .Z(
        \MC_ARK_ARC_1_3/temp3[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_4_5  ( .A1(\SB2_3_10/buf_output[0] ), .A2(
        \RI5[3][162] ), .Z(\MC_ARK_ARC_1_3/temp1[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_4_4  ( .A1(\MC_ARK_ARC_1_3/temp3[163] ), .A2(
        \MC_ARK_ARC_1_3/temp4[163] ), .Z(\MC_ARK_ARC_1_3/temp6[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_4_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[7] ), 
        .A2(n206), .Z(\MC_ARK_ARC_1_3/temp4[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_4_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[37] ), 
        .A2(\RI5[3][73] ), .Z(\MC_ARK_ARC_1_3/temp3[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_4_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[157] ), 
        .A2(\RI5[3][163] ), .Z(\MC_ARK_ARC_1_3/temp1[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_4_3  ( .A1(\RI5[3][8] ), .A2(n142), .Z(
        \MC_ARK_ARC_1_3/temp4[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_4_2  ( .A1(\RI5[3][9] ), .A2(n450), .Z(
        \MC_ARK_ARC_1_3/temp4[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_4_2  ( .A1(\RI5[3][75] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[39] ), .Z(\MC_ARK_ARC_1_3/temp3[165] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_4_2  ( .A1(\RI5[3][135] ), .A2(\RI5[3][111] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_4_1  ( .A1(\RI5[3][136] ), .A2(\RI5[3][112] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_4_1  ( .A1(\RI5[3][160] ), .A2(\RI5[3][166] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_4_0  ( .A1(\RI5[3][11] ), .A2(n448), .Z(
        \MC_ARK_ARC_1_3/temp4[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_4_0  ( .A1(\RI5[3][137] ), .A2(\RI5[3][113] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_4_0  ( .A1(\RI5[3][167] ), .A2(\RI5[3][161] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_3_5  ( .A1(\MC_ARK_ARC_1_3/temp5[168] ), .A2(
        \MC_ARK_ARC_1_3/temp6[168] ), .Z(\MC_ARK_ARC_1_3/buf_output[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_3_5  ( .A1(\MC_ARK_ARC_1_3/temp3[168] ), .A2(
        \MC_ARK_ARC_1_3/temp4[168] ), .Z(\MC_ARK_ARC_1_3/temp6[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_3_5  ( .A1(\MC_ARK_ARC_1_3/temp2[168] ), .A2(
        \MC_ARK_ARC_1_3/temp1[168] ), .Z(\MC_ARK_ARC_1_3/temp5[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_5  ( .A1(\RI5[3][12] ), .A2(n523), .Z(
        \MC_ARK_ARC_1_3/temp4[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_3_5  ( .A1(\RI5[3][42] ), .A2(\RI5[3][78] ), .Z(
        \MC_ARK_ARC_1_3/temp3[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_3_5  ( .A1(\RI5[3][114] ), .A2(\RI5[3][138] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_3_5  ( .A1(\RI5[3][162] ), .A2(\RI5[3][168] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_3_4  ( .A1(\MC_ARK_ARC_1_3/temp3[169] ), .A2(
        \MC_ARK_ARC_1_3/temp4[169] ), .Z(\MC_ARK_ARC_1_3/temp6[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_4  ( .A1(\RI5[3][13] ), .A2(n446), .Z(
        \MC_ARK_ARC_1_3/temp4[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_3_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[43] ), 
        .A2(\RI5[3][79] ), .Z(\MC_ARK_ARC_1_3/temp3[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_3_4  ( .A1(\RI5[3][139] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_3/temp2[169] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_3_4  ( .A1(\RI5[3][163] ), .A2(\RI5[3][169] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_3_2  ( .A1(\MC_ARK_ARC_1_3/temp3[171] ), .A2(
        \MC_ARK_ARC_1_3/temp4[171] ), .Z(\MC_ARK_ARC_1_3/temp6[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[15] ), 
        .A2(n444), .Z(\MC_ARK_ARC_1_3/temp4[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_3_2  ( .A1(\RI5[3][81] ), .A2(\RI5[3][45] ), .Z(
        \MC_ARK_ARC_1_3/temp3[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_1  ( .A1(\RI5[3][16] ), .A2(n79), .Z(
        \MC_ARK_ARC_1_3/temp4[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_3_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[46] ), 
        .A2(\RI5[3][82] ), .Z(\MC_ARK_ARC_1_3/temp3[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_3_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[118] ), .Z(
        \MC_ARK_ARC_1_3/temp2[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_3_0  ( .A1(\MC_ARK_ARC_1_3/temp4[173] ), .A2(
        \MC_ARK_ARC_1_3/temp3[173] ), .Z(\MC_ARK_ARC_1_3/temp6[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_0  ( .A1(\RI5[3][17] ), .A2(n49), .Z(
        \MC_ARK_ARC_1_3/temp4[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_3_0  ( .A1(\RI5[3][83] ), .A2(\RI5[3][47] ), .Z(
        \MC_ARK_ARC_1_3/temp3[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_5  ( .A1(\RI5[3][18] ), .A2(n182), .Z(
        \MC_ARK_ARC_1_3/temp4[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[19] ), 
        .A2(n172), .Z(\MC_ARK_ARC_1_3/temp4[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_2_4  ( .A1(\RI5[3][175] ), .A2(\RI5[3][169] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_2_3  ( .A1(\RI5[3][146] ), .A2(\RI5[3][122] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[21] ), 
        .A2(n97), .Z(\MC_ARK_ARC_1_3/temp4[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_2_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[147] ), 
        .A2(n575), .Z(\MC_ARK_ARC_1_3/temp2[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_1  ( .A1(\RI5[3][22] ), .A2(n121), .Z(
        \MC_ARK_ARC_1_3/temp4[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_2_1  ( .A1(\RI5[3][88] ), .A2(\RI5[3][52] ), .Z(
        \MC_ARK_ARC_1_3/temp3[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_2_1  ( .A1(\RI5[3][124] ), .A2(\RI5[3][148] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_2_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .A2(\RI5[3][172] ), .Z(\MC_ARK_ARC_1_3/temp1[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_2_0  ( .A1(\MC_ARK_ARC_1_3/temp1[179] ), .A2(
        \MC_ARK_ARC_1_3/temp2[179] ), .Z(\MC_ARK_ARC_1_3/temp5[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_0  ( .A1(\RI5[3][23] ), .A2(n96), .Z(
        \MC_ARK_ARC_1_3/temp4[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_2_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .A2(\RI5[3][89] ), .Z(\MC_ARK_ARC_1_3/temp3[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_2_0  ( .A1(\RI5[3][149] ), .A2(\RI5[3][125] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_1_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[24] ), 
        .A2(n513), .Z(\MC_ARK_ARC_1_3/temp4[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_1_5  ( .A1(\RI5[3][54] ), .A2(\RI5[3][90] ), .Z(
        \MC_ARK_ARC_1_3/temp3[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_1_4  ( .A1(\RI5[3][25] ), .A2(n435), .Z(
        \MC_ARK_ARC_1_3/temp4[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_1_4  ( .A1(\RI5[3][55] ), .A2(\RI5[3][91] ), .Z(
        \MC_ARK_ARC_1_3/temp3[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_1_4  ( .A1(\RI5[3][181] ), .A2(\RI5[3][175] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_1_3  ( .A1(\RI5[3][26] ), .A2(n106), .Z(
        \MC_ARK_ARC_1_3/temp4[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_1_1  ( .A1(\MC_ARK_ARC_1_3/temp4[184] ), .A2(
        \MC_ARK_ARC_1_3/temp3[184] ), .Z(\MC_ARK_ARC_1_3/temp6[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_1_1  ( .A1(\RI5[3][28] ), .A2(n509), .Z(
        \MC_ARK_ARC_1_3/temp4[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_1_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[94] ), 
        .A2(\RI5[3][58] ), .Z(\MC_ARK_ARC_1_3/temp3[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_1_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[184] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[178] ), .Z(
        \MC_ARK_ARC_1_3/temp1[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_1_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[29] ), 
        .A2(n101), .Z(\MC_ARK_ARC_1_3/temp4[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_1_0  ( .A1(\RI5[3][185] ), .A2(\RI5[3][179] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_0_5  ( .A1(\MC_ARK_ARC_1_3/temp5[186] ), .A2(
        \MC_ARK_ARC_1_3/temp6[186] ), .Z(\MC_ARK_ARC_1_3/buf_output[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_0_5  ( .A1(\MC_ARK_ARC_1_3/temp4[186] ), .A2(
        \MC_ARK_ARC_1_3/temp3[186] ), .Z(\MC_ARK_ARC_1_3/temp6[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_0_5  ( .A1(\MC_ARK_ARC_1_3/temp1[186] ), .A2(
        \MC_ARK_ARC_1_3/temp2[186] ), .Z(\MC_ARK_ARC_1_3/temp5[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_0_5  ( .A1(\RI5[3][30] ), .A2(n202), .Z(
        \MC_ARK_ARC_1_3/temp4[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_0_5  ( .A1(\RI5[3][60] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[96] ), .Z(\MC_ARK_ARC_1_3/temp3[186] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_0_5  ( .A1(\RI5[3][132] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[156] ), .Z(\MC_ARK_ARC_1_3/temp2[186] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_0_5  ( .A1(\RI5[3][186] ), .A2(\RI5[3][180] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_0_4  ( .A1(\RI5[3][31] ), .A2(n58), .Z(
        \MC_ARK_ARC_1_3/temp4[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_0_4  ( .A1(\RI5[3][97] ), .A2(\RI5[3][61] ), .Z(
        \MC_ARK_ARC_1_3/temp3[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_0_4  ( .A1(\RI5[3][181] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[187] ), .Z(\MC_ARK_ARC_1_3/temp1[187] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_0_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[32] ), 
        .A2(n113), .Z(\MC_ARK_ARC_1_3/temp4[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_0_3  ( .A1(n1506), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[182] ), .Z(\MC_ARK_ARC_1_3/temp1[188] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_0_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[183] ), 
        .A2(\RI5[3][189] ), .Z(\MC_ARK_ARC_1_3/temp1[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_0_1  ( .A1(\MC_ARK_ARC_1_3/temp4[190] ), .A2(
        \MC_ARK_ARC_1_3/temp3[190] ), .Z(\MC_ARK_ARC_1_3/temp6[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_0_1  ( .A1(\RI5[3][34] ), .A2(n505), .Z(
        \MC_ARK_ARC_1_3/temp4[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_0_1  ( .A1(\RI5[3][190] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[184] ), .Z(\MC_ARK_ARC_1_3/temp1[190] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_31_5  ( .A1(\RI5[4][36] ), .A2(n118), .Z(
        \MC_ARK_ARC_1_4/temp4[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_31_4  ( .A1(\MC_ARK_ARC_1_4/temp3[1] ), .A2(
        \MC_ARK_ARC_1_4/temp4[1] ), .Z(\MC_ARK_ARC_1_4/temp6[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_31_4  ( .A1(\RI5[4][37] ), .A2(n494), .Z(
        \MC_ARK_ARC_1_4/temp4[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_31_4  ( .A1(\RI5[4][187] ), .A2(\RI5[4][1] ), .Z(
        \MC_ARK_ARC_1_4/temp1[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_31_3  ( .A1(\RI5[4][38] ), .A2(n566), .Z(
        \MC_ARK_ARC_1_4/temp4[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_31_3  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[188] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[2] ), .Z(\MC_ARK_ARC_1_4/temp1[2] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_31_2  ( .A1(\MC_ARK_ARC_1_4/temp5[3] ), .A2(
        \MC_ARK_ARC_1_4/temp6[3] ), .Z(\MC_ARK_ARC_1_4/buf_output[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_31_2  ( .A1(\MC_ARK_ARC_1_4/temp3[3] ), .A2(
        \MC_ARK_ARC_1_4/temp4[3] ), .Z(\MC_ARK_ARC_1_4/temp6[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_31_2  ( .A1(\SB2_4_27/buf_output[3] ), .A2(n191), 
        .Z(\MC_ARK_ARC_1_4/temp4[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_31_2  ( .A1(\SB2_4_16/buf_output[3] ), .A2(
        \SB2_4_22/buf_output[3] ), .Z(\MC_ARK_ARC_1_4/temp3[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_31_1  ( .A1(\MC_ARK_ARC_1_4/temp6[4] ), .A2(
        \MC_ARK_ARC_1_4/temp5[4] ), .Z(\MC_ARK_ARC_1_4/buf_output[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_31_1  ( .A1(\MC_ARK_ARC_1_4/temp3[4] ), .A2(
        \MC_ARK_ARC_1_4/temp4[4] ), .Z(\MC_ARK_ARC_1_4/temp6[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_31_1  ( .A1(\MC_ARK_ARC_1_4/temp1[4] ), .A2(
        \MC_ARK_ARC_1_4/temp2[4] ), .Z(\MC_ARK_ARC_1_4/temp5[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_31_1  ( .A1(\RI5[4][40] ), .A2(n554), .Z(
        \MC_ARK_ARC_1_4/temp4[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_31_1  ( .A1(\RI5[4][106] ), .A2(\RI5[4][70] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_31_1  ( .A1(\RI5[4][166] ), .A2(\RI5[4][142] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_31_1  ( .A1(\RI5[4][4] ), .A2(\RI5[4][190] ), .Z(
        \MC_ARK_ARC_1_4/temp1[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_31_0  ( .A1(\RI5[4][41] ), .A2(n29), .Z(
        \MC_ARK_ARC_1_4/temp4[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_30_5  ( .A1(\RI5[4][42] ), .A2(n6), .Z(
        \MC_ARK_ARC_1_4/temp4[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_30_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[108] ), 
        .A2(\RI5[4][72] ), .Z(\MC_ARK_ARC_1_4/temp3[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_30_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[168] ), 
        .A2(\RI5[4][144] ), .Z(\MC_ARK_ARC_1_4/temp2[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_30_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[43] ), 
        .A2(n112), .Z(\MC_ARK_ARC_1_4/temp4[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_30_4  ( .A1(\RI5[4][109] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[73] ), .Z(\MC_ARK_ARC_1_4/temp3[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_30_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[169] ), 
        .A2(\RI5[4][145] ), .Z(\MC_ARK_ARC_1_4/temp2[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_30_4  ( .A1(\RI5[4][1] ), .A2(\RI5[4][7] ), .Z(
        \MC_ARK_ARC_1_4/temp1[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_30_3  ( .A1(\MC_ARK_ARC_1_4/temp6[8] ), .A2(
        \MC_ARK_ARC_1_4/temp5[8] ), .Z(\MC_ARK_ARC_1_4/buf_output[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_30_3  ( .A1(\RI5[4][44] ), .A2(n198), .Z(
        \MC_ARK_ARC_1_4/temp4[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_30_3  ( .A1(\RI5[4][74] ), .A2(\RI5[4][110] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_30_2  ( .A1(\MC_ARK_ARC_1_4/temp3[9] ), .A2(
        \MC_ARK_ARC_1_4/temp4[9] ), .Z(\MC_ARK_ARC_1_4/temp6[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_30_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[45] ), 
        .A2(n219), .Z(\MC_ARK_ARC_1_4/temp4[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_30_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[75] ), 
        .A2(\RI5[4][111] ), .Z(\MC_ARK_ARC_1_4/temp3[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_30_2  ( .A1(\RI5[4][147] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[171] ), .Z(\MC_ARK_ARC_1_4/temp2[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_30_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[9] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[3] ), .Z(\MC_ARK_ARC_1_4/temp1[9] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_30_1  ( .A1(\MC_ARK_ARC_1_4/temp4[10] ), .A2(
        \MC_ARK_ARC_1_4/temp3[10] ), .Z(\MC_ARK_ARC_1_4/temp6[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_30_1  ( .A1(\RI5[4][46] ), .A2(n521), .Z(
        \MC_ARK_ARC_1_4/temp4[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_30_1  ( .A1(\RI5[4][112] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_4/temp3[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_30_1  ( .A1(\RI5[4][172] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[148] ), .Z(\MC_ARK_ARC_1_4/temp2[10] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_30_1  ( .A1(\RI5[4][10] ), .A2(\RI5[4][4] ), .Z(
        \MC_ARK_ARC_1_4/temp1[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_29_5  ( .A1(\MC_ARK_ARC_1_4/temp6[12] ), .A2(
        \MC_ARK_ARC_1_4/temp5[12] ), .Z(\MC_ARK_ARC_1_4/buf_output[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_29_5  ( .A1(\MC_ARK_ARC_1_4/temp4[12] ), .A2(
        \MC_ARK_ARC_1_4/temp3[12] ), .Z(\MC_ARK_ARC_1_4/temp6[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_29_5  ( .A1(\MC_ARK_ARC_1_4/temp1[12] ), .A2(
        \MC_ARK_ARC_1_4/temp2[12] ), .Z(\MC_ARK_ARC_1_4/temp5[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_29_5  ( .A1(\RI5[4][48] ), .A2(n508), .Z(
        \MC_ARK_ARC_1_4/temp4[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_29_5  ( .A1(\RI5[4][114] ), .A2(\RI5[4][78] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_29_5  ( .A1(\RI5[4][174] ), .A2(\RI5[4][150] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_29_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[12] ), 
        .A2(\RI5[4][6] ), .Z(\MC_ARK_ARC_1_4/temp1[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_29_4  ( .A1(\MC_ARK_ARC_1_4/temp2[13] ), .A2(
        \MC_ARK_ARC_1_4/temp1[13] ), .Z(\MC_ARK_ARC_1_4/temp5[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_29_4  ( .A1(\RI5[4][49] ), .A2(n425), .Z(
        \MC_ARK_ARC_1_4/temp4[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_29_4  ( .A1(\RI5[4][79] ), .A2(\RI5[4][115] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_29_4  ( .A1(n3165), .A2(\RI5[4][151] ), .Z(
        \MC_ARK_ARC_1_4/temp2[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_29_4  ( .A1(\RI5[4][13] ), .A2(\RI5[4][7] ), .Z(
        \MC_ARK_ARC_1_4/temp1[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_29_3  ( .A1(\MC_ARK_ARC_1_4/temp6[14] ), .A2(
        \MC_ARK_ARC_1_4/temp5[14] ), .Z(\MC_ARK_ARC_1_4/buf_output[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_29_3  ( .A1(\MC_ARK_ARC_1_4/temp4[14] ), .A2(
        \MC_ARK_ARC_1_4/temp3[14] ), .Z(\MC_ARK_ARC_1_4/temp6[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_29_3  ( .A1(\RI5[4][50] ), .A2(n497), .Z(
        \MC_ARK_ARC_1_4/temp4[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_29_3  ( .A1(\RI5[4][116] ), .A2(\RI5[4][80] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_29_2  ( .A1(\RI5[4][51] ), .A2(n414), .Z(
        \MC_ARK_ARC_1_4/temp4[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_29_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[9] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[15] ), .Z(\MC_ARK_ARC_1_4/temp1[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_29_1  ( .A1(\RI5[4][52] ), .A2(n212), .Z(
        \MC_ARK_ARC_1_4/temp4[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_29_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[118] ), 
        .A2(\RI5[4][82] ), .Z(\MC_ARK_ARC_1_4/temp3[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_29_1  ( .A1(\RI5[4][178] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[154] ), .Z(\MC_ARK_ARC_1_4/temp2[16] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_29_1  ( .A1(\RI5[4][10] ), .A2(\RI5[4][16] ), .Z(
        \MC_ARK_ARC_1_4/temp1[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_29_0  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[53] ), 
        .A2(n558), .Z(\MC_ARK_ARC_1_4/temp4[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_28_5  ( .A1(\MC_ARK_ARC_1_4/temp5[18] ), .A2(
        \MC_ARK_ARC_1_4/temp6[18] ), .Z(\MC_ARK_ARC_1_4/buf_output[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_28_5  ( .A1(\MC_ARK_ARC_1_4/temp3[18] ), .A2(
        \MC_ARK_ARC_1_4/temp4[18] ), .Z(\MC_ARK_ARC_1_4/temp6[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_28_5  ( .A1(\MC_ARK_ARC_1_4/temp2[18] ), .A2(
        \MC_ARK_ARC_1_4/temp1[18] ), .Z(\MC_ARK_ARC_1_4/temp5[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_28_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[54] ), 
        .A2(n477), .Z(\MC_ARK_ARC_1_4/temp4[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_28_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[120] ), 
        .A2(\RI5[4][84] ), .Z(\MC_ARK_ARC_1_4/temp3[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_28_5  ( .A1(\RI5[4][180] ), .A2(\RI5[4][156] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_28_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[18] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[12] ), .Z(\MC_ARK_ARC_1_4/temp1[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_28_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[55] ), 
        .A2(n547), .Z(\MC_ARK_ARC_1_4/temp4[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_28_4  ( .A1(\SB2_4_21/buf_output[1] ), .A2(
        \RI5[4][121] ), .Z(\MC_ARK_ARC_1_4/temp3[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_28_3  ( .A1(\RI5[4][56] ), .A2(n63), .Z(
        \MC_ARK_ARC_1_4/temp4[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_28_2  ( .A1(\MC_ARK_ARC_1_4/temp2[21] ), .A2(
        \MC_ARK_ARC_1_4/temp1[21] ), .Z(\MC_ARK_ARC_1_4/temp5[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_28_2  ( .A1(\RI5[4][57] ), .A2(n143), .Z(
        \MC_ARK_ARC_1_4/temp4[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_28_2  ( .A1(\RI5[4][159] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[183] ), .Z(\MC_ARK_ARC_1_4/temp2[21] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_28_2  ( .A1(\RI5[4][21] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[15] ), .Z(\MC_ARK_ARC_1_4/temp1[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_28_1  ( .A1(\MC_ARK_ARC_1_4/temp1[22] ), .A2(
        \MC_ARK_ARC_1_4/temp2[22] ), .Z(\MC_ARK_ARC_1_4/temp5[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_28_1  ( .A1(\RI5[4][58] ), .A2(n209), .Z(
        \MC_ARK_ARC_1_4/temp4[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_28_1  ( .A1(\RI5[4][124] ), .A2(\RI5[4][88] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_28_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[184] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[160] ), .Z(
        \MC_ARK_ARC_1_4/temp2[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_28_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[22] ), 
        .A2(\RI5[4][16] ), .Z(\MC_ARK_ARC_1_4/temp1[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_28_0  ( .A1(\MC_ARK_ARC_1_4/temp5[23] ), .A2(
        \MC_ARK_ARC_1_4/temp6[23] ), .Z(\MC_ARK_ARC_1_4/buf_output[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_28_0  ( .A1(\RI5[4][59] ), .A2(n525), .Z(
        \MC_ARK_ARC_1_4/temp4[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_27_5  ( .A1(\RI5[4][60] ), .A2(n442), .Z(
        \MC_ARK_ARC_1_4/temp4[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_27_5  ( .A1(\RI5[4][186] ), .A2(\RI5[4][162] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_27_5  ( .A1(\RI5[4][24] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[18] ), .Z(\MC_ARK_ARC_1_4/temp1[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_27_4  ( .A1(\RI5[4][61] ), .A2(n138), .Z(
        \MC_ARK_ARC_1_4/temp4[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_27_4  ( .A1(\RI5[4][127] ), .A2(\RI5[4][91] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_27_4  ( .A1(\RI5[4][25] ), .A2(\RI5[4][19] ), .Z(
        \MC_ARK_ARC_1_4/temp1[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_27_3  ( .A1(\RI5[4][62] ), .A2(n429), .Z(
        \MC_ARK_ARC_1_4/temp4[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_27_3  ( .A1(\RI5[4][92] ), .A2(\RI5[4][128] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_27_3  ( .A1(\RI5[4][164] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[188] ), .Z(\MC_ARK_ARC_1_4/temp2[26] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_27_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[63] ), 
        .A2(n132), .Z(\MC_ARK_ARC_1_4/temp4[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_27_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[129] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[93] ), .Z(\MC_ARK_ARC_1_4/temp3[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_27_1  ( .A1(\MC_ARK_ARC_1_4/temp1[28] ), .A2(
        \MC_ARK_ARC_1_4/temp2[28] ), .Z(\MC_ARK_ARC_1_4/temp5[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_27_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[64] ), 
        .A2(n187), .Z(\MC_ARK_ARC_1_4/temp4[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_27_1  ( .A1(\RI5[4][190] ), .A2(\RI5[4][166] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_27_1  ( .A1(\RI5[4][28] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_4/temp1[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_27_0  ( .A1(\RI5[4][65] ), .A2(n156), .Z(
        \MC_ARK_ARC_1_4/temp4[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_27_0  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[167] ), 
        .A2(\RI5[4][191] ), .Z(\MC_ARK_ARC_1_4/temp2[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_27_0  ( .A1(\RI5[4][29] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[23] ), .Z(\MC_ARK_ARC_1_4/temp1[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_26_5  ( .A1(\MC_ARK_ARC_1_4/temp6[30] ), .A2(
        \MC_ARK_ARC_1_4/temp5[30] ), .Z(\MC_ARK_ARC_1_4/buf_output[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_26_5  ( .A1(\MC_ARK_ARC_1_4/temp1[30] ), .A2(
        \MC_ARK_ARC_1_4/temp2[30] ), .Z(\MC_ARK_ARC_1_4/temp5[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_26_5  ( .A1(\RI5[4][66] ), .A2(n193), .Z(
        \MC_ARK_ARC_1_4/temp4[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_26_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[132] ), 
        .A2(\RI5[4][96] ), .Z(\MC_ARK_ARC_1_4/temp3[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_26_5  ( .A1(\RI5[4][0] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[168] ), .Z(\MC_ARK_ARC_1_4/temp2[30] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_26_5  ( .A1(\RI5[4][30] ), .A2(\RI5[4][24] ), .Z(
        \MC_ARK_ARC_1_4/temp1[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_26_4  ( .A1(\MC_ARK_ARC_1_4/temp1[31] ), .A2(
        \MC_ARK_ARC_1_4/temp2[31] ), .Z(\MC_ARK_ARC_1_4/temp5[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_26_4  ( .A1(\RI5[4][67] ), .A2(n482), .Z(
        \MC_ARK_ARC_1_4/temp4[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_26_4  ( .A1(\RI5[4][133] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[97] ), .Z(\MC_ARK_ARC_1_4/temp3[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_26_4  ( .A1(\RI5[4][31] ), .A2(\RI5[4][25] ), .Z(
        \MC_ARK_ARC_1_4/temp1[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_26_3  ( .A1(\MC_ARK_ARC_1_4/temp5[32] ), .A2(
        \MC_ARK_ARC_1_4/temp6[32] ), .Z(\MC_ARK_ARC_1_4/buf_output[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_26_3  ( .A1(\SB2_4_23/buf_output[2] ), .A2(n104), 
        .Z(\MC_ARK_ARC_1_4/temp4[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_26_3  ( .A1(\RI5[4][98] ), .A2(\RI5[4][134] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_26_2  ( .A1(\RI5[4][33] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[27] ), .Z(\MC_ARK_ARC_1_4/temp1[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_26_1  ( .A1(\MC_ARK_ARC_1_4/temp6[34] ), .A2(
        \MC_ARK_ARC_1_4/temp5[34] ), .Z(\MC_ARK_ARC_1_4/buf_output[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_26_1  ( .A1(\MC_ARK_ARC_1_4/temp4[34] ), .A2(
        \MC_ARK_ARC_1_4/temp3[34] ), .Z(\MC_ARK_ARC_1_4/temp6[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_26_1  ( .A1(\MC_ARK_ARC_1_4/temp2[34] ), .A2(
        \MC_ARK_ARC_1_4/temp1[34] ), .Z(\MC_ARK_ARC_1_4/temp5[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_26_1  ( .A1(\RI5[4][70] ), .A2(n123), .Z(
        \MC_ARK_ARC_1_4/temp4[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_26_1  ( .A1(\RI5[4][136] ), .A2(\RI5[4][100] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_26_1  ( .A1(\RI5[4][4] ), .A2(\RI5[4][172] ), .Z(
        \MC_ARK_ARC_1_4/temp2[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_26_1  ( .A1(\RI5[4][28] ), .A2(\RI5[4][34] ), .Z(
        \MC_ARK_ARC_1_4/temp1[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_26_0  ( .A1(\RI5[4][71] ), .A2(n28), .Z(
        \MC_ARK_ARC_1_4/temp4[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_25_5  ( .A1(\MC_ARK_ARC_1_4/temp5[36] ), .A2(
        \MC_ARK_ARC_1_4/temp6[36] ), .Z(\MC_ARK_ARC_1_4/buf_output[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_25_5  ( .A1(\MC_ARK_ARC_1_4/temp1[36] ), .A2(
        \MC_ARK_ARC_1_4/temp2[36] ), .Z(\MC_ARK_ARC_1_4/temp5[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_25_5  ( .A1(\RI5[4][72] ), .A2(n105), .Z(
        \MC_ARK_ARC_1_4/temp4[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_25_5  ( .A1(\RI5[4][138] ), .A2(\RI5[4][102] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_25_5  ( .A1(\RI5[4][6] ), .A2(\RI5[4][174] ), .Z(
        \MC_ARK_ARC_1_4/temp2[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_25_4  ( .A1(\MC_ARK_ARC_1_4/temp6[37] ), .A2(
        \MC_ARK_ARC_1_4/temp5[37] ), .Z(\MC_ARK_ARC_1_4/buf_output[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_25_4  ( .A1(\MC_ARK_ARC_1_4/temp3[37] ), .A2(
        \MC_ARK_ARC_1_4/temp4[37] ), .Z(\MC_ARK_ARC_1_4/temp6[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_25_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[73] ), 
        .A2(n447), .Z(\MC_ARK_ARC_1_4/temp4[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_25_4  ( .A1(\RI5[4][139] ), .A2(\RI5[4][103] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_25_4  ( .A1(\RI5[4][37] ), .A2(\RI5[4][31] ), .Z(
        \MC_ARK_ARC_1_4/temp1[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_25_3  ( .A1(\SB2_4_22/buf_output[2] ), .A2(n518), 
        .Z(\MC_ARK_ARC_1_4/temp4[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_25_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[39] ), 
        .A2(\RI5[4][33] ), .Z(\MC_ARK_ARC_1_4/temp1[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_25_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[76] ), 
        .A2(n80), .Z(\MC_ARK_ARC_1_4/temp4[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_25_0  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[77] ), 
        .A2(n422), .Z(\MC_ARK_ARC_1_4/temp4[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_25_0  ( .A1(\RI5[4][107] ), .A2(\RI5[4][143] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_25_0  ( .A1(\RI5[4][35] ), .A2(\RI5[4][41] ), .Z(
        \MC_ARK_ARC_1_4/temp1[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_24_5  ( .A1(\MC_ARK_ARC_1_4/temp3[42] ), .A2(
        \MC_ARK_ARC_1_4/temp4[42] ), .Z(\MC_ARK_ARC_1_4/temp6[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_24_5  ( .A1(\RI5[4][78] ), .A2(n192), .Z(
        \MC_ARK_ARC_1_4/temp4[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_24_5  ( .A1(\RI5[4][144] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[108] ), .Z(\MC_ARK_ARC_1_4/temp3[42] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_24_5  ( .A1(\RI5[4][42] ), .A2(\RI5[4][36] ), .Z(
        \MC_ARK_ARC_1_4/temp1[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_24_4  ( .A1(\MC_ARK_ARC_1_4/temp6[43] ), .A2(
        \MC_ARK_ARC_1_4/temp5[43] ), .Z(\MC_ARK_ARC_1_4/buf_output[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_24_4  ( .A1(\MC_ARK_ARC_1_4/temp3[43] ), .A2(
        \MC_ARK_ARC_1_4/temp4[43] ), .Z(\MC_ARK_ARC_1_4/temp6[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_24_4  ( .A1(\MC_ARK_ARC_1_4/temp1[43] ), .A2(
        \MC_ARK_ARC_1_4/temp2[43] ), .Z(\MC_ARK_ARC_1_4/temp5[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_24_4  ( .A1(\RI5[4][79] ), .A2(n42), .Z(
        \MC_ARK_ARC_1_4/temp4[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_24_4  ( .A1(\RI5[4][13] ), .A2(\RI5[4][181] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_24_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[43] ), 
        .A2(\RI5[4][37] ), .Z(\MC_ARK_ARC_1_4/temp1[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_24_3  ( .A1(\RI5[4][80] ), .A2(n486), .Z(
        \MC_ARK_ARC_1_4/temp4[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_24_2  ( .A1(\MC_ARK_ARC_1_4/temp3[45] ), .A2(
        \MC_ARK_ARC_1_4/temp4[45] ), .Z(\MC_ARK_ARC_1_4/temp6[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_24_2  ( .A1(\RI5[4][81] ), .A2(n555), .Z(
        \MC_ARK_ARC_1_4/temp4[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_24_1  ( .A1(\MC_ARK_ARC_1_4/temp1[46] ), .A2(
        \MC_ARK_ARC_1_4/temp2[46] ), .Z(\MC_ARK_ARC_1_4/temp5[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_24_1  ( .A1(\RI5[4][82] ), .A2(n473), .Z(
        \MC_ARK_ARC_1_4/temp4[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_24_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[148] ), 
        .A2(\RI5[4][112] ), .Z(\MC_ARK_ARC_1_4/temp3[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_24_1  ( .A1(\RI5[4][16] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[184] ), .Z(\MC_ARK_ARC_1_4/temp2[46] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_24_0  ( .A1(\MC_ARK_ARC_1_4/temp3[47] ), .A2(
        \MC_ARK_ARC_1_4/temp4[47] ), .Z(\MC_ARK_ARC_1_4/temp6[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_24_0  ( .A1(\RI5[4][83] ), .A2(n544), .Z(
        \MC_ARK_ARC_1_4/temp4[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_23_5  ( .A1(\MC_ARK_ARC_1_4/temp3[48] ), .A2(
        \MC_ARK_ARC_1_4/temp4[48] ), .Z(\MC_ARK_ARC_1_4/temp6[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_23_5  ( .A1(\RI5[4][84] ), .A2(n461), .Z(
        \MC_ARK_ARC_1_4/temp4[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_23_5  ( .A1(\RI5[4][150] ), .A2(\RI5[4][114] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_23_4  ( .A1(\MC_ARK_ARC_1_4/temp2[49] ), .A2(
        \MC_ARK_ARC_1_4/temp1[49] ), .Z(\MC_ARK_ARC_1_4/temp5[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_23_4  ( .A1(\RI5[4][85] ), .A2(n177), .Z(
        \MC_ARK_ARC_1_4/temp4[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_23_4  ( .A1(\RI5[4][151] ), .A2(\RI5[4][115] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_23_4  ( .A1(\RI5[4][187] ), .A2(\RI5[4][19] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_23_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[43] ), 
        .A2(\RI5[4][49] ), .Z(\MC_ARK_ARC_1_4/temp1[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_23_3  ( .A1(\MC_ARK_ARC_1_4/temp3[50] ), .A2(
        \MC_ARK_ARC_1_4/temp4[50] ), .Z(\MC_ARK_ARC_1_4/temp6[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_23_3  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[86] ), 
        .A2(n206), .Z(\MC_ARK_ARC_1_4/temp4[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_23_2  ( .A1(\MC_ARK_ARC_1_4/temp5[51] ), .A2(
        \MC_ARK_ARC_1_4/temp6[51] ), .Z(\MC_ARK_ARC_1_4/buf_output[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_23_2  ( .A1(\MC_ARK_ARC_1_4/temp1[51] ), .A2(
        \MC_ARK_ARC_1_4/temp2[51] ), .Z(\MC_ARK_ARC_1_4/temp5[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_23_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[87] ), 
        .A2(n199), .Z(\MC_ARK_ARC_1_4/temp4[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_23_2  ( .A1(\RI5[4][21] ), .A2(\RI5[4][189] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_23_2  ( .A1(\RI5[4][51] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[45] ), .Z(\MC_ARK_ARC_1_4/temp1[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_23_1  ( .A1(\MC_ARK_ARC_1_4/temp5[52] ), .A2(
        \MC_ARK_ARC_1_4/temp6[52] ), .Z(\MC_ARK_ARC_1_4/buf_output[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_23_1  ( .A1(\MC_ARK_ARC_1_4/temp3[52] ), .A2(
        \MC_ARK_ARC_1_4/temp4[52] ), .Z(\MC_ARK_ARC_1_4/temp6[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_23_1  ( .A1(\MC_ARK_ARC_1_4/temp1[52] ), .A2(
        \MC_ARK_ARC_1_4/temp2[52] ), .Z(\MC_ARK_ARC_1_4/temp5[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_23_1  ( .A1(\RI5[4][88] ), .A2(n97), .Z(
        \MC_ARK_ARC_1_4/temp4[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_23_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[154] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[118] ), .Z(
        \MC_ARK_ARC_1_4/temp3[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_23_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[22] ), 
        .A2(\RI5[4][190] ), .Z(\MC_ARK_ARC_1_4/temp2[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_23_1  ( .A1(\RI5[4][52] ), .A2(\RI5[4][46] ), .Z(
        \MC_ARK_ARC_1_4/temp1[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_23_0  ( .A1(\MC_ARK_ARC_1_4/temp3[53] ), .A2(
        \MC_ARK_ARC_1_4/temp4[53] ), .Z(\MC_ARK_ARC_1_4/temp6[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_23_0  ( .A1(\RI5[4][89] ), .A2(n16), .Z(
        \MC_ARK_ARC_1_4/temp4[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_23_0  ( .A1(\RI5[4][155] ), .A2(\RI5[4][119] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_22_5  ( .A1(\MC_ARK_ARC_1_4/temp3[54] ), .A2(
        \MC_ARK_ARC_1_4/temp4[54] ), .Z(\MC_ARK_ARC_1_4/temp6[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_22_5  ( .A1(\RI5[4][90] ), .A2(n57), .Z(
        \MC_ARK_ARC_1_4/temp4[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_22_5  ( .A1(\RI5[4][156] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[120] ), .Z(\MC_ARK_ARC_1_4/temp3[54] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_22_5  ( .A1(\RI5[4][0] ), .A2(\RI5[4][24] ), .Z(
        \MC_ARK_ARC_1_4/temp2[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_22_4  ( .A1(\RI5[4][91] ), .A2(n196), .Z(
        \MC_ARK_ARC_1_4/temp4[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_22_4  ( .A1(\RI5[4][157] ), .A2(\RI5[4][121] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_22_4  ( .A1(\RI5[4][25] ), .A2(\RI5[4][1] ), .Z(
        \MC_ARK_ARC_1_4/temp2[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_22_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[55] ), 
        .A2(\RI5[4][49] ), .Z(\MC_ARK_ARC_1_4/temp1[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_22_3  ( .A1(\RI5[4][92] ), .A2(n47), .Z(
        \MC_ARK_ARC_1_4/temp4[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_22_3  ( .A1(\RI5[4][158] ), .A2(\RI5[4][122] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_22_2  ( .A1(\MC_ARK_ARC_1_4/temp3[57] ), .A2(
        \MC_ARK_ARC_1_4/temp4[57] ), .Z(\MC_ARK_ARC_1_4/temp6[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_22_2  ( .A1(\MC_ARK_ARC_1_4/temp1[57] ), .A2(
        \MC_ARK_ARC_1_4/temp2[57] ), .Z(\MC_ARK_ARC_1_4/temp5[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_22_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[93] ), 
        .A2(n213), .Z(\MC_ARK_ARC_1_4/temp4[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_22_2  ( .A1(\RI5[4][159] ), .A2(\RI5[4][123] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_22_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[3] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[27] ), .Z(\MC_ARK_ARC_1_4/temp2[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_22_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[94] ), 
        .A2(n163), .Z(\MC_ARK_ARC_1_4/temp4[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_22_1  ( .A1(\RI5[4][28] ), .A2(\RI5[4][4] ), .Z(
        \MC_ARK_ARC_1_4/temp2[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_22_1  ( .A1(\RI5[4][52] ), .A2(\RI5[4][58] ), .Z(
        \MC_ARK_ARC_1_4/temp1[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_22_0  ( .A1(\MC_ARK_ARC_1_4/temp3[59] ), .A2(
        \MC_ARK_ARC_1_4/temp4[59] ), .Z(\MC_ARK_ARC_1_4/temp6[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_22_0  ( .A1(\RI5[4][95] ), .A2(n478), .Z(
        \MC_ARK_ARC_1_4/temp4[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_21_5  ( .A1(\MC_ARK_ARC_1_4/temp3[60] ), .A2(
        \MC_ARK_ARC_1_4/temp4[60] ), .Z(\MC_ARK_ARC_1_4/temp6[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_21_5  ( .A1(\RI5[4][96] ), .A2(n146), .Z(
        \MC_ARK_ARC_1_4/temp4[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_21_5  ( .A1(\RI5[4][162] ), .A2(\RI5[4][126] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_21_5  ( .A1(\RI5[4][30] ), .A2(\RI5[4][6] ), .Z(
        \MC_ARK_ARC_1_4/temp2[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_21_5  ( .A1(\RI5[4][60] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[54] ), .Z(\MC_ARK_ARC_1_4/temp1[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_21_4  ( .A1(\MC_ARK_ARC_1_4/temp1[61] ), .A2(
        \MC_ARK_ARC_1_4/temp2[61] ), .Z(\MC_ARK_ARC_1_4/temp5[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_21_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[97] ), 
        .A2(n62), .Z(\MC_ARK_ARC_1_4/temp4[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_21_4  ( .A1(\RI5[4][127] ), .A2(\RI5[4][163] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_21_4  ( .A1(\RI5[4][61] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[55] ), .Z(\MC_ARK_ARC_1_4/temp1[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_21_3  ( .A1(\RI5[4][98] ), .A2(n210), .Z(
        \MC_ARK_ARC_1_4/temp4[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_21_2  ( .A1(\MC_ARK_ARC_1_4/temp2[63] ), .A2(
        \MC_ARK_ARC_1_4/temp1[63] ), .Z(\MC_ARK_ARC_1_4/temp5[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_21_2  ( .A1(\RI5[4][99] ), .A2(n217), .Z(
        \MC_ARK_ARC_1_4/temp4[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_21_2  ( .A1(\RI5[4][33] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[9] ), .Z(\MC_ARK_ARC_1_4/temp2[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_21_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[63] ), 
        .A2(\RI5[4][57] ), .Z(\MC_ARK_ARC_1_4/temp1[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_21_1  ( .A1(\MC_ARK_ARC_1_4/temp5[64] ), .A2(
        \MC_ARK_ARC_1_4/temp6[64] ), .Z(\MC_ARK_ARC_1_4/buf_output[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_21_1  ( .A1(\RI5[4][100] ), .A2(n526), .Z(
        \MC_ARK_ARC_1_4/temp4[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_21_1  ( .A1(\RI5[4][166] ), .A2(\RI5[4][130] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_21_1  ( .A1(\RI5[4][34] ), .A2(\RI5[4][10] ), .Z(
        \MC_ARK_ARC_1_4/temp2[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_21_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[64] ), 
        .A2(\RI5[4][58] ), .Z(\MC_ARK_ARC_1_4/temp1[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_21_0  ( .A1(\RI5[4][101] ), .A2(n443), .Z(
        \MC_ARK_ARC_1_4/temp4[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_21_0  ( .A1(\RI5[4][35] ), .A2(\RI5[4][11] ), .Z(
        \MC_ARK_ARC_1_4/temp2[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_20_5  ( .A1(\MC_ARK_ARC_1_4/temp3[66] ), .A2(
        \MC_ARK_ARC_1_4/temp4[66] ), .Z(\MC_ARK_ARC_1_4/temp6[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_20_5  ( .A1(\RI5[4][102] ), .A2(n514), .Z(
        \MC_ARK_ARC_1_4/temp4[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_20_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[168] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[132] ), .Z(
        \MC_ARK_ARC_1_4/temp3[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_20_5  ( .A1(\RI5[4][36] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[12] ), .Z(\MC_ARK_ARC_1_4/temp2[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_20_5  ( .A1(\RI5[4][66] ), .A2(\RI5[4][60] ), .Z(
        \MC_ARK_ARC_1_4/temp1[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_20_4  ( .A1(\MC_ARK_ARC_1_4/temp5[67] ), .A2(
        \MC_ARK_ARC_1_4/temp6[67] ), .Z(\MC_ARK_ARC_1_4/buf_output[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_20_4  ( .A1(\MC_ARK_ARC_1_4/temp3[67] ), .A2(
        \MC_ARK_ARC_1_4/temp4[67] ), .Z(\MC_ARK_ARC_1_4/temp6[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_20_4  ( .A1(\RI5[4][103] ), .A2(n136), .Z(
        \MC_ARK_ARC_1_4/temp4[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_20_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[169] ), 
        .A2(\RI5[4][133] ), .Z(\MC_ARK_ARC_1_4/temp3[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_20_4  ( .A1(\RI5[4][37] ), .A2(\RI5[4][13] ), .Z(
        \MC_ARK_ARC_1_4/temp2[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_20_4  ( .A1(\RI5[4][61] ), .A2(\RI5[4][67] ), .Z(
        \MC_ARK_ARC_1_4/temp1[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_20_3  ( .A1(\MC_ARK_ARC_1_4/temp5[68] ), .A2(
        \MC_ARK_ARC_1_4/temp6[68] ), .Z(\MC_ARK_ARC_1_4/buf_output[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_20_3  ( .A1(\RI5[4][104] ), .A2(n503), .Z(
        \MC_ARK_ARC_1_4/temp4[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_20_2  ( .A1(\RI5[4][105] ), .A2(n8), .Z(
        \MC_ARK_ARC_1_4/temp4[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_20_1  ( .A1(\MC_ARK_ARC_1_4/temp5[70] ), .A2(
        \MC_ARK_ARC_1_4/temp6[70] ), .Z(\MC_ARK_ARC_1_4/buf_output[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_20_1  ( .A1(\MC_ARK_ARC_1_4/temp3[70] ), .A2(
        \MC_ARK_ARC_1_4/temp4[70] ), .Z(\MC_ARK_ARC_1_4/temp6[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_20_1  ( .A1(\RI5[4][106] ), .A2(n491), .Z(
        \MC_ARK_ARC_1_4/temp4[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_20_1  ( .A1(\RI5[4][40] ), .A2(\RI5[4][16] ), .Z(
        \MC_ARK_ARC_1_4/temp2[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_20_0  ( .A1(\RI5[4][107] ), .A2(n563), .Z(
        \MC_ARK_ARC_1_4/temp4[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_20_0  ( .A1(\RI5[4][137] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[173] ), .Z(\MC_ARK_ARC_1_4/temp3[71] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_20_0  ( .A1(\RI5[4][65] ), .A2(\RI5[4][71] ), .Z(
        \MC_ARK_ARC_1_4/temp1[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_19_5  ( .A1(\MC_ARK_ARC_1_4/temp3[72] ), .A2(
        \MC_ARK_ARC_1_4/temp4[72] ), .Z(\MC_ARK_ARC_1_4/temp6[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_19_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[108] ), 
        .A2(n60), .Z(\MC_ARK_ARC_1_4/temp4[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_19_5  ( .A1(\RI5[4][174] ), .A2(\RI5[4][138] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_19_5  ( .A1(\SB2_4_29/buf_output[0] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[18] ), .Z(\MC_ARK_ARC_1_4/temp2[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_19_5  ( .A1(\RI5[4][66] ), .A2(\RI5[4][72] ), .Z(
        \MC_ARK_ARC_1_4/temp1[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_19_4  ( .A1(\MC_ARK_ARC_1_4/temp1[73] ), .A2(
        \MC_ARK_ARC_1_4/temp2[73] ), .Z(\MC_ARK_ARC_1_4/temp5[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_19_4  ( .A1(\RI5[4][109] ), .A2(
        \MC_ARK_ARC_1_3/buf_keyinput[132] ), .Z(\MC_ARK_ARC_1_4/temp4[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_19_4  ( .A1(n3166), .A2(\RI5[4][139] ), .Z(
        \MC_ARK_ARC_1_4/temp3[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_19_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[43] ), 
        .A2(\RI5[4][19] ), .Z(\MC_ARK_ARC_1_4/temp2[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_19_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[73] ), 
        .A2(\RI5[4][67] ), .Z(\MC_ARK_ARC_1_4/temp1[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_19_3  ( .A1(\RI5[4][110] ), .A2(n469), .Z(
        \MC_ARK_ARC_1_4/temp4[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_19_2  ( .A1(\RI5[4][111] ), .A2(n541), .Z(
        \MC_ARK_ARC_1_4/temp4[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_19_1  ( .A1(\MC_ARK_ARC_1_4/temp5[76] ), .A2(
        \MC_ARK_ARC_1_4/temp6[76] ), .Z(\MC_ARK_ARC_1_4/buf_output[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_19_1  ( .A1(\MC_ARK_ARC_1_4/temp3[76] ), .A2(
        \MC_ARK_ARC_1_4/temp4[76] ), .Z(\MC_ARK_ARC_1_4/temp6[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_19_1  ( .A1(\MC_ARK_ARC_1_4/temp2[76] ), .A2(
        \MC_ARK_ARC_1_4/temp1[76] ), .Z(\MC_ARK_ARC_1_4/temp5[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_19_1  ( .A1(\RI5[4][112] ), .A2(n131), .Z(
        \MC_ARK_ARC_1_4/temp4[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_19_1  ( .A1(\RI5[4][178] ), .A2(\RI5[4][142] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_19_1  ( .A1(\RI5[4][46] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_4/temp2[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_19_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[76] ), 
        .A2(\RI5[4][70] ), .Z(\MC_ARK_ARC_1_4/temp1[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_19_0  ( .A1(\RI5[4][113] ), .A2(n531), .Z(
        \MC_ARK_ARC_1_4/temp4[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_19_0  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[23] ), 
        .A2(\RI5[4][47] ), .Z(\MC_ARK_ARC_1_4/temp2[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_18_5  ( .A1(\MC_ARK_ARC_1_4/temp3[78] ), .A2(
        \MC_ARK_ARC_1_4/temp4[78] ), .Z(\MC_ARK_ARC_1_4/temp6[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_18_5  ( .A1(\RI5[4][114] ), .A2(n448), .Z(
        \MC_ARK_ARC_1_4/temp4[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_18_5  ( .A1(\RI5[4][180] ), .A2(\RI5[4][144] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_18_5  ( .A1(\RI5[4][48] ), .A2(\RI5[4][24] ), .Z(
        \MC_ARK_ARC_1_4/temp2[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_18_5  ( .A1(\RI5[4][72] ), .A2(\RI5[4][78] ), .Z(
        \MC_ARK_ARC_1_4/temp1[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_18_4  ( .A1(\MC_ARK_ARC_1_4/temp5[79] ), .A2(
        \MC_ARK_ARC_1_4/temp6[79] ), .Z(\MC_ARK_ARC_1_4/buf_output[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_18_4  ( .A1(\MC_ARK_ARC_1_4/temp3[79] ), .A2(
        \MC_ARK_ARC_1_4/temp4[79] ), .Z(\MC_ARK_ARC_1_4/temp6[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_18_4  ( .A1(\MC_ARK_ARC_1_4/temp1[79] ), .A2(
        \MC_ARK_ARC_1_4/temp2[79] ), .Z(\MC_ARK_ARC_1_4/temp5[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_18_4  ( .A1(\RI5[4][115] ), .A2(n182), .Z(
        \MC_ARK_ARC_1_4/temp4[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_18_4  ( .A1(\RI5[4][181] ), .A2(\RI5[4][145] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_18_4  ( .A1(\RI5[4][25] ), .A2(\RI5[4][49] ), .Z(
        \MC_ARK_ARC_1_4/temp2[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_18_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[73] ), 
        .A2(\RI5[4][79] ), .Z(\MC_ARK_ARC_1_4/temp1[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_18_3  ( .A1(\RI5[4][116] ), .A2(n435), .Z(
        \MC_ARK_ARC_1_4/temp4[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_18_3  ( .A1(\RI5[4][26] ), .A2(\RI5[4][50] ), .Z(
        \MC_ARK_ARC_1_4/temp2[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_18_3  ( .A1(\RI5[4][74] ), .A2(\RI5[4][80] ), .Z(
        \MC_ARK_ARC_1_4/temp1[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_18_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[117] ), 
        .A2(n200), .Z(\MC_ARK_ARC_1_4/temp4[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_18_2  ( .A1(\RI5[4][51] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[27] ), .Z(\MC_ARK_ARC_1_4/temp2[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_18_1  ( .A1(\MC_ARK_ARC_1_4/temp5[82] ), .A2(
        \MC_ARK_ARC_1_4/temp6[82] ), .Z(\MC_ARK_ARC_1_4/buf_output[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_18_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[118] ), 
        .A2(n216), .Z(\MC_ARK_ARC_1_4/temp4[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_18_1  ( .A1(\RI5[4][82] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_4/temp1[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_18_0  ( .A1(\MC_ARK_ARC_1_4/temp3[83] ), .A2(
        \MC_ARK_ARC_1_4/temp4[83] ), .Z(\MC_ARK_ARC_1_4/temp6[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_18_0  ( .A1(\MC_ARK_ARC_1_4/temp1[83] ), .A2(
        \MC_ARK_ARC_1_4/temp2[83] ), .Z(\MC_ARK_ARC_1_4/temp5[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_18_0  ( .A1(\RI5[4][119] ), .A2(n25), .Z(
        \MC_ARK_ARC_1_4/temp4[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_18_0  ( .A1(\RI5[4][29] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[53] ), .Z(\MC_ARK_ARC_1_4/temp2[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_17_5  ( .A1(\MC_ARK_ARC_1_4/temp6[84] ), .A2(
        \MC_ARK_ARC_1_4/temp5[84] ), .Z(\MC_ARK_ARC_1_4/buf_output[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_17_5  ( .A1(\MC_ARK_ARC_1_4/temp3[84] ), .A2(
        \MC_ARK_ARC_1_4/temp4[84] ), .Z(\MC_ARK_ARC_1_4/temp6[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_17_5  ( .A1(\MC_ARK_ARC_1_4/temp2[84] ), .A2(
        \MC_ARK_ARC_1_4/temp1[84] ), .Z(\MC_ARK_ARC_1_4/temp5[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_17_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[120] ), 
        .A2(n568), .Z(\MC_ARK_ARC_1_4/temp4[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_17_5  ( .A1(\RI5[4][186] ), .A2(\RI5[4][150] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_17_5  ( .A1(\RI5[4][30] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[54] ), .Z(\MC_ARK_ARC_1_4/temp2[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_17_5  ( .A1(\RI5[4][84] ), .A2(\RI5[4][78] ), .Z(
        \MC_ARK_ARC_1_4/temp1[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_17_4  ( .A1(\MC_ARK_ARC_1_4/temp3[85] ), .A2(
        \MC_ARK_ARC_1_4/temp4[85] ), .Z(\MC_ARK_ARC_1_4/temp6[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_17_4  ( .A1(\MC_ARK_ARC_1_4/temp1[85] ), .A2(
        \MC_ARK_ARC_1_4/temp2[85] ), .Z(\MC_ARK_ARC_1_4/temp5[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_17_4  ( .A1(\RI5[4][121] ), .A2(n175), .Z(
        \MC_ARK_ARC_1_4/temp4[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_17_4  ( .A1(\RI5[4][187] ), .A2(\RI5[4][151] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_17_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[55] ), 
        .A2(\RI5[4][31] ), .Z(\MC_ARK_ARC_1_4/temp2[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_17_4  ( .A1(\RI5[4][85] ), .A2(\RI5[4][79] ), .Z(
        \MC_ARK_ARC_1_4/temp1[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_17_3  ( .A1(\RI5[4][122] ), .A2(n204), .Z(
        \MC_ARK_ARC_1_4/temp4[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_17_3  ( .A1(\RI5[4][32] ), .A2(\RI5[4][56] ), .Z(
        \MC_ARK_ARC_1_4/temp2[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_17_3  ( .A1(\RI5[4][80] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[86] ), .Z(\MC_ARK_ARC_1_4/temp1[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_17_2  ( .A1(\RI5[4][123] ), .A2(n474), .Z(
        \MC_ARK_ARC_1_4/temp4[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_17_1  ( .A1(\MC_ARK_ARC_1_4/temp3[88] ), .A2(
        \MC_ARK_ARC_1_4/temp4[88] ), .Z(\MC_ARK_ARC_1_4/temp6[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_17_1  ( .A1(\RI5[4][124] ), .A2(n545), .Z(
        \MC_ARK_ARC_1_4/temp4[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_17_1  ( .A1(\RI5[4][190] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[154] ), .Z(\MC_ARK_ARC_1_4/temp3[88] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_17_0  ( .A1(\RI5[4][125] ), .A2(n462), .Z(
        \MC_ARK_ARC_1_4/temp4[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_16_5  ( .A1(\MC_ARK_ARC_1_4/temp5[90] ), .A2(
        \MC_ARK_ARC_1_4/temp6[90] ), .Z(\MC_ARK_ARC_1_4/buf_output[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_16_5  ( .A1(\MC_ARK_ARC_1_4/temp3[90] ), .A2(
        \MC_ARK_ARC_1_4/temp4[90] ), .Z(\MC_ARK_ARC_1_4/temp6[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_16_5  ( .A1(\RI5[4][126] ), .A2(n214), .Z(
        \MC_ARK_ARC_1_4/temp4[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_16_5  ( .A1(\RI5[4][0] ), .A2(\RI5[4][156] ), .Z(
        \MC_ARK_ARC_1_4/temp3[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_16_5  ( .A1(\RI5[4][60] ), .A2(\RI5[4][36] ), .Z(
        \MC_ARK_ARC_1_4/temp2[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_16_5  ( .A1(\RI5[4][90] ), .A2(\RI5[4][84] ), .Z(
        \MC_ARK_ARC_1_4/temp1[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_16_4  ( .A1(\MC_ARK_ARC_1_4/temp5[91] ), .A2(
        \MC_ARK_ARC_1_4/temp6[91] ), .Z(\MC_ARK_ARC_1_4/buf_output[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_16_4  ( .A1(\MC_ARK_ARC_1_4/temp4[91] ), .A2(
        \MC_ARK_ARC_1_4/temp3[91] ), .Z(\MC_ARK_ARC_1_4/temp6[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_16_4  ( .A1(\RI5[4][127] ), .A2(n137), .Z(
        \MC_ARK_ARC_1_4/temp4[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_16_4  ( .A1(\RI5[4][61] ), .A2(\RI5[4][37] ), .Z(
        \MC_ARK_ARC_1_4/temp2[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_16_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[129] ), 
        .A2(n440), .Z(\MC_ARK_ARC_1_4/temp4[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_16_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[87] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[93] ), .Z(\MC_ARK_ARC_1_4/temp1[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_16_1  ( .A1(\MC_ARK_ARC_1_4/temp5[94] ), .A2(
        \MC_ARK_ARC_1_4/temp6[94] ), .Z(\MC_ARK_ARC_1_4/buf_output[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_16_1  ( .A1(\MC_ARK_ARC_1_4/temp4[94] ), .A2(
        \MC_ARK_ARC_1_4/temp3[94] ), .Z(\MC_ARK_ARC_1_4/temp6[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_16_1  ( .A1(\RI5[4][130] ), .A2(n150), .Z(
        \MC_ARK_ARC_1_4/temp4[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_16_1  ( .A1(\RI5[4][4] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[160] ), .Z(\MC_ARK_ARC_1_4/temp3[94] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_16_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[64] ), 
        .A2(\RI5[4][40] ), .Z(\MC_ARK_ARC_1_4/temp2[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_16_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[94] ), 
        .A2(\RI5[4][88] ), .Z(\MC_ARK_ARC_1_4/temp1[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_16_0  ( .A1(\RI5[4][131] ), .A2(n427), .Z(
        \MC_ARK_ARC_1_4/temp4[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_15_5  ( .A1(\MC_ARK_ARC_1_4/temp5[96] ), .A2(
        \MC_ARK_ARC_1_4/temp6[96] ), .Z(\MC_ARK_ARC_1_4/buf_output[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_15_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[132] ), 
        .A2(n499), .Z(\MC_ARK_ARC_1_4/temp4[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_15_5  ( .A1(\RI5[4][6] ), .A2(\RI5[4][162] ), .Z(
        \MC_ARK_ARC_1_4/temp3[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_15_4  ( .A1(\RI5[4][133] ), .A2(n416), .Z(
        \MC_ARK_ARC_1_4/temp4[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_15_4  ( .A1(\RI5[4][7] ), .A2(\RI5[4][163] ), .Z(
        \MC_ARK_ARC_1_4/temp3[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_15_3  ( .A1(\RI5[4][134] ), .A2(n489), .Z(
        \MC_ARK_ARC_1_4/temp4[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_15_3  ( .A1(\RI5[4][92] ), .A2(\RI5[4][98] ), .Z(
        \MC_ARK_ARC_1_4/temp1[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_15_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[135] ), 
        .A2(n103), .Z(\MC_ARK_ARC_1_4/temp4[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_15_1  ( .A1(\MC_ARK_ARC_1_4/temp3[100] ), .A2(
        \MC_ARK_ARC_1_4/temp4[100] ), .Z(\MC_ARK_ARC_1_4/temp6[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_15_1  ( .A1(\RI5[4][136] ), .A2(n176), .Z(
        \MC_ARK_ARC_1_4/temp4[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_15_1  ( .A1(\RI5[4][10] ), .A2(\RI5[4][166] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_15_1  ( .A1(\RI5[4][70] ), .A2(\RI5[4][46] ), .Z(
        \MC_ARK_ARC_1_4/temp2[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_15_1  ( .A1(\RI5[4][100] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[94] ), .Z(\MC_ARK_ARC_1_4/temp1[100] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_15_0  ( .A1(\SB2_4_9/buf_output[5] ), .A2(n186), 
        .Z(\MC_ARK_ARC_1_4/temp4[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_14_5  ( .A1(\MC_ARK_ARC_1_4/temp5[102] ), .A2(
        \MC_ARK_ARC_1_4/temp6[102] ), .Z(\MC_ARK_ARC_1_4/buf_output[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_14_5  ( .A1(\MC_ARK_ARC_1_4/temp3[102] ), .A2(
        \MC_ARK_ARC_1_4/temp4[102] ), .Z(\MC_ARK_ARC_1_4/temp6[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_14_5  ( .A1(\RI5[4][138] ), .A2(n466), .Z(
        \MC_ARK_ARC_1_4/temp4[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_14_5  ( .A1(\RI5[4][102] ), .A2(\RI5[4][96] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_14_4  ( .A1(\RI5[4][139] ), .A2(n152), .Z(
        \MC_ARK_ARC_1_4/temp4[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_14_4  ( .A1(\RI5[4][13] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[169] ), .Z(\MC_ARK_ARC_1_4/temp3[103] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_14_4  ( .A1(\RI5[4][49] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[73] ), .Z(\MC_ARK_ARC_1_4/temp2[103] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_14_4  ( .A1(\RI5[4][103] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[97] ), .Z(\MC_ARK_ARC_1_4/temp1[103] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_14_3  ( .A1(\MC_ARK_ARC_1_4/temp5[104] ), .A2(
        \MC_ARK_ARC_1_4/temp6[104] ), .Z(\MC_ARK_ARC_1_4/buf_output[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_14_3  ( .A1(\MC_ARK_ARC_1_4/temp3[104] ), .A2(
        \MC_ARK_ARC_1_4/temp4[104] ), .Z(\MC_ARK_ARC_1_4/temp6[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_14_3  ( .A1(\RI5[4][140] ), .A2(n51), .Z(
        \MC_ARK_ARC_1_4/temp4[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_14_3  ( .A1(\RI5[4][14] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[170] ), .Z(\MC_ARK_ARC_1_4/temp3[104] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_14_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[141] ), 
        .A2(n142), .Z(\MC_ARK_ARC_1_4/temp4[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_14_1  ( .A1(\MC_ARK_ARC_1_4/temp2[106] ), .A2(
        \MC_ARK_ARC_1_4/temp1[106] ), .Z(\MC_ARK_ARC_1_4/temp5[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_14_1  ( .A1(\RI5[4][142] ), .A2(n35), .Z(
        \MC_ARK_ARC_1_4/temp4[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_14_1  ( .A1(\RI5[4][16] ), .A2(\RI5[4][172] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_14_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[76] ), 
        .A2(\RI5[4][52] ), .Z(\MC_ARK_ARC_1_4/temp2[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_14_1  ( .A1(\RI5[4][106] ), .A2(\RI5[4][100] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_14_0  ( .A1(\RI5[4][143] ), .A2(n515), .Z(
        \MC_ARK_ARC_1_4/temp4[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_13_5  ( .A1(\RI5[4][144] ), .A2(n431), .Z(
        \MC_ARK_ARC_1_4/temp4[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_13_5  ( .A1(\RI5[4][78] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[54] ), .Z(\MC_ARK_ARC_1_4/temp2[108] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_13_4  ( .A1(\RI5[4][145] ), .A2(n207), .Z(
        \MC_ARK_ARC_1_4/temp4[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_13_4  ( .A1(\RI5[4][79] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[55] ), .Z(\MC_ARK_ARC_1_4/temp2[109] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_13_3  ( .A1(\RI5[4][146] ), .A2(n208), .Z(
        \MC_ARK_ARC_1_4/temp4[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_13_3  ( .A1(\RI5[4][20] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[176] ), .Z(\MC_ARK_ARC_1_4/temp3[110] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_13_2  ( .A1(\SB2_4_9/buf_output[3] ), .A2(n492), 
        .Z(\MC_ARK_ARC_1_4/temp4[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_13_1  ( .A1(\MC_ARK_ARC_1_4/temp1[112] ), .A2(
        \MC_ARK_ARC_1_4/temp2[112] ), .Z(\MC_ARK_ARC_1_4/temp5[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_13_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[148] ), 
        .A2(n564), .Z(\MC_ARK_ARC_1_4/temp4[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_13_1  ( .A1(\RI5[4][82] ), .A2(\RI5[4][58] ), .Z(
        \MC_ARK_ARC_1_4/temp2[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_13_1  ( .A1(\RI5[4][112] ), .A2(\RI5[4][106] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_12_5  ( .A1(\RI5[4][150] ), .A2(n215), .Z(
        \MC_ARK_ARC_1_4/temp4[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_12_5  ( .A1(\SB2_4_6/buf_output[0] ), .A2(
        \RI5[4][24] ), .Z(\MC_ARK_ARC_1_4/temp3[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_12_4  ( .A1(\RI5[4][151] ), .A2(n147), .Z(
        \MC_ARK_ARC_1_4/temp4[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_12_4  ( .A1(\RI5[4][25] ), .A2(\RI5[4][181] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_12_3  ( .A1(\RI5[4][152] ), .A2(n201), .Z(
        \MC_ARK_ARC_1_4/temp4[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_12_2  ( .A1(\MC_ARK_ARC_1_4/temp3[117] ), .A2(
        \MC_ARK_ARC_1_4/temp4[117] ), .Z(\MC_ARK_ARC_1_4/temp6[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_12_2  ( .A1(\RI5[4][153] ), .A2(n458), .Z(
        \MC_ARK_ARC_1_4/temp4[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_12_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[183] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[27] ), .Z(
        \MC_ARK_ARC_1_4/temp3[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_12_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[117] ), 
        .A2(\RI5[4][111] ), .Z(\MC_ARK_ARC_1_4/temp1[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_12_1  ( .A1(\MC_ARK_ARC_1_4/temp3[118] ), .A2(
        \MC_ARK_ARC_1_4/temp4[118] ), .Z(\MC_ARK_ARC_1_4/temp6[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_12_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[154] ), 
        .A2(n185), .Z(\MC_ARK_ARC_1_4/temp4[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_12_1  ( .A1(\RI5[4][28] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[184] ), .Z(\MC_ARK_ARC_1_4/temp3[118] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_12_0  ( .A1(\RI5[4][155] ), .A2(n449), .Z(
        \MC_ARK_ARC_1_4/temp4[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_12_0  ( .A1(\RI5[4][185] ), .A2(\RI5[4][29] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_12_0  ( .A1(\RI5[4][65] ), .A2(\RI5[4][89] ), .Z(
        \MC_ARK_ARC_1_4/temp2[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_11_5  ( .A1(\RI5[4][156] ), .A2(n48), .Z(
        \MC_ARK_ARC_1_4/temp4[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_11_5  ( .A1(\RI5[4][30] ), .A2(\RI5[4][186] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_11_5  ( .A1(\RI5[4][66] ), .A2(\RI5[4][90] ), .Z(
        \MC_ARK_ARC_1_4/temp2[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_11_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[120] ), 
        .A2(\RI5[4][114] ), .Z(\MC_ARK_ARC_1_4/temp1[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_11_4  ( .A1(\MC_ARK_ARC_1_4/temp6[121] ), .A2(
        \MC_ARK_ARC_1_4/temp5[121] ), .Z(\MC_ARK_ARC_1_4/buf_output[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_11_4  ( .A1(\MC_ARK_ARC_1_4/temp3[121] ), .A2(
        \MC_ARK_ARC_1_4/temp4[121] ), .Z(\MC_ARK_ARC_1_4/temp6[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_11_4  ( .A1(\MC_ARK_ARC_1_4/temp2[121] ), .A2(
        \MC_ARK_ARC_1_4/temp1[121] ), .Z(\MC_ARK_ARC_1_4/temp5[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_11_4  ( .A1(\RI5[4][157] ), .A2(n183), .Z(
        \MC_ARK_ARC_1_4/temp4[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_11_4  ( .A1(\RI5[4][187] ), .A2(\RI5[4][31] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_11_4  ( .A1(\RI5[4][67] ), .A2(\RI5[4][91] ), .Z(
        \MC_ARK_ARC_1_4/temp2[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_11_4  ( .A1(\RI5[4][121] ), .A2(\RI5[4][115] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_11_3  ( .A1(\RI5[4][158] ), .A2(n507), .Z(
        \MC_ARK_ARC_1_4/temp4[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_11_2  ( .A1(\RI5[4][159] ), .A2(n124), .Z(
        \MC_ARK_ARC_1_4/temp4[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_11_2  ( .A1(\RI5[4][69] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[93] ), .Z(\MC_ARK_ARC_1_4/temp2[123] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_11_1  ( .A1(\MC_ARK_ARC_1_4/temp1[124] ), .A2(
        \MC_ARK_ARC_1_4/temp2[124] ), .Z(\MC_ARK_ARC_1_4/temp5[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_11_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[94] ), 
        .A2(\RI5[4][70] ), .Z(\MC_ARK_ARC_1_4/temp2[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_11_1  ( .A1(\RI5[4][124] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[118] ), .Z(\MC_ARK_ARC_1_4/temp1[124] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_11_0  ( .A1(\RI5[4][161] ), .A2(n569), .Z(
        \MC_ARK_ARC_1_4/temp4[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_11_0  ( .A1(\RI5[4][35] ), .A2(\RI5[4][191] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_10_5  ( .A1(\MC_ARK_ARC_1_4/temp2[126] ), .A2(
        \MC_ARK_ARC_1_4/temp1[126] ), .Z(\MC_ARK_ARC_1_4/temp5[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_10_5  ( .A1(\RI5[4][162] ), .A2(
        \MC_ARK_ARC_1_1/buf_keyinput[111] ), .Z(\MC_ARK_ARC_1_4/temp4[126] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_10_5  ( .A1(\RI5[4][36] ), .A2(\RI5[4][0] ), .Z(
        \MC_ARK_ARC_1_4/temp3[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_10_5  ( .A1(\RI5[4][96] ), .A2(\RI5[4][72] ), .Z(
        \MC_ARK_ARC_1_4/temp2[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_10_5  ( .A1(\RI5[4][126] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[120] ), .Z(\MC_ARK_ARC_1_4/temp1[126] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_10_4  ( .A1(\RI5[4][163] ), .A2(n31), .Z(
        \MC_ARK_ARC_1_4/temp4[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_10_4  ( .A1(\RI5[4][127] ), .A2(\RI5[4][121] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_10_3  ( .A1(\RI5[4][164] ), .A2(n475), .Z(
        \MC_ARK_ARC_1_4/temp4[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_10_3  ( .A1(\RI5[4][38] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[2] ), .Z(\MC_ARK_ARC_1_4/temp3[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_10_3  ( .A1(\RI5[4][74] ), .A2(\RI5[4][98] ), .Z(
        \MC_ARK_ARC_1_4/temp2[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_10_3  ( .A1(\RI5[4][122] ), .A2(\RI5[4][128] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_10_2  ( .A1(\MC_ARK_ARC_1_4/temp4[129] ), .A2(
        \MC_ARK_ARC_1_4/temp3[129] ), .Z(\MC_ARK_ARC_1_4/temp6[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_10_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[165] ), 
        .A2(n220), .Z(\MC_ARK_ARC_1_4/temp4[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_10_1  ( .A1(\RI5[4][166] ), .A2(n70), .Z(
        \MC_ARK_ARC_1_4/temp4[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_10_1  ( .A1(\RI5[4][40] ), .A2(\RI5[4][4] ), .Z(
        \MC_ARK_ARC_1_4/temp3[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_10_1  ( .A1(\RI5[4][100] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_4/temp2[130] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_10_0  ( .A1(\MC_ARK_ARC_1_4/temp6[131] ), .A2(
        \MC_ARK_ARC_1_4/temp5[131] ), .Z(\MC_ARK_ARC_1_4/buf_output[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_10_0  ( .A1(\MC_ARK_ARC_1_4/temp3[131] ), .A2(
        \MC_ARK_ARC_1_4/temp4[131] ), .Z(\MC_ARK_ARC_1_4/temp6[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_10_0  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[167] ), 
        .A2(n536), .Z(\MC_ARK_ARC_1_4/temp4[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_10_0  ( .A1(\RI5[4][5] ), .A2(\RI5[4][41] ), .Z(
        \MC_ARK_ARC_1_4/temp3[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_9_5  ( .A1(\MC_ARK_ARC_1_4/temp6[132] ), .A2(
        \MC_ARK_ARC_1_4/temp5[132] ), .Z(\MC_ARK_ARC_1_4/buf_output[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_9_5  ( .A1(\MC_ARK_ARC_1_4/temp3[132] ), .A2(
        \MC_ARK_ARC_1_4/temp4[132] ), .Z(\MC_ARK_ARC_1_4/temp6[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_9_5  ( .A1(\MC_ARK_ARC_1_4/temp2[132] ), .A2(
        \MC_ARK_ARC_1_4/temp1[132] ), .Z(\MC_ARK_ARC_1_4/temp5[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_9_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[168] ), 
        .A2(n452), .Z(\MC_ARK_ARC_1_4/temp4[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_9_5  ( .A1(\RI5[4][42] ), .A2(\RI5[4][6] ), .Z(
        \MC_ARK_ARC_1_4/temp3[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_9_5  ( .A1(\RI5[4][102] ), .A2(\RI5[4][78] ), .Z(
        \MC_ARK_ARC_1_4/temp2[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_9_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[132] ), 
        .A2(\RI5[4][126] ), .Z(\MC_ARK_ARC_1_4/temp1[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_9_4  ( .A1(\MC_ARK_ARC_1_4/temp3[133] ), .A2(
        \MC_ARK_ARC_1_4/temp4[133] ), .Z(\MC_ARK_ARC_1_4/temp6[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_9_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[169] ), 
        .A2(n154), .Z(\MC_ARK_ARC_1_4/temp4[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_9_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[43] ), 
        .A2(\RI5[4][7] ), .Z(\MC_ARK_ARC_1_4/temp3[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_9_4  ( .A1(\RI5[4][127] ), .A2(\RI5[4][133] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_9_3  ( .A1(\MC_ARK_ARC_1_4/temp3[134] ), .A2(
        \MC_ARK_ARC_1_4/temp4[134] ), .Z(\MC_ARK_ARC_1_4/temp6[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_9_3  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[170] ), 
        .A2(n172), .Z(\MC_ARK_ARC_1_4/temp4[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_9_3  ( .A1(\RI5[4][44] ), .A2(\RI5[4][8] ), .Z(
        \MC_ARK_ARC_1_4/temp3[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_9_3  ( .A1(\RI5[4][80] ), .A2(\RI5[4][104] ), .Z(
        \MC_ARK_ARC_1_4/temp2[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_9_2  ( .A1(\MC_ARK_ARC_1_4/temp5[135] ), .A2(
        \MC_ARK_ARC_1_4/temp6[135] ), .Z(\MC_ARK_ARC_1_4/buf_output[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_9_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[171] ), 
        .A2(n511), .Z(\MC_ARK_ARC_1_4/temp4[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_9_2  ( .A1(\RI5[4][105] ), .A2(\RI5[4][81] ), .Z(
        \MC_ARK_ARC_1_4/temp2[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_9_1  ( .A1(\MC_ARK_ARC_1_4/temp6[136] ), .A2(
        \MC_ARK_ARC_1_4/temp5[136] ), .Z(\MC_ARK_ARC_1_4/buf_output[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_9_1  ( .A1(\MC_ARK_ARC_1_4/temp3[136] ), .A2(
        \MC_ARK_ARC_1_4/temp4[136] ), .Z(\MC_ARK_ARC_1_4/temp6[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_9_1  ( .A1(\MC_ARK_ARC_1_4/temp2[136] ), .A2(
        \MC_ARK_ARC_1_4/temp1[136] ), .Z(\MC_ARK_ARC_1_4/temp5[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_9_1  ( .A1(\RI5[4][172] ), .A2(n428), .Z(
        \MC_ARK_ARC_1_4/temp4[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_9_1  ( .A1(\RI5[4][82] ), .A2(\RI5[4][106] ), .Z(
        \MC_ARK_ARC_1_4/temp2[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_9_1  ( .A1(\RI5[4][136] ), .A2(\RI5[4][130] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_9_0  ( .A1(\MC_ARK_ARC_1_4/temp1[137] ), .A2(
        \MC_ARK_ARC_1_4/temp2[137] ), .Z(\MC_ARK_ARC_1_4/temp5[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_9_0  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[173] ), 
        .A2(n500), .Z(\MC_ARK_ARC_1_4/temp4[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_9_0  ( .A1(\RI5[4][11] ), .A2(\RI5[4][47] ), .Z(
        \MC_ARK_ARC_1_4/temp3[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_9_0  ( .A1(\RI5[4][107] ), .A2(\RI5[4][83] ), .Z(
        \MC_ARK_ARC_1_4/temp2[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_8_5  ( .A1(\MC_ARK_ARC_1_4/temp1[138] ), .A2(
        \MC_ARK_ARC_1_4/temp2[138] ), .Z(\MC_ARK_ARC_1_4/temp5[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_8_5  ( .A1(\RI5[4][174] ), .A2(n417), .Z(
        \MC_ARK_ARC_1_4/temp4[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_8_5  ( .A1(\RI5[4][48] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[12] ), .Z(\MC_ARK_ARC_1_4/temp3[138] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_8_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[108] ), 
        .A2(\RI5[4][84] ), .Z(\MC_ARK_ARC_1_4/temp2[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_8_5  ( .A1(\RI5[4][138] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[132] ), .Z(\MC_ARK_ARC_1_4/temp1[138] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_8_4  ( .A1(n3165), .A2(n490), .Z(
        \MC_ARK_ARC_1_4/temp4[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_8_4  ( .A1(\RI5[4][139] ), .A2(\RI5[4][133] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_8_3  ( .A1(\MC_ARK_ARC_1_4/temp6[140] ), .A2(
        \MC_ARK_ARC_1_4/temp5[140] ), .Z(\MC_ARK_ARC_1_4/buf_output[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_8_3  ( .A1(\MC_ARK_ARC_1_4/temp3[140] ), .A2(
        \MC_ARK_ARC_1_4/temp4[140] ), .Z(\MC_ARK_ARC_1_4/temp6[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_8_3  ( .A1(\MC_ARK_ARC_1_4/temp2[140] ), .A2(
        \MC_ARK_ARC_1_4/temp1[140] ), .Z(\MC_ARK_ARC_1_4/temp5[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_8_3  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[176] ), 
        .A2(n561), .Z(\MC_ARK_ARC_1_4/temp4[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_8_3  ( .A1(\RI5[4][14] ), .A2(\RI5[4][50] ), .Z(
        \MC_ARK_ARC_1_4/temp3[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_8_3  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[86] ), 
        .A2(\RI5[4][110] ), .Z(\MC_ARK_ARC_1_4/temp2[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_8_3  ( .A1(\RI5[4][140] ), .A2(\RI5[4][134] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_8_2  ( .A1(\MC_ARK_ARC_1_4/temp6[141] ), .A2(
        \MC_ARK_ARC_1_4/temp5[141] ), .Z(\MC_ARK_ARC_1_4/buf_output[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_8_2  ( .A1(\MC_ARK_ARC_1_4/temp3[141] ), .A2(
        \MC_ARK_ARC_1_4/temp4[141] ), .Z(\MC_ARK_ARC_1_4/temp6[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_8_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[177] ), 
        .A2(n480), .Z(\MC_ARK_ARC_1_4/temp4[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_8_2  ( .A1(\RI5[4][51] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[15] ), .Z(\MC_ARK_ARC_1_4/temp3[141] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_8_2  ( .A1(\RI5[4][111] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[87] ), .Z(\MC_ARK_ARC_1_4/temp2[141] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_8_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[141] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[135] ), .Z(
        \MC_ARK_ARC_1_4/temp1[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_8_1  ( .A1(\MC_ARK_ARC_1_4/temp5[142] ), .A2(
        \MC_ARK_ARC_1_4/temp6[142] ), .Z(\MC_ARK_ARC_1_4/buf_output[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_8_1  ( .A1(\MC_ARK_ARC_1_4/temp3[142] ), .A2(
        \MC_ARK_ARC_1_4/temp4[142] ), .Z(\MC_ARK_ARC_1_4/temp6[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_8_1  ( .A1(\MC_ARK_ARC_1_4/temp2[142] ), .A2(
        \MC_ARK_ARC_1_4/temp1[142] ), .Z(\MC_ARK_ARC_1_4/temp5[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_8_1  ( .A1(\RI5[4][178] ), .A2(n550), .Z(
        \MC_ARK_ARC_1_4/temp4[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_8_1  ( .A1(\RI5[4][112] ), .A2(\RI5[4][88] ), .Z(
        \MC_ARK_ARC_1_4/temp2[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_8_0  ( .A1(\MC_ARK_ARC_1_4/temp6[143] ), .A2(
        \MC_ARK_ARC_1_4/temp5[143] ), .Z(\MC_ARK_ARC_1_4/buf_output[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_8_0  ( .A1(\MC_ARK_ARC_1_4/temp3[143] ), .A2(
        \MC_ARK_ARC_1_4/temp4[143] ), .Z(\MC_ARK_ARC_1_4/temp6[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_8_0  ( .A1(\MC_ARK_ARC_1_4/temp1[143] ), .A2(
        \MC_ARK_ARC_1_4/temp2[143] ), .Z(\MC_ARK_ARC_1_4/temp5[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_8_0  ( .A1(\RI5[4][179] ), .A2(n139), .Z(
        \MC_ARK_ARC_1_4/temp4[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_8_0  ( .A1(\RI5[4][17] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[53] ), .Z(\MC_ARK_ARC_1_4/temp3[143] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_8_0  ( .A1(\RI5[4][113] ), .A2(\RI5[4][89] ), .Z(
        \MC_ARK_ARC_1_4/temp2[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_8_0  ( .A1(\RI5[4][137] ), .A2(\RI5[4][143] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_7_5  ( .A1(\MC_ARK_ARC_1_4/temp5[144] ), .A2(
        \MC_ARK_ARC_1_4/temp6[144] ), .Z(\MC_ARK_ARC_1_4/buf_output[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_7_5  ( .A1(\MC_ARK_ARC_1_4/temp3[144] ), .A2(
        \MC_ARK_ARC_1_4/temp4[144] ), .Z(\MC_ARK_ARC_1_4/temp6[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_7_5  ( .A1(\MC_ARK_ARC_1_4/temp1[144] ), .A2(
        \MC_ARK_ARC_1_4/temp2[144] ), .Z(\MC_ARK_ARC_1_4/temp5[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_7_5  ( .A1(\RI5[4][180] ), .A2(n107), .Z(
        \MC_ARK_ARC_1_4/temp4[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_7_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[18] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[54] ), .Z(
        \MC_ARK_ARC_1_4/temp3[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_7_5  ( .A1(\RI5[4][114] ), .A2(\RI5[4][90] ), .Z(
        \MC_ARK_ARC_1_4/temp2[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_7_5  ( .A1(\RI5[4][144] ), .A2(\RI5[4][138] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_7_4  ( .A1(\MC_ARK_ARC_1_4/temp3[145] ), .A2(
        \MC_ARK_ARC_1_4/temp4[145] ), .Z(\MC_ARK_ARC_1_4/temp6[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_7_4  ( .A1(\RI5[4][181] ), .A2(n140), .Z(
        \MC_ARK_ARC_1_4/temp4[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_7_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[55] ), 
        .A2(\RI5[4][19] ), .Z(\MC_ARK_ARC_1_4/temp3[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_7_4  ( .A1(\RI5[4][115] ), .A2(\RI5[4][91] ), .Z(
        \MC_ARK_ARC_1_4/temp2[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_7_4  ( .A1(\RI5[4][139] ), .A2(\RI5[4][145] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_7_3  ( .A1(\MC_ARK_ARC_1_4/temp3[146] ), .A2(
        \MC_ARK_ARC_1_4/temp4[146] ), .Z(\MC_ARK_ARC_1_4/temp6[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_7_3  ( .A1(\RI5[4][182] ), .A2(n528), .Z(
        \MC_ARK_ARC_1_4/temp4[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_7_2  ( .A1(\SB2_4_3/buf_output[3] ), .A2(n445), 
        .Z(\MC_ARK_ARC_1_4/temp4[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_7_2  ( .A1(\RI5[4][147] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_4/temp1[147] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_7_1  ( .A1(\MC_ARK_ARC_1_4/temp6[148] ), .A2(
        \MC_ARK_ARC_1_4/temp5[148] ), .Z(\MC_ARK_ARC_1_4/buf_output[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_7_1  ( .A1(\MC_ARK_ARC_1_4/temp3[148] ), .A2(
        \MC_ARK_ARC_1_4/temp4[148] ), .Z(\MC_ARK_ARC_1_4/temp6[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_7_1  ( .A1(\MC_ARK_ARC_1_4/temp2[148] ), .A2(
        \MC_ARK_ARC_1_4/temp1[148] ), .Z(\MC_ARK_ARC_1_4/temp5[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_7_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[184] ), 
        .A2(n194), .Z(\MC_ARK_ARC_1_4/temp4[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_7_1  ( .A1(\RI5[4][58] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_4/temp3[148] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_7_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[148] ), 
        .A2(\RI5[4][142] ), .Z(\MC_ARK_ARC_1_4/temp1[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_7_0  ( .A1(\RI5[4][185] ), .A2(n432), .Z(
        \MC_ARK_ARC_1_4/temp4[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_6_5  ( .A1(\RI5[4][186] ), .A2(n190), .Z(
        \MC_ARK_ARC_1_4/temp4[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_6_5  ( .A1(\RI5[4][60] ), .A2(\RI5[4][24] ), .Z(
        \MC_ARK_ARC_1_4/temp3[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_6_5  ( .A1(\RI5[4][150] ), .A2(\RI5[4][144] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_6_4  ( .A1(\RI5[4][187] ), .A2(n59), .Z(
        \MC_ARK_ARC_1_4/temp4[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_6_4  ( .A1(\RI5[4][61] ), .A2(\RI5[4][25] ), .Z(
        \MC_ARK_ARC_1_4/temp3[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_6_4  ( .A1(\RI5[4][121] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[97] ), .Z(\MC_ARK_ARC_1_4/temp2[151] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_6_4  ( .A1(\RI5[4][151] ), .A2(\RI5[4][145] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_6_3  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[188] ), 
        .A2(n493), .Z(\MC_ARK_ARC_1_4/temp4[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_6_2  ( .A1(\RI5[4][189] ), .A2(n173), .Z(
        \MC_ARK_ARC_1_4/temp4[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_6_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[63] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[27] ), .Z(
        \MC_ARK_ARC_1_4/temp3[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_6_2  ( .A1(\RI5[4][99] ), .A2(\RI5[4][123] ), .Z(
        \MC_ARK_ARC_1_4/temp2[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_6_2  ( .A1(\RI5[4][147] ), .A2(\RI5[4][153] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_6_1  ( .A1(\MC_ARK_ARC_1_4/temp2[154] ), .A2(
        \MC_ARK_ARC_1_4/temp1[154] ), .Z(\MC_ARK_ARC_1_4/temp5[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_6_1  ( .A1(\RI5[4][190] ), .A2(n65), .Z(
        \MC_ARK_ARC_1_4/temp4[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_6_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[154] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[148] ), .Z(
        \MC_ARK_ARC_1_4/temp1[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_6_0  ( .A1(\RI5[4][191] ), .A2(n56), .Z(
        \MC_ARK_ARC_1_4/temp4[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_5_5  ( .A1(\MC_ARK_ARC_1_4/temp3[156] ), .A2(
        \MC_ARK_ARC_1_4/temp4[156] ), .Z(\MC_ARK_ARC_1_4/temp6[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_5_5  ( .A1(\MC_ARK_ARC_1_4/temp2[156] ), .A2(
        \MC_ARK_ARC_1_4/temp1[156] ), .Z(\MC_ARK_ARC_1_4/temp5[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_5_5  ( .A1(\RI5[4][0] ), .A2(n471), .Z(
        \MC_ARK_ARC_1_4/temp4[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_5_5  ( .A1(\RI5[4][30] ), .A2(\RI5[4][66] ), .Z(
        \MC_ARK_ARC_1_4/temp3[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_5_5  ( .A1(\RI5[4][126] ), .A2(\RI5[4][102] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_5_5  ( .A1(\RI5[4][156] ), .A2(\RI5[4][150] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_5_4  ( .A1(\MC_ARK_ARC_1_4/temp5[157] ), .A2(
        \MC_ARK_ARC_1_4/temp6[157] ), .Z(\MC_ARK_ARC_1_4/buf_output[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_5_4  ( .A1(\MC_ARK_ARC_1_4/temp3[157] ), .A2(
        \MC_ARK_ARC_1_4/temp4[157] ), .Z(\MC_ARK_ARC_1_4/temp6[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_5_4  ( .A1(\MC_ARK_ARC_1_4/temp2[157] ), .A2(
        \MC_ARK_ARC_1_4/temp1[157] ), .Z(\MC_ARK_ARC_1_4/temp5[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_5_4  ( .A1(\RI5[4][1] ), .A2(n542), .Z(
        \MC_ARK_ARC_1_4/temp4[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_5_4  ( .A1(\RI5[4][67] ), .A2(\RI5[4][31] ), .Z(
        \MC_ARK_ARC_1_4/temp3[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_5_4  ( .A1(\RI5[4][127] ), .A2(\RI5[4][103] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_5_4  ( .A1(\RI5[4][157] ), .A2(\RI5[4][151] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_5_3  ( .A1(\MC_ARK_ARC_1_4/temp1[158] ), .A2(
        \MC_ARK_ARC_1_4/temp2[158] ), .Z(\MC_ARK_ARC_1_4/temp5[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_5_3  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[2] ), 
        .A2(n459), .Z(\MC_ARK_ARC_1_4/temp4[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_5_3  ( .A1(\RI5[4][128] ), .A2(\RI5[4][104] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_5_3  ( .A1(\RI5[4][152] ), .A2(\RI5[4][158] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_5_2  ( .A1(\MC_ARK_ARC_1_4/temp1[159] ), .A2(
        \MC_ARK_ARC_1_4/temp2[159] ), .Z(\MC_ARK_ARC_1_4/temp5[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_5_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[3] ), 
        .A2(n533), .Z(\MC_ARK_ARC_1_4/temp4[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_5_2  ( .A1(\RI5[4][105] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[129] ), .Z(\MC_ARK_ARC_1_4/temp2[159] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_5_2  ( .A1(\RI5[4][159] ), .A2(\RI5[4][153] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_5_1  ( .A1(\MC_ARK_ARC_1_4/temp1[160] ), .A2(
        \MC_ARK_ARC_1_4/temp2[160] ), .Z(\MC_ARK_ARC_1_4/temp5[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_5_1  ( .A1(\RI5[4][4] ), .A2(n450), .Z(
        \MC_ARK_ARC_1_4/temp4[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_5_1  ( .A1(\RI5[4][70] ), .A2(\RI5[4][34] ), .Z(
        \MC_ARK_ARC_1_4/temp3[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_5_1  ( .A1(\RI5[4][130] ), .A2(\RI5[4][106] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_5_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[160] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[154] ), .Z(
        \MC_ARK_ARC_1_4/temp1[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_5_0  ( .A1(\MC_ARK_ARC_1_4/temp3[161] ), .A2(
        \MC_ARK_ARC_1_4/temp4[161] ), .Z(\MC_ARK_ARC_1_4/temp6[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_5_0  ( .A1(\RI5[4][5] ), .A2(n79), .Z(
        \MC_ARK_ARC_1_4/temp4[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_5_0  ( .A1(\RI5[4][107] ), .A2(\RI5[4][131] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_5_0  ( .A1(\RI5[4][161] ), .A2(\RI5[4][155] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_4_5  ( .A1(\MC_ARK_ARC_1_4/temp5[162] ), .A2(
        \MC_ARK_ARC_1_4/temp6[162] ), .Z(\MC_ARK_ARC_1_4/buf_output[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_4_5  ( .A1(\MC_ARK_ARC_1_4/temp3[162] ), .A2(
        \MC_ARK_ARC_1_4/temp4[162] ), .Z(\MC_ARK_ARC_1_4/temp6[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_4_5  ( .A1(\MC_ARK_ARC_1_4/temp1[162] ), .A2(
        \MC_ARK_ARC_1_4/temp2[162] ), .Z(\MC_ARK_ARC_1_4/temp5[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_4_5  ( .A1(\RI5[4][6] ), .A2(n437), .Z(
        \MC_ARK_ARC_1_4/temp4[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_4_5  ( .A1(\RI5[4][72] ), .A2(\RI5[4][36] ), .Z(
        \MC_ARK_ARC_1_4/temp3[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_4_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[132] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[108] ), .Z(
        \MC_ARK_ARC_1_4/temp2[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_4_5  ( .A1(\RI5[4][162] ), .A2(\RI5[4][156] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_4_4  ( .A1(\RI5[4][7] ), .A2(n202), .Z(
        \MC_ARK_ARC_1_4/temp4[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_4_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[73] ), 
        .A2(\RI5[4][37] ), .Z(\MC_ARK_ARC_1_4/temp3[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_4_4  ( .A1(\RI5[4][157] ), .A2(\RI5[4][163] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_4_3  ( .A1(\MC_ARK_ARC_1_4/temp6[164] ), .A2(
        \MC_ARK_ARC_1_4/temp5[164] ), .Z(\MC_ARK_ARC_1_4/buf_output[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_4_3  ( .A1(\MC_ARK_ARC_1_4/temp4[164] ), .A2(
        \MC_ARK_ARC_1_4/temp3[164] ), .Z(\MC_ARK_ARC_1_4/temp6[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_4_3  ( .A1(\RI5[4][8] ), .A2(n180), .Z(
        \MC_ARK_ARC_1_4/temp4[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_4_3  ( .A1(\RI5[4][38] ), .A2(\RI5[4][74] ), .Z(
        \MC_ARK_ARC_1_4/temp3[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_4_2  ( .A1(\MC_ARK_ARC_1_4/temp3[165] ), .A2(
        \MC_ARK_ARC_1_4/temp4[165] ), .Z(\MC_ARK_ARC_1_4/temp6[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_4_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[9] ), 
        .A2(n218), .Z(\MC_ARK_ARC_1_4/temp4[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_4_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[135] ), 
        .A2(\RI5[4][111] ), .Z(\MC_ARK_ARC_1_4/temp2[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_4_2  ( .A1(\RI5[4][159] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[165] ), .Z(\MC_ARK_ARC_1_4/temp1[165] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_4_1  ( .A1(\MC_ARK_ARC_1_4/temp3[166] ), .A2(
        \MC_ARK_ARC_1_4/temp4[166] ), .Z(\MC_ARK_ARC_1_4/temp6[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_4_1  ( .A1(\RI5[4][10] ), .A2(n413), .Z(
        \MC_ARK_ARC_1_4/temp4[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_4_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[76] ), 
        .A2(\RI5[4][40] ), .Z(\MC_ARK_ARC_1_4/temp3[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_4_1  ( .A1(\SB2_4_10/buf_output[4] ), .A2(
        \RI5[4][112] ), .Z(\MC_ARK_ARC_1_4/temp2[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_4_1  ( .A1(\RI5[4][166] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[160] ), .Z(\MC_ARK_ARC_1_4/temp1[166] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_4_0  ( .A1(\MC_ARK_ARC_1_4/temp3[167] ), .A2(
        \MC_ARK_ARC_1_4/temp4[167] ), .Z(\MC_ARK_ARC_1_4/temp6[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_4_0  ( .A1(\MC_ARK_ARC_1_4/temp2[167] ), .A2(
        \MC_ARK_ARC_1_4/temp1[167] ), .Z(\MC_ARK_ARC_1_4/temp5[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_4_0  ( .A1(\RI5[4][11] ), .A2(n54), .Z(
        \MC_ARK_ARC_1_4/temp4[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_4_0  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[77] ), 
        .A2(\RI5[4][41] ), .Z(\MC_ARK_ARC_1_4/temp3[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_4_0  ( .A1(\RI5[4][137] ), .A2(\RI5[4][113] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_4_0  ( .A1(\RI5[4][161] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[167] ), .Z(\MC_ARK_ARC_1_4/temp1[167] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_3_5  ( .A1(\MC_ARK_ARC_1_4/temp6[168] ), .A2(
        \MC_ARK_ARC_1_4/temp5[168] ), .Z(\MC_ARK_ARC_1_4/buf_output[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_3_5  ( .A1(\MC_ARK_ARC_1_4/temp1[168] ), .A2(
        \MC_ARK_ARC_1_4/temp2[168] ), .Z(\MC_ARK_ARC_1_4/temp5[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_3_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[12] ), 
        .A2(n24), .Z(\MC_ARK_ARC_1_4/temp4[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_3_5  ( .A1(\RI5[4][138] ), .A2(\RI5[4][114] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_3_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[168] ), 
        .A2(\RI5[4][162] ), .Z(\MC_ARK_ARC_1_4/temp1[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_3_4  ( .A1(\MC_ARK_ARC_1_4/temp6[169] ), .A2(
        \MC_ARK_ARC_1_4/temp5[169] ), .Z(\MC_ARK_ARC_1_4/buf_output[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_3_4  ( .A1(\MC_ARK_ARC_1_4/temp3[169] ), .A2(
        \MC_ARK_ARC_1_4/temp4[169] ), .Z(\MC_ARK_ARC_1_4/temp6[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_3_4  ( .A1(\MC_ARK_ARC_1_4/temp1[169] ), .A2(
        \MC_ARK_ARC_1_4/temp2[169] ), .Z(\MC_ARK_ARC_1_4/temp5[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_3_4  ( .A1(\RI5[4][13] ), .A2(n205), .Z(
        \MC_ARK_ARC_1_4/temp4[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_3_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[43] ), 
        .A2(\RI5[4][79] ), .Z(\MC_ARK_ARC_1_4/temp3[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_3_4  ( .A1(\RI5[4][139] ), .A2(\RI5[4][115] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_3_4  ( .A1(\RI5[4][163] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[169] ), .Z(\MC_ARK_ARC_1_4/temp1[169] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_3_3  ( .A1(\RI5[4][14] ), .A2(n66), .Z(
        \MC_ARK_ARC_1_4/temp4[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_3_2  ( .A1(\MC_ARK_ARC_1_4/temp2[171] ), .A2(
        \MC_ARK_ARC_1_4/temp1[171] ), .Z(\MC_ARK_ARC_1_4/temp5[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_3_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[15] ), 
        .A2(n134), .Z(\MC_ARK_ARC_1_4/temp4[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_3_2  ( .A1(\RI5[4][81] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[45] ), .Z(\MC_ARK_ARC_1_4/temp3[171] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_3_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[165] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[171] ), .Z(
        \MC_ARK_ARC_1_4/temp1[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_3_1  ( .A1(\MC_ARK_ARC_1_4/temp3[172] ), .A2(
        \MC_ARK_ARC_1_4/temp4[172] ), .Z(\MC_ARK_ARC_1_4/temp6[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_3_1  ( .A1(\MC_ARK_ARC_1_4/temp1[172] ), .A2(
        \MC_ARK_ARC_1_4/temp2[172] ), .Z(\MC_ARK_ARC_1_4/temp5[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_3_1  ( .A1(\RI5[4][16] ), .A2(n537), .Z(
        \MC_ARK_ARC_1_4/temp4[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_3_1  ( .A1(\RI5[4][46] ), .A2(\RI5[4][82] ), .Z(
        \MC_ARK_ARC_1_4/temp3[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_3_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[118] ), 
        .A2(\RI5[4][142] ), .Z(\MC_ARK_ARC_1_4/temp2[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_3_1  ( .A1(\RI5[4][172] ), .A2(\RI5[4][166] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_2_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[18] ), 
        .A2(n197), .Z(\MC_ARK_ARC_1_4/temp4[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_2_5  ( .A1(\RI5[4][144] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[120] ), .Z(\MC_ARK_ARC_1_4/temp2[174] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_2_4  ( .A1(\MC_ARK_ARC_1_4/temp3[175] ), .A2(
        \MC_ARK_ARC_1_4/temp4[175] ), .Z(\MC_ARK_ARC_1_4/temp6[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_2_4  ( .A1(\RI5[4][19] ), .A2(n441), .Z(
        \MC_ARK_ARC_1_4/temp4[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_2_4  ( .A1(\RI5[4][85] ), .A2(\RI5[4][49] ), .Z(
        \MC_ARK_ARC_1_4/temp3[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_2_4  ( .A1(\RI5[4][145] ), .A2(\RI5[4][121] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_2_4  ( .A1(n3166), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[169] ), .Z(\MC_ARK_ARC_1_4/temp1[175] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_2_3  ( .A1(\MC_ARK_ARC_1_4/temp3[176] ), .A2(
        \MC_ARK_ARC_1_4/temp4[176] ), .Z(\MC_ARK_ARC_1_4/temp6[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_2_3  ( .A1(\RI5[4][20] ), .A2(n151), .Z(
        \MC_ARK_ARC_1_4/temp4[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_2_3  ( .A1(\RI5[4][50] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[86] ), .Z(\MC_ARK_ARC_1_4/temp3[176] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_2_3  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[176] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[170] ), .Z(
        \MC_ARK_ARC_1_4/temp1[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_2_2  ( .A1(\RI5[4][21] ), .A2(n184), .Z(
        \MC_ARK_ARC_1_4/temp4[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_2_2  ( .A1(\RI5[4][51] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[87] ), .Z(\MC_ARK_ARC_1_4/temp3[177] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_2_2  ( .A1(\RI5[4][147] ), .A2(\RI5[4][123] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_2_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[171] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[177] ), .Z(
        \MC_ARK_ARC_1_4/temp1[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X7_2_1  ( .A1(\MC_ARK_ARC_1_4/temp6[178] ), .A2(
        \MC_ARK_ARC_1_4/temp5[178] ), .Z(\MC_ARK_ARC_1_4/buf_output[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_2_1  ( .A1(\MC_ARK_ARC_1_4/temp3[178] ), .A2(
        \MC_ARK_ARC_1_4/temp4[178] ), .Z(\MC_ARK_ARC_1_4/temp6[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_2_1  ( .A1(\MC_ARK_ARC_1_4/temp1[178] ), .A2(
        \MC_ARK_ARC_1_4/temp2[178] ), .Z(\MC_ARK_ARC_1_4/temp5[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_2_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[22] ), 
        .A2(n501), .Z(\MC_ARK_ARC_1_4/temp4[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_2_1  ( .A1(\RI5[4][88] ), .A2(\RI5[4][52] ), .Z(
        \MC_ARK_ARC_1_4/temp3[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_2_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[148] ), 
        .A2(\RI5[4][124] ), .Z(\MC_ARK_ARC_1_4/temp2[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_2_1  ( .A1(\RI5[4][178] ), .A2(\RI5[4][172] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_2_0  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[23] ), 
        .A2(n418), .Z(\MC_ARK_ARC_1_4/temp4[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_1_5  ( .A1(\MC_ARK_ARC_1_4/temp1[180] ), .A2(
        \MC_ARK_ARC_1_4/temp2[180] ), .Z(\MC_ARK_ARC_1_4/temp5[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_1_5  ( .A1(\RI5[4][24] ), .A2(n878), .Z(
        \MC_ARK_ARC_1_4/temp4[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_1_5  ( .A1(\RI5[4][90] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[54] ), .Z(\MC_ARK_ARC_1_4/temp3[180] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_1_5  ( .A1(\RI5[4][150] ), .A2(\RI5[4][126] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_1_5  ( .A1(\RI5[4][180] ), .A2(\RI5[4][174] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_1_4  ( .A1(\MC_ARK_ARC_1_4/temp3[181] ), .A2(
        \MC_ARK_ARC_1_4/temp4[181] ), .Z(\MC_ARK_ARC_1_4/temp6[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_1_4  ( .A1(\RI5[4][25] ), .A2(n562), .Z(
        \MC_ARK_ARC_1_4/temp4[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_1_4  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[55] ), 
        .A2(\RI5[4][91] ), .Z(\MC_ARK_ARC_1_4/temp3[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_1_4  ( .A1(\RI5[4][151] ), .A2(\RI5[4][127] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_1_4  ( .A1(n3165), .A2(\RI5[4][181] ), .Z(
        \MC_ARK_ARC_1_4/temp1[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_1_3  ( .A1(\RI5[4][26] ), .A2(n481), .Z(
        \MC_ARK_ARC_1_4/temp4[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_1_3  ( .A1(\RI5[4][56] ), .A2(\RI5[4][92] ), .Z(
        \MC_ARK_ARC_1_4/temp3[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_1_3  ( .A1(\RI5[4][152] ), .A2(\RI5[4][128] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_1_3  ( .A1(\RI5[4][182] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[176] ), .Z(\MC_ARK_ARC_1_4/temp1[182] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_1_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[27] ), 
        .A2(n188), .Z(\MC_ARK_ARC_1_4/temp4[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_1_2  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[177] ), 
        .A2(\MC_ARK_ARC_1_4/buf_datainput[183] ), .Z(
        \MC_ARK_ARC_1_4/temp1[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X5_1_1  ( .A1(\MC_ARK_ARC_1_4/temp1[184] ), .A2(
        \MC_ARK_ARC_1_4/temp2[184] ), .Z(\MC_ARK_ARC_1_4/temp5[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_1_1  ( .A1(\RI5[4][28] ), .A2(n170), .Z(
        \MC_ARK_ARC_1_4/temp4[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_1_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[94] ), 
        .A2(\RI5[4][58] ), .Z(\MC_ARK_ARC_1_4/temp3[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_1_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[154] ), 
        .A2(\RI5[4][130] ), .Z(\MC_ARK_ARC_1_4/temp2[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_1_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[184] ), 
        .A2(\RI5[4][178] ), .Z(\MC_ARK_ARC_1_4/temp1[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_0_5  ( .A1(\RI5[4][30] ), .A2(n100), .Z(
        \MC_ARK_ARC_1_4/temp4[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X3_0_5  ( .A1(\RI5[4][60] ), .A2(\RI5[4][96] ), .Z(
        \MC_ARK_ARC_1_4/temp3[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_0_5  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[132] ), 
        .A2(\RI5[4][156] ), .Z(\MC_ARK_ARC_1_4/temp2[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_0_5  ( .A1(\RI5[4][180] ), .A2(\RI5[4][186] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_0_4  ( .A1(\MC_ARK_ARC_1_4/temp3[187] ), .A2(
        \MC_ARK_ARC_1_4/temp4[187] ), .Z(\MC_ARK_ARC_1_4/temp6[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_0_4  ( .A1(\RI5[4][31] ), .A2(n529), .Z(
        \MC_ARK_ARC_1_4/temp4[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_0_4  ( .A1(\SB2_4_4/buf_output[1] ), .A2(
        \RI5[4][181] ), .Z(\MC_ARK_ARC_1_4/temp1[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_0_3  ( .A1(\SB2_4_29/buf_output[2] ), .A2(n446), 
        .Z(\MC_ARK_ARC_1_4/temp4[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X2_0_3  ( .A1(\RI5[4][158] ), .A2(\RI5[4][134] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_0_2  ( .A1(\RI5[4][33] ), .A2(n517), .Z(
        \MC_ARK_ARC_1_4/temp4[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X6_0_1  ( .A1(\MC_ARK_ARC_1_4/temp3[190] ), .A2(
        \MC_ARK_ARC_1_4/temp4[190] ), .Z(\MC_ARK_ARC_1_4/temp6[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_0_1  ( .A1(\RI5[4][34] ), .A2(
        \MC_ARK_ARC_1_3/buf_keyinput[183] ), .Z(\MC_ARK_ARC_1_4/temp4[190] )
         );
  XOR2_X1 \MC_ARK_ARC_1_4/X1_0_1  ( .A1(\MC_ARK_ARC_1_4/buf_datainput[184] ), 
        .A2(\RI5[4][190] ), .Z(\MC_ARK_ARC_1_4/temp1[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_4/X4_0_0  ( .A1(\RI5[4][35] ), .A2(n505), .Z(
        \MC_ARK_ARC_1_4/temp4[191] ) );
  INV_X1 \SB1_0_0/INV_5  ( .I(n412), .ZN(\SB1_0_0/i1_5 ) );
  INV_X1 \SB1_0_0/INV_4  ( .I(n380), .ZN(\SB1_0_0/i0[7] ) );
  INV_X1 \SB1_0_0/INV_1  ( .I(n252), .ZN(\SB1_0_0/i1_7 ) );
  INV_X1 \SB1_0_0/INV_0  ( .I(n315), .ZN(\SB1_0_0/i3[0] ) );
  INV_X1 \SB1_0_1/INV_4  ( .I(n378), .ZN(\SB1_0_1/i0[7] ) );
  INV_X1 \SB1_0_1/INV_0  ( .I(n313), .ZN(\SB1_0_1/i3[0] ) );
  INV_X1 \SB1_0_2/INV_4  ( .I(n376), .ZN(\SB1_0_2/i0[7] ) );
  INV_X1 \SB1_0_2/INV_1  ( .I(n250), .ZN(\SB1_0_2/i1_7 ) );
  INV_X1 \SB1_0_2/INV_0  ( .I(n311), .ZN(\SB1_0_2/i3[0] ) );
  INV_X1 \SB1_0_3/INV_4  ( .I(n374), .ZN(\SB1_0_3/i0[7] ) );
  INV_X1 \SB1_0_3/INV_1  ( .I(n249), .ZN(\SB1_0_3/i1_7 ) );
  INV_X1 \SB1_0_3/INV_0  ( .I(n309), .ZN(\SB1_0_3/i3[0] ) );
  INV_X1 \SB1_0_4/INV_4  ( .I(n372), .ZN(\SB1_0_4/i0[7] ) );
  INV_X1 \SB1_0_4/INV_1  ( .I(n248), .ZN(\SB1_0_4/i1_7 ) );
  INV_X1 \SB1_0_4/INV_0  ( .I(n307), .ZN(\SB1_0_4/i3[0] ) );
  INV_X1 \SB1_0_5/INV_4  ( .I(n370), .ZN(\SB1_0_5/i0[7] ) );
  INV_X1 \SB1_0_5/INV_0  ( .I(n305), .ZN(\SB1_0_5/i3[0] ) );
  INV_X1 \SB1_0_6/INV_5  ( .I(n406), .ZN(\SB1_0_6/i1_5 ) );
  INV_X1 \SB1_0_6/INV_4  ( .I(n368), .ZN(\SB1_0_6/i0[7] ) );
  INV_X1 \SB1_0_6/INV_1  ( .I(n246), .ZN(\SB1_0_6/i1_7 ) );
  INV_X1 \SB1_0_6/INV_0  ( .I(n303), .ZN(\SB1_0_6/i3[0] ) );
  INV_X1 \SB1_0_7/INV_4  ( .I(n366), .ZN(\SB1_0_7/i0[7] ) );
  INV_X1 \SB1_0_7/INV_1  ( .I(n245), .ZN(\SB1_0_7/i1_7 ) );
  INV_X1 \SB1_0_7/INV_0  ( .I(n301), .ZN(\SB1_0_7/i3[0] ) );
  INV_X1 \SB1_0_8/INV_4  ( .I(n364), .ZN(\SB1_0_8/i0[7] ) );
  INV_X1 \SB1_0_8/INV_1  ( .I(n244), .ZN(\SB1_0_8/i1_7 ) );
  INV_X1 \SB1_0_8/INV_0  ( .I(n299), .ZN(\SB1_0_8/i3[0] ) );
  INV_X1 \SB1_0_9/INV_5  ( .I(n403), .ZN(\SB1_0_9/i1_5 ) );
  INV_X1 \SB1_0_9/INV_4  ( .I(n362), .ZN(\SB1_0_9/i0[7] ) );
  INV_X1 \SB1_0_9/INV_0  ( .I(n297), .ZN(\SB1_0_9/i3[0] ) );
  INV_X1 \SB1_0_10/INV_1  ( .I(n242), .ZN(\SB1_0_10/i1_7 ) );
  INV_X1 \SB1_0_11/INV_4  ( .I(n358), .ZN(\SB1_0_11/i0[7] ) );
  INV_X1 \SB1_0_11/INV_1  ( .I(n241), .ZN(\SB1_0_11/i1_7 ) );
  INV_X1 \SB1_0_11/INV_0  ( .I(n293), .ZN(\SB1_0_11/i3[0] ) );
  INV_X1 \SB1_0_12/INV_4  ( .I(n356), .ZN(\SB1_0_12/i0[7] ) );
  INV_X1 \SB1_0_12/INV_0  ( .I(n291), .ZN(\SB1_0_12/i3[0] ) );
  INV_X1 \SB1_0_13/INV_5  ( .I(n399), .ZN(\SB1_0_13/i1_5 ) );
  INV_X1 \SB1_0_13/INV_1  ( .I(n239), .ZN(\SB1_0_13/i1_7 ) );
  INV_X1 \SB1_0_13/INV_0  ( .I(n289), .ZN(\SB1_0_13/i3[0] ) );
  INV_X1 \SB1_0_14/INV_4  ( .I(n352), .ZN(\SB1_0_14/i0[7] ) );
  INV_X1 \SB1_0_14/INV_0  ( .I(n287), .ZN(\SB1_0_14/i3[0] ) );
  INV_X1 \SB1_0_15/INV_5  ( .I(n397), .ZN(\SB1_0_15/i1_5 ) );
  INV_X1 \SB1_0_15/INV_4  ( .I(n350), .ZN(\SB1_0_15/i0[7] ) );
  INV_X1 \SB1_0_16/INV_4  ( .I(n348), .ZN(\SB1_0_16/i0[7] ) );
  INV_X1 \SB1_0_17/INV_5  ( .I(n395), .ZN(\SB1_0_17/i1_5 ) );
  INV_X1 \SB1_0_17/INV_1  ( .I(n235), .ZN(\SB1_0_17/i1_7 ) );
  INV_X1 \SB1_0_17/INV_0  ( .I(n281), .ZN(\SB1_0_17/i3[0] ) );
  INV_X1 \SB1_0_18/INV_4  ( .I(n344), .ZN(\SB1_0_18/i0[7] ) );
  INV_X1 \SB1_0_18/INV_0  ( .I(n279), .ZN(\SB1_0_18/i3[0] ) );
  INV_X1 \SB1_0_19/INV_1  ( .I(n233), .ZN(\SB1_0_19/i1_7 ) );
  INV_X1 \SB1_0_19/INV_0  ( .I(n277), .ZN(\SB1_0_19/i3[0] ) );
  INV_X1 \SB1_0_21/INV_4  ( .I(n338), .ZN(\SB1_0_21/i0[7] ) );
  INV_X1 \SB1_0_21/INV_1  ( .I(n231), .ZN(\SB1_0_21/i1_7 ) );
  INV_X1 \SB1_0_21/INV_0  ( .I(n273), .ZN(\SB1_0_21/i3[0] ) );
  INV_X1 \SB1_0_22/INV_4  ( .I(n336), .ZN(\SB1_0_22/i0[7] ) );
  INV_X1 \SB1_0_22/INV_1  ( .I(n230), .ZN(\SB1_0_22/i1_7 ) );
  INV_X1 \SB1_0_22/INV_0  ( .I(n271), .ZN(\SB1_0_22/i3[0] ) );
  INV_X1 \SB1_0_23/INV_4  ( .I(n334), .ZN(\SB1_0_23/i0[7] ) );
  INV_X1 \SB1_0_23/INV_0  ( .I(n269), .ZN(\SB1_0_23/i3[0] ) );
  INV_X1 \SB1_0_25/INV_0  ( .I(n265), .ZN(\SB1_0_25/i3[0] ) );
  INV_X1 \SB1_0_26/INV_4  ( .I(n328), .ZN(\SB1_0_26/i0[7] ) );
  INV_X1 \SB1_0_26/INV_1  ( .I(n226), .ZN(\SB1_0_26/i1_7 ) );
  INV_X1 \SB1_0_26/INV_0  ( .I(n263), .ZN(\SB1_0_26/i3[0] ) );
  INV_X1 \SB1_0_27/INV_5  ( .I(n385), .ZN(\SB1_0_27/i1_5 ) );
  INV_X1 \SB1_0_27/INV_1  ( .I(n225), .ZN(\SB1_0_27/i1_7 ) );
  INV_X1 \SB1_0_27/INV_0  ( .I(n261), .ZN(\SB1_0_27/i3[0] ) );
  INV_X1 \SB1_0_28/INV_4  ( .I(n324), .ZN(\SB1_0_28/i0[7] ) );
  INV_X1 \SB1_0_28/INV_1  ( .I(n224), .ZN(\SB1_0_28/i1_7 ) );
  INV_X1 \SB1_0_28/INV_0  ( .I(n259), .ZN(\SB1_0_28/i3[0] ) );
  INV_X1 \SB1_0_29/INV_4  ( .I(n322), .ZN(\SB1_0_29/i0[7] ) );
  INV_X1 \SB1_0_29/INV_1  ( .I(n223), .ZN(\SB1_0_29/i1_7 ) );
  INV_X1 \SB1_0_29/INV_0  ( .I(n257), .ZN(\SB1_0_29/i3[0] ) );
  INV_X1 \SB1_0_30/INV_4  ( .I(n320), .ZN(\SB1_0_30/i0[7] ) );
  INV_X1 \SB1_0_30/INV_0  ( .I(n255), .ZN(\SB1_0_30/i3[0] ) );
  INV_X1 \SB1_0_31/INV_4  ( .I(n318), .ZN(\SB1_0_31/i0[7] ) );
  INV_X1 \SB1_0_31/INV_1  ( .I(n221), .ZN(\SB1_0_31/i1_7 ) );
  INV_X1 \SB1_0_31/INV_0  ( .I(n253), .ZN(\SB1_0_31/i3[0] ) );
  INV_X1 \SB2_0_0/INV_4  ( .I(\SB1_0_1/buf_output[4] ), .ZN(\SB2_0_0/i0[7] )
         );
  INV_X1 \SB2_0_1/INV_4  ( .I(\RI3[0][184] ), .ZN(\SB2_0_1/i0[7] ) );
  INV_X1 \SB2_0_1/INV_1  ( .I(\SB1_0_5/buf_output[1] ), .ZN(\SB2_0_1/i1_7 ) );
  INV_X1 \SB2_0_2/INV_1  ( .I(\RI3[0][175] ), .ZN(\SB2_0_2/i1_7 ) );
  INV_X1 \SB2_0_2/INV_0  ( .I(\RI3[0][174] ), .ZN(\SB2_0_2/i3[0] ) );
  INV_X1 \SB2_0_3/INV_1  ( .I(\RI3[0][169] ), .ZN(\SB2_0_3/i1_7 ) );
  INV_X1 \SB2_0_4/INV_1  ( .I(\RI3[0][163] ), .ZN(\SB2_0_4/i1_7 ) );
  INV_X1 \SB2_0_5/INV_0  ( .I(\SB1_0_10/buf_output[0] ), .ZN(\SB2_0_5/i3[0] )
         );
  INV_X1 \SB2_0_6/INV_4  ( .I(\RI3[0][154] ), .ZN(\SB2_0_6/i0[7] ) );
  INV_X2 \SB2_0_6/INV_3  ( .I(\RI3[0][153] ), .ZN(\SB2_0_6/i0[8] ) );
  INV_X1 \SB2_0_6/INV_0  ( .I(\RI3[0][150] ), .ZN(\SB2_0_6/i3[0] ) );
  INV_X1 \SB2_0_8/INV_0  ( .I(\SB1_0_13/buf_output[0] ), .ZN(\SB2_0_8/i3[0] )
         );
  INV_X1 \SB2_0_9/INV_4  ( .I(\RI3[0][136] ), .ZN(\SB2_0_9/i0[7] ) );
  INV_X1 \SB2_0_11/INV_4  ( .I(\SB1_0_12/buf_output[4] ), .ZN(\SB2_0_11/i0[7] ) );
  INV_X2 \SB2_0_11/INV_3  ( .I(\RI3[0][123] ), .ZN(\SB2_0_11/i0[8] ) );
  INV_X1 \SB2_0_12/INV_0  ( .I(\RI3[0][114] ), .ZN(\SB2_0_12/i3[0] ) );
  INV_X1 \SB2_0_13/INV_4  ( .I(\SB1_0_14/buf_output[4] ), .ZN(\SB2_0_13/i0[7] ) );
  INV_X1 \SB2_0_15/INV_0  ( .I(\RI3[0][96] ), .ZN(\SB2_0_15/i3[0] ) );
  INV_X1 \SB2_0_16/INV_0  ( .I(\RI3[0][90] ), .ZN(\SB2_0_16/i3[0] ) );
  INV_X1 \SB2_0_18/INV_4  ( .I(\SB1_0_19/buf_output[4] ), .ZN(\SB2_0_18/i0[7] ) );
  INV_X1 \SB2_0_19/INV_0  ( .I(\RI3[0][72] ), .ZN(\SB2_0_19/i3[0] ) );
  INV_X1 \SB2_0_20/INV_4  ( .I(\SB1_0_21/buf_output[4] ), .ZN(\SB2_0_20/i0[7] ) );
  INV_X1 \SB2_0_21/INV_4  ( .I(\SB1_0_22/buf_output[4] ), .ZN(\SB2_0_21/i0[7] ) );
  INV_X1 \SB2_0_22/INV_0  ( .I(\SB1_0_27/buf_output[0] ), .ZN(\SB2_0_22/i3[0] ) );
  INV_X2 \SB2_0_23/INV_3  ( .I(\SB1_0_25/buf_output[3] ), .ZN(\SB2_0_23/i0[8] ) );
  INV_X2 \SB2_0_23/INV_2  ( .I(\RI3[0][50] ), .ZN(\SB2_0_23/i1[9] ) );
  INV_X1 \SB2_0_23/INV_0  ( .I(\SB1_0_28/buf_output[0] ), .ZN(\SB2_0_23/i3[0] ) );
  INV_X2 \SB2_0_24/INV_3  ( .I(\SB1_0_26/buf_output[3] ), .ZN(\SB2_0_24/i0[8] ) );
  INV_X1 \SB2_0_24/INV_1  ( .I(\SB1_0_28/buf_output[1] ), .ZN(\SB2_0_24/i1_7 )
         );
  INV_X1 \SB2_0_24/INV_0  ( .I(\SB1_0_29/buf_output[0] ), .ZN(\SB2_0_24/i3[0] ) );
  INV_X1 \SB2_0_25/INV_0  ( .I(\SB1_0_30/buf_output[0] ), .ZN(\SB2_0_25/i3[0] ) );
  INV_X1 \SB2_0_26/INV_0  ( .I(\RI3[0][30] ), .ZN(\SB2_0_26/i3[0] ) );
  INV_X1 \SB2_0_27/INV_1  ( .I(\SB1_0_31/buf_output[1] ), .ZN(\SB2_0_27/i1_7 )
         );
  INV_X1 \SB2_0_28/INV_0  ( .I(\RI3[0][18] ), .ZN(\SB2_0_28/i3[0] ) );
  INV_X2 \SB2_0_29/INV_2  ( .I(\SB1_0_0/buf_output[2] ), .ZN(\SB2_0_29/i1[9] )
         );
  INV_X1 \SB2_0_30/INV_4  ( .I(\RI3[0][10] ), .ZN(\SB2_0_30/i0[7] ) );
  INV_X1 \SB2_0_30/INV_0  ( .I(\SB1_0_3/buf_output[0] ), .ZN(\SB2_0_30/i3[0] )
         );
  INV_X1 \SB2_0_31/INV_0  ( .I(\RI3[0][0] ), .ZN(\SB2_0_31/i3[0] ) );
  INV_X1 \SB1_1_0/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[186] ), .ZN(
        \SB1_1_0/i3[0] ) );
  INV_X1 \SB1_1_1/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[184] ), .ZN(
        \SB1_1_1/i0[7] ) );
  INV_X2 \SB1_1_1/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[182] ), .ZN(
        \SB1_1_1/i1[9] ) );
  INV_X1 \SB1_1_1/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[180] ), .ZN(
        \SB1_1_1/i3[0] ) );
  INV_X1 \SB1_1_2/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[178] ), .ZN(
        \SB1_1_2/i0[7] ) );
  INV_X2 \SB1_1_2/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[177] ), .ZN(
        \SB1_1_2/i0[8] ) );
  INV_X2 \SB1_1_2/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[176] ), .ZN(
        \SB1_1_2/i1[9] ) );
  INV_X1 \SB1_1_2/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[174] ), .ZN(
        \SB1_1_2/i3[0] ) );
  INV_X1 \SB1_1_3/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[172] ), .ZN(
        \SB1_1_3/i0[7] ) );
  INV_X2 \SB1_1_4/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[164] ), .ZN(
        \SB1_1_4/i1[9] ) );
  INV_X1 \SB1_1_5/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[160] ), .ZN(
        \SB1_1_5/i0[7] ) );
  INV_X2 \SB1_1_5/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[159] ), .ZN(
        \SB1_1_5/i0[8] ) );
  INV_X1 \SB1_1_6/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[154] ), .ZN(
        \SB1_1_6/i0[7] ) );
  INV_X2 \SB1_1_6/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[153] ), .ZN(
        \SB1_1_6/i0[8] ) );
  INV_X1 \SB1_1_6/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[151] ), .ZN(
        \SB1_1_6/i1_7 ) );
  INV_X1 \SB1_1_7/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[148] ), .ZN(
        \SB1_1_7/i0[7] ) );
  INV_X1 \SB1_1_7/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[145] ), .ZN(
        \SB1_1_7/i1_7 ) );
  INV_X1 \SB1_1_8/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[139] ), .ZN(
        \SB1_1_8/i1_7 ) );
  INV_X1 \SB1_1_9/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[136] ), .ZN(
        \SB1_1_9/i0[7] ) );
  INV_X2 \SB1_1_9/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[135] ), .ZN(
        \SB1_1_9/i0[8] ) );
  INV_X2 \SB1_1_10/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[129] ), .ZN(
        \SB1_1_10/i0[8] ) );
  INV_X2 \SB1_1_10/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[128] ), .ZN(
        \SB1_1_10/i1[9] ) );
  INV_X1 \SB1_1_11/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[124] ), .ZN(
        \SB1_1_11/i0[7] ) );
  INV_X1 \SB1_1_12/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[118] ), .ZN(
        \SB1_1_12/i0[7] ) );
  INV_X2 \SB1_1_12/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[116] ), .ZN(
        \SB1_1_12/i1[9] ) );
  INV_X1 \SB1_1_13/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[112] ), .ZN(
        \SB1_1_13/i0[7] ) );
  INV_X2 \SB1_1_13/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[111] ), .ZN(
        \SB1_1_13/i0[8] ) );
  INV_X1 \SB1_1_13/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[108] ), .ZN(
        \SB1_1_13/i3[0] ) );
  INV_X1 \SB1_1_14/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[106] ), .ZN(
        \SB1_1_14/i0[7] ) );
  INV_X2 \SB1_1_14/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[105] ), .ZN(
        \SB1_1_14/i0[8] ) );
  INV_X1 \SB1_1_15/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[100] ), .ZN(
        \SB1_1_15/i0[7] ) );
  INV_X1 \SB1_1_15/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[96] ), .ZN(
        \SB1_1_15/i3[0] ) );
  INV_X2 \SB1_1_16/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[92] ), .ZN(
        \SB1_1_16/i1[9] ) );
  INV_X1 \SB1_1_16/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[90] ), .ZN(
        \SB1_1_16/i3[0] ) );
  INV_X1 \SB1_1_17/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[88] ), .ZN(
        \SB1_1_17/i0[7] ) );
  INV_X2 \SB1_1_17/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[87] ), .ZN(
        \SB1_1_17/i0[8] ) );
  INV_X1 \SB1_1_17/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[85] ), .ZN(
        \SB1_1_17/i1_7 ) );
  INV_X2 \SB1_1_18/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[80] ), .ZN(
        \SB1_1_18/i1[9] ) );
  INV_X1 \SB1_1_19/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[76] ), .ZN(
        \SB1_1_19/i0[7] ) );
  INV_X1 \SB1_1_19/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[73] ), .ZN(
        \SB1_1_19/i1_7 ) );
  INV_X1 \SB1_1_20/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[70] ), .ZN(
        \SB1_1_20/i0[7] ) );
  INV_X2 \SB1_1_20/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[69] ), .ZN(
        \SB1_1_20/i0[8] ) );
  INV_X1 \SB1_1_22/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[58] ), .ZN(
        \SB1_1_22/i0[7] ) );
  INV_X2 \SB1_1_22/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[57] ), .ZN(
        \SB1_1_22/i0[8] ) );
  INV_X2 \SB1_1_23/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[51] ), .ZN(
        \SB1_1_23/i0[8] ) );
  INV_X1 \SB1_1_24/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[46] ), .ZN(
        \SB1_1_24/i0[7] ) );
  INV_X2 \SB1_1_24/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[45] ), .ZN(
        \SB1_1_24/i0[8] ) );
  INV_X1 \SB1_1_25/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[40] ), .ZN(
        \SB1_1_25/i0[7] ) );
  INV_X1 \SB1_1_26/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[34] ), .ZN(
        \SB1_1_26/i0[7] ) );
  INV_X1 \SB1_1_27/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[28] ), .ZN(
        \SB1_1_27/i0[7] ) );
  INV_X1 \SB1_1_28/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[22] ), .ZN(
        \SB1_1_28/i0[7] ) );
  INV_X2 \SB1_1_28/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[21] ), .ZN(
        \SB1_1_28/i0[8] ) );
  INV_X1 \SB1_1_29/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[16] ), .ZN(
        \SB1_1_29/i0[7] ) );
  INV_X2 \SB1_1_29/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[15] ), .ZN(
        \SB1_1_29/i0[8] ) );
  INV_X2 \SB1_1_29/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[14] ), .ZN(
        \SB1_1_29/i1[9] ) );
  INV_X1 \SB1_1_29/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[13] ), .ZN(
        \SB1_1_29/i1_7 ) );
  INV_X2 \SB1_1_31/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[3] ), .ZN(
        \SB1_1_31/i0[8] ) );
  INV_X1 \SB1_1_31/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[0] ), .ZN(
        \SB1_1_31/i3[0] ) );
  INV_X1 \SB2_1_0/INV_0  ( .I(\SB1_1_5/buf_output[0] ), .ZN(\SB2_1_0/i3[0] )
         );
  INV_X1 \SB2_1_1/INV_4  ( .I(\SB1_1_2/buf_output[4] ), .ZN(\SB2_1_1/i0[7] )
         );
  INV_X1 \SB2_1_1/INV_0  ( .I(\SB1_1_6/buf_output[0] ), .ZN(\SB2_1_1/i3[0] )
         );
  INV_X1 \SB2_1_2/INV_0  ( .I(\SB1_1_7/buf_output[0] ), .ZN(\SB2_1_2/i3[0] )
         );
  INV_X1 \SB2_1_3/INV_4  ( .I(\SB1_1_4/buf_output[4] ), .ZN(\SB2_1_3/i0[7] )
         );
  INV_X1 \SB2_1_4/INV_4  ( .I(\SB1_1_5/buf_output[4] ), .ZN(\SB2_1_4/i0[7] )
         );
  INV_X1 \SB2_1_4/INV_0  ( .I(\SB1_1_9/buf_output[0] ), .ZN(\SB2_1_4/i3[0] )
         );
  INV_X2 \SB2_1_5/INV_2  ( .I(\SB1_1_8/buf_output[2] ), .ZN(\SB2_1_5/i1[9] )
         );
  INV_X1 \SB2_1_6/INV_4  ( .I(\SB1_1_7/buf_output[4] ), .ZN(\SB2_1_6/i0[7] )
         );
  INV_X1 \SB2_1_6/INV_0  ( .I(\SB1_1_11/buf_output[0] ), .ZN(\SB2_1_6/i3[0] )
         );
  INV_X1 \SB2_1_7/INV_0  ( .I(\SB1_1_12/buf_output[0] ), .ZN(\SB2_1_7/i3[0] )
         );
  INV_X1 \SB2_1_8/INV_0  ( .I(\SB1_1_13/buf_output[0] ), .ZN(\SB2_1_8/i3[0] )
         );
  INV_X1 \SB2_1_9/INV_4  ( .I(\SB1_1_10/buf_output[4] ), .ZN(\SB2_1_9/i0[7] )
         );
  INV_X2 \SB2_1_9/INV_3  ( .I(\SB1_1_11/buf_output[3] ), .ZN(\SB2_1_9/i0[8] )
         );
  INV_X1 \SB2_1_9/INV_0  ( .I(\SB1_1_14/buf_output[0] ), .ZN(\SB2_1_9/i3[0] )
         );
  INV_X1 \SB2_1_10/INV_4  ( .I(\SB1_1_11/buf_output[4] ), .ZN(\SB2_1_10/i0[7] ) );
  INV_X2 \SB2_1_10/INV_3  ( .I(\SB1_1_12/buf_output[3] ), .ZN(\SB2_1_10/i0[8] ) );
  INV_X1 \SB2_1_10/INV_0  ( .I(\SB1_1_15/buf_output[0] ), .ZN(\SB2_1_10/i3[0] ) );
  INV_X1 \SB2_1_11/INV_4  ( .I(\SB1_1_12/buf_output[4] ), .ZN(\SB2_1_11/i0[7] ) );
  INV_X1 \SB2_1_12/INV_4  ( .I(\SB1_1_13/buf_output[4] ), .ZN(\SB2_1_12/i0[7] ) );
  INV_X1 \SB2_1_12/INV_0  ( .I(\SB1_1_17/buf_output[0] ), .ZN(\SB2_1_12/i3[0] ) );
  INV_X1 \SB2_1_13/INV_0  ( .I(\SB1_1_18/buf_output[0] ), .ZN(\SB2_1_13/i3[0] ) );
  INV_X1 \SB2_1_14/INV_4  ( .I(\SB1_1_15/buf_output[4] ), .ZN(\SB2_1_14/i0[7] ) );
  INV_X1 \SB2_1_14/INV_0  ( .I(\SB1_1_19/buf_output[0] ), .ZN(\SB2_1_14/i3[0] ) );
  INV_X1 \SB2_1_15/INV_4  ( .I(\SB1_1_16/buf_output[4] ), .ZN(\SB2_1_15/i0[7] ) );
  INV_X1 \SB2_1_15/INV_0  ( .I(\SB1_1_20/buf_output[0] ), .ZN(\SB2_1_15/i3[0] ) );
  INV_X1 \SB2_1_16/INV_4  ( .I(\SB1_1_17/buf_output[4] ), .ZN(\SB2_1_16/i0[7] ) );
  INV_X2 \SB2_1_16/INV_2  ( .I(\SB1_1_19/buf_output[2] ), .ZN(\SB2_1_16/i1[9] ) );
  INV_X1 \SB2_1_17/INV_4  ( .I(\SB1_1_18/buf_output[4] ), .ZN(\SB2_1_17/i0[7] ) );
  INV_X2 \SB2_1_17/INV_3  ( .I(\SB1_1_19/buf_output[3] ), .ZN(\SB2_1_17/i0[8] ) );
  INV_X1 \SB2_1_17/INV_0  ( .I(\SB1_1_22/buf_output[0] ), .ZN(\SB2_1_17/i3[0] ) );
  INV_X1 \SB2_1_18/INV_4  ( .I(\SB1_1_19/buf_output[4] ), .ZN(\SB2_1_18/i0[7] ) );
  INV_X2 \SB2_1_18/INV_3  ( .I(\SB1_1_20/buf_output[3] ), .ZN(\SB2_1_18/i0[8] ) );
  INV_X1 \SB2_1_18/INV_0  ( .I(\SB1_1_23/buf_output[0] ), .ZN(\SB2_1_18/i3[0] ) );
  INV_X2 \SB2_1_20/INV_3  ( .I(\SB1_1_22/buf_output[3] ), .ZN(\SB2_1_20/i0[8] ) );
  INV_X1 \SB2_1_20/INV_0  ( .I(\SB1_1_25/buf_output[0] ), .ZN(\SB2_1_20/i3[0] ) );
  INV_X1 \SB2_1_21/INV_4  ( .I(\SB1_1_22/buf_output[4] ), .ZN(\SB2_1_21/i0[7] ) );
  INV_X1 \SB2_1_21/INV_0  ( .I(\SB1_1_26/buf_output[0] ), .ZN(\SB2_1_21/i3[0] ) );
  INV_X1 \SB2_1_22/INV_0  ( .I(\SB1_1_27/buf_output[0] ), .ZN(\SB2_1_22/i3[0] ) );
  INV_X1 \SB2_1_23/INV_4  ( .I(\SB1_1_24/buf_output[4] ), .ZN(\SB2_1_23/i0[7] ) );
  INV_X2 \SB2_1_23/INV_3  ( .I(\SB1_1_25/buf_output[3] ), .ZN(\SB2_1_23/i0[8] ) );
  INV_X1 \SB2_1_24/INV_4  ( .I(\SB1_1_25/buf_output[4] ), .ZN(\SB2_1_24/i0[7] ) );
  INV_X1 \SB2_1_24/INV_0  ( .I(\SB1_1_29/buf_output[0] ), .ZN(\SB2_1_24/i3[0] ) );
  INV_X1 \SB2_1_25/INV_4  ( .I(\SB1_1_26/buf_output[4] ), .ZN(\SB2_1_25/i0[7] ) );
  INV_X1 \SB2_1_25/INV_0  ( .I(\SB1_1_30/buf_output[0] ), .ZN(\SB2_1_25/i3[0] ) );
  INV_X1 \SB2_1_26/INV_4  ( .I(\SB1_1_27/buf_output[4] ), .ZN(\SB2_1_26/i0[7] ) );
  INV_X1 \SB2_1_26/INV_0  ( .I(\SB1_1_31/buf_output[0] ), .ZN(\SB2_1_26/i3[0] ) );
  INV_X1 \SB2_1_27/INV_4  ( .I(\SB1_1_28/buf_output[4] ), .ZN(\SB2_1_27/i0[7] ) );
  INV_X1 \SB2_1_27/INV_0  ( .I(\SB1_1_0/buf_output[0] ), .ZN(\SB2_1_27/i3[0] )
         );
  INV_X1 \SB2_1_30/INV_4  ( .I(\SB1_1_31/buf_output[4] ), .ZN(\SB2_1_30/i0[7] ) );
  INV_X1 \SB2_1_30/INV_0  ( .I(\SB1_1_3/buf_output[0] ), .ZN(\SB2_1_30/i3[0] )
         );
  INV_X1 \SB2_1_31/INV_0  ( .I(\SB1_1_4/buf_output[0] ), .ZN(\SB2_1_31/i3[0] )
         );
  INV_X1 \SB1_2_0/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[190] ), .ZN(
        \SB1_2_0/i0[7] ) );
  INV_X2 \SB1_2_0/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[189] ), .ZN(
        \SB1_2_0/i0[8] ) );
  INV_X1 \SB1_2_1/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[184] ), .ZN(
        \SB1_2_1/i0[7] ) );
  INV_X1 \SB1_2_2/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[178] ), .ZN(
        \SB1_2_2/i0[7] ) );
  INV_X2 \SB1_2_2/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[177] ), .ZN(
        \SB1_2_2/i0[8] ) );
  INV_X1 \SB1_2_2/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[174] ), .ZN(
        \SB1_2_2/i3[0] ) );
  INV_X1 \SB1_2_3/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[172] ), .ZN(
        \SB1_2_3/i0[7] ) );
  INV_X2 \SB1_2_3/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[171] ), .ZN(
        \SB1_2_3/i0[8] ) );
  INV_X2 \SB1_2_3/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[170] ), .ZN(
        \SB1_2_3/i1[9] ) );
  INV_X1 \SB1_2_4/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[166] ), .ZN(
        \SB1_2_4/i0[7] ) );
  INV_X1 \SB1_2_5/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[160] ), .ZN(
        \SB1_2_5/i0[7] ) );
  INV_X2 \SB1_2_5/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[159] ), .ZN(
        \SB1_2_5/i0[8] ) );
  INV_X1 \SB1_2_5/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[156] ), .ZN(
        \SB1_2_5/i3[0] ) );
  INV_X1 \SB1_2_6/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[154] ), .ZN(
        \SB1_2_6/i0[7] ) );
  INV_X1 \SB1_2_7/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[148] ), .ZN(
        \SB1_2_7/i0[7] ) );
  INV_X1 \SB1_2_7/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[144] ), .ZN(
        \SB1_2_7/i3[0] ) );
  INV_X1 \SB1_2_8/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[142] ), .ZN(
        \SB1_2_8/i0[7] ) );
  INV_X1 \SB1_2_9/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[136] ), .ZN(
        \SB1_2_9/i0[7] ) );
  INV_X2 \SB1_2_9/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[135] ), .ZN(
        \SB1_2_9/i0[8] ) );
  INV_X1 \SB1_2_10/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[130] ), .ZN(
        \SB1_2_10/i0[7] ) );
  INV_X2 \SB1_2_10/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[129] ), .ZN(
        \SB1_2_10/i0[8] ) );
  INV_X2 \SB1_2_10/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[128] ), .ZN(
        \SB1_2_10/i1[9] ) );
  INV_X1 \SB1_2_11/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[124] ), .ZN(
        \SB1_2_11/i0[7] ) );
  INV_X2 \SB1_2_11/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[122] ), .ZN(
        \SB1_2_11/i1[9] ) );
  INV_X1 \SB1_2_12/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[118] ), .ZN(
        \SB1_2_12/i0[7] ) );
  INV_X2 \SB1_2_12/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[117] ), .ZN(
        \SB1_2_12/i0[8] ) );
  INV_X1 \SB1_2_12/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[114] ), .ZN(
        \SB1_2_12/i3[0] ) );
  INV_X1 \SB1_2_13/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[112] ), .ZN(
        \SB1_2_13/i0[7] ) );
  INV_X1 \SB1_2_13/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[108] ), .ZN(
        \SB1_2_13/i3[0] ) );
  INV_X1 \SB1_2_14/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[106] ), .ZN(
        \SB1_2_14/i0[7] ) );
  INV_X1 \SB1_2_14/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[102] ), .ZN(
        \SB1_2_14/i3[0] ) );
  INV_X1 \SB1_2_15/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[100] ), .ZN(
        \SB1_2_15/i0[7] ) );
  INV_X2 \SB1_2_15/INV_3  ( .I(n1509), .ZN(\SB1_2_15/i0[8] ) );
  INV_X1 \SB1_2_15/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[97] ), .ZN(
        \SB1_2_15/i1_7 ) );
  INV_X1 \SB1_2_16/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[94] ), .ZN(
        \SB1_2_16/i0[7] ) );
  INV_X2 \SB1_2_16/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[92] ), .ZN(
        \SB1_2_16/i1[9] ) );
  INV_X1 \SB1_2_16/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[91] ), .ZN(
        \SB1_2_16/i1_7 ) );
  INV_X1 \SB1_2_17/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[88] ), .ZN(
        \SB1_2_17/i0[7] ) );
  INV_X2 \SB1_2_17/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[87] ), .ZN(
        \SB1_2_17/i0[8] ) );
  INV_X2 \SB1_2_18/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[81] ), .ZN(
        \SB1_2_18/i0[8] ) );
  INV_X2 \SB1_2_18/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[80] ), .ZN(
        \SB1_2_18/i1[9] ) );
  INV_X1 \SB1_2_19/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[76] ), .ZN(
        \SB1_2_19/i0[7] ) );
  INV_X2 \SB1_2_19/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[75] ), .ZN(
        \SB1_2_19/i0[8] ) );
  INV_X1 \SB1_2_20/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[70] ), .ZN(
        \SB1_2_20/i0[7] ) );
  INV_X2 \SB1_2_20/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[69] ), .ZN(
        \SB1_2_20/i0[8] ) );
  INV_X1 \SB1_2_20/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[66] ), .ZN(
        \SB1_2_20/i3[0] ) );
  INV_X1 \SB1_2_21/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[64] ), .ZN(
        \SB1_2_21/i0[7] ) );
  INV_X1 \SB1_2_22/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[58] ), .ZN(
        \SB1_2_22/i0[7] ) );
  INV_X1 \SB1_2_22/INV_0  ( .I(n6938), .ZN(\SB1_2_22/i3[0] ) );
  INV_X1 \SB1_2_23/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[52] ), .ZN(
        \SB1_2_23/i0[7] ) );
  INV_X1 \SB1_2_24/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[46] ), .ZN(
        \SB1_2_24/i0[7] ) );
  INV_X2 \SB1_2_24/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[45] ), .ZN(
        \SB1_2_24/i0[8] ) );
  INV_X2 \SB1_2_24/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[44] ), .ZN(
        \SB1_2_24/i1[9] ) );
  INV_X1 \SB1_2_25/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[40] ), .ZN(
        \SB1_2_25/i0[7] ) );
  INV_X1 \SB1_2_25/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[37] ), .ZN(
        \SB1_2_25/i1_7 ) );
  INV_X1 \SB1_2_26/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[34] ), .ZN(
        \SB1_2_26/i0[7] ) );
  INV_X2 \SB1_2_26/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[33] ), .ZN(
        \SB1_2_26/i0[8] ) );
  INV_X1 \SB1_2_27/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[28] ), .ZN(
        \SB1_2_27/i0[7] ) );
  INV_X1 \SB1_2_28/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[22] ), .ZN(
        \SB1_2_28/i0[7] ) );
  INV_X2 \SB1_2_28/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[20] ), .ZN(
        \SB1_2_28/i1[9] ) );
  INV_X1 \SB1_2_29/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[16] ), .ZN(
        \SB1_2_29/i0[7] ) );
  INV_X2 \SB1_2_29/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[15] ), .ZN(
        \SB1_2_29/i0[8] ) );
  INV_X1 \SB1_2_29/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[12] ), .ZN(
        \SB1_2_29/i3[0] ) );
  INV_X1 \SB1_2_30/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[10] ), .ZN(
        \SB1_2_30/i0[7] ) );
  INV_X2 \SB1_2_30/INV_3  ( .I(\RI1[2][9] ), .ZN(\SB1_2_30/i0[8] ) );
  INV_X1 \SB1_2_30/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[6] ), .ZN(
        \SB1_2_30/i3[0] ) );
  INV_X1 \SB1_2_31/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[4] ), .ZN(
        \SB1_2_31/i0[7] ) );
  INV_X2 \SB1_2_31/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[3] ), .ZN(
        \SB1_2_31/i0[8] ) );
  INV_X2 \SB2_2_1/INV_3  ( .I(\SB1_2_3/buf_output[3] ), .ZN(\SB2_2_1/i0[8] )
         );
  INV_X1 \SB2_2_1/INV_0  ( .I(\SB1_2_6/buf_output[0] ), .ZN(\SB2_2_1/i3[0] )
         );
  INV_X1 \SB2_2_2/INV_4  ( .I(\SB1_2_3/buf_output[4] ), .ZN(\SB2_2_2/i0[7] )
         );
  INV_X1 \SB2_2_2/INV_1  ( .I(\SB1_2_6/buf_output[1] ), .ZN(\SB2_2_2/i1_7 ) );
  INV_X1 \SB2_2_3/INV_4  ( .I(\SB1_2_4/buf_output[4] ), .ZN(\SB2_2_3/i0[7] )
         );
  INV_X1 \SB2_2_3/INV_1  ( .I(\SB1_2_7/buf_output[1] ), .ZN(\SB2_2_3/i1_7 ) );
  INV_X2 \SB2_2_4/INV_3  ( .I(\SB1_2_6/buf_output[3] ), .ZN(\SB2_2_4/i0[8] )
         );
  INV_X1 \SB2_2_4/INV_1  ( .I(\SB1_2_8/buf_output[1] ), .ZN(\SB2_2_4/i1_7 ) );
  INV_X1 \SB2_2_4/INV_0  ( .I(\SB1_2_9/buf_output[0] ), .ZN(\SB2_2_4/i3[0] )
         );
  INV_X1 \SB2_2_5/INV_4  ( .I(\SB1_2_6/buf_output[4] ), .ZN(\SB2_2_5/i0[7] )
         );
  INV_X1 \SB2_2_6/INV_4  ( .I(\SB1_2_7/buf_output[4] ), .ZN(\SB2_2_6/i0[7] )
         );
  INV_X1 \SB2_2_6/INV_0  ( .I(\SB1_2_11/buf_output[0] ), .ZN(\SB2_2_6/i3[0] )
         );
  INV_X1 \SB2_2_7/INV_4  ( .I(\SB1_2_8/buf_output[4] ), .ZN(\SB2_2_7/i0[7] )
         );
  INV_X1 \SB2_2_7/INV_0  ( .I(\SB1_2_12/buf_output[0] ), .ZN(\SB2_2_7/i3[0] )
         );
  INV_X1 \SB2_2_8/INV_4  ( .I(\SB1_2_9/buf_output[4] ), .ZN(\SB2_2_8/i0[7] )
         );
  INV_X1 \SB2_2_9/INV_4  ( .I(\SB1_2_10/buf_output[4] ), .ZN(\SB2_2_9/i0[7] )
         );
  INV_X1 \SB2_2_10/INV_4  ( .I(\SB1_2_11/buf_output[4] ), .ZN(\SB2_2_10/i0[7] ) );
  INV_X1 \SB2_2_10/INV_0  ( .I(\SB1_2_15/buf_output[0] ), .ZN(\SB2_2_10/i3[0] ) );
  INV_X1 \SB2_2_11/INV_4  ( .I(\SB1_2_12/buf_output[4] ), .ZN(\SB2_2_11/i0[7] ) );
  INV_X2 \SB2_2_11/INV_3  ( .I(\SB1_2_13/buf_output[3] ), .ZN(\SB2_2_11/i0[8] ) );
  INV_X2 \SB2_2_11/INV_2  ( .I(\SB1_2_14/buf_output[2] ), .ZN(\SB2_2_11/i1[9] ) );
  INV_X1 \SB2_2_11/INV_0  ( .I(\SB1_2_16/buf_output[0] ), .ZN(\SB2_2_11/i3[0] ) );
  INV_X1 \SB2_2_12/INV_4  ( .I(\SB1_2_13/buf_output[4] ), .ZN(\SB2_2_12/i0[7] ) );
  INV_X1 \SB2_2_12/INV_0  ( .I(\SB1_2_17/buf_output[0] ), .ZN(\SB2_2_12/i3[0] ) );
  INV_X1 \SB2_2_13/INV_4  ( .I(\SB1_2_14/buf_output[4] ), .ZN(\SB2_2_13/i0[7] ) );
  INV_X1 \SB2_2_14/INV_4  ( .I(\SB1_2_15/buf_output[4] ), .ZN(\SB2_2_14/i0[7] ) );
  INV_X1 \SB2_2_14/INV_0  ( .I(\SB1_2_19/buf_output[0] ), .ZN(\SB2_2_14/i3[0] ) );
  INV_X1 \SB2_2_15/INV_4  ( .I(\SB1_2_16/buf_output[4] ), .ZN(\SB2_2_15/i0[7] ) );
  INV_X1 \SB2_2_16/INV_4  ( .I(\SB1_2_17/buf_output[4] ), .ZN(\SB2_2_16/i0[7] ) );
  INV_X2 \SB2_2_16/INV_3  ( .I(\SB1_2_18/buf_output[3] ), .ZN(\SB2_2_16/i0[8] ) );
  INV_X1 \SB2_2_16/INV_0  ( .I(\SB1_2_21/buf_output[0] ), .ZN(\SB2_2_16/i3[0] ) );
  INV_X1 \SB2_2_17/INV_4  ( .I(\SB1_2_18/buf_output[4] ), .ZN(\SB2_2_17/i0[7] ) );
  INV_X1 \SB2_2_18/INV_0  ( .I(\SB1_2_23/buf_output[0] ), .ZN(\SB2_2_18/i3[0] ) );
  INV_X1 \SB2_2_19/INV_4  ( .I(\SB1_2_20/buf_output[4] ), .ZN(\SB2_2_19/i0[7] ) );
  INV_X1 \SB2_2_19/INV_1  ( .I(\SB1_2_23/buf_output[1] ), .ZN(\SB2_2_19/i1_7 )
         );
  INV_X1 \SB2_2_20/INV_4  ( .I(\SB1_2_21/buf_output[4] ), .ZN(\SB2_2_20/i0[7] ) );
  INV_X1 \SB2_2_20/INV_0  ( .I(\SB1_2_25/buf_output[0] ), .ZN(\SB2_2_20/i3[0] ) );
  INV_X2 \SB2_2_21/INV_3  ( .I(\SB1_2_23/buf_output[3] ), .ZN(\SB2_2_21/i0[8] ) );
  INV_X1 \SB2_2_22/INV_4  ( .I(\SB1_2_23/buf_output[4] ), .ZN(\SB2_2_22/i0[7] ) );
  INV_X1 \SB2_2_23/INV_0  ( .I(\SB1_2_28/buf_output[0] ), .ZN(\SB2_2_23/i3[0] ) );
  INV_X1 \SB2_2_24/INV_4  ( .I(\SB1_2_25/buf_output[4] ), .ZN(\SB2_2_24/i0[7] ) );
  INV_X1 \SB2_2_24/INV_1  ( .I(\SB1_2_28/buf_output[1] ), .ZN(\SB2_2_24/i1_7 )
         );
  INV_X1 \SB2_2_24/INV_0  ( .I(\SB1_2_29/buf_output[0] ), .ZN(\SB2_2_24/i3[0] ) );
  INV_X1 \SB2_2_25/INV_4  ( .I(\SB1_2_26/buf_output[4] ), .ZN(\SB2_2_25/i0[7] ) );
  INV_X1 \SB2_2_25/INV_0  ( .I(\SB1_2_30/buf_output[0] ), .ZN(\SB2_2_25/i3[0] ) );
  INV_X1 \SB2_2_27/INV_1  ( .I(\SB1_2_31/buf_output[1] ), .ZN(\SB2_2_27/i1_7 )
         );
  INV_X1 \SB2_2_27/INV_0  ( .I(\SB1_2_0/buf_output[0] ), .ZN(\SB2_2_27/i3[0] )
         );
  INV_X1 \SB2_2_28/INV_4  ( .I(\SB1_2_29/buf_output[4] ), .ZN(\SB2_2_28/i0[7] ) );
  INV_X1 \SB2_2_28/INV_0  ( .I(\SB1_2_1/buf_output[0] ), .ZN(\SB2_2_28/i3[0] )
         );
  INV_X1 \SB2_2_29/INV_4  ( .I(\SB1_2_30/buf_output[4] ), .ZN(\SB2_2_29/i0[7] ) );
  INV_X1 \SB2_2_29/INV_0  ( .I(\SB1_2_2/buf_output[0] ), .ZN(\SB2_2_29/i3[0] )
         );
  INV_X1 \SB2_2_30/INV_4  ( .I(\SB1_2_31/buf_output[4] ), .ZN(\SB2_2_30/i0[7] ) );
  INV_X1 \SB2_2_30/INV_1  ( .I(\SB1_2_2/buf_output[1] ), .ZN(\SB2_2_30/i1_7 )
         );
  INV_X1 \SB2_2_30/INV_0  ( .I(\SB1_2_3/buf_output[0] ), .ZN(\SB2_2_30/i3[0] )
         );
  INV_X1 \SB2_2_31/INV_4  ( .I(\SB1_2_0/buf_output[4] ), .ZN(\SB2_2_31/i0[7] )
         );
  INV_X1 \SB2_2_31/INV_0  ( .I(\SB1_2_4/buf_output[0] ), .ZN(\SB2_2_31/i3[0] )
         );
  INV_X1 \SB1_3_0/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[190] ), .ZN(
        \SB1_3_0/i0[7] ) );
  INV_X2 \SB1_3_0/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[189] ), .ZN(
        \SB1_3_0/i0[8] ) );
  INV_X1 \SB1_3_0/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[186] ), .ZN(
        \SB1_3_0/i3[0] ) );
  INV_X1 \SB1_3_1/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[184] ), .ZN(
        \SB1_3_1/i0[7] ) );
  INV_X1 \SB1_3_2/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[178] ), .ZN(
        \SB1_3_2/i0[7] ) );
  INV_X1 \SB1_3_2/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[174] ), .ZN(
        \SB1_3_2/i3[0] ) );
  INV_X1 \SB1_3_3/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[172] ), .ZN(
        \SB1_3_3/i0[7] ) );
  INV_X2 \SB1_3_3/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[171] ), .ZN(
        \SB1_3_3/i0[8] ) );
  INV_X1 \SB1_3_4/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[166] ), .ZN(
        \SB1_3_4/i0[7] ) );
  INV_X1 \SB1_3_5/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[160] ), .ZN(
        \SB1_3_5/i0[7] ) );
  INV_X2 \SB1_3_5/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[159] ), .ZN(
        \SB1_3_5/i0[8] ) );
  INV_X1 \SB1_3_7/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[148] ), .ZN(
        \SB1_3_7/i0[7] ) );
  INV_X1 \SB1_3_7/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[144] ), .ZN(
        \SB1_3_7/i3[0] ) );
  INV_X1 \SB1_3_8/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[142] ), .ZN(
        \SB1_3_8/i0[7] ) );
  INV_X2 \SB1_3_8/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[141] ), .ZN(
        \SB1_3_8/i0[8] ) );
  INV_X1 \SB1_3_9/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[136] ), .ZN(
        \SB1_3_9/i0[7] ) );
  INV_X1 \SB1_3_10/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[130] ), .ZN(
        \SB1_3_10/i0[7] ) );
  INV_X1 \SB1_3_11/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[124] ), .ZN(
        \SB1_3_11/i0[7] ) );
  INV_X2 \SB1_3_11/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[123] ), .ZN(
        \SB1_3_11/i0[8] ) );
  INV_X1 \SB1_3_12/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[118] ), .ZN(
        \SB1_3_12/i0[7] ) );
  INV_X1 \SB1_3_13/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[112] ), .ZN(
        \SB1_3_13/i0[7] ) );
  INV_X2 \SB1_3_13/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[111] ), .ZN(
        \SB1_3_13/i0[8] ) );
  INV_X1 \SB1_3_13/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[108] ), .ZN(
        \SB1_3_13/i3[0] ) );
  INV_X1 \SB1_3_14/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[106] ), .ZN(
        \SB1_3_14/i0[7] ) );
  INV_X1 \SB1_3_14/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[102] ), .ZN(
        \SB1_3_14/i3[0] ) );
  INV_X1 \SB1_3_15/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[100] ), .ZN(
        \SB1_3_15/i0[7] ) );
  INV_X1 \SB1_3_16/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[94] ), .ZN(
        \SB1_3_16/i0[7] ) );
  INV_X2 \SB1_3_16/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[92] ), .ZN(
        \SB1_3_16/i1[9] ) );
  INV_X1 \SB1_3_18/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[82] ), .ZN(
        \SB1_3_18/i0[7] ) );
  INV_X2 \SB1_3_18/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[81] ), .ZN(
        \SB1_3_18/i0[8] ) );
  INV_X1 \SB1_3_18/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[79] ), .ZN(
        \SB1_3_18/i1_7 ) );
  INV_X1 \SB1_3_19/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[76] ), .ZN(
        \SB1_3_19/i0[7] ) );
  INV_X1 \SB1_3_21/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[64] ), .ZN(
        \SB1_3_21/i0[7] ) );
  INV_X1 \SB1_3_22/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[58] ), .ZN(
        \SB1_3_22/i0[7] ) );
  INV_X1 \SB1_3_23/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[52] ), .ZN(
        \SB1_3_23/i0[7] ) );
  INV_X2 \SB1_3_23/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[51] ), .ZN(
        \SB1_3_23/i0[8] ) );
  INV_X1 \SB1_3_24/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[46] ), .ZN(
        \SB1_3_24/i0[7] ) );
  INV_X1 \SB1_3_25/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[40] ), .ZN(
        \SB1_3_25/i0[7] ) );
  INV_X2 \SB1_3_25/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[39] ), .ZN(
        \SB1_3_25/i0[8] ) );
  INV_X1 \SB1_3_26/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[34] ), .ZN(
        \SB1_3_26/i0[7] ) );
  INV_X1 \SB1_3_26/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[31] ), .ZN(
        \SB1_3_26/i1_7 ) );
  INV_X1 \SB1_3_28/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[22] ), .ZN(
        \SB1_3_28/i0[7] ) );
  INV_X2 \SB1_3_28/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[21] ), .ZN(
        \SB1_3_28/i0[8] ) );
  INV_X2 \SB1_3_28/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[20] ), .ZN(
        \SB1_3_28/i1[9] ) );
  INV_X1 \SB1_3_29/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[16] ), .ZN(
        \SB1_3_29/i0[7] ) );
  INV_X1 \SB1_3_30/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[10] ), .ZN(
        \SB1_3_30/i0[7] ) );
  INV_X1 \SB1_3_30/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[6] ), .ZN(
        \SB1_3_30/i3[0] ) );
  INV_X1 \SB1_3_31/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[4] ), .ZN(
        \SB1_3_31/i0[7] ) );
  INV_X1 \SB2_3_0/INV_4  ( .I(\SB1_3_1/buf_output[4] ), .ZN(\SB2_3_0/i0[7] )
         );
  INV_X1 \SB2_3_0/INV_0  ( .I(\SB1_3_5/buf_output[0] ), .ZN(\SB2_3_0/i3[0] )
         );
  INV_X1 \SB2_3_1/INV_4  ( .I(\SB1_3_2/buf_output[4] ), .ZN(\SB2_3_1/i0[7] )
         );
  INV_X1 \SB2_3_1/INV_1  ( .I(\SB1_3_5/buf_output[1] ), .ZN(\SB2_3_1/i1_7 ) );
  INV_X1 \SB2_3_2/INV_4  ( .I(\SB1_3_3/buf_output[4] ), .ZN(\SB2_3_2/i0[7] )
         );
  INV_X2 \SB2_3_3/INV_3  ( .I(\SB1_3_5/buf_output[3] ), .ZN(\SB2_3_3/i0[8] )
         );
  INV_X1 \SB2_3_3/INV_0  ( .I(\SB1_3_8/buf_output[0] ), .ZN(\SB2_3_3/i3[0] )
         );
  INV_X1 \SB2_3_4/INV_1  ( .I(\SB1_3_8/buf_output[1] ), .ZN(\SB2_3_4/i1_7 ) );
  INV_X2 \SB2_3_5/INV_3  ( .I(\SB1_3_7/buf_output[3] ), .ZN(\SB2_3_5/i0[8] )
         );
  INV_X1 \SB2_3_5/INV_0  ( .I(\SB1_3_10/buf_output[0] ), .ZN(\SB2_3_5/i3[0] )
         );
  INV_X1 \SB2_3_8/INV_4  ( .I(\SB1_3_9/buf_output[4] ), .ZN(\SB2_3_8/i0[7] )
         );
  INV_X1 \SB2_3_8/INV_0  ( .I(\SB1_3_13/buf_output[0] ), .ZN(\SB2_3_8/i3[0] )
         );
  INV_X1 \SB2_3_9/INV_0  ( .I(\SB1_3_14/buf_output[0] ), .ZN(\SB2_3_9/i3[0] )
         );
  INV_X1 \SB2_3_10/INV_0  ( .I(\SB1_3_15/buf_output[0] ), .ZN(\SB2_3_10/i3[0] ) );
  INV_X1 \SB2_3_11/INV_4  ( .I(\SB1_3_12/buf_output[4] ), .ZN(\SB2_3_11/i0[7] ) );
  INV_X2 \SB2_3_11/INV_3  ( .I(\SB1_3_13/buf_output[3] ), .ZN(\SB2_3_11/i0[8] ) );
  INV_X1 \SB2_3_13/INV_0  ( .I(\SB1_3_18/buf_output[0] ), .ZN(\SB2_3_13/i3[0] ) );
  INV_X1 \SB2_3_14/INV_4  ( .I(\SB1_3_15/buf_output[4] ), .ZN(\SB2_3_14/i0[7] ) );
  INV_X1 \SB2_3_14/INV_0  ( .I(\SB1_3_19/buf_output[0] ), .ZN(\SB2_3_14/i3[0] ) );
  INV_X1 \SB2_3_15/INV_4  ( .I(\SB1_3_16/buf_output[4] ), .ZN(\SB2_3_15/i0[7] ) );
  INV_X1 \SB2_3_15/INV_0  ( .I(\SB1_3_20/buf_output[0] ), .ZN(\SB2_3_15/i3[0] ) );
  INV_X1 \SB2_3_16/INV_4  ( .I(\SB1_3_17/buf_output[4] ), .ZN(\SB2_3_16/i0[7] ) );
  INV_X1 \SB2_3_16/INV_0  ( .I(\SB1_3_21/buf_output[0] ), .ZN(\SB2_3_16/i3[0] ) );
  INV_X1 \SB2_3_17/INV_4  ( .I(\SB1_3_18/buf_output[4] ), .ZN(\SB2_3_17/i0[7] ) );
  INV_X1 \SB2_3_17/INV_0  ( .I(\SB1_3_22/buf_output[0] ), .ZN(\SB2_3_17/i3[0] ) );
  INV_X1 \SB2_3_18/INV_4  ( .I(\SB1_3_19/buf_output[4] ), .ZN(\SB2_3_18/i0[7] ) );
  INV_X1 \SB2_3_18/INV_0  ( .I(\SB1_3_23/buf_output[0] ), .ZN(\SB2_3_18/i3[0] ) );
  INV_X1 \SB2_3_21/INV_0  ( .I(\SB1_3_26/buf_output[0] ), .ZN(\SB2_3_21/i3[0] ) );
  INV_X1 \SB2_3_22/INV_0  ( .I(\SB1_3_27/buf_output[0] ), .ZN(\SB2_3_22/i3[0] ) );
  INV_X1 \SB2_3_23/INV_4  ( .I(\SB1_3_24/buf_output[4] ), .ZN(\SB2_3_23/i0[7] ) );
  INV_X2 \SB2_3_23/INV_3  ( .I(\SB1_3_25/buf_output[3] ), .ZN(\SB2_3_23/i0[8] ) );
  INV_X1 \SB2_3_23/INV_1  ( .I(\SB1_3_27/buf_output[1] ), .ZN(\SB2_3_23/i1_7 )
         );
  INV_X1 \SB2_3_24/INV_4  ( .I(\SB1_3_25/buf_output[4] ), .ZN(\SB2_3_24/i0[7] ) );
  INV_X1 \SB2_3_25/INV_4  ( .I(\SB1_3_26/buf_output[4] ), .ZN(\SB2_3_25/i0[7] ) );
  INV_X2 \SB2_3_26/INV_3  ( .I(\SB1_3_28/buf_output[3] ), .ZN(\SB2_3_26/i0[8] ) );
  INV_X1 \SB2_3_26/INV_1  ( .I(\SB1_3_30/buf_output[1] ), .ZN(\SB2_3_26/i1_7 )
         );
  INV_X1 \SB2_3_26/INV_0  ( .I(\SB1_3_31/buf_output[0] ), .ZN(\SB2_3_26/i3[0] ) );
  INV_X1 \SB2_3_27/INV_4  ( .I(\SB1_3_28/buf_output[4] ), .ZN(\SB2_3_27/i0[7] ) );
  INV_X1 \SB2_3_27/INV_0  ( .I(\SB1_3_0/buf_output[0] ), .ZN(\SB2_3_27/i3[0] )
         );
  INV_X1 \SB2_3_28/INV_1  ( .I(\SB1_3_0/buf_output[1] ), .ZN(\SB2_3_28/i1_7 )
         );
  INV_X1 \SB2_3_28/INV_0  ( .I(\SB1_3_1/buf_output[0] ), .ZN(\SB2_3_28/i3[0] )
         );
  INV_X1 \SB2_3_29/INV_0  ( .I(\SB1_3_2/buf_output[0] ), .ZN(\SB2_3_29/i3[0] )
         );
  INV_X1 \SB2_3_30/INV_4  ( .I(\SB1_3_31/buf_output[4] ), .ZN(\SB2_3_30/i0[7] ) );
  INV_X1 \SB2_3_30/INV_0  ( .I(\SB1_3_3/buf_output[0] ), .ZN(\SB2_3_30/i3[0] )
         );
  INV_X1 \SB2_3_31/INV_4  ( .I(\SB1_3_0/buf_output[4] ), .ZN(\SB2_3_31/i0[7] )
         );
  INV_X1 \SB2_3_31/INV_0  ( .I(\SB1_3_4/buf_output[0] ), .ZN(\SB2_3_31/i3[0] )
         );
  INV_X1 \SB1_4_0/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[190] ), .ZN(
        \SB1_4_0/i0[7] ) );
  INV_X1 \SB1_4_1/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[184] ), .ZN(
        \SB1_4_1/i0[7] ) );
  INV_X1 \SB1_4_2/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[178] ), .ZN(
        \SB1_4_2/i0[7] ) );
  INV_X2 \SB1_4_2/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[177] ), .ZN(
        \SB1_4_2/i0[8] ) );
  INV_X1 \SB1_4_4/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[166] ), .ZN(
        \SB1_4_4/i0[7] ) );
  INV_X1 \SB1_4_4/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[163] ), .ZN(
        \SB1_4_4/i1_7 ) );
  INV_X1 \SB1_4_4/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[162] ), .ZN(
        \SB1_4_4/i3[0] ) );
  INV_X1 \SB1_4_5/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[160] ), .ZN(
        \SB1_4_5/i0[7] ) );
  INV_X1 \SB1_4_5/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[157] ), .ZN(
        \SB1_4_5/i1_7 ) );
  INV_X1 \SB1_4_5/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[156] ), .ZN(
        \SB1_4_5/i3[0] ) );
  INV_X1 \SB1_4_6/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[154] ), .ZN(
        \SB1_4_6/i0[7] ) );
  INV_X2 \SB1_4_6/INV_3  ( .I(n3967), .ZN(\SB1_4_6/i0[8] ) );
  INV_X1 \SB1_4_7/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[148] ), .ZN(
        \SB1_4_7/i0[7] ) );
  INV_X1 \SB1_4_7/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[145] ), .ZN(
        \SB1_4_7/i1_7 ) );
  INV_X1 \SB1_4_7/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[144] ), .ZN(
        \SB1_4_7/i3[0] ) );
  INV_X1 \SB1_4_8/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[142] ), .ZN(
        \SB1_4_8/i0[7] ) );
  INV_X1 \SB1_4_8/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[139] ), .ZN(
        \SB1_4_8/i1_7 ) );
  INV_X1 \SB1_4_9/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[136] ), .ZN(
        \SB1_4_9/i0[7] ) );
  INV_X1 \SB1_4_10/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[130] ), .ZN(
        \SB1_4_10/i0[7] ) );
  INV_X1 \SB1_4_10/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[127] ), .ZN(
        \SB1_4_10/i1_7 ) );
  INV_X1 \SB1_4_10/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[126] ), .ZN(
        \SB1_4_10/i3[0] ) );
  INV_X1 \SB1_4_11/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[124] ), .ZN(
        \SB1_4_11/i0[7] ) );
  INV_X1 \SB1_4_11/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[121] ), .ZN(
        \SB1_4_11/i1_7 ) );
  INV_X1 \SB1_4_12/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[118] ), .ZN(
        \SB1_4_12/i0[7] ) );
  INV_X2 \SB1_4_12/INV_3  ( .I(n3975), .ZN(\SB1_4_12/i0[8] ) );
  INV_X1 \SB1_4_12/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[114] ), .ZN(
        \SB1_4_12/i3[0] ) );
  INV_X1 \SB1_4_13/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[112] ), .ZN(
        \SB1_4_13/i0[7] ) );
  INV_X1 \SB1_4_13/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[108] ), .ZN(
        \SB1_4_13/i3[0] ) );
  INV_X1 \SB1_4_14/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[106] ), .ZN(
        \SB1_4_14/i0[7] ) );
  INV_X2 \SB1_4_15/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[98] ), .ZN(
        \SB1_4_15/i1[9] ) );
  INV_X1 \SB1_4_16/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[94] ), .ZN(
        \SB1_4_16/i0[7] ) );
  INV_X1 \SB1_4_17/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[88] ), .ZN(
        \SB1_4_17/i0[7] ) );
  INV_X1 \SB1_4_18/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[82] ), .ZN(
        \SB1_4_18/i0[7] ) );
  INV_X1 \SB1_4_20/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[70] ), .ZN(
        \SB1_4_20/i0[7] ) );
  INV_X1 \SB1_4_21/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[64] ), .ZN(
        \SB1_4_21/i0[7] ) );
  INV_X1 \SB1_4_21/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[60] ), .ZN(
        \SB1_4_21/i3[0] ) );
  INV_X1 \SB1_4_22/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[58] ), .ZN(
        \SB1_4_22/i0[7] ) );
  INV_X1 \SB1_4_23/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[52] ), .ZN(
        \SB1_4_23/i0[7] ) );
  INV_X2 \SB1_4_23/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[51] ), .ZN(
        \SB1_4_23/i0[8] ) );
  INV_X1 \SB1_4_24/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[46] ), .ZN(
        \SB1_4_24/i0[7] ) );
  INV_X1 \SB1_4_25/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[40] ), .ZN(
        \SB1_4_25/i0[7] ) );
  INV_X1 \SB1_4_26/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[34] ), .ZN(
        \SB1_4_26/i0[7] ) );
  INV_X1 \SB1_4_27/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[28] ), .ZN(
        \SB1_4_27/i0[7] ) );
  INV_X2 \SB1_4_27/INV_3  ( .I(n6275), .ZN(\SB1_4_27/i0[8] ) );
  INV_X1 \SB1_4_28/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[22] ), .ZN(
        \SB1_4_28/i0[7] ) );
  INV_X2 \SB1_4_28/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[20] ), .ZN(
        \SB1_4_28/i1[9] ) );
  INV_X1 \SB1_4_29/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[16] ), .ZN(
        \SB1_4_29/i0[7] ) );
  INV_X1 \SB1_4_30/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[6] ), .ZN(
        \SB1_4_30/i3[0] ) );
  INV_X1 \SB1_4_31/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[4] ), .ZN(
        \SB1_4_31/i0[7] ) );
  INV_X1 \SB2_4_0/INV_4  ( .I(\SB1_4_1/buf_output[4] ), .ZN(\SB2_4_0/i0[7] )
         );
  INV_X2 \SB2_4_0/INV_3  ( .I(\SB1_4_2/buf_output[3] ), .ZN(\SB2_4_0/i0[8] )
         );
  INV_X1 \SB2_4_1/INV_0  ( .I(\SB1_4_6/buf_output[0] ), .ZN(\SB2_4_1/i3[0] )
         );
  INV_X1 \SB2_4_2/INV_4  ( .I(\SB1_4_3/buf_output[4] ), .ZN(\SB2_4_2/i0[7] )
         );
  INV_X1 \SB2_4_2/INV_0  ( .I(\SB1_4_7/buf_output[0] ), .ZN(\SB2_4_2/i3[0] )
         );
  INV_X1 \SB2_4_3/INV_4  ( .I(\SB1_4_4/buf_output[4] ), .ZN(\SB2_4_3/i0[7] )
         );
  INV_X1 \SB2_4_3/INV_0  ( .I(\SB1_4_8/buf_output[0] ), .ZN(\SB2_4_3/i3[0] )
         );
  INV_X1 \SB2_4_4/INV_4  ( .I(\SB1_4_5/buf_output[4] ), .ZN(\SB2_4_4/i0[7] )
         );
  INV_X1 \SB2_4_4/INV_0  ( .I(\SB1_4_9/buf_output[0] ), .ZN(\SB2_4_4/i3[0] )
         );
  INV_X1 \SB2_4_5/INV_0  ( .I(\SB1_4_10/buf_output[0] ), .ZN(\SB2_4_5/i3[0] )
         );
  INV_X1 \SB2_4_6/INV_4  ( .I(\SB1_4_7/buf_output[4] ), .ZN(\SB2_4_6/i0[7] )
         );
  INV_X2 \SB2_4_6/INV_3  ( .I(\SB1_4_8/buf_output[3] ), .ZN(\SB2_4_6/i0[8] )
         );
  INV_X1 \SB2_4_6/INV_0  ( .I(\SB1_4_11/buf_output[0] ), .ZN(\SB2_4_6/i3[0] )
         );
  INV_X1 \SB2_4_7/INV_4  ( .I(\SB1_4_8/buf_output[4] ), .ZN(\SB2_4_7/i0[7] )
         );
  INV_X1 \SB2_4_7/INV_0  ( .I(\SB1_4_12/buf_output[0] ), .ZN(\SB2_4_7/i3[0] )
         );
  INV_X2 \SB2_4_8/INV_3  ( .I(\SB1_4_10/buf_output[3] ), .ZN(\SB2_4_8/i0[8] )
         );
  INV_X2 \SB2_4_8/INV_2  ( .I(\SB1_4_11/buf_output[2] ), .ZN(\SB2_4_8/i1[9] )
         );
  INV_X1 \SB2_4_8/INV_0  ( .I(\SB1_4_13/buf_output[0] ), .ZN(\SB2_4_8/i3[0] )
         );
  INV_X1 \SB2_4_9/INV_4  ( .I(\SB1_4_10/buf_output[4] ), .ZN(\SB2_4_9/i0[7] )
         );
  INV_X1 \SB2_4_10/INV_4  ( .I(\SB1_4_11/buf_output[4] ), .ZN(\SB2_4_10/i0[7] ) );
  INV_X1 \SB2_4_10/INV_0  ( .I(\SB1_4_15/buf_output[0] ), .ZN(\SB2_4_10/i3[0] ) );
  INV_X1 \SB2_4_11/INV_4  ( .I(\SB1_4_12/buf_output[4] ), .ZN(\SB2_4_11/i0[7] ) );
  INV_X2 \SB2_4_11/INV_3  ( .I(\SB1_4_13/buf_output[3] ), .ZN(\SB2_4_11/i0[8] ) );
  INV_X1 \SB2_4_13/INV_4  ( .I(\SB1_4_14/buf_output[4] ), .ZN(\SB2_4_13/i0[7] ) );
  INV_X1 \SB2_4_13/INV_0  ( .I(\SB1_4_18/buf_output[0] ), .ZN(\SB2_4_13/i3[0] ) );
  INV_X1 \SB2_4_14/INV_4  ( .I(\SB1_4_15/buf_output[4] ), .ZN(\SB2_4_14/i0[7] ) );
  INV_X1 \SB2_4_15/INV_4  ( .I(\SB1_4_16/buf_output[4] ), .ZN(\SB2_4_15/i0[7] ) );
  INV_X2 \SB2_4_15/INV_3  ( .I(\SB1_4_17/buf_output[3] ), .ZN(\SB2_4_15/i0[8] ) );
  INV_X2 \SB2_4_15/INV_2  ( .I(\SB1_4_18/buf_output[2] ), .ZN(\SB2_4_15/i1[9] ) );
  INV_X1 \SB2_4_15/INV_0  ( .I(\SB1_4_20/buf_output[0] ), .ZN(\SB2_4_15/i3[0] ) );
  INV_X1 \SB2_4_16/INV_4  ( .I(\SB1_4_17/buf_output[4] ), .ZN(\SB2_4_16/i0[7] ) );
  INV_X1 \SB2_4_16/INV_0  ( .I(\SB1_4_21/buf_output[0] ), .ZN(\SB2_4_16/i3[0] ) );
  INV_X1 \SB2_4_17/INV_4  ( .I(\SB1_4_18/buf_output[4] ), .ZN(\SB2_4_17/i0[7] ) );
  INV_X1 \SB2_4_17/INV_0  ( .I(\SB1_4_22/buf_output[0] ), .ZN(\SB2_4_17/i3[0] ) );
  INV_X1 \SB2_4_18/INV_4  ( .I(\SB1_4_19/buf_output[4] ), .ZN(\SB2_4_18/i0[7] ) );
  INV_X1 \SB2_4_18/INV_0  ( .I(\SB1_4_23/buf_output[0] ), .ZN(\SB2_4_18/i3[0] ) );
  INV_X1 \SB2_4_19/INV_4  ( .I(\SB1_4_20/buf_output[4] ), .ZN(\SB2_4_19/i0[7] ) );
  INV_X1 \SB2_4_19/INV_0  ( .I(\SB1_4_24/buf_output[0] ), .ZN(\SB2_4_19/i3[0] ) );
  INV_X1 \SB2_4_21/INV_4  ( .I(\SB1_4_22/buf_output[4] ), .ZN(\SB2_4_21/i0[7] ) );
  INV_X1 \SB2_4_21/INV_0  ( .I(\SB1_4_26/buf_output[0] ), .ZN(\SB2_4_21/i3[0] ) );
  INV_X1 \SB2_4_22/INV_4  ( .I(\SB1_4_23/buf_output[4] ), .ZN(\SB2_4_22/i0[7] ) );
  INV_X1 \SB2_4_22/INV_1  ( .I(\SB1_4_26/buf_output[1] ), .ZN(\SB2_4_22/i1_7 )
         );
  INV_X1 \SB2_4_22/INV_0  ( .I(\SB1_4_27/buf_output[0] ), .ZN(\SB2_4_22/i3[0] ) );
  INV_X1 \SB2_4_23/INV_4  ( .I(\SB1_4_24/buf_output[4] ), .ZN(\SB2_4_23/i0[7] ) );
  INV_X1 \SB2_4_23/INV_0  ( .I(\SB1_4_28/buf_output[0] ), .ZN(\SB2_4_23/i3[0] ) );
  INV_X1 \SB2_4_24/INV_4  ( .I(\SB1_4_25/buf_output[4] ), .ZN(\SB2_4_24/i0[7] ) );
  INV_X2 \SB2_4_24/INV_3  ( .I(\SB1_4_26/buf_output[3] ), .ZN(\SB2_4_24/i0[8] ) );
  INV_X1 \SB2_4_24/INV_0  ( .I(\SB1_4_29/buf_output[0] ), .ZN(\SB2_4_24/i3[0] ) );
  INV_X1 \SB2_4_25/INV_4  ( .I(\SB1_4_26/buf_output[4] ), .ZN(\SB2_4_25/i0[7] ) );
  INV_X1 \SB2_4_25/INV_0  ( .I(\SB1_4_30/buf_output[0] ), .ZN(\SB2_4_25/i3[0] ) );
  INV_X1 \SB2_4_26/INV_4  ( .I(\SB1_4_27/buf_output[4] ), .ZN(\SB2_4_26/i0[7] ) );
  INV_X1 \SB2_4_26/INV_1  ( .I(\SB1_4_30/buf_output[1] ), .ZN(\SB2_4_26/i1_7 )
         );
  INV_X1 \SB2_4_27/INV_4  ( .I(\SB1_4_28/buf_output[4] ), .ZN(\SB2_4_27/i0[7] ) );
  INV_X1 \SB2_4_27/INV_0  ( .I(\SB1_4_0/buf_output[0] ), .ZN(\SB2_4_27/i3[0] )
         );
  INV_X1 \SB2_4_28/INV_4  ( .I(\SB1_4_29/buf_output[4] ), .ZN(\SB2_4_28/i0[7] ) );
  INV_X1 \SB2_4_28/INV_0  ( .I(\SB1_4_1/buf_output[0] ), .ZN(\SB2_4_28/i3[0] )
         );
  INV_X1 \SB2_4_29/INV_4  ( .I(\SB1_4_30/buf_output[4] ), .ZN(\SB2_4_29/i0[7] ) );
  INV_X1 \SB2_4_29/INV_0  ( .I(\SB1_4_2/buf_output[0] ), .ZN(\SB2_4_29/i3[0] )
         );
  INV_X1 \SB2_4_31/INV_0  ( .I(\SB1_4_4/buf_output[0] ), .ZN(\SB2_4_31/i3[0] )
         );
  INV_X1 \SB3_0/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[190] ), .ZN(
        \SB3_0/i0[7] ) );
  INV_X1 \SB3_1/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[184] ), .ZN(
        \SB3_1/i0[7] ) );
  INV_X2 \SB3_1/INV_3  ( .I(\MC_ARK_ARC_1_4/buf_output[183] ), .ZN(
        \SB3_1/i0[8] ) );
  INV_X1 \SB3_1/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[180] ), .ZN(
        \SB3_1/i3[0] ) );
  INV_X1 \SB3_2/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[178] ), .ZN(
        \SB3_2/i0[7] ) );
  INV_X2 \SB3_2/INV_3  ( .I(\MC_ARK_ARC_1_4/buf_output[177] ), .ZN(
        \SB3_2/i0[8] ) );
  INV_X1 \SB3_3/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[172] ), .ZN(
        \SB3_3/i0[7] ) );
  INV_X1 \SB3_3/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[168] ), .ZN(
        \SB3_3/i3[0] ) );
  INV_X1 \SB3_4/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[166] ), .ZN(
        \SB3_4/i0[7] ) );
  INV_X1 \SB3_4/INV_1  ( .I(\MC_ARK_ARC_1_4/buf_output[163] ), .ZN(
        \SB3_4/i1_7 ) );
  INV_X1 \SB3_4/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[162] ), .ZN(
        \SB3_4/i3[0] ) );
  INV_X1 \SB3_5/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[160] ), .ZN(
        \SB3_5/i0[7] ) );
  INV_X1 \SB3_5/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[156] ), .ZN(
        \SB3_5/i3[0] ) );
  INV_X1 \SB3_6/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[154] ), .ZN(
        \SB3_6/i0[7] ) );
  INV_X1 \SB3_7/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[148] ), .ZN(
        \SB3_7/i0[7] ) );
  INV_X1 \SB3_8/INV_5  ( .I(\MC_ARK_ARC_1_4/buf_output[143] ), .ZN(
        \SB3_8/i1_5 ) );
  INV_X1 \SB3_8/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[142] ), .ZN(
        \SB3_8/i0[7] ) );
  INV_X1 \SB3_8/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[138] ), .ZN(
        \SB3_8/i3[0] ) );
  INV_X1 \SB3_9/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[136] ), .ZN(
        \SB3_9/i0[7] ) );
  INV_X1 \SB3_9/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[132] ), .ZN(
        \SB3_9/i3[0] ) );
  INV_X1 \SB3_10/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[130] ), .ZN(
        \SB3_10/i0[7] ) );
  INV_X1 \SB3_10/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[126] ), .ZN(
        \SB3_10/i3[0] ) );
  INV_X1 \SB3_11/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[124] ), .ZN(
        \SB3_11/i0[7] ) );
  INV_X1 \SB3_12/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[118] ), .ZN(
        \SB3_12/i0[7] ) );
  INV_X1 \SB3_13/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[112] ), .ZN(
        \SB3_13/i0[7] ) );
  INV_X1 \SB3_14/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[106] ), .ZN(
        \SB3_14/i0[7] ) );
  INV_X1 \SB3_14/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[102] ), .ZN(
        \SB3_14/i3[0] ) );
  INV_X1 \SB3_15/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[100] ), .ZN(
        \SB3_15/i0[7] ) );
  INV_X1 \SB3_15/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[96] ), .ZN(
        \SB3_15/i3[0] ) );
  INV_X1 \SB3_16/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[94] ), .ZN(
        \SB3_16/i0[7] ) );
  INV_X1 \SB3_16/INV_1  ( .I(\MC_ARK_ARC_1_4/buf_output[91] ), .ZN(
        \SB3_16/i1_7 ) );
  INV_X1 \SB3_17/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[88] ), .ZN(
        \SB3_17/i0[7] ) );
  INV_X1 \SB3_17/INV_1  ( .I(\MC_ARK_ARC_1_4/buf_output[85] ), .ZN(
        \SB3_17/i1_7 ) );
  INV_X1 \SB3_17/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[84] ), .ZN(
        \SB3_17/i3[0] ) );
  INV_X1 \SB3_18/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[82] ), .ZN(
        \SB3_18/i0[7] ) );
  INV_X1 \SB3_18/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[78] ), .ZN(
        \SB3_18/i3[0] ) );
  INV_X1 \SB3_19/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[76] ), .ZN(
        \SB3_19/i0[7] ) );
  INV_X1 \SB3_20/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[70] ), .ZN(
        \SB3_20/i0[7] ) );
  INV_X1 \SB3_21/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[64] ), .ZN(
        \SB3_21/i0[7] ) );
  INV_X1 \SB3_21/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[60] ), .ZN(
        \SB3_21/i3[0] ) );
  INV_X1 \SB3_22/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[58] ), .ZN(
        \SB3_22/i0[7] ) );
  INV_X1 \SB3_22/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[54] ), .ZN(
        \SB3_22/i3[0] ) );
  INV_X1 \SB3_23/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[52] ), .ZN(
        \SB3_23/i0[7] ) );
  INV_X1 \SB3_23/INV_1  ( .I(\MC_ARK_ARC_1_4/buf_output[49] ), .ZN(
        \SB3_23/i1_7 ) );
  INV_X1 \SB3_24/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[46] ), .ZN(
        \SB3_24/i0[7] ) );
  INV_X1 \SB3_24/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[42] ), .ZN(
        \SB3_24/i3[0] ) );
  INV_X1 \SB3_25/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[40] ), .ZN(
        \SB3_25/i0[7] ) );
  INV_X1 \SB3_26/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[34] ), .ZN(
        \SB3_26/i0[7] ) );
  INV_X1 \SB3_26/INV_1  ( .I(\MC_ARK_ARC_1_4/buf_output[31] ), .ZN(
        \SB3_26/i1_7 ) );
  INV_X1 \SB3_27/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[28] ), .ZN(
        \SB3_27/i0[7] ) );
  INV_X2 \SB3_27/INV_3  ( .I(\MC_ARK_ARC_1_4/buf_output[27] ), .ZN(
        \SB3_27/i0[8] ) );
  INV_X1 \SB3_27/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[24] ), .ZN(
        \SB3_27/i3[0] ) );
  INV_X1 \SB3_28/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[22] ), .ZN(
        \SB3_28/i0[7] ) );
  INV_X1 \SB3_29/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[16] ), .ZN(
        \SB3_29/i0[7] ) );
  INV_X1 \SB3_29/INV_1  ( .I(\MC_ARK_ARC_1_4/buf_output[13] ), .ZN(
        \SB3_29/i1_7 ) );
  INV_X1 \SB3_29/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[12] ), .ZN(
        \SB3_29/i3[0] ) );
  INV_X1 \SB3_30/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[10] ), .ZN(
        \SB3_30/i0[7] ) );
  INV_X2 \SB3_30/INV_3  ( .I(\MC_ARK_ARC_1_4/buf_output[9] ), .ZN(
        \SB3_30/i0[8] ) );
  INV_X1 \SB3_30/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[6] ), .ZN(
        \SB3_30/i3[0] ) );
  INV_X1 \SB3_31/INV_4  ( .I(\MC_ARK_ARC_1_4/buf_output[4] ), .ZN(
        \SB3_31/i0[7] ) );
  INV_X1 \SB4_0/INV_4  ( .I(\SB3_1/buf_output[4] ), .ZN(\SB4_0/i0[7] ) );
  INV_X1 \SB4_0/INV_0  ( .I(\SB3_5/buf_output[0] ), .ZN(\SB4_0/i3[0] ) );
  INV_X1 \SB4_1/INV_4  ( .I(\SB3_2/buf_output[4] ), .ZN(\SB4_1/i0[7] ) );
  INV_X1 \SB4_1/INV_0  ( .I(\SB3_6/buf_output[0] ), .ZN(\SB4_1/i3[0] ) );
  INV_X1 \SB4_2/INV_4  ( .I(\SB3_3/buf_output[4] ), .ZN(\SB4_2/i0[7] ) );
  INV_X1 \SB4_2/INV_0  ( .I(\SB3_7/buf_output[0] ), .ZN(\SB4_2/i3[0] ) );
  INV_X1 \SB4_3/INV_4  ( .I(\SB3_4/buf_output[4] ), .ZN(\SB4_3/i0[7] ) );
  INV_X1 \SB4_3/INV_0  ( .I(\SB3_8/buf_output[0] ), .ZN(\SB4_3/i3[0] ) );
  INV_X1 \SB4_4/INV_4  ( .I(\SB3_5/buf_output[4] ), .ZN(\SB4_4/i0[7] ) );
  INV_X2 \SB4_4/INV_3  ( .I(\SB3_6/buf_output[3] ), .ZN(\SB4_4/i0[8] ) );
  INV_X1 \SB4_4/INV_1  ( .I(\SB3_8/buf_output[1] ), .ZN(\SB4_4/i1_7 ) );
  INV_X1 \SB4_4/INV_0  ( .I(\SB3_9/buf_output[0] ), .ZN(\SB4_4/i3[0] ) );
  INV_X1 \SB4_5/INV_4  ( .I(\SB3_6/buf_output[4] ), .ZN(\SB4_5/i0[7] ) );
  INV_X1 \SB4_5/INV_1  ( .I(\SB3_9/buf_output[1] ), .ZN(\SB4_5/i1_7 ) );
  INV_X1 \SB4_5/INV_0  ( .I(\SB3_10/buf_output[0] ), .ZN(\SB4_5/i3[0] ) );
  INV_X1 \SB4_6/INV_4  ( .I(\SB3_7/buf_output[4] ), .ZN(\SB4_6/i0[7] ) );
  INV_X1 \SB4_6/INV_1  ( .I(\SB3_10/buf_output[1] ), .ZN(\SB4_6/i1_7 ) );
  INV_X1 \SB4_7/INV_4  ( .I(\SB3_8/buf_output[4] ), .ZN(\SB4_7/i0[7] ) );
  INV_X1 \SB4_7/INV_0  ( .I(\SB3_12/buf_output[0] ), .ZN(\SB4_7/i3[0] ) );
  INV_X1 \SB4_8/INV_4  ( .I(\SB3_9/buf_output[4] ), .ZN(\SB4_8/i0[7] ) );
  INV_X1 \SB4_8/INV_0  ( .I(\SB3_13/buf_output[0] ), .ZN(\SB4_8/i3[0] ) );
  INV_X1 \SB4_9/INV_4  ( .I(\SB3_10/buf_output[4] ), .ZN(\SB4_9/i0[7] ) );
  INV_X1 \SB4_9/INV_0  ( .I(\SB3_14/buf_output[0] ), .ZN(\SB4_9/i3[0] ) );
  INV_X1 \SB4_10/INV_4  ( .I(\SB3_11/buf_output[4] ), .ZN(\SB4_10/i0[7] ) );
  INV_X1 \SB4_11/INV_4  ( .I(\SB3_12/buf_output[4] ), .ZN(\SB4_11/i0[7] ) );
  INV_X1 \SB4_12/INV_4  ( .I(\SB3_13/buf_output[4] ), .ZN(\SB4_12/i0[7] ) );
  INV_X1 \SB4_12/INV_1  ( .I(\SB3_16/buf_output[1] ), .ZN(\SB4_12/i1_7 ) );
  INV_X1 \SB4_12/INV_0  ( .I(\SB3_17/buf_output[0] ), .ZN(\SB4_12/i3[0] ) );
  INV_X1 \SB4_13/INV_4  ( .I(\SB3_14/buf_output[4] ), .ZN(\SB4_13/i0[7] ) );
  INV_X1 \SB4_14/INV_4  ( .I(\SB3_15/buf_output[4] ), .ZN(\SB4_14/i0[7] ) );
  INV_X1 \SB4_14/INV_1  ( .I(\SB3_18/buf_output[1] ), .ZN(\SB4_14/i1_7 ) );
  INV_X1 \SB4_14/INV_0  ( .I(\SB3_19/buf_output[0] ), .ZN(\SB4_14/i3[0] ) );
  INV_X1 \SB4_15/INV_4  ( .I(\SB3_16/buf_output[4] ), .ZN(\SB4_15/i0[7] ) );
  INV_X1 \SB4_15/INV_0  ( .I(\SB3_20/buf_output[0] ), .ZN(\SB4_15/i3[0] ) );
  INV_X1 \SB4_16/INV_4  ( .I(\SB3_17/buf_output[4] ), .ZN(\SB4_16/i0[7] ) );
  INV_X1 \SB4_16/INV_0  ( .I(\SB3_21/buf_output[0] ), .ZN(\SB4_16/i3[0] ) );
  INV_X1 \SB4_17/INV_4  ( .I(\SB3_18/buf_output[4] ), .ZN(\SB4_17/i0[7] ) );
  INV_X1 \SB4_17/INV_1  ( .I(\SB3_21/buf_output[1] ), .ZN(\SB4_17/i1_7 ) );
  INV_X1 \SB4_17/INV_0  ( .I(\SB3_22/buf_output[0] ), .ZN(\SB4_17/i3[0] ) );
  INV_X1 \SB4_18/INV_4  ( .I(\SB3_19/buf_output[4] ), .ZN(\SB4_18/i0[7] ) );
  INV_X1 \SB4_18/INV_1  ( .I(\SB3_22/buf_output[1] ), .ZN(\SB4_18/i1_7 ) );
  INV_X1 \SB4_18/INV_0  ( .I(\SB3_23/buf_output[0] ), .ZN(\SB4_18/i3[0] ) );
  INV_X1 \SB4_19/INV_4  ( .I(\SB3_20/buf_output[4] ), .ZN(\SB4_19/i0[7] ) );
  INV_X1 \SB4_19/INV_1  ( .I(\RI3[5][73] ), .ZN(\SB4_19/i1_7 ) );
  INV_X1 \SB4_19/INV_0  ( .I(\SB3_24/buf_output[0] ), .ZN(\SB4_19/i3[0] ) );
  INV_X1 \SB4_20/INV_4  ( .I(\SB3_21/buf_output[4] ), .ZN(\SB4_20/i0[7] ) );
  INV_X1 \SB4_21/INV_4  ( .I(\SB3_22/buf_output[4] ), .ZN(\SB4_21/i0[7] ) );
  INV_X2 \SB4_21/INV_3  ( .I(\SB3_23/buf_output[3] ), .ZN(\SB4_21/i0[8] ) );
  INV_X1 \SB4_22/INV_4  ( .I(\SB3_23/buf_output[4] ), .ZN(\SB4_22/i0[7] ) );
  INV_X1 \SB4_22/INV_0  ( .I(\SB3_27/buf_output[0] ), .ZN(\SB4_22/i3[0] ) );
  INV_X1 \SB4_23/INV_5  ( .I(\SB3_23/buf_output[5] ), .ZN(\SB4_23/i1_5 ) );
  INV_X1 \SB4_23/INV_4  ( .I(\SB3_24/buf_output[4] ), .ZN(\SB4_23/i0[7] ) );
  INV_X1 \SB4_24/INV_4  ( .I(\SB3_25/buf_output[4] ), .ZN(\SB4_24/i0[7] ) );
  INV_X1 \SB4_25/INV_4  ( .I(\SB3_26/buf_output[4] ), .ZN(\SB4_25/i0[7] ) );
  INV_X1 \SB4_25/INV_1  ( .I(\SB3_29/buf_output[1] ), .ZN(\SB4_25/i1_7 ) );
  INV_X1 \SB4_26/INV_4  ( .I(\SB3_27/buf_output[4] ), .ZN(\SB4_26/i0[7] ) );
  INV_X1 \SB4_26/INV_0  ( .I(\SB3_31/buf_output[0] ), .ZN(\SB4_26/i3[0] ) );
  INV_X1 \SB4_27/INV_4  ( .I(\SB3_28/buf_output[4] ), .ZN(\SB4_27/i0[7] ) );
  INV_X1 \SB4_28/INV_4  ( .I(\SB3_29/buf_output[4] ), .ZN(\SB4_28/i0[7] ) );
  INV_X1 \SB4_29/INV_4  ( .I(\SB3_30/buf_output[4] ), .ZN(\SB4_29/i0[7] ) );
  INV_X1 \SB4_29/INV_0  ( .I(\SB3_2/buf_output[0] ), .ZN(\SB4_29/i3[0] ) );
  INV_X1 \SB4_30/INV_4  ( .I(\SB3_31/buf_output[4] ), .ZN(\SB4_30/i0[7] ) );
  INV_X1 \SB4_30/INV_0  ( .I(\SB3_3/buf_output[0] ), .ZN(\SB4_30/i3[0] ) );
  INV_X1 \SB4_31/INV_4  ( .I(\SB3_0/buf_output[4] ), .ZN(\SB4_31/i0[7] ) );
  INV_X1 \SB4_31/INV_0  ( .I(\SB3_4/buf_output[0] ), .ZN(\SB4_31/i3[0] ) );
  NAND3_X1 \SB1_0_0/Component_Function_3/N4  ( .A1(\SB1_0_0/i1_5 ), .A2(
        \SB1_0_0/i0[8] ), .A3(\SB1_0_0/i3[0] ), .ZN(
        \SB1_0_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_4/N2  ( .A1(\SB1_0_0/i3[0] ), .A2(
        \SB1_0_0/i0_0 ), .A3(\SB1_0_0/i1_7 ), .ZN(
        \SB1_0_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_1/Component_Function_2/N1  ( .A1(\SB1_0_1/i1_5 ), .A2(
        \SB1_0_1/i0[10] ), .A3(\SB1_0_1/i1[9] ), .ZN(
        \SB1_0_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_4/N1  ( .A1(\SB1_0_1/i0[9] ), .A2(
        \SB1_0_1/i0_0 ), .A3(\SB1_0_1/i0[8] ), .ZN(
        \SB1_0_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_2/Component_Function_2/N2  ( .A1(\SB1_0_2/i0_3 ), .A2(
        \SB1_0_2/i0[10] ), .A3(\SB1_0_2/i0[6] ), .ZN(
        \SB1_0_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_2/Component_Function_4/N4  ( .A1(\SB1_0_2/i1[9] ), .A2(
        \SB1_0_2/i1_5 ), .A3(\SB1_0_2/i0_4 ), .ZN(
        \SB1_0_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_2/Component_Function_4/N2  ( .A1(\SB1_0_2/i3[0] ), .A2(
        \SB1_0_2/i0_0 ), .A3(\SB1_0_2/i1_7 ), .ZN(
        \SB1_0_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_3/Component_Function_2/N3  ( .A1(\SB1_0_3/i0_3 ), .A2(
        \SB1_0_3/i0[8] ), .A3(\SB1_0_3/i0[9] ), .ZN(
        \SB1_0_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_3/Component_Function_3/N4  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0[8] ), .A3(\SB1_0_3/i3[0] ), .ZN(
        \SB1_0_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_3/N1  ( .A1(\SB1_0_3/i1[9] ), .A2(
        \SB1_0_3/i0_3 ), .A3(\SB1_0_3/i0[6] ), .ZN(
        \SB1_0_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_4/N4  ( .A1(\SB1_0_3/i1[9] ), .A2(
        \SB1_0_3/i1_5 ), .A3(n374), .ZN(
        \SB1_0_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_4/N3  ( .A1(\SB1_0_3/i0[9] ), .A2(
        \SB1_0_3/i0[10] ), .A3(\SB1_0_3/i0_3 ), .ZN(
        \SB1_0_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_3/Component_Function_4/N1  ( .A1(\SB1_0_3/i0[9] ), .A2(
        \SB1_0_3/i0_0 ), .A3(\SB1_0_3/i0[8] ), .ZN(
        \SB1_0_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_2/N2  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i0[10] ), .A3(\SB1_0_4/i0[6] ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_4/Component_Function_3/N4  ( .A1(\SB1_0_4/i1_5 ), .A2(
        \SB1_0_4/i0[8] ), .A3(\SB1_0_4/i3[0] ), .ZN(
        \SB1_0_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N3  ( .A1(\SB1_0_4/i0[9] ), .A2(
        \SB1_0_4/i0[10] ), .A3(\SB1_0_4/i0_3 ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N2  ( .A1(\SB1_0_4/i3[0] ), .A2(
        \SB1_0_4/i0_0 ), .A3(\SB1_0_4/i1_7 ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N1  ( .A1(\SB1_0_4/i0[9] ), .A2(
        \SB1_0_4/i0_0 ), .A3(\SB1_0_4/i0[8] ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_3/N4  ( .A1(\SB1_0_5/i1_5 ), .A2(
        \SB1_0_5/i0[8] ), .A3(\SB1_0_5/i3[0] ), .ZN(
        \SB1_0_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_5/Component_Function_4/N2  ( .A1(\SB1_0_5/i3[0] ), .A2(
        \SB1_0_5/i0_0 ), .A3(\SB1_0_5/i1_7 ), .ZN(
        \SB1_0_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_5/Component_Function_4/N1  ( .A1(\SB1_0_5/i0[9] ), .A2(
        \SB1_0_5/i0_0 ), .A3(\SB1_0_5/i0[8] ), .ZN(
        \SB1_0_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_3/N4  ( .A1(\SB1_0_6/i1_5 ), .A2(
        \SB1_0_6/i0[8] ), .A3(\SB1_0_6/i3[0] ), .ZN(
        \SB1_0_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_4/N4  ( .A1(\SB1_0_6/i1[9] ), .A2(
        \SB1_0_6/i1_5 ), .A3(\SB1_0_6/i0_4 ), .ZN(
        \SB1_0_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_3/N1  ( .A1(\SB1_0_7/i1[9] ), .A2(
        \SB1_0_7/i0_3 ), .A3(\SB1_0_7/i0[6] ), .ZN(
        \SB1_0_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_3/N4  ( .A1(\SB1_0_8/i1_5 ), .A2(
        \SB1_0_8/i0[8] ), .A3(\SB1_0_8/i3[0] ), .ZN(
        \SB1_0_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_8/Component_Function_4/N2  ( .A1(\SB1_0_8/i3[0] ), .A2(
        \SB1_0_8/i0_0 ), .A3(\SB1_0_8/i1_7 ), .ZN(
        \SB1_0_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_8/Component_Function_4/N1  ( .A1(\SB1_0_8/i0[9] ), .A2(
        \SB1_0_8/i0_0 ), .A3(\SB1_0_8/i0[8] ), .ZN(
        \SB1_0_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_2/N1  ( .A1(\SB1_0_9/i1_5 ), .A2(
        \SB1_0_9/i0[10] ), .A3(\SB1_0_9/i1[9] ), .ZN(
        \SB1_0_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_3/N4  ( .A1(\SB1_0_9/i1_5 ), .A2(
        \SB1_0_9/i0[8] ), .A3(\SB1_0_9/i3[0] ), .ZN(
        \SB1_0_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_4/N4  ( .A1(\SB1_0_9/i1[9] ), .A2(
        \SB1_0_9/i1_5 ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_4/N2  ( .A1(\SB1_0_9/i3[0] ), .A2(
        \SB1_0_9/i0_0 ), .A3(\SB1_0_9/i1_7 ), .ZN(
        \SB1_0_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_9/Component_Function_4/N1  ( .A1(\SB1_0_9/i0[9] ), .A2(
        \SB1_0_9/i0_0 ), .A3(\SB1_0_9/i0[8] ), .ZN(
        \SB1_0_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_2/N3  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i0[8] ), .A3(\SB1_0_11/i0[9] ), .ZN(
        \SB1_0_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_3/N4  ( .A1(\SB1_0_11/i1_5 ), .A2(
        \SB1_0_11/i0[8] ), .A3(\SB1_0_11/i3[0] ), .ZN(
        \SB1_0_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_11/Component_Function_3/N2  ( .A1(\SB1_0_11/i0_0 ), .A2(
        \SB1_0_11/i0_3 ), .A3(\SB1_0_11/i0_4 ), .ZN(
        \SB1_0_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_11/Component_Function_4/N4  ( .A1(\SB1_0_11/i1[9] ), .A2(
        \SB1_0_11/i1_5 ), .A3(\SB1_0_11/i0_4 ), .ZN(
        \SB1_0_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_2/N3  ( .A1(\SB1_0_12/i0_3 ), .A2(
        \SB1_0_12/i0[8] ), .A3(\SB1_0_12/i0[9] ), .ZN(
        \SB1_0_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_12/Component_Function_3/N4  ( .A1(\SB1_0_12/i1_5 ), .A2(
        \SB1_0_12/i0[8] ), .A3(\SB1_0_12/i3[0] ), .ZN(
        \SB1_0_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_3/N1  ( .A1(\SB1_0_12/i1[9] ), .A2(
        \SB1_0_12/i0_3 ), .A3(\SB1_0_12/i0[6] ), .ZN(
        \SB1_0_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_4/N4  ( .A1(\SB1_0_12/i1[9] ), .A2(
        \SB1_0_12/i1_5 ), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_3/N4  ( .A1(\SB1_0_13/i1_5 ), .A2(
        n5428), .A3(\SB1_0_13/i3[0] ), .ZN(
        \SB1_0_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_4/N2  ( .A1(\SB1_0_13/i3[0] ), .A2(
        \SB1_0_13/i0_0 ), .A3(\SB1_0_13/i1_7 ), .ZN(
        \SB1_0_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_14/Component_Function_2/N1  ( .A1(\SB1_0_14/i1_5 ), .A2(
        \SB1_0_14/i0[10] ), .A3(\SB1_0_14/i1[9] ), .ZN(
        \SB1_0_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_4/N2  ( .A1(\SB1_0_14/i3[0] ), .A2(
        \SB1_0_14/i0_0 ), .A3(\SB1_0_14/i1_7 ), .ZN(
        \SB1_0_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_14/Component_Function_4/N1  ( .A1(\SB1_0_14/i0[9] ), .A2(
        \SB1_0_14/i0_0 ), .A3(\SB1_0_14/i0[8] ), .ZN(
        \SB1_0_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_2/N1  ( .A1(\SB1_0_15/i1_5 ), .A2(
        \SB1_0_15/i0[10] ), .A3(\SB1_0_15/i1[9] ), .ZN(
        \SB1_0_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_3/N4  ( .A1(\SB1_0_15/i1_5 ), .A2(
        \SB1_0_15/i0[8] ), .A3(\SB1_0_15/i3[0] ), .ZN(
        \SB1_0_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_3/N3  ( .A1(\SB1_0_15/i1[9] ), .A2(
        \SB1_0_15/i1_7 ), .A3(\SB1_0_15/i0[10] ), .ZN(
        \SB1_0_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_15/Component_Function_4/N4  ( .A1(\SB1_0_15/i1[9] ), .A2(
        \SB1_0_15/i1_5 ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_4/N2  ( .A1(\SB1_0_15/i3[0] ), .A2(
        \SB1_0_15/i0_0 ), .A3(\SB1_0_15/i1_7 ), .ZN(
        \SB1_0_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_16/Component_Function_2/N2  ( .A1(\SB1_0_16/i0_3 ), .A2(
        \SB1_0_16/i0[10] ), .A3(\SB1_0_16/i0[6] ), .ZN(
        \SB1_0_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_16/Component_Function_4/N4  ( .A1(\SB1_0_16/i1[9] ), .A2(
        \SB1_0_16/i1_5 ), .A3(\SB1_0_16/i0_4 ), .ZN(
        \SB1_0_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_16/Component_Function_4/N2  ( .A1(\SB1_0_16/i3[0] ), .A2(
        \SB1_0_16/i0_0 ), .A3(\SB1_0_16/i1_7 ), .ZN(
        \SB1_0_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_17/Component_Function_2/N3  ( .A1(\SB1_0_17/i0_3 ), .A2(
        \SB1_0_17/i0[8] ), .A3(\SB1_0_17/i0[9] ), .ZN(
        \SB1_0_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_17/Component_Function_3/N4  ( .A1(\SB1_0_17/i1_5 ), .A2(
        \SB1_0_17/i0[8] ), .A3(\SB1_0_17/i3[0] ), .ZN(
        \SB1_0_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_3/N2  ( .A1(\SB1_0_17/i0_0 ), .A2(
        \SB1_0_17/i0_3 ), .A3(\SB1_0_17/i0_4 ), .ZN(
        \SB1_0_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_17/Component_Function_3/N1  ( .A1(\SB1_0_17/i1[9] ), .A2(
        \SB1_0_17/i0_3 ), .A3(\SB1_0_17/i0[6] ), .ZN(
        \SB1_0_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_17/Component_Function_4/N4  ( .A1(\SB1_0_17/i1[9] ), .A2(
        \SB1_0_17/i1_5 ), .A3(\SB1_0_17/i0_4 ), .ZN(
        \SB1_0_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_4/N1  ( .A1(\SB1_0_17/i0[9] ), .A2(
        \SB1_0_17/i0_0 ), .A3(\SB1_0_17/i0[8] ), .ZN(
        \SB1_0_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_2/N2  ( .A1(\SB1_0_18/i0_3 ), .A2(
        \SB1_0_18/i0[10] ), .A3(\SB1_0_18/i0[6] ), .ZN(
        \SB1_0_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_18/Component_Function_2/N1  ( .A1(\SB1_0_18/i1_5 ), .A2(
        \SB1_0_18/i0[10] ), .A3(\SB1_0_18/i1[9] ), .ZN(
        \SB1_0_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_4/N4  ( .A1(\SB1_0_18/i1[9] ), .A2(
        \SB1_0_18/i1_5 ), .A3(\SB1_0_18/i0_4 ), .ZN(
        \SB1_0_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_18/Component_Function_4/N2  ( .A1(\SB1_0_18/i3[0] ), .A2(
        n6290), .A3(\SB1_0_18/i1_7 ), .ZN(
        \SB1_0_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_19/Component_Function_2/N1  ( .A1(\SB1_0_19/i1_5 ), .A2(
        \SB1_0_19/i0[10] ), .A3(\SB1_0_19/i1[9] ), .ZN(
        \SB1_0_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_19/Component_Function_3/N3  ( .A1(\SB1_0_19/i1[9] ), .A2(
        \SB1_0_19/i1_7 ), .A3(\SB1_0_19/i0[10] ), .ZN(
        \SB1_0_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_19/Component_Function_4/N2  ( .A1(\SB1_0_19/i3[0] ), .A2(
        \SB1_0_19/i0_0 ), .A3(\SB1_0_19/i1_7 ), .ZN(
        \SB1_0_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_19/Component_Function_4/N1  ( .A1(\SB1_0_19/i0[9] ), .A2(
        \SB1_0_19/i0_0 ), .A3(\SB1_0_19/i0[8] ), .ZN(
        \SB1_0_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_2/N4  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0_0 ), .A3(\SB1_0_20/i0_4 ), .ZN(
        \SB1_0_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_20/Component_Function_3/N4  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0[8] ), .A3(\SB1_0_20/i3[0] ), .ZN(
        \SB1_0_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_20/Component_Function_4/N4  ( .A1(\SB1_0_20/i1[9] ), .A2(
        \SB1_0_20/i1_5 ), .A3(\SB1_0_20/i0_4 ), .ZN(
        \SB1_0_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_20/Component_Function_4/N2  ( .A1(\SB1_0_20/i3[0] ), .A2(
        \SB1_0_20/i0_0 ), .A3(\SB1_0_20/i1_7 ), .ZN(
        \SB1_0_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_20/Component_Function_4/N1  ( .A1(\SB1_0_20/i0[9] ), .A2(
        \SB1_0_20/i0_0 ), .A3(\SB1_0_20/i0[8] ), .ZN(
        \SB1_0_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_4/N2  ( .A1(\SB1_0_21/i3[0] ), .A2(
        \SB1_0_21/i0_0 ), .A3(\SB1_0_21/i1_7 ), .ZN(
        \SB1_0_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_22/Component_Function_2/N3  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i0[8] ), .A3(\SB1_0_22/i0[9] ), .ZN(
        \SB1_0_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_22/Component_Function_3/N4  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0[8] ), .A3(\SB1_0_22/i3[0] ), .ZN(
        \SB1_0_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_22/Component_Function_3/N3  ( .A1(\SB1_0_22/i1[9] ), .A2(
        \SB1_0_22/i1_7 ), .A3(\SB1_0_22/i0[10] ), .ZN(
        \SB1_0_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_22/Component_Function_4/N2  ( .A1(\SB1_0_22/i3[0] ), .A2(
        \SB1_0_22/i0_0 ), .A3(\SB1_0_22/i1_7 ), .ZN(
        \SB1_0_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_22/Component_Function_4/N1  ( .A1(\SB1_0_22/i0[9] ), .A2(
        \SB1_0_22/i0_0 ), .A3(\SB1_0_22/i0[8] ), .ZN(
        \SB1_0_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_2/N2  ( .A1(\SB1_0_23/i0_3 ), .A2(
        \SB1_0_23/i0[10] ), .A3(\SB1_0_23/i0[6] ), .ZN(
        \SB1_0_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_23/Component_Function_3/N4  ( .A1(\SB1_0_23/i1_5 ), .A2(
        \SB1_0_23/i0[8] ), .A3(\SB1_0_23/i3[0] ), .ZN(
        \SB1_0_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_23/Component_Function_4/N4  ( .A1(\SB1_0_23/i1[9] ), .A2(
        \SB1_0_23/i1_5 ), .A3(\SB1_0_23/i0_4 ), .ZN(
        \SB1_0_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_23/Component_Function_4/N2  ( .A1(\SB1_0_23/i3[0] ), .A2(
        \SB1_0_23/i0_0 ), .A3(\SB1_0_23/i1_7 ), .ZN(
        \SB1_0_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_23/Component_Function_4/N1  ( .A1(\SB1_0_23/i0[9] ), .A2(
        \SB1_0_23/i0_0 ), .A3(\SB1_0_23/i0[8] ), .ZN(
        \SB1_0_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_4/N2  ( .A1(\SB1_0_24/i3[0] ), .A2(
        \SB1_0_24/i0_0 ), .A3(\SB1_0_24/i1_7 ), .ZN(
        \SB1_0_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_25/Component_Function_4/N4  ( .A1(\SB1_0_25/i1[9] ), .A2(
        \SB1_0_25/i1_5 ), .A3(\SB1_0_25/i0_4 ), .ZN(
        \SB1_0_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_25/Component_Function_4/N2  ( .A1(\SB1_0_25/i3[0] ), .A2(
        \SB1_0_25/i0_0 ), .A3(\SB1_0_25/i1_7 ), .ZN(
        \SB1_0_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_25/Component_Function_4/N1  ( .A1(\SB1_0_25/i0[9] ), .A2(
        \SB1_0_25/i0_0 ), .A3(\SB1_0_25/i0[8] ), .ZN(
        \SB1_0_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_2/N1  ( .A1(\SB1_0_26/i1_5 ), .A2(
        \SB1_0_26/i0[10] ), .A3(\SB1_0_26/i1[9] ), .ZN(
        \SB1_0_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_3/N2  ( .A1(\SB1_0_26/i0_0 ), .A2(
        \SB1_0_26/i0_3 ), .A3(\SB1_0_26/i0_4 ), .ZN(
        \SB1_0_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_26/Component_Function_3/N1  ( .A1(\SB1_0_26/i1[9] ), .A2(
        \SB1_0_26/i0_3 ), .A3(\SB1_0_26/i0[6] ), .ZN(
        \SB1_0_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_4/N4  ( .A1(\SB1_0_26/i1[9] ), .A2(
        \SB1_0_26/i1_5 ), .A3(\SB1_0_26/i0_4 ), .ZN(
        \SB1_0_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_4/N3  ( .A1(\SB1_0_26/i0[9] ), .A2(
        \SB1_0_26/i0[10] ), .A3(\SB1_0_26/i0_3 ), .ZN(
        \SB1_0_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_26/Component_Function_4/N2  ( .A1(\SB1_0_26/i3[0] ), .A2(
        \SB1_0_26/i0_0 ), .A3(\SB1_0_26/i1_7 ), .ZN(
        \SB1_0_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_27/Component_Function_2/N4  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0_0 ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_2/N1  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0[10] ), .A3(\SB1_0_27/i1[9] ), .ZN(
        \SB1_0_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_3/N4  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0[8] ), .A3(\SB1_0_27/i3[0] ), .ZN(
        \SB1_0_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_3/N2  ( .A1(\SB1_0_27/i0_0 ), .A2(
        \SB1_0_27/i0_3 ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N4  ( .A1(\SB1_0_27/i1[9] ), .A2(
        \SB1_0_27/i1_5 ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_28/Component_Function_2/N3  ( .A1(\SB1_0_28/i0_3 ), .A2(
        \SB1_0_28/i0[8] ), .A3(\SB1_0_28/i0[9] ), .ZN(
        \SB1_0_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_28/Component_Function_4/N3  ( .A1(\SB1_0_28/i0[9] ), .A2(
        \SB1_0_28/i0[10] ), .A3(\SB1_0_28/i0_3 ), .ZN(
        \SB1_0_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_28/Component_Function_4/N2  ( .A1(\SB1_0_28/i3[0] ), .A2(
        \SB1_0_28/i0_0 ), .A3(\SB1_0_28/i1_7 ), .ZN(
        \SB1_0_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_28/Component_Function_4/N1  ( .A1(\SB1_0_28/i0[9] ), .A2(
        \SB1_0_28/i0_0 ), .A3(\SB1_0_28/i0[8] ), .ZN(
        \SB1_0_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_29/Component_Function_3/N4  ( .A1(\SB1_0_29/i1_5 ), .A2(
        \SB1_0_29/i0[8] ), .A3(\SB1_0_29/i3[0] ), .ZN(
        \SB1_0_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_2/N1  ( .A1(\SB1_0_30/i1_5 ), .A2(
        \SB1_0_30/i0[10] ), .A3(\SB1_0_30/i1[9] ), .ZN(
        \SB1_0_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_3/N4  ( .A1(\SB1_0_30/i1_5 ), .A2(
        \SB1_0_30/i0[8] ), .A3(\SB1_0_30/i3[0] ), .ZN(
        \SB1_0_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_2/N3  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i0[8] ), .A3(\SB1_0_31/i0[9] ), .ZN(
        \SB1_0_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_31/Component_Function_3/N4  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0[8] ), .A3(\SB1_0_31/i3[0] ), .ZN(
        \SB1_0_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_4/N2  ( .A1(\SB1_0_31/i3[0] ), .A2(
        \SB1_0_31/i0_0 ), .A3(\SB1_0_31/i1_7 ), .ZN(
        \SB1_0_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_31/Component_Function_4/N1  ( .A1(\SB1_0_31/i0[9] ), .A2(
        \SB1_0_31/i0_0 ), .A3(\SB1_0_31/i0[8] ), .ZN(
        \SB1_0_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_0/Component_Function_3/N3  ( .A1(\SB2_0_0/i1[9] ), .A2(
        \SB2_0_0/i1_7 ), .A3(\RI3[0][189] ), .ZN(
        \SB2_0_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_0/Component_Function_4/N2  ( .A1(\SB2_0_0/i3[0] ), .A2(
        \SB2_0_0/i0_0 ), .A3(\SB2_0_0/i1_7 ), .ZN(
        \SB2_0_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_1/Component_Function_3/N2  ( .A1(\SB2_0_1/i0_0 ), .A2(
        \SB2_0_1/i0_3 ), .A3(\SB2_0_1/i0_4 ), .ZN(
        \SB2_0_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_1/Component_Function_4/N2  ( .A1(n2592), .A2(\SB2_0_1/i0_0 ), 
        .A3(\SB2_0_1/i1_7 ), .ZN(\SB2_0_1/Component_Function_4/NAND4_in[1] )
         );
  NAND3_X1 \SB2_0_1/Component_Function_4/N1  ( .A1(\SB2_0_1/i0[9] ), .A2(
        \SB2_0_1/i0_0 ), .A3(\SB2_0_1/i0[8] ), .ZN(
        \SB2_0_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_4/N2  ( .A1(\SB2_0_2/i3[0] ), .A2(
        \SB2_0_2/i0_0 ), .A3(\SB2_0_2/i1_7 ), .ZN(
        \SB2_0_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_2/Component_Function_4/N1  ( .A1(\SB2_0_2/i0[9] ), .A2(
        \SB2_0_2/i0_0 ), .A3(\SB2_0_2/i0[8] ), .ZN(
        \SB2_0_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_3/Component_Function_3/N4  ( .A1(\SB2_0_3/i1_5 ), .A2(
        \SB2_0_3/i0[8] ), .A3(\SB2_0_3/i3[0] ), .ZN(
        \SB2_0_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_3/Component_Function_4/N4  ( .A1(\SB2_0_3/i1[9] ), .A2(
        \SB2_0_3/i1_5 ), .A3(\RI3[0][172] ), .ZN(
        \SB2_0_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_3/Component_Function_4/N1  ( .A1(\SB2_0_3/i0[9] ), .A2(
        \SB2_0_3/i0_0 ), .A3(\SB2_0_3/i0[8] ), .ZN(
        \SB2_0_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_4/Component_Function_3/N1  ( .A1(\SB2_0_4/i1[9] ), .A2(
        \SB2_0_4/i0_3 ), .A3(\SB2_0_4/i0[6] ), .ZN(
        \SB2_0_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_4/N2  ( .A1(\SB2_0_5/i3[0] ), .A2(
        \SB2_0_5/i0_0 ), .A3(\SB2_0_5/i1_7 ), .ZN(
        \SB2_0_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_5/Component_Function_4/N1  ( .A1(\SB2_0_5/i0[9] ), .A2(
        \SB2_0_5/i0_0 ), .A3(\SB2_0_5/i0[8] ), .ZN(
        \SB2_0_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_4/N2  ( .A1(\SB2_0_6/i3[0] ), .A2(
        \SB2_0_6/i0_0 ), .A3(\SB2_0_6/i1_7 ), .ZN(
        \SB2_0_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_6/Component_Function_4/N1  ( .A1(\SB2_0_6/i0[9] ), .A2(
        \SB2_0_6/i0_0 ), .A3(\SB2_0_6/i0[8] ), .ZN(
        \SB2_0_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_2/N2  ( .A1(\SB2_0_7/i0_3 ), .A2(
        \SB2_0_7/i0[10] ), .A3(\SB2_0_7/i0[6] ), .ZN(
        \SB2_0_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_7/Component_Function_3/N4  ( .A1(\SB2_0_7/i1_5 ), .A2(
        \SB2_0_7/i0[8] ), .A3(\SB2_0_7/i3[0] ), .ZN(
        \SB2_0_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_8/Component_Function_2/N2  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \RI3[0][141] ), .A3(\SB2_0_8/i0[6] ), .ZN(
        \SB2_0_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_8/Component_Function_4/N4  ( .A1(\SB2_0_8/i1[9] ), .A2(
        \SB2_0_8/i1_5 ), .A3(\RI3[0][142] ), .ZN(
        \SB2_0_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_9/Component_Function_3/N1  ( .A1(\SB2_0_9/i1[9] ), .A2(
        \SB2_0_9/i0_3 ), .A3(\SB2_0_9/i0[6] ), .ZN(
        \SB2_0_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_9/Component_Function_4/N1  ( .A1(\SB2_0_9/i0[9] ), .A2(n2886), .A3(\SB2_0_9/i0[8] ), .ZN(\SB2_0_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_4/N1  ( .A1(\SB2_0_10/i0[9] ), .A2(
        \RI3[0][128] ), .A3(\SB2_0_10/i0[8] ), .ZN(
        \SB2_0_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_2/N3  ( .A1(\SB2_0_11/i0_3 ), .A2(
        \SB2_0_11/i0[8] ), .A3(\SB2_0_11/i0[9] ), .ZN(
        \SB2_0_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_11/Component_Function_3/N4  ( .A1(\SB2_0_11/i1_5 ), .A2(
        \SB2_0_11/i0[8] ), .A3(\SB2_0_11/i3[0] ), .ZN(
        \SB2_0_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_11/Component_Function_4/N1  ( .A1(\SB2_0_11/i0[9] ), .A2(
        \SB2_0_11/i0_0 ), .A3(\SB2_0_11/i0[8] ), .ZN(
        \SB2_0_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_2/N3  ( .A1(\RI3[0][119] ), .A2(
        \SB2_0_12/i0[8] ), .A3(\SB2_0_12/i0[9] ), .ZN(
        \SB2_0_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_12/Component_Function_4/N2  ( .A1(\SB2_0_12/i3[0] ), .A2(
        \SB2_0_12/i0_0 ), .A3(\SB2_0_12/i1_7 ), .ZN(
        \SB2_0_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_12/Component_Function_4/N1  ( .A1(\SB2_0_12/i0[9] ), .A2(
        \SB2_0_12/i0_0 ), .A3(\SB2_0_12/i0[8] ), .ZN(
        \SB2_0_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_2/N2  ( .A1(\SB2_0_13/i0_3 ), .A2(
        \SB2_0_13/i0[10] ), .A3(\SB2_0_13/i0[6] ), .ZN(
        \SB2_0_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_13/Component_Function_4/N2  ( .A1(\SB2_0_13/i3[0] ), .A2(
        \SB2_0_13/i0_0 ), .A3(\SB2_0_13/i1_7 ), .ZN(
        \SB2_0_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_14/Component_Function_2/N2  ( .A1(\SB2_0_14/i0_3 ), .A2(
        \SB2_0_14/i0[10] ), .A3(\SB2_0_14/i0[6] ), .ZN(
        \SB2_0_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_14/Component_Function_3/N2  ( .A1(\SB2_0_14/i0_0 ), .A2(
        \SB2_0_14/i0_3 ), .A3(\SB2_0_14/i0_4 ), .ZN(
        \SB2_0_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_14/Component_Function_3/N1  ( .A1(\SB2_0_14/i1[9] ), .A2(
        \SB2_0_14/i0_3 ), .A3(\SB2_0_14/i0[6] ), .ZN(
        \SB2_0_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_14/Component_Function_4/N1  ( .A1(\SB2_0_14/i0[9] ), .A2(
        \SB2_0_14/i0_0 ), .A3(\SB2_0_14/i0[8] ), .ZN(
        \SB2_0_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_2/N1  ( .A1(\SB2_0_15/i1_5 ), .A2(
        \SB2_0_15/i0[10] ), .A3(n1508), .ZN(
        \SB2_0_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_4/N4  ( .A1(n1508), .A2(
        \SB2_0_15/i1_5 ), .A3(\RI3[0][100] ), .ZN(
        \SB2_0_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_17/Component_Function_3/N4  ( .A1(\SB2_0_17/i1_5 ), .A2(
        \SB2_0_17/i0[8] ), .A3(\SB2_0_17/i3[0] ), .ZN(
        \SB2_0_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_17/Component_Function_4/N2  ( .A1(\SB2_0_17/i3[0] ), .A2(
        \SB2_0_17/i0_0 ), .A3(\SB2_0_17/i1_7 ), .ZN(
        \SB2_0_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_17/Component_Function_4/N1  ( .A1(\SB2_0_17/i0[9] ), .A2(
        \SB2_0_17/i0_0 ), .A3(\SB2_0_17/i0[8] ), .ZN(
        \SB2_0_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_24/Component_Function_2/N3  ( .A1(\SB2_0_24/i0_3 ), .A2(
        \SB2_0_24/i0[8] ), .A3(\SB1_0_29/buf_output[0] ), .ZN(
        \SB2_0_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_3/N3  ( .A1(\SB2_0_24/i1[9] ), .A2(
        \SB2_0_24/i1_7 ), .A3(\SB2_0_24/i0[10] ), .ZN(
        \SB2_0_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_4/N4  ( .A1(\SB2_0_24/i1[9] ), .A2(
        \SB2_0_24/i1_5 ), .A3(\RI3[0][46] ), .ZN(
        \SB2_0_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_24/Component_Function_4/N3  ( .A1(\RI3[0][42] ), .A2(
        \SB2_0_24/i0[10] ), .A3(\SB2_0_24/i0_3 ), .ZN(
        \SB2_0_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_4/N2  ( .A1(\SB2_0_24/i3[0] ), .A2(
        \SB2_0_24/i0_0 ), .A3(\SB2_0_24/i1_7 ), .ZN(
        \SB2_0_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_24/Component_Function_4/N1  ( .A1(\RI3[0][42] ), .A2(
        \SB2_0_24/i0_0 ), .A3(\SB2_0_24/i0[8] ), .ZN(
        \SB2_0_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_2/N2  ( .A1(\SB2_0_26/i0_3 ), .A2(
        \RI3[0][33] ), .A3(\SB1_0_30/buf_output[1] ), .ZN(
        \SB2_0_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_26/Component_Function_3/N1  ( .A1(\SB2_0_26/i1[9] ), .A2(
        \SB2_0_26/i0_3 ), .A3(\SB2_0_26/i0[6] ), .ZN(
        \SB2_0_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_4/N4  ( .A1(\SB2_0_26/i1[9] ), .A2(
        \SB2_0_26/i1_5 ), .A3(\SB2_0_26/i0_4 ), .ZN(
        \SB2_0_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_26/Component_Function_4/N3  ( .A1(\SB2_0_26/i0[9] ), .A2(
        \RI3[0][33] ), .A3(\SB2_0_26/i0_3 ), .ZN(
        \SB2_0_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_27/Component_Function_3/N3  ( .A1(\SB2_0_27/i1[9] ), .A2(
        \SB2_0_27/i1_7 ), .A3(\SB2_0_27/i0[10] ), .ZN(
        \SB2_0_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_27/Component_Function_3/N1  ( .A1(\SB2_0_27/i1[9] ), .A2(
        \SB2_0_27/i0_3 ), .A3(\SB2_0_27/i0[6] ), .ZN(
        \SB2_0_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_2/N2  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i0[10] ), .A3(\SB2_0_28/i0[6] ), .ZN(
        \SB2_0_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_28/Component_Function_4/N2  ( .A1(\SB2_0_28/i3[0] ), .A2(
        \SB2_0_28/i0_0 ), .A3(\SB2_0_28/i1_7 ), .ZN(
        \SB2_0_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_28/Component_Function_4/N1  ( .A1(\SB2_0_28/i0[9] ), .A2(
        \SB2_0_28/i0_0 ), .A3(\SB2_0_28/i0[8] ), .ZN(
        \SB2_0_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_2/N4  ( .A1(\SB2_0_29/i1_5 ), .A2(
        \SB2_0_29/i0_0 ), .A3(\SB2_0_29/i0_4 ), .ZN(
        \SB2_0_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_29/Component_Function_4/N2  ( .A1(\SB2_0_29/i3[0] ), .A2(
        \SB2_0_29/i0_0 ), .A3(\SB2_0_29/i1_7 ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_29/Component_Function_4/N1  ( .A1(\SB2_0_29/i0[9] ), .A2(
        \SB2_0_29/i0_0 ), .A3(\SB2_0_29/i0[8] ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_2/N2  ( .A1(\SB1_0_30/buf_output[5] ), 
        .A2(\SB2_0_30/i0[10] ), .A3(\SB2_0_30/i0[6] ), .ZN(
        \SB2_0_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_30/Component_Function_2/N1  ( .A1(\SB2_0_30/i1_5 ), .A2(
        \SB2_0_30/i0[10] ), .A3(\SB2_0_30/i1[9] ), .ZN(
        \SB2_0_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_3/N1  ( .A1(\SB2_0_30/i1[9] ), .A2(
        \SB2_0_30/i0_3 ), .A3(\SB2_0_30/i0[6] ), .ZN(
        \SB2_0_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_4/N4  ( .A1(\SB2_0_30/i1[9] ), .A2(
        \SB2_0_30/i1_5 ), .A3(\SB2_0_30/i0_4 ), .ZN(
        \SB2_0_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_30/Component_Function_4/N1  ( .A1(\SB2_0_30/i0[9] ), .A2(
        \SB2_0_30/i0_0 ), .A3(\SB2_0_30/i0[8] ), .ZN(
        \SB2_0_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_2/N2  ( .A1(\SB1_1_0/i0_3 ), .A2(
        \SB1_1_0/i0[10] ), .A3(\SB1_1_0/i0[6] ), .ZN(
        \SB1_1_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_1/Component_Function_2/N3  ( .A1(\SB1_1_1/i0_3 ), .A2(
        \SB1_1_1/i0[8] ), .A3(\SB1_1_1/i0[9] ), .ZN(
        \SB1_1_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_1/Component_Function_3/N2  ( .A1(\SB1_1_1/i0_0 ), .A2(
        \SB1_1_1/i0_3 ), .A3(\SB1_1_1/i0_4 ), .ZN(
        \SB1_1_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_1/Component_Function_4/N1  ( .A1(\SB1_1_1/i0[9] ), .A2(
        \SB1_1_1/i0_0 ), .A3(\SB1_1_1/i0[8] ), .ZN(
        \SB1_1_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_4/Component_Function_4/N2  ( .A1(\SB1_1_4/i3[0] ), .A2(
        \SB1_1_4/i0_0 ), .A3(\SB1_1_4/i1_7 ), .ZN(
        \SB1_1_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_5/Component_Function_4/N1  ( .A1(\SB1_1_5/i0[9] ), .A2(
        \SB1_1_5/i0_0 ), .A3(\SB1_1_5/i0[8] ), .ZN(
        \SB1_1_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_2/N2  ( .A1(\SB1_1_6/i0_3 ), .A2(
        \SB1_1_6/i0[10] ), .A3(\SB1_1_6/i0[6] ), .ZN(
        \SB1_1_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_6/Component_Function_3/N1  ( .A1(\SB1_1_6/i1[9] ), .A2(
        \SB1_1_6/i0_3 ), .A3(\SB1_1_6/i0[6] ), .ZN(
        \SB1_1_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_2/N1  ( .A1(\SB1_1_7/i1_5 ), .A2(
        \SB1_1_7/i0[10] ), .A3(\SB1_1_7/i1[9] ), .ZN(
        \SB1_1_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_4/N2  ( .A1(\SB1_1_7/i3[0] ), .A2(
        \SB1_1_7/i0_0 ), .A3(\SB1_1_7/i1_7 ), .ZN(
        \SB1_1_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_8/Component_Function_2/N2  ( .A1(\SB1_1_8/i0_3 ), .A2(
        \SB1_1_8/i0[10] ), .A3(\SB1_1_8/i0[6] ), .ZN(
        \SB1_1_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_8/Component_Function_4/N2  ( .A1(\SB1_1_8/i3[0] ), .A2(
        \SB1_1_8/i0_0 ), .A3(\SB1_1_8/i1_7 ), .ZN(
        \SB1_1_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_8/Component_Function_4/N1  ( .A1(\SB1_1_8/i0[9] ), .A2(
        \SB1_1_8/i0_0 ), .A3(\SB1_1_8/i0[8] ), .ZN(
        \SB1_1_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_2/N3  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i0[8] ), .A3(\SB1_1_9/i0[9] ), .ZN(
        \SB1_1_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_9/Component_Function_2/N2  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i0[10] ), .A3(\SB1_1_9/i0[6] ), .ZN(
        \SB1_1_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_9/Component_Function_3/N2  ( .A1(\SB1_1_9/i0_0 ), .A2(
        \SB1_1_9/i0_3 ), .A3(\SB1_1_9/i0_4 ), .ZN(
        \SB1_1_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_10/Component_Function_2/N2  ( .A1(\SB1_1_10/i0_3 ), .A2(
        \SB1_1_10/i0[10] ), .A3(\SB1_1_10/i0[6] ), .ZN(
        \SB1_1_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_10/Component_Function_2/N1  ( .A1(\SB1_1_10/i1_5 ), .A2(
        \SB1_1_10/i0[10] ), .A3(\SB1_1_10/i1[9] ), .ZN(
        \SB1_1_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_4/N2  ( .A1(\SB1_1_10/i3[0] ), .A2(
        \SB1_1_10/i0_0 ), .A3(\SB1_1_10/i1_7 ), .ZN(
        \SB1_1_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_10/Component_Function_4/N1  ( .A1(\SB1_1_10/i0[9] ), .A2(
        \SB1_1_10/i0_0 ), .A3(\SB1_1_10/i0[8] ), .ZN(
        \SB1_1_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_3/N1  ( .A1(\SB1_1_11/i1[9] ), .A2(
        \SB1_1_11/i0_3 ), .A3(\SB1_1_11/i0[6] ), .ZN(
        \SB1_1_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_4/N4  ( .A1(\SB1_1_11/i1[9] ), .A2(
        \SB1_1_11/i1_5 ), .A3(\SB1_1_11/i0_4 ), .ZN(
        \SB1_1_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_11/Component_Function_4/N2  ( .A1(\SB1_1_11/i3[0] ), .A2(
        \SB1_1_11/i0_0 ), .A3(\SB1_1_11/i1_7 ), .ZN(
        \SB1_1_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_11/Component_Function_4/N1  ( .A1(\SB1_1_11/i0[9] ), .A2(
        \SB1_1_11/i0_0 ), .A3(\SB1_1_11/i0[8] ), .ZN(
        \SB1_1_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_12/Component_Function_2/N3  ( .A1(\SB1_1_12/i0_3 ), .A2(
        \SB1_1_12/i0[8] ), .A3(\SB1_1_12/i0[9] ), .ZN(
        \SB1_1_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_12/Component_Function_4/N2  ( .A1(\SB1_1_12/i3[0] ), .A2(
        \SB1_1_12/i0_0 ), .A3(\SB1_1_12/i1_7 ), .ZN(
        \SB1_1_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_12/Component_Function_4/N1  ( .A1(\SB1_1_12/i0[9] ), .A2(
        \SB1_1_12/i0_0 ), .A3(\SB1_1_12/i0[8] ), .ZN(
        \SB1_1_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_2/N1  ( .A1(\SB1_1_13/i1_5 ), .A2(
        \SB1_1_13/i0[10] ), .A3(\SB1_1_13/i1[9] ), .ZN(
        \SB1_1_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_3/N1  ( .A1(\SB1_1_13/i1[9] ), .A2(
        \SB1_1_13/i0_3 ), .A3(\SB1_1_13/i0[6] ), .ZN(
        \SB1_1_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_14/Component_Function_4/N2  ( .A1(\SB1_1_14/i3[0] ), .A2(
        \SB1_1_14/i0_0 ), .A3(\SB1_1_14/i1_7 ), .ZN(
        \SB1_1_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_15/Component_Function_4/N4  ( .A1(\SB1_1_15/i1[9] ), .A2(
        \SB1_1_15/i1_5 ), .A3(\SB1_1_15/i0_4 ), .ZN(
        \SB1_1_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_15/Component_Function_4/N2  ( .A1(\SB1_1_15/i3[0] ), .A2(
        \SB1_1_15/i0_0 ), .A3(\SB1_1_15/i1_7 ), .ZN(
        \SB1_1_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_16/Component_Function_2/N1  ( .A1(\SB1_1_16/i1_5 ), .A2(
        \SB1_1_16/i0[10] ), .A3(\SB1_1_16/i1[9] ), .ZN(
        \SB1_1_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_16/Component_Function_4/N2  ( .A1(\SB1_1_16/i3[0] ), .A2(
        \SB1_1_16/i0_0 ), .A3(\SB1_1_16/i1_7 ), .ZN(
        \SB1_1_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_16/Component_Function_4/N1  ( .A1(\SB1_1_16/i0[9] ), .A2(
        \SB1_1_16/i0_0 ), .A3(\SB1_1_16/i0[8] ), .ZN(
        \SB1_1_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_2/N2  ( .A1(\SB1_1_17/i0_3 ), .A2(
        \SB1_1_17/i0[10] ), .A3(\SB1_1_17/i0[6] ), .ZN(
        \SB1_1_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_19/Component_Function_2/N1  ( .A1(\SB1_1_19/i1_5 ), .A2(
        \SB1_1_19/i0[10] ), .A3(\SB1_1_19/i1[9] ), .ZN(
        \SB1_1_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_4/N2  ( .A1(\SB1_1_19/i3[0] ), .A2(
        \SB1_1_19/i0_0 ), .A3(\SB1_1_19/i1_7 ), .ZN(
        \SB1_1_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_19/Component_Function_4/N1  ( .A1(\SB1_1_19/i0[9] ), .A2(
        \SB1_1_19/i0_0 ), .A3(\SB1_1_19/i0[8] ), .ZN(
        \SB1_1_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_3/N2  ( .A1(\SB1_1_20/i0_0 ), .A2(
        \SB1_1_20/i0_3 ), .A3(\SB1_1_20/i0_4 ), .ZN(
        \SB1_1_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_20/Component_Function_4/N1  ( .A1(\SB1_1_20/i0[9] ), .A2(
        \SB1_1_20/i0_0 ), .A3(\SB1_1_20/i0[8] ), .ZN(
        \SB1_1_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_4/N1  ( .A1(\SB1_1_21/i0[9] ), .A2(
        \SB1_1_21/i0_0 ), .A3(\SB1_1_21/i0[8] ), .ZN(
        \SB1_1_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_22/Component_Function_4/N2  ( .A1(\SB1_1_22/i3[0] ), .A2(
        \SB1_1_22/i0_0 ), .A3(\SB1_1_22/i1_7 ), .ZN(
        \SB1_1_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_22/Component_Function_4/N1  ( .A1(\SB1_1_22/i0[9] ), .A2(
        \SB1_1_22/i0_0 ), .A3(\SB1_1_22/i0[8] ), .ZN(
        \SB1_1_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_24/Component_Function_4/N2  ( .A1(\SB1_1_24/i3[0] ), .A2(
        \SB1_1_24/i0_0 ), .A3(\SB1_1_24/i1_7 ), .ZN(
        \SB1_1_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_24/Component_Function_4/N1  ( .A1(\SB1_1_24/i0[9] ), .A2(
        \SB1_1_24/i0_0 ), .A3(\SB1_1_24/i0[8] ), .ZN(
        \SB1_1_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_3/N2  ( .A1(\SB1_1_25/i0_0 ), .A2(
        \SB1_1_25/i0_3 ), .A3(\SB1_1_25/i0_4 ), .ZN(
        \SB1_1_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N4  ( .A1(\SB1_1_25/i1[9] ), .A2(
        \SB1_1_25/i1_5 ), .A3(\SB1_1_25/i0_4 ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N2  ( .A1(\SB1_1_25/i3[0] ), .A2(
        \SB1_1_25/i0_0 ), .A3(\SB1_1_25/i1_7 ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N1  ( .A1(\SB1_1_25/i0[9] ), .A2(
        \SB1_1_25/i0_0 ), .A3(\SB1_1_25/i0[8] ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_3/N1  ( .A1(\SB1_1_26/i1[9] ), .A2(
        \SB1_1_26/i0_3 ), .A3(\SB1_1_26/i0[6] ), .ZN(
        \SB1_1_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_4/N2  ( .A1(\SB1_1_26/i3[0] ), .A2(
        \SB1_1_26/i0_0 ), .A3(\SB1_1_26/i1_7 ), .ZN(
        \SB1_1_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_26/Component_Function_4/N1  ( .A1(\SB1_1_26/i0[9] ), .A2(
        \SB1_1_26/i0_0 ), .A3(\SB1_1_26/i0[8] ), .ZN(
        \SB1_1_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_4/N2  ( .A1(\SB1_1_28/i3[0] ), .A2(
        \SB1_1_28/i0_0 ), .A3(\SB1_1_28/i1_7 ), .ZN(
        \SB1_1_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_28/Component_Function_4/N1  ( .A1(\SB1_1_28/i0[9] ), .A2(
        \SB1_1_28/i0_0 ), .A3(\SB1_1_28/i0[8] ), .ZN(
        \SB1_1_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_2/N2  ( .A1(\SB1_1_29/i0_3 ), .A2(
        \SB1_1_29/i0[10] ), .A3(\SB1_1_29/i0[6] ), .ZN(
        \SB1_1_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_29/Component_Function_2/N1  ( .A1(\SB1_1_29/i1_5 ), .A2(
        \SB1_1_29/i0[10] ), .A3(\SB1_1_29/i1[9] ), .ZN(
        \SB1_1_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_3/N1  ( .A1(\SB1_1_29/i1[9] ), .A2(
        \SB1_1_29/i0_3 ), .A3(\SB1_1_29/i0[6] ), .ZN(
        \SB1_1_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_4/N3  ( .A1(\SB1_1_31/i0[9] ), .A2(
        \SB1_1_31/i0[10] ), .A3(\SB1_1_31/i0_3 ), .ZN(
        \SB1_1_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_31/Component_Function_4/N2  ( .A1(\SB1_1_31/i3[0] ), .A2(
        \SB1_1_31/i0_0 ), .A3(\SB1_1_31/i1_7 ), .ZN(
        \SB1_1_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_31/Component_Function_4/N1  ( .A1(\SB1_1_31/i0[9] ), .A2(
        \SB1_1_31/i0_0 ), .A3(\SB1_1_31/i0[8] ), .ZN(
        \SB1_1_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_0/Component_Function_4/N2  ( .A1(\SB2_1_0/i3[0] ), .A2(
        \SB2_1_0/i0_0 ), .A3(\SB2_1_0/i1_7 ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_1/Component_Function_4/N3  ( .A1(\SB2_1_1/i0[9] ), .A2(
        \SB2_1_1/i0[10] ), .A3(\SB2_1_1/i0_3 ), .ZN(
        \SB2_1_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_1/Component_Function_4/N2  ( .A1(\SB2_1_1/i3[0] ), .A2(
        \SB2_1_1/i0_0 ), .A3(\SB2_1_1/i1_7 ), .ZN(
        \SB2_1_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_1/Component_Function_4/N1  ( .A1(\SB2_1_1/i0[9] ), .A2(
        \SB2_1_1/i0_0 ), .A3(\SB2_1_1/i0[8] ), .ZN(
        \SB2_1_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_4/N4  ( .A1(\SB2_1_2/i1[9] ), .A2(
        \SB2_1_2/i1_5 ), .A3(\SB2_1_2/i0_4 ), .ZN(
        \SB2_1_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_2/Component_Function_4/N2  ( .A1(\SB2_1_2/i3[0] ), .A2(
        \SB2_1_2/i0_0 ), .A3(\SB2_1_2/i1_7 ), .ZN(
        \SB2_1_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_2/Component_Function_4/N1  ( .A1(\SB2_1_2/i0[9] ), .A2(
        \SB2_1_2/i0_0 ), .A3(\SB2_1_2/i0[8] ), .ZN(
        \SB2_1_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_3/Component_Function_4/N2  ( .A1(\SB2_1_3/i3[0] ), .A2(
        \SB2_1_3/i0_0 ), .A3(\SB2_1_3/i1_7 ), .ZN(
        \SB2_1_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_3/Component_Function_4/N1  ( .A1(\SB1_1_8/buf_output[0] ), 
        .A2(\SB2_1_3/i0_0 ), .A3(\SB2_1_3/i0[8] ), .ZN(
        \SB2_1_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_4/Component_Function_4/N2  ( .A1(\SB2_1_4/i3[0] ), .A2(
        \SB2_1_4/i0_0 ), .A3(n2656), .ZN(
        \SB2_1_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_5/Component_Function_4/N2  ( .A1(\SB2_1_5/i3[0] ), .A2(
        \SB2_1_5/i0_0 ), .A3(\SB2_1_5/i1_7 ), .ZN(
        \SB2_1_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_5/Component_Function_4/N1  ( .A1(\SB2_1_5/i0[9] ), .A2(
        \SB2_1_5/i0_0 ), .A3(\SB2_1_5/i0[8] ), .ZN(
        \SB2_1_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_2/N1  ( .A1(\SB2_1_6/i1_5 ), .A2(
        \SB2_1_6/i0[10] ), .A3(\SB2_1_6/i1[9] ), .ZN(
        \SB2_1_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_4/N4  ( .A1(\SB2_1_6/i1[9] ), .A2(
        \SB2_1_6/i1_5 ), .A3(\SB2_1_6/i0_4 ), .ZN(
        \SB2_1_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_6/Component_Function_4/N2  ( .A1(\SB2_1_6/i3[0] ), .A2(
        \SB2_1_6/i0_0 ), .A3(\SB2_1_6/i1_7 ), .ZN(
        \SB2_1_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_8/Component_Function_2/N4  ( .A1(\SB2_1_8/i1_5 ), .A2(
        \SB1_1_11/buf_output[2] ), .A3(\SB1_1_9/buf_output[4] ), .ZN(
        \SB2_1_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_9/Component_Function_4/N2  ( .A1(\SB2_1_9/i3[0] ), .A2(
        \SB2_1_9/i0_0 ), .A3(\SB2_1_9/i1_7 ), .ZN(
        \SB2_1_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_9/Component_Function_4/N1  ( .A1(\SB2_1_9/i0[9] ), .A2(
        \SB2_1_9/i0_0 ), .A3(\SB2_1_9/i0[8] ), .ZN(
        \SB2_1_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_10/Component_Function_4/N2  ( .A1(\SB2_1_10/i3[0] ), .A2(
        \SB2_1_10/i0_0 ), .A3(\SB2_1_10/i1_7 ), .ZN(
        \SB2_1_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_11/Component_Function_4/N2  ( .A1(\SB2_1_11/i3[0] ), .A2(
        \SB2_1_11/i0_0 ), .A3(\SB2_1_11/i1_7 ), .ZN(
        \SB2_1_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_11/Component_Function_4/N1  ( .A1(\SB2_1_11/i0[9] ), .A2(
        \SB2_1_11/i0_0 ), .A3(\SB2_1_11/i0[8] ), .ZN(
        \SB2_1_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_12/Component_Function_4/N1  ( .A1(\SB2_1_12/i0[9] ), .A2(
        \SB2_1_12/i0_0 ), .A3(\SB2_1_12/i0[8] ), .ZN(
        \SB2_1_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_14/Component_Function_4/N4  ( .A1(\SB2_1_14/i1[9] ), .A2(
        \SB2_1_14/i1_5 ), .A3(\SB2_1_14/i0_4 ), .ZN(
        \SB2_1_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_14/Component_Function_4/N1  ( .A1(\SB2_1_14/i0[9] ), .A2(
        \SB2_1_14/i0_0 ), .A3(\SB2_1_14/i0[8] ), .ZN(
        \SB2_1_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_15/Component_Function_3/N2  ( .A1(\SB2_1_15/i0_0 ), .A2(
        \SB2_1_15/i0_3 ), .A3(\SB2_1_15/i0_4 ), .ZN(
        \SB2_1_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_15/Component_Function_4/N2  ( .A1(\SB2_1_15/i3[0] ), .A2(
        \SB2_1_15/i0_0 ), .A3(\SB2_1_15/i1_7 ), .ZN(
        \SB2_1_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_16/Component_Function_4/N2  ( .A1(\SB2_1_16/i3[0] ), .A2(
        \SB2_1_16/i0_0 ), .A3(\SB2_1_16/i1_7 ), .ZN(
        \SB2_1_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_16/Component_Function_4/N1  ( .A1(\SB2_1_16/i0[9] ), .A2(
        \SB2_1_16/i0_0 ), .A3(\SB2_1_16/i0[8] ), .ZN(
        \SB2_1_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_3/N2  ( .A1(\SB2_1_17/i0_0 ), .A2(
        \SB1_1_17/buf_output[5] ), .A3(\SB2_1_17/i0_4 ), .ZN(
        \SB2_1_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_17/Component_Function_4/N2  ( .A1(\SB2_1_17/i3[0] ), .A2(
        \SB2_1_17/i0_0 ), .A3(\SB2_1_17/i1_7 ), .ZN(
        \SB2_1_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_17/Component_Function_4/N1  ( .A1(\SB2_1_17/i0[9] ), .A2(
        \SB2_1_17/i0_0 ), .A3(\SB2_1_17/i0[8] ), .ZN(
        \SB2_1_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_4/N1  ( .A1(\SB2_1_18/i0[9] ), .A2(
        \SB2_1_18/i0_0 ), .A3(\SB2_1_18/i0[8] ), .ZN(
        \SB2_1_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_19/Component_Function_4/N1  ( .A1(\SB2_1_19/i0[9] ), .A2(
        \SB2_1_19/i0_0 ), .A3(\SB2_1_19/i0[8] ), .ZN(
        \SB2_1_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_4/N2  ( .A1(\SB2_1_22/i3[0] ), .A2(
        \SB2_1_22/i0_0 ), .A3(\SB2_1_22/i1_7 ), .ZN(
        \SB2_1_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_22/Component_Function_4/N1  ( .A1(\SB2_1_22/i0[9] ), .A2(
        \SB2_1_22/i0_0 ), .A3(n6283), .ZN(
        \SB2_1_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N2  ( .A1(\SB2_1_23/i3[0] ), .A2(
        \SB2_1_23/i0_0 ), .A3(\SB2_1_23/i1_7 ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N1  ( .A1(\SB2_1_23/i0[9] ), .A2(
        \SB2_1_23/i0_0 ), .A3(\SB2_1_23/i0[8] ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_24/Component_Function_3/N4  ( .A1(\SB2_1_24/i1_5 ), .A2(
        \SB2_1_24/i0[8] ), .A3(\SB2_1_24/i3[0] ), .ZN(
        \SB2_1_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_24/Component_Function_4/N2  ( .A1(\SB2_1_24/i3[0] ), .A2(
        \SB2_1_24/i0_0 ), .A3(\SB2_1_24/i1_7 ), .ZN(
        \SB2_1_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_24/Component_Function_4/N1  ( .A1(\SB2_1_24/i0[9] ), .A2(
        \SB2_1_24/i0_0 ), .A3(\SB2_1_24/i0[8] ), .ZN(
        \SB2_1_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_25/Component_Function_4/N2  ( .A1(\SB2_1_25/i3[0] ), .A2(
        \SB2_1_25/i0_0 ), .A3(\SB2_1_25/i1_7 ), .ZN(
        \SB2_1_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_25/Component_Function_4/N1  ( .A1(\SB2_1_25/i0[9] ), .A2(
        \SB2_1_25/i0_0 ), .A3(n3995), .ZN(
        \SB2_1_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_2/N1  ( .A1(\SB2_1_26/i1_5 ), .A2(
        \SB2_1_26/i0[10] ), .A3(\SB2_1_26/i1[9] ), .ZN(
        \SB2_1_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N4  ( .A1(\SB2_1_26/i1[9] ), .A2(
        \SB2_1_26/i1_5 ), .A3(\SB2_1_26/i0_4 ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N1  ( .A1(\SB2_1_26/i0[9] ), .A2(
        \SB2_1_26/i0_0 ), .A3(\SB2_1_26/i0[8] ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_4/N2  ( .A1(\SB2_1_27/i3[0] ), .A2(
        \RI3[1][26] ), .A3(\SB2_1_27/i1_7 ), .ZN(
        \SB2_1_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_27/Component_Function_4/N1  ( .A1(\SB2_1_27/i0[9] ), .A2(
        \RI3[1][26] ), .A3(\SB2_1_27/i0[8] ), .ZN(
        \SB2_1_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_28/Component_Function_4/N1  ( .A1(\SB2_1_28/i0[9] ), .A2(
        \SB2_1_28/i0_0 ), .A3(\SB2_1_28/i0[8] ), .ZN(
        \SB2_1_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_2/N3  ( .A1(\SB2_1_29/i0_3 ), .A2(
        \SB2_1_29/i0[8] ), .A3(\SB2_1_29/i0[9] ), .ZN(
        \SB2_1_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_29/Component_Function_3/N1  ( .A1(\SB2_1_29/i1[9] ), .A2(
        \SB2_1_29/i0_3 ), .A3(\SB2_1_29/i0[6] ), .ZN(
        \SB2_1_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_4/N2  ( .A1(\SB2_1_29/i3[0] ), .A2(
        \SB2_1_29/i0_0 ), .A3(\SB2_1_29/i1_7 ), .ZN(
        \SB2_1_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_29/Component_Function_4/N1  ( .A1(\SB2_1_29/i0[9] ), .A2(
        \SB2_1_29/i0_0 ), .A3(\SB2_1_29/i0[8] ), .ZN(
        \SB2_1_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_4/N2  ( .A1(\SB2_1_30/i3[0] ), .A2(
        \SB2_1_30/i0_0 ), .A3(\SB2_1_30/i1_7 ), .ZN(
        \SB2_1_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_30/Component_Function_4/N1  ( .A1(\SB2_1_30/i0[9] ), .A2(
        \SB2_1_30/i0_0 ), .A3(\SB2_1_30/i0[8] ), .ZN(
        \SB2_1_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_31/Component_Function_4/N1  ( .A1(\SB2_1_31/i0[9] ), .A2(
        \SB2_1_31/i0_0 ), .A3(\SB2_1_31/i0[8] ), .ZN(
        \SB2_1_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_4/N1  ( .A1(\SB1_2_0/i0[9] ), .A2(
        \SB1_2_0/i0_0 ), .A3(\SB1_2_0/i0[8] ), .ZN(
        \SB1_2_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_2/N3  ( .A1(\SB1_2_1/i0_3 ), .A2(
        \SB1_2_1/i0[8] ), .A3(\SB1_2_1/i0[9] ), .ZN(
        \SB1_2_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_2/Component_Function_3/N2  ( .A1(\SB1_2_2/i0_0 ), .A2(
        \SB1_2_2/i0_3 ), .A3(\SB1_2_2/i0_4 ), .ZN(
        \SB1_2_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_3/Component_Function_2/N1  ( .A1(\SB1_2_3/i1_5 ), .A2(
        \SB1_2_3/i0[10] ), .A3(\SB1_2_3/i1[9] ), .ZN(
        \SB1_2_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_3/N2  ( .A1(\SB1_2_4/i0_0 ), .A2(
        \SB1_2_4/i0_3 ), .A3(\SB1_2_4/i0_4 ), .ZN(
        \SB1_2_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_6/Component_Function_3/N1  ( .A1(\SB1_2_6/i1[9] ), .A2(
        \SB1_2_6/i0_3 ), .A3(\SB1_2_6/i0[6] ), .ZN(
        \SB1_2_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_4/N2  ( .A1(\SB1_2_6/i3[0] ), .A2(
        \SB1_2_6/i0_0 ), .A3(\SB1_2_6/i1_7 ), .ZN(
        \SB1_2_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_6/Component_Function_4/N1  ( .A1(\SB1_2_6/i0[9] ), .A2(
        \SB1_2_6/i0_0 ), .A3(\SB1_2_6/i0[8] ), .ZN(
        \SB1_2_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_4/N2  ( .A1(\SB1_2_7/i3[0] ), .A2(
        \SB1_2_7/i0_0 ), .A3(\SB1_2_7/i1_7 ), .ZN(
        \SB1_2_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_7/Component_Function_4/N1  ( .A1(\SB1_2_7/i0[9] ), .A2(
        \SB1_2_7/i0_0 ), .A3(n3184), .ZN(
        \SB1_2_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_2/N4  ( .A1(\SB1_2_8/i1_5 ), .A2(
        \SB1_2_8/i0_0 ), .A3(\SB1_2_8/i0_4 ), .ZN(
        \SB1_2_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_8/Component_Function_3/N2  ( .A1(\SB1_2_8/i0_0 ), .A2(
        \SB1_2_8/i0_3 ), .A3(\SB1_2_8/i0_4 ), .ZN(
        \SB1_2_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_8/Component_Function_4/N2  ( .A1(\SB1_2_8/i3[0] ), .A2(
        \SB1_2_8/i0_0 ), .A3(\SB1_2_8/i1_7 ), .ZN(
        \SB1_2_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_8/Component_Function_4/N1  ( .A1(\SB1_2_8/i0[9] ), .A2(
        \SB1_2_8/i0_0 ), .A3(\SB1_2_8/i0[8] ), .ZN(
        \SB1_2_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_4/N2  ( .A1(\SB1_2_9/i3[0] ), .A2(
        \SB1_2_9/i0_0 ), .A3(\SB1_2_9/i1_7 ), .ZN(
        \SB1_2_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_9/Component_Function_4/N1  ( .A1(\SB1_2_9/i0[9] ), .A2(
        \SB1_2_9/i0_0 ), .A3(\SB1_2_9/i0[8] ), .ZN(
        \SB1_2_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_2/N2  ( .A1(\SB1_2_10/i0_3 ), .A2(
        \SB1_2_10/i0[10] ), .A3(\SB1_2_10/i0[6] ), .ZN(
        \SB1_2_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_10/Component_Function_3/N2  ( .A1(\SB1_2_10/i0_0 ), .A2(
        \SB1_2_10/i0_3 ), .A3(\SB1_2_10/i0_4 ), .ZN(
        \SB1_2_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_10/Component_Function_4/N1  ( .A1(\SB1_2_10/i0[9] ), .A2(
        \SB1_2_10/i0_0 ), .A3(\SB1_2_10/i0[8] ), .ZN(
        \SB1_2_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_2/N1  ( .A1(\SB1_2_11/i1_5 ), .A2(
        \SB1_2_11/i0[10] ), .A3(\SB1_2_11/i1[9] ), .ZN(
        \SB1_2_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_3/N2  ( .A1(\SB1_2_11/i0_0 ), .A2(
        \SB1_2_11/i0_3 ), .A3(\SB1_2_11/i0_4 ), .ZN(
        \SB1_2_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_11/Component_Function_4/N2  ( .A1(\SB1_2_11/i3[0] ), .A2(
        \SB1_2_11/i0_0 ), .A3(\SB1_2_11/i1_7 ), .ZN(
        \SB1_2_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_13/Component_Function_4/N2  ( .A1(\SB1_2_13/i3[0] ), .A2(
        \SB1_2_13/i0_0 ), .A3(\SB1_2_13/i1_7 ), .ZN(
        \SB1_2_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_13/Component_Function_4/N1  ( .A1(\SB1_2_13/i0[9] ), .A2(
        \SB1_2_13/i0_0 ), .A3(\SB1_2_13/i0[8] ), .ZN(
        \SB1_2_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_3/N2  ( .A1(\SB1_2_14/i0_0 ), .A2(
        \RI1[2][107] ), .A3(\SB1_2_14/i0_4 ), .ZN(
        \SB1_2_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_14/Component_Function_4/N2  ( .A1(\SB1_2_14/i3[0] ), .A2(
        \SB1_2_14/i0_0 ), .A3(\SB1_2_14/i1_7 ), .ZN(
        \SB1_2_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_14/Component_Function_4/N1  ( .A1(\SB1_2_14/i0[9] ), .A2(
        \SB1_2_14/i0_0 ), .A3(\SB1_2_14/i0[8] ), .ZN(
        \SB1_2_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_16/Component_Function_4/N2  ( .A1(\SB1_2_16/i3[0] ), .A2(
        \SB1_2_16/i0_0 ), .A3(\SB1_2_16/i1_7 ), .ZN(
        \SB1_2_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_16/Component_Function_4/N1  ( .A1(\SB1_2_16/i0[9] ), .A2(
        \SB1_2_16/i0_0 ), .A3(\SB1_2_16/i0[8] ), .ZN(
        \SB1_2_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_17/Component_Function_4/N1  ( .A1(\SB1_2_17/i0[9] ), .A2(
        \SB1_2_17/i0_0 ), .A3(\SB1_2_17/i0[8] ), .ZN(
        \SB1_2_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_4/N4  ( .A1(\SB1_2_18/i1[9] ), .A2(
        \SB1_2_18/i1_5 ), .A3(\SB1_2_18/i0_4 ), .ZN(
        \SB1_2_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_18/Component_Function_4/N2  ( .A1(\SB1_2_18/i3[0] ), .A2(
        \SB1_2_18/i0_0 ), .A3(\SB1_2_18/i1_7 ), .ZN(
        \SB1_2_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_19/Component_Function_2/N3  ( .A1(\SB1_2_19/i0_3 ), .A2(
        \SB1_2_19/i0[8] ), .A3(\SB1_2_19/i0[9] ), .ZN(
        \SB1_2_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_20/Component_Function_2/N1  ( .A1(\SB1_2_20/i1_5 ), .A2(
        \SB1_2_20/i0[10] ), .A3(\SB1_2_20/i1[9] ), .ZN(
        \SB1_2_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_3/N2  ( .A1(\SB1_2_20/i0_0 ), .A2(
        \SB1_2_20/i0_3 ), .A3(\SB1_2_20/i0_4 ), .ZN(
        \SB1_2_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_20/Component_Function_4/N1  ( .A1(\SB1_2_20/i0[9] ), .A2(
        \SB1_2_20/i0_0 ), .A3(\SB1_2_20/i0[8] ), .ZN(
        \SB1_2_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_2/N2  ( .A1(\SB1_2_21/i0_3 ), .A2(
        \SB1_2_21/i0[10] ), .A3(\SB1_2_21/i0[6] ), .ZN(
        \SB1_2_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_21/Component_Function_3/N3  ( .A1(\SB1_2_21/i1[9] ), .A2(
        \SB1_2_21/i1_7 ), .A3(\SB1_2_21/i0[10] ), .ZN(
        \SB1_2_21/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_21/Component_Function_3/N1  ( .A1(\SB1_2_21/i1[9] ), .A2(
        \SB1_2_21/i0_3 ), .A3(\SB1_2_21/i0[6] ), .ZN(
        \SB1_2_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_4/N2  ( .A1(\SB1_2_21/i3[0] ), .A2(
        \SB1_2_21/i0_0 ), .A3(\SB1_2_21/i1_7 ), .ZN(
        \SB1_2_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_22/Component_Function_4/N2  ( .A1(\SB1_2_22/i3[0] ), .A2(
        \SB1_2_22/i0_0 ), .A3(\SB1_2_22/i1_7 ), .ZN(
        \SB1_2_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_2/N2  ( .A1(\SB1_2_23/i0_3 ), .A2(
        \SB1_2_23/i0[10] ), .A3(\SB1_2_23/i0[6] ), .ZN(
        \SB1_2_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_3/N3  ( .A1(\SB1_2_23/i1[9] ), .A2(
        \SB1_2_23/i1_7 ), .A3(\SB1_2_23/i0[10] ), .ZN(
        \SB1_2_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_23/Component_Function_4/N4  ( .A1(\SB1_2_23/i1[9] ), .A2(
        \SB1_2_23/i1_5 ), .A3(\SB1_2_23/i0_4 ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_23/Component_Function_4/N2  ( .A1(\SB1_2_23/i3[0] ), .A2(
        \SB1_2_23/i0_0 ), .A3(\SB1_2_23/i1_7 ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_4/N1  ( .A1(\SB1_2_23/i0[9] ), .A2(
        \SB1_2_23/i0_0 ), .A3(\SB1_2_23/i0[8] ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_4/N4  ( .A1(\SB1_2_24/i1[9] ), .A2(
        \SB1_2_24/i1_5 ), .A3(\MC_ARK_ARC_1_1/buf_output[46] ), .ZN(
        \SB1_2_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_2/N3  ( .A1(\SB1_2_25/i0_3 ), .A2(
        \SB1_2_25/i0[8] ), .A3(\SB1_2_25/i0[9] ), .ZN(
        \SB1_2_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_25/Component_Function_4/N2  ( .A1(\SB1_2_25/i3[0] ), .A2(
        \SB1_2_25/i0_0 ), .A3(\SB1_2_25/i1_7 ), .ZN(
        \SB1_2_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_25/Component_Function_4/N1  ( .A1(\SB1_2_25/i0[9] ), .A2(
        \SB1_2_25/i0_0 ), .A3(\SB1_2_25/i0[8] ), .ZN(
        \SB1_2_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_2/N2  ( .A1(\SB1_2_27/i0_3 ), .A2(
        \SB1_2_27/i0[10] ), .A3(\SB1_2_27/i0[6] ), .ZN(
        \SB1_2_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_28/Component_Function_3/N2  ( .A1(\SB1_2_28/i0_0 ), .A2(
        \SB1_2_28/i0_3 ), .A3(\SB1_2_28/i0_4 ), .ZN(
        \SB1_2_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_29/Component_Function_4/N1  ( .A1(\SB1_2_29/i0[9] ), .A2(
        \SB1_2_29/i0_0 ), .A3(\SB1_2_29/i0[8] ), .ZN(
        \SB1_2_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_4/N2  ( .A1(\SB1_2_30/i3[0] ), .A2(
        \SB1_2_30/i0_0 ), .A3(\SB1_2_30/i1_7 ), .ZN(
        \SB1_2_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_30/Component_Function_4/N1  ( .A1(\SB1_2_30/i0[9] ), .A2(
        \SB1_2_30/i0_0 ), .A3(\SB1_2_30/i0[8] ), .ZN(
        \SB1_2_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_2/N2  ( .A1(\SB1_2_31/i0_3 ), .A2(
        \SB1_2_31/i0[10] ), .A3(\SB1_2_31/i0[6] ), .ZN(
        \SB1_2_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_31/Component_Function_2/N1  ( .A1(\SB1_2_31/i1_5 ), .A2(
        \SB1_2_31/i0[10] ), .A3(\SB1_2_31/i1[9] ), .ZN(
        \SB1_2_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_4/N2  ( .A1(\SB1_2_31/i3[0] ), .A2(
        \SB1_2_31/i0_0 ), .A3(\SB1_2_31/i1_7 ), .ZN(
        \SB1_2_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_0/Component_Function_2/N1  ( .A1(\SB2_2_0/i1_5 ), .A2(
        \SB2_2_0/i0[10] ), .A3(\SB2_2_0/i1[9] ), .ZN(
        \SB2_2_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_1/Component_Function_4/N2  ( .A1(\SB2_2_1/i3[0] ), .A2(
        \SB2_2_1/i0_0 ), .A3(\SB2_2_1/i1_7 ), .ZN(
        \SB2_2_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_2/Component_Function_4/N2  ( .A1(\SB2_2_2/i3[0] ), .A2(
        \SB2_2_2/i0_0 ), .A3(\SB2_2_2/i1_7 ), .ZN(
        \SB2_2_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_2/Component_Function_4/N1  ( .A1(\SB2_2_2/i0[9] ), .A2(
        \SB2_2_2/i0_0 ), .A3(\SB2_2_2/i0[8] ), .ZN(
        \SB2_2_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_3/Component_Function_4/N2  ( .A1(\SB2_2_3/i3[0] ), .A2(
        \SB2_2_3/i0_0 ), .A3(\SB2_2_3/i1_7 ), .ZN(
        \SB2_2_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_3/Component_Function_4/N1  ( .A1(\SB2_2_3/i0[9] ), .A2(
        \SB2_2_3/i0_0 ), .A3(n3991), .ZN(
        \SB2_2_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_5/Component_Function_4/N4  ( .A1(\SB2_2_5/i1[9] ), .A2(
        \SB2_2_5/i1_5 ), .A3(\SB2_2_5/i0_4 ), .ZN(
        \SB2_2_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_5/Component_Function_4/N1  ( .A1(\SB2_2_5/i0[9] ), .A2(
        \SB2_2_5/i0_0 ), .A3(\SB2_2_5/i0[8] ), .ZN(
        \SB2_2_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_3/N4  ( .A1(\SB2_2_6/i1_5 ), .A2(
        \SB2_2_6/i0[8] ), .A3(\SB2_2_6/i3[0] ), .ZN(
        \SB2_2_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_6/Component_Function_4/N2  ( .A1(\SB2_2_6/i3[0] ), .A2(
        \SB2_2_6/i0_0 ), .A3(\SB2_2_6/i1_7 ), .ZN(
        \SB2_2_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_8/Component_Function_4/N1  ( .A1(\SB2_2_8/i0[9] ), .A2(
        \SB2_2_8/i0_0 ), .A3(\SB2_2_8/i0[8] ), .ZN(
        \SB2_2_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_9/Component_Function_4/N1  ( .A1(\SB2_2_9/i0[9] ), .A2(
        \SB2_2_9/i0_0 ), .A3(\SB2_2_9/i0[8] ), .ZN(
        \SB2_2_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_11/Component_Function_4/N2  ( .A1(\SB2_2_11/i3[0] ), .A2(
        \SB2_2_11/i0_0 ), .A3(\SB2_2_11/i1_7 ), .ZN(
        \SB2_2_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_11/Component_Function_4/N1  ( .A1(\SB2_2_11/i0[9] ), .A2(
        \SB2_2_11/i0_0 ), .A3(\SB2_2_11/i0[8] ), .ZN(
        \SB2_2_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_14/Component_Function_4/N2  ( .A1(\SB2_2_14/i3[0] ), .A2(
        \SB2_2_14/i0_0 ), .A3(\SB2_2_14/i1_7 ), .ZN(
        \SB2_2_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_14/Component_Function_4/N1  ( .A1(\SB2_2_14/i0[9] ), .A2(
        \SB2_2_14/i0_0 ), .A3(\SB2_2_14/i0[8] ), .ZN(
        \SB2_2_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_15/Component_Function_4/N4  ( .A1(\SB2_2_15/i1[9] ), .A2(
        \SB2_2_15/i1_5 ), .A3(\SB2_2_15/i0_4 ), .ZN(
        \SB2_2_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_15/Component_Function_4/N2  ( .A1(\SB2_2_15/i3[0] ), .A2(
        \SB2_2_15/i0_0 ), .A3(\SB2_2_15/i1_7 ), .ZN(
        \SB2_2_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_16/Component_Function_4/N2  ( .A1(\SB2_2_16/i3[0] ), .A2(
        \SB2_2_16/i0_0 ), .A3(\SB2_2_16/i1_7 ), .ZN(
        \SB2_2_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_16/Component_Function_4/N1  ( .A1(\SB2_2_16/i0[9] ), .A2(
        \SB2_2_16/i0_0 ), .A3(\SB2_2_16/i0[8] ), .ZN(
        \SB2_2_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_17/Component_Function_4/N1  ( .A1(\SB2_2_17/i0[9] ), .A2(
        \SB2_2_17/i0_0 ), .A3(\SB2_2_17/i0[8] ), .ZN(
        \SB2_2_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_18/Component_Function_4/N2  ( .A1(\SB2_2_18/i3[0] ), .A2(
        \SB2_2_18/i0_0 ), .A3(\SB2_2_18/i1_7 ), .ZN(
        \SB2_2_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_18/Component_Function_4/N1  ( .A1(\SB2_2_18/i0[9] ), .A2(
        \SB2_2_18/i0_0 ), .A3(\SB2_2_18/i0[8] ), .ZN(
        \SB2_2_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_4/N1  ( .A1(\SB2_2_19/i0[9] ), .A2(
        \SB2_2_19/i0_0 ), .A3(\SB2_2_19/i0[8] ), .ZN(
        \SB2_2_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_20/Component_Function_4/N2  ( .A1(\SB2_2_20/i3[0] ), .A2(
        \SB2_2_20/i0_0 ), .A3(\SB2_2_20/i1_7 ), .ZN(
        \SB2_2_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_20/Component_Function_4/N1  ( .A1(\SB2_2_20/i0[9] ), .A2(
        \SB2_2_20/i0_0 ), .A3(\SB2_2_20/i0[8] ), .ZN(
        \SB2_2_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_21/Component_Function_4/N2  ( .A1(\SB2_2_21/i3[0] ), .A2(
        \SB2_2_21/i0_0 ), .A3(\SB2_2_21/i1_7 ), .ZN(
        \SB2_2_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_21/Component_Function_4/N1  ( .A1(\SB2_2_21/i0[9] ), .A2(
        \SB2_2_21/i0_0 ), .A3(\SB2_2_21/i0[8] ), .ZN(
        \SB2_2_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_22/Component_Function_4/N4  ( .A1(\SB2_2_22/i1[9] ), .A2(
        \SB2_2_22/i1_5 ), .A3(\SB2_2_22/i0_4 ), .ZN(
        \SB2_2_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_23/Component_Function_4/N2  ( .A1(\SB2_2_23/i3[0] ), .A2(
        \SB2_2_23/i0_0 ), .A3(\SB2_2_23/i1_7 ), .ZN(
        \SB2_2_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_23/Component_Function_4/N1  ( .A1(\SB2_2_23/i0[9] ), .A2(
        \SB2_2_23/i0_0 ), .A3(\SB2_2_23/i0[8] ), .ZN(
        \SB2_2_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_24/Component_Function_4/N2  ( .A1(\SB2_2_24/i3[0] ), .A2(
        \SB2_2_24/i0_0 ), .A3(\SB2_2_24/i1_7 ), .ZN(
        \SB2_2_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_24/Component_Function_4/N1  ( .A1(\SB2_2_24/i0[9] ), .A2(
        \SB2_2_24/i0_0 ), .A3(\SB2_2_24/i0[8] ), .ZN(
        \SB2_2_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_4/N1  ( .A1(\SB2_2_25/i0[9] ), .A2(
        \SB2_2_25/i0_0 ), .A3(\SB2_2_25/i0[8] ), .ZN(
        \SB2_2_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_4/N3  ( .A1(\SB2_2_26/i0[9] ), .A2(
        \SB2_2_26/i0[10] ), .A3(\SB2_2_26/i0_3 ), .ZN(
        \SB2_2_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_26/Component_Function_4/N1  ( .A1(\SB2_2_26/i0[9] ), .A2(
        \SB2_2_26/i0_0 ), .A3(\SB2_2_26/i0[8] ), .ZN(
        \SB2_2_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_27/Component_Function_4/N1  ( .A1(\SB2_2_27/i0[9] ), .A2(
        \SB2_2_27/i0_0 ), .A3(\SB2_2_27/i0[8] ), .ZN(
        \SB2_2_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_2/N1  ( .A1(\SB2_2_29/i1_5 ), .A2(
        \SB2_2_29/i0[10] ), .A3(\SB2_2_29/i1[9] ), .ZN(
        \SB2_2_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_3/N3  ( .A1(\SB2_2_29/i1[9] ), .A2(
        \SB2_2_29/i1_7 ), .A3(\SB2_2_29/i0[10] ), .ZN(
        \SB2_2_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_29/Component_Function_4/N4  ( .A1(\SB2_2_29/i1[9] ), .A2(
        \SB2_2_29/i1_5 ), .A3(\SB2_2_29/i0_4 ), .ZN(
        \SB2_2_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_29/Component_Function_4/N1  ( .A1(\SB2_2_29/i0[9] ), .A2(
        \SB2_2_29/i0_0 ), .A3(\SB2_2_29/i0[8] ), .ZN(
        \SB2_2_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_4/N2  ( .A1(\SB2_2_30/i3[0] ), .A2(
        \SB2_2_30/i0_0 ), .A3(\SB2_2_30/i1_7 ), .ZN(
        \SB2_2_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_30/Component_Function_4/N1  ( .A1(\SB2_2_30/i0[9] ), .A2(
        \SB2_2_30/i0_0 ), .A3(\SB2_2_30/i0[8] ), .ZN(
        \SB2_2_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_31/Component_Function_4/N2  ( .A1(\SB2_2_31/i3[0] ), .A2(
        \SB2_2_31/i0_0 ), .A3(\SB2_2_31/i1_7 ), .ZN(
        \SB2_2_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_31/Component_Function_4/N1  ( .A1(\SB2_2_31/i0[9] ), .A2(
        \SB2_2_31/i0_0 ), .A3(\SB2_2_31/i0[8] ), .ZN(
        \SB2_2_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_2/N1  ( .A1(\SB1_3_0/i1_5 ), .A2(
        \SB1_3_0/i0[10] ), .A3(\SB1_3_0/i1[9] ), .ZN(
        \SB1_3_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_4/N2  ( .A1(\SB1_3_0/i3[0] ), .A2(
        \SB1_3_0/i0_0 ), .A3(\SB1_3_0/i1_7 ), .ZN(
        \SB1_3_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_0/Component_Function_4/N1  ( .A1(\SB1_3_0/i0[9] ), .A2(
        \SB1_3_0/i0_0 ), .A3(\SB1_3_0/i0[8] ), .ZN(
        \SB1_3_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_3/N1  ( .A1(\SB1_3_1/i1[9] ), .A2(
        \SB1_3_1/i0_3 ), .A3(\SB1_3_1/i0[6] ), .ZN(
        \SB1_3_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_4/N4  ( .A1(\SB1_3_1/i1[9] ), .A2(
        \SB1_3_1/i1_5 ), .A3(\SB1_3_1/i0_4 ), .ZN(
        \SB1_3_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_2/Component_Function_2/N2  ( .A1(\SB1_3_2/i0_3 ), .A2(
        \SB1_3_2/i0[10] ), .A3(\SB1_3_2/i0[6] ), .ZN(
        \SB1_3_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_4/N2  ( .A1(\SB1_3_2/i3[0] ), .A2(
        \SB1_3_2/i0_0 ), .A3(\SB1_3_2/i1_7 ), .ZN(
        \SB1_3_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_4/N1  ( .A1(\SB1_3_2/i0[9] ), .A2(
        \SB1_3_2/i0_0 ), .A3(\SB1_3_2/i0[8] ), .ZN(
        \SB1_3_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_4/N2  ( .A1(\SB1_3_3/i3[0] ), .A2(
        \SB1_3_3/i0_0 ), .A3(\SB1_3_3/i1_7 ), .ZN(
        \SB1_3_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_3/Component_Function_4/N1  ( .A1(\SB1_3_3/i0[9] ), .A2(
        \SB1_3_3/i0_0 ), .A3(\SB1_3_3/i0[8] ), .ZN(
        \SB1_3_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_4/Component_Function_3/N4  ( .A1(\SB1_3_4/i1_5 ), .A2(
        \SB1_3_4/i0[8] ), .A3(\SB1_3_4/i3[0] ), .ZN(
        \SB1_3_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_4/Component_Function_3/N1  ( .A1(\SB1_3_4/i1[9] ), .A2(
        \RI1[3][167] ), .A3(\SB1_3_4/i0[6] ), .ZN(
        \SB1_3_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_2/N1  ( .A1(\SB1_3_5/i1_5 ), .A2(
        \SB1_3_5/i0[10] ), .A3(\SB1_3_5/i1[9] ), .ZN(
        \SB1_3_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_3/N3  ( .A1(\SB1_3_5/i1[9] ), .A2(
        \SB1_3_5/i1_7 ), .A3(\SB1_3_5/i0[10] ), .ZN(
        \SB1_3_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_7/Component_Function_4/N1  ( .A1(\SB1_3_7/i0[9] ), .A2(
        \SB1_3_7/i0_0 ), .A3(\SB1_3_7/i0[8] ), .ZN(
        \SB1_3_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_8/Component_Function_4/N4  ( .A1(\SB1_3_8/i1[9] ), .A2(
        \SB1_3_8/i1_5 ), .A3(\SB1_3_8/i0_4 ), .ZN(
        \SB1_3_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_9/Component_Function_2/N3  ( .A1(\SB1_3_9/i0_3 ), .A2(
        \SB1_3_9/i0[8] ), .A3(\MC_ARK_ARC_1_2/buf_output[132] ), .ZN(
        \SB1_3_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_9/Component_Function_2/N1  ( .A1(\SB1_3_9/i1_5 ), .A2(
        \SB1_3_9/i0[10] ), .A3(\SB1_3_9/i1[9] ), .ZN(
        \SB1_3_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_4/N2  ( .A1(\SB1_3_9/i3[0] ), .A2(
        \SB1_3_9/i0_0 ), .A3(\SB1_3_9/i1_7 ), .ZN(
        \SB1_3_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_10/Component_Function_2/N4  ( .A1(\SB1_3_10/i1_5 ), .A2(
        \SB1_3_10/i0_0 ), .A3(\SB1_3_10/i0_4 ), .ZN(
        \SB1_3_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_13/Component_Function_3/N2  ( .A1(\SB1_3_13/i0_0 ), .A2(
        \SB1_3_13/i0_3 ), .A3(\SB1_3_13/i0_4 ), .ZN(
        \SB1_3_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_14/Component_Function_3/N4  ( .A1(\SB1_3_14/i1_5 ), .A2(
        \SB1_3_14/i0[8] ), .A3(\SB1_3_14/i3[0] ), .ZN(
        \SB1_3_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_15/Component_Function_4/N2  ( .A1(\SB1_3_15/i3[0] ), .A2(
        \SB1_3_15/i0_0 ), .A3(\SB1_3_15/i1_7 ), .ZN(
        \SB1_3_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_18/Component_Function_2/N2  ( .A1(\SB1_3_18/i0_3 ), .A2(
        \SB1_3_18/i0[10] ), .A3(\SB1_3_18/i0[6] ), .ZN(
        \SB1_3_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_18/Component_Function_3/N2  ( .A1(\SB1_3_18/i0_0 ), .A2(
        \SB1_3_18/i0_3 ), .A3(\SB1_3_18/i0_4 ), .ZN(
        \SB1_3_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_18/Component_Function_3/N1  ( .A1(\SB1_3_18/i1[9] ), .A2(
        \SB1_3_18/i0_3 ), .A3(\SB1_3_18/i0[6] ), .ZN(
        \SB1_3_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_4/N2  ( .A1(\SB1_3_18/i3[0] ), .A2(
        \SB1_3_18/i0_0 ), .A3(\SB1_3_18/i1_7 ), .ZN(
        \SB1_3_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_19/Component_Function_2/N1  ( .A1(\SB1_3_19/i1_5 ), .A2(
        \SB1_3_19/i0[10] ), .A3(\SB1_3_19/i1[9] ), .ZN(
        \SB1_3_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_3/N1  ( .A1(\SB1_3_19/i1[9] ), .A2(
        \SB1_3_19/i0_3 ), .A3(\SB1_3_19/i0[6] ), .ZN(
        \SB1_3_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_4/N1  ( .A1(\SB1_3_19/i0[9] ), .A2(
        \SB1_3_19/i0_0 ), .A3(\SB1_3_19/i0[8] ), .ZN(
        \SB1_3_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_4/N1  ( .A1(\SB1_3_20/i0[9] ), .A2(
        \SB1_3_20/i0_0 ), .A3(\SB1_3_20/i0[8] ), .ZN(
        \SB1_3_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_2/N2  ( .A1(n3987), .A2(
        \SB1_3_21/i0[10] ), .A3(\SB1_3_21/i0[6] ), .ZN(
        \SB1_3_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_21/Component_Function_2/N1  ( .A1(\SB1_3_21/i1_5 ), .A2(
        \SB1_3_21/i0[10] ), .A3(\SB1_3_21/i1[9] ), .ZN(
        \SB1_3_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_3/N1  ( .A1(\SB1_3_21/i1[9] ), .A2(
        \SB1_3_21/i0_3 ), .A3(\SB1_3_21/i0[6] ), .ZN(
        \SB1_3_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_22/Component_Function_2/N2  ( .A1(\SB1_3_22/i0_3 ), .A2(
        \SB1_3_22/i0[10] ), .A3(\SB1_3_22/i0[6] ), .ZN(
        \SB1_3_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_22/Component_Function_3/N1  ( .A1(\SB1_3_22/i1[9] ), .A2(
        \SB1_3_22/i0_3 ), .A3(\SB1_3_22/i0[6] ), .ZN(
        \SB1_3_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_24/Component_Function_4/N1  ( .A1(\SB1_3_24/i0[9] ), .A2(
        \SB1_3_24/i0_0 ), .A3(\SB1_3_24/i0[8] ), .ZN(
        \SB1_3_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_2/N1  ( .A1(\SB1_3_25/i1_5 ), .A2(
        \SB1_3_25/i0[10] ), .A3(\SB1_3_25/i1[9] ), .ZN(
        \SB1_3_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_3/N3  ( .A1(\SB1_3_25/i1[9] ), .A2(
        \SB1_3_25/i1_7 ), .A3(\SB1_3_25/i0[10] ), .ZN(
        \SB1_3_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_25/Component_Function_4/N1  ( .A1(\SB1_3_25/i0[9] ), .A2(
        \SB1_3_25/i0_0 ), .A3(\SB1_3_25/i0[8] ), .ZN(
        \SB1_3_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_4/N2  ( .A1(\SB1_3_26/i3[0] ), .A2(
        \SB1_3_26/i0_0 ), .A3(\SB1_3_26/i1_7 ), .ZN(
        \SB1_3_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_26/Component_Function_4/N1  ( .A1(\SB1_3_26/i0[9] ), .A2(
        \SB1_3_26/i0_0 ), .A3(\SB1_3_26/i0[8] ), .ZN(
        \SB1_3_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_2/N2  ( .A1(\SB1_3_27/i0_3 ), .A2(
        \SB1_3_27/i0[10] ), .A3(\SB1_3_27/i0[6] ), .ZN(
        \SB1_3_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N2  ( .A1(\SB1_3_28/i3[0] ), .A2(
        \SB1_3_28/i0_0 ), .A3(\SB1_3_28/i1_7 ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N1  ( .A1(\SB1_3_28/i0[9] ), .A2(
        \SB1_3_28/i0_0 ), .A3(\SB1_3_28/i0[8] ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_3/N1  ( .A1(\SB1_3_29/i1[9] ), .A2(
        \SB1_3_29/i0_3 ), .A3(\SB1_3_29/i0[6] ), .ZN(
        \SB1_3_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_2/N2  ( .A1(\SB1_3_30/i0_3 ), .A2(
        \SB1_3_30/i0[10] ), .A3(\SB1_3_30/i0[6] ), .ZN(
        \SB1_3_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_30/Component_Function_3/N2  ( .A1(\SB1_3_30/i0_0 ), .A2(
        \SB1_3_30/i0_3 ), .A3(\SB1_3_30/i0_4 ), .ZN(
        \SB1_3_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_30/Component_Function_4/N2  ( .A1(\SB1_3_30/i3[0] ), .A2(
        \SB1_3_30/i0_0 ), .A3(\SB1_3_30/i1_7 ), .ZN(
        \SB1_3_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_30/Component_Function_4/N1  ( .A1(\SB1_3_30/i0[9] ), .A2(
        \SB1_3_30/i0_0 ), .A3(\SB1_3_30/i0[8] ), .ZN(
        \SB1_3_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_3/N3  ( .A1(\SB2_3_1/i1[9] ), .A2(
        \SB2_3_1/i1_7 ), .A3(\SB2_3_1/i0[10] ), .ZN(
        \SB2_3_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_1/Component_Function_3/N1  ( .A1(\SB2_3_1/i1[9] ), .A2(
        \SB2_3_1/i0_3 ), .A3(\SB2_3_1/i0[6] ), .ZN(
        \SB2_3_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_4/N1  ( .A1(\SB2_3_1/i0[9] ), .A2(
        \SB2_3_1/i0_0 ), .A3(\SB2_3_1/i0[8] ), .ZN(
        \SB2_3_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_3/Component_Function_4/N2  ( .A1(\SB2_3_3/i3[0] ), .A2(
        \SB2_3_3/i0_0 ), .A3(\SB2_3_3/i1_7 ), .ZN(
        \SB2_3_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_4/Component_Function_2/N2  ( .A1(\SB2_3_4/i0_3 ), .A2(
        \SB2_3_4/i0[10] ), .A3(\SB2_3_4/i0[6] ), .ZN(
        \SB2_3_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_4/Component_Function_4/N4  ( .A1(\SB2_3_4/i1[9] ), .A2(
        \SB2_3_4/i1_5 ), .A3(\SB2_3_4/i0_4 ), .ZN(
        \SB2_3_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_4/Component_Function_4/N2  ( .A1(\SB2_3_4/i3[0] ), .A2(
        \SB2_3_4/i0_0 ), .A3(\SB2_3_4/i1_7 ), .ZN(
        \SB2_3_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_4/Component_Function_4/N1  ( .A1(\SB2_3_4/i0[9] ), .A2(
        \SB2_3_4/i0_0 ), .A3(\SB2_3_4/i0[8] ), .ZN(
        \SB2_3_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_5/Component_Function_3/N4  ( .A1(\SB2_3_5/i1_5 ), .A2(
        \SB2_3_5/i0[8] ), .A3(\SB2_3_5/i3[0] ), .ZN(
        \SB2_3_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_5/Component_Function_4/N2  ( .A1(\SB2_3_5/i3[0] ), .A2(
        \SB2_3_5/i0_0 ), .A3(\SB2_3_5/i1_7 ), .ZN(
        \SB2_3_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_5/Component_Function_4/N1  ( .A1(\SB2_3_5/i0[9] ), .A2(
        \SB2_3_5/i0_0 ), .A3(\SB2_3_5/i0[8] ), .ZN(
        \SB2_3_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_6/Component_Function_4/N4  ( .A1(\SB2_3_6/i1[9] ), .A2(
        \SB2_3_6/i1_5 ), .A3(\SB2_3_6/i0_4 ), .ZN(
        \SB2_3_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_6/Component_Function_4/N2  ( .A1(\SB2_3_6/i3[0] ), .A2(
        \SB2_3_6/i0_0 ), .A3(\SB2_3_6/i1_7 ), .ZN(
        \SB2_3_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_6/Component_Function_4/N1  ( .A1(\SB2_3_6/i0[9] ), .A2(
        \SB2_3_6/i0_0 ), .A3(\SB2_3_6/i0[8] ), .ZN(
        \SB2_3_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_4/N2  ( .A1(\SB2_3_7/i3[0] ), .A2(
        \SB2_3_7/i0_0 ), .A3(\SB2_3_7/i1_7 ), .ZN(
        \SB2_3_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_7/Component_Function_4/N1  ( .A1(\SB2_3_7/i0[9] ), .A2(
        \SB2_3_7/i0_0 ), .A3(\SB2_3_7/i0[8] ), .ZN(
        \SB2_3_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_8/Component_Function_4/N1  ( .A1(\SB2_3_8/i0[9] ), .A2(
        \SB2_3_8/i0_0 ), .A3(\SB2_3_8/i0[8] ), .ZN(
        \SB2_3_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_4/N4  ( .A1(\SB2_3_10/i1[9] ), .A2(
        \SB2_3_10/i1_5 ), .A3(\SB2_3_10/i0_4 ), .ZN(
        \SB2_3_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_10/Component_Function_4/N1  ( .A1(\SB2_3_10/i0[9] ), .A2(
        \SB2_3_10/i0_0 ), .A3(\SB2_3_10/i0[8] ), .ZN(
        \SB2_3_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_11/Component_Function_4/N1  ( .A1(\SB2_3_11/i0[9] ), .A2(
        \SB2_3_11/i0_0 ), .A3(\SB2_3_11/i0[8] ), .ZN(
        \SB2_3_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_4/N2  ( .A1(\SB2_3_12/i3[0] ), .A2(
        \SB2_3_12/i0_0 ), .A3(\SB2_3_12/i1_7 ), .ZN(
        \SB2_3_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_13/Component_Function_4/N1  ( .A1(\SB2_3_13/i0[9] ), .A2(
        \SB2_3_13/i0_0 ), .A3(\SB2_3_13/i0[8] ), .ZN(
        \SB2_3_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_4/N2  ( .A1(\SB2_3_14/i3[0] ), .A2(
        \SB2_3_14/i0_0 ), .A3(\SB2_3_14/i1_7 ), .ZN(
        \SB2_3_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_14/Component_Function_4/N1  ( .A1(\SB2_3_14/i0[9] ), .A2(
        \SB2_3_14/i0_0 ), .A3(\SB2_3_14/i0[8] ), .ZN(
        \SB2_3_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_4/N4  ( .A1(\SB2_3_15/i1[9] ), .A2(
        \SB2_3_15/i1_5 ), .A3(\SB1_3_16/buf_output[4] ), .ZN(
        \SB2_3_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_16/Component_Function_4/N2  ( .A1(\SB2_3_16/i3[0] ), .A2(
        \SB2_3_16/i0_0 ), .A3(\SB2_3_16/i1_7 ), .ZN(
        \SB2_3_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_16/Component_Function_4/N1  ( .A1(\SB2_3_16/i0[9] ), .A2(
        \SB2_3_16/i0_0 ), .A3(\SB2_3_16/i0[8] ), .ZN(
        \SB2_3_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_17/Component_Function_4/N1  ( .A1(\SB2_3_17/i0[9] ), .A2(
        \SB2_3_17/i0_0 ), .A3(\SB2_3_17/i0[8] ), .ZN(
        \SB2_3_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_4/N2  ( .A1(\SB2_3_18/i3[0] ), .A2(
        \SB2_3_18/i0_0 ), .A3(\SB2_3_18/i1_7 ), .ZN(
        \SB2_3_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_18/Component_Function_4/N1  ( .A1(\SB2_3_18/i0[9] ), .A2(
        \SB2_3_18/i0_0 ), .A3(\SB2_3_18/i0[8] ), .ZN(
        \SB2_3_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_19/Component_Function_4/N2  ( .A1(\SB2_3_19/i3[0] ), .A2(
        \SB2_3_19/i0_0 ), .A3(\SB2_3_19/i1_7 ), .ZN(
        \SB2_3_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_19/Component_Function_4/N1  ( .A1(\SB2_3_19/i0[9] ), .A2(
        \SB2_3_19/i0_0 ), .A3(\SB2_3_19/i0[8] ), .ZN(
        \SB2_3_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_20/Component_Function_4/N1  ( .A1(\SB2_3_20/i0[9] ), .A2(
        \SB2_3_20/i0_0 ), .A3(\SB2_3_20/i0[8] ), .ZN(
        \SB2_3_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_4/N3  ( .A1(\SB2_3_22/i0[9] ), .A2(
        \SB2_3_22/i0[10] ), .A3(\SB2_3_22/i0_3 ), .ZN(
        \SB2_3_22/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_23/Component_Function_4/N4  ( .A1(\SB2_3_23/i1[9] ), .A2(
        \SB2_3_23/i1_5 ), .A3(\SB2_3_23/i0_4 ), .ZN(
        \SB2_3_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_23/Component_Function_4/N1  ( .A1(\SB2_3_23/i0[9] ), .A2(
        \SB2_3_23/i0_0 ), .A3(\SB2_3_23/i0[8] ), .ZN(
        \SB2_3_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_24/Component_Function_4/N2  ( .A1(\SB2_3_24/i3[0] ), .A2(
        \SB2_3_24/i0_0 ), .A3(\SB2_3_24/i1_7 ), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_24/Component_Function_4/N1  ( .A1(\SB2_3_24/i0[9] ), .A2(
        \SB2_3_24/i0_0 ), .A3(\SB2_3_24/i0[8] ), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_4/N2  ( .A1(\SB2_3_26/i3[0] ), .A2(
        \SB2_3_26/i0_0 ), .A3(\SB2_3_26/i1_7 ), .ZN(
        \SB2_3_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_26/Component_Function_4/N1  ( .A1(\SB2_3_26/i0[9] ), .A2(
        \SB2_3_26/i0_0 ), .A3(\SB2_3_26/i0[8] ), .ZN(
        \SB2_3_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_4/N2  ( .A1(\SB2_3_27/i3[0] ), .A2(
        \SB2_3_27/i0_0 ), .A3(\SB2_3_27/i1_7 ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_27/Component_Function_4/N1  ( .A1(\SB2_3_27/i0[9] ), .A2(
        \SB2_3_27/i0_0 ), .A3(\SB2_3_27/i0[8] ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_29/Component_Function_4/N1  ( .A1(\SB2_3_29/i0[9] ), .A2(
        \SB2_3_29/i0_0 ), .A3(\SB2_3_29/i0[8] ), .ZN(
        \SB2_3_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_4/N2  ( .A1(\SB2_3_30/i3[0] ), .A2(
        \SB2_3_30/i0_0 ), .A3(\SB2_3_30/i1_7 ), .ZN(
        \SB2_3_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_30/Component_Function_4/N1  ( .A1(\SB2_3_30/i0[9] ), .A2(
        \SB2_3_30/i0_0 ), .A3(\SB2_3_30/i0[8] ), .ZN(
        \SB2_3_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_31/Component_Function_4/N2  ( .A1(\SB2_3_31/i3[0] ), .A2(
        \SB2_3_31/i0_0 ), .A3(\SB2_3_31/i1_7 ), .ZN(
        \SB2_3_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_1/Component_Function_2/N1  ( .A1(\SB1_4_1/i1_5 ), .A2(
        \SB1_4_1/i0[10] ), .A3(\SB1_4_1/i1[9] ), .ZN(
        \SB1_4_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_1/Component_Function_3/N1  ( .A1(\SB1_4_1/i1[9] ), .A2(
        \SB1_4_1/i0_3 ), .A3(\SB1_4_1/i0[6] ), .ZN(
        \SB1_4_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_1/Component_Function_4/N1  ( .A1(\SB1_4_1/i0[9] ), .A2(
        \SB1_4_1/i0_0 ), .A3(\SB1_4_1/i0[8] ), .ZN(
        \SB1_4_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_2/Component_Function_3/N2  ( .A1(\SB1_4_2/i0_0 ), .A2(
        \SB1_4_2/i0_3 ), .A3(\SB1_4_2/i0_4 ), .ZN(
        \SB1_4_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_3/Component_Function_2/N2  ( .A1(\SB1_4_3/i0_3 ), .A2(
        \SB1_4_3/i0[10] ), .A3(\SB1_4_3/i0[6] ), .ZN(
        \SB1_4_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_3/Component_Function_4/N2  ( .A1(\SB1_4_3/i3[0] ), .A2(
        \SB1_4_3/i0_0 ), .A3(\SB1_4_3/i1_7 ), .ZN(
        \SB1_4_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_3/Component_Function_4/N1  ( .A1(\SB1_4_3/i0[9] ), .A2(
        \SB1_4_3/i0_0 ), .A3(\SB1_4_3/i0[8] ), .ZN(
        \SB1_4_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_4/Component_Function_2/N1  ( .A1(\SB1_4_4/i1_5 ), .A2(
        \SB1_4_4/i0[10] ), .A3(\SB1_4_4/i1[9] ), .ZN(
        \SB1_4_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_4/Component_Function_3/N2  ( .A1(\SB1_4_4/i0_0 ), .A2(
        \SB1_4_4/i0_3 ), .A3(\SB1_4_4/i0_4 ), .ZN(
        \SB1_4_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_4/Component_Function_4/N2  ( .A1(\SB1_4_4/i3[0] ), .A2(
        \SB1_4_4/i0_0 ), .A3(\SB1_4_4/i1_7 ), .ZN(
        \SB1_4_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_4/Component_Function_4/N1  ( .A1(\SB1_4_4/i0[9] ), .A2(
        \SB1_4_4/i0_0 ), .A3(\SB1_4_4/i0[8] ), .ZN(
        \SB1_4_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_5/Component_Function_2/N3  ( .A1(\SB1_4_5/i0_3 ), .A2(
        \SB1_4_5/i0[8] ), .A3(\SB1_4_5/i0[9] ), .ZN(
        \SB1_4_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_5/Component_Function_2/N1  ( .A1(\SB1_4_5/i1_5 ), .A2(
        \SB1_4_5/i0[10] ), .A3(\SB1_4_5/i1[9] ), .ZN(
        \SB1_4_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_5/Component_Function_3/N2  ( .A1(\SB1_4_5/i0_0 ), .A2(
        \SB1_4_5/i0_3 ), .A3(\SB1_4_5/i0_4 ), .ZN(
        \SB1_4_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_5/Component_Function_3/N1  ( .A1(\SB1_4_5/i1[9] ), .A2(
        \SB1_4_5/i0_3 ), .A3(\SB1_4_5/i0[6] ), .ZN(
        \SB1_4_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_5/Component_Function_4/N4  ( .A1(\SB1_4_5/i1[9] ), .A2(
        \SB1_4_5/i1_5 ), .A3(\SB1_4_5/i0_4 ), .ZN(
        \SB1_4_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_5/Component_Function_4/N2  ( .A1(\SB1_4_5/i3[0] ), .A2(
        \SB1_4_5/i0_0 ), .A3(\SB1_4_5/i1_7 ), .ZN(
        \SB1_4_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_5/Component_Function_4/N1  ( .A1(\SB1_4_5/i0[9] ), .A2(
        \SB1_4_5/i0_0 ), .A3(\SB1_4_5/i0[8] ), .ZN(
        \SB1_4_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_7/Component_Function_2/N3  ( .A1(\SB1_4_7/i0_3 ), .A2(
        \SB1_4_7/i0[8] ), .A3(\SB1_4_7/i0[9] ), .ZN(
        \SB1_4_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_7/Component_Function_4/N2  ( .A1(\SB1_4_7/i3[0] ), .A2(
        \SB1_4_7/i0_0 ), .A3(\SB1_4_7/i1_7 ), .ZN(
        \SB1_4_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_7/Component_Function_4/N1  ( .A1(\SB1_4_7/i0[9] ), .A2(
        \SB1_4_7/i0_0 ), .A3(\SB1_4_7/i0[8] ), .ZN(
        \SB1_4_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_8/Component_Function_4/N4  ( .A1(\SB1_4_8/i1[9] ), .A2(
        \SB1_4_8/i1_5 ), .A3(\SB1_4_8/i0_4 ), .ZN(
        \SB1_4_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_9/Component_Function_2/N1  ( .A1(\SB1_4_9/i1_5 ), .A2(
        \SB1_4_9/i0[10] ), .A3(\SB1_4_9/i1[9] ), .ZN(
        \SB1_4_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_9/Component_Function_4/N1  ( .A1(\SB1_4_9/i0[9] ), .A2(
        \SB1_4_9/i0_0 ), .A3(\SB1_4_9/i0[8] ), .ZN(
        \SB1_4_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_10/Component_Function_3/N1  ( .A1(\SB1_4_10/i1[9] ), .A2(
        \RI1[4][131] ), .A3(\SB1_4_10/i0[6] ), .ZN(
        \SB1_4_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_10/Component_Function_4/N1  ( .A1(\SB1_4_10/i0[9] ), .A2(
        \SB1_4_10/i0_0 ), .A3(\SB1_4_10/i0[8] ), .ZN(
        \SB1_4_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_11/Component_Function_2/N1  ( .A1(\SB1_4_11/i1_5 ), .A2(
        \SB1_4_11/i0[10] ), .A3(\SB1_4_11/i1[9] ), .ZN(
        \SB1_4_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_11/Component_Function_4/N2  ( .A1(\SB1_4_11/i3[0] ), .A2(
        \SB1_4_11/i0_0 ), .A3(\SB1_4_11/i1_7 ), .ZN(
        \SB1_4_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_11/Component_Function_4/N1  ( .A1(\SB1_4_11/i0[9] ), .A2(
        \SB1_4_11/i0_0 ), .A3(\SB1_4_11/i0[8] ), .ZN(
        \SB1_4_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_13/Component_Function_2/N2  ( .A1(\SB1_4_13/i0_3 ), .A2(
        \SB1_4_13/i0[10] ), .A3(\SB1_4_13/i0[6] ), .ZN(
        \SB1_4_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_13/Component_Function_4/N4  ( .A1(\SB1_4_13/i1[9] ), .A2(
        \SB1_4_13/i1_5 ), .A3(\SB1_4_13/i0_4 ), .ZN(
        \SB1_4_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_16/Component_Function_2/N2  ( .A1(\SB1_4_16/i0_3 ), .A2(
        \SB1_4_16/i0[10] ), .A3(\SB1_4_16/i0[6] ), .ZN(
        \SB1_4_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_17/Component_Function_2/N1  ( .A1(\SB1_4_17/i1_5 ), .A2(
        \SB1_4_17/i0[10] ), .A3(\SB1_4_17/i1[9] ), .ZN(
        \SB1_4_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_17/Component_Function_3/N2  ( .A1(\SB1_4_17/i0_0 ), .A2(
        \SB1_4_17/i0_3 ), .A3(\SB1_4_17/i0_4 ), .ZN(
        \SB1_4_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_17/Component_Function_4/N1  ( .A1(\SB1_4_17/i0[9] ), .A2(
        \SB1_4_17/i0_0 ), .A3(\SB1_4_17/i0[8] ), .ZN(
        \SB1_4_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_18/Component_Function_2/N2  ( .A1(\SB1_4_18/i0_3 ), .A2(
        \SB1_4_18/i0[10] ), .A3(\SB1_4_18/i0[6] ), .ZN(
        \SB1_4_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_18/Component_Function_4/N2  ( .A1(\SB1_4_18/i3[0] ), .A2(
        \SB1_4_18/i0_0 ), .A3(\SB1_4_18/i1_7 ), .ZN(
        \SB1_4_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_19/Component_Function_4/N1  ( .A1(\SB1_4_19/i0[9] ), .A2(
        \SB1_4_19/i0_0 ), .A3(\SB1_4_19/i0[8] ), .ZN(
        \SB1_4_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_20/Component_Function_4/N2  ( .A1(\SB1_4_20/i3[0] ), .A2(
        \SB1_4_20/i0_0 ), .A3(\SB1_4_20/i1_7 ), .ZN(
        \SB1_4_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_20/Component_Function_4/N1  ( .A1(\SB1_4_20/i0[9] ), .A2(
        \SB1_4_20/i0_0 ), .A3(\SB1_4_20/i0[8] ), .ZN(
        \SB1_4_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_21/Component_Function_3/N2  ( .A1(\SB1_4_21/i0_0 ), .A2(
        \SB1_4_21/i0_3 ), .A3(\SB1_4_21/i0_4 ), .ZN(
        \SB1_4_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_21/Component_Function_3/N1  ( .A1(\SB1_4_21/i1[9] ), .A2(
        \SB1_4_21/i0_3 ), .A3(\SB1_4_21/i0[6] ), .ZN(
        \SB1_4_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_21/Component_Function_4/N2  ( .A1(\SB1_4_21/i3[0] ), .A2(
        \SB1_4_21/i0_0 ), .A3(\SB1_4_21/i1_7 ), .ZN(
        \SB1_4_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_22/Component_Function_4/N2  ( .A1(\SB1_4_22/i3[0] ), .A2(
        \SB1_4_22/i0_0 ), .A3(\SB1_4_22/i1_7 ), .ZN(
        \SB1_4_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_23/Component_Function_2/N4  ( .A1(\SB1_4_23/i1_5 ), .A2(
        \SB1_4_23/i0_0 ), .A3(\SB1_4_23/i0_4 ), .ZN(
        \SB1_4_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_23/Component_Function_2/N2  ( .A1(\SB1_4_23/i0_3 ), .A2(
        \SB1_4_23/i0[10] ), .A3(\SB1_4_23/i0[6] ), .ZN(
        \SB1_4_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_23/Component_Function_3/N2  ( .A1(\SB1_4_23/i0_0 ), .A2(
        \SB1_4_23/i0_3 ), .A3(\SB1_4_23/i0_4 ), .ZN(
        \SB1_4_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_23/Component_Function_3/N1  ( .A1(\SB1_4_23/i1[9] ), .A2(
        \SB1_4_23/i0_3 ), .A3(\SB1_4_23/i0[6] ), .ZN(
        \SB1_4_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_23/Component_Function_4/N2  ( .A1(\SB1_4_23/i3[0] ), .A2(
        \SB1_4_23/i0_0 ), .A3(\SB1_4_23/i1_7 ), .ZN(
        \SB1_4_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_26/Component_Function_4/N2  ( .A1(\SB1_4_26/i3[0] ), .A2(
        \SB1_4_26/i0_0 ), .A3(\SB1_4_26/i1_7 ), .ZN(
        \SB1_4_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_26/Component_Function_4/N1  ( .A1(\SB1_4_26/i0[9] ), .A2(
        \SB1_4_26/i0_0 ), .A3(\SB1_4_26/i0[8] ), .ZN(
        \SB1_4_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_27/Component_Function_3/N1  ( .A1(\SB1_4_27/i1[9] ), .A2(
        \SB1_4_27/i0_3 ), .A3(\SB1_4_27/i0[6] ), .ZN(
        \SB1_4_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_28/Component_Function_2/N2  ( .A1(\SB1_4_28/i0_3 ), .A2(
        \SB1_4_28/i0[10] ), .A3(\SB1_4_28/i0[6] ), .ZN(
        \SB1_4_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_28/Component_Function_4/N2  ( .A1(\SB1_4_28/i3[0] ), .A2(
        \SB1_4_28/i0_0 ), .A3(\SB1_4_28/i1_7 ), .ZN(
        \SB1_4_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_28/Component_Function_4/N1  ( .A1(\SB1_4_28/i0[9] ), .A2(
        \SB1_4_28/i0_0 ), .A3(\SB1_4_28/i0[8] ), .ZN(
        \SB1_4_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_29/Component_Function_2/N1  ( .A1(\SB1_4_29/i1_5 ), .A2(
        \SB1_4_29/i0[10] ), .A3(\SB1_4_29/i1[9] ), .ZN(
        \SB1_4_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_29/Component_Function_4/N1  ( .A1(\SB1_4_29/i0[9] ), .A2(
        \SB1_4_29/i0_0 ), .A3(\SB1_4_29/i0[8] ), .ZN(
        \SB1_4_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_30/Component_Function_4/N1  ( .A1(\SB1_4_30/i0[9] ), .A2(
        \SB1_4_30/i0_0 ), .A3(\SB1_4_30/i0[8] ), .ZN(
        \SB1_4_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_31/Component_Function_2/N1  ( .A1(\SB1_4_31/i1_5 ), .A2(
        \SB1_4_31/i0[10] ), .A3(\SB1_4_31/i1[9] ), .ZN(
        \SB1_4_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_31/Component_Function_4/N2  ( .A1(\SB1_4_31/i3[0] ), .A2(
        \SB1_4_31/i0_0 ), .A3(\SB1_4_31/i1_7 ), .ZN(
        \SB1_4_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_0/Component_Function_2/N1  ( .A1(n3978), .A2(
        \SB2_4_0/i0[10] ), .A3(\SB2_4_0/i1[9] ), .ZN(
        \SB2_4_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_0/Component_Function_3/N1  ( .A1(\SB2_4_0/i1[9] ), .A2(
        \SB1_4_0/buf_output[5] ), .A3(\SB2_4_0/i0[6] ), .ZN(
        \SB2_4_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_0/Component_Function_4/N4  ( .A1(\SB2_4_0/i1[9] ), .A2(n3978), .A3(\SB2_4_0/i0_4 ), .ZN(\SB2_4_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_0/Component_Function_4/N1  ( .A1(\SB2_4_0/i0[9] ), .A2(
        \SB2_4_0/i0_0 ), .A3(\SB2_4_0/i0[8] ), .ZN(
        \SB2_4_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_1/Component_Function_4/N2  ( .A1(\SB2_4_1/i3[0] ), .A2(
        \SB2_4_1/i0_0 ), .A3(\SB2_4_1/i1_7 ), .ZN(
        \SB2_4_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_1/Component_Function_4/N1  ( .A1(\SB2_4_1/i0[9] ), .A2(
        \SB2_4_1/i0_0 ), .A3(\SB2_4_1/i0[8] ), .ZN(
        \SB2_4_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_2/Component_Function_2/N1  ( .A1(\SB2_4_2/i1_5 ), .A2(
        \SB2_4_2/i0[10] ), .A3(\SB2_4_2/i1[9] ), .ZN(
        \SB2_4_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_2/Component_Function_4/N4  ( .A1(\SB2_4_2/i1[9] ), .A2(
        \SB2_4_2/i1_5 ), .A3(\SB2_4_2/i0_4 ), .ZN(
        \SB2_4_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_2/Component_Function_4/N2  ( .A1(\SB2_4_2/i3[0] ), .A2(
        \SB2_4_2/i0_0 ), .A3(\SB2_4_2/i1_7 ), .ZN(
        \SB2_4_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_2/Component_Function_4/N1  ( .A1(\SB2_4_2/i0[9] ), .A2(
        \SB2_4_2/i0_0 ), .A3(\SB2_4_2/i0[8] ), .ZN(
        \SB2_4_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_3/Component_Function_3/N4  ( .A1(n3988), .A2(\SB2_4_3/i0[8] ), .A3(\SB2_4_3/i3[0] ), .ZN(\SB2_4_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_3/Component_Function_4/N1  ( .A1(\SB2_4_3/i0[9] ), .A2(
        \SB2_4_3/i0_0 ), .A3(\SB2_4_3/i0[8] ), .ZN(
        \SB2_4_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_4/Component_Function_4/N2  ( .A1(\SB2_4_4/i3[0] ), .A2(
        \SB2_4_4/i0_0 ), .A3(\SB2_4_4/i1_7 ), .ZN(
        \SB2_4_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_5/Component_Function_4/N1  ( .A1(\SB2_4_5/i0[9] ), .A2(
        \SB2_4_5/i0_0 ), .A3(\SB2_4_5/i0[8] ), .ZN(
        \SB2_4_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_6/Component_Function_4/N2  ( .A1(\SB2_4_6/i3[0] ), .A2(
        \SB2_4_6/i0_0 ), .A3(\SB2_4_6/i1_7 ), .ZN(
        \SB2_4_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_7/Component_Function_4/N4  ( .A1(\SB2_4_7/i1[9] ), .A2(
        \SB2_4_7/i1_5 ), .A3(\RI3[4][148] ), .ZN(
        \SB2_4_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_7/Component_Function_4/N1  ( .A1(\SB2_4_7/i0[9] ), .A2(
        \SB2_4_7/i0_0 ), .A3(\SB2_4_7/i0[8] ), .ZN(
        \SB2_4_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_8/Component_Function_2/N1  ( .A1(\SB2_4_8/i1_5 ), .A2(
        \SB2_4_8/i0[10] ), .A3(\SB2_4_8/i1[9] ), .ZN(
        \SB2_4_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_8/Component_Function_4/N4  ( .A1(\SB2_4_8/i1[9] ), .A2(
        \SB2_4_8/i1_5 ), .A3(n3183), .ZN(
        \SB2_4_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_8/Component_Function_4/N1  ( .A1(\SB2_4_8/i0[9] ), .A2(
        \SB2_4_8/i0_0 ), .A3(\SB2_4_8/i0[8] ), .ZN(
        \SB2_4_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_9/Component_Function_4/N2  ( .A1(\SB2_4_9/i3[0] ), .A2(
        \SB2_4_9/i0_0 ), .A3(\SB2_4_9/i1_7 ), .ZN(
        \SB2_4_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_9/Component_Function_4/N1  ( .A1(\SB2_4_9/i0[9] ), .A2(
        \SB2_4_9/i0_0 ), .A3(\SB2_4_9/i0[8] ), .ZN(
        \SB2_4_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_10/Component_Function_4/N2  ( .A1(\SB2_4_10/i3[0] ), .A2(
        \SB2_4_10/i0_0 ), .A3(\SB2_4_10/i1_7 ), .ZN(
        \SB2_4_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_10/Component_Function_4/N1  ( .A1(\SB2_4_10/i0[9] ), .A2(
        \SB2_4_10/i0_0 ), .A3(\SB2_4_10/i0[8] ), .ZN(
        \SB2_4_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_11/Component_Function_4/N2  ( .A1(\SB2_4_11/i3[0] ), .A2(
        \SB2_4_11/i0_0 ), .A3(\SB2_4_11/i1_7 ), .ZN(
        \SB2_4_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_12/Component_Function_4/N1  ( .A1(\SB2_4_12/i0[9] ), .A2(
        \SB2_4_12/i0_0 ), .A3(\SB2_4_12/i0[8] ), .ZN(
        \SB2_4_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_13/Component_Function_4/N1  ( .A1(\SB2_4_13/i0[9] ), .A2(
        \SB2_4_13/i0_0 ), .A3(\SB2_4_13/i0[8] ), .ZN(
        \SB2_4_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_14/Component_Function_4/N1  ( .A1(\SB2_4_14/i0[9] ), .A2(
        \SB2_4_14/i0_0 ), .A3(\SB2_4_14/i0[8] ), .ZN(
        \SB2_4_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_15/Component_Function_4/N2  ( .A1(\SB2_4_15/i3[0] ), .A2(
        \SB2_4_15/i0_0 ), .A3(\SB2_4_15/i1_7 ), .ZN(
        \SB2_4_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_15/Component_Function_4/N1  ( .A1(\SB2_4_15/i0[9] ), .A2(
        \SB2_4_15/i0_0 ), .A3(\SB2_4_15/i0[8] ), .ZN(
        \SB2_4_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_16/Component_Function_4/N1  ( .A1(\SB2_4_16/i0[9] ), .A2(
        \SB2_4_16/i0_0 ), .A3(\SB2_4_16/i0[8] ), .ZN(
        \SB2_4_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_17/Component_Function_4/N4  ( .A1(\SB2_4_17/i1[9] ), .A2(
        \SB2_4_17/i1_5 ), .A3(\SB2_4_17/i0_4 ), .ZN(
        \SB2_4_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_17/Component_Function_4/N2  ( .A1(\SB2_4_17/i3[0] ), .A2(
        \SB2_4_17/i0_0 ), .A3(\SB2_4_17/i1_7 ), .ZN(
        \SB2_4_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_17/Component_Function_4/N1  ( .A1(\SB2_4_17/i0[9] ), .A2(
        \SB2_4_17/i0_0 ), .A3(\SB2_4_17/i0[8] ), .ZN(
        \SB2_4_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_18/Component_Function_4/N2  ( .A1(\SB2_4_18/i3[0] ), .A2(
        \SB2_4_18/i0_0 ), .A3(\SB2_4_18/i1_7 ), .ZN(
        \SB2_4_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_19/Component_Function_4/N1  ( .A1(\SB2_4_19/i0[9] ), .A2(
        \SB2_4_19/i0_0 ), .A3(\SB2_4_19/i0[8] ), .ZN(
        \SB2_4_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_20/Component_Function_4/N2  ( .A1(\SB2_4_20/i3[0] ), .A2(
        \SB2_4_20/i0_0 ), .A3(\SB2_4_20/i1_7 ), .ZN(
        \SB2_4_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_21/Component_Function_4/N1  ( .A1(\SB2_4_21/i0[9] ), .A2(
        \SB2_4_21/i0_0 ), .A3(\SB2_4_21/i0[8] ), .ZN(
        \SB2_4_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_22/Component_Function_4/N4  ( .A1(\SB2_4_22/i1[9] ), .A2(
        \SB2_4_22/i1_5 ), .A3(\SB2_4_22/i0_4 ), .ZN(
        \SB2_4_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_23/Component_Function_3/N1  ( .A1(\SB2_4_23/i1[9] ), .A2(
        \SB2_4_23/i0_3 ), .A3(\SB2_4_23/i0[6] ), .ZN(
        \SB2_4_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_24/Component_Function_4/N4  ( .A1(n5443), .A2(n6268), .A3(
        \SB2_4_24/i0_4 ), .ZN(\SB2_4_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_24/Component_Function_4/N2  ( .A1(\SB2_4_24/i3[0] ), .A2(
        \SB2_4_24/i0_0 ), .A3(\SB2_4_24/i1_7 ), .ZN(
        \SB2_4_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_24/Component_Function_4/N1  ( .A1(\SB2_4_24/i0[9] ), .A2(
        \SB2_4_24/i0_0 ), .A3(\SB2_4_24/i0[8] ), .ZN(
        \SB2_4_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_25/Component_Function_4/N1  ( .A1(\SB2_4_25/i0[9] ), .A2(
        \SB2_4_25/i0_0 ), .A3(\SB2_4_25/i0[8] ), .ZN(
        \SB2_4_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_26/Component_Function_2/N2  ( .A1(\SB2_4_26/i0_3 ), .A2(
        \SB2_4_26/i0[10] ), .A3(\SB2_4_26/i0[6] ), .ZN(
        \SB2_4_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_26/Component_Function_4/N2  ( .A1(\SB2_4_26/i3[0] ), .A2(
        \SB2_4_26/i0_0 ), .A3(\SB2_4_26/i1_7 ), .ZN(
        \SB2_4_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_26/Component_Function_4/N1  ( .A1(\SB2_4_26/i0[9] ), .A2(
        \SB2_4_26/i0_0 ), .A3(\SB2_4_26/i0[8] ), .ZN(
        \SB2_4_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_27/Component_Function_4/N4  ( .A1(\SB2_4_27/i1[9] ), .A2(
        \SB2_4_27/i1_5 ), .A3(\SB2_4_27/i0_4 ), .ZN(
        \SB2_4_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_27/Component_Function_4/N2  ( .A1(\SB2_4_27/i3[0] ), .A2(
        \SB2_4_27/i0_0 ), .A3(\SB2_4_27/i1_7 ), .ZN(
        \SB2_4_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_27/Component_Function_4/N1  ( .A1(\SB2_4_27/i0[9] ), .A2(
        \SB2_4_27/i0_0 ), .A3(\SB2_4_27/i0[8] ), .ZN(
        \SB2_4_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_28/Component_Function_4/N4  ( .A1(\SB2_4_28/i1[9] ), .A2(
        \SB2_4_28/i1_5 ), .A3(\SB2_4_28/i0_4 ), .ZN(
        \SB2_4_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_28/Component_Function_4/N2  ( .A1(\SB2_4_28/i3[0] ), .A2(
        \SB2_4_28/i0_0 ), .A3(\SB2_4_28/i1_7 ), .ZN(
        \SB2_4_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_29/Component_Function_3/N2  ( .A1(\SB2_4_29/i0_0 ), .A2(
        \SB2_4_29/i0_3 ), .A3(\SB2_4_29/i0_4 ), .ZN(
        \SB2_4_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_29/Component_Function_4/N1  ( .A1(\SB2_4_29/i0[9] ), .A2(
        \SB2_4_29/i0_0 ), .A3(\SB2_4_29/i0[8] ), .ZN(
        \SB2_4_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_30/Component_Function_4/N4  ( .A1(\SB2_4_30/i1[9] ), .A2(
        \SB2_4_30/i1_5 ), .A3(\SB1_4_31/buf_output[4] ), .ZN(
        \SB2_4_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_30/Component_Function_4/N2  ( .A1(n3983), .A2(
        \SB2_4_30/i0_0 ), .A3(\SB2_4_30/i1_7 ), .ZN(
        \SB2_4_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_30/Component_Function_4/N1  ( .A1(\SB2_4_30/i0[9] ), .A2(
        \SB2_4_30/i0_0 ), .A3(\SB2_4_30/i0[8] ), .ZN(
        \SB2_4_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_31/Component_Function_4/N1  ( .A1(\SB2_4_31/i0[9] ), .A2(
        \SB2_4_31/i0_0 ), .A3(\SB2_4_31/i0[8] ), .ZN(
        \SB2_4_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_2/N1  ( .A1(\SB3_0/i1_5 ), .A2(
        \SB3_0/i0[10] ), .A3(\SB3_0/i1[9] ), .ZN(
        \SB3_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_4/N2  ( .A1(\SB3_0/i3[0] ), .A2(
        \SB3_0/i0_0 ), .A3(\SB3_0/i1_7 ), .ZN(
        \SB3_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_0/Component_Function_4/N1  ( .A1(\SB3_0/i0[9] ), .A2(
        \SB3_0/i0_0 ), .A3(\SB3_0/i0[8] ), .ZN(
        \SB3_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_2/Component_Function_4/N2  ( .A1(\SB3_2/i3[0] ), .A2(
        \SB3_2/i0_0 ), .A3(\SB3_2/i1_7 ), .ZN(
        \SB3_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_3/Component_Function_4/N1  ( .A1(\SB3_3/i0[9] ), .A2(
        \SB3_3/i0_0 ), .A3(\SB3_3/i0[8] ), .ZN(
        \SB3_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_3/N2  ( .A1(\SB3_4/i0_0 ), .A2(
        \SB3_4/i0_3 ), .A3(\SB3_4/i0_4 ), .ZN(
        \SB3_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N4  ( .A1(\SB3_4/i1[9] ), .A2(
        \SB3_4/i1_5 ), .A3(\SB3_4/i0_4 ), .ZN(
        \SB3_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N2  ( .A1(\SB3_4/i3[0] ), .A2(
        \SB3_4/i0_0 ), .A3(\SB3_4/i1_7 ), .ZN(
        \SB3_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N1  ( .A1(\SB3_4/i0[9] ), .A2(
        \SB3_4/i0_0 ), .A3(\SB3_4/i0[8] ), .ZN(
        \SB3_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_3/N1  ( .A1(\SB3_5/i1[9] ), .A2(
        \SB3_5/i0_3 ), .A3(\SB3_5/i0[6] ), .ZN(
        \SB3_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_4/N2  ( .A1(\SB3_5/i3[0] ), .A2(
        \SB3_5/i0_0 ), .A3(\SB3_5/i1_7 ), .ZN(
        \SB3_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_5/Component_Function_4/N1  ( .A1(\SB3_5/i0[9] ), .A2(
        \SB3_5/i0_0 ), .A3(\SB3_5/i0[8] ), .ZN(
        \SB3_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_6/Component_Function_2/N1  ( .A1(\SB3_6/i1_5 ), .A2(
        \SB3_6/i0[10] ), .A3(\SB3_6/i1[9] ), .ZN(
        \SB3_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_6/Component_Function_3/N2  ( .A1(\SB3_6/i0_0 ), .A2(
        \SB3_6/i0_3 ), .A3(\SB3_6/i0_4 ), .ZN(
        \SB3_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_6/Component_Function_4/N1  ( .A1(\SB3_6/i0[9] ), .A2(
        \SB3_6/i0_0 ), .A3(\SB3_6/i0[8] ), .ZN(
        \SB3_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_2/N3  ( .A1(\SB3_8/i0_3 ), .A2(
        \SB3_8/i0[8] ), .A3(\SB3_8/i0[9] ), .ZN(
        \SB3_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_8/Component_Function_2/N1  ( .A1(\SB3_8/i1_5 ), .A2(
        \SB3_8/i0[10] ), .A3(\SB3_8/i1[9] ), .ZN(
        \SB3_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_3/N4  ( .A1(\SB3_8/i1_5 ), .A2(
        \SB3_8/i0[8] ), .A3(\SB3_8/i3[0] ), .ZN(
        \SB3_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_8/Component_Function_3/N1  ( .A1(\SB3_8/i1[9] ), .A2(
        \SB3_8/i0_3 ), .A3(\SB3_8/i0[6] ), .ZN(
        \SB3_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_4/N2  ( .A1(\SB3_8/i3[0] ), .A2(
        \SB3_8/i0_0 ), .A3(\SB3_8/i1_7 ), .ZN(
        \SB3_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_8/Component_Function_4/N1  ( .A1(\SB3_8/i0[9] ), .A2(
        \SB3_8/i0_0 ), .A3(\SB3_8/i0[8] ), .ZN(
        \SB3_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_3/N2  ( .A1(\SB3_9/i0_0 ), .A2(
        \SB3_9/i0_3 ), .A3(\SB3_9/i0_4 ), .ZN(
        \SB3_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_9/Component_Function_4/N4  ( .A1(\SB3_9/i1[9] ), .A2(
        \SB3_9/i1_5 ), .A3(\SB3_9/i0_4 ), .ZN(
        \SB3_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_9/Component_Function_4/N2  ( .A1(\SB3_9/i3[0] ), .A2(
        \SB3_9/i0_0 ), .A3(\SB3_9/i1_7 ), .ZN(
        \SB3_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_9/Component_Function_4/N1  ( .A1(\SB3_9/i0[9] ), .A2(
        \SB3_9/i0_0 ), .A3(\SB3_9/i0[8] ), .ZN(
        \SB3_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_2/N2  ( .A1(\SB3_10/i0_3 ), .A2(
        \SB3_10/i0[10] ), .A3(\SB3_10/i0[6] ), .ZN(
        \SB3_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_10/Component_Function_3/N1  ( .A1(\SB3_10/i1[9] ), .A2(
        \SB3_10/i0_3 ), .A3(\SB3_10/i0[6] ), .ZN(
        \SB3_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_4/N2  ( .A1(\SB3_10/i3[0] ), .A2(
        \SB3_10/i0_0 ), .A3(\SB3_10/i1_7 ), .ZN(
        \SB3_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_10/Component_Function_4/N1  ( .A1(\SB3_10/i0[9] ), .A2(
        \SB3_10/i0_0 ), .A3(\SB3_10/i0[8] ), .ZN(
        \SB3_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_3/N1  ( .A1(\SB3_12/i1[9] ), .A2(
        \RI1[5][119] ), .A3(\SB3_12/i0[6] ), .ZN(
        \SB3_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_4/N2  ( .A1(\SB3_12/i3[0] ), .A2(
        \SB3_12/i0_0 ), .A3(\SB3_12/i1_7 ), .ZN(
        \SB3_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_12/Component_Function_4/N1  ( .A1(\SB3_12/i0[9] ), .A2(
        \SB3_12/i0_0 ), .A3(\SB3_12/i0[8] ), .ZN(
        \SB3_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_4/N2  ( .A1(\SB3_13/i3[0] ), .A2(
        \SB3_13/i0_0 ), .A3(\SB3_13/i1_7 ), .ZN(
        \SB3_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_13/Component_Function_4/N1  ( .A1(\SB3_13/i0[9] ), .A2(
        \SB3_13/i0_0 ), .A3(\SB3_13/i0[8] ), .ZN(
        \SB3_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_2/N1  ( .A1(\SB3_14/i1_5 ), .A2(
        \SB3_14/i0[10] ), .A3(\SB3_14/i1[9] ), .ZN(
        \SB3_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_3/N3  ( .A1(\SB3_14/i1[9] ), .A2(
        \SB3_14/i1_7 ), .A3(\SB3_14/i0[10] ), .ZN(
        \SB3_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_14/Component_Function_4/N1  ( .A1(\SB3_14/i0[9] ), .A2(
        \SB3_14/i0_0 ), .A3(\SB3_14/i0[8] ), .ZN(
        \SB3_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_2/N2  ( .A1(\SB3_16/i0_3 ), .A2(
        \SB3_16/i0[10] ), .A3(\SB3_16/i0[6] ), .ZN(
        \SB3_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_16/Component_Function_2/N1  ( .A1(\SB3_16/i1_5 ), .A2(
        \SB3_16/i0[10] ), .A3(\SB3_16/i1[9] ), .ZN(
        \SB3_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_4/N2  ( .A1(\SB3_16/i3[0] ), .A2(
        \SB3_16/i0_0 ), .A3(\SB3_16/i1_7 ), .ZN(
        \SB3_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_16/Component_Function_4/N1  ( .A1(\SB3_16/i0[9] ), .A2(
        \SB3_16/i0_0 ), .A3(\SB3_16/i0[8] ), .ZN(
        \SB3_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_2/N2  ( .A1(\SB3_17/i0_3 ), .A2(
        \SB3_17/i0[10] ), .A3(\SB3_17/i0[6] ), .ZN(
        \SB3_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_17/Component_Function_3/N3  ( .A1(\SB3_17/i1[9] ), .A2(
        \SB3_17/i1_7 ), .A3(\SB3_17/i0[10] ), .ZN(
        \SB3_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_17/Component_Function_4/N4  ( .A1(\SB3_17/i1[9] ), .A2(
        \SB3_17/i1_5 ), .A3(\MC_ARK_ARC_1_4/buf_output[88] ), .ZN(
        \SB3_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_17/Component_Function_4/N2  ( .A1(\SB3_17/i3[0] ), .A2(
        \SB3_17/i0_0 ), .A3(\SB3_17/i1_7 ), .ZN(
        \SB3_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_18/Component_Function_4/N4  ( .A1(\SB3_18/i1[9] ), .A2(
        \SB3_18/i1_5 ), .A3(\SB3_18/i0_4 ), .ZN(
        \SB3_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_18/Component_Function_4/N3  ( .A1(\SB3_18/i0[9] ), .A2(
        \SB3_18/i0[10] ), .A3(\SB3_18/i0_3 ), .ZN(
        \SB3_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_18/Component_Function_4/N2  ( .A1(\SB3_18/i3[0] ), .A2(
        \SB3_18/i0_0 ), .A3(\SB3_18/i1_7 ), .ZN(
        \SB3_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_18/Component_Function_4/N1  ( .A1(\SB3_18/i0[9] ), .A2(
        \SB3_18/i0_0 ), .A3(\SB3_18/i0[8] ), .ZN(
        \SB3_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_4/N2  ( .A1(\SB3_19/i3[0] ), .A2(
        \SB3_19/i0_0 ), .A3(\SB3_19/i1_7 ), .ZN(
        \SB3_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_19/Component_Function_4/N1  ( .A1(\SB3_19/i0[9] ), .A2(
        \SB3_19/i0_0 ), .A3(\SB3_19/i0[8] ), .ZN(
        \SB3_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_2/N2  ( .A1(\SB3_20/i0_3 ), .A2(
        \SB3_20/i0[10] ), .A3(\SB3_20/i0[6] ), .ZN(
        \SB3_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_20/Component_Function_3/N1  ( .A1(\SB3_20/i1[9] ), .A2(
        \SB3_20/i0_3 ), .A3(\SB3_20/i0[6] ), .ZN(
        \SB3_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_4/N2  ( .A1(\SB3_20/i3[0] ), .A2(
        \SB3_20/i0_0 ), .A3(\SB3_20/i1_7 ), .ZN(
        \SB3_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_20/Component_Function_4/N1  ( .A1(\SB3_20/i0[9] ), .A2(
        \SB3_20/i0_0 ), .A3(\SB3_20/i0[8] ), .ZN(
        \SB3_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_4/N1  ( .A1(\SB3_21/i0[9] ), .A2(
        \SB3_21/i0_0 ), .A3(\SB3_21/i0[8] ), .ZN(
        \SB3_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_2/N2  ( .A1(\SB3_22/i0_3 ), .A2(
        \SB3_22/i0[10] ), .A3(\SB3_22/i0[6] ), .ZN(
        \SB3_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_22/Component_Function_4/N3  ( .A1(\SB3_22/i0[9] ), .A2(
        \SB3_22/i0[10] ), .A3(\SB3_22/i0_3 ), .ZN(
        \SB3_22/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_22/Component_Function_4/N2  ( .A1(\SB3_22/i3[0] ), .A2(
        \SB3_22/i0_0 ), .A3(\SB3_22/i1_7 ), .ZN(
        \SB3_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_22/Component_Function_4/N1  ( .A1(\SB3_22/i0[9] ), .A2(
        \SB3_22/i0_0 ), .A3(\SB3_22/i0[8] ), .ZN(
        \SB3_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_2/N2  ( .A1(\SB3_23/i0_3 ), .A2(
        \SB3_23/i0[10] ), .A3(\SB3_23/i0[6] ), .ZN(
        \SB3_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_23/Component_Function_3/N2  ( .A1(\SB3_23/i0_0 ), .A2(
        \RI1[5][53] ), .A3(\SB3_23/i0_4 ), .ZN(
        \SB3_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_23/Component_Function_4/N4  ( .A1(\SB3_23/i1[9] ), .A2(
        \SB3_23/i1_5 ), .A3(\SB3_23/i0_4 ), .ZN(
        \SB3_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_23/Component_Function_4/N2  ( .A1(\SB3_23/i3[0] ), .A2(
        \SB3_23/i0_0 ), .A3(\SB3_23/i1_7 ), .ZN(
        \SB3_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_24/Component_Function_4/N2  ( .A1(\SB3_24/i3[0] ), .A2(
        \SB3_24/i0_0 ), .A3(\SB3_24/i1_7 ), .ZN(
        \SB3_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_26/Component_Function_2/N1  ( .A1(\SB3_26/i1_5 ), .A2(
        \SB3_26/i0[10] ), .A3(\SB3_26/i1[9] ), .ZN(
        \SB3_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N2  ( .A1(\SB3_26/i3[0] ), .A2(
        \SB3_26/i0_0 ), .A3(\SB3_26/i1_7 ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N1  ( .A1(\SB3_26/i0[9] ), .A2(
        \SB3_26/i0_0 ), .A3(\SB3_26/i0[8] ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_4/N2  ( .A1(\SB3_27/i3[0] ), .A2(
        \SB3_27/i0_0 ), .A3(\SB3_27/i1_7 ), .ZN(
        \SB3_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_27/Component_Function_4/N1  ( .A1(\SB3_27/i0[9] ), .A2(
        \SB3_27/i0_0 ), .A3(\SB3_27/i0[8] ), .ZN(
        \SB3_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_2/N3  ( .A1(\SB3_28/i0_3 ), .A2(
        \SB3_28/i0[8] ), .A3(\SB3_28/i0[9] ), .ZN(
        \SB3_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_28/Component_Function_4/N2  ( .A1(\SB3_28/i3[0] ), .A2(
        \SB3_28/i0_0 ), .A3(\SB3_28/i1_7 ), .ZN(
        \SB3_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_28/Component_Function_4/N1  ( .A1(\SB3_28/i0[9] ), .A2(
        \SB3_28/i0_0 ), .A3(\SB3_28/i0[8] ), .ZN(
        \SB3_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_3/N2  ( .A1(\SB3_29/i0_0 ), .A2(
        \RI1[5][17] ), .A3(\SB3_29/i0_4 ), .ZN(
        \SB3_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_29/Component_Function_4/N2  ( .A1(\SB3_29/i3[0] ), .A2(
        \SB3_29/i0_0 ), .A3(\SB3_29/i1_7 ), .ZN(
        \SB3_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_30/Component_Function_4/N2  ( .A1(\SB3_30/i3[0] ), .A2(
        \SB3_30/i0_0 ), .A3(\SB3_30/i1_7 ), .ZN(
        \SB3_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_31/Component_Function_4/N2  ( .A1(\SB3_31/i3[0] ), .A2(
        \SB3_31/i0_0 ), .A3(\SB3_31/i1_7 ), .ZN(
        \SB3_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_0/Component_Function_2/N3  ( .A1(\SB4_0/i0_3 ), .A2(
        \SB4_0/i0[8] ), .A3(\SB4_0/i0[9] ), .ZN(
        \SB4_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_0/Component_Function_4/N1  ( .A1(\SB4_0/i0[9] ), .A2(
        \SB4_0/i0_0 ), .A3(\SB4_0/i0[8] ), .ZN(
        \SB4_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_2/Component_Function_2/N2  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i0[10] ), .A3(\SB4_2/i0[6] ), .ZN(
        \SB4_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_2/Component_Function_2/N1  ( .A1(\SB4_2/i1_5 ), .A2(
        \SB4_2/i0[10] ), .A3(\SB4_2/i1[9] ), .ZN(
        \SB4_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_2/Component_Function_3/N4  ( .A1(\SB4_2/i1_5 ), .A2(
        \SB4_2/i0[8] ), .A3(\SB4_2/i3[0] ), .ZN(
        \SB4_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_2/Component_Function_4/N4  ( .A1(\SB4_2/i1[9] ), .A2(
        \SB4_2/i1_5 ), .A3(\SB4_2/i0_4 ), .ZN(
        \SB4_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_3/Component_Function_2/N3  ( .A1(\SB4_3/i0_3 ), .A2(
        \SB4_3/i0[8] ), .A3(\SB4_3/i0[9] ), .ZN(
        \SB4_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_3/Component_Function_3/N4  ( .A1(\SB4_3/i1_5 ), .A2(
        \SB4_3/i0[8] ), .A3(\SB4_3/i3[0] ), .ZN(
        \SB4_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_4/Component_Function_3/N2  ( .A1(\SB4_4/i0_0 ), .A2(
        \SB4_4/i0_3 ), .A3(\SB4_4/i0_4 ), .ZN(
        \SB4_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_4/Component_Function_4/N4  ( .A1(\SB4_4/i1[9] ), .A2(
        \SB4_4/i1_5 ), .A3(\SB4_4/i0_4 ), .ZN(
        \SB4_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_5/Component_Function_3/N4  ( .A1(\SB4_5/i1_5 ), .A2(
        \SB4_5/i0[8] ), .A3(\SB4_5/i3[0] ), .ZN(
        \SB4_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_5/Component_Function_4/N1  ( .A1(\SB4_5/i0[9] ), .A2(
        \SB4_5/i0_0 ), .A3(\SB4_5/i0[8] ), .ZN(
        \SB4_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_7/Component_Function_2/N3  ( .A1(\SB4_7/i0_3 ), .A2(n3965), 
        .A3(\SB4_7/i0[9] ), .ZN(\SB4_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_7/Component_Function_3/N4  ( .A1(\SB4_7/i1_5 ), .A2(n3965), 
        .A3(\SB4_7/i3[0] ), .ZN(\SB4_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_7/Component_Function_3/N1  ( .A1(\SB4_7/i1[9] ), .A2(
        \SB4_7/i0_3 ), .A3(\SB4_7/i0[6] ), .ZN(
        \SB4_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB4_8/Component_Function_2/N3  ( .A1(\SB4_8/i0_3 ), .A2(
        \SB4_8/i0[8] ), .A3(\SB4_8/i0[9] ), .ZN(
        \SB4_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_8/Component_Function_3/N4  ( .A1(\SB4_8/i1_5 ), .A2(
        \SB4_8/i0[8] ), .A3(\SB4_8/i3[0] ), .ZN(
        \SB4_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_8/Component_Function_3/N1  ( .A1(n3996), .A2(\SB4_8/i0_3 ), 
        .A3(\SB4_8/i0[6] ), .ZN(\SB4_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB4_8/Component_Function_4/N3  ( .A1(\SB4_8/i0[9] ), .A2(
        \SB4_8/i0[10] ), .A3(\SB4_8/i0_3 ), .ZN(
        \SB4_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_9/Component_Function_2/N1  ( .A1(\SB4_9/i1_5 ), .A2(
        \SB4_9/i0[10] ), .A3(\SB4_9/i1[9] ), .ZN(
        \SB4_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_9/Component_Function_4/N4  ( .A1(\SB4_9/i1[9] ), .A2(
        \SB4_9/i1_5 ), .A3(\SB3_10/buf_output[4] ), .ZN(
        \SB4_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_12/Component_Function_2/N1  ( .A1(\SB4_12/i1_5 ), .A2(
        \SB4_12/i0[10] ), .A3(\SB4_12/i1[9] ), .ZN(
        \SB4_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_13/Component_Function_2/N3  ( .A1(\SB4_13/i0_3 ), .A2(n1498), 
        .A3(\SB4_13/i0[9] ), .ZN(\SB4_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_13/Component_Function_2/N2  ( .A1(\SB4_13/i0_3 ), .A2(
        \SB3_15/buf_output[3] ), .A3(\SB4_13/i0[6] ), .ZN(
        \SB4_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_14/Component_Function_2/N3  ( .A1(\SB4_14/i0_3 ), .A2(
        \SB4_14/i0[8] ), .A3(\SB4_14/i0[9] ), .ZN(
        \SB4_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_14/Component_Function_3/N2  ( .A1(\SB4_14/i0_0 ), .A2(
        \SB4_14/i0_3 ), .A3(\SB4_14/i0_4 ), .ZN(
        \SB4_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_14/Component_Function_3/N1  ( .A1(\SB4_14/i1[9] ), .A2(
        \SB4_14/i0_3 ), .A3(\SB4_14/i0[6] ), .ZN(
        \SB4_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB4_15/Component_Function_2/N1  ( .A1(\SB4_15/i1_5 ), .A2(
        \SB3_17/buf_output[3] ), .A3(\SB4_15/i1[9] ), .ZN(
        \SB4_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_15/Component_Function_3/N2  ( .A1(\SB4_15/i0_0 ), .A2(
        \SB4_15/i0_3 ), .A3(\SB4_15/i0_4 ), .ZN(
        \SB4_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_15/Component_Function_4/N1  ( .A1(\SB4_15/i0[9] ), .A2(
        \SB4_15/i0_0 ), .A3(n1497), .ZN(
        \SB4_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_16/Component_Function_2/N3  ( .A1(\SB4_16/i0_3 ), .A2(
        \SB4_16/i0[8] ), .A3(\SB4_16/i0[9] ), .ZN(
        \SB4_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_17/Component_Function_3/N2  ( .A1(\SB4_17/i0_0 ), .A2(
        \SB4_17/i0_3 ), .A3(\SB4_17/i0_4 ), .ZN(
        \SB4_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_17/Component_Function_4/N1  ( .A1(\SB4_17/i0[9] ), .A2(
        \SB4_17/i0_0 ), .A3(n1493), .ZN(
        \SB4_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_18/Component_Function_2/N3  ( .A1(\SB4_18/i0_3 ), .A2(
        \SB4_18/i0[8] ), .A3(\SB4_18/i0[9] ), .ZN(
        \SB4_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_18/Component_Function_2/N1  ( .A1(\SB4_18/i1_5 ), .A2(
        \SB4_18/i0[10] ), .A3(n1496), .ZN(
        \SB4_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_18/Component_Function_4/N4  ( .A1(n1496), .A2(\SB4_18/i1_5 ), 
        .A3(\SB4_18/i0_4 ), .ZN(\SB4_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_19/Component_Function_3/N1  ( .A1(\SB4_19/i1[9] ), .A2(
        \SB4_19/i0_3 ), .A3(\SB4_19/i0[6] ), .ZN(
        \SB4_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB4_19/Component_Function_4/N4  ( .A1(\SB4_19/i1[9] ), .A2(n6273), 
        .A3(\SB4_19/i0_4 ), .ZN(\SB4_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_20/Component_Function_3/N4  ( .A1(\SB4_20/i1_5 ), .A2(
        \SB4_20/i0[8] ), .A3(\SB4_20/i3[0] ), .ZN(
        \SB4_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_21/Component_Function_2/N1  ( .A1(\SB4_21/i1_5 ), .A2(
        \SB4_21/i0[10] ), .A3(n3998), .ZN(
        \SB4_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_21/Component_Function_3/N2  ( .A1(\SB3_24/buf_output[2] ), 
        .A2(\SB4_21/i0_3 ), .A3(\SB4_21/i0_4 ), .ZN(
        \SB4_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_22/Component_Function_2/N3  ( .A1(\SB4_22/i0_3 ), .A2(
        \SB4_22/i0[8] ), .A3(\SB4_22/i0[9] ), .ZN(
        \SB4_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_22/Component_Function_4/N4  ( .A1(\SB4_22/i1[9] ), .A2(
        \SB4_22/i1_5 ), .A3(\SB4_22/i0_4 ), .ZN(
        \SB4_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_23/Component_Function_3/N4  ( .A1(\SB4_23/i1_5 ), .A2(n3974), 
        .A3(\SB4_23/i3[0] ), .ZN(\SB4_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_24/Component_Function_4/N1  ( .A1(\SB4_24/i0[9] ), .A2(
        \SB4_24/i0_0 ), .A3(n1494), .ZN(
        \SB4_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_25/Component_Function_2/N4  ( .A1(\SB4_25/i1_5 ), .A2(
        \SB4_25/i0_0 ), .A3(\SB4_25/i0_4 ), .ZN(
        \SB4_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_3/N4  ( .A1(\SB4_25/i1_5 ), .A2(
        \SB4_25/i0[8] ), .A3(n5438), .ZN(
        \SB4_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_4/N4  ( .A1(\SB4_25/i1[9] ), .A2(
        \SB4_25/i1_5 ), .A3(\SB4_25/i0_4 ), .ZN(
        \SB4_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_4/N2  ( .A1(n5438), .A2(\SB4_25/i0_0 ), 
        .A3(\SB4_25/i1_7 ), .ZN(\SB4_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_26/Component_Function_2/N1  ( .A1(\SB4_26/i1_5 ), .A2(
        \SB4_26/i0[10] ), .A3(n573), .ZN(
        \SB4_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_26/Component_Function_3/N4  ( .A1(\SB4_26/i1_5 ), .A2(n3989), 
        .A3(\SB4_26/i3[0] ), .ZN(\SB4_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_27/Component_Function_2/N1  ( .A1(\SB4_27/i1_5 ), .A2(
        \SB4_27/i0[10] ), .A3(\SB4_27/i1[9] ), .ZN(
        \SB4_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_3/N2  ( .A1(\SB4_27/i0_0 ), .A2(
        \SB4_27/i0_3 ), .A3(\SB4_27/i0_4 ), .ZN(
        \SB4_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_29/Component_Function_4/N1  ( .A1(\SB4_29/i0[9] ), .A2(
        \SB4_29/i0_0 ), .A3(\SB4_29/i0[8] ), .ZN(
        \SB4_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_30/Component_Function_3/N4  ( .A1(\SB4_30/i1_5 ), .A2(
        \SB4_30/i0[8] ), .A3(\SB4_30/i3[0] ), .ZN(
        \SB4_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_30/Component_Function_4/N4  ( .A1(n3973), .A2(\SB4_30/i1_5 ), 
        .A3(\SB4_30/i0_4 ), .ZN(\SB4_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_30/Component_Function_4/N2  ( .A1(\SB4_30/i3[0] ), .A2(n5427), 
        .A3(\SB4_30/i1_7 ), .ZN(\SB4_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_31/Component_Function_4/N4  ( .A1(\SB4_31/i1[9] ), .A2(
        \SB4_31/i1_5 ), .A3(\SB4_31/i0_4 ), .ZN(
        \SB4_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_0/N4  ( .A1(\SB1_0_0/i0[7] ), .A2(
        \SB1_0_0/i0_3 ), .A3(\SB1_0_0/i0_0 ), .ZN(
        \SB1_0_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_1/N4  ( .A1(\SB1_0_0/i1_7 ), .A2(
        \SB1_0_0/i0[8] ), .A3(\SB1_0_0/i0_4 ), .ZN(
        \SB1_0_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_1/N3  ( .A1(\SB1_0_0/i1_5 ), .A2(
        \SB1_0_0/i0[6] ), .A3(\SB1_0_0/i0[9] ), .ZN(
        \SB1_0_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_0/Component_Function_1/N2  ( .A1(\SB1_0_0/i0_3 ), .A2(
        \SB1_0_0/i1_7 ), .A3(\SB1_0_0/i0[8] ), .ZN(
        \SB1_0_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_0/Component_Function_5/N3  ( .A1(\SB1_0_0/i1[9] ), .A2(n380), 
        .A3(\SB1_0_0/i0_3 ), .ZN(\SB1_0_0/Component_Function_5/NAND4_in[2] )
         );
  NAND3_X1 \SB1_0_1/Component_Function_0/N3  ( .A1(\SB1_0_1/i0[10] ), .A2(
        \SB1_0_1/i0_4 ), .A3(\SB1_0_1/i0_3 ), .ZN(
        \SB1_0_1/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_1/Component_Function_0/N1  ( .A1(\SB1_0_1/i0[10] ), .A2(
        \SB1_0_1/i0[9] ), .ZN(\SB1_0_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_1/N2  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i1_7 ), .A3(\SB1_0_1/i0[8] ), .ZN(
        \SB1_0_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_1/Component_Function_1/N1  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i1[9] ), .ZN(\SB1_0_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_5/N4  ( .A1(\SB1_0_1/i0[9] ), .A2(n251), 
        .A3(n378), .ZN(\SB1_0_1/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_2/Component_Function_0/N1  ( .A1(\SB1_0_2/i0[10] ), .A2(
        \SB1_0_2/i0[9] ), .ZN(\SB1_0_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_2/Component_Function_1/N3  ( .A1(\SB1_0_2/i1_5 ), .A2(
        \SB1_0_2/i0[6] ), .A3(\SB1_0_2/i0[9] ), .ZN(
        \SB1_0_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_3/Component_Function_0/N2  ( .A1(\SB1_0_3/i0[8] ), .A2(
        \SB1_0_3/i0[7] ), .A3(\SB1_0_3/i0[6] ), .ZN(
        \SB1_0_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_3/Component_Function_0/N1  ( .A1(\SB1_0_3/i0[10] ), .A2(
        \SB1_0_3/i0[9] ), .ZN(\SB1_0_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_1/N3  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0[6] ), .A3(\SB1_0_3/i0[9] ), .ZN(
        \SB1_0_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_3/Component_Function_1/N2  ( .A1(\SB1_0_3/i0_3 ), .A2(
        \SB1_0_3/i1_7 ), .A3(\SB1_0_3/i0[8] ), .ZN(
        \SB1_0_3/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_4/Component_Function_0/N4  ( .A1(\SB1_0_4/i0[7] ), .A2(
        \SB1_0_4/i0_3 ), .A3(\SB1_0_4/i0_0 ), .ZN(
        \SB1_0_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_0/N2  ( .A1(\SB1_0_4/i0[8] ), .A2(
        \SB1_0_4/i0[7] ), .A3(\SB1_0_4/i0[6] ), .ZN(
        \SB1_0_4/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_4/Component_Function_1/N3  ( .A1(\SB1_0_4/i1_5 ), .A2(
        \SB1_0_4/i0[6] ), .A3(\SB1_0_4/i0[9] ), .ZN(
        \SB1_0_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_5/Component_Function_1/N2  ( .A1(\SB1_0_5/i0_3 ), .A2(
        \SB1_0_5/i1_7 ), .A3(\SB1_0_5/i0[8] ), .ZN(
        \SB1_0_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_5/Component_Function_5/N4  ( .A1(n305), .A2(n247), .A3(n370), 
        .ZN(\SB1_0_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_0/N2  ( .A1(\SB1_0_6/i0[8] ), .A2(
        \SB1_0_6/i0[7] ), .A3(\SB1_0_6/i0[6] ), .ZN(
        \SB1_0_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_6/Component_Function_0/N1  ( .A1(\SB1_0_6/i0[10] ), .A2(
        \SB1_0_6/i0[9] ), .ZN(\SB1_0_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_1/N3  ( .A1(\SB1_0_6/i1_5 ), .A2(
        \SB1_0_6/i0[6] ), .A3(\SB1_0_6/i0[9] ), .ZN(
        \SB1_0_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_6/Component_Function_1/N2  ( .A1(\SB1_0_6/i0_3 ), .A2(
        \SB1_0_6/i1_7 ), .A3(\SB1_0_6/i0[8] ), .ZN(
        \SB1_0_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_6/Component_Function_1/N1  ( .A1(\SB1_0_6/i0_3 ), .A2(
        \SB1_0_6/i1[9] ), .ZN(\SB1_0_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_0/N4  ( .A1(\SB1_0_7/i0[7] ), .A2(
        \SB1_0_7/i0_3 ), .A3(\SB1_0_7/i0_0 ), .ZN(
        \SB1_0_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_0/N3  ( .A1(\SB1_0_7/i0[10] ), .A2(
        \SB1_0_7/i0_4 ), .A3(\SB1_0_7/i0_3 ), .ZN(
        \SB1_0_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_0/N2  ( .A1(\SB1_0_7/i0[8] ), .A2(
        \SB1_0_7/i0[7] ), .A3(\SB1_0_7/i0[6] ), .ZN(
        \SB1_0_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_7/Component_Function_0/N1  ( .A1(\SB1_0_7/i0[10] ), .A2(
        \SB1_0_7/i0[9] ), .ZN(\SB1_0_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_1/N4  ( .A1(\SB1_0_7/i1_7 ), .A2(
        \SB1_0_7/i0[8] ), .A3(\SB1_0_7/i0_4 ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_1/N3  ( .A1(\SB1_0_7/i1_5 ), .A2(
        \SB1_0_7/i0[6] ), .A3(\SB1_0_7/i0[9] ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_1/N2  ( .A1(\SB1_0_7/i0_3 ), .A2(
        \SB1_0_7/i1_7 ), .A3(\SB1_0_7/i0[8] ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_8/Component_Function_0/N3  ( .A1(\SB1_0_8/i0[10] ), .A2(
        \SB1_0_8/i0_4 ), .A3(\SB1_0_8/i0_3 ), .ZN(
        \SB1_0_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_8/Component_Function_0/N2  ( .A1(\SB1_0_8/i0[8] ), .A2(
        \SB1_0_8/i0[7] ), .A3(\SB1_0_8/i0[6] ), .ZN(
        \SB1_0_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_8/Component_Function_0/N1  ( .A1(\SB1_0_8/i0[10] ), .A2(
        \SB1_0_8/i0[9] ), .ZN(\SB1_0_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_1/N3  ( .A1(\SB1_0_8/i1_5 ), .A2(
        \SB1_0_8/i0[6] ), .A3(\SB1_0_8/i0[9] ), .ZN(
        \SB1_0_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_8/Component_Function_1/N2  ( .A1(\SB1_0_8/i0_3 ), .A2(
        \SB1_0_8/i1_7 ), .A3(\SB1_0_8/i0[8] ), .ZN(
        \SB1_0_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_8/Component_Function_5/N1  ( .A1(\SB1_0_8/i0_0 ), .A2(
        \SB1_0_8/i3[0] ), .ZN(\SB1_0_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_0/N3  ( .A1(\SB1_0_9/i0[10] ), .A2(
        \SB1_0_9/i0_4 ), .A3(\SB1_0_9/i0_3 ), .ZN(
        \SB1_0_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_9/Component_Function_0/N2  ( .A1(\SB1_0_9/i0[8] ), .A2(
        \SB1_0_9/i0[7] ), .A3(\SB1_0_9/i0[6] ), .ZN(
        \SB1_0_9/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_9/Component_Function_1/N4  ( .A1(\SB1_0_9/i1_7 ), .A2(
        \SB1_0_9/i0[8] ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_1/N2  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i1_7 ), .A3(\SB1_0_9/i0[8] ), .ZN(
        \SB1_0_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_9/Component_Function_1/N1  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i1[9] ), .ZN(\SB1_0_9/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_9/Component_Function_5/N1  ( .A1(\SB1_0_9/i0_0 ), .A2(
        \SB1_0_9/i3[0] ), .ZN(\SB1_0_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_0/N3  ( .A1(\SB1_0_10/i0[10] ), .A2(
        \SB1_0_10/i0_4 ), .A3(\SB1_0_10/i0_3 ), .ZN(
        \SB1_0_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_10/Component_Function_1/N2  ( .A1(\SB1_0_10/i0_3 ), .A2(
        \SB1_0_10/i1_7 ), .A3(\SB1_0_10/i0[8] ), .ZN(
        \SB1_0_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_10/Component_Function_1/N1  ( .A1(\SB1_0_10/i0_3 ), .A2(
        \SB1_0_10/i1[9] ), .ZN(\SB1_0_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_5/N2  ( .A1(\SB1_0_10/i0_0 ), .A2(
        \SB1_0_10/i0[6] ), .A3(\SB1_0_10/i0[10] ), .ZN(
        \SB1_0_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_11/Component_Function_0/N2  ( .A1(\SB1_0_11/i0[8] ), .A2(
        \SB1_0_11/i0[7] ), .A3(\SB1_0_11/i0[6] ), .ZN(
        \SB1_0_11/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_11/Component_Function_1/N4  ( .A1(\SB1_0_11/i1_7 ), .A2(
        \SB1_0_11/i0[8] ), .A3(\SB1_0_11/i0_4 ), .ZN(
        \SB1_0_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_11/Component_Function_1/N3  ( .A1(\SB1_0_11/i1_5 ), .A2(
        \SB1_0_11/i0[6] ), .A3(n293), .ZN(
        \SB1_0_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_1/N2  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i1_7 ), .A3(\SB1_0_11/i0[8] ), .ZN(
        \SB1_0_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_11/Component_Function_1/N1  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i1[9] ), .ZN(\SB1_0_11/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_11/Component_Function_5/N1  ( .A1(\SB1_0_11/i0_0 ), .A2(
        \SB1_0_11/i3[0] ), .ZN(\SB1_0_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_0/N3  ( .A1(\SB1_0_12/i0[10] ), .A2(
        \SB1_0_12/i0_4 ), .A3(\SB1_0_12/i0_3 ), .ZN(
        \SB1_0_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_12/Component_Function_0/N2  ( .A1(\SB1_0_12/i0[8] ), .A2(
        \SB1_0_12/i0[7] ), .A3(\SB1_0_12/i0[6] ), .ZN(
        \SB1_0_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_12/Component_Function_0/N1  ( .A1(\SB1_0_12/i0[10] ), .A2(
        \SB1_0_12/i0[9] ), .ZN(\SB1_0_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_1/N4  ( .A1(\SB1_0_12/i1_7 ), .A2(
        \SB1_0_12/i0[8] ), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_1/N3  ( .A1(\SB1_0_12/i1_5 ), .A2(
        \SB1_0_12/i0[6] ), .A3(\SB1_0_12/i0[9] ), .ZN(
        \SB1_0_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_12/Component_Function_1/N2  ( .A1(\SB1_0_12/i0_3 ), .A2(
        \SB1_0_12/i1_7 ), .A3(\SB1_0_12/i0[8] ), .ZN(
        \SB1_0_12/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_13/Component_Function_0/N3  ( .A1(\SB1_0_13/i0[10] ), .A2(
        \SB1_0_13/i0_4 ), .A3(\SB1_0_13/i0_3 ), .ZN(
        \SB1_0_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_13/Component_Function_0/N2  ( .A1(n5428), .A2(
        \SB1_0_13/i0[7] ), .A3(\SB1_0_13/i0[6] ), .ZN(
        \SB1_0_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_13/Component_Function_0/N1  ( .A1(\SB1_0_13/i0[10] ), .A2(
        \SB1_0_13/i0[9] ), .ZN(\SB1_0_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_5/N2  ( .A1(\SB1_0_13/i0_0 ), .A2(
        \SB1_0_13/i0[6] ), .A3(\SB1_0_13/i0[10] ), .ZN(
        \SB1_0_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_14/Component_Function_0/N4  ( .A1(\SB1_0_14/i0[7] ), .A2(
        \SB1_0_14/i0_3 ), .A3(\SB1_0_14/i0_0 ), .ZN(
        \SB1_0_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_14/Component_Function_1/N3  ( .A1(\SB1_0_14/i1_5 ), .A2(
        \SB1_0_14/i0[6] ), .A3(\SB1_0_14/i0[9] ), .ZN(
        \SB1_0_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_14/Component_Function_1/N2  ( .A1(\SB1_0_14/i0_3 ), .A2(
        \SB1_0_14/i1_7 ), .A3(\SB1_0_14/i0[8] ), .ZN(
        \SB1_0_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_15/Component_Function_0/N3  ( .A1(\SB1_0_15/i0[10] ), .A2(
        \SB1_0_15/i0_4 ), .A3(\SB1_0_15/i0_3 ), .ZN(
        \SB1_0_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_16/Component_Function_0/N3  ( .A1(\SB1_0_16/i0[10] ), .A2(
        \SB1_0_16/i0_4 ), .A3(\SB1_0_16/i0_3 ), .ZN(
        \SB1_0_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_16/Component_Function_0/N2  ( .A1(\SB1_0_16/i0[8] ), .A2(
        \SB1_0_16/i0[7] ), .A3(\SB1_0_16/i0[6] ), .ZN(
        \SB1_0_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_16/Component_Function_0/N1  ( .A1(\SB1_0_16/i0[10] ), .A2(
        \SB1_0_16/i0[9] ), .ZN(\SB1_0_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_1/N4  ( .A1(\SB1_0_16/i1_7 ), .A2(
        \SB1_0_16/i0[8] ), .A3(\SB1_0_16/i0_4 ), .ZN(
        \SB1_0_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_16/Component_Function_5/N2  ( .A1(\SB1_0_16/i0_0 ), .A2(
        \SB1_0_16/i0[6] ), .A3(\SB1_0_16/i0[10] ), .ZN(
        \SB1_0_16/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_17/Component_Function_0/N4  ( .A1(\SB1_0_17/i0[7] ), .A2(
        \SB1_0_17/i0_3 ), .A3(\SB1_0_17/i0_0 ), .ZN(
        \SB1_0_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_0/N3  ( .A1(\SB1_0_17/i0[10] ), .A2(
        \SB1_0_17/i0_4 ), .A3(\SB1_0_17/i0_3 ), .ZN(
        \SB1_0_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_17/Component_Function_0/N2  ( .A1(\SB1_0_17/i0[8] ), .A2(
        \SB1_0_17/i0[7] ), .A3(\SB1_0_17/i0[6] ), .ZN(
        \SB1_0_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_17/Component_Function_0/N1  ( .A1(\SB1_0_17/i0[10] ), .A2(
        \SB1_0_17/i0[9] ), .ZN(\SB1_0_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_17/Component_Function_1/N4  ( .A1(\SB1_0_17/i1_7 ), .A2(
        \SB1_0_17/i0[8] ), .A3(\SB1_0_17/i0_4 ), .ZN(
        \SB1_0_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_1/N3  ( .A1(\SB1_0_17/i1_5 ), .A2(
        \SB1_0_17/i0[6] ), .A3(\SB1_0_17/i0[9] ), .ZN(
        \SB1_0_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_17/Component_Function_1/N2  ( .A1(\SB1_0_17/i0_3 ), .A2(
        \SB1_0_17/i1_7 ), .A3(\SB1_0_17/i0[8] ), .ZN(
        \SB1_0_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_17/Component_Function_1/N1  ( .A1(\SB1_0_17/i0_3 ), .A2(
        \SB1_0_17/i1[9] ), .ZN(\SB1_0_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_0/N3  ( .A1(\SB1_0_18/i0[10] ), .A2(
        \SB1_0_18/i0_4 ), .A3(\SB1_0_18/i0_3 ), .ZN(
        \SB1_0_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_19/Component_Function_0/N3  ( .A1(\SB1_0_19/i0[10] ), .A2(
        \SB1_0_19/i0_4 ), .A3(\SB1_0_19/i0_3 ), .ZN(
        \SB1_0_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_19/Component_Function_1/N3  ( .A1(\SB1_0_19/i1_5 ), .A2(
        \SB1_0_19/i0[6] ), .A3(\SB1_0_19/i0[9] ), .ZN(
        \SB1_0_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_20/Component_Function_0/N3  ( .A1(\SB1_0_20/i0[10] ), .A2(
        \SB1_0_20/i0_4 ), .A3(\SB1_0_20/i0_3 ), .ZN(
        \SB1_0_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_20/Component_Function_1/N3  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0[6] ), .A3(\SB1_0_20/i0[9] ), .ZN(
        \SB1_0_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_20/Component_Function_1/N2  ( .A1(\SB1_0_20/i0_3 ), .A2(
        \SB1_0_20/i1_7 ), .A3(\SB1_0_20/i0[8] ), .ZN(
        \SB1_0_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_21/Component_Function_0/N3  ( .A1(\SB1_0_21/i0[10] ), .A2(
        \SB1_0_21/i0_4 ), .A3(\SB1_0_21/i0_3 ), .ZN(
        \SB1_0_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_21/Component_Function_0/N2  ( .A1(\SB1_0_21/i0[8] ), .A2(
        \SB1_0_21/i0[7] ), .A3(\SB1_0_21/i0[6] ), .ZN(
        \SB1_0_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_21/Component_Function_1/N2  ( .A1(\SB1_0_21/i0_3 ), .A2(
        \SB1_0_21/i1_7 ), .A3(\SB1_0_21/i0[8] ), .ZN(
        \SB1_0_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_21/Component_Function_1/N1  ( .A1(\SB1_0_21/i0_3 ), .A2(
        \SB1_0_21/i1[9] ), .ZN(\SB1_0_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_0/N2  ( .A1(\SB1_0_22/i0[8] ), .A2(
        \SB1_0_22/i0[7] ), .A3(\SB1_0_22/i0[6] ), .ZN(
        \SB1_0_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_22/Component_Function_0/N1  ( .A1(\SB1_0_22/i0[10] ), .A2(
        \SB1_0_22/i0[9] ), .ZN(\SB1_0_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_1/N4  ( .A1(\SB1_0_22/i1_7 ), .A2(
        \SB1_0_22/i0[8] ), .A3(\SB1_0_22/i0_4 ), .ZN(
        \SB1_0_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_22/Component_Function_1/N3  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0[6] ), .A3(\SB1_0_22/i0[9] ), .ZN(
        \SB1_0_22/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_22/Component_Function_1/N1  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i1[9] ), .ZN(\SB1_0_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_0/N4  ( .A1(\SB1_0_23/i0[7] ), .A2(
        \SB1_0_23/i0_3 ), .A3(\SB1_0_23/i0_0 ), .ZN(
        \SB1_0_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_23/Component_Function_0/N2  ( .A1(\SB1_0_23/i0[8] ), .A2(
        \SB1_0_23/i0[7] ), .A3(\SB1_0_23/i0[6] ), .ZN(
        \SB1_0_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_23/Component_Function_0/N1  ( .A1(\SB1_0_23/i0[10] ), .A2(
        \SB1_0_23/i0[9] ), .ZN(\SB1_0_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_1/N2  ( .A1(\SB1_0_23/i0_3 ), .A2(
        \SB1_0_23/i1_7 ), .A3(\SB1_0_23/i0[8] ), .ZN(
        \SB1_0_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_23/Component_Function_5/N2  ( .A1(\SB1_0_23/i0_0 ), .A2(
        \SB1_0_23/i0[6] ), .A3(\SB1_0_23/i0[10] ), .ZN(
        \SB1_0_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_24/Component_Function_1/N2  ( .A1(\SB1_0_24/i0_3 ), .A2(
        \SB1_0_24/i1_7 ), .A3(\SB1_0_24/i0[8] ), .ZN(
        \SB1_0_24/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_25/Component_Function_0/N2  ( .A1(\SB1_0_25/i0[8] ), .A2(
        \SB1_0_25/i0[7] ), .A3(\SB1_0_25/i0[6] ), .ZN(
        \SB1_0_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_25/Component_Function_0/N1  ( .A1(\SB1_0_25/i0[10] ), .A2(
        \SB1_0_25/i0[9] ), .ZN(\SB1_0_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_1/N4  ( .A1(\SB1_0_25/i1_7 ), .A2(
        \SB1_0_25/i0[8] ), .A3(n330), .ZN(
        \SB1_0_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_0/N4  ( .A1(\SB1_0_26/i0[7] ), .A2(
        \SB1_0_26/i0_3 ), .A3(\SB1_0_26/i0_0 ), .ZN(
        \SB1_0_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_0/N3  ( .A1(\SB1_0_26/i0[10] ), .A2(
        \SB1_0_26/i0_4 ), .A3(\SB1_0_26/i0_3 ), .ZN(
        \SB1_0_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_26/Component_Function_0/N2  ( .A1(\SB1_0_26/i0[8] ), .A2(
        \SB1_0_26/i0[7] ), .A3(\SB1_0_26/i0[6] ), .ZN(
        \SB1_0_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_26/Component_Function_0/N1  ( .A1(\SB1_0_26/i0[10] ), .A2(
        \SB1_0_26/i0[9] ), .ZN(\SB1_0_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_1/N4  ( .A1(\SB1_0_26/i1_7 ), .A2(
        \SB1_0_26/i0[8] ), .A3(\SB1_0_26/i0_4 ), .ZN(
        \SB1_0_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_1/N2  ( .A1(\SB1_0_26/i0_3 ), .A2(
        \SB1_0_26/i1_7 ), .A3(\SB1_0_26/i0[8] ), .ZN(
        \SB1_0_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_26/Component_Function_1/N1  ( .A1(\SB1_0_26/i0_3 ), .A2(
        \SB1_0_26/i1[9] ), .ZN(\SB1_0_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_5/N2  ( .A1(\SB1_0_26/i0_0 ), .A2(
        \SB1_0_26/i0[6] ), .A3(\SB1_0_26/i0[10] ), .ZN(
        \SB1_0_26/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_27/Component_Function_0/N4  ( .A1(\SB1_0_27/i0[7] ), .A2(
        \SB1_0_27/i0_3 ), .A3(\SB1_0_27/i0_0 ), .ZN(
        \SB1_0_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_0/N3  ( .A1(\SB1_0_27/i0[10] ), .A2(
        \SB1_0_27/i0_4 ), .A3(\SB1_0_27/i0_3 ), .ZN(
        \SB1_0_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_27/Component_Function_0/N2  ( .A1(\SB1_0_27/i0[8] ), .A2(
        \SB1_0_27/i0[7] ), .A3(\SB1_0_27/i0[6] ), .ZN(
        \SB1_0_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_27/Component_Function_0/N1  ( .A1(\SB1_0_27/i0[10] ), .A2(
        \SB1_0_27/i0[9] ), .ZN(\SB1_0_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_1/N3  ( .A1(\SB1_0_27/i1_5 ), .A2(n225), .A3(n261), .ZN(\SB1_0_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_27/Component_Function_1/N2  ( .A1(\SB1_0_27/i0_3 ), .A2(
        \SB1_0_27/i1_7 ), .A3(\SB1_0_27/i0[8] ), .ZN(
        \SB1_0_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_27/Component_Function_1/N1  ( .A1(\SB1_0_27/i0_3 ), .A2(
        \SB1_0_27/i1[9] ), .ZN(\SB1_0_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_5/N4  ( .A1(\SB1_0_27/i0[9] ), .A2(
        \SB1_0_27/i0[6] ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_27/Component_Function_5/N1  ( .A1(\SB1_0_27/i0_0 ), .A2(
        \SB1_0_27/i3[0] ), .ZN(\SB1_0_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_0/N2  ( .A1(\SB1_0_28/i0[8] ), .A2(
        \SB1_0_28/i0[7] ), .A3(\SB1_0_28/i0[6] ), .ZN(
        \SB1_0_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_28/Component_Function_0/N1  ( .A1(\SB1_0_28/i0[10] ), .A2(
        \SB1_0_28/i0[9] ), .ZN(\SB1_0_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_1/N3  ( .A1(\SB1_0_28/i1_5 ), .A2(
        \SB1_0_28/i0[6] ), .A3(\SB1_0_28/i0[9] ), .ZN(
        \SB1_0_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_28/Component_Function_1/N2  ( .A1(\SB1_0_28/i0_3 ), .A2(
        \SB1_0_28/i1_7 ), .A3(\SB1_0_28/i0[8] ), .ZN(
        \SB1_0_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_28/Component_Function_1/N1  ( .A1(\SB1_0_28/i0_3 ), .A2(
        \SB1_0_28/i1[9] ), .ZN(\SB1_0_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_5/N2  ( .A1(\SB1_0_28/i0_0 ), .A2(
        \SB1_0_28/i0[6] ), .A3(\SB1_0_28/i0[10] ), .ZN(
        \SB1_0_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_29/Component_Function_0/N2  ( .A1(\SB1_0_29/i0[8] ), .A2(
        \SB1_0_29/i0[7] ), .A3(\SB1_0_29/i0[6] ), .ZN(
        \SB1_0_29/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_29/Component_Function_1/N4  ( .A1(\SB1_0_29/i1_7 ), .A2(
        \SB1_0_29/i0[8] ), .A3(\SB1_0_29/i0_4 ), .ZN(
        \SB1_0_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_29/Component_Function_1/N3  ( .A1(\SB1_0_29/i1_5 ), .A2(
        \SB1_0_29/i0[6] ), .A3(\SB1_0_29/i0[9] ), .ZN(
        \SB1_0_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_29/Component_Function_1/N2  ( .A1(\SB1_0_29/i0_3 ), .A2(
        \SB1_0_29/i1_7 ), .A3(\SB1_0_29/i0[8] ), .ZN(
        \SB1_0_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_29/Component_Function_1/N1  ( .A1(\SB1_0_29/i0_3 ), .A2(
        \SB1_0_29/i1[9] ), .ZN(\SB1_0_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_0/N2  ( .A1(\SB1_0_30/i0[8] ), .A2(
        \SB1_0_30/i0[7] ), .A3(\SB1_0_30/i0[6] ), .ZN(
        \SB1_0_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_30/Component_Function_0/N1  ( .A1(\SB1_0_30/i0[10] ), .A2(
        \SB1_0_30/i0[9] ), .ZN(\SB1_0_30/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_30/Component_Function_1/N1  ( .A1(\SB1_0_30/i0_3 ), .A2(
        \SB1_0_30/i1[9] ), .ZN(\SB1_0_30/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_30/Component_Function_5/N1  ( .A1(\SB1_0_30/i0_0 ), .A2(
        \SB1_0_30/i3[0] ), .ZN(\SB1_0_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_0/N2  ( .A1(\SB1_0_31/i0[8] ), .A2(
        \SB1_0_31/i0[7] ), .A3(\SB1_0_31/i0[6] ), .ZN(
        \SB1_0_31/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_31/Component_Function_1/N3  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0[6] ), .A3(\SB1_0_31/i0[9] ), .ZN(
        \SB1_0_31/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_31/Component_Function_1/N1  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i1[9] ), .ZN(\SB1_0_31/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_31/Component_Function_5/N1  ( .A1(\SB1_0_31/i0_0 ), .A2(
        \SB1_0_31/i3[0] ), .ZN(\SB1_0_31/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_0/Component_Function_5/N1  ( .A1(\SB2_0_0/i0_0 ), .A2(
        \SB2_0_0/i3[0] ), .ZN(\SB2_0_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_0/N4  ( .A1(\SB2_0_1/i0[7] ), .A2(
        \SB2_0_1/i0_3 ), .A3(\SB2_0_1/i0_0 ), .ZN(
        \SB2_0_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_1/Component_Function_0/N2  ( .A1(\SB2_0_1/i0[8] ), .A2(
        \SB2_0_1/i0[7] ), .A3(\SB2_0_1/i0[6] ), .ZN(
        \SB2_0_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_1/Component_Function_0/N1  ( .A1(\SB2_0_1/i0[10] ), .A2(
        \SB2_0_1/i0[9] ), .ZN(\SB2_0_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_1/N3  ( .A1(\SB2_0_1/i1_5 ), .A2(
        \SB2_0_1/i0[6] ), .A3(\SB2_0_1/i0[9] ), .ZN(
        \SB2_0_1/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_1/Component_Function_1/N1  ( .A1(\SB2_0_1/i0_3 ), .A2(
        \SB2_0_1/i1[9] ), .ZN(\SB2_0_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_0/N2  ( .A1(\SB2_0_2/i0[8] ), .A2(
        \SB2_0_2/i0[7] ), .A3(\SB2_0_2/i0[6] ), .ZN(
        \SB2_0_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_2/Component_Function_0/N1  ( .A1(\SB2_0_2/i0[10] ), .A2(
        \SB2_0_2/i0[9] ), .ZN(\SB2_0_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_1/N4  ( .A1(\SB2_0_2/i1_7 ), .A2(
        \SB2_0_2/i0[8] ), .A3(\RI3[0][178] ), .ZN(
        \SB2_0_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_2/Component_Function_1/N3  ( .A1(\SB2_0_2/i1_5 ), .A2(
        \SB2_0_2/i0[6] ), .A3(\SB2_0_2/i0[9] ), .ZN(
        \SB2_0_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_2/Component_Function_1/N2  ( .A1(\SB2_0_2/i0_3 ), .A2(
        \SB2_0_2/i1_7 ), .A3(\SB2_0_2/i0[8] ), .ZN(
        \SB2_0_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_2/Component_Function_1/N1  ( .A1(\SB2_0_2/i0_3 ), .A2(
        \SB2_0_2/i1[9] ), .ZN(\SB2_0_2/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_2/Component_Function_5/N1  ( .A1(\SB2_0_2/i0_0 ), .A2(
        \SB2_0_2/i3[0] ), .ZN(\SB2_0_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_3/Component_Function_1/N4  ( .A1(\SB2_0_3/i1_7 ), .A2(
        \SB2_0_3/i0[8] ), .A3(\RI3[0][172] ), .ZN(
        \SB2_0_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_3/Component_Function_1/N2  ( .A1(\SB2_0_3/i0_3 ), .A2(
        \SB2_0_3/i1_7 ), .A3(\SB2_0_3/i0[8] ), .ZN(
        \SB2_0_3/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_4/Component_Function_0/N2  ( .A1(\SB2_0_4/i0[8] ), .A2(
        \SB2_0_4/i0[7] ), .A3(\SB2_0_4/i0[6] ), .ZN(
        \SB2_0_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_4/Component_Function_0/N1  ( .A1(\SB2_0_4/i0[10] ), .A2(
        \SB2_0_4/i0[9] ), .ZN(\SB2_0_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_4/Component_Function_1/N3  ( .A1(\SB2_0_4/i1_5 ), .A2(
        \SB2_0_4/i0[6] ), .A3(\SB2_0_4/i0[9] ), .ZN(
        \SB2_0_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_4/Component_Function_1/N2  ( .A1(\SB2_0_4/i0_3 ), .A2(
        \SB2_0_4/i1_7 ), .A3(\SB2_0_4/i0[8] ), .ZN(
        \SB2_0_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_4/Component_Function_1/N1  ( .A1(\SB2_0_4/i0_3 ), .A2(
        \SB2_0_4/i1[9] ), .ZN(\SB2_0_4/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_4/Component_Function_5/N1  ( .A1(\SB2_0_4/i0_0 ), .A2(n630), 
        .ZN(\SB2_0_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_0/N3  ( .A1(\SB2_0_5/i0[10] ), .A2(
        \SB2_0_5/i0_4 ), .A3(\SB2_0_5/i0_3 ), .ZN(
        \SB2_0_5/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_5/Component_Function_0/N1  ( .A1(\SB2_0_5/i0[10] ), .A2(
        \SB2_0_5/i0[9] ), .ZN(\SB2_0_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_1/N3  ( .A1(n6282), .A2(\SB2_0_5/i0[6] ), .A3(\SB2_0_5/i0[9] ), .ZN(\SB2_0_5/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_5/Component_Function_1/N1  ( .A1(\SB2_0_5/i0_3 ), .A2(
        \SB2_0_5/i1[9] ), .ZN(\SB2_0_5/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_5/Component_Function_5/N1  ( .A1(\SB2_0_5/i0_0 ), .A2(
        \SB2_0_5/i3[0] ), .ZN(\SB2_0_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_1/N3  ( .A1(\SB2_0_6/i1_5 ), .A2(
        \SB2_0_6/i0[6] ), .A3(\RI3[0][150] ), .ZN(
        \SB2_0_6/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_6/Component_Function_1/N1  ( .A1(\SB2_0_6/i0_3 ), .A2(
        \SB2_0_6/i1[9] ), .ZN(\SB2_0_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_0/N3  ( .A1(\SB2_0_7/i0[10] ), .A2(
        \RI3[0][148] ), .A3(\SB2_0_7/i0_3 ), .ZN(
        \SB2_0_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_7/Component_Function_0/N2  ( .A1(\SB2_0_7/i0[8] ), .A2(
        \SB2_0_7/i0[7] ), .A3(\SB2_0_7/i0[6] ), .ZN(
        \SB2_0_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_7/Component_Function_0/N1  ( .A1(\SB2_0_7/i0[10] ), .A2(
        \SB2_0_7/i0[9] ), .ZN(\SB2_0_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_1/N3  ( .A1(\SB2_0_7/i1_5 ), .A2(
        \SB2_0_7/i0[6] ), .A3(\SB2_0_7/i0[9] ), .ZN(
        \SB2_0_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_7/Component_Function_1/N2  ( .A1(\SB2_0_7/i0_3 ), .A2(
        \SB2_0_7/i1_7 ), .A3(\SB2_0_7/i0[8] ), .ZN(
        \SB2_0_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_7/Component_Function_1/N1  ( .A1(\SB2_0_7/i0_3 ), .A2(
        \SB2_0_7/i1[9] ), .ZN(\SB2_0_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_8/Component_Function_0/N4  ( .A1(\SB2_0_8/i0[7] ), .A2(
        \SB2_0_8/i0_3 ), .A3(\RI3[0][140] ), .ZN(
        \SB2_0_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_8/Component_Function_1/N3  ( .A1(\SB2_0_8/i1_5 ), .A2(
        \RI3[0][139] ), .A3(\SB2_0_8/i0[9] ), .ZN(
        \SB2_0_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_8/Component_Function_1/N2  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \SB2_0_8/i1_7 ), .A3(\SB2_0_8/i0[8] ), .ZN(
        \SB2_0_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_9/Component_Function_0/N3  ( .A1(\SB2_0_9/i0[10] ), .A2(
        \SB2_0_9/i0_4 ), .A3(\SB2_0_9/i0_3 ), .ZN(
        \SB2_0_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_9/Component_Function_0/N2  ( .A1(\SB2_0_9/i0[8] ), .A2(
        \SB2_0_9/i0[7] ), .A3(\SB2_0_9/i0[6] ), .ZN(
        \SB2_0_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_9/Component_Function_0/N1  ( .A1(\SB2_0_9/i0[10] ), .A2(
        \SB2_0_9/i0[9] ), .ZN(\SB2_0_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_9/Component_Function_1/N4  ( .A1(\SB2_0_9/i1_7 ), .A2(
        \SB2_0_9/i0[8] ), .A3(\RI3[0][136] ), .ZN(
        \SB2_0_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_9/Component_Function_1/N3  ( .A1(\SB2_0_9/i1_5 ), .A2(
        \SB2_0_9/i0[6] ), .A3(\SB2_0_9/i0[9] ), .ZN(
        \SB2_0_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_9/Component_Function_1/N2  ( .A1(\SB2_0_9/i0_3 ), .A2(
        \SB2_0_9/i1_7 ), .A3(\SB2_0_9/i0[8] ), .ZN(
        \SB2_0_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_9/Component_Function_1/N1  ( .A1(\SB2_0_9/i0_3 ), .A2(
        \SB2_0_9/i1[9] ), .ZN(\SB2_0_9/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_9/Component_Function_5/N1  ( .A1(n2886), .A2(\SB2_0_9/i3[0] ), .ZN(\SB2_0_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_0/N3  ( .A1(\SB2_0_10/i0[10] ), .A2(
        \SB2_0_10/i0_4 ), .A3(\SB2_0_10/i0_3 ), .ZN(
        \SB2_0_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_10/Component_Function_0/N2  ( .A1(\SB2_0_10/i0[8] ), .A2(
        n2965), .A3(\SB2_0_10/i0[6] ), .ZN(
        \SB2_0_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_10/Component_Function_0/N1  ( .A1(\SB2_0_10/i0[10] ), .A2(
        \SB2_0_10/i0[9] ), .ZN(\SB2_0_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_1/N2  ( .A1(\SB2_0_10/i0_3 ), .A2(
        \SB2_0_10/i1_7 ), .A3(\SB2_0_10/i0[8] ), .ZN(
        \SB2_0_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_10/Component_Function_1/N1  ( .A1(\SB2_0_10/i0_3 ), .A2(
        \SB2_0_10/i1[9] ), .ZN(\SB2_0_10/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_10/Component_Function_5/N1  ( .A1(\RI3[0][128] ), .A2(
        \SB2_0_10/i3[0] ), .ZN(\SB2_0_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_0/N2  ( .A1(\SB2_0_11/i0[8] ), .A2(
        \SB2_0_11/i0[7] ), .A3(\SB2_0_11/i0[6] ), .ZN(
        \SB2_0_11/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_11/Component_Function_1/N3  ( .A1(\SB2_0_11/i1_5 ), .A2(
        \RI3[0][121] ), .A3(\SB2_0_11/i0[9] ), .ZN(
        \SB2_0_11/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_11/Component_Function_1/N1  ( .A1(\SB2_0_11/i0_3 ), .A2(
        \SB2_0_11/i1[9] ), .ZN(\SB2_0_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_0/N4  ( .A1(\SB2_0_12/i0[7] ), .A2(
        \RI3[0][119] ), .A3(\SB2_0_12/i0_0 ), .ZN(
        \SB2_0_12/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_12/Component_Function_0/N1  ( .A1(\SB2_0_12/i0[10] ), .A2(
        \SB2_0_12/i0[9] ), .ZN(\SB2_0_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_1/N4  ( .A1(\SB2_0_12/i1_7 ), .A2(
        \SB2_0_12/i0[8] ), .A3(\RI3[0][118] ), .ZN(
        \SB2_0_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_12/Component_Function_1/N2  ( .A1(\RI3[0][119] ), .A2(
        \SB2_0_12/i1_7 ), .A3(\SB2_0_12/i0[8] ), .ZN(
        \SB2_0_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_12/Component_Function_1/N1  ( .A1(\RI3[0][119] ), .A2(
        \SB2_0_12/i1[9] ), .ZN(\SB2_0_12/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_12/Component_Function_5/N1  ( .A1(\SB2_0_12/i0_0 ), .A2(
        \SB2_0_12/i3[0] ), .ZN(\SB2_0_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_0/N3  ( .A1(\SB2_0_13/i0[10] ), .A2(
        \RI3[0][112] ), .A3(\SB2_0_13/i0_3 ), .ZN(
        \SB2_0_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_13/Component_Function_0/N2  ( .A1(\SB2_0_13/i0[8] ), .A2(
        \SB2_0_13/i0[7] ), .A3(\SB2_0_13/i0[6] ), .ZN(
        \SB2_0_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_13/Component_Function_0/N1  ( .A1(\SB2_0_13/i0[10] ), .A2(
        \SB2_0_13/i0[9] ), .ZN(\SB2_0_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_1/N4  ( .A1(\SB2_0_13/i1_7 ), .A2(
        \SB2_0_13/i0[8] ), .A3(\SB1_0_14/buf_output[4] ), .ZN(
        \SB2_0_13/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_13/Component_Function_1/N1  ( .A1(\SB2_0_13/i0_3 ), .A2(
        \SB2_0_13/i1[9] ), .ZN(\SB2_0_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_14/Component_Function_0/N4  ( .A1(n2822), .A2(
        \SB2_0_14/i0_3 ), .A3(\SB2_0_14/i0_0 ), .ZN(
        \SB2_0_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_14/Component_Function_0/N3  ( .A1(\SB2_0_14/i0[10] ), .A2(
        \SB2_0_14/i0_4 ), .A3(\SB2_0_14/i0_3 ), .ZN(
        \SB2_0_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_14/Component_Function_0/N2  ( .A1(\SB2_0_14/i0[8] ), .A2(
        n2822), .A3(\SB2_0_14/i0[6] ), .ZN(
        \SB2_0_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_14/Component_Function_0/N1  ( .A1(\SB2_0_14/i0[10] ), .A2(
        \SB2_0_14/i0[9] ), .ZN(\SB2_0_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_14/Component_Function_1/N2  ( .A1(\SB2_0_14/i0_3 ), .A2(
        \SB2_0_14/i1_7 ), .A3(\SB2_0_14/i0[8] ), .ZN(
        \SB2_0_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_14/Component_Function_1/N1  ( .A1(\SB2_0_14/i0_3 ), .A2(
        \SB2_0_14/i1[9] ), .ZN(\SB2_0_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_0/N4  ( .A1(\SB2_0_15/i0[7] ), .A2(
        \SB2_0_15/i0_3 ), .A3(\SB1_0_18/buf_output[2] ), .ZN(
        \SB2_0_15/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_15/Component_Function_0/N1  ( .A1(\SB2_0_15/i0[10] ), .A2(
        \SB2_0_15/i0[9] ), .ZN(\SB2_0_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_1/N4  ( .A1(\SB2_0_15/i1_7 ), .A2(
        \SB2_0_15/i0[8] ), .A3(\RI3[0][100] ), .ZN(
        \SB2_0_15/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_15/Component_Function_5/N1  ( .A1(\SB1_0_18/buf_output[2] ), 
        .A2(\SB2_0_15/i3[0] ), .ZN(\SB2_0_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_16/Component_Function_0/N2  ( .A1(\SB2_0_16/i0[8] ), .A2(
        \SB2_0_16/i0[7] ), .A3(\SB2_0_16/i0[6] ), .ZN(
        \SB2_0_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_16/Component_Function_0/N1  ( .A1(\RI3[0][93] ), .A2(
        \SB2_0_16/i0[9] ), .ZN(\SB2_0_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_17/Component_Function_0/N2  ( .A1(\SB2_0_17/i0[8] ), .A2(
        \SB2_0_17/i0[7] ), .A3(\SB2_0_17/i0[6] ), .ZN(
        \SB2_0_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_17/Component_Function_0/N1  ( .A1(\SB2_0_17/i0[10] ), .A2(
        \SB2_0_17/i0[9] ), .ZN(\SB2_0_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_17/Component_Function_1/N4  ( .A1(\SB2_0_17/i1_7 ), .A2(
        \SB2_0_17/i0[8] ), .A3(\RI3[0][88] ), .ZN(
        \SB2_0_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_17/Component_Function_1/N2  ( .A1(\SB2_0_17/i0_3 ), .A2(
        \SB2_0_17/i1_7 ), .A3(\SB2_0_17/i0[8] ), .ZN(
        \SB2_0_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_17/Component_Function_1/N1  ( .A1(\SB2_0_17/i0_3 ), .A2(
        \SB2_0_17/i1[9] ), .ZN(\SB2_0_17/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_18/Component_Function_0/N1  ( .A1(\SB2_0_18/i0[10] ), .A2(
        \SB2_0_18/i0[9] ), .ZN(\SB2_0_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_19/Component_Function_0/N1  ( .A1(\RI3[0][75] ), .A2(
        \SB2_0_19/i0[9] ), .ZN(\SB2_0_19/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_19/Component_Function_1/N1  ( .A1(\RI3[0][77] ), .A2(
        \SB2_0_19/i1[9] ), .ZN(\SB2_0_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_19/Component_Function_5/N1  ( .A1(\SB1_0_22/buf_output[2] ), 
        .A2(\SB2_0_19/i3[0] ), .ZN(\SB2_0_19/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_20/Component_Function_0/N1  ( .A1(\SB2_0_20/i0[10] ), .A2(
        \SB2_0_20/i0[9] ), .ZN(\SB2_0_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_20/Component_Function_1/N1  ( .A1(\SB2_0_20/i0_3 ), .A2(
        \SB2_0_20/i1[9] ), .ZN(\SB2_0_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_21/Component_Function_0/N3  ( .A1(\SB2_0_21/i0[10] ), .A2(
        \SB2_0_21/i0_4 ), .A3(\SB2_0_21/i0_3 ), .ZN(
        \SB2_0_21/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_21/Component_Function_0/N1  ( .A1(\SB2_0_21/i0[10] ), .A2(
        \SB2_0_21/i0[9] ), .ZN(\SB2_0_21/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_21/Component_Function_5/N1  ( .A1(\RI3[0][62] ), .A2(
        \SB2_0_21/i3[0] ), .ZN(\SB2_0_21/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_22/Component_Function_5/N1  ( .A1(\SB2_0_22/i0_0 ), .A2(
        \SB2_0_22/i3[0] ), .ZN(\SB2_0_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_23/Component_Function_0/N4  ( .A1(\SB2_0_23/i0[7] ), .A2(
        \SB2_0_23/i0_3 ), .A3(\SB2_0_23/i0_0 ), .ZN(
        \SB2_0_23/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_23/Component_Function_0/N1  ( .A1(\SB2_0_23/i0[10] ), .A2(
        \SB2_0_23/i0[9] ), .ZN(\SB2_0_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_23/Component_Function_1/N2  ( .A1(\SB2_0_23/i0_3 ), .A2(
        \SB2_0_23/i1_7 ), .A3(\SB2_0_23/i0[8] ), .ZN(
        \SB2_0_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_24/Component_Function_0/N4  ( .A1(\SB2_0_24/i0[7] ), .A2(
        \SB2_0_24/i0_3 ), .A3(\SB2_0_24/i0_0 ), .ZN(
        \SB2_0_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_24/Component_Function_0/N3  ( .A1(\SB2_0_24/i0[10] ), .A2(
        \RI3[0][46] ), .A3(\SB2_0_24/i0_3 ), .ZN(
        \SB2_0_24/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_24/Component_Function_0/N1  ( .A1(\SB2_0_24/i0[10] ), .A2(
        \RI3[0][42] ), .ZN(\SB2_0_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_24/Component_Function_1/N4  ( .A1(\SB2_0_24/i1_7 ), .A2(
        \SB2_0_24/i0[8] ), .A3(\RI3[0][46] ), .ZN(
        \SB2_0_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_24/Component_Function_1/N3  ( .A1(\SB2_0_24/i1_5 ), .A2(
        \SB2_0_24/i0[6] ), .A3(\RI3[0][42] ), .ZN(
        \SB2_0_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_1/N2  ( .A1(\SB2_0_24/i0_3 ), .A2(
        \SB2_0_24/i1_7 ), .A3(\SB2_0_24/i0[8] ), .ZN(
        \SB2_0_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_24/Component_Function_1/N1  ( .A1(\SB2_0_24/i0_3 ), .A2(
        \SB2_0_24/i1[9] ), .ZN(\SB2_0_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_25/Component_Function_0/N2  ( .A1(\SB2_0_25/i0[8] ), .A2(
        n2978), .A3(\SB2_0_25/i0[6] ), .ZN(
        \SB2_0_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_25/Component_Function_0/N1  ( .A1(\SB2_0_25/i0[10] ), .A2(
        \SB2_0_25/i0[9] ), .ZN(\SB2_0_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_25/Component_Function_1/N4  ( .A1(\SB2_0_25/i1_7 ), .A2(
        \SB2_0_25/i0[8] ), .A3(\SB2_0_25/i0_4 ), .ZN(
        \SB2_0_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_25/Component_Function_1/N2  ( .A1(\SB2_0_25/i0_3 ), .A2(
        \SB2_0_25/i1_7 ), .A3(\SB2_0_25/i0[8] ), .ZN(
        \SB2_0_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_25/Component_Function_1/N1  ( .A1(\SB2_0_25/i0_3 ), .A2(
        \SB2_0_25/i1[9] ), .ZN(\SB2_0_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_0/N3  ( .A1(\RI3[0][33] ), .A2(
        \SB2_0_26/i0_4 ), .A3(\SB2_0_26/i0_3 ), .ZN(
        \SB2_0_26/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_26/Component_Function_0/N1  ( .A1(\RI3[0][33] ), .A2(
        \SB2_0_26/i0[9] ), .ZN(\SB2_0_26/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_26/Component_Function_1/N1  ( .A1(\SB2_0_26/i0_3 ), .A2(
        \SB2_0_26/i1[9] ), .ZN(\SB2_0_26/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_26/Component_Function_5/N1  ( .A1(\SB2_0_26/i0_0 ), .A2(
        \SB2_0_26/i3[0] ), .ZN(\SB2_0_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_27/Component_Function_0/N4  ( .A1(\SB2_0_27/i0[7] ), .A2(
        \SB2_0_27/i0_3 ), .A3(\SB2_0_27/i0_0 ), .ZN(
        \SB2_0_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_27/Component_Function_0/N3  ( .A1(\SB2_0_27/i0[10] ), .A2(
        \RI3[0][28] ), .A3(\SB2_0_27/i0_3 ), .ZN(
        \SB2_0_27/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_27/Component_Function_0/N1  ( .A1(\SB2_0_27/i0[10] ), .A2(
        \SB2_0_27/i0[9] ), .ZN(\SB2_0_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_27/Component_Function_1/N3  ( .A1(\SB2_0_27/i1_5 ), .A2(
        \SB2_0_27/i0[6] ), .A3(\SB2_0_27/i0[9] ), .ZN(
        \SB2_0_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_27/Component_Function_1/N2  ( .A1(\SB2_0_27/i0_3 ), .A2(
        \SB2_0_27/i1_7 ), .A3(\SB2_0_27/i0[8] ), .ZN(
        \SB2_0_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_27/Component_Function_1/N1  ( .A1(\SB2_0_27/i0_3 ), .A2(
        \SB2_0_27/i1[9] ), .ZN(\SB2_0_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_0/N2  ( .A1(\SB2_0_28/i0[8] ), .A2(
        \SB2_0_28/i0[7] ), .A3(\SB2_0_28/i0[6] ), .ZN(
        \SB2_0_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_28/Component_Function_0/N1  ( .A1(\SB2_0_28/i0[10] ), .A2(
        \SB2_0_28/i0[9] ), .ZN(\SB2_0_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_1/N4  ( .A1(\SB2_0_28/i1_7 ), .A2(
        \SB2_0_28/i0[8] ), .A3(\SB2_0_28/i0_4 ), .ZN(
        \SB2_0_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_28/Component_Function_1/N2  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i1_7 ), .A3(\SB2_0_28/i0[8] ), .ZN(
        \SB2_0_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_28/Component_Function_1/N1  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i1[9] ), .ZN(\SB2_0_28/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_28/Component_Function_5/N1  ( .A1(\SB2_0_28/i0_0 ), .A2(
        \SB2_0_28/i3[0] ), .ZN(\SB2_0_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_0/N4  ( .A1(n2657), .A2(
        \SB2_0_29/i0_3 ), .A3(\SB2_0_29/i0_0 ), .ZN(
        \SB2_0_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_29/Component_Function_0/N2  ( .A1(\SB2_0_29/i0[8] ), .A2(
        n2657), .A3(\SB2_0_29/i0[6] ), .ZN(
        \SB2_0_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_29/Component_Function_0/N1  ( .A1(\SB2_0_29/i0[10] ), .A2(
        \SB2_0_29/i0[9] ), .ZN(\SB2_0_29/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_29/Component_Function_1/N1  ( .A1(\SB2_0_29/i0_3 ), .A2(
        \SB2_0_29/i1[9] ), .ZN(\SB2_0_29/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_29/Component_Function_5/N1  ( .A1(\SB2_0_29/i0_0 ), .A2(
        \SB2_0_29/i3[0] ), .ZN(\SB2_0_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_0/N2  ( .A1(\SB2_0_30/i0[8] ), .A2(
        \SB2_0_30/i0[7] ), .A3(\SB2_0_30/i0[6] ), .ZN(
        \SB2_0_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_30/Component_Function_0/N1  ( .A1(\SB2_0_30/i0[10] ), .A2(
        \SB2_0_30/i0[9] ), .ZN(\SB2_0_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_1/N3  ( .A1(\SB2_0_30/i1_5 ), .A2(
        \SB2_0_30/i0[6] ), .A3(\SB2_0_30/i0[9] ), .ZN(
        \SB2_0_30/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_30/Component_Function_1/N1  ( .A1(\SB2_0_30/i0_3 ), .A2(
        \SB2_0_30/i1[9] ), .ZN(\SB2_0_30/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_30/Component_Function_5/N1  ( .A1(\SB2_0_30/i0_0 ), .A2(
        \SB2_0_30/i3[0] ), .ZN(\SB2_0_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_0/N3  ( .A1(\SB2_0_31/i0[10] ), .A2(
        \RI3[0][4] ), .A3(\SB2_0_31/i0_3 ), .ZN(
        \SB2_0_31/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_31/Component_Function_0/N1  ( .A1(\SB2_0_31/i0[10] ), .A2(
        \SB2_0_31/i0[9] ), .ZN(\SB2_0_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_1/N4  ( .A1(\SB2_0_31/i1_7 ), .A2(
        \SB2_0_31/i0[8] ), .A3(\RI3[0][4] ), .ZN(
        \SB2_0_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_31/Component_Function_1/N2  ( .A1(\SB2_0_31/i0_3 ), .A2(
        \SB2_0_31/i1_7 ), .A3(\SB2_0_31/i0[8] ), .ZN(
        \SB2_0_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_31/Component_Function_1/N1  ( .A1(\SB2_0_31/i0_3 ), .A2(
        \SB2_0_31/i1[9] ), .ZN(\SB2_0_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_0/N3  ( .A1(\SB1_1_0/i0[10] ), .A2(
        \SB1_1_0/i0_4 ), .A3(\SB1_1_0/i0_3 ), .ZN(
        \SB1_1_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_0/Component_Function_0/N2  ( .A1(\SB1_1_0/i0[8] ), .A2(
        \SB1_1_0/i0[7] ), .A3(\SB1_1_0/i0[6] ), .ZN(
        \SB1_1_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_0/Component_Function_0/N1  ( .A1(\SB1_1_0/i0[10] ), .A2(
        \SB1_1_0/i0[9] ), .ZN(\SB1_1_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_1/Component_Function_0/N2  ( .A1(\SB1_1_1/i0[8] ), .A2(
        \SB1_1_1/i0[7] ), .A3(\SB1_1_1/i0[6] ), .ZN(
        \SB1_1_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_1/Component_Function_0/N1  ( .A1(\SB1_1_1/i0[10] ), .A2(
        \SB1_1_1/i0[9] ), .ZN(\SB1_1_1/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_1/Component_Function_1/N1  ( .A1(\SB1_1_1/i0_3 ), .A2(
        \SB1_1_1/i1[9] ), .ZN(\SB1_1_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_2/Component_Function_0/N2  ( .A1(\SB1_1_2/i0[8] ), .A2(
        \SB1_1_2/i0[7] ), .A3(\SB1_1_2/i0[6] ), .ZN(
        \SB1_1_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_2/Component_Function_0/N1  ( .A1(\SB1_1_2/i0[10] ), .A2(
        \SB1_1_2/i0[9] ), .ZN(\SB1_1_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_2/Component_Function_1/N2  ( .A1(\SB1_1_2/i0_3 ), .A2(
        \SB1_1_2/i1_7 ), .A3(\SB1_1_2/i0[8] ), .ZN(
        \SB1_1_2/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_3/Component_Function_0/N4  ( .A1(\SB1_1_3/i0[7] ), .A2(
        \SB1_1_3/i0_3 ), .A3(\SB1_1_3/i0_0 ), .ZN(
        \SB1_1_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_3/Component_Function_0/N2  ( .A1(\SB1_1_3/i0[8] ), .A2(
        \SB1_1_3/i0[7] ), .A3(\SB1_1_3/i0[6] ), .ZN(
        \SB1_1_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_3/Component_Function_0/N1  ( .A1(\SB1_1_3/i0[10] ), .A2(
        \SB1_1_3/i0[9] ), .ZN(\SB1_1_3/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_4/Component_Function_0/N1  ( .A1(\SB1_1_4/i0[10] ), .A2(
        \SB1_1_4/i0[9] ), .ZN(\SB1_1_4/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_4/Component_Function_1/N1  ( .A1(\SB1_1_4/i0_3 ), .A2(
        \SB1_1_4/i1[9] ), .ZN(\SB1_1_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_0/N4  ( .A1(\SB1_1_5/i0[7] ), .A2(
        \SB1_1_5/i0_3 ), .A3(\SB1_1_5/i0_0 ), .ZN(
        \SB1_1_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_5/Component_Function_0/N3  ( .A1(\SB1_1_5/i0[10] ), .A2(
        \SB1_1_5/i0_4 ), .A3(\SB1_1_5/i0_3 ), .ZN(
        \SB1_1_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_5/Component_Function_0/N2  ( .A1(\SB1_1_5/i0[8] ), .A2(
        \SB1_1_5/i0[7] ), .A3(\SB1_1_5/i0[6] ), .ZN(
        \SB1_1_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_5/Component_Function_0/N1  ( .A1(\SB1_1_5/i0[10] ), .A2(
        \SB1_1_5/i0[9] ), .ZN(\SB1_1_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_1/N2  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i1_7 ), .A3(\SB1_1_5/i0[8] ), .ZN(
        \SB1_1_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_5/Component_Function_1/N1  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i1[9] ), .ZN(\SB1_1_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_0/N2  ( .A1(\SB1_1_6/i0[8] ), .A2(
        \SB1_1_6/i0[7] ), .A3(\SB1_1_6/i0[6] ), .ZN(
        \SB1_1_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_6/Component_Function_0/N1  ( .A1(\SB1_1_6/i0[10] ), .A2(
        \SB1_1_6/i0[9] ), .ZN(\SB1_1_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_1/N2  ( .A1(\SB1_1_6/i0_3 ), .A2(
        \SB1_1_6/i1_7 ), .A3(\SB1_1_6/i0[8] ), .ZN(
        \SB1_1_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_6/Component_Function_1/N1  ( .A1(\SB1_1_6/i0_3 ), .A2(
        \SB1_1_6/i1[9] ), .ZN(\SB1_1_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_0/N2  ( .A1(\SB1_1_7/i0[8] ), .A2(
        \SB1_1_7/i0[7] ), .A3(\SB1_1_7/i0[6] ), .ZN(
        \SB1_1_7/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_7/Component_Function_1/N2  ( .A1(\SB1_1_7/i0_3 ), .A2(
        \SB1_1_7/i1_7 ), .A3(\SB1_1_7/i0[8] ), .ZN(
        \SB1_1_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_8/Component_Function_1/N4  ( .A1(\SB1_1_8/i1_7 ), .A2(
        \SB1_1_8/i0[8] ), .A3(\SB1_1_8/i0_4 ), .ZN(
        \SB1_1_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_8/Component_Function_1/N2  ( .A1(\SB1_1_8/i0_3 ), .A2(
        \SB1_1_8/i1_7 ), .A3(\SB1_1_8/i0[8] ), .ZN(
        \SB1_1_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_9/Component_Function_0/N2  ( .A1(\SB1_1_9/i0[8] ), .A2(
        \SB1_1_9/i0[7] ), .A3(\SB1_1_9/i0[6] ), .ZN(
        \SB1_1_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_9/Component_Function_0/N1  ( .A1(\SB1_1_9/i0[10] ), .A2(
        \SB1_1_9/i0[9] ), .ZN(\SB1_1_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_1/N2  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i1_7 ), .A3(\SB1_1_9/i0[8] ), .ZN(
        \SB1_1_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_9/Component_Function_1/N1  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i1[9] ), .ZN(\SB1_1_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_0/N3  ( .A1(\SB1_1_10/i0[10] ), .A2(
        \SB1_1_10/i0_4 ), .A3(\SB1_1_10/i0_3 ), .ZN(
        \SB1_1_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_10/Component_Function_0/N2  ( .A1(\SB1_1_10/i0[8] ), .A2(
        \SB1_1_10/i0[7] ), .A3(\SB1_1_10/i0[6] ), .ZN(
        \SB1_1_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_10/Component_Function_0/N1  ( .A1(\SB1_1_10/i0[10] ), .A2(
        \SB1_1_10/i0[9] ), .ZN(\SB1_1_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_10/Component_Function_1/N1  ( .A1(\SB1_1_10/i0_3 ), .A2(
        \SB1_1_10/i1[9] ), .ZN(\SB1_1_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_5/N2  ( .A1(\SB1_1_10/i0_0 ), .A2(
        \SB1_1_10/i0[6] ), .A3(\SB1_1_10/i0[10] ), .ZN(
        \SB1_1_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_11/Component_Function_0/N4  ( .A1(\SB1_1_11/i0[7] ), .A2(
        \SB1_1_11/i0_3 ), .A3(\SB1_1_11/i0_0 ), .ZN(
        \SB1_1_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_11/Component_Function_0/N2  ( .A1(\SB1_1_11/i0[8] ), .A2(
        \SB1_1_11/i0[7] ), .A3(\SB1_1_11/i0[6] ), .ZN(
        \SB1_1_11/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_12/Component_Function_0/N2  ( .A1(\SB1_1_12/i0[8] ), .A2(
        \SB1_1_12/i0[7] ), .A3(\SB1_1_12/i0[6] ), .ZN(
        \SB1_1_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_12/Component_Function_0/N1  ( .A1(\SB1_1_12/i0[10] ), .A2(
        \SB1_1_12/i0[9] ), .ZN(\SB1_1_12/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_12/Component_Function_1/N1  ( .A1(\SB1_1_12/i0_3 ), .A2(
        \SB1_1_12/i1[9] ), .ZN(\SB1_1_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_0/N3  ( .A1(\SB1_1_13/i0[10] ), .A2(
        \SB1_1_13/i0_4 ), .A3(\SB1_1_13/i0_3 ), .ZN(
        \SB1_1_13/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_13/Component_Function_0/N1  ( .A1(\SB1_1_13/i0[10] ), .A2(
        \SB1_1_13/i0[9] ), .ZN(\SB1_1_13/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_13/Component_Function_1/N1  ( .A1(\SB1_1_13/i0_3 ), .A2(
        \SB1_1_13/i1[9] ), .ZN(\SB1_1_13/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_14/Component_Function_0/N1  ( .A1(\SB1_1_14/i0[10] ), .A2(
        \SB1_1_14/i0[9] ), .ZN(\SB1_1_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_0/N2  ( .A1(\SB1_1_15/i0[8] ), .A2(
        \SB1_1_15/i0[7] ), .A3(\SB1_1_15/i0[6] ), .ZN(
        \SB1_1_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_15/Component_Function_0/N1  ( .A1(\SB1_1_15/i0[10] ), .A2(
        \SB1_1_15/i0[9] ), .ZN(\SB1_1_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_1/N2  ( .A1(\SB1_1_15/i0_3 ), .A2(
        \SB1_1_15/i1_7 ), .A3(\SB1_1_15/i0[8] ), .ZN(
        \SB1_1_15/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_16/Component_Function_0/N3  ( .A1(\SB1_1_16/i0[10] ), .A2(
        \SB1_1_16/i0_4 ), .A3(\SB1_1_16/i0_3 ), .ZN(
        \SB1_1_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_16/Component_Function_0/N2  ( .A1(\SB1_1_16/i0[8] ), .A2(
        \SB1_1_16/i0[7] ), .A3(\SB1_1_16/i0[6] ), .ZN(
        \SB1_1_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_16/Component_Function_0/N1  ( .A1(\SB1_1_16/i0[10] ), .A2(
        \SB1_1_16/i0[9] ), .ZN(\SB1_1_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_0/N2  ( .A1(\SB1_1_17/i0[8] ), .A2(
        \SB1_1_17/i0[7] ), .A3(\SB1_1_17/i0[6] ), .ZN(
        \SB1_1_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_17/Component_Function_0/N1  ( .A1(\SB1_1_17/i0[10] ), .A2(
        \SB1_1_17/i0[9] ), .ZN(\SB1_1_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_0/N3  ( .A1(\SB1_1_18/i0[10] ), .A2(
        \SB1_1_18/i0_4 ), .A3(\SB1_1_18/i0_3 ), .ZN(
        \SB1_1_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_18/Component_Function_0/N2  ( .A1(\SB1_1_18/i0[8] ), .A2(
        \SB1_1_18/i0[7] ), .A3(\SB1_1_18/i0[6] ), .ZN(
        \SB1_1_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_18/Component_Function_0/N1  ( .A1(\SB1_1_18/i0[10] ), .A2(
        \SB1_1_18/i0[9] ), .ZN(\SB1_1_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_18/Component_Function_1/N1  ( .A1(\SB1_1_18/i0_3 ), .A2(
        \SB1_1_18/i1[9] ), .ZN(\SB1_1_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_0/N3  ( .A1(\SB1_1_19/i0[10] ), .A2(
        \SB1_1_19/i0_4 ), .A3(\SB1_1_19/i0_3 ), .ZN(
        \SB1_1_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_19/Component_Function_0/N2  ( .A1(\SB1_1_19/i0[8] ), .A2(
        \SB1_1_19/i0[7] ), .A3(\SB1_1_19/i0[6] ), .ZN(
        \SB1_1_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_19/Component_Function_0/N1  ( .A1(\SB1_1_19/i0[10] ), .A2(
        \SB1_1_19/i0[9] ), .ZN(\SB1_1_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_1/N2  ( .A1(\SB1_1_19/i0_3 ), .A2(
        \SB1_1_19/i1_7 ), .A3(\SB1_1_19/i0[8] ), .ZN(
        \SB1_1_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_19/Component_Function_1/N1  ( .A1(\SB1_1_19/i0_3 ), .A2(
        \SB1_1_19/i1[9] ), .ZN(\SB1_1_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_0/N4  ( .A1(\SB1_1_20/i0[7] ), .A2(
        \SB1_1_20/i0_3 ), .A3(\SB1_1_20/i0_0 ), .ZN(
        \SB1_1_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_20/Component_Function_0/N3  ( .A1(\SB1_1_20/i0[10] ), .A2(
        \SB1_1_20/i0_4 ), .A3(\SB1_1_20/i0_3 ), .ZN(
        \SB1_1_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_20/Component_Function_0/N2  ( .A1(\SB1_1_20/i0[8] ), .A2(
        \SB1_1_20/i0[7] ), .A3(\SB1_1_20/i0[6] ), .ZN(
        \SB1_1_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_20/Component_Function_0/N1  ( .A1(\SB1_1_20/i0[10] ), .A2(
        \SB1_1_20/i0[9] ), .ZN(\SB1_1_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_20/Component_Function_1/N1  ( .A1(\SB1_1_20/i0_3 ), .A2(
        \SB1_1_20/i1[9] ), .ZN(\SB1_1_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_0/N3  ( .A1(\SB1_1_21/i0[10] ), .A2(
        \SB1_1_21/i0_4 ), .A3(\SB1_1_21/i0_3 ), .ZN(
        \SB1_1_21/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_21/Component_Function_0/N1  ( .A1(\SB1_1_21/i0[10] ), .A2(
        \SB1_1_21/i0[9] ), .ZN(\SB1_1_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_1/N2  ( .A1(\SB1_1_21/i0_3 ), .A2(
        \SB1_1_21/i1_7 ), .A3(\SB1_1_21/i0[8] ), .ZN(
        \SB1_1_21/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_22/Component_Function_0/N2  ( .A1(\SB1_1_22/i0[8] ), .A2(
        \SB1_1_22/i0[7] ), .A3(\SB1_1_22/i0[6] ), .ZN(
        \SB1_1_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_22/Component_Function_1/N1  ( .A1(\SB1_1_22/i0_3 ), .A2(
        \SB1_1_22/i1[9] ), .ZN(\SB1_1_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_23/Component_Function_0/N3  ( .A1(\SB1_1_23/i0[10] ), .A2(
        \SB1_1_23/i0_4 ), .A3(\SB1_1_23/i0_3 ), .ZN(
        \SB1_1_23/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_23/Component_Function_0/N1  ( .A1(\SB1_1_23/i0[10] ), .A2(
        \SB1_1_23/i0[9] ), .ZN(\SB1_1_23/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_24/Component_Function_0/N1  ( .A1(\SB1_1_24/i0[10] ), .A2(
        \SB1_1_24/i0[9] ), .ZN(\SB1_1_24/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_25/Component_Function_0/N1  ( .A1(\SB1_1_25/i0[10] ), .A2(
        \SB1_1_25/i0[9] ), .ZN(\SB1_1_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_1/N2  ( .A1(\SB1_1_25/i0_3 ), .A2(
        \SB1_1_25/i1_7 ), .A3(\SB1_1_25/i0[8] ), .ZN(
        \SB1_1_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_25/Component_Function_1/N1  ( .A1(\SB1_1_25/i0_3 ), .A2(
        \SB1_1_25/i1[9] ), .ZN(\SB1_1_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_0/N4  ( .A1(\SB1_1_26/i0[7] ), .A2(
        \SB1_1_26/i0_3 ), .A3(\SB1_1_26/i0_0 ), .ZN(
        \SB1_1_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_26/Component_Function_0/N2  ( .A1(\SB1_1_26/i0[8] ), .A2(
        \SB1_1_26/i0[7] ), .A3(\SB1_1_26/i0[6] ), .ZN(
        \SB1_1_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_26/Component_Function_0/N1  ( .A1(\SB1_1_26/i0[10] ), .A2(
        \SB1_1_26/i0[9] ), .ZN(\SB1_1_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_27/Component_Function_1/N2  ( .A1(\SB1_1_27/i0_3 ), .A2(
        \SB1_1_27/i1_7 ), .A3(\SB1_1_27/i0[8] ), .ZN(
        \SB1_1_27/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_28/Component_Function_0/N3  ( .A1(\SB1_1_28/i0[10] ), .A2(
        \SB1_1_28/i0_4 ), .A3(\SB1_1_28/i0_3 ), .ZN(
        \SB1_1_28/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_28/Component_Function_0/N1  ( .A1(\SB1_1_28/i0[10] ), .A2(
        \SB1_1_28/i0[9] ), .ZN(\SB1_1_28/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_28/Component_Function_1/N1  ( .A1(\SB1_1_28/i0_3 ), .A2(
        \SB1_1_28/i1[9] ), .ZN(\SB1_1_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_0/N3  ( .A1(\SB1_1_29/i0[10] ), .A2(
        \SB1_1_29/i0_4 ), .A3(\SB1_1_29/i0_3 ), .ZN(
        \SB1_1_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_29/Component_Function_0/N2  ( .A1(\SB1_1_29/i0[8] ), .A2(
        \SB1_1_29/i0[7] ), .A3(\SB1_1_29/i0[6] ), .ZN(
        \SB1_1_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_29/Component_Function_0/N1  ( .A1(\SB1_1_29/i0[10] ), .A2(
        \SB1_1_29/i0[9] ), .ZN(\SB1_1_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_30/Component_Function_0/N3  ( .A1(\SB1_1_30/i0[10] ), .A2(
        \SB1_1_30/i0_4 ), .A3(\SB1_1_30/i0_3 ), .ZN(
        \SB1_1_30/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_30/Component_Function_0/N1  ( .A1(\SB1_1_30/i0[10] ), .A2(
        \SB1_1_30/i0[9] ), .ZN(\SB1_1_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_30/Component_Function_1/N3  ( .A1(\SB1_1_30/i1_5 ), .A2(
        \SB1_1_30/i0[6] ), .A3(\SB1_1_30/i0[9] ), .ZN(
        \SB1_1_30/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_30/Component_Function_1/N1  ( .A1(\SB1_1_30/i0_3 ), .A2(
        \SB1_1_30/i1[9] ), .ZN(\SB1_1_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_0/N3  ( .A1(\SB1_1_31/i0[10] ), .A2(
        \SB1_1_31/i0_4 ), .A3(\SB1_1_31/i0_3 ), .ZN(
        \SB1_1_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_31/Component_Function_1/N2  ( .A1(\SB1_1_31/i0_3 ), .A2(
        \SB1_1_31/i1_7 ), .A3(\SB1_1_31/i0[8] ), .ZN(
        \SB1_1_31/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_31/Component_Function_5/N2  ( .A1(\SB1_1_31/i0_0 ), .A2(
        \SB1_1_31/i0[6] ), .A3(\MC_ARK_ARC_1_0/buf_output[3] ), .ZN(
        \SB1_1_31/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_0/Component_Function_1/N1  ( .A1(\SB2_1_0/i0_3 ), .A2(
        \SB2_1_0/i1[9] ), .ZN(\SB2_1_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_1/Component_Function_0/N2  ( .A1(\SB2_1_1/i0[8] ), .A2(
        \SB2_1_1/i0[7] ), .A3(\SB2_1_1/i0[6] ), .ZN(
        \SB2_1_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_1/Component_Function_0/N1  ( .A1(\SB2_1_1/i0[10] ), .A2(
        \SB2_1_1/i0[9] ), .ZN(\SB2_1_1/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_2/Component_Function_0/N1  ( .A1(\SB2_1_2/i0[10] ), .A2(
        \SB2_1_2/i0[9] ), .ZN(\SB2_1_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_1/N3  ( .A1(\SB2_1_2/i1_5 ), .A2(
        \SB2_1_2/i0[6] ), .A3(\SB2_1_2/i0[9] ), .ZN(
        \SB2_1_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_2/Component_Function_1/N2  ( .A1(\SB2_1_2/i0_3 ), .A2(
        \SB2_1_2/i1_7 ), .A3(\SB2_1_2/i0[8] ), .ZN(
        \SB2_1_2/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_3/Component_Function_0/N2  ( .A1(\SB2_1_3/i0[8] ), .A2(
        \SB2_1_3/i0[7] ), .A3(\SB2_1_3/i0[6] ), .ZN(
        \SB2_1_3/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_3/Component_Function_1/N2  ( .A1(\SB2_1_3/i0_3 ), .A2(
        \SB2_1_3/i1_7 ), .A3(\SB2_1_3/i0[8] ), .ZN(
        \SB2_1_3/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_4/Component_Function_0/N2  ( .A1(\SB2_1_4/i0[8] ), .A2(
        \SB2_1_4/i0[7] ), .A3(\SB1_1_8/buf_output[1] ), .ZN(
        \SB2_1_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_4/Component_Function_0/N1  ( .A1(\SB2_1_4/i0[10] ), .A2(
        \SB2_1_4/i0[9] ), .ZN(\SB2_1_4/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_4/Component_Function_1/N1  ( .A1(\SB2_1_4/i0_3 ), .A2(
        \SB2_1_4/i1[9] ), .ZN(\SB2_1_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_0/N2  ( .A1(\SB2_1_5/i0[8] ), .A2(
        \SB2_1_5/i0[7] ), .A3(\SB2_1_5/i0[6] ), .ZN(
        \SB2_1_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_6/Component_Function_0/N4  ( .A1(\SB2_1_6/i0[7] ), .A2(
        \SB2_1_6/i0_3 ), .A3(\SB2_1_6/i0_0 ), .ZN(
        \SB2_1_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_6/Component_Function_1/N3  ( .A1(\SB2_1_6/i1_5 ), .A2(
        \SB2_1_6/i0[6] ), .A3(\SB1_1_11/buf_output[0] ), .ZN(
        \SB2_1_6/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_6/Component_Function_1/N1  ( .A1(\SB2_1_6/i0_3 ), .A2(
        \SB2_1_6/i1[9] ), .ZN(\SB2_1_6/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_6/Component_Function_5/N1  ( .A1(\SB2_1_6/i0_0 ), .A2(
        \SB2_1_6/i3[0] ), .ZN(\SB2_1_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_0/N4  ( .A1(\SB2_1_7/i0[7] ), .A2(
        \SB2_1_7/i0_3 ), .A3(\SB2_1_7/i0_0 ), .ZN(
        \SB2_1_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_7/Component_Function_0/N2  ( .A1(\SB2_1_7/i0[8] ), .A2(
        \SB2_1_7/i0[7] ), .A3(\SB2_1_7/i0[6] ), .ZN(
        \SB2_1_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_7/Component_Function_0/N1  ( .A1(\SB2_1_7/i0[10] ), .A2(
        \SB2_1_7/i0[9] ), .ZN(\SB2_1_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_1/N2  ( .A1(\SB2_1_7/i0_3 ), .A2(
        \SB2_1_7/i1_7 ), .A3(\SB2_1_7/i0[8] ), .ZN(
        \SB2_1_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_7/Component_Function_1/N1  ( .A1(\SB2_1_7/i0_3 ), .A2(
        \SB2_1_7/i1[9] ), .ZN(\SB2_1_7/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_8/Component_Function_0/N1  ( .A1(\SB2_1_8/i0[10] ), .A2(
        \SB2_1_8/i0[9] ), .ZN(\SB2_1_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_8/Component_Function_1/N3  ( .A1(\SB2_1_8/i1_5 ), .A2(
        \SB2_1_8/i0[6] ), .A3(\SB2_1_8/i0[9] ), .ZN(
        \SB2_1_8/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_8/Component_Function_1/N1  ( .A1(\SB2_1_8/i0_3 ), .A2(
        \SB2_1_8/i1[9] ), .ZN(\SB2_1_8/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_8/Component_Function_5/N1  ( .A1(\SB2_1_8/i0_0 ), .A2(
        \SB2_1_8/i3[0] ), .ZN(\SB2_1_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_9/Component_Function_0/N2  ( .A1(\SB2_1_9/i0[8] ), .A2(
        \SB2_1_9/i0[7] ), .A3(\SB2_1_9/i0[6] ), .ZN(
        \SB2_1_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_9/Component_Function_0/N1  ( .A1(\SB2_1_9/i0[10] ), .A2(
        \SB2_1_9/i0[9] ), .ZN(\SB2_1_9/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_9/Component_Function_5/N1  ( .A1(\SB2_1_9/i0_0 ), .A2(
        \SB2_1_9/i3[0] ), .ZN(\SB2_1_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_10/Component_Function_1/N4  ( .A1(\SB2_1_10/i1_7 ), .A2(
        \SB2_1_10/i0[8] ), .A3(\SB2_1_10/i0_4 ), .ZN(
        \SB2_1_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_10/Component_Function_1/N3  ( .A1(\SB2_1_10/i1_5 ), .A2(
        \SB2_1_10/i0[6] ), .A3(\SB2_1_10/i0[9] ), .ZN(
        \SB2_1_10/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_11/Component_Function_0/N1  ( .A1(\SB2_1_11/i0[10] ), .A2(
        \SB2_1_11/i0[9] ), .ZN(\SB2_1_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_11/Component_Function_1/N2  ( .A1(\SB2_1_11/i0_3 ), .A2(
        \SB2_1_11/i1_7 ), .A3(\SB2_1_11/i0[8] ), .ZN(
        \SB2_1_11/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_12/Component_Function_0/N2  ( .A1(\SB2_1_12/i0[8] ), .A2(
        \SB2_1_12/i0[7] ), .A3(\SB2_1_12/i0[6] ), .ZN(
        \SB2_1_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_12/Component_Function_0/N1  ( .A1(\SB2_1_12/i0[10] ), .A2(
        \SB2_1_12/i0[9] ), .ZN(\SB2_1_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_12/Component_Function_1/N2  ( .A1(\SB2_1_12/i0_3 ), .A2(
        \SB2_1_12/i1_7 ), .A3(\SB2_1_12/i0[8] ), .ZN(
        \SB2_1_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_12/Component_Function_1/N1  ( .A1(\SB2_1_12/i0_3 ), .A2(
        \SB2_1_12/i1[9] ), .ZN(\SB2_1_12/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_13/Component_Function_0/N1  ( .A1(\SB2_1_13/i0[10] ), .A2(
        \SB2_1_13/i0[9] ), .ZN(\SB2_1_13/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_13/Component_Function_1/N1  ( .A1(\SB2_1_13/i0_3 ), .A2(
        \SB2_1_13/i1[9] ), .ZN(\SB2_1_13/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_14/Component_Function_0/N1  ( .A1(\SB2_1_14/i0[10] ), .A2(
        \SB2_1_14/i0[9] ), .ZN(\SB2_1_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_14/Component_Function_1/N3  ( .A1(\SB2_1_14/i1_5 ), .A2(
        \SB2_1_14/i0[6] ), .A3(\SB2_1_14/i0[9] ), .ZN(
        \SB2_1_14/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_14/Component_Function_1/N1  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i1[9] ), .ZN(\SB2_1_14/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_15/Component_Function_0/N1  ( .A1(\SB2_1_15/i0[10] ), .A2(
        \SB2_1_15/i0[9] ), .ZN(\SB2_1_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_15/Component_Function_1/N3  ( .A1(\SB2_1_15/i1_5 ), .A2(
        \SB2_1_15/i0[6] ), .A3(\SB2_1_15/i0[9] ), .ZN(
        \SB2_1_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_16/Component_Function_1/N2  ( .A1(\SB2_1_16/i0_3 ), .A2(
        \SB2_1_16/i1_7 ), .A3(\SB2_1_16/i0[8] ), .ZN(
        \SB2_1_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_16/Component_Function_1/N1  ( .A1(\SB2_1_16/i0_3 ), .A2(
        \SB2_1_16/i1[9] ), .ZN(\SB2_1_16/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_16/Component_Function_5/N1  ( .A1(\SB2_1_16/i0_0 ), .A2(
        \SB2_1_16/i3[0] ), .ZN(\SB2_1_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_0/N4  ( .A1(\SB2_1_17/i0[7] ), .A2(
        \SB2_1_17/i0_3 ), .A3(\SB2_1_17/i0_0 ), .ZN(
        \SB2_1_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_17/Component_Function_0/N2  ( .A1(\SB2_1_17/i0[8] ), .A2(
        \SB2_1_17/i0[7] ), .A3(\SB2_1_17/i0[6] ), .ZN(
        \SB2_1_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_17/Component_Function_0/N1  ( .A1(\SB2_1_17/i0[10] ), .A2(
        \SB2_1_17/i0[9] ), .ZN(\SB2_1_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_1/N4  ( .A1(\SB2_1_17/i1_7 ), .A2(
        \SB2_1_17/i0[8] ), .A3(\SB2_1_17/i0_4 ), .ZN(
        \SB2_1_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_17/Component_Function_1/N2  ( .A1(\SB2_1_17/i0_3 ), .A2(
        \SB2_1_17/i1_7 ), .A3(\SB2_1_17/i0[8] ), .ZN(
        \SB2_1_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_18/Component_Function_0/N1  ( .A1(\SB2_1_18/i0[10] ), .A2(
        \SB2_1_18/i0[9] ), .ZN(\SB2_1_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_18/Component_Function_1/N1  ( .A1(\SB2_1_18/i0_3 ), .A2(
        \SB2_1_18/i1[9] ), .ZN(\SB2_1_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_19/Component_Function_0/N3  ( .A1(\SB2_1_19/i0[10] ), .A2(
        \SB2_1_19/i0_4 ), .A3(\SB2_1_19/i0_3 ), .ZN(
        \SB2_1_19/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_20/Component_Function_0/N1  ( .A1(\SB2_1_20/i0[10] ), .A2(
        \SB2_1_20/i0[9] ), .ZN(\SB2_1_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_20/Component_Function_1/N1  ( .A1(\SB2_1_20/i0_3 ), .A2(
        \SB2_1_20/i1[9] ), .ZN(\SB2_1_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_21/Component_Function_0/N2  ( .A1(\SB2_1_21/i0[8] ), .A2(
        \SB2_1_21/i0[7] ), .A3(\SB2_1_21/i0[6] ), .ZN(
        \SB2_1_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_21/Component_Function_1/N1  ( .A1(\SB2_1_21/i0_3 ), .A2(
        \SB2_1_21/i1[9] ), .ZN(\SB2_1_21/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_21/Component_Function_5/N1  ( .A1(\SB2_1_21/i0_0 ), .A2(
        \SB2_1_21/i3[0] ), .ZN(\SB2_1_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_0/N3  ( .A1(\SB2_1_22/i0[10] ), .A2(
        \SB2_1_22/i0_4 ), .A3(\SB2_1_22/i0_3 ), .ZN(
        \SB2_1_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_22/Component_Function_0/N2  ( .A1(n6283), .A2(
        \SB2_1_22/i0[7] ), .A3(\SB2_1_22/i0[6] ), .ZN(
        \SB2_1_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_22/Component_Function_0/N1  ( .A1(\SB2_1_22/i0[10] ), .A2(
        \SB2_1_22/i0[9] ), .ZN(\SB2_1_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_1/N2  ( .A1(\SB2_1_22/i0_3 ), .A2(
        \SB2_1_22/i1_7 ), .A3(n6283), .ZN(
        \SB2_1_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_22/Component_Function_1/N1  ( .A1(\SB2_1_22/i0_3 ), .A2(
        \SB2_1_22/i1[9] ), .ZN(\SB2_1_22/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_22/Component_Function_5/N1  ( .A1(\SB2_1_22/i0_0 ), .A2(
        \SB2_1_22/i3[0] ), .ZN(\SB2_1_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_0/N2  ( .A1(\SB2_1_23/i0[8] ), .A2(
        \SB2_1_23/i0[7] ), .A3(\SB2_1_23/i0[6] ), .ZN(
        \SB2_1_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_23/Component_Function_0/N1  ( .A1(\SB2_1_23/i0[10] ), .A2(
        \SB2_1_23/i0[9] ), .ZN(\SB2_1_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_24/Component_Function_0/N2  ( .A1(\SB2_1_24/i0[8] ), .A2(
        \SB2_1_24/i0[7] ), .A3(\SB2_1_24/i0[6] ), .ZN(
        \SB2_1_24/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_24/Component_Function_1/N3  ( .A1(\SB2_1_24/i1_5 ), .A2(
        \SB2_1_24/i0[6] ), .A3(\SB2_1_24/i0[9] ), .ZN(
        \SB2_1_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_25/Component_Function_0/N2  ( .A1(n3995), .A2(
        \SB2_1_25/i0[7] ), .A3(\SB2_1_25/i0[6] ), .ZN(
        \SB2_1_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_25/Component_Function_1/N2  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB2_1_25/i1_7 ), .A3(n3995), .ZN(
        \SB2_1_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_25/Component_Function_1/N1  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB2_1_25/i1[9] ), .ZN(\SB2_1_25/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_25/Component_Function_5/N1  ( .A1(\SB2_1_25/i0_0 ), .A2(
        \SB2_1_25/i3[0] ), .ZN(\SB2_1_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_0/N2  ( .A1(\SB2_1_26/i0[8] ), .A2(
        \SB2_1_26/i0[7] ), .A3(\SB2_1_26/i0[6] ), .ZN(
        \SB2_1_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_27/Component_Function_5/N1  ( .A1(\RI3[1][26] ), .A2(
        \SB2_1_27/i3[0] ), .ZN(\SB2_1_27/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_28/Component_Function_0/N1  ( .A1(\SB2_1_28/i0[10] ), .A2(
        \SB2_1_28/i0[9] ), .ZN(\SB2_1_28/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_28/Component_Function_1/N1  ( .A1(\SB2_1_28/i0_3 ), .A2(
        \SB2_1_28/i1[9] ), .ZN(\SB2_1_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_0/N4  ( .A1(n6612), .A2(
        \SB2_1_29/i0_3 ), .A3(\SB2_1_29/i0_0 ), .ZN(
        \SB2_1_29/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_29/Component_Function_0/N1  ( .A1(\SB2_1_29/i0[10] ), .A2(
        \SB2_1_29/i0[9] ), .ZN(\SB2_1_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_1/N4  ( .A1(\SB2_1_29/i1_7 ), .A2(
        \SB2_1_29/i0[8] ), .A3(\SB2_1_29/i0_4 ), .ZN(
        \SB2_1_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_29/Component_Function_1/N3  ( .A1(\SB2_1_29/i1_5 ), .A2(
        \SB2_1_29/i0[6] ), .A3(\SB2_1_29/i0[9] ), .ZN(
        \SB2_1_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_29/Component_Function_1/N2  ( .A1(\SB2_1_29/i0_3 ), .A2(
        \SB2_1_29/i1_7 ), .A3(\SB2_1_29/i0[8] ), .ZN(
        \SB2_1_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_29/Component_Function_1/N1  ( .A1(\SB2_1_29/i0_3 ), .A2(
        \SB2_1_29/i1[9] ), .ZN(\SB2_1_29/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_30/Component_Function_0/N1  ( .A1(\SB2_1_30/i0[10] ), .A2(
        \SB2_1_30/i0[9] ), .ZN(\SB2_1_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_1/N2  ( .A1(\SB2_1_30/i0_3 ), .A2(
        \SB2_1_30/i1_7 ), .A3(\SB2_1_30/i0[8] ), .ZN(
        \SB2_1_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_31/Component_Function_1/N2  ( .A1(\SB2_1_31/i0_3 ), .A2(
        \SB2_1_31/i1_7 ), .A3(\SB2_1_31/i0[8] ), .ZN(
        \SB2_1_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_31/Component_Function_1/N1  ( .A1(\SB2_1_31/i0_3 ), .A2(
        \SB2_1_31/i1[9] ), .ZN(\SB2_1_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_0/N3  ( .A1(\SB1_2_0/i0[10] ), .A2(
        \SB1_2_0/i0_4 ), .A3(\RI1[2][191] ), .ZN(
        \SB1_2_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_0/Component_Function_0/N2  ( .A1(\SB1_2_0/i0[8] ), .A2(
        \SB1_2_0/i0[7] ), .A3(\SB1_2_0/i0[6] ), .ZN(
        \SB1_2_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_0/Component_Function_0/N1  ( .A1(\SB1_2_0/i0[10] ), .A2(
        \SB1_2_0/i0[9] ), .ZN(\SB1_2_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_0/N3  ( .A1(\SB1_2_1/i0[10] ), .A2(
        \SB1_2_1/i0_4 ), .A3(\SB1_2_1/i0_3 ), .ZN(
        \SB1_2_1/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_1/Component_Function_0/N1  ( .A1(\SB1_2_1/i0[10] ), .A2(
        \SB1_2_1/i0[9] ), .ZN(\SB1_2_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_1/N2  ( .A1(\SB1_2_1/i0_3 ), .A2(
        \SB1_2_1/i1_7 ), .A3(\SB1_2_1/i0[8] ), .ZN(
        \SB1_2_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_1/Component_Function_1/N1  ( .A1(\SB1_2_1/i0_3 ), .A2(
        \SB1_2_1/i1[9] ), .ZN(\SB1_2_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_2/Component_Function_0/N2  ( .A1(\SB1_2_2/i0[8] ), .A2(
        \SB1_2_2/i0[7] ), .A3(\SB1_2_2/i0[6] ), .ZN(
        \SB1_2_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_2/Component_Function_0/N1  ( .A1(\SB1_2_2/i0[10] ), .A2(
        \SB1_2_2/i0[9] ), .ZN(\SB1_2_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_2/Component_Function_1/N4  ( .A1(\SB1_2_2/i1_7 ), .A2(
        \SB1_2_2/i0[8] ), .A3(\SB1_2_2/i0_4 ), .ZN(
        \SB1_2_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_1/N2  ( .A1(\SB1_2_2/i0_3 ), .A2(
        \SB1_2_2/i1_7 ), .A3(\SB1_2_2/i0[8] ), .ZN(
        \SB1_2_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_2/Component_Function_1/N1  ( .A1(\SB1_2_2/i0_3 ), .A2(
        \SB1_2_2/i1[9] ), .ZN(\SB1_2_2/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_2/Component_Function_5/N1  ( .A1(\SB1_2_2/i0_0 ), .A2(
        \SB1_2_2/i3[0] ), .ZN(\SB1_2_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_3/Component_Function_0/N2  ( .A1(\SB1_2_3/i0[8] ), .A2(
        \SB1_2_3/i0[7] ), .A3(\SB1_2_3/i0[6] ), .ZN(
        \SB1_2_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_3/Component_Function_0/N1  ( .A1(\SB1_2_3/i0[10] ), .A2(
        \SB1_2_3/i0[9] ), .ZN(\SB1_2_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_3/Component_Function_1/N2  ( .A1(\SB1_2_3/i0_3 ), .A2(
        \SB1_2_3/i1_7 ), .A3(\SB1_2_3/i0[8] ), .ZN(
        \SB1_2_3/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_4/Component_Function_0/N2  ( .A1(\SB1_2_4/i0[8] ), .A2(
        \SB1_2_4/i0[7] ), .A3(\SB1_2_4/i0[6] ), .ZN(
        \SB1_2_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_4/Component_Function_1/N1  ( .A1(\SB1_2_4/i0_3 ), .A2(
        \SB1_2_4/i1[9] ), .ZN(\SB1_2_4/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_5/Component_Function_0/N1  ( .A1(\SB1_2_5/i0[10] ), .A2(
        \SB1_2_5/i0[9] ), .ZN(\SB1_2_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_0/N3  ( .A1(\SB1_2_6/i0[10] ), .A2(
        \SB1_2_6/i0_4 ), .A3(\SB1_2_6/i0_3 ), .ZN(
        \SB1_2_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_6/Component_Function_0/N2  ( .A1(\SB1_2_6/i0[8] ), .A2(
        \SB1_2_6/i0[7] ), .A3(\SB1_2_6/i0[6] ), .ZN(
        \SB1_2_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_6/Component_Function_0/N1  ( .A1(\SB1_2_6/i0[10] ), .A2(
        \SB1_2_6/i0[9] ), .ZN(\SB1_2_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_1/N2  ( .A1(\SB1_2_6/i0_3 ), .A2(
        \SB1_2_6/i1_7 ), .A3(\SB1_2_6/i0[8] ), .ZN(
        \SB1_2_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_6/Component_Function_1/N1  ( .A1(\SB1_2_6/i0_3 ), .A2(
        \SB1_2_6/i1[9] ), .ZN(\SB1_2_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_0/N2  ( .A1(n3184), .A2(\SB1_2_7/i0[7] ), .A3(\SB1_2_7/i0[6] ), .ZN(\SB1_2_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_7/Component_Function_0/N1  ( .A1(\SB1_2_7/i0[10] ), .A2(
        \SB1_2_7/i0[9] ), .ZN(\SB1_2_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_1/N4  ( .A1(\SB1_2_7/i1_7 ), .A2(n3184), 
        .A3(\SB1_2_7/i0_4 ), .ZN(\SB1_2_7/Component_Function_1/NAND4_in[3] )
         );
  NAND2_X1 \SB1_2_7/Component_Function_1/N1  ( .A1(\RI1[2][149] ), .A2(
        \SB1_2_7/i1[9] ), .ZN(\SB1_2_7/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_8/Component_Function_0/N1  ( .A1(\SB1_2_8/i0[10] ), .A2(
        \SB1_2_8/i0[9] ), .ZN(\SB1_2_8/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_8/Component_Function_1/N1  ( .A1(\SB1_2_8/i0_3 ), .A2(
        \SB1_2_8/i1[9] ), .ZN(\SB1_2_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_0/N2  ( .A1(\SB1_2_9/i0[8] ), .A2(
        \SB1_2_9/i0[7] ), .A3(\SB1_2_9/i0[6] ), .ZN(
        \SB1_2_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_9/Component_Function_0/N1  ( .A1(\SB1_2_9/i0[10] ), .A2(
        \SB1_2_9/i0[9] ), .ZN(\SB1_2_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_1/N2  ( .A1(\SB1_2_9/i0_3 ), .A2(
        \SB1_2_9/i1_7 ), .A3(\SB1_2_9/i0[8] ), .ZN(
        \SB1_2_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_9/Component_Function_1/N1  ( .A1(\SB1_2_9/i0_3 ), .A2(
        \SB1_2_9/i1[9] ), .ZN(\SB1_2_9/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_10/Component_Function_0/N1  ( .A1(\SB1_2_10/i0[10] ), .A2(
        \SB1_2_10/i0[9] ), .ZN(\SB1_2_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_10/Component_Function_1/N1  ( .A1(\SB1_2_10/i0_3 ), .A2(
        \SB1_2_10/i1[9] ), .ZN(\SB1_2_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_0/N3  ( .A1(\SB1_2_11/i0[10] ), .A2(
        \SB1_2_11/i0_4 ), .A3(\SB1_2_11/i0_3 ), .ZN(
        \SB1_2_11/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_11/Component_Function_0/N1  ( .A1(\SB1_2_11/i0[10] ), .A2(
        \SB1_2_11/i0[9] ), .ZN(\SB1_2_11/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_11/Component_Function_5/N1  ( .A1(\SB1_2_11/i0_0 ), .A2(
        \SB1_2_11/i3[0] ), .ZN(\SB1_2_11/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_12/Component_Function_0/N1  ( .A1(\SB1_2_12/i0[10] ), .A2(
        \MC_ARK_ARC_1_1/buf_output[114] ), .ZN(
        \SB1_2_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_12/Component_Function_1/N4  ( .A1(\SB1_2_12/i1_7 ), .A2(
        \SB1_2_12/i0[8] ), .A3(\SB1_2_12/i0_4 ), .ZN(
        \SB1_2_12/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_12/Component_Function_5/N1  ( .A1(\RI1[2][116] ), .A2(
        \SB1_2_12/i3[0] ), .ZN(\SB1_2_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_13/Component_Function_0/N4  ( .A1(\SB1_2_13/i0[7] ), .A2(
        \SB1_2_13/i0_3 ), .A3(\SB1_2_13/i0_0 ), .ZN(
        \SB1_2_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_13/Component_Function_0/N3  ( .A1(\SB1_2_13/i0[10] ), .A2(
        \SB1_2_13/i0_4 ), .A3(\SB1_2_13/i0_3 ), .ZN(
        \SB1_2_13/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_13/Component_Function_0/N1  ( .A1(\SB1_2_13/i0[10] ), .A2(
        \SB1_2_13/i0[9] ), .ZN(\SB1_2_13/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_13/Component_Function_1/N1  ( .A1(\SB1_2_13/i0_3 ), .A2(
        \SB1_2_13/i1[9] ), .ZN(\SB1_2_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_0/N2  ( .A1(\SB1_2_14/i0[8] ), .A2(
        \SB1_2_14/i0[7] ), .A3(\SB1_2_14/i0[6] ), .ZN(
        \SB1_2_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_14/Component_Function_0/N1  ( .A1(\SB1_2_14/i0[10] ), .A2(
        \SB1_2_14/i0[9] ), .ZN(\SB1_2_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_1/N2  ( .A1(\RI1[2][107] ), .A2(
        \SB1_2_14/i1_7 ), .A3(\SB1_2_14/i0[8] ), .ZN(
        \SB1_2_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_15/Component_Function_0/N3  ( .A1(\SB1_2_15/i0[10] ), .A2(
        \SB1_2_15/i0_4 ), .A3(\RI1[2][101] ), .ZN(
        \SB1_2_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_15/Component_Function_0/N2  ( .A1(\SB1_2_15/i0[8] ), .A2(
        \SB1_2_15/i0[7] ), .A3(\SB1_2_15/i0[6] ), .ZN(
        \SB1_2_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_15/Component_Function_0/N1  ( .A1(\SB1_2_15/i0[10] ), .A2(
        \SB1_2_15/i0[9] ), .ZN(\SB1_2_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_15/Component_Function_1/N4  ( .A1(\SB1_2_15/i1_7 ), .A2(
        \SB1_2_15/i0[8] ), .A3(\SB1_2_15/i0_4 ), .ZN(
        \SB1_2_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_16/Component_Function_0/N3  ( .A1(\SB1_2_16/i0[10] ), .A2(
        \SB1_2_16/i0_4 ), .A3(\SB1_2_16/i0_3 ), .ZN(
        \SB1_2_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_16/Component_Function_0/N2  ( .A1(\SB1_2_16/i0[8] ), .A2(
        \SB1_2_16/i0[7] ), .A3(\SB1_2_16/i0[6] ), .ZN(
        \SB1_2_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_16/Component_Function_0/N1  ( .A1(\SB1_2_16/i0[10] ), .A2(
        \SB1_2_16/i0[9] ), .ZN(\SB1_2_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_16/Component_Function_1/N3  ( .A1(\SB1_2_16/i1_5 ), .A2(
        \SB1_2_16/i0[6] ), .A3(\SB1_2_16/i0[9] ), .ZN(
        \SB1_2_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_16/Component_Function_1/N2  ( .A1(\SB1_2_16/i0_3 ), .A2(
        \SB1_2_16/i1_7 ), .A3(\SB1_2_16/i0[8] ), .ZN(
        \SB1_2_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_17/Component_Function_0/N1  ( .A1(\SB1_2_17/i0[10] ), .A2(
        \SB1_2_17/i0[9] ), .ZN(\SB1_2_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_17/Component_Function_1/N2  ( .A1(\SB1_2_17/i0_3 ), .A2(
        \SB1_2_17/i1_7 ), .A3(\SB1_2_17/i0[8] ), .ZN(
        \SB1_2_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_17/Component_Function_1/N1  ( .A1(\SB1_2_17/i0_3 ), .A2(
        \SB1_2_17/i1[9] ), .ZN(\SB1_2_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_0/N3  ( .A1(\SB1_2_18/i0[10] ), .A2(
        \SB1_2_18/i0_4 ), .A3(\SB1_2_18/i0_3 ), .ZN(
        \SB1_2_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_18/Component_Function_0/N2  ( .A1(\SB1_2_18/i0[8] ), .A2(
        \SB1_2_18/i0[7] ), .A3(\SB1_2_18/i0[6] ), .ZN(
        \SB1_2_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_18/Component_Function_0/N1  ( .A1(\SB1_2_18/i0[10] ), .A2(
        \SB1_2_18/i0[9] ), .ZN(\SB1_2_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_18/Component_Function_1/N1  ( .A1(\SB1_2_18/i0_3 ), .A2(
        \SB1_2_18/i1[9] ), .ZN(\SB1_2_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_0/N4  ( .A1(\SB1_2_19/i0[7] ), .A2(
        \SB1_2_19/i0_3 ), .A3(\SB1_2_19/i0_0 ), .ZN(
        \SB1_2_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_0/N3  ( .A1(\SB1_2_19/i0[10] ), .A2(
        \SB1_2_19/i0_4 ), .A3(\SB1_2_19/i0_3 ), .ZN(
        \SB1_2_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_19/Component_Function_0/N2  ( .A1(\SB1_2_19/i0[8] ), .A2(
        \SB1_2_19/i0[7] ), .A3(\SB1_2_19/i0[6] ), .ZN(
        \SB1_2_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_19/Component_Function_0/N1  ( .A1(\SB1_2_19/i0[10] ), .A2(
        \SB1_2_19/i0[9] ), .ZN(\SB1_2_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_1/N4  ( .A1(\SB1_2_19/i1_7 ), .A2(
        \SB1_2_19/i0[8] ), .A3(\SB1_2_19/i0_4 ), .ZN(
        \SB1_2_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_1/N3  ( .A1(\SB1_2_19/i1_5 ), .A2(
        \SB1_2_19/i0[6] ), .A3(\SB1_2_19/i0[9] ), .ZN(
        \SB1_2_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_20/Component_Function_0/N4  ( .A1(\SB1_2_20/i0[7] ), .A2(
        \SB1_2_20/i0_3 ), .A3(\SB1_2_20/i0_0 ), .ZN(
        \SB1_2_20/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_20/Component_Function_0/N1  ( .A1(\SB1_2_20/i0[10] ), .A2(
        \SB1_2_20/i0[9] ), .ZN(\SB1_2_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_1/N4  ( .A1(\SB1_2_20/i1_7 ), .A2(
        \SB1_2_20/i0[8] ), .A3(\SB1_2_20/i0_4 ), .ZN(
        \SB1_2_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_20/Component_Function_1/N2  ( .A1(\SB1_2_20/i0_3 ), .A2(
        \SB1_2_20/i1_7 ), .A3(\SB1_2_20/i0[8] ), .ZN(
        \SB1_2_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_20/Component_Function_1/N1  ( .A1(\SB1_2_20/i0_3 ), .A2(
        \SB1_2_20/i1[9] ), .ZN(\SB1_2_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_1/N2  ( .A1(\SB1_2_21/i0_3 ), .A2(
        \SB1_2_21/i1_7 ), .A3(\SB1_2_21/i0[8] ), .ZN(
        \SB1_2_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_21/Component_Function_1/N1  ( .A1(\SB1_2_21/i0_3 ), .A2(
        \SB1_2_21/i1[9] ), .ZN(\SB1_2_21/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_22/Component_Function_5/N1  ( .A1(\SB1_2_22/i0_0 ), .A2(
        \SB1_2_22/i3[0] ), .ZN(\SB1_2_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_0/N3  ( .A1(\SB1_2_23/i0[10] ), .A2(
        \SB1_2_23/i0_4 ), .A3(\SB1_2_23/i0_3 ), .ZN(
        \SB1_2_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_23/Component_Function_0/N2  ( .A1(\SB1_2_23/i0[8] ), .A2(
        \SB1_2_23/i0[7] ), .A3(\SB1_2_23/i0[6] ), .ZN(
        \SB1_2_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_23/Component_Function_0/N1  ( .A1(\SB1_2_23/i0[10] ), .A2(
        \SB1_2_23/i0[9] ), .ZN(\SB1_2_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_1/N3  ( .A1(\SB1_2_23/i1_5 ), .A2(
        \SB1_2_23/i0[6] ), .A3(\SB1_2_23/i0[9] ), .ZN(
        \SB1_2_23/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_23/Component_Function_1/N1  ( .A1(\SB1_2_23/i0_3 ), .A2(
        \SB1_2_23/i1[9] ), .ZN(\SB1_2_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_0/N3  ( .A1(\SB1_2_24/i0[10] ), .A2(
        \SB1_2_24/i0_4 ), .A3(\SB1_2_24/i0_3 ), .ZN(
        \SB1_2_24/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_24/Component_Function_1/N1  ( .A1(\SB1_2_24/i0_3 ), .A2(
        \SB1_2_24/i1[9] ), .ZN(\SB1_2_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_25/Component_Function_0/N4  ( .A1(\SB1_2_25/i0[7] ), .A2(
        \SB1_2_25/i0_3 ), .A3(\SB1_2_25/i0_0 ), .ZN(
        \SB1_2_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_0/N3  ( .A1(\SB1_2_25/i0[10] ), .A2(
        \SB1_2_25/i0_4 ), .A3(\SB1_2_25/i0_3 ), .ZN(
        \SB1_2_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_25/Component_Function_0/N2  ( .A1(\SB1_2_25/i0[8] ), .A2(
        \SB1_2_25/i0[7] ), .A3(\SB1_2_25/i0[6] ), .ZN(
        \SB1_2_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_25/Component_Function_0/N1  ( .A1(\SB1_2_25/i0[10] ), .A2(
        \SB1_2_25/i0[9] ), .ZN(\SB1_2_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_25/Component_Function_1/N4  ( .A1(\SB1_2_25/i1_7 ), .A2(
        \SB1_2_25/i0[8] ), .A3(\SB1_2_25/i0_4 ), .ZN(
        \SB1_2_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_1/N3  ( .A1(\SB1_2_25/i1_5 ), .A2(
        \SB1_2_25/i0[6] ), .A3(\SB1_2_25/i0[9] ), .ZN(
        \SB1_2_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_25/Component_Function_1/N2  ( .A1(\SB1_2_25/i0_3 ), .A2(
        \SB1_2_25/i1_7 ), .A3(\SB1_2_25/i0[8] ), .ZN(
        \SB1_2_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_26/Component_Function_1/N1  ( .A1(\SB1_2_26/i0_3 ), .A2(
        \SB1_2_26/i1[9] ), .ZN(\SB1_2_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_0/N3  ( .A1(\SB1_2_27/i0[10] ), .A2(
        \SB1_2_27/i0_4 ), .A3(\SB1_2_27/i0_3 ), .ZN(
        \SB1_2_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_27/Component_Function_0/N2  ( .A1(\SB1_2_27/i0[8] ), .A2(
        \SB1_2_27/i0[7] ), .A3(\SB1_2_27/i0[6] ), .ZN(
        \SB1_2_27/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_27/Component_Function_1/N4  ( .A1(\SB1_2_27/i1_7 ), .A2(
        \SB1_2_27/i0[8] ), .A3(\SB1_2_27/i0_4 ), .ZN(
        \SB1_2_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_27/Component_Function_1/N2  ( .A1(\SB1_2_27/i0_3 ), .A2(
        \SB1_2_27/i1_7 ), .A3(\SB1_2_27/i0[8] ), .ZN(
        \SB1_2_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_27/Component_Function_1/N1  ( .A1(\SB1_2_27/i0_3 ), .A2(
        \SB1_2_27/i1[9] ), .ZN(\SB1_2_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_0/N3  ( .A1(\SB1_2_28/i0[10] ), .A2(
        \SB1_2_28/i0_4 ), .A3(\SB1_2_28/i0_3 ), .ZN(
        \SB1_2_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_28/Component_Function_0/N2  ( .A1(\SB1_2_28/i0[8] ), .A2(
        \SB1_2_28/i0[7] ), .A3(\SB1_2_28/i0[6] ), .ZN(
        \SB1_2_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_28/Component_Function_0/N1  ( .A1(\SB1_2_28/i0[10] ), .A2(
        \SB1_2_28/i0[9] ), .ZN(\SB1_2_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_1/N3  ( .A1(\SB1_2_28/i1_5 ), .A2(
        \SB1_2_28/i0[6] ), .A3(\SB1_2_28/i0[9] ), .ZN(
        \SB1_2_28/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_29/Component_Function_1/N1  ( .A1(\RI1[2][17] ), .A2(
        \SB1_2_29/i1[9] ), .ZN(\SB1_2_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_0/N3  ( .A1(\SB1_2_30/i0[10] ), .A2(
        \SB1_2_30/i0_4 ), .A3(\SB1_2_30/i0_3 ), .ZN(
        \SB1_2_30/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_30/Component_Function_0/N1  ( .A1(\SB1_2_30/i0[10] ), .A2(
        \SB1_2_30/i0[9] ), .ZN(\SB1_2_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_1/N2  ( .A1(\SB1_2_30/i0_3 ), .A2(
        \SB1_2_30/i1_7 ), .A3(\SB1_2_30/i0[8] ), .ZN(
        \SB1_2_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_30/Component_Function_1/N1  ( .A1(\SB1_2_30/i0_3 ), .A2(
        \SB1_2_30/i1[9] ), .ZN(\SB1_2_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_0/N2  ( .A1(\SB1_2_31/i0[8] ), .A2(
        \SB1_2_31/i0[7] ), .A3(\SB1_2_31/i0[6] ), .ZN(
        \SB1_2_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_31/Component_Function_0/N1  ( .A1(\SB1_2_31/i0[10] ), .A2(
        \SB1_2_31/i0[9] ), .ZN(\SB1_2_31/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_0/Component_Function_0/N1  ( .A1(\SB2_2_0/i0[10] ), .A2(
        \SB2_2_0/i0[9] ), .ZN(\SB2_2_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_1/Component_Function_0/N2  ( .A1(\SB2_2_1/i0[8] ), .A2(n2748), .A3(\SB2_2_1/i0[6] ), .ZN(\SB2_2_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_1/Component_Function_0/N1  ( .A1(\SB2_2_1/i0[10] ), .A2(
        \SB2_2_1/i0[9] ), .ZN(\SB2_2_1/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_2/Component_Function_0/N1  ( .A1(\SB2_2_2/i0[10] ), .A2(
        \SB2_2_2/i0[9] ), .ZN(\SB2_2_2/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_2/Component_Function_1/N1  ( .A1(\SB2_2_2/i0_3 ), .A2(n6267), 
        .ZN(\SB2_2_2/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_3/Component_Function_0/N1  ( .A1(\SB2_2_3/i0[10] ), .A2(
        \SB2_2_3/i0[9] ), .ZN(\SB2_2_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_3/Component_Function_1/N2  ( .A1(\SB2_2_3/i0_3 ), .A2(
        \SB2_2_3/i1_7 ), .A3(n3991), .ZN(
        \SB2_2_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_4/Component_Function_0/N1  ( .A1(\SB2_2_4/i0[10] ), .A2(
        \SB2_2_4/i0[9] ), .ZN(\SB2_2_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_4/Component_Function_1/N2  ( .A1(\SB2_2_4/i0_3 ), .A2(
        \SB2_2_4/i1_7 ), .A3(\SB2_2_4/i0[8] ), .ZN(
        \SB2_2_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_5/Component_Function_1/N1  ( .A1(\SB2_2_5/i0_3 ), .A2(
        \SB2_2_5/i1[9] ), .ZN(\SB2_2_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_0/N2  ( .A1(\SB2_2_6/i0[8] ), .A2(
        \SB2_2_6/i0[7] ), .A3(\SB2_2_6/i0[6] ), .ZN(
        \SB2_2_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_6/Component_Function_0/N1  ( .A1(\SB2_2_6/i0[10] ), .A2(
        \SB2_2_6/i0[9] ), .ZN(\SB2_2_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_1/N2  ( .A1(\SB2_2_6/i0_3 ), .A2(
        \SB2_2_6/i1_7 ), .A3(\SB2_2_6/i0[8] ), .ZN(
        \SB2_2_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_7/Component_Function_1/N1  ( .A1(\SB2_2_7/i0_3 ), .A2(
        \SB2_2_7/i1[9] ), .ZN(\SB2_2_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_8/Component_Function_0/N3  ( .A1(\SB2_2_8/i0[10] ), .A2(
        \SB2_2_8/i0_4 ), .A3(\SB2_2_8/i0_3 ), .ZN(
        \SB2_2_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_8/Component_Function_0/N2  ( .A1(\SB2_2_8/i0[8] ), .A2(
        \SB2_2_8/i0[7] ), .A3(\SB2_2_8/i0[6] ), .ZN(
        \SB2_2_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_8/Component_Function_0/N1  ( .A1(\SB2_2_8/i0[10] ), .A2(
        \SB2_2_8/i0[9] ), .ZN(\SB2_2_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_8/Component_Function_1/N2  ( .A1(\SB2_2_8/i0_3 ), .A2(
        \SB2_2_8/i1_7 ), .A3(\SB2_2_8/i0[8] ), .ZN(
        \SB2_2_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_8/Component_Function_1/N1  ( .A1(\SB2_2_8/i0_3 ), .A2(
        \SB2_2_8/i1[9] ), .ZN(\SB2_2_8/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_9/Component_Function_0/N1  ( .A1(\SB2_2_9/i0[10] ), .A2(
        \SB2_2_9/i0[9] ), .ZN(\SB2_2_9/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_10/Component_Function_0/N1  ( .A1(\SB2_2_10/i0[10] ), .A2(
        \SB2_2_10/i0[9] ), .ZN(\SB2_2_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_10/Component_Function_1/N1  ( .A1(\SB2_2_10/i0_3 ), .A2(
        \SB2_2_10/i1[9] ), .ZN(\SB2_2_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_11/Component_Function_0/N2  ( .A1(\SB2_2_11/i0[8] ), .A2(
        \SB2_2_11/i0[7] ), .A3(\SB2_2_11/i0[6] ), .ZN(
        \SB2_2_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_11/Component_Function_0/N1  ( .A1(\SB2_2_11/i0[10] ), .A2(
        \SB2_2_11/i0[9] ), .ZN(\SB2_2_11/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_11/Component_Function_1/N1  ( .A1(\SB2_2_11/i0_3 ), .A2(
        \SB2_2_11/i1[9] ), .ZN(\SB2_2_11/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_12/Component_Function_0/N1  ( .A1(\SB2_2_12/i0[10] ), .A2(
        \SB2_2_12/i0[9] ), .ZN(\SB2_2_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_12/Component_Function_1/N3  ( .A1(\SB2_2_12/i1_5 ), .A2(
        \SB2_2_12/i0[6] ), .A3(\SB2_2_12/i0[9] ), .ZN(
        \SB2_2_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_13/Component_Function_0/N2  ( .A1(\SB2_2_13/i0[8] ), .A2(
        \SB2_2_13/i0[7] ), .A3(\SB2_2_13/i0[6] ), .ZN(
        \SB2_2_13/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_13/Component_Function_1/N4  ( .A1(\SB2_2_13/i1_7 ), .A2(
        \SB2_2_13/i0[8] ), .A3(\SB2_2_13/i0_4 ), .ZN(
        \SB2_2_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_13/Component_Function_1/N2  ( .A1(\SB2_2_13/i0_3 ), .A2(
        \SB2_2_13/i1_7 ), .A3(\SB2_2_13/i0[8] ), .ZN(
        \SB2_2_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_14/Component_Function_0/N2  ( .A1(\SB2_2_14/i0[8] ), .A2(
        \SB2_2_14/i0[7] ), .A3(\SB2_2_14/i0[6] ), .ZN(
        \SB2_2_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_14/Component_Function_1/N1  ( .A1(\SB2_2_14/i0_3 ), .A2(
        \SB2_2_14/i1[9] ), .ZN(\SB2_2_14/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_15/Component_Function_0/N1  ( .A1(\SB2_2_15/i0[10] ), .A2(
        \SB2_2_15/i0[9] ), .ZN(\SB2_2_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_0/N2  ( .A1(\SB2_2_16/i0[8] ), .A2(
        \SB2_2_16/i0[7] ), .A3(\SB2_2_16/i0[6] ), .ZN(
        \SB2_2_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_17/Component_Function_5/N1  ( .A1(\SB2_2_17/i0_0 ), .A2(
        \SB2_2_17/i3[0] ), .ZN(\SB2_2_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_18/Component_Function_0/N4  ( .A1(n1102), .A2(
        \SB2_2_18/i0_3 ), .A3(\SB2_2_18/i0_0 ), .ZN(
        \SB2_2_18/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_18/Component_Function_0/N1  ( .A1(\SB2_2_18/i0[10] ), .A2(
        \SB2_2_18/i0[9] ), .ZN(\SB2_2_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_0/N3  ( .A1(\SB2_2_19/i0[10] ), .A2(
        \SB2_2_19/i0_4 ), .A3(\SB2_2_19/i0_3 ), .ZN(
        \SB2_2_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_19/Component_Function_0/N2  ( .A1(\SB2_2_19/i0[8] ), .A2(
        \SB2_2_19/i0[7] ), .A3(\SB2_2_19/i0[6] ), .ZN(
        \SB2_2_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_19/Component_Function_0/N1  ( .A1(\SB2_2_19/i0[10] ), .A2(
        \SB2_2_19/i0[9] ), .ZN(\SB2_2_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_1/N2  ( .A1(\SB2_2_19/i0_3 ), .A2(
        \SB2_2_19/i1_7 ), .A3(\SB2_2_19/i0[8] ), .ZN(
        \SB2_2_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_19/Component_Function_1/N1  ( .A1(\SB2_2_19/i0_3 ), .A2(
        \SB2_2_19/i1[9] ), .ZN(\SB2_2_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_19/Component_Function_5/N1  ( .A1(\SB2_2_19/i0_0 ), .A2(
        \SB2_2_19/i3[0] ), .ZN(\SB2_2_19/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_20/Component_Function_0/N1  ( .A1(\SB2_2_20/i0[10] ), .A2(
        \SB2_2_20/i0[9] ), .ZN(\SB2_2_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_21/Component_Function_0/N2  ( .A1(\SB2_2_21/i0[8] ), .A2(
        n7225), .A3(\SB2_2_21/i0[6] ), .ZN(
        \SB2_2_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_21/Component_Function_1/N3  ( .A1(\SB2_2_21/i1_5 ), .A2(
        \SB2_2_21/i0[6] ), .A3(\SB1_2_26/buf_output[0] ), .ZN(
        \SB2_2_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_22/Component_Function_1/N4  ( .A1(\SB2_2_22/i1_7 ), .A2(
        \SB2_2_22/i0[8] ), .A3(\SB2_2_22/i0_4 ), .ZN(
        \SB2_2_22/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_22/Component_Function_1/N1  ( .A1(\SB2_2_22/i0_3 ), .A2(
        \SB2_2_22/i1[9] ), .ZN(\SB2_2_22/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_23/Component_Function_0/N1  ( .A1(\SB2_2_23/i0[10] ), .A2(
        \SB2_2_23/i0[9] ), .ZN(\SB2_2_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_23/Component_Function_1/N2  ( .A1(\SB2_2_23/i0_3 ), .A2(
        \SB2_2_23/i1_7 ), .A3(\SB2_2_23/i0[8] ), .ZN(
        \SB2_2_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_23/Component_Function_1/N1  ( .A1(\SB2_2_23/i0_3 ), .A2(
        \SB2_2_23/i1[9] ), .ZN(\SB2_2_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_24/Component_Function_0/N2  ( .A1(\SB2_2_24/i0[8] ), .A2(
        \SB2_2_24/i0[7] ), .A3(\SB2_2_24/i0[6] ), .ZN(
        \SB2_2_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_24/Component_Function_0/N1  ( .A1(\SB2_2_24/i0[10] ), .A2(
        \SB2_2_24/i0[9] ), .ZN(\SB2_2_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_24/Component_Function_1/N4  ( .A1(\SB2_2_24/i1_7 ), .A2(
        \SB2_2_24/i0[8] ), .A3(\SB2_2_24/i0_4 ), .ZN(
        \SB2_2_24/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_25/Component_Function_0/N1  ( .A1(\SB2_2_25/i0[10] ), .A2(
        \SB2_2_25/i0[9] ), .ZN(\SB2_2_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_1/N2  ( .A1(\SB2_2_25/i0_3 ), .A2(
        \SB2_2_25/i1_7 ), .A3(\SB2_2_25/i0[8] ), .ZN(
        \SB2_2_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_26/Component_Function_1/N1  ( .A1(\SB2_2_26/i0_3 ), .A2(
        \SB2_2_26/i1[9] ), .ZN(\SB2_2_26/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_27/Component_Function_5/N1  ( .A1(\SB2_2_27/i0_0 ), .A2(
        \SB2_2_27/i3[0] ), .ZN(\SB2_2_27/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_28/Component_Function_0/N1  ( .A1(\SB2_2_28/i0[10] ), .A2(
        \SB2_2_28/i0[9] ), .ZN(\SB2_2_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_28/Component_Function_1/N3  ( .A1(\SB2_2_28/i1_5 ), .A2(
        \SB2_2_28/i0[6] ), .A3(\SB2_2_28/i0[9] ), .ZN(
        \SB2_2_28/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_28/Component_Function_1/N1  ( .A1(\SB2_2_28/i0_3 ), .A2(
        \SB2_2_28/i1[9] ), .ZN(\SB2_2_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_0/N3  ( .A1(\SB2_2_29/i0[10] ), .A2(
        \SB2_2_29/i0_4 ), .A3(\SB2_2_29/i0_3 ), .ZN(
        \SB2_2_29/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_29/Component_Function_0/N1  ( .A1(\SB2_2_29/i0[10] ), .A2(
        \SB2_2_29/i0[9] ), .ZN(\SB2_2_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_1/N4  ( .A1(\SB2_2_29/i1_7 ), .A2(
        \SB2_2_29/i0[8] ), .A3(\SB2_2_29/i0_4 ), .ZN(
        \SB2_2_29/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_29/Component_Function_1/N1  ( .A1(\SB2_2_29/i0_3 ), .A2(
        \SB2_2_29/i1[9] ), .ZN(\SB2_2_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_0/N2  ( .A1(\SB2_2_30/i0[8] ), .A2(
        \SB2_2_30/i0[7] ), .A3(\SB2_2_30/i0[6] ), .ZN(
        \SB2_2_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_30/Component_Function_0/N1  ( .A1(\SB2_2_30/i0[10] ), .A2(
        \SB2_2_30/i0[9] ), .ZN(\SB2_2_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_1/N2  ( .A1(\SB2_2_30/i0_3 ), .A2(
        \SB2_2_30/i1_7 ), .A3(\SB2_2_30/i0[8] ), .ZN(
        \SB2_2_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_31/Component_Function_1/N2  ( .A1(\SB2_2_31/i0_3 ), .A2(
        \SB2_2_31/i1_7 ), .A3(\SB2_2_31/i0[8] ), .ZN(
        \SB2_2_31/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_0/Component_Function_0/N2  ( .A1(\SB1_3_0/i0[8] ), .A2(
        \SB1_3_0/i0[7] ), .A3(\SB1_3_0/i0[6] ), .ZN(
        \SB1_3_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_0/Component_Function_0/N1  ( .A1(\SB1_3_0/i0[10] ), .A2(
        \SB1_3_0/i0[9] ), .ZN(\SB1_3_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_1/N2  ( .A1(\SB1_3_0/i0_3 ), .A2(
        \SB1_3_0/i1_7 ), .A3(\SB1_3_0/i0[8] ), .ZN(
        \SB1_3_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_0/Component_Function_1/N1  ( .A1(\SB1_3_0/i0_3 ), .A2(
        \SB1_3_0/i1[9] ), .ZN(\SB1_3_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_0/N3  ( .A1(\SB1_3_1/i0[10] ), .A2(
        \SB1_3_1/i0_4 ), .A3(\SB1_3_1/i0_3 ), .ZN(
        \SB1_3_1/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_1/Component_Function_0/N1  ( .A1(\SB1_3_1/i0[10] ), .A2(
        \SB1_3_1/i0[9] ), .ZN(\SB1_3_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_0/N4  ( .A1(\SB1_3_3/i0[7] ), .A2(
        \SB1_3_3/i0_3 ), .A3(\SB1_3_3/i0_0 ), .ZN(
        \SB1_3_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_3/Component_Function_0/N3  ( .A1(\SB1_3_3/i0[10] ), .A2(
        \SB1_3_3/i0_4 ), .A3(\SB1_3_3/i0_3 ), .ZN(
        \SB1_3_3/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_3/Component_Function_0/N1  ( .A1(\SB1_3_3/i0[10] ), .A2(
        \SB1_3_3/i0[9] ), .ZN(\SB1_3_3/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_3/Component_Function_1/N1  ( .A1(\SB1_3_3/i0_3 ), .A2(
        \SB1_3_3/i1[9] ), .ZN(\SB1_3_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_4/Component_Function_0/N2  ( .A1(\SB1_3_4/i0[8] ), .A2(
        \SB1_3_4/i0[7] ), .A3(\SB1_3_4/i0[6] ), .ZN(
        \SB1_3_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_4/Component_Function_0/N1  ( .A1(\SB1_3_4/i0[10] ), .A2(
        \SB1_3_4/i0[9] ), .ZN(\SB1_3_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_4/Component_Function_1/N4  ( .A1(\SB1_3_4/i1_7 ), .A2(
        \SB1_3_4/i0[8] ), .A3(\SB1_3_4/i0_4 ), .ZN(
        \SB1_3_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_4/Component_Function_1/N3  ( .A1(\SB1_3_4/i1_5 ), .A2(
        \SB1_3_4/i0[6] ), .A3(\SB1_3_4/i0[9] ), .ZN(
        \SB1_3_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_5/Component_Function_0/N3  ( .A1(\SB1_3_5/i0[10] ), .A2(
        \SB1_3_5/i0_4 ), .A3(\SB1_3_5/i0_3 ), .ZN(
        \SB1_3_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_5/Component_Function_0/N2  ( .A1(\SB1_3_5/i0[8] ), .A2(
        \SB1_3_5/i0[7] ), .A3(\SB1_3_5/i0[6] ), .ZN(
        \SB1_3_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_5/Component_Function_0/N1  ( .A1(\SB1_3_5/i0[10] ), .A2(
        \SB1_3_5/i0[9] ), .ZN(\SB1_3_5/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_5/Component_Function_1/N1  ( .A1(\SB1_3_5/i0_3 ), .A2(
        \SB1_3_5/i1[9] ), .ZN(\SB1_3_5/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_5/Component_Function_5/N1  ( .A1(\SB1_3_5/i0_0 ), .A2(
        \SB1_3_5/i3[0] ), .ZN(\SB1_3_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_0/N2  ( .A1(\SB1_3_6/i0[8] ), .A2(
        \SB1_3_6/i0[7] ), .A3(\SB1_3_6/i0[6] ), .ZN(
        \SB1_3_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_6/Component_Function_0/N1  ( .A1(\SB1_3_6/i0[10] ), .A2(
        \SB1_3_6/i0[9] ), .ZN(\SB1_3_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_7/Component_Function_0/N3  ( .A1(\SB1_3_7/i0[10] ), .A2(
        \SB1_3_7/i0_4 ), .A3(\SB1_3_7/i0_3 ), .ZN(
        \SB1_3_7/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_7/Component_Function_0/N1  ( .A1(\SB1_3_7/i0[10] ), .A2(
        \SB1_3_7/i0[9] ), .ZN(\SB1_3_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_7/Component_Function_1/N2  ( .A1(\SB1_3_7/i0_3 ), .A2(
        \SB1_3_7/i1_7 ), .A3(\SB1_3_7/i0[8] ), .ZN(
        \SB1_3_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_7/Component_Function_1/N1  ( .A1(\SB1_3_7/i0_3 ), .A2(
        \SB1_3_7/i1[9] ), .ZN(\SB1_3_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_8/Component_Function_0/N3  ( .A1(\SB1_3_8/i0[10] ), .A2(
        \SB1_3_8/i0_4 ), .A3(\SB1_3_8/i0_3 ), .ZN(
        \SB1_3_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_8/Component_Function_0/N2  ( .A1(\SB1_3_8/i0[8] ), .A2(
        \SB1_3_8/i0[7] ), .A3(\SB1_3_8/i0[6] ), .ZN(
        \SB1_3_8/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_8/Component_Function_1/N2  ( .A1(\SB1_3_8/i0_3 ), .A2(
        \SB1_3_8/i1_7 ), .A3(\SB1_3_8/i0[8] ), .ZN(
        \SB1_3_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_8/Component_Function_1/N1  ( .A1(\SB1_3_8/i0_3 ), .A2(
        \SB1_3_8/i1[9] ), .ZN(\SB1_3_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_0/N4  ( .A1(\SB1_3_9/i0[7] ), .A2(
        \SB1_3_9/i0_3 ), .A3(\SB1_3_9/i0_0 ), .ZN(
        \SB1_3_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_9/Component_Function_0/N3  ( .A1(\SB1_3_9/i0[10] ), .A2(
        \SB1_3_9/i0_4 ), .A3(\SB1_3_9/i0_3 ), .ZN(
        \SB1_3_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_9/Component_Function_0/N2  ( .A1(\SB1_3_9/i0[8] ), .A2(
        \SB1_3_9/i0[7] ), .A3(\SB1_3_9/i0[6] ), .ZN(
        \SB1_3_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_9/Component_Function_0/N1  ( .A1(\SB1_3_9/i0[10] ), .A2(
        n3979), .ZN(\SB1_3_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_1/N3  ( .A1(\SB1_3_9/i1_5 ), .A2(
        \SB1_3_9/i0[6] ), .A3(n3979), .ZN(
        \SB1_3_9/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_9/Component_Function_1/N1  ( .A1(\SB1_3_9/i0_3 ), .A2(
        \SB1_3_9/i1[9] ), .ZN(\SB1_3_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_10/Component_Function_0/N2  ( .A1(\SB1_3_10/i0[8] ), .A2(
        \SB1_3_10/i0[7] ), .A3(\SB1_3_10/i0[6] ), .ZN(
        \SB1_3_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_10/Component_Function_0/N1  ( .A1(\SB1_3_10/i0[10] ), .A2(
        \SB1_3_10/i0[9] ), .ZN(\SB1_3_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_11/Component_Function_0/N4  ( .A1(\SB1_3_11/i0[7] ), .A2(
        \SB1_3_11/i0_3 ), .A3(\SB1_3_11/i0_0 ), .ZN(
        \SB1_3_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_11/Component_Function_0/N3  ( .A1(\SB1_3_11/i0[10] ), .A2(
        \SB1_3_11/i0_4 ), .A3(\SB1_3_11/i0_3 ), .ZN(
        \SB1_3_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_11/Component_Function_0/N2  ( .A1(\SB1_3_11/i0[8] ), .A2(
        \SB1_3_11/i0[7] ), .A3(\SB1_3_11/i0[6] ), .ZN(
        \SB1_3_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_11/Component_Function_0/N1  ( .A1(\SB1_3_11/i0[10] ), .A2(
        \SB1_3_11/i0[9] ), .ZN(\SB1_3_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_11/Component_Function_1/N2  ( .A1(\SB1_3_11/i0_3 ), .A2(
        \SB1_3_11/i1_7 ), .A3(\SB1_3_11/i0[8] ), .ZN(
        \SB1_3_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_11/Component_Function_1/N1  ( .A1(\SB1_3_11/i0_3 ), .A2(
        \SB1_3_11/i1[9] ), .ZN(\SB1_3_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_12/Component_Function_0/N4  ( .A1(\SB1_3_12/i0[7] ), .A2(
        \SB1_3_12/i0_3 ), .A3(\SB1_3_12/i0_0 ), .ZN(
        \SB1_3_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_12/Component_Function_0/N3  ( .A1(\SB1_3_12/i0[10] ), .A2(
        \SB1_3_12/i0_4 ), .A3(\SB1_3_12/i0_3 ), .ZN(
        \SB1_3_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_0/N3  ( .A1(\SB1_3_13/i0[10] ), .A2(
        \SB1_3_13/i0_4 ), .A3(\SB1_3_13/i0_3 ), .ZN(
        \SB1_3_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_0/N2  ( .A1(\SB1_3_13/i0[8] ), .A2(
        \SB1_3_13/i0[7] ), .A3(\SB1_3_13/i0[6] ), .ZN(
        \SB1_3_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_13/Component_Function_1/N1  ( .A1(\SB1_3_13/i0_3 ), .A2(
        \SB1_3_13/i1[9] ), .ZN(\SB1_3_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_0/N3  ( .A1(\SB1_3_14/i0[10] ), .A2(
        \SB1_3_14/i0_4 ), .A3(\RI1[3][107] ), .ZN(
        \SB1_3_14/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_14/Component_Function_0/N1  ( .A1(\SB1_3_14/i0[10] ), .A2(
        \SB1_3_14/i0[9] ), .ZN(\SB1_3_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_1/N2  ( .A1(\RI1[3][107] ), .A2(
        \SB1_3_14/i1_7 ), .A3(\SB1_3_14/i0[8] ), .ZN(
        \SB1_3_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_14/Component_Function_1/N1  ( .A1(\RI1[3][107] ), .A2(
        \SB1_3_14/i1[9] ), .ZN(\SB1_3_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_15/Component_Function_0/N4  ( .A1(\SB1_3_15/i0[7] ), .A2(
        \SB1_3_15/i0_3 ), .A3(\SB1_3_15/i0_0 ), .ZN(
        \SB1_3_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_15/Component_Function_0/N2  ( .A1(\SB1_3_15/i0[8] ), .A2(
        \SB1_3_15/i0[7] ), .A3(\SB1_3_15/i0[6] ), .ZN(
        \SB1_3_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_15/Component_Function_0/N1  ( .A1(\SB1_3_15/i0[10] ), .A2(
        \SB1_3_15/i0[9] ), .ZN(\SB1_3_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_15/Component_Function_1/N2  ( .A1(\SB1_3_15/i0_3 ), .A2(
        \SB1_3_15/i1_7 ), .A3(\SB1_3_15/i0[8] ), .ZN(
        \SB1_3_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_15/Component_Function_1/N1  ( .A1(\SB1_3_15/i0_3 ), .A2(
        n5431), .ZN(\SB1_3_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_0/N4  ( .A1(\SB1_3_16/i0[7] ), .A2(
        \SB1_3_16/i0_3 ), .A3(\SB1_3_16/i0_0 ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_16/Component_Function_0/N2  ( .A1(\SB1_3_16/i0[8] ), .A2(
        \SB1_3_16/i0[7] ), .A3(\SB1_3_16/i0[6] ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_16/Component_Function_0/N1  ( .A1(\SB1_3_16/i0[10] ), .A2(
        \MC_ARK_ARC_1_2/buf_output[90] ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_17/Component_Function_0/N3  ( .A1(\SB1_3_17/i0[10] ), .A2(
        \SB1_3_17/i0_4 ), .A3(\SB1_3_17/i0_3 ), .ZN(
        \SB1_3_17/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_17/Component_Function_0/N1  ( .A1(\SB1_3_17/i0[10] ), .A2(
        \SB1_3_17/i0[9] ), .ZN(\SB1_3_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_0/N3  ( .A1(\SB1_3_18/i0[10] ), .A2(
        \SB1_3_18/i0_4 ), .A3(\SB1_3_18/i0_3 ), .ZN(
        \SB1_3_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_18/Component_Function_0/N2  ( .A1(\SB1_3_18/i0[8] ), .A2(
        \SB1_3_18/i0[7] ), .A3(\SB1_3_18/i0[6] ), .ZN(
        \SB1_3_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_18/Component_Function_0/N1  ( .A1(\SB1_3_18/i0[10] ), .A2(
        \SB1_3_18/i0[9] ), .ZN(\SB1_3_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_18/Component_Function_1/N1  ( .A1(\SB1_3_18/i0_3 ), .A2(
        \SB1_3_18/i1[9] ), .ZN(\SB1_3_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_0/N3  ( .A1(\SB1_3_19/i0[10] ), .A2(
        \SB1_3_19/i0_4 ), .A3(\SB1_3_19/i0_3 ), .ZN(
        \SB1_3_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_19/Component_Function_0/N2  ( .A1(\SB1_3_19/i0[8] ), .A2(
        \SB1_3_19/i0[7] ), .A3(\SB1_3_19/i0[6] ), .ZN(
        \SB1_3_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_19/Component_Function_0/N1  ( .A1(\SB1_3_19/i0[10] ), .A2(
        \SB1_3_19/i0[9] ), .ZN(\SB1_3_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_1/N3  ( .A1(\SB1_3_19/i1_5 ), .A2(
        \SB1_3_19/i0[6] ), .A3(\SB1_3_19/i0[9] ), .ZN(
        \SB1_3_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_20/Component_Function_0/N3  ( .A1(\SB1_3_20/i0[10] ), .A2(
        \SB1_3_20/i0_4 ), .A3(\SB1_3_20/i0_3 ), .ZN(
        \SB1_3_20/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_20/Component_Function_0/N1  ( .A1(\SB1_3_20/i0[10] ), .A2(
        \SB1_3_20/i0[9] ), .ZN(\SB1_3_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_1/N2  ( .A1(\SB1_3_20/i0_3 ), .A2(
        \SB1_3_20/i1_7 ), .A3(\SB1_3_20/i0[8] ), .ZN(
        \SB1_3_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_21/Component_Function_0/N3  ( .A1(\SB1_3_21/i0[10] ), .A2(
        \SB1_3_21/i0_4 ), .A3(\SB1_3_21/i0_3 ), .ZN(
        \SB1_3_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_21/Component_Function_0/N2  ( .A1(\SB1_3_21/i0[8] ), .A2(
        \SB1_3_21/i0[7] ), .A3(\SB1_3_21/i0[6] ), .ZN(
        \SB1_3_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_21/Component_Function_0/N1  ( .A1(\SB1_3_21/i0[10] ), .A2(
        \SB1_3_21/i0[9] ), .ZN(\SB1_3_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_1/N2  ( .A1(\SB1_3_21/i0_3 ), .A2(
        \SB1_3_21/i1_7 ), .A3(\SB1_3_21/i0[8] ), .ZN(
        \SB1_3_21/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_22/Component_Function_0/N2  ( .A1(\SB1_3_22/i0[8] ), .A2(
        \SB1_3_22/i0[7] ), .A3(\SB1_3_22/i0[6] ), .ZN(
        \SB1_3_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_22/Component_Function_0/N1  ( .A1(\SB1_3_22/i0[10] ), .A2(
        \SB1_3_22/i0[9] ), .ZN(\SB1_3_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_23/Component_Function_0/N2  ( .A1(\SB1_3_23/i0[8] ), .A2(
        \SB1_3_23/i0[7] ), .A3(\SB1_3_23/i0[6] ), .ZN(
        \SB1_3_23/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_24/Component_Function_0/N2  ( .A1(\SB1_3_24/i0[8] ), .A2(
        \SB1_3_24/i0[7] ), .A3(\SB1_3_24/i0[6] ), .ZN(
        \SB1_3_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_24/Component_Function_0/N1  ( .A1(\SB1_3_24/i0[10] ), .A2(
        \SB1_3_24/i0[9] ), .ZN(\SB1_3_24/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_24/Component_Function_1/N1  ( .A1(\SB1_3_24/i0_3 ), .A2(
        \SB1_3_24/i1[9] ), .ZN(\SB1_3_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_0/N3  ( .A1(\SB1_3_25/i0[10] ), .A2(
        \SB1_3_25/i0_4 ), .A3(\SB1_3_25/i0_3 ), .ZN(
        \SB1_3_25/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_25/Component_Function_1/N1  ( .A1(\SB1_3_25/i0_3 ), .A2(
        \SB1_3_25/i1[9] ), .ZN(\SB1_3_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_0/N2  ( .A1(\SB1_3_26/i0[8] ), .A2(
        \SB1_3_26/i0[7] ), .A3(\SB1_3_26/i0[6] ), .ZN(
        \SB1_3_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_26/Component_Function_0/N1  ( .A1(\SB1_3_26/i0[10] ), .A2(
        \SB1_3_26/i0[9] ), .ZN(\SB1_3_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_1/N2  ( .A1(\SB1_3_26/i0_3 ), .A2(
        \SB1_3_26/i1_7 ), .A3(\SB1_3_26/i0[8] ), .ZN(
        \SB1_3_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_26/Component_Function_1/N1  ( .A1(\SB1_3_26/i0_3 ), .A2(
        \SB1_3_26/i1[9] ), .ZN(\SB1_3_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_0/N4  ( .A1(\SB1_3_27/i0[7] ), .A2(
        \SB1_3_27/i0_3 ), .A3(\SB1_3_27/i0_0 ), .ZN(
        \SB1_3_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_27/Component_Function_0/N3  ( .A1(\SB1_3_27/i0[10] ), .A2(
        \SB1_3_27/i0_4 ), .A3(\SB1_3_27/i0_3 ), .ZN(
        \SB1_3_27/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_27/Component_Function_0/N1  ( .A1(\SB1_3_27/i0[10] ), .A2(
        \SB1_3_27/i0[9] ), .ZN(\SB1_3_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_1/N2  ( .A1(\SB1_3_27/i0_3 ), .A2(
        \SB1_3_27/i1_7 ), .A3(\SB1_3_27/i0[8] ), .ZN(
        \SB1_3_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_28/Component_Function_1/N1  ( .A1(\SB1_3_28/i0_3 ), .A2(
        \SB1_3_28/i1[9] ), .ZN(\SB1_3_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_0/N3  ( .A1(\SB1_3_29/i0[10] ), .A2(
        \SB1_3_29/i0_4 ), .A3(\SB1_3_29/i0_3 ), .ZN(
        \SB1_3_29/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_29/Component_Function_0/N1  ( .A1(\SB1_3_29/i0[10] ), .A2(
        \SB1_3_29/i0[9] ), .ZN(\SB1_3_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_1/N3  ( .A1(\SB1_3_30/i1_5 ), .A2(
        \SB1_3_30/i0[6] ), .A3(\SB1_3_30/i0[9] ), .ZN(
        \SB1_3_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_30/Component_Function_1/N2  ( .A1(\SB1_3_30/i0_3 ), .A2(
        \SB1_3_30/i1_7 ), .A3(\SB1_3_30/i0[8] ), .ZN(
        \SB1_3_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_30/Component_Function_1/N1  ( .A1(\SB1_3_30/i0_3 ), .A2(
        \SB1_3_30/i1[9] ), .ZN(\SB1_3_30/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_30/Component_Function_5/N1  ( .A1(\SB1_3_30/i0_0 ), .A2(
        \SB1_3_30/i3[0] ), .ZN(\SB1_3_30/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_31/Component_Function_1/N1  ( .A1(\SB1_3_31/i0_3 ), .A2(
        \SB1_3_31/i1[9] ), .ZN(\SB1_3_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_0/N2  ( .A1(\SB2_3_0/i0[8] ), .A2(
        \SB2_3_0/i0[7] ), .A3(\SB2_3_0/i0[6] ), .ZN(
        \SB2_3_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_0/Component_Function_1/N3  ( .A1(\SB2_3_0/i1_5 ), .A2(
        \SB2_3_0/i0[6] ), .A3(\SB2_3_0/i0[9] ), .ZN(
        \SB2_3_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_0/Component_Function_1/N2  ( .A1(\SB2_3_0/i0_3 ), .A2(
        \SB2_3_0/i1_7 ), .A3(\SB2_3_0/i0[8] ), .ZN(
        \SB2_3_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_0/Component_Function_1/N1  ( .A1(\SB2_3_0/i0_3 ), .A2(
        \SB2_3_0/i1[9] ), .ZN(\SB2_3_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_0/N2  ( .A1(\SB2_3_1/i0[8] ), .A2(
        \SB2_3_1/i0[7] ), .A3(\SB2_3_1/i0[6] ), .ZN(
        \SB2_3_1/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_1/Component_Function_1/N2  ( .A1(\SB2_3_1/i0_3 ), .A2(
        \SB2_3_1/i1_7 ), .A3(\SB2_3_1/i0[8] ), .ZN(
        \SB2_3_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_2/Component_Function_1/N1  ( .A1(\SB2_3_2/i0_3 ), .A2(
        \SB2_3_2/i1[9] ), .ZN(\SB2_3_2/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_3/Component_Function_0/N1  ( .A1(\SB2_3_3/i0[10] ), .A2(
        \SB2_3_3/i0[9] ), .ZN(\SB2_3_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_3/Component_Function_1/N4  ( .A1(\SB2_3_3/i1_7 ), .A2(
        \SB2_3_3/i0[8] ), .A3(\SB1_3_4/buf_output[4] ), .ZN(
        \SB2_3_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_3/Component_Function_1/N2  ( .A1(\SB2_3_3/i0_3 ), .A2(
        \SB2_3_3/i1_7 ), .A3(\SB2_3_3/i0[8] ), .ZN(
        \SB2_3_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_3/Component_Function_1/N1  ( .A1(\SB2_3_3/i0_3 ), .A2(
        \SB2_3_3/i1[9] ), .ZN(\SB2_3_3/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_4/Component_Function_0/N1  ( .A1(\SB2_3_4/i0[10] ), .A2(
        \SB2_3_4/i0[9] ), .ZN(\SB2_3_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_4/Component_Function_1/N3  ( .A1(\SB2_3_4/i1_5 ), .A2(
        \SB2_3_4/i0[6] ), .A3(\SB2_3_4/i0[9] ), .ZN(
        \SB2_3_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_4/Component_Function_1/N2  ( .A1(\SB2_3_4/i0_3 ), .A2(
        \SB2_3_4/i1_7 ), .A3(\SB2_3_4/i0[8] ), .ZN(
        \SB2_3_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_4/Component_Function_1/N1  ( .A1(\SB2_3_4/i0_3 ), .A2(
        \SB2_3_4/i1[9] ), .ZN(\SB2_3_4/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_5/Component_Function_5/N1  ( .A1(\SB2_3_5/i0_0 ), .A2(
        \SB2_3_5/i3[0] ), .ZN(\SB2_3_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_6/Component_Function_0/N2  ( .A1(\SB2_3_6/i0[8] ), .A2(
        \SB2_3_6/i0[7] ), .A3(\SB2_3_6/i0[6] ), .ZN(
        \SB2_3_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_6/Component_Function_0/N1  ( .A1(\SB2_3_6/i0[10] ), .A2(
        \SB2_3_6/i0[9] ), .ZN(\SB2_3_6/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_6/Component_Function_1/N1  ( .A1(\SB2_3_6/i0_3 ), .A2(
        \SB2_3_6/i1[9] ), .ZN(\SB2_3_6/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_7/Component_Function_0/N1  ( .A1(\SB2_3_7/i0[10] ), .A2(
        \SB2_3_7/i0[9] ), .ZN(\SB2_3_7/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_7/Component_Function_1/N1  ( .A1(\SB2_3_7/i0_3 ), .A2(
        \SB2_3_7/i1[9] ), .ZN(\SB2_3_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_8/Component_Function_0/N4  ( .A1(\SB2_3_8/i0[7] ), .A2(
        \SB2_3_8/i0_3 ), .A3(\SB2_3_8/i0_0 ), .ZN(
        \SB2_3_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_8/Component_Function_0/N3  ( .A1(\SB2_3_8/i0[10] ), .A2(
        \SB2_3_8/i0_4 ), .A3(\SB2_3_8/i0_3 ), .ZN(
        \SB2_3_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_8/Component_Function_1/N4  ( .A1(\SB2_3_8/i1_7 ), .A2(
        \SB2_3_8/i0[8] ), .A3(\SB2_3_8/i0_4 ), .ZN(
        \SB2_3_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_8/Component_Function_1/N2  ( .A1(\SB2_3_8/i0_3 ), .A2(
        \SB2_3_8/i1_7 ), .A3(\SB2_3_8/i0[8] ), .ZN(
        \SB2_3_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_8/Component_Function_1/N1  ( .A1(\SB2_3_8/i0_3 ), .A2(
        \SB2_3_8/i1[9] ), .ZN(\SB2_3_8/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_9/Component_Function_0/N1  ( .A1(\SB2_3_9/i0[10] ), .A2(
        \SB2_3_9/i0[9] ), .ZN(\SB2_3_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_1/N2  ( .A1(\SB2_3_10/i0_3 ), .A2(
        \SB2_3_10/i1_7 ), .A3(\SB2_3_10/i0[8] ), .ZN(
        \SB2_3_10/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_11/Component_Function_0/N4  ( .A1(\SB2_3_11/i0[7] ), .A2(
        \SB2_3_11/i0_3 ), .A3(\SB2_3_11/i0_0 ), .ZN(
        \SB2_3_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_11/Component_Function_0/N2  ( .A1(\SB2_3_11/i0[8] ), .A2(
        \SB2_3_11/i0[7] ), .A3(\SB2_3_11/i0[6] ), .ZN(
        \SB2_3_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_11/Component_Function_0/N1  ( .A1(\SB2_3_11/i0[10] ), .A2(
        \SB2_3_11/i0[9] ), .ZN(\SB2_3_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_11/Component_Function_1/N4  ( .A1(\SB2_3_11/i1_7 ), .A2(
        \SB2_3_11/i0[8] ), .A3(\SB2_3_11/i0_4 ), .ZN(
        \SB2_3_11/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_12/Component_Function_5/N1  ( .A1(\SB2_3_12/i0_0 ), .A2(
        \SB2_3_12/i3[0] ), .ZN(\SB2_3_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_1/N2  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i1_7 ), .A3(\SB2_3_13/i0[8] ), .ZN(
        \SB2_3_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_13/Component_Function_1/N1  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i1[9] ), .ZN(\SB2_3_13/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_14/Component_Function_0/N1  ( .A1(\SB2_3_14/i0[10] ), .A2(
        \SB2_3_14/i0[9] ), .ZN(\SB2_3_14/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_14/Component_Function_1/N1  ( .A1(\SB2_3_14/i0_3 ), .A2(
        \SB2_3_14/i1[9] ), .ZN(\SB2_3_14/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_15/Component_Function_0/N1  ( .A1(\SB2_3_15/i0[10] ), .A2(
        \SB2_3_15/i0[9] ), .ZN(\SB2_3_15/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_15/Component_Function_5/N1  ( .A1(\SB2_3_15/i0_0 ), .A2(
        \SB2_3_15/i3[0] ), .ZN(\SB2_3_15/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_16/Component_Function_0/N1  ( .A1(\SB2_3_16/i0[10] ), .A2(
        \SB2_3_16/i0[9] ), .ZN(\SB2_3_16/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_16/Component_Function_1/N1  ( .A1(\SB2_3_16/i0_3 ), .A2(
        \SB2_3_16/i1[9] ), .ZN(\SB2_3_16/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_17/Component_Function_0/N1  ( .A1(\SB2_3_17/i0[10] ), .A2(
        \SB2_3_17/i0[9] ), .ZN(\SB2_3_17/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_17/Component_Function_1/N1  ( .A1(\SB2_3_17/i0_3 ), .A2(
        \SB2_3_17/i1[9] ), .ZN(\SB2_3_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_0/N3  ( .A1(\SB2_3_18/i0[10] ), .A2(
        \SB2_3_18/i0_4 ), .A3(\SB2_3_18/i0_3 ), .ZN(
        \SB2_3_18/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_18/Component_Function_0/N1  ( .A1(\SB2_3_18/i0[10] ), .A2(
        \SB2_3_18/i0[9] ), .ZN(\SB2_3_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_18/Component_Function_1/N1  ( .A1(\SB2_3_18/i0_3 ), .A2(
        \SB2_3_18/i1[9] ), .ZN(\SB2_3_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_20/Component_Function_0/N2  ( .A1(\SB2_3_20/i0[8] ), .A2(
        n6819), .A3(\SB2_3_20/i0[6] ), .ZN(
        \SB2_3_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_20/Component_Function_0/N1  ( .A1(\SB2_3_20/i0[10] ), .A2(
        \SB2_3_20/i0[9] ), .ZN(\SB2_3_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_20/Component_Function_1/N1  ( .A1(\SB2_3_20/i0_3 ), .A2(
        \SB2_3_20/i1[9] ), .ZN(\SB2_3_20/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_21/Component_Function_0/N1  ( .A1(\SB2_3_21/i0[10] ), .A2(
        \SB2_3_21/i0[9] ), .ZN(\SB2_3_21/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_21/Component_Function_1/N1  ( .A1(\SB2_3_21/i0_3 ), .A2(
        \SB2_3_21/i1[9] ), .ZN(\SB2_3_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_1/N2  ( .A1(\SB2_3_22/i0_3 ), .A2(
        \SB2_3_22/i1_7 ), .A3(\SB2_3_22/i0[8] ), .ZN(
        \SB2_3_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_22/Component_Function_5/N1  ( .A1(\SB2_3_22/i0_0 ), .A2(
        \SB2_3_22/i3[0] ), .ZN(\SB2_3_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_0/N2  ( .A1(\SB2_3_23/i0[8] ), .A2(
        \SB2_3_23/i0[7] ), .A3(\SB2_3_23/i0[6] ), .ZN(
        \SB2_3_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_23/Component_Function_0/N1  ( .A1(\SB2_3_23/i0[10] ), .A2(
        \SB2_3_23/i0[9] ), .ZN(\SB2_3_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_1/N2  ( .A1(\SB2_3_23/i0_3 ), .A2(
        \SB2_3_23/i1_7 ), .A3(\SB2_3_23/i0[8] ), .ZN(
        \SB2_3_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_24/Component_Function_0/N4  ( .A1(\SB2_3_24/i0[7] ), .A2(
        \SB2_3_24/i0_3 ), .A3(\SB2_3_24/i0_0 ), .ZN(
        \SB2_3_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_24/Component_Function_0/N2  ( .A1(\SB2_3_24/i0[8] ), .A2(
        \SB2_3_24/i0[7] ), .A3(\SB2_3_24/i0[6] ), .ZN(
        \SB2_3_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_24/Component_Function_0/N1  ( .A1(\SB2_3_24/i0[10] ), .A2(
        \SB2_3_24/i0[9] ), .ZN(\SB2_3_24/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_26/Component_Function_0/N1  ( .A1(\SB2_3_26/i0[10] ), .A2(
        \SB2_3_26/i0[9] ), .ZN(\SB2_3_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_1/N3  ( .A1(\SB2_3_26/i1_5 ), .A2(
        \SB2_3_26/i0[6] ), .A3(\SB2_3_26/i0[9] ), .ZN(
        \SB2_3_26/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_26/Component_Function_1/N1  ( .A1(\SB2_3_26/i0_3 ), .A2(
        \SB2_3_26/i1[9] ), .ZN(\SB2_3_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_0/N2  ( .A1(\SB2_3_27/i0[8] ), .A2(
        \SB2_3_27/i0[7] ), .A3(\SB2_3_27/i0[6] ), .ZN(
        \SB2_3_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_27/Component_Function_0/N1  ( .A1(\SB2_3_27/i0[10] ), .A2(
        \SB2_3_27/i0[9] ), .ZN(\SB2_3_27/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_28/Component_Function_0/N1  ( .A1(\SB2_3_28/i0[10] ), .A2(
        \SB2_3_28/i0[9] ), .ZN(\SB2_3_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_28/Component_Function_1/N2  ( .A1(\SB2_3_28/i0_3 ), .A2(
        \SB2_3_28/i1_7 ), .A3(\SB2_3_28/i0[8] ), .ZN(
        \SB2_3_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_29/Component_Function_0/N3  ( .A1(\SB2_3_29/i0[10] ), .A2(
        \SB2_3_29/i0_4 ), .A3(\SB2_3_29/i0_3 ), .ZN(
        \SB2_3_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_29/Component_Function_1/N2  ( .A1(\SB2_3_29/i0_3 ), .A2(
        \SB2_3_29/i1_7 ), .A3(\SB2_3_29/i0[8] ), .ZN(
        \SB2_3_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_29/Component_Function_1/N1  ( .A1(\SB2_3_29/i0_3 ), .A2(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_0/N3  ( .A1(\SB2_3_30/i0[10] ), .A2(
        \SB2_3_30/i0_4 ), .A3(\SB2_3_30/i0_3 ), .ZN(
        \SB2_3_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_30/Component_Function_0/N2  ( .A1(\SB2_3_30/i0[8] ), .A2(
        \SB2_3_30/i0[7] ), .A3(\SB2_3_30/i0[6] ), .ZN(
        \SB2_3_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_30/Component_Function_0/N1  ( .A1(\SB2_3_30/i0[10] ), .A2(
        \SB2_3_30/i0[9] ), .ZN(\SB2_3_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_1/N2  ( .A1(\SB2_3_30/i0_3 ), .A2(
        \SB2_3_30/i1_7 ), .A3(\SB2_3_30/i0[8] ), .ZN(
        \SB2_3_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_30/Component_Function_1/N1  ( .A1(\SB2_3_30/i0_3 ), .A2(
        \SB2_3_30/i1[9] ), .ZN(\SB2_3_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_31/Component_Function_0/N2  ( .A1(\SB2_3_31/i0[8] ), .A2(
        \SB2_3_31/i0[7] ), .A3(\SB1_3_3/buf_output[1] ), .ZN(
        \SB2_3_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_31/Component_Function_0/N1  ( .A1(\SB2_3_31/i0[10] ), .A2(
        \SB2_3_31/i0[9] ), .ZN(\SB2_3_31/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_31/Component_Function_1/N1  ( .A1(\SB2_3_31/i0_3 ), .A2(
        \SB2_3_31/i1[9] ), .ZN(\SB2_3_31/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_31/Component_Function_5/N1  ( .A1(\SB2_3_31/i0_0 ), .A2(
        \SB2_3_31/i3[0] ), .ZN(\SB2_3_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_0/Component_Function_0/N2  ( .A1(\SB1_4_0/i0[8] ), .A2(
        \SB1_4_0/i0[7] ), .A3(\SB1_4_0/i0[6] ), .ZN(
        \SB1_4_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_1/Component_Function_0/N3  ( .A1(\SB1_4_1/i0[10] ), .A2(
        \SB1_4_1/i0_4 ), .A3(\SB1_4_1/i0_3 ), .ZN(
        \SB1_4_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_1/Component_Function_1/N2  ( .A1(\SB1_4_1/i0_3 ), .A2(
        \SB1_4_1/i1_7 ), .A3(\SB1_4_1/i0[8] ), .ZN(
        \SB1_4_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_2/Component_Function_0/N4  ( .A1(\SB1_4_2/i0[7] ), .A2(
        \SB1_4_2/i0_3 ), .A3(\SB1_4_2/i0_0 ), .ZN(
        \SB1_4_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_2/Component_Function_0/N3  ( .A1(\SB1_4_2/i0[10] ), .A2(
        \SB1_4_2/i0_4 ), .A3(\SB1_4_2/i0_3 ), .ZN(
        \SB1_4_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_2/Component_Function_0/N2  ( .A1(\SB1_4_2/i0[8] ), .A2(
        \SB1_4_2/i0[7] ), .A3(\SB1_4_2/i0[6] ), .ZN(
        \SB1_4_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_2/Component_Function_0/N1  ( .A1(\SB1_4_2/i0[10] ), .A2(
        \SB1_4_2/i0[9] ), .ZN(\SB1_4_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_3/Component_Function_0/N2  ( .A1(\SB1_4_3/i0[8] ), .A2(
        \SB1_4_3/i0[7] ), .A3(\SB1_4_3/i0[6] ), .ZN(
        \SB1_4_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_3/Component_Function_0/N1  ( .A1(\SB1_4_3/i0[10] ), .A2(
        \SB1_4_3/i0[9] ), .ZN(\SB1_4_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_3/Component_Function_1/N2  ( .A1(\SB1_4_3/i0_3 ), .A2(
        \SB1_4_3/i1_7 ), .A3(\SB1_4_3/i0[8] ), .ZN(
        \SB1_4_3/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_4/Component_Function_0/N4  ( .A1(\SB1_4_4/i0[7] ), .A2(
        \SB1_4_4/i0_3 ), .A3(\SB1_4_4/i0_0 ), .ZN(
        \SB1_4_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_4/Component_Function_0/N2  ( .A1(\SB1_4_4/i0[8] ), .A2(
        \SB1_4_4/i0[7] ), .A3(\SB1_4_4/i0[6] ), .ZN(
        \SB1_4_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_4/Component_Function_0/N1  ( .A1(\SB1_4_4/i0[10] ), .A2(
        \SB1_4_4/i0[9] ), .ZN(\SB1_4_4/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_4/Component_Function_1/N1  ( .A1(\SB1_4_4/i0_3 ), .A2(
        \SB1_4_4/i1[9] ), .ZN(\SB1_4_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_5/Component_Function_0/N2  ( .A1(\SB1_4_5/i0[8] ), .A2(
        \SB1_4_5/i0[7] ), .A3(\SB1_4_5/i0[6] ), .ZN(
        \SB1_4_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_5/Component_Function_0/N1  ( .A1(\SB1_4_5/i0[10] ), .A2(
        \SB1_4_5/i0[9] ), .ZN(\SB1_4_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_5/Component_Function_1/N4  ( .A1(\SB1_4_5/i1_7 ), .A2(
        \SB1_4_5/i0[8] ), .A3(\SB1_4_5/i0_4 ), .ZN(
        \SB1_4_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_5/Component_Function_1/N3  ( .A1(\SB1_4_5/i1_5 ), .A2(
        \SB1_4_5/i0[6] ), .A3(\SB1_4_5/i0[9] ), .ZN(
        \SB1_4_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_5/Component_Function_1/N2  ( .A1(\SB1_4_5/i0_3 ), .A2(
        \SB1_4_5/i1_7 ), .A3(\SB1_4_5/i0[8] ), .ZN(
        \SB1_4_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_5/Component_Function_1/N1  ( .A1(\SB1_4_5/i0_3 ), .A2(
        \SB1_4_5/i1[9] ), .ZN(\SB1_4_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_7/Component_Function_0/N2  ( .A1(\SB1_4_7/i0[8] ), .A2(
        \SB1_4_7/i0[7] ), .A3(\SB1_4_7/i0[6] ), .ZN(
        \SB1_4_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_7/Component_Function_0/N1  ( .A1(\SB1_4_7/i0[10] ), .A2(
        \SB1_4_7/i0[9] ), .ZN(\SB1_4_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_7/Component_Function_1/N3  ( .A1(\SB1_4_7/i1_5 ), .A2(
        \SB1_4_7/i0[6] ), .A3(\SB1_4_7/i0[9] ), .ZN(
        \SB1_4_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_7/Component_Function_1/N2  ( .A1(\SB1_4_7/i0_3 ), .A2(
        \SB1_4_7/i1_7 ), .A3(\SB1_4_7/i0[8] ), .ZN(
        \SB1_4_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_7/Component_Function_1/N1  ( .A1(\SB1_4_7/i0_3 ), .A2(
        \SB1_4_7/i1[9] ), .ZN(\SB1_4_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_8/Component_Function_0/N3  ( .A1(\SB1_4_8/i0[10] ), .A2(
        \SB1_4_8/i0_4 ), .A3(\SB1_4_8/i0_3 ), .ZN(
        \SB1_4_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_8/Component_Function_0/N2  ( .A1(\SB1_4_8/i0[8] ), .A2(
        \SB1_4_8/i0[7] ), .A3(\SB1_4_8/i0[6] ), .ZN(
        \SB1_4_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_8/Component_Function_0/N1  ( .A1(\SB1_4_8/i0[10] ), .A2(
        \SB1_4_8/i0[9] ), .ZN(\SB1_4_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_8/Component_Function_1/N2  ( .A1(\SB1_4_8/i0_3 ), .A2(
        \SB1_4_8/i1_7 ), .A3(\SB1_4_8/i0[8] ), .ZN(
        \SB1_4_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_9/Component_Function_0/N3  ( .A1(\SB1_4_9/i0[10] ), .A2(
        \SB1_4_9/i0_4 ), .A3(\SB1_4_9/i0_3 ), .ZN(
        \SB1_4_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_9/Component_Function_0/N2  ( .A1(\SB1_4_9/i0[8] ), .A2(
        \SB1_4_9/i0[7] ), .A3(\SB1_4_9/i0[6] ), .ZN(
        \SB1_4_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_9/Component_Function_0/N1  ( .A1(\SB1_4_9/i0[10] ), .A2(
        \SB1_4_9/i0[9] ), .ZN(\SB1_4_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_9/Component_Function_1/N2  ( .A1(\SB1_4_9/i0_3 ), .A2(
        \SB1_4_9/i1_7 ), .A3(\SB1_4_9/i0[8] ), .ZN(
        \SB1_4_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_9/Component_Function_1/N1  ( .A1(\SB1_4_9/i0_3 ), .A2(
        \SB1_4_9/i1[9] ), .ZN(\SB1_4_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_10/Component_Function_0/N2  ( .A1(\SB1_4_10/i0[8] ), .A2(
        \SB1_4_10/i0[7] ), .A3(\SB1_4_10/i0[6] ), .ZN(
        \SB1_4_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_10/Component_Function_0/N1  ( .A1(\SB1_4_10/i0[10] ), .A2(
        \SB1_4_10/i0[9] ), .ZN(\SB1_4_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_10/Component_Function_1/N1  ( .A1(\RI1[4][131] ), .A2(
        \SB1_4_10/i1[9] ), .ZN(\SB1_4_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_11/Component_Function_0/N3  ( .A1(\SB1_4_11/i0[10] ), .A2(
        \SB1_4_11/i0_4 ), .A3(\SB1_4_11/i0_3 ), .ZN(
        \SB1_4_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_11/Component_Function_0/N2  ( .A1(\SB1_4_11/i0[8] ), .A2(
        \SB1_4_11/i0[7] ), .A3(\SB1_4_11/i0[6] ), .ZN(
        \SB1_4_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_11/Component_Function_0/N1  ( .A1(\SB1_4_11/i0[10] ), .A2(
        \SB1_4_11/i0[9] ), .ZN(\SB1_4_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_11/Component_Function_1/N4  ( .A1(\SB1_4_11/i1_7 ), .A2(
        \SB1_4_11/i0[8] ), .A3(\SB1_4_11/i0_4 ), .ZN(
        \SB1_4_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_11/Component_Function_1/N2  ( .A1(\SB1_4_11/i0_3 ), .A2(
        \SB1_4_11/i1_7 ), .A3(\SB1_4_11/i0[8] ), .ZN(
        \SB1_4_11/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_12/Component_Function_0/N2  ( .A1(\SB1_4_12/i0[8] ), .A2(
        \SB1_4_12/i0[7] ), .A3(\SB1_4_12/i0[6] ), .ZN(
        \SB1_4_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_12/Component_Function_0/N1  ( .A1(\SB1_4_12/i0[10] ), .A2(
        \SB1_4_12/i0[9] ), .ZN(\SB1_4_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_13/Component_Function_0/N4  ( .A1(\SB1_4_13/i0[7] ), .A2(
        \SB1_4_13/i0_3 ), .A3(\SB1_4_13/i0_0 ), .ZN(
        \SB1_4_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_13/Component_Function_0/N2  ( .A1(\SB1_4_13/i0[8] ), .A2(
        \SB1_4_13/i0[7] ), .A3(\SB1_4_13/i0[6] ), .ZN(
        \SB1_4_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_13/Component_Function_0/N1  ( .A1(\SB1_4_13/i0[10] ), .A2(
        \SB1_4_13/i0[9] ), .ZN(\SB1_4_13/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_13/Component_Function_1/N1  ( .A1(\SB1_4_13/i0_3 ), .A2(
        \SB1_4_13/i1[9] ), .ZN(\SB1_4_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_15/Component_Function_0/N3  ( .A1(\SB1_4_15/i0[10] ), .A2(
        \SB1_4_15/i0_4 ), .A3(\SB1_4_15/i0_3 ), .ZN(
        \SB1_4_15/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_4_15/Component_Function_0/N1  ( .A1(\SB1_4_15/i0[10] ), .A2(
        \SB1_4_15/i0[9] ), .ZN(\SB1_4_15/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_15/Component_Function_1/N1  ( .A1(\SB1_4_15/i0_3 ), .A2(
        \SB1_4_15/i1[9] ), .ZN(\SB1_4_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_15/Component_Function_5/N2  ( .A1(\SB1_4_15/i0_0 ), .A2(
        \SB1_4_15/i0[6] ), .A3(\SB1_4_15/i0[10] ), .ZN(
        \SB1_4_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_15/Component_Function_5/N1  ( .A1(\SB1_4_15/i0_0 ), .A2(
        \SB1_4_15/i3[0] ), .ZN(\SB1_4_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_16/Component_Function_0/N2  ( .A1(\SB1_4_16/i0[8] ), .A2(
        \SB1_4_16/i0[7] ), .A3(\SB1_4_16/i0[6] ), .ZN(
        \SB1_4_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_16/Component_Function_0/N1  ( .A1(\SB1_4_16/i0[10] ), .A2(
        \SB1_4_16/i0[9] ), .ZN(\SB1_4_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_17/Component_Function_0/N2  ( .A1(\SB1_4_17/i0[8] ), .A2(
        \SB1_4_17/i0[7] ), .A3(\SB1_4_17/i0[6] ), .ZN(
        \SB1_4_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_18/Component_Function_0/N4  ( .A1(\SB1_4_18/i0[7] ), .A2(
        \SB1_4_18/i0_3 ), .A3(\SB1_4_18/i0_0 ), .ZN(
        \SB1_4_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_18/Component_Function_0/N2  ( .A1(\SB1_4_18/i0[8] ), .A2(
        \SB1_4_18/i0[7] ), .A3(\SB1_4_18/i0[6] ), .ZN(
        \SB1_4_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_18/Component_Function_0/N1  ( .A1(\SB1_4_18/i0[10] ), .A2(
        \SB1_4_18/i0[9] ), .ZN(\SB1_4_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_18/Component_Function_1/N1  ( .A1(\SB1_4_18/i0_3 ), .A2(
        \SB1_4_18/i1[9] ), .ZN(\SB1_4_18/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_19/Component_Function_0/N1  ( .A1(\SB1_4_19/i0[10] ), .A2(
        \SB1_4_19/i0[9] ), .ZN(\SB1_4_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_19/Component_Function_1/N4  ( .A1(\SB1_4_19/i1_7 ), .A2(
        \SB1_4_19/i0[8] ), .A3(\SB1_4_19/i0_4 ), .ZN(
        \SB1_4_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_20/Component_Function_0/N3  ( .A1(\SB1_4_20/i0[10] ), .A2(
        \SB1_4_20/i0_4 ), .A3(\SB1_4_20/i0_3 ), .ZN(
        \SB1_4_20/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_4_20/Component_Function_0/N1  ( .A1(\SB1_4_20/i0[10] ), .A2(
        \SB1_4_20/i0[9] ), .ZN(\SB1_4_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_20/Component_Function_1/N1  ( .A1(\SB1_4_20/i0_3 ), .A2(
        \SB1_4_20/i1[9] ), .ZN(\SB1_4_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_21/Component_Function_0/N4  ( .A1(\SB1_4_21/i0[7] ), .A2(
        \SB1_4_21/i0_3 ), .A3(\SB1_4_21/i0_0 ), .ZN(
        \SB1_4_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_21/Component_Function_0/N3  ( .A1(\SB1_4_21/i0[10] ), .A2(
        \SB1_4_21/i0_4 ), .A3(\SB1_4_21/i0_3 ), .ZN(
        \SB1_4_21/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_4_21/Component_Function_0/N1  ( .A1(\SB1_4_21/i0[10] ), .A2(
        \SB1_4_21/i0[9] ), .ZN(\SB1_4_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_22/Component_Function_0/N2  ( .A1(\SB1_4_22/i0[8] ), .A2(
        \SB1_4_22/i0[7] ), .A3(\SB1_4_22/i0[6] ), .ZN(
        \SB1_4_22/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_23/Component_Function_0/N3  ( .A1(\SB1_4_23/i0[10] ), .A2(
        \SB1_4_23/i0_4 ), .A3(\SB1_4_23/i0_3 ), .ZN(
        \SB1_4_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_23/Component_Function_0/N2  ( .A1(\SB1_4_23/i0[8] ), .A2(
        \SB1_4_23/i0[7] ), .A3(\SB1_4_23/i0[6] ), .ZN(
        \SB1_4_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_23/Component_Function_0/N1  ( .A1(\SB1_4_23/i0[10] ), .A2(
        \SB1_4_23/i0[9] ), .ZN(\SB1_4_23/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_23/Component_Function_1/N1  ( .A1(\SB1_4_23/i0_3 ), .A2(
        \SB1_4_23/i1[9] ), .ZN(\SB1_4_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_24/Component_Function_0/N3  ( .A1(\SB1_4_24/i0[10] ), .A2(
        \SB1_4_24/i0_4 ), .A3(\SB1_4_24/i0_3 ), .ZN(
        \SB1_4_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_24/Component_Function_0/N2  ( .A1(\SB1_4_24/i0[8] ), .A2(
        \SB1_4_24/i0[7] ), .A3(\SB1_4_24/i0[6] ), .ZN(
        \SB1_4_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_24/Component_Function_0/N1  ( .A1(\SB1_4_24/i0[10] ), .A2(
        \SB1_4_24/i0[9] ), .ZN(\SB1_4_24/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_25/Component_Function_0/N1  ( .A1(\SB1_4_25/i0[10] ), .A2(
        \SB1_4_25/i0[9] ), .ZN(\SB1_4_25/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_25/Component_Function_1/N1  ( .A1(\SB1_4_25/i0_3 ), .A2(
        \SB1_4_25/i1[9] ), .ZN(\SB1_4_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_26/Component_Function_0/N3  ( .A1(\SB1_4_26/i0[10] ), .A2(
        \SB1_4_26/i0_4 ), .A3(\SB1_4_26/i0_3 ), .ZN(
        \SB1_4_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_26/Component_Function_0/N2  ( .A1(\SB1_4_26/i0[8] ), .A2(
        \SB1_4_26/i0[7] ), .A3(\SB1_4_26/i0[6] ), .ZN(
        \SB1_4_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_26/Component_Function_0/N1  ( .A1(\SB1_4_26/i0[10] ), .A2(
        \SB1_4_26/i0[9] ), .ZN(\SB1_4_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_26/Component_Function_1/N4  ( .A1(\SB1_4_26/i1_7 ), .A2(
        \SB1_4_26/i0[8] ), .A3(\SB1_4_26/i0_4 ), .ZN(
        \SB1_4_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_27/Component_Function_0/N4  ( .A1(\SB1_4_27/i0[7] ), .A2(
        \SB1_4_27/i0_3 ), .A3(\RI1[4][26] ), .ZN(
        \SB1_4_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_27/Component_Function_0/N2  ( .A1(\SB1_4_27/i0[8] ), .A2(
        \SB1_4_27/i0[7] ), .A3(\SB1_4_27/i0[6] ), .ZN(
        \SB1_4_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_28/Component_Function_0/N1  ( .A1(\SB1_4_28/i0[10] ), .A2(
        \SB1_4_28/i0[9] ), .ZN(\SB1_4_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_29/Component_Function_0/N3  ( .A1(\SB1_4_29/i0[10] ), .A2(
        \SB1_4_29/i0_4 ), .A3(\RI1[4][17] ), .ZN(
        \SB1_4_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_29/Component_Function_0/N2  ( .A1(\SB1_4_29/i0[8] ), .A2(
        \SB1_4_29/i0[7] ), .A3(\SB1_4_29/i0[6] ), .ZN(
        \SB1_4_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_29/Component_Function_1/N1  ( .A1(\RI1[4][17] ), .A2(
        \SB1_4_29/i1[9] ), .ZN(\SB1_4_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_30/Component_Function_0/N3  ( .A1(\SB1_4_30/i0[10] ), .A2(
        \SB1_4_30/i0_4 ), .A3(\SB1_4_30/i0_3 ), .ZN(
        \SB1_4_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_30/Component_Function_0/N2  ( .A1(\SB1_4_30/i0[8] ), .A2(
        \SB1_4_30/i0[7] ), .A3(\SB1_4_30/i0[6] ), .ZN(
        \SB1_4_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_30/Component_Function_0/N1  ( .A1(\SB1_4_30/i0[10] ), .A2(
        \SB1_4_30/i0[9] ), .ZN(\SB1_4_30/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_30/Component_Function_1/N1  ( .A1(\SB1_4_30/i0_3 ), .A2(
        \SB1_4_30/i1[9] ), .ZN(\SB1_4_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_31/Component_Function_0/N2  ( .A1(\SB1_4_31/i0[8] ), .A2(
        \SB1_4_31/i0[7] ), .A3(\SB1_4_31/i0[6] ), .ZN(
        \SB1_4_31/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_0/Component_Function_0/N4  ( .A1(\SB2_4_0/i0[7] ), .A2(
        \SB2_4_0/i0_3 ), .A3(\SB2_4_0/i0_0 ), .ZN(
        \SB2_4_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_0/Component_Function_0/N3  ( .A1(\SB2_4_0/i0[10] ), .A2(
        \SB2_4_0/i0_4 ), .A3(\SB2_4_0/i0_3 ), .ZN(
        \SB2_4_0/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_0/Component_Function_0/N1  ( .A1(\SB2_4_0/i0[10] ), .A2(
        \SB2_4_0/i0[9] ), .ZN(\SB2_4_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_0/Component_Function_1/N3  ( .A1(n3978), .A2(\SB2_4_0/i0[6] ), .A3(\SB2_4_0/i0[9] ), .ZN(\SB2_4_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_0/Component_Function_1/N2  ( .A1(\SB2_4_0/i0_3 ), .A2(
        \SB2_4_0/i1_7 ), .A3(\SB2_4_0/i0[8] ), .ZN(
        \SB2_4_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_0/Component_Function_1/N1  ( .A1(\SB2_4_0/i0_3 ), .A2(
        \SB2_4_0/i1[9] ), .ZN(\SB2_4_0/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_1/Component_Function_0/N1  ( .A1(\SB2_4_1/i0[10] ), .A2(
        \SB2_4_1/i0[9] ), .ZN(\SB2_4_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_1/Component_Function_1/N2  ( .A1(\SB2_4_1/i0_3 ), .A2(
        \SB2_4_1/i1_7 ), .A3(\SB2_4_1/i0[8] ), .ZN(
        \SB2_4_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_1/Component_Function_1/N1  ( .A1(\SB2_4_1/i0_3 ), .A2(
        \SB2_4_1/i1[9] ), .ZN(\SB2_4_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_2/Component_Function_0/N2  ( .A1(\SB2_4_2/i0[8] ), .A2(
        \SB2_4_2/i0[7] ), .A3(\SB2_4_2/i0[6] ), .ZN(
        \SB2_4_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_2/Component_Function_0/N1  ( .A1(\SB2_4_2/i0[10] ), .A2(
        \SB2_4_2/i0[9] ), .ZN(\SB2_4_2/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_2/Component_Function_1/N1  ( .A1(\SB2_4_2/i0_3 ), .A2(
        \SB2_4_2/i1[9] ), .ZN(\SB2_4_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_3/Component_Function_0/N2  ( .A1(\SB2_4_3/i0[8] ), .A2(
        \SB2_4_3/i0[7] ), .A3(\SB2_4_3/i0[6] ), .ZN(
        \SB2_4_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_3/Component_Function_0/N1  ( .A1(\SB2_4_3/i0[10] ), .A2(
        \SB2_4_3/i0[9] ), .ZN(\SB2_4_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_3/Component_Function_1/N3  ( .A1(n3988), .A2(\SB2_4_3/i0[6] ), .A3(\SB2_4_3/i0[9] ), .ZN(\SB2_4_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_3/Component_Function_1/N2  ( .A1(\SB2_4_3/i0_3 ), .A2(
        \SB2_4_3/i1_7 ), .A3(\SB2_4_3/i0[8] ), .ZN(
        \SB2_4_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_3/Component_Function_1/N1  ( .A1(\SB2_4_3/i0_3 ), .A2(
        \SB2_4_3/i1[9] ), .ZN(\SB2_4_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_4/Component_Function_0/N2  ( .A1(\SB2_4_4/i0[8] ), .A2(
        \SB2_4_4/i0[7] ), .A3(\SB2_4_4/i0[6] ), .ZN(
        \SB2_4_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_4/Component_Function_0/N1  ( .A1(\SB2_4_4/i0[10] ), .A2(
        \SB2_4_4/i0[9] ), .ZN(\SB2_4_4/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_4/Component_Function_1/N1  ( .A1(\SB2_4_4/i0_3 ), .A2(
        \SB2_4_4/i1[9] ), .ZN(\SB2_4_4/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_5/Component_Function_0/N1  ( .A1(\SB2_4_5/i0[10] ), .A2(
        \SB2_4_5/i0[9] ), .ZN(\SB2_4_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_6/Component_Function_0/N3  ( .A1(\SB2_4_6/i0[10] ), .A2(
        \SB2_4_6/i0_4 ), .A3(\SB2_4_6/i0_3 ), .ZN(
        \SB2_4_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_6/Component_Function_0/N2  ( .A1(\SB2_4_6/i0[8] ), .A2(
        \SB2_4_6/i0[7] ), .A3(\SB2_4_6/i0[6] ), .ZN(
        \SB2_4_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_6/Component_Function_0/N1  ( .A1(\SB2_4_6/i0[10] ), .A2(
        \SB2_4_6/i0[9] ), .ZN(\SB2_4_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_6/Component_Function_1/N3  ( .A1(\SB2_4_6/i1_5 ), .A2(
        \SB2_4_6/i0[6] ), .A3(\SB2_4_6/i0[9] ), .ZN(
        \SB2_4_6/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_6/Component_Function_1/N1  ( .A1(\SB2_4_6/i0_3 ), .A2(
        \SB2_4_6/i1[9] ), .ZN(\SB2_4_6/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_6/Component_Function_5/N1  ( .A1(\SB2_4_6/i0_0 ), .A2(
        \SB2_4_6/i3[0] ), .ZN(\SB2_4_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_7/Component_Function_0/N3  ( .A1(\SB2_4_7/i0[10] ), .A2(
        \RI3[4][148] ), .A3(\SB2_4_7/i0_3 ), .ZN(
        \SB2_4_7/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_7/Component_Function_0/N1  ( .A1(\SB2_4_7/i0[10] ), .A2(
        \SB2_4_7/i0[9] ), .ZN(\SB2_4_7/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_7/Component_Function_1/N1  ( .A1(\SB2_4_7/i0_3 ), .A2(
        \SB2_4_7/i1[9] ), .ZN(\SB2_4_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_8/Component_Function_0/N4  ( .A1(\SB2_4_8/i0[7] ), .A2(
        \SB2_4_8/i0_3 ), .A3(\SB2_4_8/i0_0 ), .ZN(
        \SB2_4_8/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_4_8/Component_Function_0/N1  ( .A1(\SB2_4_8/i0[10] ), .A2(
        \SB2_4_8/i0[9] ), .ZN(\SB2_4_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_8/Component_Function_1/N4  ( .A1(\SB2_4_8/i1_7 ), .A2(
        \SB2_4_8/i0[8] ), .A3(n3183), .ZN(
        \SB2_4_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_8/Component_Function_1/N3  ( .A1(\SB2_4_8/i1_5 ), .A2(
        \SB2_4_8/i0[6] ), .A3(\SB1_4_13/buf_output[0] ), .ZN(
        \SB2_4_8/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_8/Component_Function_1/N1  ( .A1(\SB2_4_8/i0_3 ), .A2(
        \SB2_4_8/i1[9] ), .ZN(\SB2_4_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_9/Component_Function_0/N2  ( .A1(\SB2_4_9/i0[8] ), .A2(
        \SB2_4_9/i0[7] ), .A3(\SB2_4_9/i0[6] ), .ZN(
        \SB2_4_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_9/Component_Function_0/N1  ( .A1(\SB2_4_9/i0[10] ), .A2(
        \SB2_4_9/i0[9] ), .ZN(\SB2_4_9/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_9/Component_Function_1/N1  ( .A1(\SB2_4_9/i0_3 ), .A2(
        \SB2_4_9/i1[9] ), .ZN(\SB2_4_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_10/Component_Function_0/N4  ( .A1(\SB2_4_10/i0[7] ), .A2(
        \SB2_4_10/i0_3 ), .A3(\SB2_4_10/i0_0 ), .ZN(
        \SB2_4_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_10/Component_Function_0/N3  ( .A1(\SB2_4_10/i0[10] ), .A2(
        \SB2_4_10/i0_4 ), .A3(\SB2_4_10/i0_3 ), .ZN(
        \SB2_4_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_10/Component_Function_0/N2  ( .A1(\SB2_4_10/i0[8] ), .A2(
        \SB2_4_10/i0[7] ), .A3(\SB2_4_10/i0[6] ), .ZN(
        \SB2_4_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_10/Component_Function_0/N1  ( .A1(\SB2_4_10/i0[10] ), .A2(
        \SB2_4_10/i0[9] ), .ZN(\SB2_4_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_10/Component_Function_1/N3  ( .A1(n6269), .A2(
        \SB2_4_10/i0[6] ), .A3(\SB2_4_10/i0[9] ), .ZN(
        \SB2_4_10/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_10/Component_Function_1/N1  ( .A1(\SB2_4_10/i0_3 ), .A2(
        \SB2_4_10/i1[9] ), .ZN(\SB2_4_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_11/Component_Function_0/N3  ( .A1(\SB2_4_11/i0[10] ), .A2(
        \SB2_4_11/i0_4 ), .A3(\SB2_4_11/i0_3 ), .ZN(
        \SB2_4_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_11/Component_Function_0/N2  ( .A1(\SB2_4_11/i0[8] ), .A2(
        \SB2_4_11/i0[7] ), .A3(\SB2_4_11/i0[6] ), .ZN(
        \SB2_4_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_11/Component_Function_0/N1  ( .A1(\SB2_4_11/i0[10] ), .A2(
        \SB2_4_11/i0[9] ), .ZN(\SB2_4_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_11/Component_Function_1/N2  ( .A1(\SB2_4_11/i0_3 ), .A2(
        \SB2_4_11/i1_7 ), .A3(\SB2_4_11/i0[8] ), .ZN(
        \SB2_4_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_12/Component_Function_0/N1  ( .A1(\SB2_4_12/i0[10] ), .A2(
        \SB2_4_12/i0[9] ), .ZN(\SB2_4_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_12/Component_Function_1/N4  ( .A1(\SB2_4_12/i1_7 ), .A2(
        \SB2_4_12/i0[8] ), .A3(\SB2_4_12/i0_4 ), .ZN(
        \SB2_4_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_12/Component_Function_1/N2  ( .A1(\SB2_4_12/i0_3 ), .A2(
        \SB2_4_12/i1_7 ), .A3(\SB2_4_12/i0[8] ), .ZN(
        \SB2_4_12/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_13/Component_Function_0/N2  ( .A1(\SB2_4_13/i0[8] ), .A2(
        \SB2_4_13/i0[7] ), .A3(\SB2_4_13/i0[6] ), .ZN(
        \SB2_4_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_13/Component_Function_0/N1  ( .A1(\SB2_4_13/i0[10] ), .A2(
        \SB2_4_13/i0[9] ), .ZN(\SB2_4_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_13/Component_Function_1/N3  ( .A1(\SB2_4_13/i1_5 ), .A2(
        \SB2_4_13/i0[6] ), .A3(\SB2_4_13/i0[9] ), .ZN(
        \SB2_4_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_13/Component_Function_1/N2  ( .A1(\SB2_4_13/i0_3 ), .A2(
        \SB2_4_13/i1_7 ), .A3(\SB2_4_13/i0[8] ), .ZN(
        \SB2_4_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_14/Component_Function_0/N2  ( .A1(\SB2_4_14/i0[8] ), .A2(
        \SB2_4_14/i0[7] ), .A3(\SB2_4_14/i0[6] ), .ZN(
        \SB2_4_14/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_14/Component_Function_1/N4  ( .A1(\SB2_4_14/i1_7 ), .A2(
        \SB2_4_14/i0[8] ), .A3(\SB1_4_15/buf_output[4] ), .ZN(
        \SB2_4_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_14/Component_Function_1/N3  ( .A1(\SB2_4_14/i1_5 ), .A2(
        \SB2_4_14/i0[6] ), .A3(\SB2_4_14/i0[9] ), .ZN(
        \SB2_4_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_14/Component_Function_1/N2  ( .A1(\SB2_4_14/i0_3 ), .A2(
        \SB2_4_14/i1_7 ), .A3(\SB2_4_14/i0[8] ), .ZN(
        \SB2_4_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_15/Component_Function_0/N3  ( .A1(\SB2_4_15/i0[10] ), .A2(
        \SB2_4_15/i0_4 ), .A3(\SB2_4_15/i0_3 ), .ZN(
        \SB2_4_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_15/Component_Function_0/N2  ( .A1(\SB2_4_15/i0[8] ), .A2(
        \SB2_4_15/i0[7] ), .A3(\SB2_4_15/i0[6] ), .ZN(
        \SB2_4_15/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_15/Component_Function_1/N3  ( .A1(\SB2_4_15/i1_5 ), .A2(
        \SB2_4_15/i0[6] ), .A3(\SB2_4_15/i0[9] ), .ZN(
        \SB2_4_15/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_15/Component_Function_1/N1  ( .A1(\SB2_4_15/i0_3 ), .A2(
        \SB2_4_15/i1[9] ), .ZN(\SB2_4_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_16/Component_Function_0/N3  ( .A1(\SB2_4_16/i0[10] ), .A2(
        \SB2_4_16/i0_4 ), .A3(\SB2_4_16/i0_3 ), .ZN(
        \SB2_4_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_16/Component_Function_0/N2  ( .A1(\SB2_4_16/i0[8] ), .A2(
        \SB2_4_16/i0[7] ), .A3(\SB2_4_16/i0[6] ), .ZN(
        \SB2_4_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_16/Component_Function_0/N1  ( .A1(\SB2_4_16/i0[10] ), .A2(
        \SB2_4_16/i0[9] ), .ZN(\SB2_4_16/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_16/Component_Function_1/N1  ( .A1(\SB2_4_16/i0_3 ), .A2(
        \SB2_4_16/i1[9] ), .ZN(\SB2_4_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_17/Component_Function_0/N3  ( .A1(\SB2_4_17/i0[10] ), .A2(
        \SB2_4_17/i0_4 ), .A3(\SB2_4_17/i0_3 ), .ZN(
        \SB2_4_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_17/Component_Function_0/N2  ( .A1(\SB2_4_17/i0[8] ), .A2(
        \SB2_4_17/i0[7] ), .A3(\SB2_4_17/i0[6] ), .ZN(
        \SB2_4_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_17/Component_Function_0/N1  ( .A1(\SB2_4_17/i0[10] ), .A2(
        \SB2_4_17/i0[9] ), .ZN(\SB2_4_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_17/Component_Function_1/N4  ( .A1(\SB2_4_17/i1_7 ), .A2(
        \SB2_4_17/i0[8] ), .A3(\SB1_4_18/buf_output[4] ), .ZN(
        \SB2_4_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_18/Component_Function_0/N4  ( .A1(\SB2_4_18/i0[7] ), .A2(
        \SB2_4_18/i0_3 ), .A3(\SB2_4_18/i0_0 ), .ZN(
        \SB2_4_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_18/Component_Function_0/N2  ( .A1(\SB2_4_18/i0[8] ), .A2(
        \SB2_4_18/i0[7] ), .A3(\SB2_4_18/i0[6] ), .ZN(
        \SB2_4_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_18/Component_Function_0/N1  ( .A1(\SB2_4_18/i0[10] ), .A2(
        \SB2_4_18/i0[9] ), .ZN(\SB2_4_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_19/Component_Function_0/N2  ( .A1(\SB2_4_19/i0[8] ), .A2(
        \SB2_4_19/i0[7] ), .A3(\SB2_4_19/i0[6] ), .ZN(
        \SB2_4_19/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_19/Component_Function_1/N4  ( .A1(\SB2_4_19/i1_7 ), .A2(
        \SB2_4_19/i0[8] ), .A3(\SB1_4_20/buf_output[4] ), .ZN(
        \SB2_4_19/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_4_19/Component_Function_1/N1  ( .A1(\SB2_4_19/i0_3 ), .A2(
        \SB2_4_19/i1[9] ), .ZN(\SB2_4_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_20/Component_Function_0/N1  ( .A1(\SB2_4_20/i0[10] ), .A2(
        \SB2_4_20/i0[9] ), .ZN(\SB2_4_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_20/Component_Function_1/N1  ( .A1(\SB2_4_20/i0_3 ), .A2(
        \SB2_4_20/i1[9] ), .ZN(\SB2_4_20/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_21/Component_Function_0/N1  ( .A1(\SB2_4_21/i0[10] ), .A2(
        \SB2_4_21/i0[9] ), .ZN(\SB2_4_21/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_21/Component_Function_1/N1  ( .A1(\SB2_4_21/i0_3 ), .A2(
        \SB2_4_21/i1[9] ), .ZN(\SB2_4_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_22/Component_Function_0/N2  ( .A1(\SB2_4_22/i0[8] ), .A2(
        \SB2_4_22/i0[7] ), .A3(\SB2_4_22/i0[6] ), .ZN(
        \SB2_4_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_22/Component_Function_0/N1  ( .A1(\SB2_4_22/i0[10] ), .A2(
        \SB2_4_22/i0[9] ), .ZN(\SB2_4_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_22/Component_Function_1/N2  ( .A1(\SB2_4_22/i0_3 ), .A2(
        \SB2_4_22/i1_7 ), .A3(\SB2_4_22/i0[8] ), .ZN(
        \SB2_4_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_22/Component_Function_1/N1  ( .A1(\SB2_4_22/i0_3 ), .A2(
        \SB2_4_22/i1[9] ), .ZN(\SB2_4_22/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_22/Component_Function_5/N1  ( .A1(\SB2_4_22/i0_0 ), .A2(
        \SB2_4_22/i3[0] ), .ZN(\SB2_4_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_23/Component_Function_0/N3  ( .A1(\SB2_4_23/i0[10] ), .A2(
        \SB2_4_23/i0_4 ), .A3(\SB2_4_23/i0_3 ), .ZN(
        \SB2_4_23/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_23/Component_Function_0/N1  ( .A1(\SB2_4_23/i0[10] ), .A2(
        \SB2_4_23/i0[9] ), .ZN(\SB2_4_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_23/Component_Function_1/N2  ( .A1(\SB2_4_23/i0_3 ), .A2(
        \SB2_4_23/i1_7 ), .A3(\SB2_4_23/i0[8] ), .ZN(
        \SB2_4_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_23/Component_Function_1/N1  ( .A1(\SB2_4_23/i0_3 ), .A2(
        \SB2_4_23/i1[9] ), .ZN(\SB2_4_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_24/Component_Function_0/N4  ( .A1(\SB2_4_24/i0[7] ), .A2(
        \SB2_4_24/i0_3 ), .A3(\SB2_4_24/i0_0 ), .ZN(
        \SB2_4_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_24/Component_Function_0/N2  ( .A1(\SB2_4_24/i0[8] ), .A2(
        \SB2_4_24/i0[7] ), .A3(\SB2_4_24/i0[6] ), .ZN(
        \SB2_4_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_24/Component_Function_0/N1  ( .A1(\SB2_4_24/i0[10] ), .A2(
        \SB2_4_24/i0[9] ), .ZN(\SB2_4_24/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_24/Component_Function_1/N1  ( .A1(\SB2_4_24/i0_3 ), .A2(
        n5443), .ZN(\SB2_4_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_26/Component_Function_0/N2  ( .A1(\SB2_4_26/i0[8] ), .A2(
        \SB2_4_26/i0[7] ), .A3(\SB2_4_26/i0[6] ), .ZN(
        \SB2_4_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_26/Component_Function_1/N2  ( .A1(\SB2_4_26/i0_3 ), .A2(
        \SB2_4_26/i1_7 ), .A3(\SB2_4_26/i0[8] ), .ZN(
        \SB2_4_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_26/Component_Function_5/N1  ( .A1(\SB2_4_26/i0_0 ), .A2(
        \SB2_4_26/i3[0] ), .ZN(\SB2_4_26/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_27/Component_Function_0/N1  ( .A1(\SB2_4_27/i0[10] ), .A2(
        \SB2_4_27/i0[9] ), .ZN(\SB2_4_27/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_27/Component_Function_1/N1  ( .A1(\SB2_4_27/i0_3 ), .A2(
        \SB2_4_27/i1[9] ), .ZN(\SB2_4_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_28/Component_Function_0/N4  ( .A1(\SB2_4_28/i0[7] ), .A2(
        \SB2_4_28/i0_3 ), .A3(\SB2_4_28/i0_0 ), .ZN(
        \SB2_4_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_28/Component_Function_0/N2  ( .A1(n4000), .A2(
        \SB2_4_28/i0[7] ), .A3(\SB2_4_28/i0[6] ), .ZN(
        \SB2_4_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_28/Component_Function_0/N1  ( .A1(\SB2_4_28/i0[10] ), .A2(
        \SB2_4_28/i0[9] ), .ZN(\SB2_4_28/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_28/Component_Function_1/N1  ( .A1(\SB2_4_28/i0_3 ), .A2(
        \SB2_4_28/i1[9] ), .ZN(\SB2_4_28/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_28/Component_Function_5/N1  ( .A1(\SB2_4_28/i0_0 ), .A2(
        \SB2_4_28/i3[0] ), .ZN(\SB2_4_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_29/Component_Function_0/N2  ( .A1(\SB2_4_29/i0[8] ), .A2(
        \SB2_4_29/i0[7] ), .A3(\SB2_4_29/i0[6] ), .ZN(
        \SB2_4_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_29/Component_Function_0/N1  ( .A1(\SB2_4_29/i0[10] ), .A2(
        \SB2_4_29/i0[9] ), .ZN(\SB2_4_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_29/Component_Function_1/N3  ( .A1(\SB2_4_29/i1_5 ), .A2(
        \SB2_4_29/i0[6] ), .A3(\SB2_4_29/i0[9] ), .ZN(
        \SB2_4_29/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_29/Component_Function_1/N1  ( .A1(\SB2_4_29/i0_3 ), .A2(
        \SB2_4_29/i1[9] ), .ZN(\SB2_4_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_30/Component_Function_0/N3  ( .A1(\SB2_4_30/i0[10] ), .A2(
        \SB1_4_31/buf_output[4] ), .A3(\SB2_4_30/i0_3 ), .ZN(
        \SB2_4_30/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_30/Component_Function_0/N1  ( .A1(\SB2_4_30/i0[10] ), .A2(
        \SB2_4_30/i0[9] ), .ZN(\SB2_4_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_30/Component_Function_1/N2  ( .A1(\SB2_4_30/i0_3 ), .A2(
        \SB2_4_30/i1_7 ), .A3(\SB2_4_30/i0[8] ), .ZN(
        \SB2_4_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_30/Component_Function_1/N1  ( .A1(\SB2_4_30/i0_3 ), .A2(
        \SB2_4_30/i1[9] ), .ZN(\SB2_4_30/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_31/Component_Function_0/N1  ( .A1(\SB2_4_31/i0[10] ), .A2(
        \SB2_4_31/i0[9] ), .ZN(\SB2_4_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_31/Component_Function_1/N4  ( .A1(\SB2_4_31/i1_7 ), .A2(
        \SB2_4_31/i0[8] ), .A3(\SB2_4_31/i0_4 ), .ZN(
        \SB2_4_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_31/Component_Function_1/N3  ( .A1(\SB2_4_31/i1_5 ), .A2(
        \SB2_4_31/i0[6] ), .A3(\SB2_4_31/i0[9] ), .ZN(
        \SB2_4_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_31/Component_Function_1/N2  ( .A1(\SB2_4_31/i0_3 ), .A2(
        \SB2_4_31/i1_7 ), .A3(\SB2_4_31/i0[8] ), .ZN(
        \SB2_4_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_31/Component_Function_1/N1  ( .A1(\SB2_4_31/i0_3 ), .A2(
        \SB2_4_31/i1[9] ), .ZN(\SB2_4_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_0/N4  ( .A1(\SB3_0/i0[7] ), .A2(
        \SB3_0/i0_3 ), .A3(\SB3_0/i0_0 ), .ZN(
        \SB3_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_0/Component_Function_0/N2  ( .A1(\SB3_0/i0[8] ), .A2(
        \SB3_0/i0[7] ), .A3(\SB3_0/i0[6] ), .ZN(
        \SB3_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB3_1/Component_Function_0/N2  ( .A1(\SB3_1/i0[8] ), .A2(
        \SB3_1/i0[7] ), .A3(\SB3_1/i0[6] ), .ZN(
        \SB3_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_1/Component_Function_0/N1  ( .A1(\SB3_1/i0[10] ), .A2(
        \SB3_1/i0[9] ), .ZN(\SB3_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_1/Component_Function_1/N2  ( .A1(\SB3_1/i0_3 ), .A2(
        \SB3_1/i1_7 ), .A3(\SB3_1/i0[8] ), .ZN(
        \SB3_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB3_2/Component_Function_0/N3  ( .A1(\SB3_2/i0[10] ), .A2(
        \SB3_2/i0_4 ), .A3(\SB3_2/i0_3 ), .ZN(
        \SB3_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_3/Component_Function_1/N2  ( .A1(\SB3_3/i0_3 ), .A2(
        \SB3_3/i1_7 ), .A3(\SB3_3/i0[8] ), .ZN(
        \SB3_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_3/Component_Function_1/N1  ( .A1(\SB3_3/i0_3 ), .A2(
        \SB3_3/i1[9] ), .ZN(\SB3_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_0/N4  ( .A1(\SB3_4/i0[7] ), .A2(
        \SB3_4/i0_3 ), .A3(\SB3_4/i0_0 ), .ZN(
        \SB3_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_4/Component_Function_0/N3  ( .A1(\SB3_4/i0[10] ), .A2(
        \SB3_4/i0_4 ), .A3(\SB3_4/i0_3 ), .ZN(
        \SB3_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_4/Component_Function_0/N2  ( .A1(\SB3_4/i0[8] ), .A2(
        \SB3_4/i0[7] ), .A3(\SB3_4/i0[6] ), .ZN(
        \SB3_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_4/Component_Function_0/N1  ( .A1(\SB3_4/i0[10] ), .A2(
        \SB3_4/i0[9] ), .ZN(\SB3_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_1/N3  ( .A1(\SB3_4/i1_5 ), .A2(
        \SB3_4/i0[6] ), .A3(\SB3_4/i0[9] ), .ZN(
        \SB3_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_4/Component_Function_1/N2  ( .A1(\SB3_4/i0_3 ), .A2(
        \SB3_4/i1_7 ), .A3(\SB3_4/i0[8] ), .ZN(
        \SB3_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_4/Component_Function_1/N1  ( .A1(\SB3_4/i0_3 ), .A2(
        \SB3_4/i1[9] ), .ZN(\SB3_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_5/N2  ( .A1(\SB3_4/i0_0 ), .A2(
        \SB3_4/i0[6] ), .A3(\SB3_4/i0[10] ), .ZN(
        \SB3_4/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_4/Component_Function_5/N1  ( .A1(\SB3_4/i0_0 ), .A2(
        \SB3_4/i3[0] ), .ZN(\SB3_4/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB3_5/Component_Function_0/N1  ( .A1(\SB3_5/i0[10] ), .A2(
        \SB3_5/i0[9] ), .ZN(\SB3_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_1/N4  ( .A1(\SB3_5/i1_7 ), .A2(
        \SB3_5/i0[8] ), .A3(\SB3_5/i0_4 ), .ZN(
        \SB3_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_6/Component_Function_0/N3  ( .A1(\SB3_6/i0[10] ), .A2(
        \SB3_6/i0_4 ), .A3(\SB3_6/i0_3 ), .ZN(
        \SB3_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_6/Component_Function_0/N2  ( .A1(\SB3_6/i0[8] ), .A2(
        \SB3_6/i0[7] ), .A3(\SB3_6/i0[6] ), .ZN(
        \SB3_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_6/Component_Function_0/N1  ( .A1(\SB3_6/i0[10] ), .A2(
        \SB3_6/i0[9] ), .ZN(\SB3_6/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB3_6/Component_Function_1/N1  ( .A1(\SB3_6/i0_3 ), .A2(
        \SB3_6/i1[9] ), .ZN(\SB3_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_0/N3  ( .A1(\SB3_7/i0[10] ), .A2(
        \SB3_7/i0_4 ), .A3(\SB3_7/i0_3 ), .ZN(
        \SB3_7/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_7/Component_Function_0/N1  ( .A1(\SB3_7/i0[10] ), .A2(
        \SB3_7/i0[9] ), .ZN(\SB3_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_1/N3  ( .A1(\SB3_7/i1_5 ), .A2(
        \SB3_7/i0[6] ), .A3(\SB3_7/i0[9] ), .ZN(
        \SB3_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_8/Component_Function_0/N2  ( .A1(\SB3_8/i0[8] ), .A2(
        \SB3_8/i0[7] ), .A3(\SB3_8/i0[6] ), .ZN(
        \SB3_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_8/Component_Function_0/N1  ( .A1(\SB3_8/i0[10] ), .A2(
        \SB3_8/i0[9] ), .ZN(\SB3_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_1/N4  ( .A1(\SB3_8/i1_7 ), .A2(
        \SB3_8/i0[8] ), .A3(\SB3_8/i0_4 ), .ZN(
        \SB3_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_8/Component_Function_1/N3  ( .A1(\SB3_8/i1_5 ), .A2(
        \SB3_8/i0[6] ), .A3(\SB3_8/i0[9] ), .ZN(
        \SB3_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_8/Component_Function_1/N2  ( .A1(\SB3_8/i0_3 ), .A2(
        \SB3_8/i1_7 ), .A3(\SB3_8/i0[8] ), .ZN(
        \SB3_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_8/Component_Function_1/N1  ( .A1(\SB3_8/i0_3 ), .A2(
        \SB3_8/i1[9] ), .ZN(\SB3_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_0/N4  ( .A1(\SB3_9/i0[7] ), .A2(
        \SB3_9/i0_3 ), .A3(\SB3_9/i0_0 ), .ZN(
        \SB3_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_9/Component_Function_0/N3  ( .A1(\SB3_9/i0[10] ), .A2(
        \SB3_9/i0_4 ), .A3(\SB3_9/i0_3 ), .ZN(
        \SB3_9/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_9/Component_Function_0/N1  ( .A1(\SB3_9/i0[10] ), .A2(
        \SB3_9/i0[9] ), .ZN(\SB3_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_1/N3  ( .A1(\SB3_9/i1_5 ), .A2(
        \SB3_9/i0[6] ), .A3(\SB3_9/i0[9] ), .ZN(
        \SB3_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_9/Component_Function_1/N2  ( .A1(\SB3_9/i0_3 ), .A2(
        \SB3_9/i1_7 ), .A3(\SB3_9/i0[8] ), .ZN(
        \SB3_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_9/Component_Function_1/N1  ( .A1(\SB3_9/i0_3 ), .A2(
        \SB3_9/i1[9] ), .ZN(\SB3_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_5/N2  ( .A1(\SB3_9/i0_0 ), .A2(
        \SB3_9/i0[6] ), .A3(\SB3_9/i0[10] ), .ZN(
        \SB3_9/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB3_9/Component_Function_5/N1  ( .A1(\SB3_9/i0_0 ), .A2(
        \SB3_9/i3[0] ), .ZN(\SB3_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_0/N3  ( .A1(\SB3_10/i0[10] ), .A2(
        \SB3_10/i0_4 ), .A3(\SB3_10/i0_3 ), .ZN(
        \SB3_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_10/Component_Function_0/N2  ( .A1(\SB3_10/i0[8] ), .A2(
        \SB3_10/i0[7] ), .A3(\SB3_10/i0[6] ), .ZN(
        \SB3_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_10/Component_Function_0/N1  ( .A1(\SB3_10/i0[10] ), .A2(
        \SB3_10/i0[9] ), .ZN(\SB3_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_1/N3  ( .A1(\SB3_10/i1_5 ), .A2(
        \SB3_10/i0[6] ), .A3(\SB3_10/i0[9] ), .ZN(
        \SB3_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_10/Component_Function_1/N2  ( .A1(\SB3_10/i0_3 ), .A2(
        \SB3_10/i1_7 ), .A3(\SB3_10/i0[8] ), .ZN(
        \SB3_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_10/Component_Function_1/N1  ( .A1(\SB3_10/i0_3 ), .A2(
        \SB3_10/i1[9] ), .ZN(\SB3_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_11/Component_Function_1/N2  ( .A1(\SB3_11/i0_3 ), .A2(
        \SB3_11/i1_7 ), .A3(\SB3_11/i0[8] ), .ZN(
        \SB3_11/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB3_12/Component_Function_0/N2  ( .A1(\SB3_12/i0[8] ), .A2(
        \SB3_12/i0[7] ), .A3(\SB3_12/i0[6] ), .ZN(
        \SB3_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_12/Component_Function_0/N1  ( .A1(\SB3_12/i0[10] ), .A2(
        \SB3_12/i0[9] ), .ZN(\SB3_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_1/N4  ( .A1(\SB3_12/i1_7 ), .A2(
        \SB3_12/i0[8] ), .A3(\SB3_12/i0_4 ), .ZN(
        \SB3_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_13/Component_Function_1/N2  ( .A1(\SB3_13/i0_3 ), .A2(
        \SB3_13/i1_7 ), .A3(\SB3_13/i0[8] ), .ZN(
        \SB3_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB3_14/Component_Function_0/N3  ( .A1(\SB3_14/i0[10] ), .A2(
        \SB3_14/i0_4 ), .A3(\SB3_14/i0_3 ), .ZN(
        \SB3_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_14/Component_Function_0/N2  ( .A1(\SB3_14/i0[8] ), .A2(
        \SB3_14/i0[7] ), .A3(\SB3_14/i0[6] ), .ZN(
        \SB3_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_14/Component_Function_0/N1  ( .A1(\SB3_14/i0[10] ), .A2(
        \SB3_14/i0[9] ), .ZN(\SB3_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_1/N3  ( .A1(\SB3_14/i1_5 ), .A2(
        \SB3_14/i0[6] ), .A3(\SB3_14/i0[9] ), .ZN(
        \SB3_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_15/Component_Function_0/N3  ( .A1(\SB3_15/i0[10] ), .A2(
        \SB3_15/i0_4 ), .A3(\SB3_15/i0_3 ), .ZN(
        \SB3_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_15/Component_Function_1/N2  ( .A1(\SB3_15/i0_3 ), .A2(
        \SB3_15/i1_7 ), .A3(\SB3_15/i0[8] ), .ZN(
        \SB3_15/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB3_16/Component_Function_0/N4  ( .A1(\SB3_16/i0[7] ), .A2(
        \SB3_16/i0_3 ), .A3(\SB3_16/i0_0 ), .ZN(
        \SB3_16/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB3_16/Component_Function_0/N1  ( .A1(\SB3_16/i0[10] ), .A2(
        \SB3_16/i0[9] ), .ZN(\SB3_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_1/N2  ( .A1(\SB3_16/i0_3 ), .A2(
        \SB3_16/i1_7 ), .A3(\SB3_16/i0[8] ), .ZN(
        \SB3_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_16/Component_Function_1/N1  ( .A1(\SB3_16/i0_3 ), .A2(
        \SB3_16/i1[9] ), .ZN(\SB3_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_0/N2  ( .A1(\SB3_17/i0[8] ), .A2(
        \SB3_17/i0[7] ), .A3(\SB3_17/i0[6] ), .ZN(
        \SB3_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_17/Component_Function_0/N1  ( .A1(\SB3_17/i0[10] ), .A2(
        \SB3_17/i0[9] ), .ZN(\SB3_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_1/N3  ( .A1(\SB3_17/i1_5 ), .A2(
        \SB3_17/i0[6] ), .A3(\SB3_17/i0[9] ), .ZN(
        \SB3_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_18/Component_Function_0/N3  ( .A1(\SB3_18/i0[10] ), .A2(
        \SB3_18/i0_4 ), .A3(\SB3_18/i0_3 ), .ZN(
        \SB3_18/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_18/Component_Function_0/N1  ( .A1(\SB3_18/i0[10] ), .A2(
        \SB3_18/i0[9] ), .ZN(\SB3_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_18/Component_Function_1/N2  ( .A1(\SB3_18/i0_3 ), .A2(
        \SB3_18/i1_7 ), .A3(\SB3_18/i0[8] ), .ZN(
        \SB3_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_18/Component_Function_1/N1  ( .A1(\SB3_18/i0_3 ), .A2(
        \SB3_18/i1[9] ), .ZN(\SB3_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_0/N3  ( .A1(\SB3_19/i0[10] ), .A2(
        \SB3_19/i0_4 ), .A3(\SB3_19/i0_3 ), .ZN(
        \SB3_19/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_19/Component_Function_0/N1  ( .A1(\SB3_19/i0[10] ), .A2(
        \SB3_19/i0[9] ), .ZN(\SB3_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_1/N2  ( .A1(\SB3_19/i0_3 ), .A2(
        \SB3_19/i1_7 ), .A3(\SB3_19/i0[8] ), .ZN(
        \SB3_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_19/Component_Function_1/N1  ( .A1(\SB3_19/i0_3 ), .A2(
        \SB3_19/i1[9] ), .ZN(\SB3_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_0/N2  ( .A1(\SB3_20/i0[8] ), .A2(
        \SB3_20/i0[7] ), .A3(\SB3_20/i0[6] ), .ZN(
        \SB3_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_20/Component_Function_0/N1  ( .A1(\SB3_20/i0[10] ), .A2(
        \SB3_20/i0[9] ), .ZN(\SB3_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB3_21/Component_Function_0/N1  ( .A1(\SB3_21/i0[10] ), .A2(
        \SB3_21/i0[9] ), .ZN(\SB3_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_1/N2  ( .A1(\SB3_21/i0_3 ), .A2(
        \SB3_21/i1_7 ), .A3(\SB3_21/i0[8] ), .ZN(
        \SB3_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_21/Component_Function_1/N1  ( .A1(\SB3_21/i0_3 ), .A2(
        \SB3_21/i1[9] ), .ZN(\SB3_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_0/N3  ( .A1(\SB3_22/i0[10] ), .A2(
        \SB3_22/i0_4 ), .A3(\SB3_22/i0_3 ), .ZN(
        \SB3_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_22/Component_Function_0/N2  ( .A1(\SB3_22/i0[8] ), .A2(
        \SB3_22/i0[7] ), .A3(\SB3_22/i0[6] ), .ZN(
        \SB3_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_22/Component_Function_0/N1  ( .A1(\SB3_22/i0[10] ), .A2(
        \SB3_22/i0[9] ), .ZN(\SB3_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_1/N2  ( .A1(\SB3_22/i0_3 ), .A2(
        \SB3_22/i1_7 ), .A3(\SB3_22/i0[8] ), .ZN(
        \SB3_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_22/Component_Function_1/N1  ( .A1(\SB3_22/i0_3 ), .A2(
        \SB3_22/i1[9] ), .ZN(\SB3_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_0/N3  ( .A1(\SB3_23/i0[10] ), .A2(
        \SB3_23/i0_4 ), .A3(\SB3_23/i0_3 ), .ZN(
        \SB3_23/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_23/Component_Function_0/N1  ( .A1(\SB3_23/i0[10] ), .A2(
        \SB3_23/i0[9] ), .ZN(\SB3_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_1/N4  ( .A1(\SB3_23/i1_7 ), .A2(
        \SB3_23/i0[8] ), .A3(\SB3_23/i0_4 ), .ZN(
        \SB3_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_23/Component_Function_1/N2  ( .A1(\SB3_23/i0_3 ), .A2(
        \SB3_23/i1_7 ), .A3(\SB3_23/i0[8] ), .ZN(
        \SB3_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB3_24/Component_Function_0/N2  ( .A1(\SB3_24/i0[8] ), .A2(
        \SB3_24/i0[7] ), .A3(\SB3_24/i0[6] ), .ZN(
        \SB3_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_24/Component_Function_0/N1  ( .A1(\SB3_24/i0[10] ), .A2(
        \SB3_24/i0[9] ), .ZN(\SB3_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_24/Component_Function_1/N3  ( .A1(\SB3_24/i1_5 ), .A2(
        \SB3_24/i0[6] ), .A3(\SB3_24/i0[9] ), .ZN(
        \SB3_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_24/Component_Function_1/N2  ( .A1(\SB3_24/i0_3 ), .A2(
        \SB3_24/i1_7 ), .A3(\SB3_24/i0[8] ), .ZN(
        \SB3_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_24/Component_Function_1/N1  ( .A1(\SB3_24/i0_3 ), .A2(
        \SB3_24/i1[9] ), .ZN(\SB3_24/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB3_25/Component_Function_1/N1  ( .A1(\SB3_25/i0_3 ), .A2(
        \SB3_25/i1[9] ), .ZN(\SB3_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_0/N2  ( .A1(\SB3_26/i0[8] ), .A2(
        \SB3_26/i0[7] ), .A3(\SB3_26/i0[6] ), .ZN(
        \SB3_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB3_26/Component_Function_1/N4  ( .A1(\SB3_26/i1_7 ), .A2(
        \SB3_26/i0[8] ), .A3(\SB3_26/i0_4 ), .ZN(
        \SB3_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_26/Component_Function_1/N2  ( .A1(\SB3_26/i0_3 ), .A2(
        \SB3_26/i1_7 ), .A3(\SB3_26/i0[8] ), .ZN(
        \SB3_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_26/Component_Function_1/N1  ( .A1(\SB3_26/i0_3 ), .A2(
        \SB3_26/i1[9] ), .ZN(\SB3_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_0/N4  ( .A1(\SB3_27/i0[7] ), .A2(
        \SB3_27/i0_3 ), .A3(\SB3_27/i0_0 ), .ZN(
        \SB3_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_27/Component_Function_0/N3  ( .A1(\SB3_27/i0[10] ), .A2(
        \SB3_27/i0_4 ), .A3(\SB3_27/i0_3 ), .ZN(
        \SB3_27/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_27/Component_Function_0/N1  ( .A1(\SB3_27/i0[10] ), .A2(
        \SB3_27/i0[9] ), .ZN(\SB3_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_0/N3  ( .A1(\SB3_28/i0[10] ), .A2(
        \SB3_28/i0_4 ), .A3(\SB3_28/i0_3 ), .ZN(
        \SB3_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_28/Component_Function_0/N2  ( .A1(\SB3_28/i0[8] ), .A2(
        \SB3_28/i0[7] ), .A3(\SB3_28/i0[6] ), .ZN(
        \SB3_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_28/Component_Function_0/N1  ( .A1(\SB3_28/i0[10] ), .A2(
        \SB3_28/i0[9] ), .ZN(\SB3_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_1/N4  ( .A1(\SB3_28/i1_7 ), .A2(
        \SB3_28/i0[8] ), .A3(\SB3_28/i0_4 ), .ZN(
        \SB3_28/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB3_28/Component_Function_1/N1  ( .A1(\SB3_28/i0_3 ), .A2(
        \SB3_28/i1[9] ), .ZN(\SB3_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_0/N3  ( .A1(\SB3_29/i0[10] ), .A2(
        \SB3_29/i0_4 ), .A3(n3976), .ZN(
        \SB3_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_29/Component_Function_0/N2  ( .A1(\SB3_29/i0[8] ), .A2(
        \SB3_29/i0[7] ), .A3(\SB3_29/i0[6] ), .ZN(
        \SB3_29/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB3_29/Component_Function_1/N4  ( .A1(\SB3_29/i1_7 ), .A2(
        \SB3_29/i0[8] ), .A3(\SB3_29/i0_4 ), .ZN(
        \SB3_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_29/Component_Function_1/N3  ( .A1(\SB3_29/i1_5 ), .A2(
        \SB3_29/i0[6] ), .A3(\SB3_29/i0[9] ), .ZN(
        \SB3_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_29/Component_Function_1/N2  ( .A1(\RI1[5][17] ), .A2(
        \SB3_29/i1_7 ), .A3(\SB3_29/i0[8] ), .ZN(
        \SB3_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_29/Component_Function_1/N1  ( .A1(\RI1[5][17] ), .A2(
        \SB3_29/i1[9] ), .ZN(\SB3_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_0/N2  ( .A1(\SB3_30/i0[8] ), .A2(
        \SB3_30/i0[7] ), .A3(\SB3_30/i0[6] ), .ZN(
        \SB3_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_30/Component_Function_0/N1  ( .A1(\SB3_30/i0[10] ), .A2(
        \SB3_30/i0[9] ), .ZN(\SB3_30/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB3_30/Component_Function_1/N1  ( .A1(\SB3_30/i0_3 ), .A2(
        \SB3_30/i1[9] ), .ZN(\SB3_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_31/Component_Function_1/N4  ( .A1(\SB3_31/i1_7 ), .A2(
        \SB3_31/i0[8] ), .A3(\SB3_31/i0_4 ), .ZN(
        \SB3_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_0/Component_Function_0/N2  ( .A1(\SB4_0/i0[8] ), .A2(
        \SB4_0/i0[7] ), .A3(\SB4_0/i0[6] ), .ZN(
        \SB4_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_0/Component_Function_1/N2  ( .A1(\SB4_0/i0_3 ), .A2(
        \SB4_0/i1_7 ), .A3(\SB4_0/i0[8] ), .ZN(
        \SB4_0/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_0/Component_Function_5/N1  ( .A1(\SB4_0/i0_0 ), .A2(
        \SB4_0/i3[0] ), .ZN(\SB4_0/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB4_1/Component_Function_0/N1  ( .A1(\SB4_1/i0[10] ), .A2(
        \SB4_1/i0[9] ), .ZN(\SB4_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_1/Component_Function_1/N2  ( .A1(\SB4_1/i0_3 ), .A2(
        \SB4_1/i1_7 ), .A3(\SB4_1/i0[8] ), .ZN(
        \SB4_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_1/Component_Function_5/N4  ( .A1(\SB4_1/i0[9] ), .A2(
        \SB4_1/i0[6] ), .A3(\SB4_1/i0_4 ), .ZN(
        \SB4_1/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_1/Component_Function_5/N1  ( .A1(\SB4_1/i0_0 ), .A2(
        \SB4_1/i3[0] ), .ZN(\SB4_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_2/Component_Function_0/N2  ( .A1(\SB4_2/i0[8] ), .A2(
        \SB4_2/i0[7] ), .A3(\SB4_2/i0[6] ), .ZN(
        \SB4_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_2/Component_Function_0/N1  ( .A1(\SB4_2/i0[10] ), .A2(
        \SB4_2/i0[9] ), .ZN(\SB4_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_2/Component_Function_1/N4  ( .A1(\SB4_2/i1_7 ), .A2(
        \SB4_2/i0[8] ), .A3(\SB4_2/i0_4 ), .ZN(
        \SB4_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_2/Component_Function_1/N3  ( .A1(\SB4_2/i1_5 ), .A2(
        \SB4_2/i0[6] ), .A3(\SB4_2/i0[9] ), .ZN(
        \SB4_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_2/Component_Function_1/N2  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i1_7 ), .A3(\SB4_2/i0[8] ), .ZN(
        \SB4_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_2/Component_Function_1/N1  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i1[9] ), .ZN(\SB4_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_2/Component_Function_5/N4  ( .A1(\SB4_2/i0[9] ), .A2(
        \SB4_2/i0[6] ), .A3(\SB4_2/i0_4 ), .ZN(
        \SB4_2/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_2/Component_Function_5/N1  ( .A1(\SB4_2/i0_0 ), .A2(
        \SB4_2/i3[0] ), .ZN(\SB4_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_3/Component_Function_1/N2  ( .A1(\SB4_3/i0_3 ), .A2(
        \SB4_3/i1_7 ), .A3(\SB4_3/i0[8] ), .ZN(
        \SB4_3/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_4/Component_Function_0/N2  ( .A1(\SB4_4/i0[8] ), .A2(
        \SB4_4/i0[7] ), .A3(\SB4_4/i0[6] ), .ZN(
        \SB4_4/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_4/Component_Function_1/N3  ( .A1(\SB4_4/i1_5 ), .A2(
        \SB4_4/i0[6] ), .A3(\SB4_4/i0[9] ), .ZN(
        \SB4_4/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB4_4/Component_Function_1/N1  ( .A1(\SB4_4/i0_3 ), .A2(
        \SB4_4/i1[9] ), .ZN(\SB4_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_4/Component_Function_5/N3  ( .A1(\SB4_4/i1[9] ), .A2(
        \SB4_4/i0_4 ), .A3(\SB4_4/i0_3 ), .ZN(
        \SB4_4/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_5/Component_Function_0/N3  ( .A1(\SB4_5/i0[10] ), .A2(
        \SB4_5/i0_4 ), .A3(\SB4_5/i0_3 ), .ZN(
        \SB4_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_5/Component_Function_0/N2  ( .A1(\SB4_5/i0[8] ), .A2(
        \SB4_5/i0[7] ), .A3(\SB4_5/i0[6] ), .ZN(
        \SB4_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_5/Component_Function_0/N1  ( .A1(\SB4_5/i0[10] ), .A2(
        \SB4_5/i0[9] ), .ZN(\SB4_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_5/Component_Function_1/N4  ( .A1(\SB4_5/i1_7 ), .A2(
        \SB4_5/i0[8] ), .A3(\SB4_5/i0_4 ), .ZN(
        \SB4_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_5/Component_Function_1/N3  ( .A1(\SB4_5/i1_5 ), .A2(
        \SB4_5/i0[6] ), .A3(\SB3_10/buf_output[0] ), .ZN(
        \SB4_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_5/Component_Function_1/N2  ( .A1(\SB4_5/i0_3 ), .A2(
        \SB4_5/i1_7 ), .A3(\SB4_5/i0[8] ), .ZN(
        \SB4_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_5/Component_Function_1/N1  ( .A1(\SB4_5/i0_3 ), .A2(
        \SB4_5/i1[9] ), .ZN(\SB4_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_5/Component_Function_5/N3  ( .A1(\SB4_5/i1[9] ), .A2(
        \SB4_5/i0_4 ), .A3(\SB4_5/i0_3 ), .ZN(
        \SB4_5/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB4_5/Component_Function_5/N1  ( .A1(\SB4_5/i0_0 ), .A2(
        \SB4_5/i3[0] ), .ZN(\SB4_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_6/Component_Function_0/N2  ( .A1(\SB4_6/i0[8] ), .A2(
        \SB4_6/i0[7] ), .A3(\SB4_6/i0[6] ), .ZN(
        \SB4_6/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_6/Component_Function_1/N3  ( .A1(\SB4_6/i1_5 ), .A2(
        \SB4_6/i0[6] ), .A3(\SB4_6/i0[9] ), .ZN(
        \SB4_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_6/Component_Function_5/N4  ( .A1(\SB4_6/i0[9] ), .A2(
        \SB4_6/i0[6] ), .A3(\SB4_6/i0_4 ), .ZN(
        \SB4_6/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_6/Component_Function_5/N1  ( .A1(\SB4_6/i0_0 ), .A2(
        \SB4_6/i3[0] ), .ZN(\SB4_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_7/Component_Function_0/N2  ( .A1(n3965), .A2(\SB4_7/i0[7] ), 
        .A3(\SB4_7/i0[6] ), .ZN(\SB4_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_7/Component_Function_0/N1  ( .A1(\SB3_9/buf_output[3] ), .A2(
        \SB4_7/i0[9] ), .ZN(\SB4_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_7/Component_Function_1/N4  ( .A1(\SB4_7/i1_7 ), .A2(n3965), 
        .A3(\SB4_7/i0_4 ), .ZN(\SB4_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_7/Component_Function_1/N2  ( .A1(\SB4_7/i0_3 ), .A2(
        \SB4_7/i1_7 ), .A3(n3965), .ZN(
        \SB4_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_8/Component_Function_0/N2  ( .A1(\SB4_8/i0[8] ), .A2(
        \SB4_8/i0[7] ), .A3(\SB4_8/i0[6] ), .ZN(
        \SB4_8/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_8/Component_Function_1/N4  ( .A1(\SB4_8/i1_7 ), .A2(
        \SB4_8/i0[8] ), .A3(\SB4_8/i0_4 ), .ZN(
        \SB4_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_8/Component_Function_1/N3  ( .A1(\SB4_8/i1_5 ), .A2(
        \SB4_8/i0[6] ), .A3(\SB3_13/buf_output[0] ), .ZN(
        \SB4_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_8/Component_Function_1/N2  ( .A1(\SB4_8/i0_3 ), .A2(
        \SB4_8/i1_7 ), .A3(\SB4_8/i0[8] ), .ZN(
        \SB4_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_8/Component_Function_5/N1  ( .A1(\SB4_8/i0_0 ), .A2(
        \SB4_8/i3[0] ), .ZN(\SB4_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_9/Component_Function_0/N4  ( .A1(\SB4_9/i0[7] ), .A2(
        \SB4_9/i0_3 ), .A3(\SB4_9/i0_0 ), .ZN(
        \SB4_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_9/Component_Function_0/N3  ( .A1(\SB4_9/i0[10] ), .A2(n6272), 
        .A3(\SB4_9/i0_3 ), .ZN(\SB4_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_9/Component_Function_1/N2  ( .A1(\SB4_9/i0_3 ), .A2(
        \SB4_9/i1_7 ), .A3(n1499), .ZN(
        \SB4_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_9/Component_Function_1/N1  ( .A1(\SB4_9/i0_3 ), .A2(
        \SB4_9/i1[9] ), .ZN(\SB4_9/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB4_9/Component_Function_5/N1  ( .A1(\SB4_9/i0_0 ), .A2(
        \SB4_9/i3[0] ), .ZN(\SB4_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_11/Component_Function_1/N3  ( .A1(\SB4_11/i1_5 ), .A2(
        \SB4_11/i0[6] ), .A3(\SB4_11/i0[9] ), .ZN(
        \SB4_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_11/Component_Function_1/N2  ( .A1(\SB4_11/i0_3 ), .A2(
        \SB4_11/i1_7 ), .A3(\SB4_11/i0[8] ), .ZN(
        \SB4_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_11/Component_Function_1/N1  ( .A1(\SB4_11/i0_3 ), .A2(
        \SB4_11/i1[9] ), .ZN(\SB4_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_11/Component_Function_5/N2  ( .A1(\SB4_11/i0_0 ), .A2(
        \SB4_11/i0[6] ), .A3(\SB4_11/i0[10] ), .ZN(
        \SB4_11/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB4_12/Component_Function_1/N2  ( .A1(\SB4_12/i0_3 ), .A2(
        \SB4_12/i1_7 ), .A3(\SB4_12/i0[8] ), .ZN(
        \SB4_12/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_12/Component_Function_5/N3  ( .A1(\SB4_12/i1[9] ), .A2(
        \SB4_12/i0_4 ), .A3(\SB4_12/i0_3 ), .ZN(
        \SB4_12/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_13/Component_Function_1/N2  ( .A1(\SB4_13/i0_3 ), .A2(
        \SB4_13/i1_7 ), .A3(n1498), .ZN(
        \SB4_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_13/Component_Function_1/N1  ( .A1(\SB4_13/i0_3 ), .A2(
        \SB4_13/i1[9] ), .ZN(\SB4_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_14/Component_Function_0/N3  ( .A1(\SB4_14/i0[10] ), .A2(
        \SB4_14/i0_4 ), .A3(\SB4_14/i0_3 ), .ZN(
        \SB4_14/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB4_14/Component_Function_0/N1  ( .A1(\SB4_14/i0[10] ), .A2(
        \SB4_14/i0[9] ), .ZN(\SB4_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_14/Component_Function_1/N4  ( .A1(\SB4_14/i1_7 ), .A2(
        \SB4_14/i0[8] ), .A3(\SB4_14/i0_4 ), .ZN(
        \SB4_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_14/Component_Function_1/N3  ( .A1(n1495), .A2(\SB4_14/i0[6] ), 
        .A3(\SB4_14/i0[9] ), .ZN(\SB4_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_14/Component_Function_1/N2  ( .A1(\SB4_14/i0_3 ), .A2(
        \SB4_14/i1_7 ), .A3(\SB4_14/i0[8] ), .ZN(
        \SB4_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_14/Component_Function_1/N1  ( .A1(\SB4_14/i0_3 ), .A2(
        \SB4_14/i1[9] ), .ZN(\SB4_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_14/Component_Function_5/N3  ( .A1(\SB4_14/i1[9] ), .A2(
        \SB4_14/i0_4 ), .A3(\SB4_14/i0_3 ), .ZN(
        \SB4_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_14/Component_Function_5/N2  ( .A1(\SB4_14/i0_0 ), .A2(
        \SB4_14/i0[6] ), .A3(\SB4_14/i0[10] ), .ZN(
        \SB4_14/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB4_15/Component_Function_0/N2  ( .A1(n1497), .A2(\SB4_15/i0[7] ), 
        .A3(\SB4_15/i0[6] ), .ZN(\SB4_15/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_15/Component_Function_1/N3  ( .A1(\SB4_15/i1_5 ), .A2(
        \SB4_15/i0[6] ), .A3(\SB4_15/i0[9] ), .ZN(
        \SB4_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_15/Component_Function_1/N2  ( .A1(\SB4_15/i0_3 ), .A2(
        \SB4_15/i1_7 ), .A3(n1497), .ZN(
        \SB4_15/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_15/Component_Function_5/N4  ( .A1(\SB4_15/i0[9] ), .A2(
        \SB4_15/i0[6] ), .A3(\SB4_15/i0_4 ), .ZN(
        \SB4_15/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_15/Component_Function_5/N1  ( .A1(\SB4_15/i0_0 ), .A2(
        \SB4_15/i3[0] ), .ZN(\SB4_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_16/Component_Function_0/N3  ( .A1(\SB4_16/i0[10] ), .A2(
        \SB4_16/i0_4 ), .A3(\SB4_16/i0_3 ), .ZN(
        \SB4_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_16/Component_Function_0/N2  ( .A1(\SB4_16/i0[8] ), .A2(
        \SB4_16/i0[7] ), .A3(\SB4_16/i0[6] ), .ZN(
        \SB4_16/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_17/Component_Function_0/N2  ( .A1(n1493), .A2(\SB4_17/i0[7] ), 
        .A3(\SB4_17/i0[6] ), .ZN(\SB4_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_17/Component_Function_1/N4  ( .A1(\SB4_17/i1_7 ), .A2(n1493), 
        .A3(\SB4_17/i0_4 ), .ZN(\SB4_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_17/Component_Function_1/N3  ( .A1(n3984), .A2(\SB4_17/i0[6] ), 
        .A3(\SB4_17/i0[9] ), .ZN(\SB4_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_17/Component_Function_1/N2  ( .A1(\SB4_17/i0_3 ), .A2(
        \SB4_17/i1_7 ), .A3(n1493), .ZN(
        \SB4_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_17/Component_Function_5/N4  ( .A1(\SB4_17/i0[9] ), .A2(
        \SB4_17/i0[6] ), .A3(\SB4_17/i0_4 ), .ZN(
        \SB4_17/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_17/Component_Function_5/N2  ( .A1(\SB4_17/i0_0 ), .A2(
        \SB4_17/i0[6] ), .A3(\SB4_17/i0[10] ), .ZN(
        \SB4_17/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_17/Component_Function_5/N1  ( .A1(\SB4_17/i0_0 ), .A2(
        \SB4_17/i3[0] ), .ZN(\SB4_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_18/Component_Function_0/N3  ( .A1(\SB4_18/i0[10] ), .A2(
        \SB4_18/i0_4 ), .A3(\SB4_18/i0_3 ), .ZN(
        \SB4_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_18/Component_Function_0/N2  ( .A1(\SB4_18/i0[8] ), .A2(
        \SB4_18/i0[7] ), .A3(\SB4_18/i0[6] ), .ZN(
        \SB4_18/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_18/Component_Function_1/N4  ( .A1(\SB4_18/i1_7 ), .A2(
        \SB4_18/i0[8] ), .A3(\SB4_18/i0_4 ), .ZN(
        \SB4_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_18/Component_Function_1/N2  ( .A1(\SB4_18/i0_3 ), .A2(
        \SB4_18/i1_7 ), .A3(\SB4_18/i0[8] ), .ZN(
        \SB4_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_18/Component_Function_5/N4  ( .A1(\SB4_18/i0[9] ), .A2(
        \SB4_18/i0[6] ), .A3(\SB4_18/i0_4 ), .ZN(
        \SB4_18/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_18/Component_Function_5/N1  ( .A1(\SB4_18/i0_0 ), .A2(
        \SB4_18/i3[0] ), .ZN(\SB4_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_19/Component_Function_0/N3  ( .A1(\SB4_19/i0[10] ), .A2(
        \SB4_19/i0_4 ), .A3(\SB4_19/i0_3 ), .ZN(
        \SB4_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_1/N4  ( .A1(\SB4_19/i1_7 ), .A2(
        \SB4_19/i0[8] ), .A3(\SB4_19/i0_4 ), .ZN(
        \SB4_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_19/Component_Function_5/N2  ( .A1(\SB4_19/i0_0 ), .A2(
        \SB4_19/i0[6] ), .A3(\SB4_19/i0[10] ), .ZN(
        \SB4_19/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_19/Component_Function_5/N1  ( .A1(\SB4_19/i0_0 ), .A2(
        \SB4_19/i3[0] ), .ZN(\SB4_19/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB4_20/Component_Function_0/N1  ( .A1(\SB4_20/i0[10] ), .A2(
        \SB4_20/i0[9] ), .ZN(\SB4_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_20/Component_Function_1/N4  ( .A1(\SB4_20/i1_7 ), .A2(
        \SB4_20/i0[8] ), .A3(\SB4_20/i0_4 ), .ZN(
        \SB4_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_20/Component_Function_1/N2  ( .A1(\SB4_20/i0_3 ), .A2(
        \SB4_20/i1_7 ), .A3(\SB4_20/i0[8] ), .ZN(
        \SB4_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_20/Component_Function_5/N4  ( .A1(\SB4_20/i0[9] ), .A2(
        \SB4_20/i0[6] ), .A3(\SB3_21/buf_output[4] ), .ZN(
        \SB4_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_20/Component_Function_5/N3  ( .A1(\SB4_20/i1[9] ), .A2(
        \SB4_20/i0_4 ), .A3(\SB4_20/i0_3 ), .ZN(
        \SB4_20/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_21/Component_Function_5/N4  ( .A1(\SB4_21/i0[9] ), .A2(
        \SB4_21/i0[6] ), .A3(\SB4_21/i0_4 ), .ZN(
        \SB4_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_22/Component_Function_0/N3  ( .A1(\SB4_22/i0[10] ), .A2(
        \SB4_22/i0_4 ), .A3(\SB4_22/i0_3 ), .ZN(
        \SB4_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_22/Component_Function_0/N2  ( .A1(\SB4_22/i0[8] ), .A2(
        \SB4_22/i0[7] ), .A3(\SB4_22/i0[6] ), .ZN(
        \SB4_22/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_22/Component_Function_1/N4  ( .A1(\SB4_22/i1_7 ), .A2(
        \SB4_22/i0[8] ), .A3(\SB4_22/i0_4 ), .ZN(
        \SB4_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_22/Component_Function_1/N2  ( .A1(\SB4_22/i0_3 ), .A2(
        \SB4_22/i1_7 ), .A3(\SB4_22/i0[8] ), .ZN(
        \SB4_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_22/Component_Function_1/N1  ( .A1(\SB4_22/i0_3 ), .A2(
        \SB4_22/i1[9] ), .ZN(\SB4_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_23/Component_Function_0/N3  ( .A1(\SB4_23/i0[10] ), .A2(
        \SB4_23/i0_4 ), .A3(\SB4_23/i0_3 ), .ZN(
        \SB4_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_23/Component_Function_0/N2  ( .A1(n3974), .A2(\SB4_23/i0[7] ), 
        .A3(\SB3_27/buf_output[1] ), .ZN(
        \SB4_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_23/Component_Function_1/N1  ( .A1(\SB4_23/i0_3 ), .A2(
        \SB4_23/i1[9] ), .ZN(\SB4_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_24/Component_Function_1/N3  ( .A1(\SB4_24/i1_5 ), .A2(
        \SB4_24/i0[6] ), .A3(\SB4_24/i0[9] ), .ZN(
        \SB4_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_24/Component_Function_1/N2  ( .A1(\SB4_24/i0_3 ), .A2(
        \SB4_24/i1_7 ), .A3(n1494), .ZN(
        \SB4_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_24/Component_Function_1/N1  ( .A1(\SB4_24/i0_3 ), .A2(
        \SB4_24/i1[9] ), .ZN(\SB4_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_24/Component_Function_5/N2  ( .A1(\SB4_24/i0_0 ), .A2(
        \SB4_24/i0[6] ), .A3(\SB3_26/buf_output[3] ), .ZN(
        \SB4_24/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB4_25/Component_Function_0/N4  ( .A1(\SB4_25/i0[7] ), .A2(
        \SB4_25/i0_3 ), .A3(\SB4_25/i0_0 ), .ZN(
        \SB4_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_0/N3  ( .A1(\SB4_25/i0[10] ), .A2(
        \SB4_25/i0_4 ), .A3(\SB4_25/i0_3 ), .ZN(
        \SB4_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_25/Component_Function_0/N2  ( .A1(\SB4_25/i0[8] ), .A2(
        \SB4_25/i0[7] ), .A3(\SB4_25/i0[6] ), .ZN(
        \SB4_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_25/Component_Function_1/N4  ( .A1(\SB4_25/i1_7 ), .A2(
        \SB4_25/i0[8] ), .A3(\SB4_25/i0_4 ), .ZN(
        \SB4_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_5/N2  ( .A1(\SB4_25/i0_0 ), .A2(
        \SB4_25/i0[6] ), .A3(\SB4_25/i0[10] ), .ZN(
        \SB4_25/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_25/Component_Function_5/N1  ( .A1(\SB4_25/i0_0 ), .A2(n5438), 
        .ZN(\SB4_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_26/Component_Function_0/N3  ( .A1(\SB4_26/i0[10] ), .A2(
        \SB4_26/i0_4 ), .A3(\SB4_26/i0_3 ), .ZN(
        \SB4_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_26/Component_Function_1/N4  ( .A1(\SB4_26/i1_7 ), .A2(n3989), 
        .A3(\SB3_27/buf_output[4] ), .ZN(
        \SB4_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_26/Component_Function_5/N4  ( .A1(\SB4_26/i0[9] ), .A2(
        \SB4_26/i0[6] ), .A3(\SB4_26/i0_4 ), .ZN(
        \SB4_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_26/Component_Function_5/N3  ( .A1(n573), .A2(\SB4_26/i0_4 ), 
        .A3(\SB4_26/i0_3 ), .ZN(\SB4_26/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB4_26/Component_Function_5/N1  ( .A1(\SB3_29/buf_output[2] ), 
        .A2(\SB4_26/i3[0] ), .ZN(\SB4_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_0/N3  ( .A1(\SB4_27/i0[10] ), .A2(
        \SB4_27/i0_4 ), .A3(\SB4_27/i0_3 ), .ZN(
        \SB4_27/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB4_27/Component_Function_0/N1  ( .A1(\SB4_27/i0[10] ), .A2(
        \SB4_27/i0[9] ), .ZN(\SB4_27/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB4_27/Component_Function_1/N1  ( .A1(\SB4_27/i0_3 ), .A2(
        \SB4_27/i1[9] ), .ZN(\SB4_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_5/N4  ( .A1(\SB4_27/i0[9] ), .A2(
        \SB4_27/i0[6] ), .A3(\SB4_27/i0_4 ), .ZN(
        \SB4_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_27/Component_Function_5/N3  ( .A1(\SB4_27/i1[9] ), .A2(
        \SB4_27/i0_4 ), .A3(\SB4_27/i0_3 ), .ZN(
        \SB4_27/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_27/Component_Function_5/N2  ( .A1(\SB4_27/i0_0 ), .A2(
        \SB4_27/i0[6] ), .A3(\SB4_27/i0[10] ), .ZN(
        \SB4_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB4_28/Component_Function_1/N4  ( .A1(\SB4_28/i1_7 ), .A2(
        \SB4_28/i0[8] ), .A3(\SB4_28/i0_4 ), .ZN(
        \SB4_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_28/Component_Function_1/N2  ( .A1(\SB4_28/i0_3 ), .A2(
        \SB4_28/i1_7 ), .A3(\SB4_28/i0[8] ), .ZN(
        \SB4_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_29/Component_Function_1/N3  ( .A1(\SB4_29/i1_5 ), .A2(
        \SB4_29/i0[6] ), .A3(\SB4_29/i0[9] ), .ZN(
        \SB4_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_29/Component_Function_1/N2  ( .A1(\SB4_29/i0_3 ), .A2(
        \SB4_29/i1_7 ), .A3(\SB4_29/i0[8] ), .ZN(
        \SB4_29/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_29/Component_Function_5/N3  ( .A1(\SB4_29/i1[9] ), .A2(
        \SB4_29/i0_4 ), .A3(\SB4_29/i0_3 ), .ZN(
        \SB4_29/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB4_29/Component_Function_5/N1  ( .A1(\SB4_29/i0_0 ), .A2(
        \SB4_29/i3[0] ), .ZN(\SB4_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_30/Component_Function_1/N4  ( .A1(\SB4_30/i1_7 ), .A2(
        \SB4_30/i0[8] ), .A3(\SB4_30/i0_4 ), .ZN(
        \SB4_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_30/Component_Function_1/N2  ( .A1(\SB4_30/i0_3 ), .A2(
        \SB4_30/i1_7 ), .A3(\SB4_30/i0[8] ), .ZN(
        \SB4_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_30/Component_Function_1/N1  ( .A1(\SB4_30/i0_3 ), .A2(n3973), 
        .ZN(\SB4_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_30/Component_Function_5/N2  ( .A1(n5427), .A2(\SB4_30/i0[6] ), 
        .A3(\SB4_30/i0[10] ), .ZN(\SB4_30/Component_Function_5/NAND4_in[1] )
         );
  NAND2_X1 \SB4_30/Component_Function_5/N1  ( .A1(n5427), .A2(\SB4_30/i3[0] ), 
        .ZN(\SB4_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_31/Component_Function_1/N4  ( .A1(\SB4_31/i1_7 ), .A2(
        \SB4_31/i0[8] ), .A3(\SB4_31/i0_4 ), .ZN(
        \SB4_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_31/Component_Function_1/N3  ( .A1(\SB4_31/i1_5 ), .A2(
        \SB4_31/i0[6] ), .A3(\SB4_31/i0[9] ), .ZN(
        \SB4_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_31/Component_Function_1/N2  ( .A1(\SB4_31/i0_3 ), .A2(
        \SB4_31/i1_7 ), .A3(\SB4_31/i0[8] ), .ZN(
        \SB4_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_31/Component_Function_1/N1  ( .A1(\SB4_31/i0_3 ), .A2(
        \SB4_31/i1[9] ), .ZN(\SB4_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_31/Component_Function_5/N2  ( .A1(\SB4_31/i0_0 ), .A2(
        \SB4_31/i0[6] ), .A3(\SB4_31/i0[10] ), .ZN(
        \SB4_31/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_31/Component_Function_5/N1  ( .A1(\SB4_31/i0_0 ), .A2(
        \SB4_31/i3[0] ), .ZN(\SB4_31/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_0_0/BUF_5  ( .I(\SB1_0_0/buf_output[5] ), .Z(\SB2_0_0/i0_3 ) );
  BUF_X4 \SB2_0_26/BUF_5  ( .I(\RI3[0][35] ), .Z(\SB2_0_26/i0_3 ) );
  BUF_X4 \SB1_1_0/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[191] ), .Z(
        \SB1_1_0/i0_3 ) );
  BUF_X4 \SB1_1_5/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[161] ), .Z(
        \SB1_1_5/i0_3 ) );
  BUF_X4 \SB1_1_8/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[143] ), .Z(
        \SB1_1_8/i0_3 ) );
  BUF_X4 \SB1_1_10/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[131] ), .Z(
        \SB1_1_10/i0_3 ) );
  BUF_X4 \SB1_1_13/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[113] ), .Z(
        \SB1_1_13/i0_3 ) );
  BUF_X4 \SB1_1_14/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[107] ), .Z(
        \SB1_1_14/i0_3 ) );
  BUF_X4 \SB1_1_16/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[95] ), .Z(
        \SB1_1_16/i0_3 ) );
  BUF_X4 \SB1_1_17/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[89] ), .Z(
        \SB1_1_17/i0_3 ) );
  BUF_X4 \SB1_1_19/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[77] ), .Z(
        \SB1_1_19/i0_3 ) );
  BUF_X4 \SB1_1_25/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[41] ), .Z(
        \SB1_1_25/i0_3 ) );
  BUF_X4 \SB1_1_27/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[29] ), .Z(
        \SB1_1_27/i0_3 ) );
  BUF_X4 \SB2_1_0/BUF_5  ( .I(\SB1_1_0/buf_output[5] ), .Z(\SB2_1_0/i0_3 ) );
  BUF_X4 \SB2_1_3/BUF_5  ( .I(\SB1_1_3/buf_output[5] ), .Z(\SB2_1_3/i0_3 ) );
  BUF_X4 \SB2_1_5/BUF_5  ( .I(\SB1_1_5/buf_output[5] ), .Z(\SB2_1_5/i0_3 ) );
  BUF_X4 \SB2_1_6/BUF_5  ( .I(\SB1_1_6/buf_output[5] ), .Z(\SB2_1_6/i0_3 ) );
  BUF_X4 \SB2_1_14/BUF_5  ( .I(\SB1_1_14/buf_output[5] ), .Z(\SB2_1_14/i0_3 )
         );
  BUF_X4 \SB2_1_18/BUF_5  ( .I(\SB1_1_18/buf_output[5] ), .Z(\SB2_1_18/i0_3 )
         );
  BUF_X4 \SB2_1_19/BUF_5  ( .I(\SB1_1_19/buf_output[5] ), .Z(\SB2_1_19/i0_3 )
         );
  BUF_X4 \SB2_1_25/BUF_5  ( .I(\SB1_1_25/buf_output[5] ), .Z(\SB2_1_25/i0_3 )
         );
  BUF_X4 \SB1_2_9/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[137] ), .Z(
        \SB1_2_9/i0_3 ) );
  BUF_X4 \SB1_2_17/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[89] ), .Z(
        \SB1_2_17/i0_3 ) );
  BUF_X4 \SB1_2_19/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[77] ), .Z(
        \SB1_2_19/i0_3 ) );
  BUF_X4 \SB1_2_20/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[71] ), .Z(
        \SB1_2_20/i0_3 ) );
  BUF_X4 \SB1_2_24/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[47] ), .Z(
        \SB1_2_24/i0_3 ) );
  BUF_X4 \SB1_2_27/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[29] ), .Z(
        \SB1_2_27/i0_3 ) );
  BUF_X4 \SB2_2_1/BUF_5  ( .I(\SB1_2_1/buf_output[5] ), .Z(\SB2_2_1/i0_3 ) );
  BUF_X4 \SB2_2_6/BUF_5  ( .I(\SB1_2_6/buf_output[5] ), .Z(\SB2_2_6/i0_3 ) );
  BUF_X4 \SB2_2_20/BUF_5  ( .I(\SB1_2_20/buf_output[5] ), .Z(\SB2_2_20/i0_3 )
         );
  BUF_X4 \SB2_2_24/BUF_5  ( .I(\SB1_2_24/buf_output[5] ), .Z(\SB2_2_24/i0_3 )
         );
  BUF_X4 \SB2_2_25/BUF_5  ( .I(\SB1_2_25/buf_output[5] ), .Z(\SB2_2_25/i0_3 )
         );
  BUF_X4 \SB2_2_27/BUF_5  ( .I(\SB1_2_27/buf_output[5] ), .Z(\SB2_2_27/i0_3 )
         );
  BUF_X4 \SB1_3_1/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[185] ), .Z(
        \SB1_3_1/i0_3 ) );
  BUF_X4 \SB1_3_8/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[143] ), .Z(
        \SB1_3_8/i0_3 ) );
  BUF_X4 \SB1_3_11/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[125] ), .Z(
        \SB1_3_11/i0_3 ) );
  BUF_X4 \SB1_3_17/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[89] ), .Z(
        \SB1_3_17/i0_3 ) );
  BUF_X4 \SB1_3_20/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[71] ), .Z(
        \SB1_3_20/i0_3 ) );
  BUF_X4 \SB1_3_23/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[53] ), .Z(
        \SB1_3_23/i0_3 ) );
  BUF_X4 \SB1_3_25/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[41] ), .Z(
        \SB1_3_25/i0_3 ) );
  BUF_X4 \SB2_3_0/BUF_5  ( .I(\SB1_3_0/buf_output[5] ), .Z(\SB2_3_0/i0_3 ) );
  BUF_X4 \SB2_3_11/BUF_5  ( .I(\SB1_3_11/buf_output[5] ), .Z(\SB2_3_11/i0_3 )
         );
  BUF_X4 \SB2_3_18/BUF_5  ( .I(\SB1_3_18/buf_output[5] ), .Z(\SB2_3_18/i0_3 )
         );
  BUF_X4 \SB2_3_19/BUF_5  ( .I(\SB1_3_19/buf_output[5] ), .Z(\SB2_3_19/i0_3 )
         );
  BUF_X4 \SB2_3_22/BUF_5  ( .I(\SB1_3_22/buf_output[5] ), .Z(\SB2_3_22/i0_3 )
         );
  BUF_X4 \SB1_4_5/BUF_5  ( .I(\MC_ARK_ARC_1_3/buf_output[161] ), .Z(
        \SB1_4_5/i0_3 ) );
  BUF_X4 \SB1_4_26/BUF_5  ( .I(\MC_ARK_ARC_1_3/buf_output[35] ), .Z(
        \SB1_4_26/i0_3 ) );
  BUF_X4 \SB2_4_1/BUF_5  ( .I(\SB1_4_1/buf_output[5] ), .Z(\SB2_4_1/i0_3 ) );
  BUF_X4 \SB2_4_2/BUF_5  ( .I(\SB1_4_2/buf_output[5] ), .Z(\SB2_4_2/i0_3 ) );
  BUF_X4 \SB2_4_5/BUF_5  ( .I(\SB1_4_5/buf_output[5] ), .Z(\SB2_4_5/i0_3 ) );
  BUF_X4 \SB3_27/BUF_5  ( .I(\MC_ARK_ARC_1_4/buf_output[29] ), .Z(
        \SB3_27/i0_3 ) );
  BUF_X4 \SB4_13/BUF_5  ( .I(\SB3_13/buf_output[5] ), .Z(\SB4_13/i0_3 ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_21  ( .I(\SB2_3_30/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[21] ) );
  INV_X2 \SB2_3_2/INV_3  ( .I(\SB1_3_4/buf_output[3] ), .ZN(\SB2_3_2/i0[8] )
         );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_12  ( .I(\SB2_4_2/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[12] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_113  ( .I(\SB2_0_13/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[113] ) );
  INV_X2 \SB2_3_16/INV_3  ( .I(\SB1_3_18/buf_output[3] ), .ZN(\SB2_3_16/i0[8] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_19  ( .I(\SB2_3_0/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[19] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_115  ( .I(\SB2_2_16/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[115] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_125  ( .I(\SB2_1_11/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[125] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_55  ( .I(\SB2_2_26/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[55] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_7  ( .I(\SB2_2_2/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[7] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_43  ( .I(\SB2_4_28/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[43] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_54  ( .I(\SB2_4_27/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[54] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_173  ( .I(\RI5[0][173] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[173] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_121  ( .I(\SB2_2_15/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[121] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_53  ( .I(\SB2_3_23/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[53] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_143  ( .I(\SB2_3_8/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[143] ) );
  INV_X2 \SB4_11/INV_3  ( .I(\SB3_13/buf_output[3] ), .ZN(\SB4_11/i0[8] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_155  ( .I(\SB2_3_6/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[155] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_151  ( .I(\SB2_1_10/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[151] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_83  ( .I(\SB2_1_18/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[83] ) );
  NAND3_X1 \SB1_4_10/Component_Function_1/N2  ( .A1(\RI1[4][131] ), .A2(
        \SB1_4_10/i1_7 ), .A3(\SB1_4_10/i0[8] ), .ZN(
        \SB1_4_10/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_71  ( .I(\SB2_3_20/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[71] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_179  ( .I(\SB2_2_2/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[179] ) );
  INV_X2 \SB1_4_20/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[69] ), .ZN(
        \SB1_4_20/i0[8] ) );
  INV_X2 \SB1_4_22/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[57] ), .ZN(
        \SB1_4_22/i0[8] ) );
  INV_X2 \SB1_4_0/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[189] ), .ZN(
        \SB1_4_0/i0[8] ) );
  INV_X2 \SB1_3_15/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[99] ), .ZN(
        \SB1_3_15/i0[8] ) );
  INV_X2 \SB1_4_17/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[87] ), .ZN(
        \SB1_4_17/i0[8] ) );
  NAND3_X1 \SB1_3_10/Component_Function_4/N4  ( .A1(\SB1_3_10/i1[9] ), .A2(
        \SB1_3_10/i1_5 ), .A3(\SB1_3_10/i0_4 ), .ZN(
        \SB1_3_10/Component_Function_4/NAND4_in[3] ) );
  INV_X2 \SB1_4_13/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[111] ), .ZN(
        \SB1_4_13/i0[8] ) );
  INV_X2 \SB3_14/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[104] ), .ZN(
        \SB3_14/i1[9] ) );
  INV_X2 \SB3_28/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[20] ), .ZN(
        \SB3_28/i1[9] ) );
  INV_X2 \SB1_4_30/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[9] ), .ZN(
        \SB1_4_30/i0[8] ) );
  INV_X2 \SB1_3_6/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[153] ), .ZN(
        \SB1_3_6/i0[8] ) );
  INV_X2 \SB1_4_31/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[3] ), .ZN(
        \SB1_4_31/i0[8] ) );
  INV_X2 \SB1_3_14/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[104] ), .ZN(
        \SB1_3_14/i1[9] ) );
  INV_X2 \SB1_4_3/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[171] ), .ZN(
        \SB1_4_3/i0[8] ) );
  INV_X2 \SB1_4_28/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[21] ), .ZN(
        \SB1_4_28/i0[8] ) );
  INV_X2 \SB1_4_20/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[68] ), .ZN(
        \SB1_4_20/i1[9] ) );
  INV_X2 \SB2_4_30/INV_2  ( .I(\SB1_4_1/buf_output[2] ), .ZN(\SB2_4_30/i1[9] )
         );
  INV_X2 \SB1_3_17/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[87] ), .ZN(
        \SB1_3_17/i0[8] ) );
  INV_X2 \SB2_1_3/INV_3  ( .I(\SB1_1_5/buf_output[3] ), .ZN(\SB2_1_3/i0[8] )
         );
  CLKBUF_X4 \SB2_2_30/BUF_2  ( .I(\SB1_2_1/buf_output[2] ), .Z(\SB2_2_30/i0_0 ) );
  INV_X2 \SB1_3_29/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[15] ), .ZN(
        \SB1_3_29/i0[8] ) );
  INV_X2 \SB2_3_2/INV_2  ( .I(\SB1_3_5/buf_output[2] ), .ZN(\SB2_3_2/i1[9] )
         );
  INV_X2 \SB1_2_4/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[165] ), .ZN(
        \SB1_2_4/i0[8] ) );
  CLKBUF_X4 \SB2_1_0/BUF_2  ( .I(\SB1_1_3/buf_output[2] ), .Z(\SB2_1_0/i0_0 )
         );
  INV_X2 \SB1_3_9/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[134] ), .ZN(
        \SB1_3_9/i1[9] ) );
  INV_X2 \SB1_1_4/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[165] ), .ZN(
        \SB1_1_4/i0[8] ) );
  INV_X2 \SB3_17/INV_3  ( .I(\MC_ARK_ARC_1_4/buf_output[87] ), .ZN(
        \SB3_17/i0[8] ) );
  NAND3_X1 \SB1_1_15/Component_Function_3/N2  ( .A1(\SB1_1_15/i0_0 ), .A2(
        \SB1_1_15/i0_3 ), .A3(\SB1_1_15/i0_4 ), .ZN(
        \SB1_1_15/Component_Function_3/NAND4_in[1] ) );
  INV_X2 \SB3_23/INV_3  ( .I(\MC_ARK_ARC_1_4/buf_output[51] ), .ZN(
        \SB3_23/i0[8] ) );
  INV_X2 \SB1_3_14/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[105] ), .ZN(
        \SB1_3_14/i0[8] ) );
  INV_X2 \SB1_3_22/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[56] ), .ZN(
        \SB1_3_22/i1[9] ) );
  INV_X1 \SB1_0_3/INV_5  ( .I(n409), .ZN(\SB1_0_3/i1_5 ) );
  INV_X2 \SB1_4_30/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[8] ), .ZN(
        \SB1_4_30/i1[9] ) );
  INV_X2 \SB1_3_22/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[57] ), .ZN(
        \SB1_3_22/i0[8] ) );
  INV_X2 \SB1_1_5/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[158] ), .ZN(
        \SB1_1_5/i1[9] ) );
  INV_X2 \SB1_1_30/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[9] ), .ZN(
        \SB1_1_30/i0[8] ) );
  NAND3_X1 \SB2_1_14/Component_Function_0/N4  ( .A1(\SB2_1_14/i0[7] ), .A2(
        \SB2_1_14/i0_3 ), .A3(\SB2_1_14/i0_0 ), .ZN(
        \SB2_1_14/Component_Function_0/NAND4_in[3] ) );
  INV_X2 \SB1_3_2/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[176] ), .ZN(
        \SB1_3_2/i1[9] ) );
  INV_X2 \SB1_3_17/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[86] ), .ZN(
        \SB1_3_17/i1[9] ) );
  INV_X2 \SB1_3_9/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[135] ), .ZN(
        \SB1_3_9/i0[8] ) );
  INV_X2 \SB1_1_16/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[93] ), .ZN(
        \SB1_1_16/i0[8] ) );
  INV_X2 \SB3_26/INV_3  ( .I(\MC_ARK_ARC_1_4/buf_output[33] ), .ZN(
        \SB3_26/i0[8] ) );
  INV_X2 \SB1_2_16/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[93] ), .ZN(
        \SB1_2_16/i0[8] ) );
  INV_X2 \SB1_2_8/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[140] ), .ZN(
        \SB1_2_8/i1[9] ) );
  INV_X2 \SB1_4_22/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[56] ), .ZN(
        \SB1_4_22/i1[9] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_111_0  ( .I(Key[103]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[111] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_2/BUF_79_0  ( .I(n128), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[79] ) );
  BUF_X4 \SB1_0_12/BUF_5  ( .I(n400), .Z(\SB1_0_12/i0_3 ) );
  BUF_X4 \SB2_1_21/BUF_4  ( .I(\SB1_1_22/buf_output[4] ), .Z(\SB2_1_21/i0_4 )
         );
  BUF_X4 \SB1_3_5/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[160] ), .Z(
        \SB1_3_5/i0_4 ) );
  BUF_X4 \SB2_1_24/BUF_4  ( .I(\SB1_1_25/buf_output[4] ), .Z(\SB2_1_24/i0_4 )
         );
  BUF_X4 \SB1_0_24/BUF_5  ( .I(n388), .Z(\SB1_0_24/i0_3 ) );
  BUF_X4 \SB1_2_4/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[166] ), .Z(
        \SB1_2_4/i0_4 ) );
  BUF_X4 \SB2_0_31/BUF_5  ( .I(\RI3[0][5] ), .Z(\SB2_0_31/i0_3 ) );
  BUF_X4 \SB2_1_27/BUF_4  ( .I(\SB1_1_28/buf_output[4] ), .Z(\SB2_1_27/i0_4 )
         );
  BUF_X4 \SB1_0_30/BUF_5  ( .I(n382), .Z(\SB1_0_30/i0_3 ) );
  BUF_X4 \SB1_3_21/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[64] ), .Z(
        \SB1_3_21/i0_4 ) );
  BUF_X4 \SB2_0_6/BUF_5  ( .I(\RI3[0][155] ), .Z(\SB2_0_6/i0_3 ) );
  BUF_X4 \SB1_3_29/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[16] ), .Z(
        \SB1_3_29/i0_4 ) );
  NAND4_X2 \SB1_2_25/Component_Function_0/N5  ( .A1(
        \SB1_2_25/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_25/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_25/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_25/buf_output[0] ) );
  BUF_X4 \SB1_0_17/BUF_5  ( .I(n395), .Z(\SB1_0_17/i0_3 ) );
  NAND4_X2 \SB3_8/Component_Function_4/N5  ( .A1(
        \SB3_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_8/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_8/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_8/buf_output[4] )
         );
  BUF_X4 \SB1_4_27/BUF_5  ( .I(\MC_ARK_ARC_1_3/buf_output[29] ), .Z(
        \SB1_4_27/i0_3 ) );
  BUF_X4 \SB1_1_8/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[142] ), .Z(
        \SB1_1_8/i0_4 ) );
  BUF_X4 \SB1_2_26/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[35] ), .Z(
        \SB1_2_26/i0_3 ) );
  INV_X2 \SB1_2_10/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[131] ), .ZN(
        \SB1_2_10/i1_5 ) );
  BUF_X4 \SB2_3_27/BUF_2  ( .I(\SB1_3_30/buf_output[2] ), .Z(\SB2_3_27/i0_0 )
         );
  INV_X2 \SB2_2_13/INV_2  ( .I(\SB1_2_16/buf_output[2] ), .ZN(\SB2_2_13/i1[9] ) );
  BUF_X4 \SB2_0_18/BUF_3  ( .I(\RI3[0][81] ), .Z(\SB2_0_18/i0[10] ) );
  BUF_X4 \SB1_3_31/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[4] ), .Z(
        \SB1_3_31/i0_4 ) );
  BUF_X4 \SB1_2_27/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[28] ), .Z(
        \SB1_2_27/i0_4 ) );
  INV_X2 \SB1_1_15/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[99] ), .ZN(
        \SB1_1_15/i0[8] ) );
  INV_X2 \SB1_3_4/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[164] ), .ZN(
        \SB1_3_4/i1[9] ) );
  INV_X2 \SB1_1_7/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[147] ), .ZN(
        \SB1_1_7/i0[8] ) );
  INV_X2 \SB2_2_1/INV_2  ( .I(\SB1_2_4/buf_output[2] ), .ZN(\SB2_2_1/i1[9] )
         );
  NAND4_X2 \SB1_3_18/Component_Function_0/N5  ( .A1(
        \SB1_3_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_18/buf_output[0] ) );
  INV_X2 \SB1_0_26/INV_3  ( .I(n327), .ZN(\SB1_0_26/i0[8] ) );
  BUF_X4 \SB1_3_2/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[179] ), .Z(
        \SB1_3_2/i0_3 ) );
  INV_X2 \SB1_2_23/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[53] ), .ZN(
        \SB1_2_23/i1_5 ) );
  INV_X2 \SB2_2_17/INV_2  ( .I(\SB1_2_20/buf_output[2] ), .ZN(\SB2_2_17/i1[9] ) );
  BUF_X4 \SB1_4_19/BUF_5  ( .I(\MC_ARK_ARC_1_3/buf_output[77] ), .Z(
        \SB1_4_19/i0_3 ) );
  INV_X2 \SB1_3_21/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[62] ), .ZN(
        \SB1_3_21/i1[9] ) );
  INV_X2 \SB1_2_20/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[68] ), .ZN(
        \SB1_2_20/i1[9] ) );
  INV_X2 \SB2_4_18/INV_3  ( .I(\SB1_4_20/buf_output[3] ), .ZN(\SB2_4_18/i0[8] ) );
  INV_X2 \SB1_3_1/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[183] ), .ZN(
        \SB1_3_1/i0[8] ) );
  NAND4_X2 \SB1_4_26/Component_Function_0/N5  ( .A1(
        \SB1_4_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_4_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_26/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_4_26/buf_output[0] ) );
  INV_X2 \SB1_3_19/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[75] ), .ZN(
        \SB1_3_19/i0[8] ) );
  BUF_X4 \SB2_1_17/BUF_5  ( .I(\SB1_1_17/buf_output[5] ), .Z(\SB2_1_17/i0_3 )
         );
  INV_X2 \SB1_1_0/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[189] ), .ZN(
        \SB1_1_0/i0[8] ) );
  BUF_X4 \SB2_1_31/BUF_5  ( .I(\SB1_1_31/buf_output[5] ), .Z(\SB2_1_31/i0_3 )
         );
  INV_X2 \SB1_3_29/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[14] ), .ZN(
        \SB1_3_29/i1[9] ) );
  INV_X2 \SB2_4_10/INV_2  ( .I(\SB1_4_13/buf_output[2] ), .ZN(\SB2_4_10/i1[9] ) );
  BUF_X4 \SB1_2_26/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[32] ), .Z(
        \SB1_2_26/i0_0 ) );
  INV_X2 \SB2_0_14/INV_2  ( .I(\SB1_0_17/buf_output[2] ), .ZN(\SB2_0_14/i1[9] ) );
  INV_X2 \SB2_2_14/INV_3  ( .I(\SB1_2_16/buf_output[3] ), .ZN(\SB2_2_14/i0[8] ) );
  NAND4_X2 \SB1_3_9/Component_Function_0/N5  ( .A1(
        \SB1_3_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_9/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_9/buf_output[0] ) );
  INV_X2 \SB3_18/INV_2  ( .I(\RI1[5][80] ), .ZN(\SB3_18/i1[9] ) );
  BUF_X4 \SB1_2_30/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[11] ), .Z(
        \SB1_2_30/i0_3 ) );
  BUF_X4 \SB2_3_24/BUF_5  ( .I(\SB1_3_24/buf_output[5] ), .Z(\SB2_3_24/i0_3 )
         );
  INV_X2 \SB1_1_21/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[63] ), .ZN(
        \SB1_1_21/i0[8] ) );
  INV_X2 \SB1_2_21/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[62] ), .ZN(
        \SB1_2_21/i1[9] ) );
  INV_X2 \SB2_0_19/INV_2  ( .I(\SB1_0_22/buf_output[2] ), .ZN(\SB2_0_19/i1[9] ) );
  BUF_X4 \SB1_3_13/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[113] ), .Z(
        \SB1_3_13/i0_3 ) );
  NAND4_X2 \SB1_3_24/Component_Function_0/N5  ( .A1(
        \SB1_3_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_24/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_24/buf_output[0] ) );
  INV_X2 \SB1_2_17/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[86] ), .ZN(
        \SB1_2_17/i1[9] ) );
  NAND3_X2 \SB1_1_30/Component_Function_2/N3  ( .A1(\SB1_1_30/i0_3 ), .A2(
        \SB1_1_30/i0[8] ), .A3(\SB1_1_30/i0[9] ), .ZN(
        \SB1_1_30/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB1_2_30/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[8] ), .ZN(
        \SB1_2_30/i1[9] ) );
  INV_X2 \SB1_2_7/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[146] ), .ZN(
        \SB1_2_7/i1[9] ) );
  INV_X2 \SB1_3_18/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[80] ), .ZN(
        \SB1_3_18/i1[9] ) );
  INV_X2 \SB1_4_6/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[152] ), .ZN(
        \SB1_4_6/i1[9] ) );
  INV_X2 \SB1_1_8/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[141] ), .ZN(
        \SB1_1_8/i0[8] ) );
  INV_X2 \SB1_0_17/INV_2  ( .I(n282), .ZN(\SB1_0_17/i1[9] ) );
  INV_X2 \SB2_1_28/INV_2  ( .I(\SB1_1_31/buf_output[2] ), .ZN(\SB2_1_28/i1[9] ) );
  INV_X2 \SB1_2_31/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[2] ), .ZN(
        \SB1_2_31/i1[9] ) );
  INV_X2 \SB1_3_23/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[50] ), .ZN(
        \SB1_3_23/i1[9] ) );
  INV_X2 \SB2_1_13/INV_2  ( .I(\SB1_1_16/buf_output[2] ), .ZN(\SB2_1_13/i1[9] ) );
  BUF_X4 \SB2_2_28/BUF_5  ( .I(\SB1_2_28/buf_output[5] ), .Z(\SB2_2_28/i0_3 )
         );
  INV_X2 \SB1_4_26/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[33] ), .ZN(
        \SB1_4_26/i0[8] ) );
  INV_X2 \SB1_1_24/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[44] ), .ZN(
        \SB1_1_24/i1[9] ) );
  INV_X2 \SB1_3_1/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[182] ), .ZN(
        \SB1_3_1/i1[9] ) );
  INV_X2 \SB1_2_1/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[183] ), .ZN(
        \SB1_2_1/i0[8] ) );
  BUF_X4 \SB2_2_8/BUF_5  ( .I(\SB1_2_8/buf_output[5] ), .Z(\SB2_2_8/i0_3 ) );
  INV_X2 \SB1_2_6/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[155] ), .ZN(
        \SB1_2_6/i1_5 ) );
  INV_X2 \SB1_4_7/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[146] ), .ZN(
        \SB1_4_7/i1[9] ) );
  INV_X2 \SB1_2_0/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[188] ), .ZN(
        \SB1_2_0/i1[9] ) );
  INV_X2 \SB1_4_13/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[110] ), .ZN(
        \SB1_4_13/i1[9] ) );
  INV_X2 \SB1_3_12/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[116] ), .ZN(
        \SB1_3_12/i1[9] ) );
  INV_X2 \SB1_1_28/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[20] ), .ZN(
        \SB1_1_28/i1[9] ) );
  INV_X2 \SB1_1_6/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[155] ), .ZN(
        \SB1_1_6/i1_5 ) );
  INV_X2 \SB2_2_6/INV_3  ( .I(\SB1_2_8/buf_output[3] ), .ZN(\SB2_2_6/i0[8] )
         );
  BUF_X4 \SB2_2_31/BUF_1  ( .I(\SB1_2_3/buf_output[1] ), .Z(\SB2_2_31/i0[6] )
         );
  INV_X2 \SB1_3_20/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[68] ), .ZN(
        \SB1_3_20/i1[9] ) );
  INV_X2 \SB3_23/INV_5  ( .I(\RI1[5][53] ), .ZN(\SB3_23/i1_5 ) );
  BUF_X4 \SB1_1_23/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[51] ), .Z(
        \SB1_1_23/i0[10] ) );
  INV_X2 \SB2_2_24/INV_5  ( .I(\SB1_2_24/buf_output[5] ), .ZN(\SB2_2_24/i1_5 )
         );
  INV_X2 \SB1_4_31/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[2] ), .ZN(
        \SB1_4_31/i1[9] ) );
  INV_X2 \SB1_1_0/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[188] ), .ZN(
        \SB1_1_0/i1[9] ) );
  BUF_X4 \SB1_1_10/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[130] ), .Z(
        \SB1_1_10/i0_4 ) );
  INV_X2 \SB1_2_27/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[26] ), .ZN(
        \SB1_2_27/i1[9] ) );
  NAND3_X1 \SB3_8/Component_Function_0/N3  ( .A1(\SB3_8/i0[10] ), .A2(
        \SB3_8/i0_4 ), .A3(\SB3_8/i0_3 ), .ZN(
        \SB3_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_23/Component_Function_4/N4  ( .A1(\SB1_4_23/i1[9] ), .A2(
        \SB1_4_23/i1_5 ), .A3(\SB1_4_23/i0_4 ), .ZN(
        \SB1_4_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_2/N4  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0_0 ), .A3(n1105), .ZN(
        \SB1_0_31/Component_Function_2/NAND4_in[3] ) );
  INV_X2 \SB1_2_2/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[176] ), .ZN(
        \SB1_2_2/i1[9] ) );
  INV_X2 \SB2_4_19/INV_3  ( .I(\SB1_4_21/buf_output[3] ), .ZN(\SB2_4_19/i0[8] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_41  ( .I(\SB2_0_25/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[41] ) );
  INV_X2 \SB1_0_24/INV_2  ( .I(n268), .ZN(\SB1_0_24/i1[9] ) );
  INV_X2 \SB1_2_1/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[182] ), .ZN(
        \SB1_2_1/i1[9] ) );
  INV_X2 \SB1_3_19/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[74] ), .ZN(
        \SB1_3_19/i1[9] ) );
  BUF_X2 \SB1_0_27/BUF_2  ( .I(n262), .Z(\SB1_0_27/i0_0 ) );
  BUF_X4 \SB2_1_28/BUF_5  ( .I(\SB1_1_28/buf_output[5] ), .Z(\SB2_1_28/i0_3 )
         );
  BUF_X4 \SB1_4_0/BUF_2  ( .I(\MC_ARK_ARC_1_3/buf_output[188] ), .Z(
        \SB1_4_0/i0_0 ) );
  INV_X2 \SB1_3_11/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[122] ), .ZN(
        \SB1_3_11/i1[9] ) );
  INV_X2 \SB2_1_21/INV_3  ( .I(\SB1_1_23/buf_output[3] ), .ZN(\SB2_1_21/i0[8] ) );
  INV_X2 \SB1_1_7/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[146] ), .ZN(
        \SB1_1_7/i1[9] ) );
  BUF_X4 \SB2_3_17/BUF_4  ( .I(\SB1_3_18/buf_output[4] ), .Z(\SB2_3_17/i0_4 )
         );
  INV_X2 \SB3_1/INV_5  ( .I(\RI1[5][185] ), .ZN(\SB3_1/i1_5 ) );
  INV_X2 \SB2_1_24/INV_3  ( .I(\SB1_1_26/buf_output[3] ), .ZN(\SB2_1_24/i0[8] ) );
  INV_X2 \SB1_1_13/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[110] ), .ZN(
        \SB1_1_13/i1[9] ) );
  INV_X2 \SB2_2_9/INV_2  ( .I(\SB1_2_12/buf_output[2] ), .ZN(\SB2_2_9/i1[9] )
         );
  BUF_X4 \SB1_3_14/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[106] ), .Z(
        \SB1_3_14/i0_4 ) );
  INV_X2 \SB1_1_25/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[38] ), .ZN(
        \SB1_1_25/i1[9] ) );
  INV_X2 \SB3_31/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[2] ), .ZN(
        \SB3_31/i1[9] ) );
  INV_X2 \SB1_0_7/INV_2  ( .I(n302), .ZN(\SB1_0_7/i1[9] ) );
  INV_X2 \SB1_1_20/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[68] ), .ZN(
        \SB1_1_20/i1[9] ) );
  NAND3_X2 \SB1_2_10/Component_Function_5/N3  ( .A1(\SB1_2_10/i1[9] ), .A2(
        \SB1_2_10/i0_4 ), .A3(\SB1_2_10/i0_3 ), .ZN(
        \SB1_2_10/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 \SB1_1_9/Component_Function_1/N5  ( .A1(
        \SB1_1_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_9/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_9/buf_output[1] ) );
  NAND4_X1 \SB2_0_9/Component_Function_1/N5  ( .A1(
        \SB2_0_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_9/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_9/buf_output[1] ) );
  INV_X2 \SB1_1_14/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[104] ), .ZN(
        \SB1_1_14/i1[9] ) );
  INV_X2 \SB1_1_15/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[98] ), .ZN(
        \SB1_1_15/i1[9] ) );
  INV_X2 \SB2_3_17/INV_5  ( .I(\SB1_3_17/buf_output[5] ), .ZN(\SB2_3_17/i1_5 )
         );
  INV_X2 \SB1_4_26/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[32] ), .ZN(
        \SB1_4_26/i1[9] ) );
  INV_X2 \SB2_1_7/INV_3  ( .I(\SB1_1_9/buf_output[3] ), .ZN(\SB2_1_7/i0[8] )
         );
  INV_X2 \SB1_1_9/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[134] ), .ZN(
        \SB1_1_9/i1[9] ) );
  INV_X2 \SB1_0_23/INV_3  ( .I(n333), .ZN(\SB1_0_23/i0[8] ) );
  INV_X2 \SB2_0_20/INV_2  ( .I(\RI3[0][68] ), .ZN(\SB2_0_20/i1[9] ) );
  BUF_X4 \SB2_0_17/BUF_5  ( .I(\RI3[0][89] ), .Z(\SB2_0_17/i0_3 ) );
  INV_X2 \SB3_23/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[50] ), .ZN(
        \SB3_23/i1[9] ) );
  INV_X2 \SB1_0_9/INV_2  ( .I(n298), .ZN(\SB1_0_9/i1[9] ) );
  BUF_X2 \SB1_0_1/BUF_0  ( .I(n313), .Z(\SB1_0_1/i0[9] ) );
  INV_X2 \SB1_2_27/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[27] ), .ZN(
        \SB1_2_27/i0[8] ) );
  INV_X2 \SB1_2_25/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[41] ), .ZN(
        \SB1_2_25/i1_5 ) );
  INV_X2 \SB4_3/INV_2  ( .I(\SB3_6/buf_output[2] ), .ZN(\SB4_3/i1[9] ) );
  INV_X2 \SB2_0_13/INV_2  ( .I(\RI3[0][110] ), .ZN(\SB2_0_13/i1[9] ) );
  INV_X2 \SB1_2_6/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[152] ), .ZN(
        \SB1_2_6/i1[9] ) );
  INV_X2 \SB2_2_31/INV_2  ( .I(\SB1_2_2/buf_output[2] ), .ZN(\SB2_2_31/i1[9] )
         );
  INV_X2 \SB2_3_29/INV_2  ( .I(\SB1_3_0/buf_output[2] ), .ZN(\SB2_3_29/i1[9] )
         );
  INV_X2 \SB1_1_11/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[122] ), .ZN(
        \SB1_1_11/i1[9] ) );
  INV_X2 \SB1_2_13/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[111] ), .ZN(
        \SB1_2_13/i0[8] ) );
  BUF_X2 \SB1_0_4/BUF_1  ( .I(n248), .Z(\SB1_0_4/i0[6] ) );
  BUF_X2 \SB1_0_29/BUF_0  ( .I(n257), .Z(\SB1_0_29/i0[9] ) );
  BUF_X2 \SB1_0_12/BUF_0  ( .I(n291), .Z(\SB1_0_12/i0[9] ) );
  INV_X2 \SB1_2_23/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[50] ), .ZN(
        \SB1_2_23/i1[9] ) );
  INV_X2 \SB3_2/INV_5  ( .I(\RI1[5][179] ), .ZN(\SB3_2/i1_5 ) );
  INV_X2 \SB2_3_6/INV_2  ( .I(\SB1_3_9/buf_output[2] ), .ZN(\SB2_3_6/i1[9] )
         );
  NAND3_X2 \SB2_4_22/Component_Function_5/N4  ( .A1(\SB2_4_22/i0[9] ), .A2(
        \SB2_4_22/i0[6] ), .A3(\SB2_4_22/i0_4 ), .ZN(
        \SB2_4_22/Component_Function_5/NAND4_in[3] ) );
  INV_X2 \SB2_0_23/INV_5  ( .I(\RI3[0][53] ), .ZN(\SB2_0_23/i1_5 ) );
  INV_X2 \SB2_1_23/INV_5  ( .I(\SB1_1_23/buf_output[5] ), .ZN(\SB2_1_23/i1_5 )
         );
  INV_X2 \SB1_0_22/INV_2  ( .I(n272), .ZN(\SB1_0_22/i1[9] ) );
  INV_X2 \SB1_1_3/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[170] ), .ZN(
        \SB1_1_3/i1[9] ) );
  NAND3_X2 \SB2_0_19/Component_Function_5/N3  ( .A1(\SB2_0_19/i1[9] ), .A2(
        \RI3[0][76] ), .A3(\RI3[0][77] ), .ZN(
        \SB2_0_19/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB1_4_12/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[116] ), .ZN(
        \SB1_4_12/i1[9] ) );
  INV_X2 \SB2_0_13/INV_5  ( .I(\RI3[0][113] ), .ZN(\SB2_0_13/i1_5 ) );
  INV_X2 \SB1_1_17/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[86] ), .ZN(
        \SB1_1_17/i1[9] ) );
  INV_X2 \SB1_1_8/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[140] ), .ZN(
        \SB1_1_8/i1[9] ) );
  INV_X2 \SB1_0_4/INV_2  ( .I(n308), .ZN(\SB1_0_4/i1[9] ) );
  INV_X2 \SB3_12/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[116] ), .ZN(
        \SB3_12/i1[9] ) );
  INV_X2 \SB1_4_1/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[182] ), .ZN(
        \SB1_4_1/i1[9] ) );
  INV_X2 \SB1_1_21/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[62] ), .ZN(
        \SB1_1_21/i1[9] ) );
  INV_X2 \SB1_0_23/INV_2  ( .I(n270), .ZN(\SB1_0_23/i1[9] ) );
  INV_X2 \SB1_2_5/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[158] ), .ZN(
        \SB1_2_5/i1[9] ) );
  INV_X2 \SB1_4_29/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[14] ), .ZN(
        \SB1_4_29/i1[9] ) );
  INV_X2 \SB1_3_5/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[158] ), .ZN(
        \SB1_3_5/i1[9] ) );
  BUF_X2 \SB1_0_4/BUF_0  ( .I(n307), .Z(\SB1_0_4/i0[9] ) );
  INV_X2 \SB1_1_26/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[35] ), .ZN(
        \SB1_1_26/i1_5 ) );
  INV_X2 \SB2_0_9/INV_2  ( .I(\SB2_0_9/i0_0 ), .ZN(\SB2_0_9/i1[9] ) );
  INV_X2 \SB3_30/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[8] ), .ZN(
        \SB3_30/i1[9] ) );
  INV_X2 \SB2_0_21/INV_3  ( .I(\RI3[0][63] ), .ZN(\SB2_0_21/i0[8] ) );
  INV_X2 \SB3_27/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[26] ), .ZN(
        \SB3_27/i1[9] ) );
  INV_X2 \SB1_4_14/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[104] ), .ZN(
        \SB1_4_14/i1[9] ) );
  INV_X2 \SB1_3_13/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[110] ), .ZN(
        \SB1_3_13/i1[9] ) );
  INV_X2 \SB1_2_26/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[32] ), .ZN(
        \SB1_2_26/i1[9] ) );
  INV_X2 \SB1_4_19/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[74] ), .ZN(
        \SB1_4_19/i1[9] ) );
  BUF_X2 \SB1_0_10/BUF_1  ( .I(n242), .Z(\SB1_0_10/i0[6] ) );
  INV_X2 \SB1_1_27/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[26] ), .ZN(
        \SB1_1_27/i1[9] ) );
  BUF_X4 \SB2_0_12/BUF_0  ( .I(\RI3[0][114] ), .Z(\SB2_0_12/i0[9] ) );
  INV_X2 \SB1_2_25/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[38] ), .ZN(
        \SB1_2_25/i1[9] ) );
  INV_X2 \SB1_3_27/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[27] ), .ZN(
        \SB1_3_27/i0[8] ) );
  INV_X2 \SB2_0_0/INV_5  ( .I(\SB1_0_0/buf_output[5] ), .ZN(\SB2_0_0/i1_5 ) );
  INV_X2 \SB2_2_25/INV_2  ( .I(\SB1_2_28/buf_output[2] ), .ZN(\SB2_2_25/i1[9] ) );
  BUF_X2 \SB1_0_26/BUF_1  ( .I(n226), .Z(\SB1_0_26/i0[6] ) );
  INV_X2 \SB1_2_19/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[74] ), .ZN(
        \SB1_2_19/i1[9] ) );
  INV_X2 \SB1_0_16/INV_3  ( .I(n347), .ZN(\SB1_0_16/i0[8] ) );
  BUF_X4 \SB1_0_7/BUF_5  ( .I(n405), .Z(\SB1_0_7/i0_3 ) );
  INV_X2 \SB4_0/INV_5  ( .I(\SB3_0/buf_output[5] ), .ZN(\SB4_0/i1_5 ) );
  INV_X2 \SB1_3_25/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[38] ), .ZN(
        \SB1_3_25/i1[9] ) );
  INV_X2 \SB1_1_15/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[101] ), .ZN(
        \SB1_1_15/i1_5 ) );
  INV_X2 \SB3_7/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[146] ), .ZN(
        \SB3_7/i1[9] ) );
  INV_X2 \SB1_3_6/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[152] ), .ZN(
        \SB1_3_6/i1[9] ) );
  INV_X2 \SB2_3_18/INV_2  ( .I(\SB1_3_21/buf_output[2] ), .ZN(\SB2_3_18/i1[9] ) );
  INV_X2 \SB1_3_21/INV_5  ( .I(n3987), .ZN(\SB1_3_21/i1_5 ) );
  INV_X2 \SB1_3_7/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[147] ), .ZN(
        \SB1_3_7/i0[8] ) );
  INV_X2 \SB1_3_7/INV_2  ( .I(n1510), .ZN(\SB1_3_7/i1[9] ) );
  INV_X2 \SB1_2_4/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[164] ), .ZN(
        \SB1_2_4/i1[9] ) );
  INV_X2 \SB1_4_10/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[128] ), .ZN(
        \SB1_4_10/i1[9] ) );
  INV_X2 \SB1_4_20/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[71] ), .ZN(
        \SB1_4_20/i1_5 ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_97  ( .I(\SB2_4_19/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[97] ) );
  INV_X2 \SB1_0_19/INV_3  ( .I(n341), .ZN(\SB1_0_19/i0[8] ) );
  INV_X2 \SB2_3_31/INV_2  ( .I(\SB1_3_2/buf_output[2] ), .ZN(\SB2_3_31/i1[9] )
         );
  NAND4_X2 \SB1_2_2/Component_Function_2/N5  ( .A1(
        \SB1_2_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_2/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_2/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_2/buf_output[2] ) );
  NAND3_X2 \SB2_1_6/Component_Function_5/N4  ( .A1(\SB2_1_6/i0[9] ), .A2(
        \SB2_1_6/i0[6] ), .A3(\SB2_1_6/i0_4 ), .ZN(
        \SB2_1_6/Component_Function_5/NAND4_in[3] ) );
  INV_X2 \SB1_2_14/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[104] ), .ZN(
        \SB1_2_14/i1[9] ) );
  INV_X2 \SB2_0_18/INV_5  ( .I(\RI3[0][83] ), .ZN(\SB2_0_18/i1_5 ) );
  INV_X2 \SB2_4_19/INV_2  ( .I(\SB1_4_22/buf_output[2] ), .ZN(\SB2_4_19/i1[9] ) );
  BUF_X4 \SB2_3_3/BUF_4  ( .I(\SB1_3_4/buf_output[4] ), .Z(\SB2_3_3/i0_4 ) );
  INV_X2 \SB3_30/INV_5  ( .I(\RI1[5][11] ), .ZN(\SB3_30/i1_5 ) );
  INV_X2 \SB1_4_25/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[38] ), .ZN(
        \SB1_4_25/i1[9] ) );
  INV_X2 \SB2_1_20/INV_2  ( .I(\SB1_1_23/buf_output[2] ), .ZN(\SB2_1_20/i1[9] ) );
  INV_X2 \SB2_1_30/INV_5  ( .I(\SB1_1_30/buf_output[5] ), .ZN(\SB2_1_30/i1_5 )
         );
  INV_X2 \SB3_0/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[188] ), .ZN(
        \SB3_0/i1[9] ) );
  INV_X2 \SB2_2_16/INV_5  ( .I(\RI3[2][95] ), .ZN(\SB2_2_16/i1_5 ) );
  INV_X2 \SB1_3_8/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[140] ), .ZN(
        \SB1_3_8/i1[9] ) );
  INV_X2 \SB1_0_20/INV_2  ( .I(n276), .ZN(\SB1_0_20/i1[9] ) );
  INV_X2 \SB2_2_14/INV_5  ( .I(\SB1_2_14/buf_output[5] ), .ZN(\SB2_2_14/i1_5 )
         );
  INV_X2 \SB2_1_26/INV_2  ( .I(\SB1_1_29/buf_output[2] ), .ZN(\SB2_1_26/i1[9] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_64  ( .I(\SB2_0_22/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[64] ) );
  INV_X2 \SB1_2_9/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[134] ), .ZN(
        \SB1_2_9/i1[9] ) );
  INV_X2 \SB3_7/INV_5  ( .I(n6270), .ZN(\SB3_7/i1_5 ) );
  INV_X2 \SB1_4_0/INV_2  ( .I(n3977), .ZN(\SB1_4_0/i1[9] ) );
  INV_X2 \SB1_3_20/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[69] ), .ZN(
        \SB1_3_20/i0[8] ) );
  INV_X2 \SB1_3_31/INV_2  ( .I(n3982), .ZN(\SB1_3_31/i1[9] ) );
  INV_X2 \SB1_3_27/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[26] ), .ZN(
        \SB1_3_27/i1[9] ) );
  INV_X2 \SB1_4_25/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[39] ), .ZN(
        \SB1_4_25/i0[8] ) );
  INV_X2 \SB2_0_21/INV_5  ( .I(\RI3[0][65] ), .ZN(\SB2_0_21/i1_5 ) );
  INV_X2 \SB1_1_31/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[2] ), .ZN(
        \SB1_1_31/i1[9] ) );
  NAND4_X2 \SB2_4_23/Component_Function_2/N5  ( .A1(
        \SB2_4_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_23/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_4_23/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_4_23/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_4_23/buf_output[2] ) );
  NAND3_X1 \SB1_0_21/Component_Function_2/N3  ( .A1(\SB1_0_21/i0_3 ), .A2(
        \SB1_0_21/i0[8] ), .A3(\SB1_0_21/i0[9] ), .ZN(
        \SB1_0_21/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB1_0_8/INV_2  ( .I(n300), .ZN(\SB1_0_8/i1[9] ) );
  NAND4_X2 \SB1_3_5/Component_Function_2/N5  ( .A1(
        \SB1_3_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_5/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_3_5/buf_output[2] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_21  ( .I(\SB2_1_30/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[21] ) );
  INV_X2 \SB2_3_24/INV_5  ( .I(\SB1_3_24/buf_output[5] ), .ZN(\SB2_3_24/i1_5 )
         );
  NAND3_X1 \SB4_9/Component_Function_1/N4  ( .A1(\SB4_9/i1_7 ), .A2(n1499), 
        .A3(n6272), .ZN(\SB4_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_23/Component_Function_5/N3  ( .A1(\SB4_23/i1[9] ), .A2(
        \SB4_23/i0_4 ), .A3(\SB4_23/i0_3 ), .ZN(
        \SB4_23/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_22/Component_Function_1/N4  ( .A1(\SB2_4_22/i1_7 ), .A2(
        \SB2_4_22/i0[8] ), .A3(\SB2_4_22/i0_4 ), .ZN(
        \SB2_4_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_16/Component_Function_3/N4  ( .A1(\SB1_0_16/i1_5 ), .A2(
        \SB1_0_16/i0[8] ), .A3(\SB1_0_16/i3[0] ), .ZN(
        \SB1_0_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_2/N3  ( .A1(\SB1_0_7/i0_3 ), .A2(
        \SB1_0_7/i0[8] ), .A3(\SB1_0_7/i0[9] ), .ZN(
        \SB1_0_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_14/Component_Function_3/N3  ( .A1(\SB1_0_14/i1[9] ), .A2(
        \SB1_0_14/i1_7 ), .A3(\SB1_0_14/i0[10] ), .ZN(
        \SB1_0_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_23/Component_Function_3/N2  ( .A1(\SB1_0_23/i0_0 ), .A2(
        \SB1_0_23/i0_3 ), .A3(\SB1_0_23/i0_4 ), .ZN(
        \SB1_0_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_21/Component_Function_5/N4  ( .A1(\SB1_0_21/i0[9] ), .A2(
        \SB1_0_21/i0[6] ), .A3(\SB1_0_21/i0_4 ), .ZN(
        \SB1_0_21/Component_Function_5/NAND4_in[3] ) );
  BUF_X2 \SB1_0_18/BUF_0  ( .I(n279), .Z(\SB1_0_18/i0[9] ) );
  BUF_X2 \SB1_0_25/BUF_0  ( .I(n265), .Z(\SB1_0_25/i0[9] ) );
  BUF_X2 \SB1_0_23/BUF_0  ( .I(n269), .Z(\SB1_0_23/i0[9] ) );
  NAND3_X1 \SB4_21/Component_Function_1/N4  ( .A1(\SB4_21/i1_7 ), .A2(
        \SB4_21/i0[8] ), .A3(\SB4_21/i0_4 ), .ZN(
        \SB4_21/Component_Function_1/NAND4_in[3] ) );
  BUF_X2 \SB1_0_27/BUF_1  ( .I(n225), .Z(\SB1_0_27/i0[6] ) );
  INV_X2 \SB2_4_31/INV_2  ( .I(\SB1_4_2/buf_output[2] ), .ZN(\SB2_4_31/i1[9] )
         );
  INV_X2 \SB1_0_2/INV_2  ( .I(n312), .ZN(\SB1_0_2/i1[9] ) );
  NAND3_X2 \SB2_0_20/Component_Function_1/N4  ( .A1(\SB2_0_20/i1_7 ), .A2(
        \SB2_0_20/i0[8] ), .A3(\RI3[0][70] ), .ZN(
        \SB2_0_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 \SB1_1_2/Component_Function_5/N3  ( .A1(\SB1_1_2/i1[9] ), .A2(
        \SB1_1_2/i0_4 ), .A3(\SB1_1_2/i0_3 ), .ZN(
        \SB1_1_2/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB1_0_30/INV_2  ( .I(n256), .ZN(\SB1_0_30/i1[9] ) );
  BUF_X4 \SB2_1_18/BUF_4  ( .I(\SB1_1_19/buf_output[4] ), .Z(\SB2_1_18/i0_4 )
         );
  BUF_X4 \SB1_0_21/BUF_5  ( .I(n391), .Z(\SB1_0_21/i0_3 ) );
  NAND4_X2 \SB1_2_2/Component_Function_5/N5  ( .A1(
        \SB1_2_2/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_2_2/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_2/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_2_2/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_2_2/buf_output[5] ) );
  INV_X2 \SB1_0_13/INV_2  ( .I(n290), .ZN(\SB1_0_13/i1[9] ) );
  INV_X2 \SB2_3_31/INV_5  ( .I(\SB1_3_31/buf_output[5] ), .ZN(\SB2_3_31/i1_5 )
         );
  INV_X2 \SB1_0_30/INV_3  ( .I(n319), .ZN(\SB1_0_30/i0[8] ) );
  BUF_X4 \SB1_2_26/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[34] ), .Z(
        \SB1_2_26/i0_4 ) );
  BUF_X4 \SB1_2_24/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[45] ), .Z(
        \SB1_2_24/i0[10] ) );
  INV_X2 \SB2_1_4/INV_5  ( .I(\SB1_1_4/buf_output[5] ), .ZN(\SB2_1_4/i1_5 ) );
  NAND4_X2 \SB1_0_30/Component_Function_0/N5  ( .A1(
        \SB1_0_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_30/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_30/buf_output[0] ) );
  BUF_X4 \SB1_2_12/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[117] ), .Z(
        \SB1_2_12/i0[10] ) );
  NAND4_X2 \SB1_2_8/Component_Function_1/N5  ( .A1(
        \SB1_2_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_8/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_8/buf_output[1] ) );
  INV_X2 \SB2_2_5/INV_5  ( .I(\SB1_2_5/buf_output[5] ), .ZN(\SB2_2_5/i1_5 ) );
  INV_X2 \SB2_2_0/INV_2  ( .I(\SB1_2_3/buf_output[2] ), .ZN(\SB2_2_0/i1[9] )
         );
  INV_X2 \SB2_0_10/INV_3  ( .I(\RI3[0][129] ), .ZN(\SB2_0_10/i0[8] ) );
  NAND4_X1 \SB2_0_29/Component_Function_1/N5  ( .A1(
        \SB2_0_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_29/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_29/buf_output[1] ) );
  INV_X2 \SB1_0_5/INV_2  ( .I(n306), .ZN(\SB1_0_5/i1[9] ) );
  NAND4_X2 \SB2_2_5/Component_Function_0/N5  ( .A1(
        \SB2_2_5/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_5/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_5/buf_output[0] ) );
  BUF_X2 \SB1_0_28/BUF_1  ( .I(n224), .Z(\SB1_0_28/i0[6] ) );
  BUF_X4 \SB1_1_9/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[135] ), .Z(
        \SB1_1_9/i0[10] ) );
  INV_X2 \SB3_17/INV_5  ( .I(\RI1[5][89] ), .ZN(\SB3_17/i1_5 ) );
  INV_X2 \SB1_4_11/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[122] ), .ZN(
        \SB1_4_11/i1[9] ) );
  INV_X2 \SB3_13/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[110] ), .ZN(
        \SB3_13/i1[9] ) );
  NAND3_X2 \SB1_4_10/Component_Function_5/N3  ( .A1(\SB1_4_10/i1[9] ), .A2(
        \SB1_4_10/i0_4 ), .A3(\RI1[4][131] ), .ZN(
        \SB1_4_10/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB1_0_12/INV_2  ( .I(n292), .ZN(\SB1_0_12/i1[9] ) );
  BUF_X4 \SB1_1_23/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[52] ), .Z(
        \SB1_1_23/i0_4 ) );
  INV_X2 \SB1_4_16/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[92] ), .ZN(
        \SB1_4_16/i1[9] ) );
  NAND3_X2 \SB2_2_8/Component_Function_5/N3  ( .A1(\SB2_2_8/i1[9] ), .A2(
        \SB2_2_8/i0_4 ), .A3(\SB2_2_8/i0_3 ), .ZN(
        \SB2_2_8/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB1_0_24/INV_3  ( .I(n331), .ZN(\SB1_0_24/i0[8] ) );
  INV_X2 \SB1_2_9/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[137] ), .ZN(
        \SB1_2_9/i1_5 ) );
  NAND3_X2 \SB1_3_9/Component_Function_5/N3  ( .A1(\SB1_3_9/i1[9] ), .A2(
        \SB1_3_9/i0_4 ), .A3(\SB1_3_9/i0_3 ), .ZN(
        \SB1_3_9/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB2_0_29/INV_3  ( .I(\RI3[0][15] ), .ZN(\SB2_0_29/i0[8] ) );
  BUF_X2 \SB2_0_28/BUF_3_0  ( .I(\SB2_0_28/buf_output[3] ), .Z(\RI5[0][33] )
         );
  NAND4_X2 \SB2_0_6/Component_Function_3/N5  ( .A1(
        \SB2_0_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_6/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_6/buf_output[3] ) );
  NAND4_X2 \SB1_3_0/Component_Function_4/N5  ( .A1(
        \SB1_3_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_3_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_0/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_3_0/buf_output[4] ) );
  INV_X2 \SB3_31/INV_5  ( .I(n3981), .ZN(\SB3_31/i1_5 ) );
  NAND4_X2 \SB1_3_25/Component_Function_4/N5  ( .A1(
        \SB1_3_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_25/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_25/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_25/buf_output[4] ) );
  INV_X2 \SB2_2_28/INV_5  ( .I(\SB1_2_28/buf_output[5] ), .ZN(\SB2_2_28/i1_5 )
         );
  NAND4_X2 \SB1_4_4/Component_Function_4/N5  ( .A1(
        \SB1_4_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_4_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_4_4/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_4_4/buf_output[4] ) );
  INV_X2 \SB1_3_7/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[149] ), .ZN(
        \SB1_3_7/i1_5 ) );
  NAND4_X2 \SB1_1_12/Component_Function_0/N5  ( .A1(
        \SB1_1_12/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_12/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_12/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_12/buf_output[0] ) );
  NAND3_X2 \SB1_3_22/Component_Function_5/N4  ( .A1(\SB1_3_22/i0[9] ), .A2(
        \SB1_3_22/i0[6] ), .A3(\SB1_3_22/i0_4 ), .ZN(
        \SB1_3_22/Component_Function_5/NAND4_in[3] ) );
  INV_X2 \SB2_0_24/INV_2  ( .I(\RI3[0][44] ), .ZN(\SB2_0_24/i1[9] ) );
  BUF_X2 \SB1_0_27/BUF_0  ( .I(n261), .Z(\SB1_0_27/i0[9] ) );
  INV_X2 \SB2_1_11/INV_5  ( .I(\SB1_1_11/buf_output[5] ), .ZN(\SB2_1_11/i1_5 )
         );
  INV_X2 \SB2_0_17/INV_5  ( .I(\RI3[0][89] ), .ZN(\SB2_0_17/i1_5 ) );
  NAND4_X2 \SB2_1_18/Component_Function_4/N5  ( .A1(
        \SB2_1_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_18/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_18/buf_output[4] ) );
  INV_X2 \SB1_4_3/INV_5  ( .I(\RI1[4][173] ), .ZN(\SB1_4_3/i1_5 ) );
  BUF_X2 \SB1_0_24/BUF_3_0  ( .I(\SB1_0_24/buf_output[3] ), .Z(\RI3[0][57] )
         );
  INV_X2 \SB2_3_27/INV_5  ( .I(\SB1_3_27/buf_output[5] ), .ZN(\SB2_3_27/i1_5 )
         );
  INV_X2 \SB2_1_31/INV_2  ( .I(\SB1_1_2/buf_output[2] ), .ZN(\SB2_1_31/i1[9] )
         );
  NAND4_X2 \SB1_3_11/Component_Function_0/N5  ( .A1(
        \SB1_3_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_11/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_11/buf_output[0] ) );
  NAND3_X2 \SB2_2_5/Component_Function_5/N2  ( .A1(\SB2_2_5/i0_0 ), .A2(
        \SB2_2_5/i0[6] ), .A3(\SB2_2_5/i0[10] ), .ZN(
        \SB2_2_5/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB2_2_30/INV_5  ( .I(\SB1_2_30/buf_output[5] ), .ZN(\SB2_2_30/i1_5 )
         );
  INV_X2 \SB2_2_23/INV_5  ( .I(\SB1_2_23/buf_output[5] ), .ZN(\SB2_2_23/i1_5 )
         );
  NAND4_X2 \SB1_3_24/Component_Function_1/N5  ( .A1(
        \SB1_3_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_24/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_24/buf_output[1] ) );
  NAND4_X2 \SB1_0_27/Component_Function_0/N5  ( .A1(
        \SB1_0_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_27/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_27/buf_output[0] ) );
  NAND4_X2 \SB2_2_14/Component_Function_1/N5  ( .A1(
        \SB2_2_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_14/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_2_14/buf_output[1] ) );
  INV_X2 \SB2_3_30/INV_5  ( .I(\SB1_3_30/buf_output[5] ), .ZN(\SB2_3_30/i1_5 )
         );
  NAND4_X2 \SB1_4_5/Component_Function_0/N5  ( .A1(
        \SB1_4_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_4_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_5/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_4_5/buf_output[0] ) );
  NAND4_X2 \SB2_1_21/Component_Function_4/N5  ( .A1(
        \SB2_1_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_21/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_21/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_21/buf_output[4] ) );
  BUF_X2 \SB1_0_16/BUF_0  ( .I(n283), .Z(\SB1_0_16/i0[9] ) );
  BUF_X2 \SB1_0_3/BUF_1  ( .I(n249), .Z(\SB1_0_3/i0[6] ) );
  BUF_X2 \SB1_0_26/BUF_0  ( .I(n263), .Z(\SB1_0_26/i0[9] ) );
  CLKBUF_X4 \SB1_0_10/BUF_3  ( .I(n359), .Z(\SB1_0_10/i0[10] ) );
  CLKBUF_X4 \SB1_0_24/BUF_2  ( .I(n268), .Z(\SB1_0_24/i0_0 ) );
  CLKBUF_X4 \SB1_0_23/BUF_3  ( .I(n333), .Z(\SB1_0_23/i0[10] ) );
  BUF_X2 \SB1_0_17/BUF_0  ( .I(n281), .Z(\SB1_0_17/i0[9] ) );
  BUF_X2 \SB1_0_20/BUF_0  ( .I(n275), .Z(\SB1_0_20/i0[9] ) );
  BUF_X2 \SB1_0_22/BUF_0  ( .I(n271), .Z(\SB1_0_22/i0[9] ) );
  BUF_X2 \SB1_0_8/BUF_1  ( .I(n244), .Z(\SB1_0_8/i0[6] ) );
  BUF_X2 \SB1_0_8/BUF_0  ( .I(n299), .Z(\SB1_0_8/i0[9] ) );
  BUF_X2 \SB1_0_31/BUF_0  ( .I(n253), .Z(\SB1_0_31/i0[9] ) );
  CLKBUF_X4 \SB1_0_5/BUF_4  ( .I(n370), .Z(\SB1_0_5/i0_4 ) );
  CLKBUF_X4 \SB1_0_28/BUF_3  ( .I(n323), .Z(\SB1_0_28/i0[10] ) );
  BUF_X2 \SB1_0_6/BUF_0  ( .I(n303), .Z(\SB1_0_6/i0[9] ) );
  CLKBUF_X4 \SB1_0_7/BUF_2  ( .I(n302), .Z(\SB1_0_7/i0_0 ) );
  CLKBUF_X4 \SB1_0_1/BUF_3  ( .I(n377), .Z(\SB1_0_1/i0[10] ) );
  CLKBUF_X4 \SB1_0_1/BUF_4  ( .I(n378), .Z(\SB1_0_1/i0_4 ) );
  CLKBUF_X4 \SB1_0_30/BUF_3  ( .I(n319), .Z(\SB1_0_30/i0[10] ) );
  BUF_X2 \SB1_0_2/BUF_1  ( .I(n250), .Z(\SB1_0_2/i0[6] ) );
  BUF_X2 \SB1_0_2/BUF_0  ( .I(n311), .Z(\SB1_0_2/i0[9] ) );
  INV_X2 \SB2_0_23/INV_1  ( .I(\RI3[0][49] ), .ZN(\SB2_0_23/i1_7 ) );
  INV_X2 \SB2_0_9/INV_3  ( .I(\SB1_0_11/buf_output[3] ), .ZN(\SB2_0_9/i0[8] )
         );
  CLKBUF_X4 \SB2_0_22/BUF_0  ( .I(\SB1_0_27/buf_output[0] ), .Z(
        \SB2_0_22/i0[9] ) );
  CLKBUF_X4 \SB2_0_29/BUF_2  ( .I(\SB1_0_0/buf_output[2] ), .Z(\SB2_0_29/i0_0 ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_31  ( .I(\SB2_0_30/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[31] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_139  ( .I(\SB2_0_12/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[139] ) );
  CLKBUF_X4 \SB1_1_27/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[24] ), .Z(
        \SB1_1_27/i0[9] ) );
  CLKBUF_X4 \SB1_1_21/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[60] ), .Z(
        \SB1_1_21/i0[9] ) );
  CLKBUF_X4 \SB1_1_13/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[108] ), .Z(
        \SB1_1_13/i0[9] ) );
  CLKBUF_X4 \SB1_1_3/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[169] ), .Z(
        \SB1_1_3/i0[6] ) );
  BUF_X4 \SB1_1_11/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[125] ), .Z(
        \SB1_1_11/i0_3 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_168  ( .I(\SB2_1_8/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[168] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_103  ( .I(\SB2_1_18/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[103] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_187  ( .I(\SB2_1_4/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[187] ) );
  CLKBUF_X4 \SB1_2_27/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[25] ), .Z(
        \SB1_2_27/i0[6] ) );
  CLKBUF_X4 \SB1_2_9/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[133] ), .Z(
        \SB1_2_9/i0[6] ) );
  CLKBUF_X4 \SB2_2_30/BUF_1  ( .I(\SB1_2_2/buf_output[1] ), .Z(
        \SB2_2_30/i0[6] ) );
  CLKBUF_X4 \SB1_3_15/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[97] ), .Z(
        \SB1_3_15/i0[6] ) );
  BUF_X4 \SB1_3_6/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[153] ), .Z(
        \SB1_3_6/i0[10] ) );
  CLKBUF_X4 \SB2_3_7/BUF_1  ( .I(\SB1_3_11/buf_output[1] ), .Z(\SB2_3_7/i0[6] ) );
  CLKBUF_X4 \SB2_3_7/BUF_0  ( .I(\SB1_3_12/buf_output[0] ), .Z(\SB2_3_7/i0[9] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_1  ( .I(\SB2_3_3/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[1] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_115  ( .I(\SB2_3_16/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[115] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_133  ( .I(\SB2_3_13/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[133] ) );
  CLKBUF_X4 \SB1_4_13/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[108] ), .Z(
        \SB1_4_13/i0[9] ) );
  CLKBUF_X4 \SB1_4_18/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[78] ), .Z(
        \SB1_4_18/i0[9] ) );
  BUF_X4 \SB2_4_0/BUF_5  ( .I(\SB1_4_0/buf_output[5] ), .Z(\SB2_4_0/i0_3 ) );
  CLKBUF_X4 \SB4_18/BUF_0  ( .I(\SB3_23/buf_output[0] ), .Z(\SB4_18/i0[9] ) );
  NAND4_X2 \SB2_1_26/Component_Function_3/N5  ( .A1(
        \SB2_1_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_26/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_26/buf_output[3] ) );
  INV_X1 \SB1_0_30/INV_5  ( .I(n382), .ZN(\SB1_0_30/i1_5 ) );
  NAND4_X2 \SB1_0_9/Component_Function_5/N5  ( .A1(
        \SB1_0_9/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_0_9/buf_output[5] ) );
  NAND3_X2 \SB2_1_21/Component_Function_4/N4  ( .A1(\SB2_1_21/i1[9] ), .A2(
        \SB2_1_21/i1_5 ), .A3(\SB2_1_21/i0_4 ), .ZN(
        \SB2_1_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_17/Component_Function_2/N4  ( .A1(n3984), .A2(\SB4_17/i0_0 ), 
        .A3(\SB4_17/i0_4 ), .ZN(\SB4_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_24/Component_Function_4/N4  ( .A1(\SB3_24/i1[9] ), .A2(
        \SB3_24/i1_5 ), .A3(\SB3_24/i0_4 ), .ZN(
        \SB3_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N3  ( .A1(\SB3_26/i0[9] ), .A2(
        \SB3_26/i0[10] ), .A3(\SB3_26/i0_3 ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N3  ( .A1(\SB3_4/i0[9] ), .A2(
        \SB3_4/i0[10] ), .A3(\SB3_4/i0_3 ), .ZN(
        \SB3_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_29/Component_Function_1/N3  ( .A1(\SB1_4_29/i1_5 ), .A2(
        \SB1_4_29/i0[6] ), .A3(\SB1_4_29/i0[9] ), .ZN(
        \SB1_4_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_10/Component_Function_3/N2  ( .A1(\SB1_4_10/i0_0 ), .A2(
        \RI1[4][131] ), .A3(\SB1_4_10/i0_4 ), .ZN(
        \SB1_4_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_23/Component_Function_1/N4  ( .A1(\SB2_1_23/i1_7 ), .A2(
        \SB2_1_23/i0[8] ), .A3(\SB2_1_23/i0_4 ), .ZN(
        \SB2_1_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_30/Component_Function_4/N3  ( .A1(\SB2_1_30/i0[9] ), .A2(
        \SB2_1_30/i0[10] ), .A3(\SB2_1_30/i0_3 ), .ZN(
        \SB2_1_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_2/Component_Function_5/N4  ( .A1(\SB2_0_2/i0[9] ), .A2(
        \SB2_0_2/i0[6] ), .A3(\RI3[0][178] ), .ZN(
        \SB2_0_2/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_11/Component_Function_3/N2  ( .A1(\SB2_0_11/i0_0 ), .A2(
        \RI3[0][125] ), .A3(\SB2_0_11/i0_4 ), .ZN(
        \SB2_0_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_25/Component_Function_1/N3  ( .A1(\SB2_0_25/i1_5 ), .A2(
        \SB2_0_25/i0[6] ), .A3(\SB2_0_25/i0[9] ), .ZN(
        \SB2_0_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_9/Component_Function_2/N4  ( .A1(\SB2_0_9/i1_5 ), .A2(
        \SB2_0_9/i0_0 ), .A3(\SB2_0_9/i0_4 ), .ZN(
        \SB2_0_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_10/Component_Function_1/N4  ( .A1(\SB2_0_10/i1_7 ), .A2(
        \SB2_0_10/i0[8] ), .A3(\SB2_0_10/i0_4 ), .ZN(
        \SB2_0_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_11/Component_Function_0/N3  ( .A1(\SB2_0_11/i0[10] ), .A2(
        \SB2_0_11/i0_4 ), .A3(\SB2_0_11/i0_3 ), .ZN(
        \SB2_0_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_20/Component_Function_4/N4  ( .A1(\SB2_0_20/i1[9] ), .A2(
        \SB2_0_20/i1_5 ), .A3(\RI3[0][70] ), .ZN(
        \SB2_0_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_5/N4  ( .A1(\SB1_0_17/i0[9] ), .A2(
        n235), .A3(n346), .ZN(\SB1_0_17/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_3/N4  ( .A1(\SB1_0_7/i1_5 ), .A2(
        \SB1_0_7/i0[8] ), .A3(\SB1_0_7/i3[0] ), .ZN(
        \SB1_0_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N3  ( .A1(\SB1_0_27/i0[9] ), .A2(
        \SB1_0_27/i0[10] ), .A3(\SB1_0_27/i0_3 ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_30/Component_Function_4/N1  ( .A1(\SB1_0_30/i0[9] ), .A2(
        \SB1_0_30/i0_0 ), .A3(\SB1_0_30/i0[8] ), .ZN(
        \SB1_0_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_5/N4  ( .A1(\SB1_0_3/i0[9] ), .A2(n249), 
        .A3(n374), .ZN(\SB1_0_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_5/N4  ( .A1(n289), .A2(n239), .A3(n354), .ZN(\SB1_0_13/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_3/N3  ( .A1(\SB1_0_30/i1[9] ), .A2(
        \SB1_0_30/i1_7 ), .A3(\SB1_0_30/i0[10] ), .ZN(
        \SB1_0_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_2/Component_Function_5/N4  ( .A1(\SB1_0_2/i0[9] ), .A2(n250), 
        .A3(n376), .ZN(\SB1_0_2/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 \SB3_9/Component_Function_3/N5  ( .A1(
        \SB3_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_3/NAND4_in[3] ), .ZN(\SB3_9/buf_output[3] )
         );
  NAND3_X1 \SB2_2_8/Component_Function_4/N4  ( .A1(\SB2_2_8/i1[9] ), .A2(
        \SB2_2_8/i1_5 ), .A3(\SB2_2_8/i0_4 ), .ZN(
        \SB2_2_8/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 \SB1_3_14/Component_Function_0/N5  ( .A1(
        \SB1_3_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_14/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_14/buf_output[0] ) );
  NAND3_X2 \SB1_0_13/Component_Function_5/N3  ( .A1(\SB1_0_13/i1[9] ), .A2(
        \SB1_0_13/i0_4 ), .A3(\SB1_0_13/i0_3 ), .ZN(
        \SB1_0_13/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 \SB2_0_21/Component_Function_1/N5  ( .A1(
        \SB2_0_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_21/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_21/buf_output[1] ) );
  NAND4_X2 \SB2_4_10/Component_Function_4/N5  ( .A1(
        \SB2_4_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_4_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_4_10/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_4_10/buf_output[4] ) );
  BUF_X4 \SB1_0_19/BUF_4  ( .I(n342), .Z(\SB1_0_19/i0_4 ) );
  BUF_X4 \SB1_0_8/BUF_5  ( .I(n404), .Z(\SB1_0_8/i0_3 ) );
  INV_X2 \SB1_0_15/INV_2  ( .I(n286), .ZN(\SB1_0_15/i1[9] ) );
  NAND4_X2 \SB2_0_13/Component_Function_2/N5  ( .A1(
        \SB2_0_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_13/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_13/buf_output[2] ) );
  NAND4_X2 \SB1_1_11/Component_Function_4/N5  ( .A1(
        \SB1_1_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_11/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_11/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_11/buf_output[4] ) );
  INV_X2 \SB2_2_27/INV_5  ( .I(\SB1_2_27/buf_output[5] ), .ZN(\SB2_2_27/i1_5 )
         );
  NAND4_X2 \SB3_19/Component_Function_4/N5  ( .A1(
        \SB3_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_19/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_19/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_19/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_19/buf_output[4] ) );
  NAND4_X2 \SB2_1_11/Component_Function_4/N5  ( .A1(
        \SB2_1_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_11/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_11/buf_output[4] ) );
  NAND4_X2 \SB2_4_30/Component_Function_4/N5  ( .A1(
        \SB2_4_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_4_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_4_30/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_4_30/buf_output[4] ) );
  BUF_X4 \SB1_0_15/BUF_5  ( .I(n397), .Z(\SB1_0_15/i0_3 ) );
  NAND4_X2 \SB2_0_7/Component_Function_1/N5  ( .A1(
        \SB2_0_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_7/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_7/buf_output[1] ) );
  BUF_X4 \SB1_0_19/BUF_5  ( .I(n393), .Z(\SB1_0_19/i0_3 ) );
  BUF_X4 \SB2_4_3/BUF_4_0  ( .I(\SB2_4_3/buf_output[4] ), .Z(\RI5[4][178] ) );
  NAND4_X1 \SB2_0_31/Component_Function_2/N5  ( .A1(
        \SB2_0_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_31/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_31/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_31/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_31/buf_output[2] ) );
  NAND3_X2 \SB2_3_17/Component_Function_5/N2  ( .A1(\SB2_3_17/i0_0 ), .A2(
        \SB2_3_17/i0[6] ), .A3(\SB2_3_17/i0[10] ), .ZN(
        \SB2_3_17/Component_Function_5/NAND4_in[1] ) );
  INV_X1 \SB1_0_1/INV_5  ( .I(n411), .ZN(\SB1_0_1/i1_5 ) );
  INV_X1 \SB1_0_12/INV_5  ( .I(n400), .ZN(\SB1_0_12/i1_5 ) );
  NAND3_X1 \SB1_0_1/Component_Function_3/N3  ( .A1(\SB1_0_1/i1[9] ), .A2(
        \SB1_0_1/i1_7 ), .A3(\SB1_0_1/i0[10] ), .ZN(
        \SB1_0_1/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 \SB2_1_14/Component_Function_3/N5  ( .A1(
        \SB2_1_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_14/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_14/buf_output[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_4/N2  ( .A1(\SB1_0_17/i3[0] ), .A2(
        \SB1_0_17/i0_0 ), .A3(\SB1_0_17/i1_7 ), .ZN(
        \SB1_0_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_17/Component_Function_5/N2  ( .A1(\SB1_0_17/i0_0 ), .A2(
        \SB1_0_17/i0[6] ), .A3(\SB1_0_17/i0[10] ), .ZN(
        \SB1_0_17/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_1/Component_Function_2/N3  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i0[8] ), .A3(\SB1_0_1/i0[9] ), .ZN(
        \SB1_0_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_9/Component_Function_4/N3  ( .A1(\SB3_9/i0[9] ), .A2(
        \SB3_9/i0[10] ), .A3(\SB3_9/i0_3 ), .ZN(
        \SB3_9/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 \SB3_0/Component_Function_4/N5  ( .A1(
        \SB3_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_0/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_0/buf_output[4] )
         );
  NAND3_X1 \SB1_0_12/Component_Function_3/N2  ( .A1(\SB1_0_12/i0_0 ), .A2(
        \SB1_0_12/i0_3 ), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_12/Component_Function_4/N1  ( .A1(\SB1_0_12/i0[9] ), .A2(
        \SB1_0_12/i0_0 ), .A3(\SB1_0_12/i0[8] ), .ZN(
        \SB1_0_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_4/N2  ( .A1(\SB1_0_12/i3[0] ), .A2(
        \SB1_0_12/i0_0 ), .A3(\SB1_0_12/i1_7 ), .ZN(
        \SB1_0_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_19/Component_Function_1/N3  ( .A1(n6273), .A2(\SB4_19/i0[6] ), 
        .A3(\SB4_19/i0[9] ), .ZN(\SB4_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_11/Component_Function_4/N2  ( .A1(\SB2_3_11/i3[0] ), .A2(
        \SB2_3_11/i0_0 ), .A3(\SB2_3_11/i1_7 ), .ZN(
        \SB2_3_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_3/Component_Function_4/N3  ( .A1(\SB3_3/i0[9] ), .A2(
        \SB3_3/i0[10] ), .A3(\SB3_3/i0_3 ), .ZN(
        \SB3_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_6/Component_Function_0/N4  ( .A1(\SB4_6/i0[7] ), .A2(
        \SB4_6/i0_3 ), .A3(\SB4_6/i0_0 ), .ZN(
        \SB4_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_20/Component_Function_1/N3  ( .A1(\SB2_4_20/i1_5 ), .A2(
        \SB2_4_20/i0[6] ), .A3(\SB2_4_20/i0[9] ), .ZN(
        \SB2_4_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB1_4_31/Component_Function_5/N4  ( .A1(\SB1_4_31/i0[9] ), .A2(
        \SB1_4_31/i0[6] ), .A3(\SB1_4_31/i0_4 ), .ZN(
        \SB1_4_31/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 \SB2_1_11/Component_Function_3/N5  ( .A1(
        \SB2_1_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_11/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_11/buf_output[3] ) );
  NAND4_X2 \SB3_29/Component_Function_2/N5  ( .A1(
        \SB3_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_29/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_29/buf_output[2] ) );
  NAND4_X2 \SB2_0_17/Component_Function_4/N5  ( .A1(
        \SB2_0_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_17/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_17/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_17/buf_output[4] ) );
  NAND4_X2 \SB2_4_2/Component_Function_0/N5  ( .A1(
        \SB2_4_2/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_4_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_4_2/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_4_2/buf_output[0] ) );
  NAND3_X2 \SB2_0_17/Component_Function_4/N4  ( .A1(\SB2_0_17/i1[9] ), .A2(
        \SB2_0_17/i1_5 ), .A3(\RI3[0][88] ), .ZN(
        \SB2_0_17/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 \SB1_3_19/Component_Function_4/N5  ( .A1(
        \SB1_3_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_19/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_19/buf_output[4] ) );
  NAND4_X2 \SB1_2_16/Component_Function_2/N5  ( .A1(
        \SB1_2_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_16/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_16/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_16/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_16/buf_output[2] ) );
  NAND3_X2 \SB1_1_17/Component_Function_5/N4  ( .A1(\SB1_1_17/i0[9] ), .A2(
        \SB1_1_17/i0[6] ), .A3(\SB1_1_17/i0_4 ), .ZN(
        \SB1_1_17/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \SB2_3_8/BUF_4_0  ( .I(\SB2_3_8/buf_output[4] ), .Z(\RI5[3][148] ) );
  NAND4_X2 \SB1_3_28/Component_Function_4/N5  ( .A1(
        \SB1_3_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_28/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_28/buf_output[4] ) );
  NAND4_X2 \SB2_1_24/Component_Function_4/N5  ( .A1(
        \SB2_1_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_24/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_24/buf_output[4] ) );
  BUF_X4 \SB2_1_24/BUF_4_0  ( .I(\SB2_1_24/buf_output[4] ), .Z(\RI5[1][52] )
         );
  INV_X2 \SB1_2_28/INV_5  ( .I(n6291), .ZN(\SB1_2_28/i1_5 ) );
  NAND4_X2 \SB1_1_28/Component_Function_4/N5  ( .A1(
        \SB1_1_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_28/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_28/buf_output[4] ) );
  NAND4_X2 \SB2_2_19/Component_Function_4/N5  ( .A1(
        \SB2_2_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_19/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_19/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_2_19/buf_output[4] ) );
  NAND4_X2 \SB1_4_20/Component_Function_4/N5  ( .A1(
        \SB1_4_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_4_20/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_4_20/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_4_20/buf_output[4] ) );
  NAND4_X2 \SB2_4_11/Component_Function_4/N5  ( .A1(
        \SB2_4_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_4_11/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_4_11/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_4_11/buf_output[4] ) );
  NAND4_X2 \SB2_4_20/Component_Function_2/N5  ( .A1(
        \SB2_4_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_20/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_4_20/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_4_20/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_4_20/buf_output[2] ) );
  NAND4_X2 \SB2_2_25/Component_Function_4/N5  ( .A1(
        \SB2_2_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_25/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_25/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_2_25/buf_output[4] ) );
  NAND4_X2 \SB3_22/Component_Function_0/N5  ( .A1(
        \SB3_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_22/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_22/buf_output[0] ) );
  NAND4_X2 \SB1_2_24/Component_Function_1/N5  ( .A1(
        \SB1_2_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_24/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_24/buf_output[1] ) );
  NAND4_X2 \SB1_3_4/Component_Function_0/N5  ( .A1(
        \SB1_3_4/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_4/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_4/buf_output[0] ) );
  NAND4_X2 \SB1_1_22/Component_Function_1/N5  ( .A1(
        \SB1_1_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_22/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_22/buf_output[1] ) );
  NAND4_X2 \SB1_3_9/Component_Function_2/N5  ( .A1(
        \SB1_3_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_9/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_9/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_9/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_3_9/buf_output[2] ) );
  NAND4_X2 \SB1_2_20/Component_Function_2/N5  ( .A1(
        \SB1_2_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_20/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_20/buf_output[2] ) );
  INV_X1 \SB1_0_12/INV_1  ( .I(n240), .ZN(\SB1_0_12/i1_7 ) );
  BUF_X2 \SB1_0_11/BUF_0  ( .I(n293), .Z(\SB1_0_11/i0[9] ) );
  BUF_X2 \SB1_0_17/BUF_1  ( .I(n235), .Z(\SB1_0_17/i0[6] ) );
  INV_X1 \SB1_0_19/INV_5  ( .I(n393), .ZN(\SB1_0_19/i1_5 ) );
  NAND3_X1 \SB1_0_22/Component_Function_4/N4  ( .A1(\SB1_0_22/i1[9] ), .A2(
        \SB1_0_22/i1_5 ), .A3(\SB1_0_22/i0_4 ), .ZN(
        \SB1_0_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_4/N3  ( .A1(\SB1_0_24/i0[9] ), .A2(
        \SB1_0_24/i0[10] ), .A3(\SB1_0_24/i0_3 ), .ZN(
        \SB1_0_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_30/Component_Function_1/N2  ( .A1(\SB1_0_30/i0_3 ), .A2(
        \SB1_0_30/i1_7 ), .A3(\SB1_0_30/i0[8] ), .ZN(
        \SB1_0_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_11/Component_Function_0/N4  ( .A1(\SB1_0_11/i0[7] ), .A2(
        \SB1_0_11/i0_3 ), .A3(\SB1_0_11/i0_0 ), .ZN(
        \SB1_0_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_11/Component_Function_5/N4  ( .A1(\SB1_0_11/i0[9] ), .A2(
        \SB1_0_11/i0[6] ), .A3(\SB1_0_11/i0_4 ), .ZN(
        \SB1_0_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_22/Component_Function_5/N2  ( .A1(\SB1_0_22/i0_0 ), .A2(
        \SB1_0_22/i0[6] ), .A3(\SB1_0_22/i0[10] ), .ZN(
        \SB1_0_22/Component_Function_5/NAND4_in[1] ) );
  INV_X1 \SB2_0_7/INV_0  ( .I(\RI3[0][144] ), .ZN(\SB2_0_7/i3[0] ) );
  BUF_X2 \SB2_0_8/BUF_2  ( .I(\RI3[0][140] ), .Z(\SB2_0_8/i0_0 ) );
  INV_X1 \SB2_0_18/INV_0  ( .I(\RI3[0][78] ), .ZN(\SB2_0_18/i3[0] ) );
  INV_X1 \SB2_0_10/INV_0  ( .I(\RI3[0][126] ), .ZN(\SB2_0_10/i3[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_3/N2  ( .A1(\SB2_0_19/i0_0 ), .A2(
        \RI3[0][77] ), .A3(\RI3[0][76] ), .ZN(
        \SB2_0_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_26/Component_Function_1/N3  ( .A1(\SB2_0_26/i1_5 ), .A2(
        \SB2_0_26/i0[6] ), .A3(\SB2_0_26/i0[9] ), .ZN(
        \SB2_0_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_9/Component_Function_5/N3  ( .A1(\SB2_0_9/i1[9] ), .A2(
        \SB2_0_9/i0_4 ), .A3(\SB2_0_9/i0_3 ), .ZN(
        \SB2_0_9/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_28/Component_Function_5/N2  ( .A1(\SB2_0_28/i0_0 ), .A2(
        \SB2_0_28/i0[6] ), .A3(\SB2_0_28/i0[10] ), .ZN(
        \SB2_0_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_3/Component_Function_5/N4  ( .A1(\SB1_0_8/buf_output[0] ), 
        .A2(\SB2_0_3/i0[6] ), .A3(\RI3[0][172] ), .ZN(
        \SB2_0_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_31/Component_Function_4/N3  ( .A1(\SB2_0_31/i0[9] ), .A2(
        \SB2_0_31/i0[10] ), .A3(\SB2_0_31/i0_3 ), .ZN(
        \SB2_0_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_8/Component_Function_4/N3  ( .A1(\SB2_0_8/i0[9] ), .A2(
        \SB2_0_8/i0[10] ), .A3(\SB2_0_8/i0_3 ), .ZN(
        \SB2_0_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_17/Component_Function_5/N4  ( .A1(\SB2_0_17/i0[9] ), .A2(
        \SB2_0_17/i0[6] ), .A3(\RI3[0][88] ), .ZN(
        \SB2_0_17/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_11/Component_Function_1/N4  ( .A1(\SB2_0_11/i1_7 ), .A2(
        \SB2_0_11/i0[8] ), .A3(\SB2_0_11/i0_4 ), .ZN(
        \SB2_0_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_14/Component_Function_4/N4  ( .A1(\SB2_0_14/i1[9] ), .A2(
        \SB2_0_14/i1_5 ), .A3(\SB2_0_14/i0_4 ), .ZN(
        \SB2_0_14/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_75  ( .I(\SB2_0_21/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[75] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_137  ( .I(\SB2_0_9/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[137] ) );
  INV_X1 \SB1_1_16/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[91] ), .ZN(
        \SB1_1_16/i1_7 ) );
  BUF_X4 \SB1_1_15/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[101] ), .Z(
        \SB1_1_15/i0_3 ) );
  BUF_X4 \SB1_1_26/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[35] ), .Z(
        \SB1_1_26/i0_3 ) );
  BUF_X2 \SB1_1_0/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[186] ), .Z(
        \SB1_1_0/i0[9] ) );
  NAND3_X1 \SB1_1_17/Component_Function_2/N4  ( .A1(\SB1_1_17/i1_5 ), .A2(
        \SB1_1_17/i0_0 ), .A3(\MC_ARK_ARC_1_0/buf_output[88] ), .ZN(
        \SB1_1_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_10/Component_Function_0/N4  ( .A1(\SB1_1_10/i0[7] ), .A2(
        \SB1_1_10/i0_3 ), .A3(\SB1_1_10/i0_0 ), .ZN(
        \SB1_1_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_22/Component_Function_2/N4  ( .A1(\SB1_1_22/i1_5 ), .A2(
        \SB1_1_22/i0_0 ), .A3(\SB1_1_22/i0_4 ), .ZN(
        \SB1_1_22/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_28/Component_Function_1/N4  ( .A1(\SB1_1_28/i1_7 ), .A2(
        \SB1_1_28/i0[8] ), .A3(\SB1_1_28/i0_4 ), .ZN(
        \SB1_1_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_12/Component_Function_4/N4  ( .A1(\SB1_1_12/i1[9] ), .A2(
        \SB1_1_12/i1_5 ), .A3(\SB1_1_12/i0_4 ), .ZN(
        \SB1_1_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_6/Component_Function_5/N4  ( .A1(\SB1_1_6/i0[9] ), .A2(
        \SB1_1_6/i0[6] ), .A3(\SB1_1_6/i0_4 ), .ZN(
        \SB1_1_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_11/Component_Function_5/N2  ( .A1(\SB1_1_11/i0_0 ), .A2(
        \SB1_1_11/i0[6] ), .A3(\SB1_1_11/i0[10] ), .ZN(
        \SB1_1_11/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_4/Component_Function_2/N2  ( .A1(\SB1_1_4/i0_3 ), .A2(
        \SB1_1_4/i0[10] ), .A3(\SB1_1_4/i0[6] ), .ZN(
        \SB1_1_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_22/Component_Function_4/N4  ( .A1(\SB1_1_22/i1[9] ), .A2(
        \SB1_1_22/i1_5 ), .A3(\SB1_1_22/i0_4 ), .ZN(
        \SB1_1_22/Component_Function_4/NAND4_in[3] ) );
  BUF_X2 \SB2_1_2/BUF_0  ( .I(\SB1_1_7/buf_output[0] ), .Z(\SB2_1_2/i0[9] ) );
  INV_X1 \SB2_1_29/INV_0  ( .I(\SB1_1_2/buf_output[0] ), .ZN(\SB2_1_29/i3[0] )
         );
  INV_X1 \SB2_1_8/INV_1  ( .I(\SB1_1_12/buf_output[1] ), .ZN(\SB2_1_8/i1_7 )
         );
  NAND3_X1 \SB2_1_9/Component_Function_4/N4  ( .A1(\SB2_1_9/i1[9] ), .A2(
        \SB2_1_9/i1_5 ), .A3(\SB2_1_9/i0_4 ), .ZN(
        \SB2_1_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_15/Component_Function_5/N4  ( .A1(\SB2_1_15/i0[9] ), .A2(
        \SB2_1_15/i0[6] ), .A3(\SB2_1_15/i0_4 ), .ZN(
        \SB2_1_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_21/Component_Function_4/N1  ( .A1(\SB2_1_21/i0[9] ), .A2(
        \SB2_1_21/i0_0 ), .A3(\SB2_1_21/i0[8] ), .ZN(
        \SB2_1_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_5/N4  ( .A1(\SB1_1_27/buf_output[0] ), 
        .A2(\SB2_1_22/i0[6] ), .A3(\SB2_1_22/i0_4 ), .ZN(
        \SB2_1_22/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_22  ( .I(\SB2_1_29/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[22] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_45  ( .I(\SB2_1_26/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[45] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_189  ( .I(\SB2_1_2/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[189] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_110  ( .I(\SB2_1_16/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[110] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_32  ( .I(\SB2_1_29/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[32] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_150  ( .I(\SB2_1_11/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[150] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_72  ( .I(\SB2_1_24/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[72] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_36  ( .I(\SB2_1_30/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[36] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_163  ( .I(\SB2_1_8/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[163] ) );
  INV_X1 \SB1_2_7/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[145] ), .ZN(
        \SB1_2_7/i1_7 ) );
  NAND3_X1 \SB1_2_14/Component_Function_4/N3  ( .A1(\SB1_2_14/i0[9] ), .A2(
        \SB1_2_14/i0[10] ), .A3(\RI1[2][107] ), .ZN(
        \SB1_2_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_7/Component_Function_3/N1  ( .A1(\SB1_2_7/i1[9] ), .A2(
        \RI1[2][149] ), .A3(\SB1_2_7/i0[6] ), .ZN(
        \SB1_2_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_4/N3  ( .A1(\SB1_2_23/i0[9] ), .A2(
        \SB1_2_23/i0[10] ), .A3(\SB1_2_23/i0_3 ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[2] ) );
  INV_X1 \SB2_2_16/INV_1  ( .I(\SB1_2_20/buf_output[1] ), .ZN(\SB2_2_16/i1_7 )
         );
  NAND3_X1 \SB2_2_17/Component_Function_4/N4  ( .A1(\SB2_2_17/i1[9] ), .A2(
        \SB2_2_17/i1_5 ), .A3(\SB1_2_18/buf_output[4] ), .ZN(
        \SB2_2_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_9/Component_Function_4/N2  ( .A1(\SB2_2_9/i3[0] ), .A2(
        \SB2_2_9/i0_0 ), .A3(\SB2_2_9/i1_7 ), .ZN(
        \SB2_2_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_13/Component_Function_4/N4  ( .A1(\SB2_2_13/i1[9] ), .A2(
        \SB2_2_13/i1_5 ), .A3(\SB2_2_13/i0_4 ), .ZN(
        \SB2_2_13/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_99  ( .I(\SB2_2_17/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[99] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_68  ( .I(\SB2_2_23/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[68] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_92  ( .I(\SB2_2_19/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[92] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_120  ( .I(\SB2_2_16/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[120] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_89  ( .I(\SB2_2_17/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[89] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_151  ( .I(\SB2_2_10/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[151] ) );
  NAND3_X1 \SB1_3_14/Component_Function_1/N4  ( .A1(\SB1_3_14/i1_7 ), .A2(
        \SB1_3_14/i0[8] ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_8/Component_Function_1/N4  ( .A1(\SB1_3_8/i1_7 ), .A2(
        \SB1_3_8/i0[8] ), .A3(\SB1_3_8/i0_4 ), .ZN(
        \SB1_3_8/Component_Function_1/NAND4_in[3] ) );
  INV_X1 \SB2_3_11/INV_0  ( .I(\SB1_3_16/buf_output[0] ), .ZN(\SB2_3_11/i3[0] ) );
  INV_X1 \SB2_3_6/INV_0  ( .I(\SB1_3_11/buf_output[0] ), .ZN(\SB2_3_6/i3[0] )
         );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_129  ( .I(\SB2_3_12/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[129] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_69  ( .I(\SB2_3_22/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[69] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_128  ( .I(\SB2_3_13/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[128] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_20  ( .I(\SB2_3_31/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[20] ) );
  NAND3_X1 \SB1_4_24/Component_Function_4/N3  ( .A1(\SB1_4_24/i0[9] ), .A2(
        \SB1_4_24/i0[10] ), .A3(\SB1_4_24/i0_3 ), .ZN(
        \SB1_4_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_10/Component_Function_3/N3  ( .A1(\SB2_4_10/i1[9] ), .A2(
        \SB2_4_10/i1_7 ), .A3(\SB2_4_10/i0[10] ), .ZN(
        \SB2_4_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_9/Component_Function_1/N4  ( .A1(\SB2_4_9/i1_7 ), .A2(
        \SB2_4_9/i0[8] ), .A3(\SB2_4_9/i0_4 ), .ZN(
        \SB2_4_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_23/Component_Function_4/N4  ( .A1(\SB2_4_23/i1[9] ), .A2(
        \SB2_4_23/i1_5 ), .A3(\SB2_4_23/i0_4 ), .ZN(
        \SB2_4_23/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_171  ( .I(\SB2_4_5/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[171] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_188  ( .I(\SB2_4_3/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[188] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_168  ( .I(\SB2_4_8/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[168] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_53  ( .I(\SB2_4_23/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[53] ) );
  NAND3_X1 \SB3_19/Component_Function_4/N4  ( .A1(\SB3_19/i1[9] ), .A2(
        \SB3_19/i1_5 ), .A3(\SB3_19/i0_4 ), .ZN(
        \SB3_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_6/Component_Function_4/N3  ( .A1(\SB3_6/i0[9] ), .A2(
        \SB3_6/i0[10] ), .A3(\SB3_6/i0_3 ), .ZN(
        \SB3_6/Component_Function_4/NAND4_in[2] ) );
  INV_X1 \SB4_4/INV_5  ( .I(\SB3_4/buf_output[5] ), .ZN(\SB4_4/i1_5 ) );
  NAND3_X1 \SB4_26/Component_Function_1/N2  ( .A1(\SB4_26/i0_3 ), .A2(
        \SB4_26/i1_7 ), .A3(n3989), .ZN(
        \SB4_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_6/Component_Function_2/N3  ( .A1(\SB4_6/i0_3 ), .A2(
        \SB4_6/i0[8] ), .A3(\SB4_6/i0[9] ), .ZN(
        \SB4_6/Component_Function_2/NAND4_in[2] ) );
  INV_X1 U1 ( .I(n209), .ZN(n454) );
  INV_X1 U4 ( .I(n21), .ZN(n492) );
  INV_X1 U8 ( .I(n11), .ZN(n417) );
  INV_X1 U9 ( .I(n5), .ZN(n448) );
  INV_X1 U10 ( .I(n549), .ZN(n186) );
  CLKBUF_X2 U11 ( .I(Key[143]), .Z(n209) );
  BUF_X2 U12 ( .I(Key[47]), .Z(n185) );
  BUF_X2 U13 ( .I(Key[88]), .Z(n218) );
  BUF_X2 U14 ( .I(Key[183]), .Z(n208) );
  BUF_X2 U17 ( .I(Key[86]), .Z(n196) );
  CLKBUF_X2 U65 ( .I(Key[2]), .Z(n42) );
  CLKBUF_X2 U66 ( .I(Key[90]), .Z(n25) );
  CLKBUF_X2 U67 ( .I(Key[0]), .Z(n37) );
  CLKBUF_X2 U68 ( .I(Key[31]), .Z(n6) );
  CLKBUF_X2 U71 ( .I(Key[187]), .Z(n11) );
  CLKBUF_X2 U72 ( .I(Key[114]), .Z(n83) );
  CLKBUF_X2 U74 ( .I(Key[162]), .Z(n43) );
  CLKBUF_X2 U75 ( .I(Key[72]), .Z(n16) );
  CLKBUF_X2 U77 ( .I(Key[36]), .Z(n7) );
  CLKBUF_X2 U78 ( .I(Key[78]), .Z(n71) );
  CLKBUF_X2 U80 ( .I(Key[151]), .Z(n5) );
  CLKBUF_X2 U81 ( .I(Key[186]), .Z(n2) );
  BUF_X2 U83 ( .I(Key[19]), .Z(n215) );
  CLKBUF_X2 U84 ( .I(Key[84]), .Z(n74) );
  CLKBUF_X2 U86 ( .I(Key[174]), .Z(n39) );
  CLKBUF_X2 U87 ( .I(Key[48]), .Z(n67) );
  BUF_X2 U88 ( .I(Key[185]), .Z(n187) );
  BUF_X2 U90 ( .I(Key[7]), .Z(n193) );
  INV_X1 U91 ( .I(n452), .ZN(n1) );
  BUF_X2 U93 ( .I(Key[65]), .Z(n194) );
  BUF_X2 U96 ( .I(Key[158]), .Z(n3) );
  BUF_X2 U97 ( .I(Key[98]), .Z(n4) );
  CLKBUF_X2 U98 ( .I(Key[42]), .Z(n10) );
  BUF_X2 U99 ( .I(Key[124]), .Z(n12) );
  BUF_X2 U100 ( .I(Key[153]), .Z(n14) );
  BUF_X2 U101 ( .I(Key[117]), .Z(n15) );
  BUF_X2 U102 ( .I(Key[99]), .Z(n17) );
  BUF_X2 U103 ( .I(Key[127]), .Z(n18) );
  BUF_X2 U104 ( .I(Key[176]), .Z(n19) );
  BUF_X2 U105 ( .I(Key[94]), .Z(n21) );
  BUF_X2 U106 ( .I(Key[92]), .Z(n22) );
  BUF_X2 U107 ( .I(Key[160]), .Z(n23) );
  BUF_X2 U108 ( .I(Key[13]), .Z(n24) );
  BUF_X2 U109 ( .I(Key[53]), .Z(n26) );
  BUF_X2 U110 ( .I(Key[121]), .Z(n27) );
  BUF_X2 U112 ( .I(Key[14]), .Z(n31) );
  BUF_X2 U113 ( .I(Key[133]), .Z(n32) );
  BUF_X2 U114 ( .I(Key[166]), .Z(n34) );
  BUF_X2 U115 ( .I(Key[155]), .Z(n35) );
  BUF_X2 U116 ( .I(Key[50]), .Z(n36) );
  BUF_X2 U117 ( .I(Key[64]), .Z(n40) );
  BUF_X2 U118 ( .I(Key[5]), .Z(n41) );
  BUF_X2 U119 ( .I(Key[189]), .Z(n47) );
  BUF_X2 U121 ( .I(Key[157]), .Z(n49) );
  BUF_X2 U122 ( .I(Key[108]), .Z(n52) );
  BUF_X2 U123 ( .I(Key[144]), .Z(n53) );
  BUF_X2 U125 ( .I(Key[132]), .Z(n55) );
  BUF_X2 U126 ( .I(Key[175]), .Z(n57) );
  BUF_X2 U127 ( .I(Key[171]), .Z(n58) );
  BUF_X2 U128 ( .I(Key[182]), .Z(n59) );
  BUF_X2 U129 ( .I(Key[109]), .Z(n60) );
  BUF_X2 U130 ( .I(Key[136]), .Z(n61) );
  BUF_X2 U131 ( .I(Key[128]), .Z(n62) );
  BUF_X2 U132 ( .I(Key[129]), .Z(n63) );
  BUF_X2 U133 ( .I(Key[107]), .Z(n65) );
  BUF_X2 U134 ( .I(Key[27]), .Z(n66) );
  XOR2_X1 U135 ( .A1(Plaintext[144]), .A2(Key[144]), .Z(n301) );
  BUF_X2 U136 ( .I(Key[73]), .Z(n68) );
  BUF_X2 U137 ( .I(Key[112]), .Z(n69) );
  BUF_X2 U138 ( .I(Key[131]), .Z(n70) );
  BUF_X2 U139 ( .I(Key[57]), .Z(n72) );
  BUF_X2 U140 ( .I(Key[93]), .Z(n73) );
  BUF_X2 U141 ( .I(Key[87]), .Z(n75) );
  BUF_X2 U142 ( .I(Key[149]), .Z(n76) );
  BUF_X2 U143 ( .I(Key[41]), .Z(n77) );
  BUF_X2 U144 ( .I(Key[60]), .Z(n79) );
  BUF_X2 U145 ( .I(Key[77]), .Z(n80) );
  BUF_X2 U146 ( .I(Key[115]), .Z(n81) );
  BUF_X2 U147 ( .I(Key[156]), .Z(n82) );
  BUF_X2 U148 ( .I(Key[81]), .Z(n85) );
  BUF_X2 U150 ( .I(Key[150]), .Z(n88) );
  BUF_X2 U151 ( .I(Key[23]), .Z(n91) );
  BUF_X2 U152 ( .I(Key[17]), .Z(n92) );
  BUF_X2 U154 ( .I(Key[163]), .Z(n96) );
  BUF_X2 U155 ( .I(Key[161]), .Z(n97) );
  BUF_X2 U159 ( .I(Key[10]), .Z(n103) );
  BUF_X2 U160 ( .I(Key[21]), .Z(n104) );
  BUF_X2 U161 ( .I(Key[49]), .Z(n105) );
  BUF_X2 U164 ( .I(Key[37]), .Z(n107) );
  BUF_X2 U165 ( .I(Key[29]), .Z(n108) );
  BUF_X2 U167 ( .I(Key[63]), .Z(n110) );
  BUF_X2 U168 ( .I(Key[180]), .Z(n111) );
  BUF_X2 U171 ( .I(Key[134]), .Z(n112) );
  BUF_X2 U174 ( .I(Key[51]), .Z(n117) );
  BUF_X2 U176 ( .I(Key[168]), .Z(n119) );
  BUF_X2 U177 ( .I(Key[105]), .Z(n120) );
  XOR2_X1 U178 ( .A1(Plaintext[10]), .A2(Key[10]), .Z(n320) );
  BUF_X2 U179 ( .I(Key[66]), .Z(n121) );
  BUF_X2 U180 ( .I(Key[190]), .Z(n122) );
  BUF_X2 U182 ( .I(Key[178]), .Z(n124) );
  BUF_X2 U183 ( .I(Key[167]), .Z(n125) );
  BUF_X2 U184 ( .I(Key[16]), .Z(n126) );
  BUF_X2 U185 ( .I(Key[118]), .Z(n128) );
  BUF_X2 U186 ( .I(Key[135]), .Z(n129) );
  BUF_X2 U187 ( .I(Key[32]), .Z(n130) );
  BUF_X2 U189 ( .I(Key[82]), .Z(n132) );
  BUF_X2 U193 ( .I(Key[170]), .Z(n136) );
  BUF_X2 U202 ( .I(Key[25]), .Z(n146) );
  BUF_X2 U203 ( .I(Key[122]), .Z(n147) );
  BUF_X2 U206 ( .I(Key[69]), .Z(n151) );
  BUF_X2 U209 ( .I(Key[26]), .Z(n155) );
  BUF_X2 U211 ( .I(Key[8]), .Z(n157) );
  BUF_X2 U213 ( .I(Key[95]), .Z(n160) );
  BUF_X2 U215 ( .I(Key[20]), .Z(n162) );
  BUF_X2 U218 ( .I(Key[188]), .Z(n166) );
  BUF_X2 U220 ( .I(Key[3]), .Z(n169) );
  BUF_X2 U223 ( .I(Key[4]), .Z(n173) );
  BUF_X2 U224 ( .I(Key[191]), .Z(n174) );
  BUF_X2 U229 ( .I(Key[111]), .Z(n179) );
  BUF_X2 U230 ( .I(Key[177]), .Z(n180) );
  XOR2_X1 U231 ( .A1(Plaintext[97]), .A2(Key[97]), .Z(n237) );
  XOR2_X1 U232 ( .A1(Plaintext[3]), .A2(Key[3]), .Z(n317) );
  XOR2_X1 U233 ( .A1(Plaintext[96]), .A2(Key[96]), .Z(n285) );
  XOR2_X1 U237 ( .A1(Plaintext[126]), .A2(Key[126]), .Z(n295) );
  XOR2_X1 U238 ( .A1(Plaintext[7]), .A2(Key[7]), .Z(n222) );
  XOR2_X1 U242 ( .A1(Plaintext[52]), .A2(Key[52]), .Z(n334) );
  XOR2_X1 U246 ( .A1(Key[76]), .A2(Plaintext[76]), .Z(n342) );
  INV_X1 U249 ( .I(Key[28]), .ZN(n158) );
  INV_X1 U251 ( .I(n195), .ZN(n8) );
  INV_X1 U252 ( .I(n203), .ZN(n51) );
  INV_X1 U253 ( .I(n130), .ZN(n542) );
  INV_X1 U254 ( .I(n210), .ZN(n148) );
  INV_X1 U255 ( .I(n208), .ZN(n9) );
  INV_X1 U256 ( .I(n149), .ZN(n482) );
  INV_X1 U257 ( .I(n157), .ZN(n562) );
  INV_X1 U258 ( .I(n110), .ZN(n518) );
  INV_X1 U260 ( .I(n212), .ZN(n89) );
  INV_X1 U262 ( .I(n219), .ZN(n44) );
  INV_X1 U263 ( .I(n166), .ZN(n416) );
  INV_X1 U264 ( .I(n129), .ZN(n459) );
  INV_X1 U265 ( .I(n133), .ZN(n561) );
  INV_X1 U266 ( .I(n159), .ZN(n473) );
  INV_X1 U267 ( .I(n111), .ZN(n422) );
  INV_X1 U268 ( .I(n135), .ZN(n514) );
  INV_X1 U269 ( .I(n215), .ZN(n167) );
  INV_X1 U271 ( .I(n214), .ZN(n145) );
  INV_X1 U272 ( .I(n189), .ZN(n541) );
  INV_X1 U273 ( .I(n200), .ZN(n113) );
  INV_X1 U274 ( .I(n82), .ZN(n443) );
  INV_X1 U275 ( .I(\MC_ARK_ARC_1_1/buf_keyinput[111] ), .ZN(n87) );
  INV_X1 U276 ( .I(n184), .ZN(n20) );
  INV_X1 U277 ( .I(n211), .ZN(n445) );
  INV_X1 U278 ( .I(n173), .ZN(n565) );
  INV_X1 U279 ( .I(n141), .ZN(n507) );
  INV_X1 U280 ( .I(n139), .ZN(n64) );
  INV_X1 U281 ( .I(n88), .ZN(n449) );
  INV_X1 U282 ( .I(n78), .ZN(n568) );
  INV_X1 U283 ( .I(n180), .ZN(n424) );
  INV_X1 U284 ( .I(n109), .ZN(n435) );
  INV_X1 U285 ( .I(n85), .ZN(n503) );
  INV_X1 U286 ( .I(n91), .ZN(n550) );
  INV_X1 U287 ( .I(n72), .ZN(n522) );
  INV_X1 U288 ( .I(n75), .ZN(n497) );
  INV_X1 U290 ( .I(n146), .ZN(n548) );
  INV_X1 U292 ( .I(n37), .ZN(n569) );
  INV_X1 U294 ( .I(n144), .ZN(n521) );
  INV_X1 U295 ( .I(n71), .ZN(n505) );
  INV_X1 U296 ( .I(n152), .ZN(n538) );
  INV_X1 U297 ( .I(n112), .ZN(n460) );
  INV_X1 U298 ( .I(n174), .ZN(n413) );
  INV_X1 U299 ( .I(n202), .ZN(n115) );
  INV_X1 U300 ( .I(n114), .ZN(n447) );
  INV_X1 U301 ( .I(n155), .ZN(n547) );
  INV_X1 U302 ( .I(n108), .ZN(n545) );
  INV_X1 U303 ( .I(n213), .ZN(n90) );
  INV_X1 U305 ( .I(n217), .ZN(n50) );
  INV_X1 U306 ( .I(n216), .ZN(n13) );
  INV_X1 U307 ( .I(n181), .ZN(n533) );
  INV_X1 U308 ( .I(n69), .ZN(n480) );
  INV_X1 U309 ( .I(n154), .ZN(n523) );
  INV_X1 U310 ( .I(n160), .ZN(n491) );
  INV_X1 U311 ( .I(n103), .ZN(n560) );
  INV_X1 U312 ( .I(n190), .ZN(n504) );
  INV_X1 U315 ( .I(n106), .ZN(n511) );
  INV_X1 U316 ( .I(n24), .ZN(n557) );
  INV_X1 U317 ( .I(n128), .ZN(n474) );
  INV_X1 U318 ( .I(n196), .ZN(n498) );
  INV_X1 U319 ( .I(n205), .ZN(n476) );
  INV_X1 U320 ( .I(n137), .ZN(n451) );
  INV_X1 U321 ( .I(n68), .ZN(n508) );
  INV_X1 U323 ( .I(n163), .ZN(n559) );
  INV_X1 U324 ( .I(n206), .ZN(n45) );
  INV_X1 U325 ( .I(n187), .ZN(n419) );
  INV_X1 U327 ( .I(n119), .ZN(n432) );
  INV_X1 U328 ( .I(n100), .ZN(n456) );
  INV_X1 U329 ( .I(n118), .ZN(n421) );
  INV_X1 U330 ( .I(n77), .ZN(n537) );
  INV_X1 U331 ( .I(n107), .ZN(n539) );
  INV_X1 U332 ( .I(n138), .ZN(n513) );
  INV_X1 U334 ( .I(n162), .ZN(n552) );
  INV_X1 U335 ( .I(n175), .ZN(n487) );
  INV_X1 U336 ( .I(n39), .ZN(n427) );
  INV_X1 U338 ( .I(n43), .ZN(n438) );
  INV_X1 U339 ( .I(n197), .ZN(n524) );
  INV_X1 U340 ( .I(n169), .ZN(n566) );
  INV_X1 U341 ( .I(n172), .ZN(n33) );
  INV_X1 U342 ( .I(n49), .ZN(n442) );
  INV_X1 U343 ( .I(n63), .ZN(n464) );
  INV_X1 U344 ( .I(n53), .ZN(n453) );
  INV_X1 U345 ( .I(n96), .ZN(n437) );
  INV_X1 U346 ( .I(n204), .ZN(n171) );
  INV_X1 U347 ( .I(n58), .ZN(n429) );
  INV_X1 U348 ( .I(n95), .ZN(n558) );
  INV_X1 U349 ( .I(n47), .ZN(n415) );
  INV_X1 U350 ( .I(n151), .ZN(n512) );
  INV_X1 U352 ( .I(n25), .ZN(n495) );
  INV_X1 U353 ( .I(n201), .ZN(n153) );
  INV_X1 U354 ( .I(n156), .ZN(n94) );
  INV_X1 U355 ( .I(n179), .ZN(n481) );
  INV_X1 U356 ( .I(Key[24]), .ZN(n549) );
  INV_X1 U357 ( .I(n74), .ZN(n500) );
  INV_X1 U358 ( .I(n185), .ZN(n532) );
  INV_X1 U359 ( .I(n83), .ZN(n478) );
  INV_X1 U360 ( .I(n165), .ZN(n428) );
  INV_X1 U362 ( .I(n56), .ZN(n553) );
  INV_X1 U363 ( .I(n92), .ZN(n554) );
  INV_X1 U364 ( .I(n10), .ZN(n536) );
  INV_X1 U365 ( .I(n150), .ZN(n510) );
  INV_X1 U366 ( .I(n79), .ZN(n520) );
  INV_X1 U368 ( .I(n38), .ZN(n525) );
  INV_X1 U369 ( .I(n140), .ZN(n455) );
  INV_X1 U370 ( .I(n105), .ZN(n530) );
  INV_X1 U371 ( .I(n136), .ZN(n430) );
  INV_X1 U372 ( .I(n120), .ZN(n486) );
  INV_X1 U373 ( .I(n182), .ZN(n127) );
  INV_X1 U374 ( .I(n116), .ZN(n499) );
  INV_X1 U375 ( .I(n104), .ZN(n551) );
  INV_X1 U377 ( .I(n177), .ZN(n535) );
  INV_X1 U378 ( .I(n126), .ZN(n555) );
  INV_X1 U379 ( .I(n198), .ZN(n534) );
  INV_X1 U380 ( .I(n183), .ZN(n436) );
  INV_X1 U381 ( .I(Key[22]), .ZN(n164) );
  INV_X1 U382 ( .I(n218), .ZN(n102) );
  INV_X1 U383 ( .I(n191), .ZN(n84) );
  INV_X1 U384 ( .I(n142), .ZN(n527) );
  INV_X1 U386 ( .I(n124), .ZN(n423) );
  INV_X1 U387 ( .I(n48), .ZN(n519) );
  XOR2_X1 U388 ( .A1(Key[0]), .A2(Plaintext[0]), .Z(n253) );
  XOR2_X1 U389 ( .A1(Key[1]), .A2(Plaintext[1]), .Z(n221) );
  XOR2_X1 U390 ( .A1(Key[2]), .A2(Plaintext[2]), .Z(n254) );
  XOR2_X1 U391 ( .A1(Key[4]), .A2(Plaintext[4]), .Z(n318) );
  XOR2_X1 U392 ( .A1(Key[5]), .A2(Plaintext[5]), .Z(n381) );
  XOR2_X1 U393 ( .A1(Key[6]), .A2(Plaintext[6]), .Z(n255) );
  XOR2_X1 U394 ( .A1(Key[8]), .A2(Plaintext[8]), .Z(n256) );
  XOR2_X1 U395 ( .A1(Key[9]), .A2(Plaintext[9]), .Z(n319) );
  XOR2_X1 U396 ( .A1(Key[11]), .A2(Plaintext[11]), .Z(n382) );
  XOR2_X1 U397 ( .A1(Key[12]), .A2(Plaintext[12]), .Z(n257) );
  XOR2_X1 U398 ( .A1(Key[13]), .A2(Plaintext[13]), .Z(n223) );
  XOR2_X1 U399 ( .A1(Key[14]), .A2(Plaintext[14]), .Z(n258) );
  XOR2_X1 U400 ( .A1(Key[15]), .A2(Plaintext[15]), .Z(n321) );
  XOR2_X1 U401 ( .A1(Key[16]), .A2(Plaintext[16]), .Z(n322) );
  XOR2_X1 U402 ( .A1(Key[17]), .A2(Plaintext[17]), .Z(n383) );
  XOR2_X1 U403 ( .A1(Key[18]), .A2(Plaintext[18]), .Z(n259) );
  XOR2_X1 U404 ( .A1(Key[19]), .A2(Plaintext[19]), .Z(n224) );
  XOR2_X1 U405 ( .A1(Key[20]), .A2(Plaintext[20]), .Z(n260) );
  XOR2_X1 U406 ( .A1(Key[21]), .A2(Plaintext[21]), .Z(n323) );
  XOR2_X1 U407 ( .A1(Key[22]), .A2(Plaintext[22]), .Z(n324) );
  XOR2_X1 U408 ( .A1(Key[23]), .A2(Plaintext[23]), .Z(n384) );
  XOR2_X1 U409 ( .A1(Key[24]), .A2(Plaintext[24]), .Z(n261) );
  XOR2_X1 U410 ( .A1(Key[25]), .A2(Plaintext[25]), .Z(n225) );
  XOR2_X1 U411 ( .A1(Key[26]), .A2(Plaintext[26]), .Z(n262) );
  XOR2_X1 U412 ( .A1(Key[27]), .A2(Plaintext[27]), .Z(n325) );
  XOR2_X1 U413 ( .A1(Key[28]), .A2(Plaintext[28]), .Z(n326) );
  XOR2_X1 U414 ( .A1(Key[29]), .A2(Plaintext[29]), .Z(n385) );
  XOR2_X1 U415 ( .A1(Key[30]), .A2(Plaintext[30]), .Z(n263) );
  XOR2_X1 U416 ( .A1(Key[31]), .A2(Plaintext[31]), .Z(n226) );
  XOR2_X1 U417 ( .A1(Key[32]), .A2(Plaintext[32]), .Z(n264) );
  XOR2_X1 U418 ( .A1(Key[33]), .A2(Plaintext[33]), .Z(n327) );
  XOR2_X1 U419 ( .A1(Key[34]), .A2(Plaintext[34]), .Z(n328) );
  XOR2_X1 U420 ( .A1(Key[35]), .A2(Plaintext[35]), .Z(n386) );
  XOR2_X1 U421 ( .A1(Key[36]), .A2(Plaintext[36]), .Z(n265) );
  XOR2_X1 U422 ( .A1(Key[37]), .A2(Plaintext[37]), .Z(n227) );
  XOR2_X1 U423 ( .A1(Key[38]), .A2(Plaintext[38]), .Z(n266) );
  XOR2_X1 U424 ( .A1(Key[39]), .A2(Plaintext[39]), .Z(n329) );
  XOR2_X1 U425 ( .A1(Key[40]), .A2(Plaintext[40]), .Z(n330) );
  XOR2_X1 U426 ( .A1(Key[41]), .A2(Plaintext[41]), .Z(n387) );
  XOR2_X1 U427 ( .A1(Key[42]), .A2(Plaintext[42]), .Z(n267) );
  XOR2_X1 U428 ( .A1(Key[43]), .A2(Plaintext[43]), .Z(n228) );
  XOR2_X1 U429 ( .A1(Key[44]), .A2(Plaintext[44]), .Z(n268) );
  XOR2_X1 U430 ( .A1(Key[45]), .A2(Plaintext[45]), .Z(n331) );
  XOR2_X1 U431 ( .A1(Key[46]), .A2(Plaintext[46]), .Z(n332) );
  XOR2_X1 U432 ( .A1(Key[47]), .A2(Plaintext[47]), .Z(n388) );
  XOR2_X1 U433 ( .A1(Key[48]), .A2(Plaintext[48]), .Z(n269) );
  XOR2_X1 U434 ( .A1(Key[49]), .A2(Plaintext[49]), .Z(n229) );
  XOR2_X1 U435 ( .A1(Key[50]), .A2(Plaintext[50]), .Z(n270) );
  XOR2_X1 U436 ( .A1(Key[51]), .A2(Plaintext[51]), .Z(n333) );
  XOR2_X1 U437 ( .A1(Key[53]), .A2(Plaintext[53]), .Z(n389) );
  XOR2_X1 U438 ( .A1(Key[54]), .A2(Plaintext[54]), .Z(n271) );
  XOR2_X1 U439 ( .A1(Key[55]), .A2(Plaintext[55]), .Z(n230) );
  XOR2_X1 U440 ( .A1(Key[56]), .A2(Plaintext[56]), .Z(n272) );
  XOR2_X1 U441 ( .A1(Key[57]), .A2(Plaintext[57]), .Z(n335) );
  XOR2_X1 U442 ( .A1(Key[58]), .A2(Plaintext[58]), .Z(n336) );
  XOR2_X1 U443 ( .A1(Key[59]), .A2(Plaintext[59]), .Z(n390) );
  XOR2_X1 U444 ( .A1(Key[60]), .A2(Plaintext[60]), .Z(n273) );
  XOR2_X1 U445 ( .A1(Key[61]), .A2(Plaintext[61]), .Z(n231) );
  XOR2_X1 U446 ( .A1(Key[62]), .A2(Plaintext[62]), .Z(n274) );
  XOR2_X1 U447 ( .A1(Key[63]), .A2(Plaintext[63]), .Z(n337) );
  XOR2_X1 U448 ( .A1(Key[64]), .A2(Plaintext[64]), .Z(n338) );
  XOR2_X1 U449 ( .A1(Key[65]), .A2(Plaintext[65]), .Z(n391) );
  XOR2_X1 U450 ( .A1(Key[66]), .A2(Plaintext[66]), .Z(n275) );
  XOR2_X1 U451 ( .A1(Key[67]), .A2(Plaintext[67]), .Z(n232) );
  XOR2_X1 U452 ( .A1(Key[68]), .A2(Plaintext[68]), .Z(n276) );
  XOR2_X1 U453 ( .A1(Key[69]), .A2(Plaintext[69]), .Z(n339) );
  XOR2_X1 U454 ( .A1(Key[70]), .A2(Plaintext[70]), .Z(n340) );
  XOR2_X1 U455 ( .A1(Key[71]), .A2(Plaintext[71]), .Z(n392) );
  XOR2_X1 U456 ( .A1(Key[72]), .A2(Plaintext[72]), .Z(n277) );
  XOR2_X1 U457 ( .A1(Key[73]), .A2(Plaintext[73]), .Z(n233) );
  XOR2_X1 U458 ( .A1(Key[74]), .A2(Plaintext[74]), .Z(n278) );
  XOR2_X1 U459 ( .A1(Key[75]), .A2(Plaintext[75]), .Z(n341) );
  XOR2_X1 U460 ( .A1(Key[77]), .A2(Plaintext[77]), .Z(n393) );
  XOR2_X1 U461 ( .A1(Key[78]), .A2(Plaintext[78]), .Z(n279) );
  XOR2_X1 U462 ( .A1(Key[79]), .A2(Plaintext[79]), .Z(n234) );
  XOR2_X1 U463 ( .A1(Key[80]), .A2(Plaintext[80]), .Z(n280) );
  XOR2_X1 U464 ( .A1(Key[81]), .A2(Plaintext[81]), .Z(n343) );
  XOR2_X1 U465 ( .A1(Key[82]), .A2(Plaintext[82]), .Z(n344) );
  XOR2_X1 U466 ( .A1(Key[83]), .A2(Plaintext[83]), .Z(n394) );
  XOR2_X1 U467 ( .A1(Key[84]), .A2(Plaintext[84]), .Z(n281) );
  XOR2_X1 U468 ( .A1(Key[85]), .A2(Plaintext[85]), .Z(n235) );
  XOR2_X1 U469 ( .A1(Key[86]), .A2(Plaintext[86]), .Z(n282) );
  XOR2_X1 U470 ( .A1(Key[87]), .A2(Plaintext[87]), .Z(n345) );
  XOR2_X1 U471 ( .A1(Key[88]), .A2(Plaintext[88]), .Z(n346) );
  XOR2_X1 U472 ( .A1(Key[89]), .A2(Plaintext[89]), .Z(n395) );
  XOR2_X1 U473 ( .A1(Key[90]), .A2(Plaintext[90]), .Z(n283) );
  XOR2_X1 U474 ( .A1(Key[91]), .A2(Plaintext[91]), .Z(n236) );
  XOR2_X1 U475 ( .A1(Key[92]), .A2(Plaintext[92]), .Z(n284) );
  XOR2_X1 U476 ( .A1(Key[93]), .A2(Plaintext[93]), .Z(n347) );
  XOR2_X1 U477 ( .A1(Key[94]), .A2(Plaintext[94]), .Z(n348) );
  XOR2_X1 U478 ( .A1(Key[95]), .A2(Plaintext[95]), .Z(n396) );
  XOR2_X1 U479 ( .A1(Key[98]), .A2(Plaintext[98]), .Z(n286) );
  XOR2_X1 U480 ( .A1(Key[99]), .A2(Plaintext[99]), .Z(n349) );
  XOR2_X1 U481 ( .A1(Key[100]), .A2(Plaintext[100]), .Z(n350) );
  XOR2_X1 U482 ( .A1(Key[101]), .A2(Plaintext[101]), .Z(n397) );
  XOR2_X1 U483 ( .A1(Key[102]), .A2(Plaintext[102]), .Z(n287) );
  XOR2_X1 U484 ( .A1(Key[103]), .A2(Plaintext[103]), .Z(n238) );
  XOR2_X1 U485 ( .A1(Key[104]), .A2(Plaintext[104]), .Z(n288) );
  XOR2_X1 U486 ( .A1(Key[105]), .A2(Plaintext[105]), .Z(n351) );
  XOR2_X1 U487 ( .A1(Key[106]), .A2(Plaintext[106]), .Z(n352) );
  XOR2_X1 U488 ( .A1(Key[107]), .A2(Plaintext[107]), .Z(n398) );
  XOR2_X1 U489 ( .A1(Key[108]), .A2(Plaintext[108]), .Z(n289) );
  XOR2_X1 U490 ( .A1(Key[109]), .A2(Plaintext[109]), .Z(n239) );
  XOR2_X1 U491 ( .A1(Key[110]), .A2(Plaintext[110]), .Z(n290) );
  XOR2_X1 U492 ( .A1(Key[111]), .A2(Plaintext[111]), .Z(n353) );
  XOR2_X1 U493 ( .A1(Key[112]), .A2(Plaintext[112]), .Z(n354) );
  XOR2_X1 U494 ( .A1(Key[113]), .A2(Plaintext[113]), .Z(n399) );
  XOR2_X1 U495 ( .A1(Key[114]), .A2(Plaintext[114]), .Z(n291) );
  XOR2_X1 U496 ( .A1(Key[115]), .A2(Plaintext[115]), .Z(n240) );
  XOR2_X1 U497 ( .A1(Key[116]), .A2(Plaintext[116]), .Z(n292) );
  XOR2_X1 U498 ( .A1(Key[117]), .A2(Plaintext[117]), .Z(n355) );
  XOR2_X1 U499 ( .A1(Key[118]), .A2(Plaintext[118]), .Z(n356) );
  XOR2_X1 U500 ( .A1(Key[119]), .A2(Plaintext[119]), .Z(n400) );
  XOR2_X1 U501 ( .A1(Key[120]), .A2(Plaintext[120]), .Z(n293) );
  XOR2_X1 U502 ( .A1(Key[121]), .A2(Plaintext[121]), .Z(n241) );
  XOR2_X1 U503 ( .A1(Key[122]), .A2(Plaintext[122]), .Z(n294) );
  XOR2_X1 U504 ( .A1(Key[123]), .A2(Plaintext[123]), .Z(n357) );
  XOR2_X1 U505 ( .A1(Key[124]), .A2(Plaintext[124]), .Z(n358) );
  XOR2_X1 U506 ( .A1(Key[125]), .A2(Plaintext[125]), .Z(n401) );
  XOR2_X1 U507 ( .A1(Key[127]), .A2(Plaintext[127]), .Z(n242) );
  XOR2_X1 U508 ( .A1(Key[128]), .A2(Plaintext[128]), .Z(n296) );
  XOR2_X1 U509 ( .A1(Key[129]), .A2(Plaintext[129]), .Z(n359) );
  XOR2_X1 U510 ( .A1(Key[130]), .A2(Plaintext[130]), .Z(n360) );
  XOR2_X1 U511 ( .A1(Key[131]), .A2(Plaintext[131]), .Z(n402) );
  XOR2_X1 U512 ( .A1(Key[132]), .A2(Plaintext[132]), .Z(n297) );
  XOR2_X1 U513 ( .A1(Key[133]), .A2(Plaintext[133]), .Z(n243) );
  XOR2_X1 U514 ( .A1(Key[134]), .A2(Plaintext[134]), .Z(n298) );
  XOR2_X1 U515 ( .A1(Key[135]), .A2(Plaintext[135]), .Z(n361) );
  XOR2_X1 U516 ( .A1(Key[136]), .A2(Plaintext[136]), .Z(n362) );
  XOR2_X1 U517 ( .A1(Key[137]), .A2(Plaintext[137]), .Z(n403) );
  XOR2_X1 U518 ( .A1(Key[138]), .A2(Plaintext[138]), .Z(n299) );
  XOR2_X1 U519 ( .A1(Key[139]), .A2(Plaintext[139]), .Z(n244) );
  XOR2_X1 U520 ( .A1(Key[140]), .A2(Plaintext[140]), .Z(n300) );
  XOR2_X1 U521 ( .A1(Key[141]), .A2(Plaintext[141]), .Z(n363) );
  XOR2_X1 U522 ( .A1(Key[142]), .A2(Plaintext[142]), .Z(n364) );
  XOR2_X1 U523 ( .A1(Key[143]), .A2(Plaintext[143]), .Z(n404) );
  XOR2_X1 U524 ( .A1(Key[145]), .A2(Plaintext[145]), .Z(n245) );
  XOR2_X1 U525 ( .A1(Key[146]), .A2(Plaintext[146]), .Z(n302) );
  XOR2_X1 U526 ( .A1(Key[147]), .A2(Plaintext[147]), .Z(n365) );
  XOR2_X1 U527 ( .A1(Key[148]), .A2(Plaintext[148]), .Z(n366) );
  XOR2_X1 U528 ( .A1(Key[149]), .A2(Plaintext[149]), .Z(n405) );
  XOR2_X1 U529 ( .A1(Key[150]), .A2(Plaintext[150]), .Z(n303) );
  XOR2_X1 U530 ( .A1(Key[151]), .A2(Plaintext[151]), .Z(n246) );
  XOR2_X1 U531 ( .A1(Key[152]), .A2(Plaintext[152]), .Z(n304) );
  XOR2_X1 U532 ( .A1(Key[153]), .A2(Plaintext[153]), .Z(n367) );
  XOR2_X1 U533 ( .A1(Key[154]), .A2(Plaintext[154]), .Z(n368) );
  XOR2_X1 U534 ( .A1(Key[155]), .A2(Plaintext[155]), .Z(n406) );
  XOR2_X1 U535 ( .A1(Key[156]), .A2(Plaintext[156]), .Z(n305) );
  XOR2_X1 U536 ( .A1(Key[157]), .A2(Plaintext[157]), .Z(n247) );
  XOR2_X1 U537 ( .A1(Key[158]), .A2(Plaintext[158]), .Z(n306) );
  XOR2_X1 U538 ( .A1(Key[159]), .A2(Plaintext[159]), .Z(n369) );
  XOR2_X1 U539 ( .A1(Key[160]), .A2(Plaintext[160]), .Z(n370) );
  XOR2_X1 U540 ( .A1(Key[161]), .A2(Plaintext[161]), .Z(n407) );
  XOR2_X1 U541 ( .A1(Key[162]), .A2(Plaintext[162]), .Z(n307) );
  XOR2_X1 U542 ( .A1(Key[163]), .A2(Plaintext[163]), .Z(n248) );
  XOR2_X1 U543 ( .A1(Key[164]), .A2(Plaintext[164]), .Z(n308) );
  XOR2_X1 U544 ( .A1(Key[165]), .A2(Plaintext[165]), .Z(n371) );
  XOR2_X1 U545 ( .A1(Key[166]), .A2(Plaintext[166]), .Z(n372) );
  XOR2_X1 U546 ( .A1(Key[167]), .A2(Plaintext[167]), .Z(n408) );
  XOR2_X1 U547 ( .A1(Key[168]), .A2(Plaintext[168]), .Z(n309) );
  XOR2_X1 U548 ( .A1(Key[169]), .A2(Plaintext[169]), .Z(n249) );
  XOR2_X1 U549 ( .A1(Key[170]), .A2(Plaintext[170]), .Z(n310) );
  XOR2_X1 U550 ( .A1(Key[171]), .A2(Plaintext[171]), .Z(n373) );
  XOR2_X1 U551 ( .A1(Key[172]), .A2(Plaintext[172]), .Z(n374) );
  XOR2_X1 U552 ( .A1(Key[173]), .A2(Plaintext[173]), .Z(n409) );
  XOR2_X1 U553 ( .A1(Key[174]), .A2(Plaintext[174]), .Z(n311) );
  XOR2_X1 U554 ( .A1(Key[175]), .A2(Plaintext[175]), .Z(n250) );
  XOR2_X1 U555 ( .A1(Key[176]), .A2(Plaintext[176]), .Z(n312) );
  XOR2_X1 U556 ( .A1(Key[177]), .A2(Plaintext[177]), .Z(n375) );
  XOR2_X1 U557 ( .A1(Key[178]), .A2(Plaintext[178]), .Z(n376) );
  XOR2_X1 U558 ( .A1(Key[179]), .A2(Plaintext[179]), .Z(n410) );
  XOR2_X1 U559 ( .A1(Key[180]), .A2(Plaintext[180]), .Z(n313) );
  XOR2_X1 U560 ( .A1(Key[181]), .A2(Plaintext[181]), .Z(n251) );
  XOR2_X1 U561 ( .A1(Key[182]), .A2(Plaintext[182]), .Z(n314) );
  XOR2_X1 U562 ( .A1(Key[183]), .A2(Plaintext[183]), .Z(n377) );
  XOR2_X1 U563 ( .A1(Key[184]), .A2(Plaintext[184]), .Z(n378) );
  XOR2_X1 U564 ( .A1(Key[185]), .A2(Plaintext[185]), .Z(n411) );
  XOR2_X1 U565 ( .A1(Key[186]), .A2(Plaintext[186]), .Z(n315) );
  XOR2_X1 U566 ( .A1(Key[187]), .A2(Plaintext[187]), .Z(n252) );
  XOR2_X1 U567 ( .A1(Key[188]), .A2(Plaintext[188]), .Z(n316) );
  XOR2_X1 U568 ( .A1(Key[189]), .A2(Plaintext[189]), .Z(n379) );
  XOR2_X1 U569 ( .A1(Key[190]), .A2(Plaintext[190]), .Z(n380) );
  XOR2_X1 U570 ( .A1(Key[191]), .A2(Plaintext[191]), .Z(n412) );
  BUF_X4 \SB2_3_12/BUF_5_0  ( .I(\SB2_3_12/buf_output[5] ), .Z(\RI5[3][119] )
         );
  BUF_X4 \SB2_2_23/BUF_5_0  ( .I(\SB2_2_23/buf_output[5] ), .Z(\RI5[2][53] )
         );
  NAND4_X2 \SB2_1_22/Component_Function_5/N5  ( .A1(
        \SB2_1_22/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_1_22/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_22/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_1_22/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_1_22/buf_output[5] ) );
  BUF_X4 \SB2_2_7/BUF_5_0  ( .I(\SB2_2_7/buf_output[5] ), .Z(\RI5[2][149] ) );
  INV_X2 \SB1_1_7/INV_5  ( .I(\RI1[1][149] ), .ZN(\SB1_1_7/i1_5 ) );
  BUF_X4 \SB2_2_30/BUF_5_0  ( .I(\SB2_2_30/buf_output[5] ), .Z(\RI5[2][11] )
         );
  BUF_X4 \SB2_4_8/BUF_5_0  ( .I(\SB2_4_8/buf_output[5] ), .Z(\RI5[4][143] ) );
  NAND4_X2 \SB2_1_5/Component_Function_3/N5  ( .A1(
        \SB2_1_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_5/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_5/buf_output[3] ) );
  BUF_X4 \SB2_1_5/BUF_5_0  ( .I(\SB2_1_5/buf_output[5] ), .Z(\RI5[1][161] ) );
  BUF_X4 \SB2_1_7/BUF_5_0  ( .I(\SB2_1_7/buf_output[5] ), .Z(\RI5[1][149] ) );
  BUF_X4 \SB2_2_7/BUF_3_0  ( .I(\SB2_2_7/buf_output[3] ), .Z(\RI5[2][159] ) );
  BUF_X4 \SB2_1_23/BUF_3_0  ( .I(\SB2_1_23/buf_output[3] ), .Z(\RI5[1][63] )
         );
  NAND4_X2 \SB2_1_23/Component_Function_3/N5  ( .A1(
        \SB2_1_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_23/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_23/buf_output[3] ) );
  BUF_X4 \SB2_2_12/BUF_2_0  ( .I(\SB2_2_12/buf_output[2] ), .Z(\RI5[2][134] )
         );
  INV_X2 \SB2_3_2/INV_5  ( .I(n6280), .ZN(\SB2_3_2/i1_5 ) );
  BUF_X4 \SB2_4_12/BUF_5_0  ( .I(\SB2_4_12/buf_output[5] ), .Z(\RI5[4][119] )
         );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_58  ( .I(\SB2_1_23/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[58] ) );
  BUF_X4 \SB2_3_26/BUF_5_0  ( .I(\SB2_3_26/buf_output[5] ), .Z(\RI5[3][35] )
         );
  BUF_X4 \SB2_1_23/BUF_5_0  ( .I(\SB2_1_23/buf_output[5] ), .Z(\RI5[1][53] )
         );
  NAND3_X2 \SB1_2_10/Component_Function_5/N4  ( .A1(\SB1_2_10/i0[9] ), .A2(
        \SB1_2_10/i0[6] ), .A3(\SB1_2_10/i0_4 ), .ZN(
        \SB1_2_10/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_5  ( .I(\SB2_3_31/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[5] ) );
  BUF_X4 \SB2_2_20/BUF_5_0  ( .I(\SB2_2_20/buf_output[5] ), .Z(\RI5[2][71] )
         );
  BUF_X4 \SB2_4_2/BUF_3_0  ( .I(\SB2_4_2/buf_output[3] ), .Z(\RI5[4][189] ) );
  BUF_X4 \SB2_3_26/BUF_2_0  ( .I(\SB2_3_26/buf_output[2] ), .Z(\RI5[3][50] )
         );
  NAND4_X2 \SB1_0_1/Component_Function_1/N5  ( .A1(
        \SB1_0_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_1/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_1/buf_output[1] ) );
  INV_X2 \SB2_4_29/INV_3  ( .I(\SB1_4_31/buf_output[3] ), .ZN(\SB2_4_29/i0[8] ) );
  INV_X2 \SB1_4_31/INV_5  ( .I(\RI1[4][5] ), .ZN(\SB1_4_31/i1_5 ) );
  BUF_X2 \SB2_0_28/BUF_0  ( .I(\RI3[0][18] ), .Z(\SB2_0_28/i0[9] ) );
  NAND3_X2 \SB2_2_28/Component_Function_2/N3  ( .A1(\SB2_2_28/i0_3 ), .A2(
        \SB2_2_28/i0[8] ), .A3(\SB2_2_28/i0[9] ), .ZN(
        \SB2_2_28/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 \SB2_1_9/Component_Function_3/N5  ( .A1(
        \SB2_1_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_9/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_9/buf_output[3] ) );
  BUF_X4 \SB2_2_30/BUF_4_0  ( .I(\SB2_2_30/buf_output[4] ), .Z(\RI5[2][16] )
         );
  BUF_X4 \SB2_1_8/BUF_3_0  ( .I(\SB2_1_8/buf_output[3] ), .Z(\RI5[1][153] ) );
  INV_X2 \SB1_0_28/INV_3  ( .I(n323), .ZN(\SB1_0_28/i0[8] ) );
  BUF_X4 \SB2_3_20/BUF_2_0  ( .I(\SB2_3_20/buf_output[2] ), .Z(\RI5[3][86] )
         );
  BUF_X4 \SB2_3_19/BUF_5_0  ( .I(\SB2_3_19/buf_output[5] ), .Z(\RI5[3][77] )
         );
  NAND3_X2 \SB1_2_5/Component_Function_5/N2  ( .A1(\SB1_2_5/i0_0 ), .A2(
        \SB1_2_5/i0[6] ), .A3(\SB1_2_5/i0[10] ), .ZN(
        \SB1_2_5/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB2_3_6/INV_5  ( .I(\SB1_3_6/buf_output[5] ), .ZN(\SB2_3_6/i1_5 ) );
  INV_X2 \SB2_3_15/INV_2  ( .I(\SB1_3_18/buf_output[2] ), .ZN(\SB2_3_15/i1[9] ) );
  BUF_X4 \SB2_3_6/BUF_3_0  ( .I(\SB2_3_6/buf_output[3] ), .Z(\RI5[3][165] ) );
  INV_X2 \SB2_3_6/INV_3  ( .I(\SB1_3_8/buf_output[3] ), .ZN(\SB2_3_6/i0[8] )
         );
  BUF_X4 \SB2_4_4/BUF_4_0  ( .I(\SB2_4_4/buf_output[4] ), .Z(\RI5[4][172] ) );
  BUF_X4 \SB2_3_6/BUF_1_0  ( .I(\SB2_3_6/buf_output[1] ), .Z(\RI5[3][175] ) );
  BUF_X4 \SB2_3_0/BUF_2_0  ( .I(\SB2_3_0/buf_output[2] ), .Z(\RI5[3][14] ) );
  NAND4_X2 \SB1_4_8/Component_Function_4/N5  ( .A1(
        \SB1_4_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_8/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_4_8/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_4_8/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_4_8/buf_output[4] ) );
  INV_X2 \SB1_3_3/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[173] ), .ZN(
        \SB1_3_3/i1_5 ) );
  BUF_X4 \SB2_3_16/BUF_5_0  ( .I(\SB2_3_16/buf_output[5] ), .Z(\RI5[3][95] )
         );
  NAND4_X2 \SB2_1_21/Component_Function_3/N5  ( .A1(
        \SB2_1_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_21/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_21/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_21/buf_output[3] ) );
  NAND4_X2 \SB2_4_22/Component_Function_5/N5  ( .A1(
        \SB2_4_22/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_4_22/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_4_22/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_4_22/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_4_22/buf_output[5] ) );
  BUF_X4 \SB2_2_3/BUF_4_0  ( .I(\SB2_2_3/buf_output[4] ), .Z(\RI5[2][178] ) );
  INV_X2 \SB2_1_24/INV_5  ( .I(\SB1_1_24/buf_output[5] ), .ZN(\SB2_1_24/i1_5 )
         );
  INV_X2 \SB1_2_28/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[21] ), .ZN(
        \SB1_2_28/i0[8] ) );
  NAND3_X2 \SB1_2_13/Component_Function_5/N2  ( .A1(\SB1_2_13/i0_0 ), .A2(
        \SB1_2_13/i0[6] ), .A3(\SB1_2_13/i0[10] ), .ZN(
        \SB1_2_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_3_2/Component_Function_3/N1  ( .A1(\SB2_3_2/i1[9] ), .A2(
        \SB2_3_2/i0_3 ), .A3(\SB2_3_2/i0[6] ), .ZN(
        \SB2_3_2/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_0_11/BUF_5_0  ( .I(\SB2_0_11/buf_output[5] ), .Z(\RI5[0][125] )
         );
  NAND3_X2 \SB2_1_23/Component_Function_2/N3  ( .A1(\SB2_1_23/i0_3 ), .A2(
        \SB2_1_23/i0[8] ), .A3(\SB2_1_23/i0[9] ), .ZN(
        \SB2_1_23/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_173  ( .I(\SB2_4_3/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[173] ) );
  BUF_X4 \SB2_3_18/BUF_0_0  ( .I(\SB2_3_18/buf_output[0] ), .Z(\RI5[3][108] )
         );
  BUF_X4 \SB2_2_12/BUF_0_0  ( .I(\SB2_2_12/buf_output[0] ), .Z(\RI5[2][144] )
         );
  INV_X2 \SB1_0_10/INV_3  ( .I(n359), .ZN(\SB1_0_10/i0[8] ) );
  INV_X2 \SB2_3_31/INV_3  ( .I(\SB1_3_1/buf_output[3] ), .ZN(\SB2_3_31/i0[8] )
         );
  INV_X2 \SB1_0_1/INV_3  ( .I(n377), .ZN(\SB1_0_1/i0[8] ) );
  BUF_X4 \SB2_3_10/BUF_5_0  ( .I(\SB2_3_10/buf_output[5] ), .Z(\RI5[3][131] )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_23  ( .I(\SB2_2_28/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[23] ) );
  BUF_X4 \SB1_3_7/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[149] ), .Z(
        \SB1_3_7/i0_3 ) );
  BUF_X4 \SB2_1_28/BUF_3_0  ( .I(\SB2_1_28/buf_output[3] ), .Z(\RI5[1][33] )
         );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_39  ( .I(\SB2_3_27/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[39] ) );
  BUF_X4 \SB2_3_27/BUF_5  ( .I(\SB1_3_27/buf_output[5] ), .Z(\SB2_3_27/i0_3 )
         );
  NAND3_X1 \SB1_4_14/Component_Function_1/N4  ( .A1(\SB1_4_14/i1_7 ), .A2(
        \SB1_4_14/i0[8] ), .A3(\MC_ARK_ARC_1_3/buf_output[106] ), .ZN(
        \SB1_4_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 \SB2_3_19/Component_Function_3/N4  ( .A1(\SB2_3_19/i1_5 ), .A2(
        \SB2_3_19/i0[8] ), .A3(\SB2_3_19/i3[0] ), .ZN(
        \SB2_3_19/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_3_19/BUF_3_0  ( .I(\SB2_3_19/buf_output[3] ), .Z(\RI5[3][87] )
         );
  NAND4_X2 \SB2_3_24/Component_Function_4/N5  ( .A1(
        \SB2_3_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_24/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_3_24/buf_output[4] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_65  ( .I(\SB2_2_21/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[65] ) );
  BUF_X4 \SB2_4_10/BUF_1_0  ( .I(\SB2_4_10/buf_output[1] ), .Z(\RI5[4][151] )
         );
  BUF_X4 \SB1_2_25/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[41] ), .Z(
        \SB1_2_25/i0_3 ) );
  BUF_X4 \SB2_3_14/BUF_5_0  ( .I(\SB2_3_14/buf_output[5] ), .Z(\RI5[3][107] )
         );
  BUF_X4 \SB2_1_27/BUF_1_0  ( .I(\SB2_1_27/buf_output[1] ), .Z(\RI5[1][49] )
         );
  INV_X2 \SB2_4_7/INV_3  ( .I(\SB1_4_9/buf_output[3] ), .ZN(\SB2_4_7/i0[8] )
         );
  INV_X2 \SB2_1_27/INV_5  ( .I(\SB1_1_27/buf_output[5] ), .ZN(\SB2_1_27/i1_5 )
         );
  BUF_X4 \SB2_3_15/BUF_5_0  ( .I(\SB2_3_15/buf_output[5] ), .Z(\RI5[3][101] )
         );
  INV_X2 \SB4_11/INV_2  ( .I(\SB3_14/buf_output[2] ), .ZN(\SB4_11/i1[9] ) );
  NAND4_X2 \SB2_4_10/Component_Function_0/N5  ( .A1(
        \SB2_4_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_4_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_4_10/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_4_10/buf_output[0] ) );
  INV_X2 \SB1_0_4/INV_3  ( .I(n371), .ZN(\SB1_0_4/i0[8] ) );
  BUF_X4 \SB2_2_23/BUF_0_0  ( .I(\SB2_2_23/buf_output[0] ), .Z(\RI5[2][78] )
         );
  BUF_X4 \SB1_2_23/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[53] ), .Z(
        \SB1_2_23/i0_3 ) );
  BUF_X4 \SB2_4_3/BUF_5  ( .I(\SB1_4_3/buf_output[5] ), .Z(\SB2_4_3/i0_3 ) );
  BUF_X2 \SB3_15/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[96] ), .Z(
        \SB3_15/i0[9] ) );
  CLKBUF_X4 \SB4_12/BUF_2  ( .I(\SB3_15/buf_output[2] ), .Z(\SB4_12/i0_0 ) );
  BUF_X4 \SB2_4_27/BUF_4_0  ( .I(\SB2_4_27/buf_output[4] ), .Z(\RI5[4][34] )
         );
  INV_X4 \SB1_1_21/INV_4  ( .I(\SB1_1_21/i0_4 ), .ZN(\SB1_1_21/i0[7] ) );
  BUF_X4 \SB2_3_14/BUF_4_0  ( .I(\SB2_3_14/buf_output[4] ), .Z(\RI5[3][112] )
         );
  NAND4_X2 \SB2_3_14/Component_Function_4/N5  ( .A1(
        \SB2_3_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_14/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_14/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_3_14/buf_output[4] ) );
  NAND3_X2 \SB2_4_26/Component_Function_5/N2  ( .A1(\SB2_4_26/i0_0 ), .A2(
        \SB2_4_26/i0[6] ), .A3(\SB2_4_26/i0[10] ), .ZN(
        \SB2_4_26/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_3_11/BUF_5_0  ( .I(\SB2_3_11/buf_output[5] ), .Z(\RI5[3][125] )
         );
  BUF_X4 \SB2_3_31/BUF_0_0  ( .I(\SB2_3_31/buf_output[0] ), .Z(\RI5[3][30] )
         );
  BUF_X4 \SB2_4_26/BUF_4_0  ( .I(\SB2_4_26/buf_output[4] ), .Z(\RI5[4][40] )
         );
  BUF_X4 \SB2_1_5/BUF_3_0  ( .I(\SB2_1_5/buf_output[3] ), .Z(\RI5[1][171] ) );
  INV_X2 \SB1_2_1/INV_5  ( .I(\RI1[2][185] ), .ZN(\SB1_2_1/i1_5 ) );
  NAND4_X2 \SB2_4_2/Component_Function_3/N5  ( .A1(
        \SB2_4_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_4_2/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_4_2/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_4_2/buf_output[3] ) );
  NAND4_X2 \SB2_1_8/Component_Function_4/N5  ( .A1(
        \SB2_1_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_8/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_8/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_8/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_8/buf_output[4] ) );
  BUF_X4 \SB2_4_0/BUF_4_0  ( .I(\SB2_4_0/buf_output[4] ), .Z(\RI5[4][4] ) );
  NAND3_X2 \SB1_2_13/Component_Function_1/N3  ( .A1(\SB1_2_13/i1_5 ), .A2(
        \SB1_2_13/i0[6] ), .A3(\SB1_2_13/i0[9] ), .ZN(
        \SB1_2_13/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 \SB2_3_11/BUF_4_0  ( .I(\SB2_3_11/buf_output[4] ), .Z(\RI5[3][130] )
         );
  NAND3_X2 \SB1_1_21/Component_Function_0/N4  ( .A1(\SB1_1_21/i0[7] ), .A2(
        \SB1_1_21/i0_3 ), .A3(\SB1_1_21/i0_0 ), .ZN(
        \SB1_1_21/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 \SB2_1_23/BUF_0_0  ( .I(\SB2_1_23/buf_output[0] ), .Z(\RI5[1][78] )
         );
  INV_X2 \SB1_1_25/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[39] ), .ZN(
        \SB1_1_25/i0[8] ) );
  BUF_X4 \SB1_0_12/BUF_5_0  ( .I(\SB1_0_12/buf_output[5] ), .Z(\RI3[0][119] )
         );
  BUF_X4 \SB2_3_2/BUF_5  ( .I(\SB1_3_2/buf_output[5] ), .Z(\SB2_3_2/i0_3 ) );
  INV_X2 \SB2_0_7/INV_4  ( .I(\RI3[0][148] ), .ZN(\SB2_0_7/i0[7] ) );
  BUF_X4 \SB1_0_9/BUF_5  ( .I(n403), .Z(\SB1_0_9/i0_3 ) );
  BUF_X4 \SB1_3_26/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[35] ), .Z(
        \SB1_3_26/i0_3 ) );
  NAND3_X2 \SB2_3_21/Component_Function_5/N2  ( .A1(\SB2_3_21/i0_0 ), .A2(
        \SB2_3_21/i0[6] ), .A3(\SB2_3_21/i0[10] ), .ZN(
        \SB2_3_21/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_1_8/BUF_5  ( .I(\SB1_1_8/buf_output[5] ), .Z(\SB2_1_8/i0_3 ) );
  BUF_X4 \SB2_1_22/BUF_5  ( .I(\SB1_1_22/buf_output[5] ), .Z(\SB2_1_22/i0_3 )
         );
  BUF_X4 \SB2_2_23/BUF_5  ( .I(\SB1_2_23/buf_output[5] ), .Z(\SB2_2_23/i0_3 )
         );
  BUF_X4 \SB1_1_22/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[59] ), .Z(
        \SB1_1_22/i0_3 ) );
  INV_X2 \SB4_3/INV_3  ( .I(\RI3[5][171] ), .ZN(\SB4_3/i0[8] ) );
  BUF_X4 \SB1_0_25/BUF_5  ( .I(n387), .Z(\SB1_0_25/i0_3 ) );
  CLKBUF_X4 \SB1_3_20/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[69] ), .Z(
        \SB1_3_20/i0[10] ) );
  BUF_X4 \SB2_0_13/BUF_2_0  ( .I(\SB2_0_13/buf_output[2] ), .Z(\RI5[0][128] )
         );
  BUF_X4 \SB1_3_3/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[173] ), .Z(
        \SB1_3_3/i0_3 ) );
  BUF_X4 \SB2_3_1/BUF_3_0  ( .I(\SB2_3_1/buf_output[3] ), .Z(\RI5[3][3] ) );
  BUF_X4 \SB2_0_30/BUF_5_0  ( .I(\SB2_0_30/buf_output[5] ), .Z(\RI5[0][11] )
         );
  BUF_X4 \SB2_4_0/BUF_2_0  ( .I(\SB2_4_0/buf_output[2] ), .Z(\RI5[4][14] ) );
  BUF_X4 \SB1_4_3/BUF_5  ( .I(\RI1[4][173] ), .Z(\SB1_4_3/i0_3 ) );
  BUF_X4 \SB2_1_8/BUF_4_0  ( .I(\SB2_1_8/buf_output[4] ), .Z(\RI5[1][148] ) );
  BUF_X4 \SB2_2_9/BUF_4_0  ( .I(\SB2_2_9/buf_output[4] ), .Z(\RI5[2][142] ) );
  NAND4_X2 \SB2_2_9/Component_Function_4/N5  ( .A1(
        \SB2_2_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_9/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_2_9/buf_output[4] ) );
  CLKBUF_X4 \SB1_0_29/BUF_2  ( .I(n258), .Z(\SB1_0_29/i0_0 ) );
  BUF_X4 \SB2_0_27/BUF_5_0  ( .I(\SB2_0_27/buf_output[5] ), .Z(\RI5[0][29] )
         );
  INV_X2 \SB1_1_9/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[137] ), .ZN(
        \SB1_1_9/i1_5 ) );
  NAND3_X2 \SB1_1_21/Component_Function_0/N2  ( .A1(\SB1_1_21/i0[8] ), .A2(
        \SB1_1_21/i0[7] ), .A3(\SB1_1_21/i0[6] ), .ZN(
        \SB1_1_21/Component_Function_0/NAND4_in[1] ) );
  INV_X2 \SB3_9/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[134] ), .ZN(
        \SB3_9/i1[9] ) );
  BUF_X4 \SB2_1_0/BUF_0_0  ( .I(\SB2_1_0/buf_output[0] ), .Z(\RI5[1][24] ) );
  BUF_X4 \SB2_0_23/BUF_2_0  ( .I(\SB2_0_23/buf_output[2] ), .Z(\RI5[0][68] )
         );
  BUF_X4 \SB2_1_21/BUF_1_0  ( .I(\SB2_1_21/buf_output[1] ), .Z(\RI5[1][85] )
         );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_182  ( .I(\SB2_1_4/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[182] ) );
  BUF_X4 \SB2_1_4/BUF_5  ( .I(\SB1_1_4/buf_output[5] ), .Z(\SB2_1_4/i0_3 ) );
  BUF_X4 \SB2_0_8/BUF_4_0  ( .I(\SB2_0_8/buf_output[4] ), .Z(\RI5[0][148] ) );
  NAND3_X2 \SB1_3_25/Component_Function_2/N3  ( .A1(\SB1_3_25/i0_3 ), .A2(
        \SB1_3_25/i0[8] ), .A3(\SB1_3_25/i0[9] ), .ZN(
        \SB1_3_25/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 \SB2_0_5/Component_Function_3/N5  ( .A1(
        \SB2_0_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_5/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_5/buf_output[3] ) );
  INV_X2 \SB2_1_19/INV_5  ( .I(\SB1_1_19/buf_output[5] ), .ZN(\SB2_1_19/i1_5 )
         );
  NAND4_X2 \SB2_3_6/Component_Function_1/N5  ( .A1(
        \SB2_3_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_6/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_6/buf_output[1] ) );
  NAND4_X2 \SB2_1_9/Component_Function_4/N5  ( .A1(
        \SB2_1_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_9/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_9/buf_output[4] ) );
  INV_X2 \SB1_4_19/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[77] ), .ZN(
        \SB1_4_19/i1_5 ) );
  BUF_X4 \SB2_1_25/BUF_4_0  ( .I(\SB2_1_25/buf_output[4] ), .Z(\RI5[1][46] )
         );
  BUF_X4 \SB2_0_25/BUF_0_0  ( .I(\SB2_0_25/buf_output[0] ), .Z(\RI5[0][66] )
         );
  BUF_X4 \SB2_1_7/BUF_3_0  ( .I(\SB2_1_7/buf_output[3] ), .Z(\RI5[1][159] ) );
  INV_X4 \SB2_0_21/INV_2  ( .I(\RI3[0][62] ), .ZN(\SB2_0_21/i1[9] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_77  ( .I(\SB2_4_19/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[77] ) );
  BUF_X4 \SB2_2_19/BUF_5  ( .I(\SB1_2_19/buf_output[5] ), .Z(\SB2_2_19/i0_3 )
         );
  INV_X2 \SB2_4_3/INV_3  ( .I(\SB1_4_5/buf_output[3] ), .ZN(\SB2_4_3/i0[8] )
         );
  CLKBUF_X4 \SB1_0_26/BUF_2  ( .I(n264), .Z(\SB1_0_26/i0_0 ) );
  NAND3_X2 \SB1_2_19/Component_Function_5/N3  ( .A1(\SB1_2_19/i1[9] ), .A2(
        \SB1_2_19/i0_4 ), .A3(\SB1_2_19/i0_3 ), .ZN(
        \SB1_2_19/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 \SB4_12/BUF_3  ( .I(\SB3_14/buf_output[3] ), .Z(\SB4_12/i0[10] )
         );
  NAND4_X2 \SB2_3_18/Component_Function_4/N5  ( .A1(
        \SB2_3_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_18/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_3_18/buf_output[4] ) );
  BUF_X4 \SB2_2_27/BUF_4_0  ( .I(\SB2_2_27/buf_output[4] ), .Z(\RI5[2][34] )
         );
  NAND4_X2 \SB2_2_27/Component_Function_4/N5  ( .A1(
        \SB2_2_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_27/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_27/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_27/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_2_27/buf_output[4] ) );
  BUF_X4 \SB2_0_8/BUF_2_0  ( .I(\SB2_0_8/buf_output[2] ), .Z(\RI5[0][158] ) );
  NAND4_X2 \SB1_0_13/Component_Function_0/N5  ( .A1(
        \SB1_0_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_13/buf_output[0] ) );
  BUF_X4 \SB2_4_7/BUF_0_0  ( .I(\SB2_4_7/buf_output[0] ), .Z(\RI5[4][174] ) );
  BUF_X4 \SB2_0_10/BUF_3_0  ( .I(\SB2_0_10/buf_output[3] ), .Z(\RI5[0][141] )
         );
  BUF_X4 \SB2_3_25/BUF_1_0  ( .I(\SB2_3_25/buf_output[1] ), .Z(\RI5[3][61] )
         );
  INV_X2 \SB1_4_0/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[187] ), .ZN(
        \SB1_4_0/i1_7 ) );
  INV_X2 \SB1_1_11/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[125] ), .ZN(
        \SB1_1_11/i1_5 ) );
  INV_X2 \SB1_1_12/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[117] ), .ZN(
        \SB1_1_12/i0[8] ) );
  BUF_X4 \SB2_0_16/BUF_4_0  ( .I(\SB2_0_16/buf_output[4] ), .Z(\RI5[0][100] )
         );
  NAND3_X2 \SB2_1_27/Component_Function_3/N4  ( .A1(\SB2_1_27/i1_5 ), .A2(
        \SB2_1_27/i0[8] ), .A3(\SB2_1_27/i3[0] ), .ZN(
        \SB2_1_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_3_16/Component_Function_5/N3  ( .A1(\SB1_3_16/i1[9] ), .A2(
        \SB1_3_16/i0_4 ), .A3(\SB1_3_16/i0_3 ), .ZN(
        \SB1_3_16/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB1_0_20/INV_5  ( .I(n392), .ZN(\SB1_0_20/i1_5 ) );
  BUF_X4 \SB2_0_15/BUF_5_0  ( .I(\SB2_0_15/buf_output[5] ), .Z(\RI5[0][101] )
         );
  INV_X2 \SB2_2_0/INV_4  ( .I(n5444), .ZN(\SB2_2_0/i0[7] ) );
  NAND3_X2 \SB2_2_30/Component_Function_2/N3  ( .A1(\SB2_2_30/i0_3 ), .A2(
        \SB2_2_30/i0[8] ), .A3(\SB2_2_30/i0[9] ), .ZN(
        \SB2_2_30/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB2_0_8/BUF_5_0  ( .I(\SB2_0_8/buf_output[5] ), .Z(\RI5[0][143] ) );
  NAND3_X2 \SB2_0_18/Component_Function_2/N1  ( .A1(\SB2_0_18/i1_5 ), .A2(
        \SB2_0_18/i0[10] ), .A3(\SB2_0_18/i1[9] ), .ZN(
        \SB2_0_18/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_0_16/BUF_3_0  ( .I(\SB2_0_16/buf_output[3] ), .Z(\RI5[0][105] )
         );
  BUF_X4 \SB2_0_16/BUF_5_0  ( .I(\SB2_0_16/buf_output[5] ), .Z(\RI5[0][95] )
         );
  INV_X2 \SB1_4_29/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[15] ), .ZN(
        \SB1_4_29/i0[8] ) );
  BUF_X4 \SB2_1_13/BUF_4_0  ( .I(\SB2_1_13/buf_output[4] ), .Z(\RI5[1][118] )
         );
  NAND4_X2 \SB2_1_14/Component_Function_1/N5  ( .A1(
        \SB2_1_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_14/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_1_14/buf_output[1] ) );
  BUF_X4 \SB2_0_8/BUF_3_0  ( .I(\SB2_0_8/buf_output[3] ), .Z(\RI5[0][153] ) );
  INV_X2 \SB1_0_3/INV_2  ( .I(n310), .ZN(\SB1_0_3/i1[9] ) );
  NAND3_X2 \SB1_2_28/Component_Function_2/N3  ( .A1(\SB1_2_28/i0_3 ), .A2(
        \SB1_2_28/i0[8] ), .A3(\SB1_2_28/i0[9] ), .ZN(
        \SB1_2_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_25/Component_Function_3/N1  ( .A1(\SB2_2_25/i1[9] ), .A2(
        \SB2_2_25/i0_3 ), .A3(\SB2_2_25/i0[6] ), .ZN(
        \SB2_2_25/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_0_0/BUF_5_0  ( .I(\SB2_0_0/buf_output[5] ), .Z(\RI5[0][191] ) );
  INV_X2 \SB1_0_2/INV_5  ( .I(n410), .ZN(\SB1_0_2/i1_5 ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_87  ( .I(\SB2_4_19/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[87] ) );
  BUF_X4 \SB3_19/BUF_5  ( .I(\RI1[5][77] ), .Z(\SB3_19/i0_3 ) );
  CLKBUF_X4 \SB2_2_21/BUF_2  ( .I(\SB1_2_24/buf_output[2] ), .Z(
        \SB2_2_21/i0_0 ) );
  BUF_X4 \SB1_0_2/BUF_5  ( .I(n410), .Z(\SB1_0_2/i0_3 ) );
  INV_X2 \SB2_4_11/INV_5  ( .I(\SB1_4_11/buf_output[5] ), .ZN(\SB2_4_11/i1_5 )
         );
  BUF_X4 \SB2_3_30/BUF_4_0  ( .I(\SB2_3_30/buf_output[4] ), .Z(\RI5[3][16] )
         );
  BUF_X4 \SB2_0_7/BUF_1_0  ( .I(\SB2_0_7/buf_output[1] ), .Z(\RI5[0][169] ) );
  NAND3_X2 \SB2_2_22/Component_Function_5/N2  ( .A1(\SB2_2_22/i0_0 ), .A2(
        \SB2_2_22/i0[6] ), .A3(\SB2_2_22/i0[10] ), .ZN(
        \SB2_2_22/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB1_1_6/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[155] ), .Z(
        \SB1_1_6/i0_3 ) );
  BUF_X4 \SB1_0_24/BUF_2_0  ( .I(\SB1_0_24/buf_output[2] ), .Z(\RI3[0][62] )
         );
  BUF_X2 \SB2_1_8/BUF_2  ( .I(\SB1_1_11/buf_output[2] ), .Z(\SB2_1_8/i0_0 ) );
  BUF_X4 \SB2_1_19/BUF_5_0  ( .I(\SB2_1_19/buf_output[5] ), .Z(\RI5[1][77] )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_131  ( .I(\SB2_2_10/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[131] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_177  ( .I(\SB2_4_4/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[177] ) );
  NAND3_X2 \SB2_1_11/Component_Function_5/N2  ( .A1(\SB2_1_11/i0_0 ), .A2(
        \SB2_1_11/i0[6] ), .A3(\SB2_1_11/i0[10] ), .ZN(
        \SB2_1_11/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB1_0_28/INV_2  ( .I(n260), .ZN(\SB1_0_28/i1[9] ) );
  NAND3_X2 \SB1_1_4/Component_Function_0/N4  ( .A1(\SB1_1_4/i0[7] ), .A2(
        \SB1_1_4/i0_3 ), .A3(\SB1_1_4/i0_0 ), .ZN(
        \SB1_1_4/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 \SB2_0_23/BUF_5_0  ( .I(\SB2_0_23/buf_output[5] ), .Z(\RI5[0][53] )
         );
  NAND4_X2 \SB2_1_6/Component_Function_4/N5  ( .A1(
        \SB2_1_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_6/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_6/buf_output[4] ) );
  BUF_X4 \SB2_0_23/BUF_0_0  ( .I(\SB2_0_23/buf_output[0] ), .Z(\RI5[0][78] )
         );
  NAND3_X2 \SB2_4_4/Component_Function_2/N2  ( .A1(\SB2_4_4/i0_3 ), .A2(
        \SB2_4_4/i0[10] ), .A3(\SB2_4_4/i0[6] ), .ZN(
        \SB2_4_4/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB1_0_13/BUF_5  ( .I(n399), .Z(\SB1_0_13/i0_3 ) );
  NAND3_X2 \SB2_1_9/Component_Function_2/N3  ( .A1(\SB2_1_9/i0_3 ), .A2(
        \SB2_1_9/i0[8] ), .A3(\SB2_1_9/i0[9] ), .ZN(
        \SB2_1_9/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB1_1_30/BUF_2_0  ( .I(\SB1_1_30/buf_output[2] ), .Z(\RI3[1][26] )
         );
  INV_X2 \SB1_2_26/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[35] ), .ZN(
        \SB1_2_26/i1_5 ) );
  INV_X2 \SB1_1_20/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[71] ), .ZN(
        \SB1_1_20/i1_5 ) );
  NAND4_X2 \SB2_3_18/Component_Function_1/N5  ( .A1(
        \SB2_3_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_18/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_18/buf_output[1] ) );
  BUF_X4 \SB2_0_5/BUF_3_0  ( .I(\SB2_0_5/buf_output[3] ), .Z(\RI5[0][171] ) );
  INV_X2 \SB1_2_19/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[77] ), .ZN(
        \SB1_2_19/i1_5 ) );
  BUF_X4 \SB2_2_17/BUF_4_0  ( .I(\SB2_2_17/buf_output[4] ), .Z(\RI5[2][94] )
         );
  BUF_X4 \SB1_0_18/BUF_5  ( .I(n394), .Z(\SB1_0_18/i0_3 ) );
  INV_X2 \SB1_1_13/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[113] ), .ZN(
        \SB1_1_13/i1_5 ) );
  NAND2_X2 \SB2_2_25/Component_Function_5/N1  ( .A1(\SB2_2_25/i0_0 ), .A2(
        \SB2_2_25/i3[0] ), .ZN(\SB2_2_25/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_3_6/BUF_5  ( .I(\SB1_3_6/buf_output[5] ), .Z(\SB2_3_6/i0_3 ) );
  BUF_X4 \SB1_2_10/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[131] ), .Z(
        \SB1_2_10/i0_3 ) );
  BUF_X4 \SB2_2_30/BUF_5  ( .I(\SB1_2_30/buf_output[5] ), .Z(\SB2_2_30/i0_3 )
         );
  INV_X2 \SB2_1_18/INV_5  ( .I(\SB1_1_18/buf_output[5] ), .ZN(\SB2_1_18/i1_5 )
         );
  CLKBUF_X4 \SB4_29/BUF_4  ( .I(\SB3_30/buf_output[4] ), .Z(\SB4_29/i0_4 ) );
  NAND4_X2 \SB2_2_10/Component_Function_0/N5  ( .A1(
        \SB2_2_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_10/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_2_10/buf_output[0] ) );
  NAND3_X2 \SB2_2_30/Component_Function_5/N4  ( .A1(\SB2_2_30/i0[9] ), .A2(
        \SB2_2_30/i0[6] ), .A3(\SB2_2_30/i0_4 ), .ZN(
        \SB2_2_30/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_31/Component_Function_2/N1  ( .A1(\SB2_2_31/i1_5 ), .A2(
        \SB2_2_31/i0[10] ), .A3(\SB2_2_31/i1[9] ), .ZN(
        \SB2_2_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_8/Component_Function_5/N2  ( .A1(\SB2_1_8/i0_0 ), .A2(
        \SB2_1_8/i0[6] ), .A3(\SB2_1_8/i0[10] ), .ZN(
        \SB2_1_8/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_0_21/BUF_2_0  ( .I(\SB2_0_21/buf_output[2] ), .Z(\RI5[0][80] )
         );
  INV_X8 \SB2_1_27/INV_2  ( .I(\RI3[1][26] ), .ZN(\SB2_1_27/i1[9] ) );
  BUF_X4 \SB2_3_5/BUF_4_0  ( .I(\SB2_3_5/buf_output[4] ), .Z(\RI5[3][166] ) );
  INV_X2 \SB1_2_24/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[43] ), .ZN(
        \SB1_2_24/i1_7 ) );
  BUF_X4 \SB2_0_28/BUF_0_0  ( .I(\SB2_0_28/buf_output[0] ), .Z(\RI5[0][48] )
         );
  INV_X2 \SB1_1_3/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[169] ), .ZN(
        \SB1_1_3/i1_7 ) );
  NAND4_X2 \SB2_1_21/Component_Function_1/N5  ( .A1(
        \SB2_1_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_21/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_1_21/buf_output[1] ) );
  BUF_X4 \SB2_3_8/BUF_0_0  ( .I(\SB2_3_8/buf_output[0] ), .Z(\RI5[3][168] ) );
  BUF_X2 \SB1_0_23/BUF_2  ( .I(n270), .Z(\SB1_0_23/i0_0 ) );
  BUF_X4 \SB2_0_12/BUF_5_0  ( .I(\SB2_0_12/buf_output[5] ), .Z(\RI5[0][119] )
         );
  BUF_X4 \SB2_1_15/BUF_5_0  ( .I(\SB2_1_15/buf_output[5] ), .Z(\RI5[1][101] )
         );
  NAND3_X2 \SB2_1_6/Component_Function_2/N3  ( .A1(\SB2_1_6/i0_3 ), .A2(
        \SB2_1_6/i0[8] ), .A3(\SB2_1_6/i0[9] ), .ZN(
        \SB2_1_6/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 \SB1_0_31/Component_Function_1/N5  ( .A1(
        \SB1_0_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_31/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_31/buf_output[1] ) );
  INV_X2 \SB1_3_6/INV_5  ( .I(n4004), .ZN(\SB1_3_6/i1_5 ) );
  INV_X2 \SB2_2_20/INV_5  ( .I(\SB1_2_20/buf_output[5] ), .ZN(\SB2_2_20/i1_5 )
         );
  BUF_X4 \SB2_1_16/BUF_5  ( .I(\SB1_1_16/buf_output[5] ), .Z(\SB2_1_16/i0_3 )
         );
  NAND4_X2 \SB1_0_3/Component_Function_0/N5  ( .A1(
        \SB1_0_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_3/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_3/buf_output[0] ) );
  NAND2_X2 \SB1_0_2/Component_Function_5/N1  ( .A1(\SB1_0_2/i0_0 ), .A2(
        \SB1_0_2/i3[0] ), .ZN(\SB1_0_2/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_0_10/BUF_4_0  ( .I(\SB2_0_10/buf_output[4] ), .Z(\RI5[0][136] )
         );
  NAND3_X2 \SB2_2_18/Component_Function_2/N3  ( .A1(\SB2_2_18/i0_3 ), .A2(
        \SB2_2_18/i0[8] ), .A3(\SB2_2_18/i0[9] ), .ZN(
        \SB2_2_18/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 \SB2_4_31/Component_Function_2/N5  ( .A1(
        \SB2_4_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_31/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_4_31/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_4_31/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_4_31/buf_output[2] ) );
  NAND4_X2 \SB2_0_26/Component_Function_5/N5  ( .A1(
        \SB2_0_26/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_0_26/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_26/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_0_26/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_0_26/buf_output[5] ) );
  BUF_X4 \SB2_3_11/BUF_0_0  ( .I(\SB2_3_11/buf_output[0] ), .Z(\RI5[3][150] )
         );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_9  ( .I(\SB2_4_0/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[9] ) );
  NAND4_X2 \SB2_4_0/Component_Function_1/N5  ( .A1(
        \SB2_4_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_0/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_4_0/buf_output[1] ) );
  INV_X2 \SB1_0_20/INV_1  ( .I(n232), .ZN(\SB1_0_20/i1_7 ) );
  INV_X2 \SB2_1_14/INV_5  ( .I(\SB1_1_14/buf_output[5] ), .ZN(\SB2_1_14/i1_5 )
         );
  BUF_X4 \SB2_3_28/BUF_3_0  ( .I(\SB2_3_28/buf_output[3] ), .Z(\RI5[3][33] )
         );
  INV_X2 \SB3_27/INV_5  ( .I(\MC_ARK_ARC_1_4/buf_output[29] ), .ZN(
        \SB3_27/i1_5 ) );
  NAND3_X2 \SB1_1_31/Component_Function_0/N4  ( .A1(\SB1_1_31/i0[7] ), .A2(
        \SB1_1_31/i0_3 ), .A3(\SB1_1_31/i0_0 ), .ZN(
        \SB1_1_31/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_149  ( .I(\RI5[0][149] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[149] ) );
  NAND3_X2 \SB3_17/Component_Function_3/N2  ( .A1(\SB3_17/i0_0 ), .A2(
        \SB3_17/i0_3 ), .A3(\SB3_17/i0_4 ), .ZN(
        \SB3_17/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 \SB1_0_26/BUF_1_0  ( .I(\SB1_0_26/buf_output[1] ), .Z(\RI3[0][55] )
         );
  INV_X2 \SB1_1_4/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[167] ), .ZN(
        \SB1_1_4/i1_5 ) );
  NAND4_X2 \SB2_2_22/Component_Function_3/N5  ( .A1(
        \SB2_2_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_22/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_2_22/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_2_22/buf_output[3] ) );
  NAND4_X2 \SB2_2_0/Component_Function_3/N5  ( .A1(
        \SB2_2_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_0/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_0/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_0/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_0/buf_output[3] ) );
  BUF_X4 \SB2_0_30/BUF_2_0  ( .I(\SB2_0_30/buf_output[2] ), .Z(\RI5[0][26] )
         );
  BUF_X2 \SB2_0_3/BUF_0_0  ( .I(\SB2_0_3/buf_output[0] ), .Z(\RI5[0][6] ) );
  BUF_X4 \SB2_2_2/BUF_4_0  ( .I(\SB2_2_2/buf_output[4] ), .Z(\RI5[2][184] ) );
  BUF_X4 \SB1_3_19/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[77] ), .Z(
        \SB1_3_19/i0_3 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_71  ( .I(\SB2_1_20/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[71] ) );
  BUF_X4 \SB2_4_12/BUF_2_0  ( .I(\SB2_4_12/buf_output[2] ), .Z(\RI5[4][134] )
         );
  NAND4_X2 \SB1_0_10/Component_Function_0/N5  ( .A1(
        \SB1_0_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_10/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_10/buf_output[0] ) );
  BUF_X4 \SB2_0_13/BUF_1_0  ( .I(\SB2_0_13/buf_output[1] ), .Z(\RI5[0][133] )
         );
  BUF_X4 \SB2_0_11/BUF_2_0  ( .I(\SB2_0_11/buf_output[2] ), .Z(\RI5[0][140] )
         );
  BUF_X4 \SB2_0_6/BUF_3_0  ( .I(\SB2_0_6/buf_output[3] ), .Z(\RI5[0][165] ) );
  NAND3_X2 \SB2_3_22/Component_Function_2/N3  ( .A1(\SB2_3_22/i0_3 ), .A2(
        \SB2_3_22/i0[8] ), .A3(\SB2_3_22/i0[9] ), .ZN(
        \SB2_3_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_12/Component_Function_2/N3  ( .A1(\SB2_2_12/i0_3 ), .A2(
        \SB2_2_12/i0[8] ), .A3(\SB2_2_12/i0[9] ), .ZN(
        \SB2_2_12/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB2_3_14/BUF_0_0  ( .I(\SB2_3_14/buf_output[0] ), .Z(\RI5[3][132] )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_29  ( .I(\SB2_2_27/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[29] ) );
  BUF_X4 \SB2_4_4/BUF_5  ( .I(\SB1_4_4/buf_output[5] ), .Z(\SB2_4_4/i0_3 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_164  ( .I(\SB2_1_7/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[164] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_98  ( .I(\SB2_2_18/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[98] ) );
  CLKBUF_X4 \SB2_0_4/BUF_2  ( .I(\SB1_0_7/buf_output[2] ), .Z(\SB2_0_4/i0_0 )
         );
  CLKBUF_X4 \SB4_6/BUF_2  ( .I(\SB3_9/buf_output[2] ), .Z(\SB4_6/i0_0 ) );
  CLKBUF_X4 \SB2_4_8/BUF_3  ( .I(\SB1_4_10/buf_output[3] ), .Z(
        \SB2_4_8/i0[10] ) );
  BUF_X4 \SB2_0_6/BUF_5_0  ( .I(\SB2_0_6/buf_output[5] ), .Z(\RI5[0][155] ) );
  BUF_X4 \SB2_0_1/BUF_3_0  ( .I(\SB2_0_1/buf_output[3] ), .Z(\RI5[0][3] ) );
  NAND4_X2 \SB2_4_10/Component_Function_1/N5  ( .A1(
        \SB2_4_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_10/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_4_10/buf_output[1] ) );
  BUF_X4 \SB2_4_13/BUF_0_0  ( .I(\SB2_4_13/buf_output[0] ), .Z(\RI5[4][138] )
         );
  BUF_X4 \SB2_2_25/BUF_0_0  ( .I(\SB2_2_25/buf_output[0] ), .Z(\RI5[2][66] )
         );
  BUF_X4 \SB2_0_23/BUF_1_0  ( .I(\SB2_0_23/buf_output[1] ), .Z(\RI5[0][73] )
         );
  NAND3_X2 \SB2_1_12/Component_Function_5/N3  ( .A1(\SB2_1_12/i1[9] ), .A2(
        \SB2_1_12/i0_4 ), .A3(\SB2_1_12/i0_3 ), .ZN(
        \SB2_1_12/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_0_6/BUF_4_0  ( .I(\SB2_0_6/buf_output[4] ), .Z(\RI5[0][160] ) );
  BUF_X2 \SB2_0_6/BUF_0  ( .I(\RI3[0][150] ), .Z(\SB2_0_6/i0[9] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_108  ( .I(\SB2_1_18/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[108] ) );
  BUF_X4 \SB1_2_31/BUF_5  ( .I(\RI1[2][5] ), .Z(\SB1_2_31/i0_3 ) );
  BUF_X4 \SB1_2_3/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[173] ), .Z(
        \SB1_2_3/i0_3 ) );
  NAND3_X1 \SB2_4_8/Component_Function_5/N3  ( .A1(\SB2_4_8/i1[9] ), .A2(n3183), .A3(\SB1_4_8/buf_output[5] ), .ZN(\SB2_4_8/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_31/Component_Function_0/N2  ( .A1(\SB1_1_31/i0[8] ), .A2(
        \SB1_1_31/i0[7] ), .A3(\SB1_1_31/i0[6] ), .ZN(
        \SB1_1_31/Component_Function_0/NAND4_in[1] ) );
  BUF_X4 \SB2_1_0/BUF_5_0  ( .I(\SB2_1_0/buf_output[5] ), .Z(\RI5[1][191] ) );
  BUF_X4 \SB2_0_23/BUF_5  ( .I(\RI3[0][53] ), .Z(\SB2_0_23/i0_3 ) );
  INV_X2 \SB2_3_18/INV_5  ( .I(\SB1_3_18/buf_output[5] ), .ZN(\SB2_3_18/i1_5 )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_35  ( .I(\SB2_2_26/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[35] ) );
  BUF_X4 \SB1_2_1/BUF_5  ( .I(\RI1[2][185] ), .Z(\SB1_2_1/i0_3 ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_176  ( .I(\SB2_4_5/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[176] ) );
  BUF_X4 \SB3_25/BUF_5  ( .I(\RI1[5][41] ), .Z(\SB3_25/i0_3 ) );
  CLKBUF_X4 \SB2_4_5/BUF_3  ( .I(\SB1_4_7/buf_output[3] ), .Z(\SB2_4_5/i0[10] ) );
  CLKBUF_X4 \SB2_1_18/BUF_3  ( .I(\SB1_1_20/buf_output[3] ), .Z(
        \SB2_1_18/i0[10] ) );
  CLKBUF_X4 \SB3_29/BUF_2  ( .I(\MC_ARK_ARC_1_4/buf_output[14] ), .Z(
        \SB3_29/i0_0 ) );
  BUF_X4 \SB2_1_15/BUF_4_0  ( .I(\SB2_1_15/buf_output[4] ), .Z(\RI5[1][106] )
         );
  INV_X2 \SB2_3_25/INV_5  ( .I(\SB1_3_25/buf_output[5] ), .ZN(\SB2_3_25/i1_5 )
         );
  INV_X1 \SB1_4_8/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[143] ), .ZN(
        \SB1_4_8/i1_5 ) );
  BUF_X4 \SB2_0_4/BUF_4_0  ( .I(\SB2_0_4/buf_output[4] ), .Z(\RI5[0][172] ) );
  INV_X2 \SB2_0_15/INV_3  ( .I(\RI3[0][99] ), .ZN(\SB2_0_15/i0[8] ) );
  BUF_X4 \SB2_2_11/BUF_2_0  ( .I(\SB2_2_11/buf_output[2] ), .Z(\RI5[2][140] )
         );
  BUF_X4 \SB2_3_24/BUF_0_0  ( .I(\SB2_3_24/buf_output[0] ), .Z(\RI5[3][72] )
         );
  INV_X2 \SB1_1_14/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[107] ), .ZN(
        \SB1_1_14/i1_5 ) );
  INV_X2 \SB2_1_18/INV_1  ( .I(\SB1_1_22/buf_output[1] ), .ZN(\SB2_1_18/i1_7 )
         );
  BUF_X4 \SB2_0_30/BUF_0_0  ( .I(\SB2_0_30/buf_output[0] ), .Z(\RI5[0][36] )
         );
  INV_X2 \SB1_4_14/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[107] ), .ZN(
        \SB1_4_14/i1_5 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_62  ( .I(\SB2_1_24/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[62] ) );
  BUF_X2 U616 ( .I(Key[164]), .Z(n183) );
  BUF_X4 \SB2_4_26/BUF_0_0  ( .I(\SB2_4_26/buf_output[0] ), .Z(\RI5[4][60] )
         );
  INV_X2 \SB3_15/INV_5  ( .I(\MC_ARK_ARC_1_4/buf_output[101] ), .ZN(
        \SB3_15/i1_5 ) );
  INV_X2 \SB1_0_0/INV_3  ( .I(n379), .ZN(\SB1_0_0/i0[8] ) );
  INV_X2 \SB1_3_23/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[53] ), .ZN(
        \SB1_3_23/i1_5 ) );
  BUF_X4 \SB1_0_0/BUF_3  ( .I(n379), .Z(\SB1_0_0/i0[10] ) );
  NAND3_X2 \SB1_1_13/Component_Function_2/N3  ( .A1(\SB1_1_13/i0_3 ), .A2(
        \SB1_1_13/i0[8] ), .A3(\SB1_1_13/i0[9] ), .ZN(
        \SB1_1_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_8/Component_Function_0/N4  ( .A1(\SB1_1_8/i0[7] ), .A2(
        \SB1_1_8/i0_3 ), .A3(\SB1_1_8/i0_0 ), .ZN(
        \SB1_1_8/Component_Function_0/NAND4_in[3] ) );
  NAND2_X2 \SB1_1_16/Component_Function_5/N1  ( .A1(\SB1_1_16/i0_0 ), .A2(
        \SB1_1_16/i3[0] ), .ZN(\SB1_1_16/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_0_29/BUF_3_0  ( .I(\SB2_0_29/buf_output[3] ), .Z(\RI5[0][27] )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_100  ( .I(\SB2_2_16/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[100] ) );
  BUF_X4 \SB2_2_5/BUF_5  ( .I(\SB1_2_5/buf_output[5] ), .Z(\SB2_2_5/i0_3 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_38  ( .I(\SB2_1_28/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[38] ) );
  BUF_X4 \SB1_0_20/BUF_5_0  ( .I(\SB1_0_20/buf_output[5] ), .Z(\RI3[0][71] )
         );
  NAND3_X2 \SB2_1_28/Component_Function_2/N2  ( .A1(\SB2_1_28/i0_3 ), .A2(
        \SB2_1_28/i0[10] ), .A3(\SB2_1_28/i0[6] ), .ZN(
        \SB2_1_28/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_1_6/BUF_4_0  ( .I(\SB2_1_6/buf_output[4] ), .Z(\RI5[1][160] ) );
  INV_X2 \SB2_0_3/INV_4  ( .I(\RI3[0][172] ), .ZN(\SB2_0_3/i0[7] ) );
  BUF_X4 \SB2_2_20/BUF_4_0  ( .I(\SB2_2_20/buf_output[4] ), .Z(\RI5[2][76] )
         );
  BUF_X4 \SB1_4_21/BUF_5  ( .I(\RI1[4][65] ), .Z(\SB1_4_21/i0_3 ) );
  BUF_X4 \SB2_0_18/BUF_5  ( .I(\RI3[0][83] ), .Z(\SB2_0_18/i0_3 ) );
  BUF_X4 \SB2_0_13/BUF_4_0  ( .I(\SB2_0_13/buf_output[4] ), .Z(\RI5[0][118] )
         );
  BUF_X4 \SB2_2_17/BUF_0_0  ( .I(\SB2_2_17/buf_output[0] ), .Z(\RI5[2][114] )
         );
  NAND4_X2 \SB2_0_2/Component_Function_1/N5  ( .A1(
        \SB2_0_2/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_2/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_2/buf_output[1] ) );
  BUF_X4 \SB2_0_31/BUF_5_0  ( .I(\SB2_0_31/buf_output[5] ), .Z(\RI5[0][5] ) );
  BUF_X4 \SB2_3_2/BUF_2_0  ( .I(\SB2_3_2/buf_output[2] ), .Z(\RI5[3][2] ) );
  NAND3_X2 \SB2_1_14/Component_Function_2/N2  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i0[10] ), .A3(\SB2_1_14/i0[6] ), .ZN(
        \SB2_1_14/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_4_19/BUF_5  ( .I(\SB1_4_19/buf_output[5] ), .Z(\SB2_4_19/i0_3 )
         );
  BUF_X4 \SB2_3_25/BUF_0_0  ( .I(\SB2_3_25/buf_output[0] ), .Z(\RI5[3][66] )
         );
  BUF_X4 \SB2_0_11/BUF_0_0  ( .I(\SB2_0_11/buf_output[0] ), .Z(\RI5[0][150] )
         );
  BUF_X4 \SB2_0_22/BUF_3_0  ( .I(\SB2_0_22/buf_output[3] ), .Z(\RI5[0][69] )
         );
  NAND2_X2 \SB1_4_13/Component_Function_5/N1  ( .A1(\SB1_4_13/i0_0 ), .A2(
        \SB1_4_13/i3[0] ), .ZN(\SB1_4_13/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_1_19/BUF_0_0  ( .I(\SB2_1_19/buf_output[0] ), .Z(\RI5[1][102] )
         );
  INV_X2 \SB1_3_13/INV_5  ( .I(n4005), .ZN(\SB1_3_13/i1_5 ) );
  NAND4_X2 \SB2_0_10/Component_Function_1/N5  ( .A1(
        \SB2_0_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_10/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_10/buf_output[1] ) );
  NAND2_X2 \SB1_0_19/Component_Function_0/N1  ( .A1(\SB1_0_19/i0[10] ), .A2(
        \SB1_0_19/i0[9] ), .ZN(\SB1_0_19/Component_Function_0/NAND4_in[0] ) );
  NAND2_X2 \SB1_1_3/Component_Function_5/N1  ( .A1(\SB1_1_3/i0_0 ), .A2(
        \SB1_1_3/i3[0] ), .ZN(\SB1_1_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_19/Component_Function_2/N3  ( .A1(\SB2_3_19/i0_3 ), .A2(
        \SB2_3_19/i0[8] ), .A3(\SB2_3_19/i0[9] ), .ZN(
        \SB2_3_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_28/Component_Function_2/N2  ( .A1(\SB2_2_28/i0_3 ), .A2(
        \SB2_2_28/i0[10] ), .A3(\SB2_2_28/i0[6] ), .ZN(
        \SB2_2_28/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_162  ( .I(\SB2_2_9/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[162] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_97  ( .I(\SB2_0_19/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[97] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_86  ( .I(\SB2_4_20/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[86] ) );
  BUF_X4 \SB2_2_7/BUF_5  ( .I(\SB1_2_7/buf_output[5] ), .Z(\SB2_2_7/i0_3 ) );
  BUF_X4 \SB2_1_21/BUF_5  ( .I(\SB1_1_21/buf_output[5] ), .Z(\SB2_1_21/i0_3 )
         );
  BUF_X4 \SB2_3_7/BUF_0_0  ( .I(\SB2_3_7/buf_output[0] ), .Z(\RI5[3][174] ) );
  NAND2_X2 \SB1_2_6/Component_Function_5/N1  ( .A1(\SB1_2_6/i0_0 ), .A2(
        \SB1_2_6/i3[0] ), .ZN(\SB1_2_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_20/Component_Function_2/N3  ( .A1(\SB2_2_20/i0_3 ), .A2(
        \SB2_2_20/i0[8] ), .A3(\SB2_2_20/i0[9] ), .ZN(
        \SB2_2_20/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB2_2_0/BUF_4_0  ( .I(\SB2_2_0/buf_output[4] ), .Z(\RI5[2][4] ) );
  NAND4_X2 \SB2_4_3/Component_Function_1/N5  ( .A1(
        \SB2_4_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_3/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_4_3/buf_output[1] ) );
  INV_X2 \SB2_3_2/INV_1  ( .I(\SB1_3_6/buf_output[1] ), .ZN(\SB2_3_2/i1_7 ) );
  BUF_X4 \SB2_0_2/BUF_2_0  ( .I(\SB2_0_2/buf_output[2] ), .Z(\RI5[0][2] ) );
  BUF_X4 \SB2_1_18/BUF_2_0  ( .I(\SB2_1_18/buf_output[2] ), .Z(\RI5[1][98] )
         );
  NAND4_X2 \SB2_0_2/Component_Function_4/N5  ( .A1(
        \SB2_0_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_2/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_2/buf_output[4] ) );
  NAND4_X2 \SB2_0_2/Component_Function_3/N5  ( .A1(
        \SB2_0_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_0_2/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_0_2/buf_output[3] ) );
  BUF_X4 \SB2_4_5/BUF_4_0  ( .I(\SB2_4_5/buf_output[4] ), .Z(\RI5[4][166] ) );
  NAND2_X2 \SB1_0_12/Component_Function_5/N1  ( .A1(\SB1_0_12/i0_0 ), .A2(
        \SB1_0_12/i3[0] ), .ZN(\SB1_0_12/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_4_6/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[151] ), .ZN(
        \SB1_4_6/i1_7 ) );
  NAND3_X2 \SB2_3_25/Component_Function_2/N2  ( .A1(\SB2_3_25/i0_3 ), .A2(
        \SB2_3_25/i0[10] ), .A3(\SB2_3_25/i0[6] ), .ZN(
        \SB2_3_25/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_102  ( .I(\SB2_0_19/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[102] ) );
  BUF_X4 \SB2_2_18/BUF_5  ( .I(\SB1_2_18/buf_output[5] ), .Z(\SB2_2_18/i0_3 )
         );
  NAND3_X2 \SB2_1_21/Component_Function_3/N1  ( .A1(\SB2_1_21/i1[9] ), .A2(
        \SB2_1_21/i0_3 ), .A3(\SB2_1_21/i0[6] ), .ZN(
        \SB2_1_21/Component_Function_3/NAND4_in[0] ) );
  CLKBUF_X4 \SB2_0_6/BUF_2  ( .I(\RI3[0][152] ), .Z(\SB2_0_6/i0_0 ) );
  NAND4_X2 \SB2_3_16/Component_Function_4/N5  ( .A1(
        \SB2_3_16/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_16/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_16/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_16/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_3_16/buf_output[4] ) );
  BUF_X4 \SB2_0_0/BUF_2_0  ( .I(\SB2_0_0/buf_output[2] ), .Z(\RI5[0][14] ) );
  BUF_X4 \SB2_3_16/BUF_4_0  ( .I(\SB2_3_16/buf_output[4] ), .Z(\RI5[3][100] )
         );
  BUF_X4 \SB2_3_19/BUF_2_0  ( .I(\SB2_3_19/buf_output[2] ), .Z(\RI5[3][92] )
         );
  NAND4_X2 \SB2_3_12/Component_Function_4/N5  ( .A1(
        \SB2_3_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_12/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_12/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_3_12/buf_output[4] ) );
  BUF_X4 \SB2_1_2/BUF_4_0  ( .I(\SB2_1_2/buf_output[4] ), .Z(\RI5[1][184] ) );
  INV_X2 \SB2_1_2/INV_4  ( .I(\SB2_1_2/i0_4 ), .ZN(\SB2_1_2/i0[7] ) );
  NAND4_X2 \SB2_4_16/Component_Function_1/N5  ( .A1(
        \SB2_4_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_16/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_4_16/buf_output[1] ) );
  INV_X2 \SB1_0_25/INV_3  ( .I(n329), .ZN(\SB1_0_25/i0[8] ) );
  BUF_X4 \SB2_2_14/BUF_5  ( .I(\SB1_2_14/buf_output[5] ), .Z(\SB2_2_14/i0_3 )
         );
  NAND3_X2 \SB2_1_31/Component_Function_2/N1  ( .A1(\SB2_1_31/i1_5 ), .A2(
        \SB2_1_31/i0[10] ), .A3(\SB2_1_31/i1[9] ), .ZN(
        \SB2_1_31/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_2_18/BUF_1_0  ( .I(\SB2_2_18/buf_output[1] ), .Z(\RI5[2][103] )
         );
  NAND3_X2 \SB1_0_13/Component_Function_3/N1  ( .A1(\SB1_0_13/i1[9] ), .A2(
        \SB1_0_13/i0_3 ), .A3(\SB1_0_13/i0[6] ), .ZN(
        \SB1_0_13/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 \SB2_0_20/Component_Function_3/N5  ( .A1(
        \SB2_0_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_20/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_20/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_20/buf_output[3] ) );
  NAND3_X2 \SB2_1_11/Component_Function_2/N1  ( .A1(\SB2_1_11/i1_5 ), .A2(
        \SB2_1_11/i0[10] ), .A3(\SB2_1_11/i1[9] ), .ZN(
        \SB2_1_11/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_1_14/BUF_0_0  ( .I(\SB2_1_14/buf_output[0] ), .Z(\RI5[1][132] )
         );
  BUF_X4 \SB2_0_24/BUF_0_0  ( .I(\SB2_0_24/buf_output[0] ), .Z(\RI5[0][72] )
         );
  NAND3_X2 \SB2_1_28/Component_Function_2/N1  ( .A1(\SB2_1_28/i1_5 ), .A2(
        \SB2_1_28/i0[10] ), .A3(\SB2_1_28/i1[9] ), .ZN(
        \SB2_1_28/Component_Function_2/NAND4_in[0] ) );
  INV_X2 \SB1_3_18/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[83] ), .ZN(
        \SB1_3_18/i1_5 ) );
  NAND2_X2 \SB2_2_12/Component_Function_5/N1  ( .A1(\SB2_2_12/i0_0 ), .A2(
        \SB2_2_12/i3[0] ), .ZN(\SB2_2_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_11/Component_Function_2/N2  ( .A1(\SB2_1_11/i0_3 ), .A2(
        \SB2_1_11/i0[10] ), .A3(\SB2_1_11/i0[6] ), .ZN(
        \SB2_1_11/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_52  ( .I(\SB2_2_24/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[52] ) );
  NAND3_X2 \SB2_3_8/Component_Function_2/N3  ( .A1(\SB2_3_8/i0_3 ), .A2(
        \SB2_3_8/i0[8] ), .A3(\SB2_3_8/i0[9] ), .ZN(
        \SB2_3_8/Component_Function_2/NAND4_in[2] ) );
  INV_X4 \SB3_6/INV_5  ( .I(\SB3_6/i0_3 ), .ZN(\SB3_6/i1_5 ) );
  INV_X2 \SB1_0_15/INV_3  ( .I(n349), .ZN(\SB1_0_15/i0[8] ) );
  NAND2_X1 \SB1_2_3/Component_Function_5/N1  ( .A1(\SB1_2_3/i0_0 ), .A2(
        \SB1_2_3/i3[0] ), .ZN(\SB1_2_3/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 \SB2_0_25/Component_Function_2/N5  ( .A1(
        \SB2_0_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_25/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_25/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_25/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_25/buf_output[2] ) );
  INV_X2 \SB1_2_17/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[89] ), .ZN(
        \SB1_2_17/i1_5 ) );
  BUF_X4 \SB2_0_24/BUF_3_0  ( .I(\SB2_0_24/buf_output[3] ), .Z(\RI5[0][57] )
         );
  INV_X2 \SB1_1_0/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[191] ), .ZN(
        \SB1_1_0/i1_5 ) );
  NAND3_X2 \SB2_2_9/Component_Function_5/N4  ( .A1(\SB2_2_9/i0[9] ), .A2(
        \SB2_2_9/i0[6] ), .A3(\SB2_2_9/i0_4 ), .ZN(
        \SB2_2_9/Component_Function_5/NAND4_in[3] ) );
  INV_X2 \SB1_0_21/INV_3  ( .I(n337), .ZN(\SB1_0_21/i0[8] ) );
  NAND3_X2 \SB1_2_3/Component_Function_2/N2  ( .A1(\SB1_2_3/i0_3 ), .A2(
        \SB1_2_3/i0[10] ), .A3(\SB1_2_3/i0[6] ), .ZN(
        \SB1_2_3/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 \SB2_0_26/Component_Function_4/N5  ( .A1(
        \SB2_0_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_26/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_26/buf_output[4] ) );
  BUF_X4 \SB2_0_16/BUF_2_0  ( .I(\SB2_0_16/buf_output[2] ), .Z(\RI5[0][110] )
         );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_154  ( .I(\SB2_4_7/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[154] ) );
  BUF_X4 \SB2_0_26/BUF_0_0  ( .I(\SB2_0_26/buf_output[0] ), .Z(\RI5[0][60] )
         );
  NAND3_X2 \SB2_2_0/Component_Function_0/N4  ( .A1(\SB2_2_0/i0[7] ), .A2(
        \SB2_2_0/i0_3 ), .A3(\SB2_2_0/i0_0 ), .ZN(
        \SB2_2_0/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 \SB2_0_26/BUF_4_0  ( .I(\SB2_0_26/buf_output[4] ), .Z(\RI5[0][40] )
         );
  BUF_X4 \SB1_0_28/BUF_3_0  ( .I(\SB1_0_28/buf_output[3] ), .Z(\RI3[0][33] )
         );
  BUF_X4 \SB2_2_3/BUF_5  ( .I(\SB1_2_3/buf_output[5] ), .Z(\SB2_2_3/i0_3 ) );
  BUF_X4 \SB1_4_20/BUF_5  ( .I(\MC_ARK_ARC_1_3/buf_output[71] ), .Z(
        \SB1_4_20/i0_3 ) );
  CLKBUF_X4 \SB1_2_17/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[87] ), .Z(
        \SB1_2_17/i0[10] ) );
  BUF_X4 \SB2_0_2/BUF_1_0  ( .I(\SB2_0_2/buf_output[1] ), .Z(\RI5[0][7] ) );
  BUF_X4 \SB2_1_15/BUF_3_0  ( .I(\SB2_1_15/buf_output[3] ), .Z(\RI5[1][111] )
         );
  BUF_X4 \SB2_2_19/BUF_1_0  ( .I(\SB2_2_19/buf_output[1] ), .Z(\RI5[2][97] )
         );
  NAND4_X2 \SB2_4_30/Component_Function_0/N5  ( .A1(
        \SB2_4_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_4_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_4_30/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_4_30/buf_output[0] ) );
  BUF_X4 \SB1_0_6/BUF_5  ( .I(n406), .Z(\SB1_0_6/i0_3 ) );
  NAND2_X2 \SB2_2_6/Component_Function_5/N1  ( .A1(\SB2_2_6/i0_0 ), .A2(
        \SB2_2_6/i3[0] ), .ZN(\SB2_2_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_28/Component_Function_3/N1  ( .A1(\SB2_2_28/i1[9] ), .A2(
        \SB2_2_28/i0_3 ), .A3(\SB2_2_28/i0[6] ), .ZN(
        \SB2_2_28/Component_Function_3/NAND4_in[0] ) );
  INV_X2 \SB1_0_1/INV_2  ( .I(n314), .ZN(\SB1_0_1/i1[9] ) );
  NAND4_X2 \SB2_1_1/Component_Function_0/N5  ( .A1(
        \SB2_1_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_1/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_1_1/buf_output[0] ) );
  BUF_X4 \SB2_0_15/BUF_4_0  ( .I(\SB2_0_15/buf_output[4] ), .Z(\RI5[0][106] )
         );
  BUF_X4 \SB2_1_25/BUF_0_0  ( .I(\SB2_1_25/buf_output[0] ), .Z(\RI5[1][66] )
         );
  BUF_X4 \SB2_1_24/BUF_3_0  ( .I(\SB2_1_24/buf_output[3] ), .Z(\RI5[1][57] )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_24  ( .I(\SB2_2_0/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[24] ) );
  INV_X2 \SB2_3_22/INV_5  ( .I(\SB1_3_22/buf_output[5] ), .ZN(\SB2_3_22/i1_5 )
         );
  BUF_X4 \SB2_0_29/BUF_5_0  ( .I(\SB2_0_29/buf_output[5] ), .Z(\RI5[0][17] )
         );
  BUF_X4 \SB2_0_31/BUF_0_0  ( .I(\SB2_0_31/buf_output[0] ), .Z(\RI5[0][30] )
         );
  INV_X2 \SB2_0_31/INV_4  ( .I(\RI3[0][4] ), .ZN(\SB2_0_31/i0[7] ) );
  BUF_X4 \SB2_3_17/BUF_5  ( .I(\SB1_3_17/buf_output[5] ), .Z(\SB2_3_17/i0_3 )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_164  ( .I(\SB2_2_7/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[164] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_170  ( .I(\SB2_3_6/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[170] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_178  ( .I(\SB2_1_3/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[178] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_141  ( .I(\SB2_3_10/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[141] ) );
  NAND4_X2 \SB2_3_31/Component_Function_1/N5  ( .A1(
        \SB2_3_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_31/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_31/buf_output[1] ) );
  NAND3_X2 \SB2_3_18/Component_Function_3/N1  ( .A1(\SB2_3_18/i1[9] ), .A2(
        \SB2_3_18/i0_3 ), .A3(\SB2_3_18/i0[6] ), .ZN(
        \SB2_3_18/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 \SB2_3_26/Component_Function_3/N5  ( .A1(
        \SB2_3_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_26/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_26/buf_output[3] ) );
  NAND4_X2 \SB2_0_20/Component_Function_1/N5  ( .A1(
        \SB2_0_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_20/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_20/buf_output[1] ) );
  INV_X2 \SB1_1_27/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[25] ), .ZN(
        \SB1_1_27/i1_7 ) );
  BUF_X4 \SB2_2_6/BUF_3_0  ( .I(\SB2_2_6/buf_output[3] ), .Z(\RI5[2][165] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_22  ( .I(\SB2_4_29/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[22] ) );
  INV_X2 \SB1_3_31/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[1] ), .ZN(
        \SB1_3_31/i1_7 ) );
  BUF_X4 \SB1_0_0/BUF_5  ( .I(n412), .Z(\SB1_0_0/i0_3 ) );
  NAND4_X2 \SB2_0_30/Component_Function_1/N5  ( .A1(
        \SB2_0_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_30/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_30/buf_output[1] ) );
  NAND4_X2 \SB2_0_7/Component_Function_4/N5  ( .A1(
        \SB2_0_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_7/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_7/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_7/buf_output[4] ) );
  BUF_X4 \SB2_0_25/BUF_2_0  ( .I(\SB2_0_25/buf_output[2] ), .Z(\RI5[0][56] )
         );
  NAND3_X2 \SB3_25/Component_Function_1/N4  ( .A1(\SB3_25/i1_7 ), .A2(
        \SB3_25/i0[8] ), .A3(\SB3_25/i0_4 ), .ZN(
        \SB3_25/Component_Function_1/NAND4_in[3] ) );
  INV_X8 \SB2_0_12/INV_5  ( .I(\RI3[0][119] ), .ZN(\SB2_0_12/i1_5 ) );
  INV_X2 \SB2_4_6/INV_5  ( .I(\SB1_4_6/buf_output[5] ), .ZN(\SB2_4_6/i1_5 ) );
  NAND3_X2 \SB2_2_8/Component_Function_2/N1  ( .A1(\SB2_2_8/i1_5 ), .A2(
        \SB2_2_8/i0[10] ), .A3(\SB2_2_8/i1[9] ), .ZN(
        \SB2_2_8/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_152  ( .I(\SB2_1_9/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[152] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_146  ( .I(\SB2_2_10/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[146] ) );
  CLKBUF_X4 \SB2_4_12/BUF_2  ( .I(\SB1_4_15/buf_output[2] ), .Z(
        \SB2_4_12/i0_0 ) );
  BUF_X4 \SB2_1_3/BUF_3_0  ( .I(\SB2_1_3/buf_output[3] ), .Z(\RI5[1][183] ) );
  BUF_X4 \SB2_3_25/BUF_2_0  ( .I(\SB2_3_25/buf_output[2] ), .Z(\RI5[3][56] )
         );
  BUF_X4 \SB2_2_20/BUF_0_0  ( .I(\SB2_2_20/buf_output[0] ), .Z(\RI5[2][96] )
         );
  BUF_X4 \SB2_3_1/BUF_0_0  ( .I(\SB2_3_1/buf_output[0] ), .Z(\RI5[3][18] ) );
  BUF_X4 \SB2_2_12/BUF_3_0  ( .I(\SB2_2_12/buf_output[3] ), .Z(\RI5[2][129] )
         );
  NAND2_X2 \SB1_1_4/Component_Function_5/N1  ( .A1(\SB1_1_4/i0_0 ), .A2(
        \SB1_1_4/i3[0] ), .ZN(\SB1_1_4/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 \SB2_1_25/Component_Function_1/N5  ( .A1(
        \SB2_1_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_25/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_1_25/buf_output[1] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_74  ( .I(\SB2_2_22/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[74] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_191_1  ( .I(\MC_ARK_ARC_1_3/buf_output[191] ), 
        .Z(\RI1[4][191] ) );
  NAND3_X2 \SB2_2_3/Component_Function_2/N3  ( .A1(\SB2_2_3/i0_3 ), .A2(n3991), 
        .A3(\SB2_2_3/i0[9] ), .ZN(\SB2_2_3/Component_Function_2/NAND4_in[2] )
         );
  BUF_X4 \SB2_0_25/BUF_1_0  ( .I(\SB2_0_25/buf_output[1] ), .Z(\RI5[0][61] )
         );
  NAND4_X2 \SB2_0_25/Component_Function_1/N5  ( .A1(
        \SB2_0_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_25/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_25/buf_output[1] ) );
  BUF_X4 \SB2_2_1/BUF_0_0  ( .I(\SB2_2_1/buf_output[0] ), .Z(\RI5[2][18] ) );
  INV_X4 \SB1_4_22/INV_5  ( .I(\RI1[4][59] ), .ZN(\SB1_4_22/i1_5 ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_63  ( .I(\SB2_2_23/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[63] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_105  ( .I(\SB2_3_16/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[105] ) );
  INV_X2 \SB2_1_13/INV_4  ( .I(n2156), .ZN(\SB2_1_13/i0[7] ) );
  NAND3_X2 \SB1_1_21/Component_Function_2/N3  ( .A1(\SB1_1_21/i0_3 ), .A2(
        \SB1_1_21/i0[8] ), .A3(\SB1_1_21/i0[9] ), .ZN(
        \SB1_1_21/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_122  ( .I(\SB2_2_14/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[122] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_56  ( .I(\SB2_2_25/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[56] ) );
  NAND3_X2 \SB2_2_7/Component_Function_3/N1  ( .A1(\SB2_2_7/i1[9] ), .A2(
        \SB2_2_7/i0_3 ), .A3(\SB2_2_7/i0[6] ), .ZN(
        \SB2_2_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_28/Component_Function_2/N1  ( .A1(\SB2_3_28/i1_5 ), .A2(
        \SB2_3_28/i0[10] ), .A3(\SB2_3_28/i1[9] ), .ZN(
        \SB2_3_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_4_21/Component_Function_3/N3  ( .A1(\SB2_4_21/i1[9] ), .A2(
        \SB2_4_21/i1_7 ), .A3(\SB2_4_21/i0[10] ), .ZN(
        \SB2_4_21/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_4  ( .I(\SB2_1_0/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[4] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_75  ( .I(\SB2_4_21/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[75] ) );
  BUF_X4 \SB1_0_19/BUF_4_0  ( .I(\SB1_0_19/buf_output[4] ), .Z(\RI3[0][82] )
         );
  INV_X2 \SB1_1_25/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[41] ), .ZN(
        \SB1_1_25/i1_5 ) );
  NAND3_X2 \SB1_0_2/Component_Function_2/N1  ( .A1(\SB1_0_2/i1_5 ), .A2(
        \SB1_0_2/i0[10] ), .A3(\SB1_0_2/i1[9] ), .ZN(
        \SB1_0_2/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_0_7/BUF_0_0  ( .I(\SB2_0_7/buf_output[0] ), .Z(\RI5[0][174] ) );
  BUF_X4 \SB2_1_25/BUF_1_0  ( .I(\SB2_1_25/buf_output[1] ), .Z(\RI5[1][61] )
         );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_176  ( .I(\SB2_3_5/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[176] ) );
  BUF_X4 \SB2_2_10/BUF_4_0  ( .I(\SB2_2_10/buf_output[4] ), .Z(\RI5[2][136] )
         );
  BUF_X4 \SB2_1_5/BUF_4_0  ( .I(\SB2_1_5/buf_output[4] ), .Z(\RI5[1][166] ) );
  INV_X2 \SB1_2_24/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[47] ), .ZN(
        \SB1_2_24/i1_5 ) );
  BUF_X4 \SB1_1_2/BUF_5  ( .I(\RI1[1][179] ), .Z(\SB1_1_2/i0_3 ) );
  CLKBUF_X4 \SB1_0_26/BUF_3  ( .I(n327), .Z(\SB1_0_26/i0[10] ) );
  INV_X2 \SB1_0_10/INV_2  ( .I(n296), .ZN(\SB1_0_10/i1[9] ) );
  BUF_X4 \SB2_0_28/BUF_5_0  ( .I(\SB2_0_28/buf_output[5] ), .Z(\RI5[0][23] )
         );
  INV_X4 \SB2_0_20/INV_5  ( .I(\RI3[0][71] ), .ZN(\SB2_0_20/i1_5 ) );
  NAND3_X2 \SB2_1_25/Component_Function_5/N4  ( .A1(\SB2_1_25/i0[9] ), .A2(
        \SB2_1_25/i0[6] ), .A3(\SB2_1_25/i0_4 ), .ZN(
        \SB2_1_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB1_4_31/Component_Function_5/N2  ( .A1(\SB1_4_31/i0_0 ), .A2(
        \SB1_4_31/i0[6] ), .A3(\SB1_4_31/i0[10] ), .ZN(
        \SB1_4_31/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_2_8/BUF_4_0  ( .I(\SB2_2_8/buf_output[4] ), .Z(\RI5[2][148] ) );
  BUF_X4 \SB2_4_20/BUF_1_0  ( .I(\SB2_4_20/buf_output[1] ), .Z(\RI5[4][91] )
         );
  BUF_X4 \SB2_3_16/BUF_0_0  ( .I(\SB2_3_16/buf_output[0] ), .Z(\RI5[3][120] )
         );
  NAND3_X2 \SB1_2_24/Component_Function_4/N3  ( .A1(\SB1_2_24/i0[9] ), .A2(
        \SB1_2_24/i0[10] ), .A3(\SB1_2_24/i0_3 ), .ZN(
        \SB1_2_24/Component_Function_4/NAND4_in[2] ) );
  INV_X2 \SB1_4_25/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[37] ), .ZN(
        \SB1_4_25/i1_7 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_0  ( .I(\SB2_1_4/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[0] ) );
  CLKBUF_X4 \SB2_1_16/BUF_0  ( .I(\SB1_1_21/buf_output[0] ), .Z(
        \SB2_1_16/i0[9] ) );
  NAND3_X2 \SB2_3_25/Component_Function_2/N4  ( .A1(\SB2_3_25/i1_5 ), .A2(
        \SB2_3_25/i0_0 ), .A3(\SB2_3_25/i0_4 ), .ZN(
        \SB2_3_25/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_117  ( .I(\SB2_1_14/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[117] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_146  ( .I(\SB2_1_10/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[146] ) );
  BUF_X4 \SB1_0_20/BUF_4_0  ( .I(\SB1_0_20/buf_output[4] ), .Z(\RI3[0][76] )
         );
  NAND3_X2 \SB2_2_12/Component_Function_2/N2  ( .A1(\SB2_2_12/i0_3 ), .A2(
        \SB2_2_12/i0[10] ), .A3(\SB2_2_12/i0[6] ), .ZN(
        \SB2_2_12/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 \SB1_3_30/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[7] ), .Z(
        \SB1_3_30/i0[6] ) );
  BUF_X4 \SB2_0_29/BUF_4_0  ( .I(\SB2_0_29/buf_output[4] ), .Z(\RI5[0][22] )
         );
  NAND4_X2 \SB2_0_29/Component_Function_4/N5  ( .A1(
        \SB2_0_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_29/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_29/buf_output[4] ) );
  BUF_X4 \SB2_1_3/BUF_0_0  ( .I(\SB2_1_3/buf_output[0] ), .Z(\RI5[1][6] ) );
  NAND2_X2 \SB2_4_18/Component_Function_5/N1  ( .A1(\SB2_4_18/i0_0 ), .A2(
        \SB2_4_18/i3[0] ), .ZN(\SB2_4_18/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_0_6/INV_3  ( .I(n367), .ZN(\SB1_0_6/i0[8] ) );
  BUF_X4 \SB2_3_1/BUF_2_0  ( .I(\SB2_3_1/buf_output[2] ), .Z(\RI5[3][8] ) );
  NAND4_X2 \SB2_0_12/Component_Function_1/N5  ( .A1(
        \SB2_0_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_12/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_12/buf_output[1] ) );
  NAND3_X2 \SB2_0_12/Component_Function_1/N3  ( .A1(\SB2_0_12/i1_5 ), .A2(
        \SB2_0_12/i0[6] ), .A3(\SB2_0_12/i0[9] ), .ZN(
        \SB2_0_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_17/Component_Function_3/N3  ( .A1(\SB2_2_17/i1[9] ), .A2(
        \SB2_2_17/i1_7 ), .A3(\SB2_2_17/i0[10] ), .ZN(
        \SB2_2_17/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_70  ( .I(\SB2_0_21/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[70] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_141  ( .I(\SB2_1_10/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[141] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_159  ( .I(\SB2_3_7/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[159] ) );
  NAND3_X2 \SB1_1_31/Component_Function_5/N3  ( .A1(\SB1_1_31/i1[9] ), .A2(
        \SB1_1_31/i0_4 ), .A3(\SB1_1_31/i0_3 ), .ZN(
        \SB1_1_31/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_17/Component_Function_3/N1  ( .A1(\SB2_3_17/i1[9] ), .A2(
        \SB2_3_17/i0_3 ), .A3(\SB2_3_17/i0[6] ), .ZN(
        \SB2_3_17/Component_Function_3/NAND4_in[0] ) );
  INV_X2 \SB1_3_8/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[143] ), .ZN(
        \SB1_3_8/i1_5 ) );
  CLKBUF_X4 \SB2_1_1/BUF_2  ( .I(\SB1_1_4/buf_output[2] ), .Z(\SB2_1_1/i0_0 )
         );
  NAND3_X2 \SB3_2/Component_Function_4/N3  ( .A1(\SB3_2/i0[9] ), .A2(
        \SB3_2/i0[10] ), .A3(\SB3_2/i0_3 ), .ZN(
        \SB3_2/Component_Function_4/NAND4_in[2] ) );
  INV_X2 \SB1_2_27/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[29] ), .ZN(
        \SB1_2_27/i1_5 ) );
  NAND4_X2 \SB2_2_15/Component_Function_2/N5  ( .A1(
        \SB2_2_15/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_15/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_15/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_2_15/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_2_15/buf_output[2] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_160  ( .I(\SB2_4_6/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[160] ) );
  NAND3_X2 \SB2_0_20/Component_Function_1/N2  ( .A1(\SB2_0_20/i0_3 ), .A2(
        \SB2_0_20/i1_7 ), .A3(\SB2_0_20/i0[8] ), .ZN(
        \SB2_0_20/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \SB2_1_27/BUF_0_0  ( .I(\SB2_1_27/buf_output[0] ), .Z(\RI5[1][54] )
         );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_7  ( .I(\SB2_3_2/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[7] ) );
  NAND4_X2 \SB1_0_9/Component_Function_4/N5  ( .A1(
        \SB1_0_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_0_9/buf_output[4] ) );
  BUF_X4 \SB2_0_8/BUF_0_0  ( .I(\SB2_0_8/buf_output[0] ), .Z(\RI5[0][168] ) );
  BUF_X4 \SB2_1_0/BUF_1_0  ( .I(\SB2_1_0/buf_output[1] ), .Z(\RI5[1][19] ) );
  BUF_X2 \SB2_0_9/BUF_1_0  ( .I(\SB2_0_9/buf_output[1] ), .Z(\RI5[0][157] ) );
  NAND3_X2 \SB1_1_17/Component_Function_5/N2  ( .A1(\SB1_1_17/i0_0 ), .A2(
        \SB1_1_17/i0[6] ), .A3(\SB1_1_17/i0[10] ), .ZN(
        \SB1_1_17/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB1_2_13/Component_Function_1/N4  ( .A1(\SB1_2_13/i1_7 ), .A2(
        \SB1_2_13/i0[8] ), .A3(\SB1_2_13/i0_4 ), .ZN(
        \SB1_2_13/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 \SB2_0_6/BUF_0_0  ( .I(\SB2_0_6/buf_output[0] ), .Z(\RI5[0][180] ) );
  INV_X2 \SB2_2_25/INV_5  ( .I(\SB1_2_25/buf_output[5] ), .ZN(\SB2_2_25/i1_5 )
         );
  BUF_X4 \SB2_0_24/BUF_4_0  ( .I(\SB2_0_24/buf_output[4] ), .Z(\RI5[0][52] )
         );
  NAND4_X2 \SB2_0_24/Component_Function_4/N5  ( .A1(
        \SB2_0_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_24/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_24/buf_output[4] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_22  ( .I(\SB2_2_29/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[22] ) );
  NAND4_X2 \SB1_0_3/Component_Function_4/N5  ( .A1(
        \SB1_0_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_3/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_3/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_0_3/buf_output[4] ) );
  NAND4_X2 \SB2_0_24/Component_Function_0/N5  ( .A1(
        \SB2_0_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_24/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_0_24/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_0_24/buf_output[0] ) );
  NAND2_X2 \SB3_12/Component_Function_5/N1  ( .A1(\SB3_12/i0_0 ), .A2(
        \SB3_12/i3[0] ), .ZN(\SB3_12/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_2_11/BUF_3_0  ( .I(\SB2_2_11/buf_output[3] ), .Z(\RI5[2][135] )
         );
  BUF_X4 \SB2_4_22/BUF_0_0  ( .I(\SB2_4_22/buf_output[0] ), .Z(\RI5[4][84] )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_28  ( .I(\SB2_2_28/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[28] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_158  ( .I(\SB2_3_8/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[158] ) );
  INV_X1 \SB3_31/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[0] ), .ZN(
        \SB3_31/i3[0] ) );
  NAND3_X2 \SB2_0_21/Component_Function_4/N1  ( .A1(\SB2_0_21/i0[9] ), .A2(
        \SB2_0_21/i0_0 ), .A3(\SB2_0_21/i0[8] ), .ZN(
        \SB2_0_21/Component_Function_4/NAND4_in[0] ) );
  INV_X4 \SB1_2_15/INV_5  ( .I(\RI1[2][101] ), .ZN(\SB1_2_15/i1_5 ) );
  BUF_X4 \SB2_0_4/BUF_5_0  ( .I(\SB2_0_4/buf_output[5] ), .Z(\RI5[0][167] ) );
  BUF_X4 \SB2_1_20/BUF_3_0  ( .I(\SB2_1_20/buf_output[3] ), .Z(\RI5[1][81] )
         );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_124  ( .I(\SB2_1_12/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[124] ) );
  NAND4_X2 \SB1_0_9/Component_Function_1/N5  ( .A1(
        \SB1_0_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_9/buf_output[1] ) );
  NAND2_X2 \SB2_1_28/Component_Function_5/N1  ( .A1(\SB2_1_28/i0_0 ), .A2(
        \SB2_1_28/i3[0] ), .ZN(\SB2_1_28/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB2_0_11/INV_5  ( .I(\RI3[0][125] ), .ZN(\SB2_0_11/i1_5 ) );
  NAND2_X2 \SB2_2_13/Component_Function_5/N1  ( .A1(\SB2_2_13/i0_0 ), .A2(
        \SB2_2_13/i3[0] ), .ZN(\SB2_2_13/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 \SB2_0_28/BUF_2  ( .I(\SB1_0_31/buf_output[2] ), .Z(
        \SB2_0_28/i0_0 ) );
  NAND3_X2 \SB2_2_19/Component_Function_3/N2  ( .A1(\SB2_2_19/i0_0 ), .A2(
        \SB2_2_19/i0_3 ), .A3(\SB2_2_19/i0_4 ), .ZN(
        \SB2_2_19/Component_Function_3/NAND4_in[1] ) );
  NAND2_X2 \SB1_3_4/Component_Function_5/N1  ( .A1(\SB1_3_4/i0_0 ), .A2(
        \SB1_3_4/i3[0] ), .ZN(\SB1_3_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_0_22/Component_Function_2/N4  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0_0 ), .A3(\SB1_0_22/i0_4 ), .ZN(
        \SB1_0_22/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 \SB2_3_16/Component_Function_1/N5  ( .A1(
        \SB2_3_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_16/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_16/buf_output[1] ) );
  NAND3_X2 \SB1_2_7/Component_Function_3/N3  ( .A1(\SB1_2_7/i1[9] ), .A2(
        \SB1_2_7/i1_7 ), .A3(\SB1_2_7/i0[10] ), .ZN(
        \SB1_2_7/Component_Function_3/NAND4_in[2] ) );
  NAND2_X2 \SB1_0_20/Component_Function_5/N1  ( .A1(\SB1_0_20/i0_0 ), .A2(
        \SB1_0_20/i3[0] ), .ZN(\SB1_0_20/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_2_1/BUF_1_0  ( .I(\SB2_2_1/buf_output[1] ), .Z(\RI5[2][13] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_71  ( .I(\SB2_0_20/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[71] ) );
  INV_X2 \SB2_4_14/INV_5  ( .I(\SB1_4_14/buf_output[5] ), .ZN(\SB2_4_14/i1_5 )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_10  ( .I(\SB2_2_31/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[10] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_150  ( .I(\SB2_2_11/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[150] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_15  ( .I(\SB2_4_31/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[15] ) );
  INV_X8 \SB1_2_12/INV_5  ( .I(\RI1[2][119] ), .ZN(\SB1_2_12/i1_5 ) );
  INV_X4 \SB1_4_0/INV_5  ( .I(\RI1[4][191] ), .ZN(\SB1_4_0/i1_5 ) );
  NAND3_X2 \SB2_1_17/Component_Function_2/N4  ( .A1(n3990), .A2(
        \SB2_1_17/i0_0 ), .A3(\SB2_1_17/i0_4 ), .ZN(
        \SB2_1_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_4_30/Component_Function_5/N3  ( .A1(\SB2_4_30/i1[9] ), .A2(
        \SB1_4_31/buf_output[4] ), .A3(\SB2_4_30/i0_3 ), .ZN(
        \SB2_4_30/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 \SB2_0_17/Component_Function_0/N5  ( .A1(
        \SB2_0_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_17/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_0_17/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_0_17/buf_output[0] ) );
  BUF_X4 \SB2_0_22/BUF_5_0  ( .I(\SB2_0_22/buf_output[5] ), .Z(\RI5[0][59] )
         );
  NAND3_X2 \SB2_0_18/Component_Function_1/N2  ( .A1(\SB2_0_18/i0_3 ), .A2(
        \SB2_0_18/i1_7 ), .A3(\SB2_0_18/i0[8] ), .ZN(
        \SB2_0_18/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_61  ( .I(\SB2_2_25/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[61] ) );
  BUF_X4 \SB2_3_7/BUF_4_0  ( .I(\SB2_3_7/buf_output[4] ), .Z(\RI5[3][154] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_94  ( .I(\SB2_3_17/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[94] ) );
  BUF_X4 \SB2_0_23/BUF_3_0  ( .I(\SB2_0_23/buf_output[3] ), .Z(\RI5[0][63] )
         );
  NAND2_X2 \SB1_1_12/Component_Function_5/N1  ( .A1(\SB1_1_12/i0_0 ), .A2(
        \SB1_1_12/i3[0] ), .ZN(\SB1_1_12/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_0_27/INV_3  ( .I(n325), .ZN(\SB1_0_27/i0[8] ) );
  BUF_X2 \SB1_0_27/BUF_1_0  ( .I(\SB1_0_27/buf_output[1] ), .Z(\RI3[0][49] )
         );
  NAND2_X2 \SB1_2_25/Component_Function_5/N1  ( .A1(\SB1_2_25/i0_0 ), .A2(
        \SB1_2_25/i3[0] ), .ZN(\SB1_2_25/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_3_6/BUF_4_0  ( .I(\SB2_3_6/buf_output[4] ), .Z(\RI5[3][160] ) );
  NAND3_X2 \SB3_17/Component_Function_0/N3  ( .A1(\SB3_17/i0[10] ), .A2(
        \SB3_17/i0_4 ), .A3(\SB3_17/i0_3 ), .ZN(
        \SB3_17/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 \SB2_0_2/BUF_5_0  ( .I(\SB2_0_2/buf_output[5] ), .Z(\RI5[0][179] ) );
  NAND3_X2 \SB2_3_15/Component_Function_1/N4  ( .A1(\SB2_3_15/i1_7 ), .A2(
        \SB2_3_15/i0[8] ), .A3(\SB2_3_15/i0_4 ), .ZN(
        \SB2_3_15/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 \SB2_2_2/BUF_0  ( .I(\SB1_2_7/buf_output[0] ), .Z(\SB2_2_2/i0[9] )
         );
  BUF_X4 \SB2_2_8/BUF_2_0  ( .I(\SB2_2_8/buf_output[2] ), .Z(\RI5[2][158] ) );
  BUF_X4 \SB2_0_7/BUF_2  ( .I(\SB1_0_10/buf_output[2] ), .Z(\SB2_0_7/i0_0 ) );
  NAND3_X2 \SB2_2_4/Component_Function_3/N4  ( .A1(\SB2_2_4/i1_5 ), .A2(
        \SB2_2_4/i0[8] ), .A3(\SB2_2_4/i3[0] ), .ZN(
        \SB2_2_4/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_177  ( .I(\SB2_1_4/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[177] ) );
  NAND3_X2 \SB2_2_3/Component_Function_2/N2  ( .A1(\SB2_2_3/i0_3 ), .A2(
        \SB2_2_3/i0[10] ), .A3(\SB2_2_3/i0[6] ), .ZN(
        \SB2_2_3/Component_Function_2/NAND4_in[1] ) );
  NAND2_X2 \SB1_3_2/Component_Function_5/N1  ( .A1(\SB1_3_2/i0_0 ), .A2(
        \SB1_3_2/i3[0] ), .ZN(\SB1_3_2/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_0_0/BUF_0_0  ( .I(\SB2_0_0/buf_output[0] ), .Z(\RI5[0][24] ) );
  INV_X2 \SB1_1_27/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[29] ), .ZN(
        \SB1_1_27/i1_5 ) );
  NAND3_X2 \SB1_1_27/Component_Function_3/N2  ( .A1(\SB1_1_27/i0_0 ), .A2(
        \SB1_1_27/i0_3 ), .A3(\SB1_1_27/i0_4 ), .ZN(
        \SB1_1_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_17/Component_Function_2/N1  ( .A1(\SB2_0_17/i1_5 ), .A2(
        \SB2_0_17/i0[10] ), .A3(\SB2_0_17/i1[9] ), .ZN(
        \SB2_0_17/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_143  ( .I(\SB2_2_8/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[143] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_140  ( .I(\SB2_3_11/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[140] ) );
  NAND4_X2 \SB1_0_21/Component_Function_1/N5  ( .A1(
        \SB1_0_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_21/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_21/buf_output[1] ) );
  NAND2_X2 \SB1_1_9/Component_Function_5/N1  ( .A1(\SB1_1_9/i0_0 ), .A2(
        \SB1_1_9/i3[0] ), .ZN(\SB1_1_9/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_3_11/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[125] ), .ZN(
        \SB1_3_11/i1_5 ) );
  INV_X2 \SB1_3_25/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[41] ), .ZN(
        \SB1_3_25/i1_5 ) );
  NAND2_X2 \SB2_0_16/Component_Function_5/N1  ( .A1(\SB2_0_16/i0_0 ), .A2(
        \SB2_0_16/i3[0] ), .ZN(\SB2_0_16/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 \SB2_4_10/BUF_0  ( .I(\SB1_4_15/buf_output[0] ), .Z(
        \SB2_4_10/i0[9] ) );
  BUF_X4 \SB2_0_19/BUF_3_0  ( .I(\SB2_0_19/buf_output[3] ), .Z(\RI5[0][87] )
         );
  NAND3_X2 \SB2_1_15/Component_Function_3/N3  ( .A1(\SB2_1_15/i1[9] ), .A2(
        \SB2_1_15/i1_7 ), .A3(\SB2_1_15/i0[10] ), .ZN(
        \SB2_1_15/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB2_4_0/BUF_0_0  ( .I(\SB2_4_0/buf_output[0] ), .Z(\RI5[4][24] ) );
  BUF_X4 \SB2_2_0/BUF_3_0  ( .I(\SB2_2_0/buf_output[3] ), .Z(\RI5[2][9] ) );
  NAND4_X2 \SB2_0_28/Component_Function_0/N5  ( .A1(
        \SB2_0_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_0_28/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_0_28/buf_output[0] ) );
  NAND3_X2 \SB2_3_6/Component_Function_2/N3  ( .A1(\SB2_3_6/i0_3 ), .A2(
        \SB2_3_6/i0[8] ), .A3(\SB2_3_6/i0[9] ), .ZN(
        \SB2_3_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB3_7/Component_Function_2/N2  ( .A1(\SB3_7/i0_3 ), .A2(
        \SB3_7/i0[10] ), .A3(\SB3_7/i0[6] ), .ZN(
        \SB3_7/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 \SB2_0_13/Component_Function_1/N5  ( .A1(
        \SB2_0_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_13/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_13/buf_output[1] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_110  ( .I(\SB2_2_16/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[110] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_3/BUF_156  ( .I(\SB2_3_10/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[156] ) );
  BUF_X4 \SB2_2_19/BUF_0_0  ( .I(\SB2_2_19/buf_output[0] ), .Z(\RI5[2][102] )
         );
  NAND3_X2 \SB1_3_7/Component_Function_3/N2  ( .A1(\SB1_3_7/i0_0 ), .A2(
        \SB1_3_7/i0_3 ), .A3(\SB1_3_7/i0_4 ), .ZN(
        \SB1_3_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_15/Component_Function_2/N1  ( .A1(\SB2_1_15/i1_5 ), .A2(
        \SB2_1_15/i0[10] ), .A3(\SB2_1_15/i1[9] ), .ZN(
        \SB2_1_15/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_14  ( .I(\SB2_2_0/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[14] ) );
  CLKBUF_X4 \SB2_4_20/BUF_2  ( .I(\SB1_4_23/buf_output[2] ), .Z(
        \SB2_4_20/i0_0 ) );
  CLKBUF_X4 \SB2_1_6/BUF_2  ( .I(\RI3[1][152] ), .Z(\SB2_1_6/i0_0 ) );
  INV_X2 \SB1_0_16/INV_2  ( .I(n284), .ZN(\SB1_0_16/i1[9] ) );
  NAND3_X2 \SB1_1_14/Component_Function_2/N2  ( .A1(\SB1_1_14/i0_3 ), .A2(
        \SB1_1_14/i0[10] ), .A3(\SB1_1_14/i0[6] ), .ZN(
        \SB1_1_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB1_2_20/Component_Function_3/N1  ( .A1(\SB1_2_20/i1[9] ), .A2(
        \SB1_2_20/i0_3 ), .A3(\SB1_2_20/i0[6] ), .ZN(
        \SB1_2_20/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_116  ( .I(\SB2_3_15/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[116] ) );
  BUF_X4 \SB2_1_15/BUF_5  ( .I(\SB1_1_15/buf_output[5] ), .Z(\SB2_1_15/i0_3 )
         );
  CLKBUF_X4 \SB2_3_24/BUF_2  ( .I(\SB1_3_27/buf_output[2] ), .Z(
        \SB2_3_24/i0_0 ) );
  NAND2_X2 \SB1_2_27/Component_Function_5/N1  ( .A1(\SB1_2_27/i0_0 ), .A2(
        \SB1_2_27/i3[0] ), .ZN(\SB1_2_27/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB1_0_24/BUF_4  ( .I(n332), .Z(\SB1_0_24/i0_4 ) );
  NAND3_X2 \SB2_1_30/Component_Function_2/N3  ( .A1(\SB2_1_30/i0_3 ), .A2(
        \SB2_1_30/i0[8] ), .A3(\SB2_1_30/i0[9] ), .ZN(
        \SB2_1_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB1_0_24/Component_Function_0/N4  ( .A1(\SB1_0_24/i0[7] ), .A2(
        \SB1_0_24/i0_3 ), .A3(\SB1_0_24/i0_0 ), .ZN(
        \SB1_0_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_1/Component_Function_3/N1  ( .A1(\SB2_2_1/i1[9] ), .A2(
        \SB2_2_1/i0_3 ), .A3(\SB2_2_1/i0[6] ), .ZN(
        \SB2_2_1/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_2_29/BUF_3_0  ( .I(\SB2_2_29/buf_output[3] ), .Z(\RI5[2][27] )
         );
  INV_X2 \SB1_0_31/INV_2  ( .I(n254), .ZN(\SB1_0_31/i1[9] ) );
  INV_X4 \SB1_0_24/INV_4  ( .I(\SB1_0_24/i0_4 ), .ZN(\SB1_0_24/i0[7] ) );
  NAND2_X2 \SB1_3_3/Component_Function_5/N1  ( .A1(\SB1_3_3/i0_0 ), .A2(
        \SB1_3_3/i3[0] ), .ZN(\SB1_3_3/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB1_1_30/BUF_5  ( .I(\RI1[1][11] ), .Z(\SB1_1_30/i0_3 ) );
  CLKBUF_X4 \SB2_0_24/BUF_3  ( .I(\SB1_0_26/buf_output[3] ), .Z(
        \SB2_0_24/i0[10] ) );
  CLKBUF_X4 \SB1_0_27/BUF_3  ( .I(n325), .Z(\SB1_0_27/i0[10] ) );
  NAND4_X2 \SB2_2_19/Component_Function_1/N5  ( .A1(
        \SB2_2_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_19/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_2_19/buf_output[1] ) );
  NAND2_X2 \SB2_3_20/Component_Function_5/N1  ( .A1(\SB2_3_20/i0_0 ), .A2(
        \SB2_3_20/i3[0] ), .ZN(\SB2_3_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_22/Component_Function_2/N1  ( .A1(\SB2_2_22/i1_5 ), .A2(
        \SB2_2_22/i0[10] ), .A3(\SB2_2_22/i1[9] ), .ZN(
        \SB2_2_22/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_172  ( .I(\SB2_2_4/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[172] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_108  ( .I(\SB2_4_18/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[108] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_62  ( .I(\SB2_3_24/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[62] ) );
  NAND4_X2 \SB2_0_19/Component_Function_3/N5  ( .A1(
        \SB2_0_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_19/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_19/buf_output[3] ) );
  NAND4_X2 \SB2_0_6/Component_Function_1/N5  ( .A1(
        \SB2_0_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_6/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_6/buf_output[1] ) );
  NAND3_X2 \SB2_4_17/Component_Function_2/N3  ( .A1(\SB2_4_17/i0_3 ), .A2(
        \SB2_4_17/i0[8] ), .A3(\SB2_4_17/i0[9] ), .ZN(
        \SB2_4_17/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB1_3_17/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[89] ), .ZN(
        \SB1_3_17/i1_5 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_162  ( .I(\SB2_1_9/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[162] ) );
  INV_X2 \SB1_0_3/INV_3  ( .I(n373), .ZN(\SB1_0_3/i0[8] ) );
  INV_X2 \SB1_0_2/INV_3  ( .I(n375), .ZN(\SB1_0_2/i0[8] ) );
  NAND4_X2 \SB2_2_29/Component_Function_1/N5  ( .A1(
        \SB2_2_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_29/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_2_29/buf_output[1] ) );
  BUF_X4 \SB2_3_15/BUF_3_0  ( .I(\SB2_3_15/buf_output[3] ), .Z(\RI5[3][111] )
         );
  BUF_X4 \SB2_0_26/BUF_2_0  ( .I(\SB2_0_26/buf_output[2] ), .Z(\RI5[0][50] )
         );
  INV_X4 \SB1_2_7/INV_5  ( .I(\RI1[2][149] ), .ZN(\SB1_2_7/i1_5 ) );
  BUF_X4 \SB2_3_4/BUF_4_0  ( .I(\SB2_3_4/buf_output[4] ), .Z(\RI5[3][172] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_45  ( .I(\SB2_4_26/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[45] ) );
  BUF_X4 \SB1_0_18/BUF_3_0  ( .I(\SB1_0_18/buf_output[3] ), .Z(\RI3[0][93] )
         );
  BUF_X4 \SB2_3_15/BUF_4_0  ( .I(\SB2_3_15/buf_output[4] ), .Z(\RI5[3][106] )
         );
  NAND3_X2 \SB2_3_14/Component_Function_2/N3  ( .A1(\SB2_3_14/i0_3 ), .A2(
        \SB2_3_14/i0[8] ), .A3(\SB2_3_14/i0[9] ), .ZN(
        \SB2_3_14/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_4/BUF_11_1  ( .I(\MC_ARK_ARC_1_4/buf_output[11] ), 
        .Z(\RI1[5][11] ) );
  CLKBUF_X2 U111 ( .I(Key[138]), .Z(n28) );
  CLKBUF_X2 U157 ( .I(Key[139]), .Z(n100) );
  INV_X1 U28 ( .I(n52), .ZN(n484) );
  CLKBUF_X1 \MC_ARK_ARC_1_0/BUF_57_0  ( .I(n162), .Z(
        \MC_ARK_ARC_1_0/buf_keyinput[57] ) );
  INV_X1 U48 ( .I(n12), .ZN(n468) );
  INV_X1 U33 ( .I(n61), .ZN(n458) );
  INV_X1 U46 ( .I(n19), .ZN(n425) );
  CLKBUF_X2 \MC_ARK_ARC_1_1/BUF_119_0  ( .I(n179), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[119] ) );
  CLKBUF_X4 \SB1_0_8/BUF_3  ( .I(n363), .Z(\SB1_0_8/i0[10] ) );
  INV_X1 U27 ( .I(n161), .ZN(n469) );
  CLKBUF_X4 \SB1_0_18/BUF_4  ( .I(n344), .Z(\SB1_0_18/i0_4 ) );
  CLKBUF_X4 \SB1_0_12/BUF_1  ( .I(n240), .Z(\SB1_0_12/i0[6] ) );
  CLKBUF_X4 \SB1_0_14/BUF_2  ( .I(n288), .Z(\SB1_0_14/i0_0 ) );
  INV_X1 U25 ( .I(n70), .ZN(n463) );
  CLKBUF_X4 \SB1_0_7/BUF_4  ( .I(n366), .Z(\SB1_0_7/i0_4 ) );
  CLKBUF_X4 \SB1_0_29/BUF_4  ( .I(n322), .Z(\SB1_0_29/i0_4 ) );
  CLKBUF_X4 \SB1_0_16/BUF_4  ( .I(n348), .Z(\SB1_0_16/i0_4 ) );
  INV_X1 U61 ( .I(n80), .ZN(n506) );
  INV_X1 U63 ( .I(n97), .ZN(n439) );
  CLKBUF_X4 \SB1_0_15/BUF_2  ( .I(n286), .Z(\SB1_0_15/i0_0 ) );
  CLKBUF_X4 \SB1_0_9/BUF_2  ( .I(n298), .Z(\SB1_0_9/i0_0 ) );
  CLKBUF_X4 \SB1_0_15/BUF_3  ( .I(n349), .Z(\SB1_0_15/i0[10] ) );
  CLKBUF_X4 \SB1_0_22/BUF_2  ( .I(n272), .Z(\SB1_0_22/i0_0 ) );
  CLKBUF_X4 \SB1_0_22/BUF_4  ( .I(n336), .Z(\SB1_0_22/i0_4 ) );
  INV_X1 U41 ( .I(n17), .ZN(n489) );
  INV_X1 U57 ( .I(n59), .ZN(n420) );
  CLKBUF_X4 \SB1_0_26/BUF_4  ( .I(n328), .Z(\SB1_0_26/i0_4 ) );
  CLKBUF_X4 \SB2_0_9/BUF_4  ( .I(\RI3[0][136] ), .Z(\SB2_0_9/i0_4 ) );
  CLKBUF_X4 \SB2_0_1/BUF_2  ( .I(\RI3[0][182] ), .Z(\SB2_0_1/i0_0 ) );
  CLKBUF_X4 \SB2_0_9/BUF_1  ( .I(\RI3[0][133] ), .Z(\SB2_0_9/i0[6] ) );
  CLKBUF_X4 \SB2_0_9/BUF_3  ( .I(\SB1_0_11/buf_output[3] ), .Z(
        \SB2_0_9/i0[10] ) );
  CLKBUF_X4 \SB2_0_30/BUF_2  ( .I(\RI3[0][8] ), .Z(\SB2_0_30/i0_0 ) );
  CLKBUF_X4 \SB2_0_29/BUF_0  ( .I(\SB1_0_2/buf_output[0] ), .Z(
        \SB2_0_29/i0[9] ) );
  CLKBUF_X4 \SB2_0_31/BUF_3  ( .I(\RI3[0][3] ), .Z(\SB2_0_31/i0[10] ) );
  CLKBUF_X4 \SB2_0_8/BUF_5  ( .I(\RI3[0][143] ), .Z(\SB2_0_8/i0_3 ) );
  BUF_X4 \SB1_0_13/BUF_4_0  ( .I(\SB1_0_13/buf_output[4] ), .Z(\RI3[0][118] )
         );
  CLKBUF_X4 \SB2_0_5/BUF_2  ( .I(\RI3[0][158] ), .Z(\SB2_0_5/i0_0 ) );
  CLKBUF_X4 \SB2_0_11/BUF_4  ( .I(\SB1_0_12/buf_output[4] ), .Z(
        \SB2_0_11/i0_4 ) );
  CLKBUF_X4 \SB2_0_10/BUF_3  ( .I(\RI3[0][129] ), .Z(\SB2_0_10/i0[10] ) );
  CLKBUF_X4 \SB2_0_31/BUF_1  ( .I(\RI3[0][1] ), .Z(\SB2_0_31/i0[6] ) );
  CLKBUF_X4 \SB2_0_16/BUF_1  ( .I(\RI3[0][91] ), .Z(\SB2_0_16/i0[6] ) );
  CLKBUF_X4 \SB2_0_6/BUF_3  ( .I(\RI3[0][153] ), .Z(\SB2_0_6/i0[10] ) );
  CLKBUF_X4 \SB2_0_15/BUF_0  ( .I(\RI3[0][96] ), .Z(\SB2_0_15/i0[9] ) );
  CLKBUF_X4 \SB2_0_3/BUF_4_0  ( .I(\SB2_0_3/buf_output[4] ), .Z(\RI5[0][178] )
         );
  CLKBUF_X4 \SB2_0_13/BUF_0_0  ( .I(\SB2_0_13/buf_output[0] ), .Z(
        \RI5[0][138] ) );
  BUF_X4 \SB2_0_9/BUF_3_0  ( .I(\SB2_0_9/buf_output[3] ), .Z(\RI5[0][147] ) );
  BUF_X4 \SB2_0_25/BUF_3_0  ( .I(\SB2_0_25/buf_output[3] ), .Z(\RI5[0][51] )
         );
  BUF_X4 \SB2_0_12/BUF_3_0  ( .I(\SB2_0_12/buf_output[3] ), .Z(\RI5[0][129] )
         );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_108  ( .I(\SB2_0_18/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[108] ) );
  CLKBUF_X4 \SB2_0_24/BUF_5_0  ( .I(\SB2_0_24/buf_output[5] ), .Z(\RI5[0][47] ) );
  CLKBUF_X4 \SB1_1_24/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[43] ), .Z(
        \SB1_1_24/i0[6] ) );
  CLKBUF_X4 \SB1_1_8/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[140] ), .Z(
        \SB1_1_8/i0_0 ) );
  CLKBUF_X4 \SB1_1_18/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[79] ), .Z(
        \SB1_1_18/i0[6] ) );
  CLKBUF_X4 \SB1_1_11/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[122] ), .Z(
        \SB1_1_11/i0_0 ) );
  CLKBUF_X4 \SB1_1_12/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[114] ), .Z(
        \SB1_1_12/i0[9] ) );
  CLKBUF_X4 \SB1_1_16/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[90] ), .Z(
        \SB1_1_16/i0[9] ) );
  CLKBUF_X4 \SB2_1_26/BUF_2  ( .I(\SB1_1_29/buf_output[2] ), .Z(
        \SB2_1_26/i0_0 ) );
  CLKBUF_X4 \SB2_1_15/BUF_0  ( .I(\SB1_1_20/buf_output[0] ), .Z(
        \SB2_1_15/i0[9] ) );
  CLKBUF_X4 \SB2_1_12/BUF_4  ( .I(\SB1_1_13/buf_output[4] ), .Z(
        \SB2_1_12/i0_4 ) );
  CLKBUF_X4 \SB2_1_5/BUF_2  ( .I(\SB1_1_8/buf_output[2] ), .Z(\SB2_1_5/i0_0 )
         );
  CLKBUF_X4 \SB2_1_4/BUF_3  ( .I(\SB1_1_6/buf_output[3] ), .Z(\SB2_1_4/i0[10] ) );
  CLKBUF_X4 \SB2_1_28/BUF_1  ( .I(\SB1_1_0/buf_output[1] ), .Z(
        \SB2_1_28/i0[6] ) );
  CLKBUF_X4 \SB2_1_7/BUF_0  ( .I(\SB1_1_12/buf_output[0] ), .Z(\SB2_1_7/i0[9] ) );
  CLKBUF_X4 \SB2_1_25/BUF_2  ( .I(\SB1_1_28/buf_output[2] ), .Z(
        \SB2_1_25/i0_0 ) );
  CLKBUF_X4 \SB2_1_10/BUF_2  ( .I(\SB1_1_13/buf_output[2] ), .Z(
        \SB2_1_10/i0_0 ) );
  CLKBUF_X4 \SB2_1_14/BUF_4  ( .I(\SB1_1_15/buf_output[4] ), .Z(
        \SB2_1_14/i0_4 ) );
  CLKBUF_X4 \SB2_1_27/BUF_0  ( .I(\SB1_1_0/buf_output[0] ), .Z(
        \SB2_1_27/i0[9] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_145  ( .I(\SB2_1_11/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[145] ) );
  BUF_X4 \SB2_1_0/BUF_3_0  ( .I(\SB2_1_0/buf_output[3] ), .Z(\RI5[1][9] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_84  ( .I(\SB2_1_22/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[84] ) );
  CLKBUF_X4 \SB1_2_0/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[188] ), .Z(
        \SB1_2_0/i0_0 ) );
  CLKBUF_X4 \SB1_2_24/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[46] ), .Z(
        \SB1_2_24/i0_4 ) );
  CLKBUF_X4 \SB1_2_20/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[67] ), .Z(
        \SB1_2_20/i0[6] ) );
  BUF_X2 \SB1_2_23/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[49] ), .Z(
        \SB1_2_23/i0[6] ) );
  CLKBUF_X4 \SB1_2_1/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[183] ), .Z(
        \SB1_2_1/i0[10] ) );
  CLKBUF_X4 \SB1_2_23/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[52] ), .Z(
        \SB1_2_23/i0_4 ) );
  CLKBUF_X4 \SB1_2_30/BUF_3  ( .I(\RI1[2][9] ), .Z(\SB1_2_30/i0[10] ) );
  CLKBUF_X4 \SB1_2_21/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[62] ), .Z(
        \SB1_2_21/i0_0 ) );
  CLKBUF_X4 \SB2_2_12/BUF_0  ( .I(\SB1_2_17/buf_output[0] ), .Z(
        \SB2_2_12/i0[9] ) );
  CLKBUF_X4 \SB2_2_28/BUF_3  ( .I(\SB1_2_30/buf_output[3] ), .Z(
        \SB2_2_28/i0[10] ) );
  CLKBUF_X4 \SB2_2_16/BUF_2  ( .I(\SB1_2_19/buf_output[2] ), .Z(
        \SB2_2_16/i0_0 ) );
  CLKBUF_X4 \SB2_2_3/BUF_4  ( .I(\SB1_2_4/buf_output[4] ), .Z(\SB2_2_3/i0_4 )
         );
  CLKBUF_X4 \SB2_2_18/BUF_3  ( .I(\SB1_2_20/buf_output[3] ), .Z(
        \SB2_2_18/i0[10] ) );
  CLKBUF_X4 \SB2_2_21/BUF_3  ( .I(\SB1_2_23/buf_output[3] ), .Z(
        \SB2_2_21/i0[10] ) );
  CLKBUF_X4 \SB2_2_18/BUF_2  ( .I(\SB1_2_21/buf_output[2] ), .Z(
        \SB2_2_18/i0_0 ) );
  CLKBUF_X4 \SB2_2_1/BUF_0  ( .I(\SB1_2_6/buf_output[0] ), .Z(\SB2_2_1/i0[9] )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_106  ( .I(\SB2_2_15/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[106] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_112  ( .I(\SB2_2_14/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[112] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_49  ( .I(\SB2_2_27/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[49] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_171  ( .I(\SB2_2_5/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[171] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_70  ( .I(\SB2_2_21/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[70] ) );
  CLKBUF_X4 \SB1_3_24/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[42] ), .Z(
        \SB1_3_24/i0[9] ) );
  CLKBUF_X4 \SB1_3_27/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[27] ), .Z(
        \SB1_3_27/i0[10] ) );
  CLKBUF_X4 \SB1_3_9/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[135] ), .Z(
        \SB1_3_9/i0[10] ) );
  CLKBUF_X4 \SB1_3_10/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[130] ), .Z(
        \SB1_3_10/i0_4 ) );
  CLKBUF_X4 \SB1_3_18/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[82] ), .Z(
        \SB1_3_18/i0_4 ) );
  CLKBUF_X4 \SB1_3_11/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[124] ), .Z(
        \SB1_3_11/i0_4 ) );
  CLKBUF_X4 \SB1_3_15/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[100] ), .Z(
        \SB1_3_15/i0_4 ) );
  CLKBUF_X4 \SB1_3_5/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[156] ), .Z(
        \SB1_3_5/i0[9] ) );
  CLKBUF_X4 \SB1_3_13/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[109] ), .Z(
        \SB1_3_13/i0[6] ) );
  CLKBUF_X4 \SB1_3_19/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[76] ), .Z(
        \SB1_3_19/i0_4 ) );
  CLKBUF_X4 \SB2_3_2/BUF_1  ( .I(\SB1_3_6/buf_output[1] ), .Z(\SB2_3_2/i0[6] )
         );
  CLKBUF_X4 \SB2_3_16/BUF_2  ( .I(\SB1_3_19/buf_output[2] ), .Z(
        \SB2_3_16/i0_0 ) );
  CLKBUF_X4 \SB2_3_31/BUF_0  ( .I(\SB1_3_4/buf_output[0] ), .Z(
        \SB2_3_31/i0[9] ) );
  CLKBUF_X4 \SB2_3_20/BUF_3  ( .I(\SB1_3_22/buf_output[3] ), .Z(
        \SB2_3_20/i0[10] ) );
  CLKBUF_X4 \SB2_3_11/BUF_0  ( .I(\SB1_3_16/buf_output[0] ), .Z(
        \SB2_3_11/i0[9] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_147  ( .I(\SB2_3_9/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[147] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_157  ( .I(\SB2_3_9/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[157] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_3/BUF_109  ( .I(\SB2_3_17/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[109] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_118  ( .I(\SB2_3_13/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[118] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_96  ( .I(\SB2_3_20/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[96] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_182  ( .I(\SB2_3_4/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[182] ) );
  CLKBUF_X4 \SB1_4_10/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[127] ), .Z(
        \SB1_4_10/i0[6] ) );
  CLKBUF_X4 \SB1_4_16/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[94] ), .Z(
        \SB1_4_16/i0_4 ) );
  CLKBUF_X4 \SB1_4_20/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[70] ), .Z(
        \SB1_4_20/i0_4 ) );
  CLKBUF_X4 \SB1_4_30/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[10] ), .Z(
        \SB1_4_30/i0_4 ) );
  CLKBUF_X4 \SB1_4_26/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[34] ), .Z(
        \SB1_4_26/i0_4 ) );
  CLKBUF_X4 \SB1_4_22/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[54] ), .Z(
        \SB1_4_22/i0[9] ) );
  CLKBUF_X4 \SB1_4_4/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[162] ), .Z(
        \SB1_4_4/i0[9] ) );
  CLKBUF_X4 \SB2_4_19/BUF_3  ( .I(\SB1_4_21/buf_output[3] ), .Z(
        \SB2_4_19/i0[10] ) );
  CLKBUF_X4 \SB2_4_9/BUF_3  ( .I(\SB1_4_11/buf_output[3] ), .Z(
        \SB2_4_9/i0[10] ) );
  CLKBUF_X4 \SB2_4_30/BUF_2  ( .I(\SB1_4_1/buf_output[2] ), .Z(\SB2_4_30/i0_0 ) );
  CLKBUF_X4 \SB2_4_23/BUF_1  ( .I(\SB1_4_27/buf_output[1] ), .Z(
        \SB2_4_23/i0[6] ) );
  CLKBUF_X4 \SB2_4_26/BUF_0  ( .I(\SB1_4_31/buf_output[0] ), .Z(
        \SB2_4_26/i0[9] ) );
  CLKBUF_X4 \SB2_4_3/BUF_0  ( .I(\SB1_4_8/buf_output[0] ), .Z(\SB2_4_3/i0[9] )
         );
  CLKBUF_X4 \SB2_4_27/BUF_0  ( .I(\SB1_4_0/buf_output[0] ), .Z(
        \SB2_4_27/i0[9] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_93  ( .I(\SB2_4_18/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[93] ) );
  BUF_X4 \SB2_4_24/BUF_3_0  ( .I(\SB2_4_24/buf_output[3] ), .Z(\RI5[4][57] )
         );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_118  ( .I(\SB2_4_13/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[118] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_2  ( .I(\SB2_4_2/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[2] ) );
  BUF_X4 \MC_ARK_ARC_1_4/BUF_55  ( .I(\SB2_4_26/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[55] ) );
  CLKBUF_X4 \SB3_9/BUF_2  ( .I(\MC_ARK_ARC_1_4/buf_output[134] ), .Z(
        \SB3_9/i0_0 ) );
  INV_X1 \SB3_20/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[66] ), .ZN(
        \SB3_20/i3[0] ) );
  BUF_X2 \SB3_20/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[66] ), .Z(
        \SB3_20/i0[9] ) );
  CLKBUF_X4 \SB4_19/BUF_4  ( .I(\SB3_20/buf_output[4] ), .Z(\SB4_19/i0_4 ) );
  BUF_X4 \SB2_0_25/BUF_4_0  ( .I(\SB2_0_25/buf_output[4] ), .Z(\RI5[0][46] )
         );
  BUF_X4 \SB2_1_6/BUF_4  ( .I(\SB1_1_7/buf_output[4] ), .Z(\SB2_1_6/i0_4 ) );
  BUF_X2 \SB1_0_0/BUF_0  ( .I(n315), .Z(\SB1_0_0/i0[9] ) );
  INV_X1 \SB1_0_24/INV_1  ( .I(n228), .ZN(\SB1_0_24/i1_7 ) );
  BUF_X2 \SB1_0_9/BUF_0  ( .I(n297), .Z(\SB1_0_9/i0[9] ) );
  NAND3_X1 \SB1_0_0/Component_Function_0/N2  ( .A1(\SB1_0_0/i0[8] ), .A2(
        \SB1_0_0/i0[7] ), .A3(\SB1_0_0/i0[6] ), .ZN(
        \SB1_0_0/Component_Function_0/NAND4_in[1] ) );
  BUF_X2 \SB1_0_11/BUF_4  ( .I(n358), .Z(\SB1_0_11/i0_4 ) );
  INV_X1 \SB1_0_25/INV_4  ( .I(n330), .ZN(\SB1_0_25/i0[7] ) );
  BUF_X2 \SB1_0_22/BUF_1  ( .I(n230), .Z(\SB1_0_22/i0[6] ) );
  INV_X1 \SB1_0_16/INV_1  ( .I(n236), .ZN(\SB1_0_16/i1_7 ) );
  INV_X1 \SB1_0_8/INV_5  ( .I(n404), .ZN(\SB1_0_8/i1_5 ) );
  INV_X1 \SB1_0_7/INV_3  ( .I(n365), .ZN(\SB1_0_7/i0[8] ) );
  NAND3_X1 \SB1_0_14/Component_Function_0/N2  ( .A1(\SB1_0_14/i0[8] ), .A2(
        \SB1_0_14/i0[7] ), .A3(\SB1_0_14/i0[6] ), .ZN(
        \SB1_0_14/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_12/Component_Function_0/N4  ( .A1(\SB1_0_12/i0[7] ), .A2(
        \SB1_0_12/i0_3 ), .A3(\SB1_0_12/i0_0 ), .ZN(
        \SB1_0_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_0/N3  ( .A1(\SB1_0_31/i0[10] ), .A2(
        \SB1_0_31/i0_4 ), .A3(\SB1_0_31/i0_3 ), .ZN(
        \SB1_0_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_6/Component_Function_4/N2  ( .A1(\SB1_0_6/i3[0] ), .A2(
        \SB1_0_6/i0_0 ), .A3(\SB1_0_6/i1_7 ), .ZN(
        \SB1_0_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_1/Component_Function_4/N2  ( .A1(\SB1_0_1/i3[0] ), .A2(
        \SB1_0_1/i0_0 ), .A3(\SB1_0_1/i1_7 ), .ZN(
        \SB1_0_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_22/Component_Function_1/N2  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i1_7 ), .A3(\SB1_0_22/i0[8] ), .ZN(
        \SB1_0_22/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_8/Component_Function_1/N4  ( .A1(\SB1_0_8/i1_7 ), .A2(
        \SB1_0_8/i0[8] ), .A3(\SB1_0_8/i0_4 ), .ZN(
        \SB1_0_8/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_25/Component_Function_5/N1  ( .A1(\SB1_0_25/i0_0 ), .A2(
        \SB1_0_25/i3[0] ), .ZN(\SB1_0_25/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_18/Component_Function_5/N1  ( .A1(n280), .A2(
        \SB1_0_18/i3[0] ), .ZN(\SB1_0_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_0/N4  ( .A1(\SB1_0_13/i0[7] ), .A2(
        \SB1_0_13/i0_3 ), .A3(\SB1_0_13/i0_0 ), .ZN(
        \SB1_0_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_3/N1  ( .A1(\SB1_0_0/i1[9] ), .A2(
        \SB1_0_0/i0_3 ), .A3(\SB1_0_0/i0[6] ), .ZN(
        \SB1_0_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_0/N4  ( .A1(\SB1_0_15/i0[7] ), .A2(
        \SB1_0_15/i0_3 ), .A3(\SB1_0_15/i0_0 ), .ZN(
        \SB1_0_15/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_14/Component_Function_1/N1  ( .A1(\SB1_0_14/i0_3 ), .A2(
        \SB1_0_14/i1[9] ), .ZN(\SB1_0_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_2/N2  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i0[10] ), .A3(\SB1_0_9/i0[6] ), .ZN(
        \SB1_0_9/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_20/Component_Function_0/N1  ( .A1(\SB1_0_20/i0[10] ), .A2(
        \SB1_0_20/i0[9] ), .ZN(\SB1_0_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_24/Component_Function_1/N1  ( .A1(\SB1_0_24/i0_3 ), .A2(
        \SB1_0_24/i1[9] ), .ZN(\SB1_0_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_5/N2  ( .A1(\SB1_0_15/i0_0 ), .A2(
        \SB1_0_15/i0[6] ), .A3(\SB1_0_15/i0[10] ), .ZN(
        \SB1_0_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_12/Component_Function_1/N1  ( .A1(\SB1_0_12/i0_3 ), .A2(
        \SB1_0_12/i1[9] ), .ZN(\SB1_0_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_1/N4  ( .A1(\SB1_0_14/i1_7 ), .A2(
        \SB1_0_14/i0[8] ), .A3(n352), .ZN(
        \SB1_0_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_4/N4  ( .A1(\SB1_0_31/i1[9] ), .A2(
        \SB1_0_31/i1_5 ), .A3(\SB1_0_31/i0_4 ), .ZN(
        \SB1_0_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_4/N3  ( .A1(\SB1_0_10/i0[9] ), .A2(
        \SB1_0_10/i0[10] ), .A3(\SB1_0_10/i0_3 ), .ZN(
        \SB1_0_10/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_31/Component_Function_0/N1  ( .A1(\SB1_0_31/i0[10] ), .A2(
        \SB1_0_31/i0[9] ), .ZN(\SB1_0_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_4/N3  ( .A1(\SB1_0_12/i0[9] ), .A2(
        \SB1_0_12/i0[10] ), .A3(\SB1_0_12/i0_3 ), .ZN(
        \SB1_0_12/Component_Function_4/NAND4_in[2] ) );
  BUF_X2 \SB2_0_4/BUF_1  ( .I(\RI3[0][163] ), .Z(\SB2_0_4/i0[6] ) );
  INV_X1 \SB2_0_13/INV_0  ( .I(\SB1_0_18/buf_output[0] ), .ZN(\SB2_0_13/i3[0] ) );
  INV_X1 \SB2_0_28/INV_1  ( .I(\RI3[0][19] ), .ZN(\SB2_0_28/i1_7 ) );
  BUF_X2 \SB2_0_3/BUF_0  ( .I(\SB1_0_8/buf_output[0] ), .Z(\SB2_0_3/i0[9] ) );
  BUF_X2 \SB2_0_5/BUF_1  ( .I(\SB1_0_9/buf_output[1] ), .Z(\SB2_0_5/i0[6] ) );
  BUF_X2 \SB2_0_13/BUF_0  ( .I(\SB1_0_18/buf_output[0] ), .Z(\SB2_0_13/i0[9] )
         );
  INV_X1 \SB2_0_8/INV_1  ( .I(\RI3[0][139] ), .ZN(\SB2_0_8/i1_7 ) );
  INV_X1 \SB2_0_5/INV_1  ( .I(\SB1_0_9/buf_output[1] ), .ZN(\SB2_0_5/i1_7 ) );
  INV_X1 \SB2_0_13/INV_1  ( .I(\RI3[0][109] ), .ZN(\SB2_0_13/i1_7 ) );
  INV_X1 \SB2_0_11/INV_1  ( .I(\RI3[0][121] ), .ZN(\SB2_0_11/i1_7 ) );
  INV_X1 \SB2_0_10/INV_1  ( .I(\RI3[0][127] ), .ZN(\SB2_0_10/i1_7 ) );
  INV_X1 \SB2_0_20/INV_1  ( .I(\RI3[0][67] ), .ZN(\SB2_0_20/i1_7 ) );
  NAND3_X1 \SB2_0_9/Component_Function_3/N2  ( .A1(n2886), .A2(\SB2_0_9/i0_3 ), 
        .A3(\SB2_0_9/i0_4 ), .ZN(\SB2_0_9/Component_Function_3/NAND4_in[1] )
         );
  NAND3_X1 \SB2_0_10/Component_Function_4/N2  ( .A1(\SB2_0_10/i3[0] ), .A2(
        \RI3[0][128] ), .A3(\SB2_0_10/i1_7 ), .ZN(
        \SB2_0_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_0/Component_Function_4/N4  ( .A1(\SB2_0_0/i1[9] ), .A2(
        \SB2_0_0/i1_5 ), .A3(\RI3[0][190] ), .ZN(
        \SB2_0_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_13/Component_Function_4/N1  ( .A1(\SB2_0_13/i0[9] ), .A2(
        \SB2_0_13/i0_0 ), .A3(\SB2_0_13/i0[8] ), .ZN(
        \SB2_0_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_4/N3  ( .A1(\SB2_0_10/i0[9] ), .A2(
        \SB2_0_10/i0[10] ), .A3(\SB2_0_10/i0_3 ), .ZN(
        \SB2_0_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_25/Component_Function_5/N4  ( .A1(\SB2_0_25/i0[9] ), .A2(
        \SB2_0_25/i0[6] ), .A3(\SB2_0_25/i0_4 ), .ZN(
        \SB2_0_25/Component_Function_5/NAND4_in[3] ) );
  INV_X1 \SB2_0_17/INV_0  ( .I(\SB1_0_22/buf_output[0] ), .ZN(\SB2_0_17/i3[0] ) );
  BUF_X2 \SB2_0_20/BUF_1  ( .I(\RI3[0][67] ), .Z(\SB2_0_20/i0[6] ) );
  INV_X1 \SB2_0_23/INV_4  ( .I(\SB1_0_24/buf_output[4] ), .ZN(\SB2_0_23/i0[7] ) );
  NAND3_X1 \SB2_0_30/Component_Function_3/N4  ( .A1(\SB2_0_30/i1_5 ), .A2(
        \SB2_0_30/i0[8] ), .A3(\SB2_0_30/i3[0] ), .ZN(
        \SB2_0_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_10/Component_Function_5/N2  ( .A1(\RI3[0][128] ), .A2(
        \SB2_0_10/i0[6] ), .A3(\SB2_0_10/i0[10] ), .ZN(
        \SB2_0_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_10/Component_Function_3/N4  ( .A1(\SB2_0_10/i1_5 ), .A2(
        \SB2_0_10/i0[8] ), .A3(\SB2_0_10/i3[0] ), .ZN(
        \SB2_0_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_18/Component_Function_4/N2  ( .A1(\SB2_0_18/i3[0] ), .A2(
        \SB2_0_18/i0_0 ), .A3(\SB2_0_18/i1_7 ), .ZN(
        \SB2_0_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_24/Component_Function_2/N1  ( .A1(\SB2_0_24/i1_5 ), .A2(
        \SB2_0_24/i0[10] ), .A3(\SB2_0_24/i1[9] ), .ZN(
        \SB2_0_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_2/N3  ( .A1(\SB2_0_7/i0_3 ), .A2(
        \SB2_0_7/i0[8] ), .A3(\SB2_0_7/i0[9] ), .ZN(
        \SB2_0_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_18/Component_Function_1/N3  ( .A1(\SB2_0_18/i1_5 ), .A2(
        \SB2_0_18/i0[6] ), .A3(\SB2_0_18/i0[9] ), .ZN(
        \SB2_0_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_20/Component_Function_2/N2  ( .A1(\RI3[0][71] ), .A2(
        \SB2_0_20/i0[10] ), .A3(\SB2_0_20/i0[6] ), .ZN(
        \SB2_0_20/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_8/Component_Function_1/N1  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \SB2_0_8/i1[9] ), .ZN(\SB2_0_8/Component_Function_1/NAND4_in[0] ) );
  BUF_X2 \SB2_0_12/BUF_0_0  ( .I(\SB2_0_12/buf_output[0] ), .Z(\RI5[0][144] )
         );
  INV_X1 U60 ( .I(n14), .ZN(n446) );
  BUF_X2 \SB1_1_29/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[13] ), .Z(
        \SB1_1_29/i0[6] ) );
  INV_X1 \SB1_1_14/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[103] ), .ZN(
        \SB1_1_14/i1_7 ) );
  INV_X1 \SB1_1_5/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[157] ), .ZN(
        \SB1_1_5/i1_7 ) );
  INV_X1 \SB1_1_31/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[1] ), .ZN(
        \SB1_1_31/i1_7 ) );
  BUF_X2 \SB1_1_1/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[180] ), .Z(
        \SB1_1_1/i0[9] ) );
  NAND3_X1 \SB1_1_18/Component_Function_4/N4  ( .A1(\SB1_1_18/i1[9] ), .A2(
        \SB1_1_18/i1_5 ), .A3(\SB1_1_18/i0_4 ), .ZN(
        \SB1_1_18/Component_Function_4/NAND4_in[3] ) );
  INV_X1 \SB1_1_9/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[132] ), .ZN(
        \SB1_1_9/i3[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_4/N4  ( .A1(\SB1_1_28/i1[9] ), .A2(
        \SB1_1_28/i1_5 ), .A3(\SB1_1_28/i0_4 ), .ZN(
        \SB1_1_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_14/Component_Function_4/N4  ( .A1(\SB1_1_14/i1[9] ), .A2(
        \SB1_1_14/i1_5 ), .A3(\SB1_1_14/i0_4 ), .ZN(
        \SB1_1_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_7/Component_Function_4/N4  ( .A1(\SB1_1_7/i1[9] ), .A2(
        \SB1_1_7/i1_5 ), .A3(\SB1_1_7/i0_4 ), .ZN(
        \SB1_1_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_18/Component_Function_0/N4  ( .A1(\SB1_1_18/i0[7] ), .A2(
        \SB1_1_18/i0_3 ), .A3(\SB1_1_18/i0_0 ), .ZN(
        \SB1_1_18/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_22/Component_Function_0/N1  ( .A1(\SB1_1_22/i0[10] ), .A2(
        \SB1_1_22/i0[9] ), .ZN(\SB1_1_22/Component_Function_0/NAND4_in[0] ) );
  INV_X1 \SB1_1_25/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[36] ), .ZN(
        \SB1_1_25/i3[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_4/N1  ( .A1(\SB1_1_18/i0[9] ), .A2(
        \SB1_1_18/i0_0 ), .A3(\SB1_1_18/i0[8] ), .ZN(
        \SB1_1_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_4/N4  ( .A1(\SB1_1_19/i1[9] ), .A2(
        \SB1_1_19/i1_5 ), .A3(\SB1_1_19/i0_4 ), .ZN(
        \SB1_1_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_25/Component_Function_2/N1  ( .A1(\SB1_1_25/i1_5 ), .A2(
        \SB1_1_25/i0[10] ), .A3(\SB1_1_25/i1[9] ), .ZN(
        \SB1_1_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_1/N2  ( .A1(\SB1_1_20/i0_3 ), .A2(
        \SB1_1_20/i1_7 ), .A3(\SB1_1_20/i0[8] ), .ZN(
        \SB1_1_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_26/Component_Function_1/N2  ( .A1(\SB1_1_26/i0_3 ), .A2(
        \SB1_1_26/i1_7 ), .A3(\SB1_1_26/i0[8] ), .ZN(
        \SB1_1_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_9/Component_Function_4/N2  ( .A1(\SB1_1_9/i3[0] ), .A2(
        \SB1_1_9/i0_0 ), .A3(\SB1_1_9/i1_7 ), .ZN(
        \SB1_1_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_1/Component_Function_1/N3  ( .A1(\SB1_1_1/i1_5 ), .A2(
        \SB1_1_1/i0[6] ), .A3(\SB1_1_1/i0[9] ), .ZN(
        \SB1_1_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_20/Component_Function_4/N4  ( .A1(\SB1_1_20/i1[9] ), .A2(
        \SB1_1_20/i1_5 ), .A3(\SB1_1_20/i0_4 ), .ZN(
        \SB1_1_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_28/Component_Function_2/N2  ( .A1(\SB1_1_28/i0_3 ), .A2(
        \SB1_1_28/i0[10] ), .A3(\SB1_1_28/i0[6] ), .ZN(
        \SB1_1_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_7/Component_Function_0/N3  ( .A1(\SB1_1_7/i0[10] ), .A2(
        \SB1_1_7/i0_4 ), .A3(\SB1_1_7/i0_3 ), .ZN(
        \SB1_1_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_4/Component_Function_3/N2  ( .A1(\SB1_1_4/i0_0 ), .A2(
        \SB1_1_4/i0_3 ), .A3(\SB1_1_4/i0_4 ), .ZN(
        \SB1_1_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_3/Component_Function_2/N2  ( .A1(\SB1_1_3/i0_3 ), .A2(
        \SB1_1_3/i0[10] ), .A3(\SB1_1_3/i0[6] ), .ZN(
        \SB1_1_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_4/Component_Function_0/N2  ( .A1(\SB1_1_4/i0[8] ), .A2(
        \SB1_1_4/i0[7] ), .A3(\SB1_1_4/i0[6] ), .ZN(
        \SB1_1_4/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_12/Component_Function_3/N3  ( .A1(\SB1_1_12/i1[9] ), .A2(
        \SB1_1_12/i1_7 ), .A3(\SB1_1_12/i0[10] ), .ZN(
        \SB1_1_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_26/Component_Function_3/N4  ( .A1(\SB1_1_26/i1_5 ), .A2(
        \SB1_1_26/i0[8] ), .A3(\SB1_1_26/i3[0] ), .ZN(
        \SB1_1_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_10/Component_Function_4/N4  ( .A1(\SB1_1_10/i1[9] ), .A2(
        \SB1_1_10/i1_5 ), .A3(\MC_ARK_ARC_1_0/buf_output[130] ), .ZN(
        \SB1_1_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_6/Component_Function_4/N1  ( .A1(\SB1_1_6/i0[9] ), .A2(
        \SB1_1_6/i0_0 ), .A3(\SB1_1_6/i0[8] ), .ZN(
        \SB1_1_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_3/N2  ( .A1(\SB1_1_0/i0_0 ), .A2(
        \SB1_1_0/i0_3 ), .A3(\SB1_1_0/i0_4 ), .ZN(
        \SB1_1_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_18/Component_Function_3/N2  ( .A1(\SB1_1_18/i0_0 ), .A2(
        \SB1_1_18/i0_3 ), .A3(\SB1_1_18/i0_4 ), .ZN(
        \SB1_1_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N3  ( .A1(\SB1_1_25/i0[9] ), .A2(
        \SB1_1_25/i0[10] ), .A3(\SB1_1_25/i0_3 ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_9/Component_Function_4/N1  ( .A1(\SB1_1_9/i0[9] ), .A2(
        \SB1_1_9/i0_0 ), .A3(\SB1_1_9/i0[8] ), .ZN(
        \SB1_1_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_16/Component_Function_3/N3  ( .A1(\SB1_1_16/i1[9] ), .A2(
        \SB1_1_16/i1_7 ), .A3(\SB1_1_16/i0[10] ), .ZN(
        \SB1_1_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_24/Component_Function_0/N2  ( .A1(\SB1_1_24/i0[8] ), .A2(
        \SB1_1_24/i0[7] ), .A3(\SB1_1_24/i0[6] ), .ZN(
        \SB1_1_24/Component_Function_0/NAND4_in[1] ) );
  INV_X1 \SB2_1_5/INV_1  ( .I(\SB1_1_9/buf_output[1] ), .ZN(\SB2_1_5/i1_7 ) );
  NAND3_X1 \SB2_1_11/Component_Function_1/N4  ( .A1(\SB2_1_11/i1_7 ), .A2(
        \SB2_1_11/i0[8] ), .A3(\SB2_1_11/i0_4 ), .ZN(
        \SB2_1_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_5/Component_Function_1/N4  ( .A1(\SB2_1_5/i1_7 ), .A2(
        \SB2_1_5/i0[8] ), .A3(\SB2_1_5/i0_4 ), .ZN(
        \SB2_1_5/Component_Function_1/NAND4_in[3] ) );
  BUF_X2 \SB2_1_14/BUF_0  ( .I(\SB1_1_19/buf_output[0] ), .Z(\SB2_1_14/i0[9] )
         );
  NAND3_X1 \SB2_1_18/Component_Function_1/N2  ( .A1(\SB2_1_18/i0_3 ), .A2(
        \SB2_1_18/i1_7 ), .A3(\SB2_1_18/i0[8] ), .ZN(
        \SB2_1_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_16/Component_Function_0/N2  ( .A1(\SB2_1_16/i0[8] ), .A2(
        \SB2_1_16/i0[7] ), .A3(\SB2_1_16/i0[6] ), .ZN(
        \SB2_1_16/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_28/Component_Function_4/N2  ( .A1(\SB2_1_28/i3[0] ), .A2(
        \SB2_1_28/i0_0 ), .A3(\SB2_1_28/i1_7 ), .ZN(
        \SB2_1_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_19/Component_Function_3/N4  ( .A1(\SB2_1_19/i1_5 ), .A2(
        \SB2_1_19/i0[8] ), .A3(\SB2_1_19/i3[0] ), .ZN(
        \SB2_1_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_23/Component_Function_1/N2  ( .A1(\SB2_1_23/i0_3 ), .A2(
        \SB2_1_23/i1_7 ), .A3(\SB2_1_23/i0[8] ), .ZN(
        \SB2_1_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_22/Component_Function_2/N1  ( .A1(\SB2_1_22/i1_5 ), .A2(
        \SB2_1_22/i0[10] ), .A3(\SB2_1_22/i1[9] ), .ZN(
        \SB2_1_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_1/N3  ( .A1(\SB2_1_26/i1_5 ), .A2(
        \SB2_1_26/i0[6] ), .A3(\SB2_1_26/i0[9] ), .ZN(
        \SB2_1_26/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_27/Component_Function_1/N1  ( .A1(\SB2_1_27/i0_3 ), .A2(
        \SB2_1_27/i1[9] ), .ZN(\SB2_1_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_0/N2  ( .A1(\SB2_1_27/i0[8] ), .A2(
        \SB2_1_27/i0[7] ), .A3(\SB2_1_27/i0[6] ), .ZN(
        \SB2_1_27/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_1/Component_Function_3/N1  ( .A1(\SB2_1_1/i1[9] ), .A2(
        \SB2_1_1/i0_3 ), .A3(\SB2_1_1/i0[6] ), .ZN(
        \SB2_1_1/Component_Function_3/NAND4_in[0] ) );
  INV_X1 \SB1_2_24/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[42] ), .ZN(
        \SB1_2_24/i3[0] ) );
  INV_X1 \SB1_2_31/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[0] ), .ZN(
        \SB1_2_31/i3[0] ) );
  BUF_X2 \SB1_2_12/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[114] ), .Z(
        \SB1_2_12/i0[9] ) );
  INV_X1 \SB1_2_4/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[162] ), .ZN(
        \SB1_2_4/i3[0] ) );
  INV_X1 \SB1_2_6/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[150] ), .ZN(
        \SB1_2_6/i3[0] ) );
  INV_X1 \SB1_2_28/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[19] ), .ZN(
        \SB1_2_28/i1_7 ) );
  BUF_X2 \SB1_2_20/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[66] ), .Z(
        \SB1_2_20/i0[9] ) );
  INV_X1 \SB1_2_2/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[175] ), .ZN(
        \SB1_2_2/i1_7 ) );
  BUF_X2 \SB1_2_23/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[48] ), .Z(
        \SB1_2_23/i0[9] ) );
  INV_X1 \SB1_2_31/INV_5  ( .I(\RI1[2][5] ), .ZN(\SB1_2_31/i1_5 ) );
  BUF_X2 \SB1_2_28/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[19] ), .Z(
        \SB1_2_28/i0[6] ) );
  NAND3_X1 \SB1_2_17/Component_Function_3/N3  ( .A1(\SB1_2_17/i1[9] ), .A2(
        \SB1_2_17/i1_7 ), .A3(\SB1_2_17/i0[10] ), .ZN(
        \SB1_2_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_4/Component_Function_4/N2  ( .A1(\SB1_2_4/i3[0] ), .A2(
        \SB1_2_4/i0_0 ), .A3(\SB1_2_4/i1_7 ), .ZN(
        \SB1_2_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_20/Component_Function_4/N2  ( .A1(\SB1_2_20/i3[0] ), .A2(
        \SB1_2_20/i0_0 ), .A3(\SB1_2_20/i1_7 ), .ZN(
        \SB1_2_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_12/Component_Function_3/N4  ( .A1(\SB1_2_12/i1_5 ), .A2(
        \SB1_2_12/i0[8] ), .A3(\SB1_2_12/i3[0] ), .ZN(
        \SB1_2_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_4/N1  ( .A1(\SB1_2_2/i0[9] ), .A2(
        \SB1_2_2/i0_0 ), .A3(\SB1_2_2/i0[8] ), .ZN(
        \SB1_2_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_16/Component_Function_4/N4  ( .A1(\SB1_2_16/i1[9] ), .A2(
        \SB1_2_16/i1_5 ), .A3(\SB1_2_16/i0_4 ), .ZN(
        \SB1_2_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_4/N4  ( .A1(\SB1_2_19/i1[9] ), .A2(
        \SB1_2_19/i1_5 ), .A3(\SB1_2_19/i0_4 ), .ZN(
        \SB1_2_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_4/N2  ( .A1(\SB1_2_19/i3[0] ), .A2(
        \SB1_2_19/i0_0 ), .A3(\SB1_2_19/i1_7 ), .ZN(
        \SB1_2_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_2/Component_Function_2/N1  ( .A1(\SB1_2_2/i1_5 ), .A2(
        \SB1_2_2/i0[10] ), .A3(\SB1_2_2/i1[9] ), .ZN(
        \SB1_2_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_5/N2  ( .A1(\SB1_2_31/i0_0 ), .A2(
        \SB1_2_31/i0[6] ), .A3(\SB1_2_31/i0[10] ), .ZN(
        \SB1_2_31/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_2/Component_Function_2/N2  ( .A1(\SB1_2_2/i0_3 ), .A2(
        \SB1_2_2/i0[10] ), .A3(\SB1_2_2/i0[6] ), .ZN(
        \SB1_2_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_19/Component_Function_4/N1  ( .A1(\SB1_2_19/i0[9] ), .A2(
        \SB1_2_19/i0_0 ), .A3(\SB1_2_19/i0[8] ), .ZN(
        \SB1_2_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_0/N2  ( .A1(\SB1_2_8/i0[8] ), .A2(
        \SB1_2_8/i0[7] ), .A3(\SB1_2_8/i0[6] ), .ZN(
        \SB1_2_8/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_31/Component_Function_1/N3  ( .A1(\SB1_2_31/i1_5 ), .A2(
        \SB1_2_31/i0[6] ), .A3(\SB1_2_31/i0[9] ), .ZN(
        \SB1_2_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_8/Component_Function_1/N3  ( .A1(\SB1_2_8/i1_5 ), .A2(
        \SB1_2_8/i0[6] ), .A3(\SB1_2_8/i0[9] ), .ZN(
        \SB1_2_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_6/Component_Function_1/N3  ( .A1(\SB1_2_6/i1_5 ), .A2(
        \SB1_2_6/i0[6] ), .A3(\SB1_2_6/i0[9] ), .ZN(
        \SB1_2_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_2/Component_Function_1/N3  ( .A1(\SB1_2_2/i1_5 ), .A2(
        \SB1_2_2/i0[6] ), .A3(\SB1_2_2/i0[9] ), .ZN(
        \SB1_2_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_15/Component_Function_2/N4  ( .A1(\SB1_2_15/i1_5 ), .A2(
        \SB1_2_15/i0_0 ), .A3(\SB1_2_15/i0_4 ), .ZN(
        \SB1_2_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_12/Component_Function_0/N4  ( .A1(\SB1_2_12/i0[7] ), .A2(
        \RI1[2][119] ), .A3(\RI1[2][116] ), .ZN(
        \SB1_2_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_31/Component_Function_4/N1  ( .A1(\SB1_2_31/i0[9] ), .A2(
        \SB1_2_31/i0_0 ), .A3(\SB1_2_31/i0[8] ), .ZN(
        \SB1_2_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_12/Component_Function_0/N3  ( .A1(\SB1_2_12/i0[10] ), .A2(
        \SB1_2_12/i0_4 ), .A3(\RI1[2][119] ), .ZN(
        \SB1_2_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_15/Component_Function_1/N3  ( .A1(\SB1_2_15/i1_5 ), .A2(
        \SB1_2_15/i0[6] ), .A3(\SB1_2_15/i0[9] ), .ZN(
        \SB1_2_15/Component_Function_1/NAND4_in[2] ) );
  BUF_X2 \SB2_2_10/BUF_0  ( .I(\SB1_2_15/buf_output[0] ), .Z(\SB2_2_10/i0[9] )
         );
  INV_X1 \SB2_2_19/INV_0  ( .I(\SB1_2_24/buf_output[0] ), .ZN(\SB2_2_19/i3[0] ) );
  BUF_X2 \SB2_2_27/BUF_1  ( .I(\SB1_2_31/buf_output[1] ), .Z(\SB2_2_27/i0[6] )
         );
  BUF_X2 \SB2_2_0/BUF_0  ( .I(\SB1_2_5/buf_output[0] ), .Z(\SB2_2_0/i0[9] ) );
  NAND3_X1 \SB2_2_26/Component_Function_4/N2  ( .A1(\SB2_2_26/i3[0] ), .A2(
        \SB2_2_26/i0_0 ), .A3(\SB2_2_26/i1_7 ), .ZN(
        \SB2_2_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_2/Component_Function_0/N4  ( .A1(\SB2_2_2/i0[7] ), .A2(
        \SB2_2_2/i0_3 ), .A3(\SB2_2_2/i0_0 ), .ZN(
        \SB2_2_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_24/Component_Function_1/N3  ( .A1(\SB2_2_24/i1_5 ), .A2(
        \SB2_2_24/i0[6] ), .A3(\SB2_2_24/i0[9] ), .ZN(
        \SB2_2_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_20/Component_Function_0/N4  ( .A1(\SB2_2_20/i0[7] ), .A2(
        \SB2_2_20/i0_3 ), .A3(\SB2_2_20/i0_0 ), .ZN(
        \SB2_2_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_19/Component_Function_3/N4  ( .A1(\SB2_2_19/i1_5 ), .A2(
        \SB2_2_19/i0[8] ), .A3(\SB2_2_19/i3[0] ), .ZN(
        \SB2_2_19/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_31/Component_Function_1/N1  ( .A1(\SB2_2_31/i0_3 ), .A2(
        \SB2_2_31/i1[9] ), .ZN(\SB2_2_31/Component_Function_1/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_124  ( .I(\SB2_2_12/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[124] ) );
  INV_X1 \SB1_3_6/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[150] ), .ZN(
        \SB1_3_6/i3[0] ) );
  INV_X1 \SB1_3_3/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[169] ), .ZN(
        \SB1_3_3/i1_7 ) );
  NAND3_X1 \SB1_3_5/Component_Function_4/N4  ( .A1(\SB1_3_5/i1[9] ), .A2(
        \SB1_3_5/i1_5 ), .A3(\SB1_3_5/i0_4 ), .ZN(
        \SB1_3_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_5/Component_Function_4/N1  ( .A1(\SB1_3_5/i0[9] ), .A2(
        \SB1_3_5/i0_0 ), .A3(\SB1_3_5/i0[8] ), .ZN(
        \SB1_3_5/Component_Function_4/NAND4_in[0] ) );
  BUF_X2 \SB1_3_18/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[79] ), .Z(
        \SB1_3_18/i0[6] ) );
  BUF_X2 \SB1_3_18/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[78] ), .Z(
        \SB1_3_18/i0[9] ) );
  INV_X1 \SB1_3_21/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[61] ), .ZN(
        \SB1_3_21/i1_7 ) );
  NAND3_X1 \SB1_3_22/Component_Function_4/N2  ( .A1(\SB1_3_22/i3[0] ), .A2(
        \SB1_3_22/i0_0 ), .A3(\SB1_3_22/i1_7 ), .ZN(
        \SB1_3_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_6/Component_Function_4/N2  ( .A1(\SB1_3_6/i3[0] ), .A2(
        \SB1_3_6/i0_0 ), .A3(\SB1_3_6/i1_7 ), .ZN(
        \SB1_3_6/Component_Function_4/NAND4_in[1] ) );
  INV_X1 \SB1_3_24/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[42] ), .ZN(
        \SB1_3_24/i3[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_0/N2  ( .A1(\SB1_3_25/i0[8] ), .A2(
        \SB1_3_25/i0[7] ), .A3(\SB1_3_25/i0[6] ), .ZN(
        \SB1_3_25/Component_Function_0/NAND4_in[1] ) );
  INV_X1 \SB1_3_18/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[78] ), .ZN(
        \SB1_3_18/i3[0] ) );
  INV_X1 \SB1_3_19/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[72] ), .ZN(
        \SB1_3_19/i3[0] ) );
  INV_X1 \SB1_3_25/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[37] ), .ZN(
        \SB1_3_25/i1_7 ) );
  NAND3_X1 \SB1_3_29/Component_Function_1/N2  ( .A1(\SB1_3_29/i0_3 ), .A2(
        \SB1_3_29/i1_7 ), .A3(\SB1_3_29/i0[8] ), .ZN(
        \SB1_3_29/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_27/Component_Function_3/N1  ( .A1(\SB1_3_27/i1[9] ), .A2(
        \SB1_3_27/i0_3 ), .A3(\SB1_3_27/i0[6] ), .ZN(
        \SB1_3_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_1/N4  ( .A1(\SB1_3_29/i1_7 ), .A2(
        \SB1_3_29/i0[8] ), .A3(\SB1_3_29/i0_4 ), .ZN(
        \SB1_3_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_9/Component_Function_4/N4  ( .A1(\SB1_3_9/i1[9] ), .A2(
        \SB1_3_9/i1_5 ), .A3(\SB1_3_9/i0_4 ), .ZN(
        \SB1_3_9/Component_Function_4/NAND4_in[3] ) );
  BUF_X2 \SB1_3_21/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[61] ), .Z(
        \SB1_3_21/i0[6] ) );
  NAND3_X1 \SB1_3_4/Component_Function_0/N3  ( .A1(\SB1_3_4/i0[10] ), .A2(
        \SB1_3_4/i0_4 ), .A3(\RI1[3][167] ), .ZN(
        \SB1_3_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_21/Component_Function_4/N4  ( .A1(\SB1_3_21/i1[9] ), .A2(
        \SB1_3_21/i1_5 ), .A3(\SB1_3_21/i0_4 ), .ZN(
        \SB1_3_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_12/Component_Function_4/N4  ( .A1(\SB1_3_12/i1[9] ), .A2(
        \SB1_3_12/i1_5 ), .A3(\SB1_3_12/i0_4 ), .ZN(
        \SB1_3_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_30/Component_Function_2/N4  ( .A1(\SB1_3_30/i1_5 ), .A2(
        \SB1_3_30/i0_0 ), .A3(\SB1_3_30/i0_4 ), .ZN(
        \SB1_3_30/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_22/Component_Function_0/N4  ( .A1(\SB1_3_22/i0[7] ), .A2(
        \SB1_3_22/i0_3 ), .A3(\SB1_3_22/i0_0 ), .ZN(
        \SB1_3_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_17/Component_Function_0/N2  ( .A1(\SB1_3_17/i0[8] ), .A2(
        \SB1_3_17/i0[7] ), .A3(\SB1_3_17/i0[6] ), .ZN(
        \SB1_3_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_18/Component_Function_4/N1  ( .A1(\SB1_3_18/i0[9] ), .A2(
        \SB1_3_18/i0_0 ), .A3(\SB1_3_18/i0[8] ), .ZN(
        \SB1_3_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_1/N3  ( .A1(\SB1_3_21/i1_5 ), .A2(
        \SB1_3_21/i0[6] ), .A3(\SB1_3_21/i0[9] ), .ZN(
        \SB1_3_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_19/Component_Function_2/N4  ( .A1(\SB1_3_19/i1_5 ), .A2(
        \SB1_3_19/i0_0 ), .A3(\SB1_3_19/i0_4 ), .ZN(
        \SB1_3_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_16/Component_Function_1/N3  ( .A1(\SB1_3_16/i1_5 ), .A2(
        \SB1_3_16/i0[6] ), .A3(\MC_ARK_ARC_1_2/buf_output[90] ), .ZN(
        \SB1_3_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_17/Component_Function_4/N1  ( .A1(\SB1_3_17/i0[9] ), .A2(
        \SB1_3_17/i0_0 ), .A3(\SB1_3_17/i0[8] ), .ZN(
        \SB1_3_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_8/Component_Function_3/N2  ( .A1(\SB1_3_8/i0_0 ), .A2(
        \SB1_3_8/i0_3 ), .A3(\SB1_3_8/i0_4 ), .ZN(
        \SB1_3_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_4/Component_Function_2/N2  ( .A1(\RI1[3][167] ), .A2(
        \SB1_3_4/i0[10] ), .A3(\SB1_3_4/i0[6] ), .ZN(
        \SB1_3_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_13/Component_Function_3/N1  ( .A1(\SB1_3_13/i1[9] ), .A2(
        \SB1_3_13/i0_3 ), .A3(\SB1_3_13/i0[6] ), .ZN(
        \SB1_3_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_3/N2  ( .A1(\SB1_3_14/i0_0 ), .A2(
        \RI1[3][107] ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_19/Component_Function_5/N4  ( .A1(\SB1_3_19/i0[9] ), .A2(
        \SB1_3_19/i0[6] ), .A3(\SB1_3_19/i0_4 ), .ZN(
        \SB1_3_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_24/Component_Function_2/N2  ( .A1(\SB1_3_24/i0_3 ), .A2(
        \SB1_3_24/i0[10] ), .A3(\SB1_3_24/i0[6] ), .ZN(
        \SB1_3_24/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_12/Component_Function_0/N1  ( .A1(\SB1_3_12/i0[10] ), .A2(
        \SB1_3_12/i0[9] ), .ZN(\SB1_3_12/Component_Function_0/NAND4_in[0] ) );
  INV_X1 \SB2_3_9/INV_1  ( .I(\SB1_3_13/buf_output[1] ), .ZN(\SB2_3_9/i1_7 )
         );
  INV_X1 \SB2_3_19/INV_0  ( .I(\SB1_3_24/buf_output[0] ), .ZN(\SB2_3_19/i3[0] ) );
  INV_X1 \SB2_3_7/INV_0  ( .I(\SB1_3_12/buf_output[0] ), .ZN(\SB2_3_7/i3[0] )
         );
  NAND3_X1 \SB2_3_25/Component_Function_4/N2  ( .A1(\SB2_3_25/i3[0] ), .A2(
        \SB2_3_25/i0_0 ), .A3(\SB2_3_25/i1_7 ), .ZN(
        \SB2_3_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_15/Component_Function_4/N2  ( .A1(\SB2_3_15/i3[0] ), .A2(
        \SB2_3_15/i0_0 ), .A3(\SB2_3_15/i1_7 ), .ZN(
        \SB2_3_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_25/Component_Function_4/N4  ( .A1(\SB2_3_25/i1[9] ), .A2(
        \SB2_3_25/i1_5 ), .A3(\SB1_3_26/buf_output[4] ), .ZN(
        \SB2_3_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_30/Component_Function_4/N4  ( .A1(\SB2_3_30/i1[9] ), .A2(
        \SB2_3_30/i1_5 ), .A3(\SB2_3_30/i0_4 ), .ZN(
        \SB2_3_30/Component_Function_4/NAND4_in[3] ) );
  INV_X1 \SB2_3_10/INV_4  ( .I(\SB2_3_10/i0_4 ), .ZN(\SB2_3_10/i0[7] ) );
  NAND3_X1 \SB2_3_19/Component_Function_0/N2  ( .A1(\SB2_3_19/i0[8] ), .A2(
        n2998), .A3(\SB2_3_19/i0[6] ), .ZN(
        \SB2_3_19/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_4/Component_Function_3/N3  ( .A1(\SB2_3_4/i1[9] ), .A2(
        \SB2_3_4/i1_7 ), .A3(\SB2_3_4/i0[10] ), .ZN(
        \SB2_3_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_31/Component_Function_1/N3  ( .A1(\SB2_3_31/i1_5 ), .A2(
        \SB2_3_31/i0[6] ), .A3(\SB2_3_31/i0[9] ), .ZN(
        \SB2_3_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_11/Component_Function_1/N3  ( .A1(\SB2_3_11/i1_5 ), .A2(
        \SB2_3_11/i0[6] ), .A3(\SB2_3_11/i0[9] ), .ZN(
        \SB2_3_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_2/Component_Function_0/N2  ( .A1(\SB2_3_2/i0[8] ), .A2(
        \SB2_3_2/i0[7] ), .A3(\SB2_3_2/i0[6] ), .ZN(
        \SB2_3_2/Component_Function_0/NAND4_in[1] ) );
  INV_X1 \SB1_4_26/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[30] ), .ZN(
        \SB1_4_26/i3[0] ) );
  INV_X1 \SB1_4_13/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[109] ), .ZN(
        \SB1_4_13/i1_7 ) );
  INV_X1 \SB1_4_15/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[101] ), .ZN(
        \SB1_4_15/i1_5 ) );
  BUF_X2 \SB1_4_30/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[6] ), .Z(
        \SB1_4_30/i0[9] ) );
  NAND3_X1 \SB1_4_21/Component_Function_4/N4  ( .A1(\SB1_4_21/i1[9] ), .A2(
        \SB1_4_21/i1_5 ), .A3(\SB1_4_21/i0_4 ), .ZN(
        \SB1_4_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_6/Component_Function_3/N2  ( .A1(\SB1_4_6/i0_0 ), .A2(
        \RI1[4][155] ), .A3(\SB1_4_6/i0_4 ), .ZN(
        \SB1_4_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_28/Component_Function_1/N4  ( .A1(\SB1_4_28/i1_7 ), .A2(
        \SB1_4_28/i0[8] ), .A3(\SB1_4_28/i0_4 ), .ZN(
        \SB1_4_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_26/Component_Function_4/N4  ( .A1(\SB1_4_26/i1[9] ), .A2(
        \SB1_4_26/i1_5 ), .A3(\SB1_4_26/i0_4 ), .ZN(
        \SB1_4_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_2/Component_Function_5/N3  ( .A1(\SB1_4_2/i1[9] ), .A2(
        \SB1_4_2/i0_4 ), .A3(\SB1_4_2/i0_3 ), .ZN(
        \SB1_4_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_21/Component_Function_2/N2  ( .A1(\SB1_4_21/i0_3 ), .A2(
        \SB1_4_21/i0[10] ), .A3(\SB1_4_21/i0[6] ), .ZN(
        \SB1_4_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_16/Component_Function_1/N2  ( .A1(\SB1_4_16/i0_3 ), .A2(
        \SB1_4_16/i1_7 ), .A3(\SB1_4_16/i0[8] ), .ZN(
        \SB1_4_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_12/Component_Function_0/N3  ( .A1(\SB1_4_12/i0[10] ), .A2(
        \SB1_4_12/i0_4 ), .A3(\RI1[4][119] ), .ZN(
        \SB1_4_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_21/Component_Function_1/N2  ( .A1(\SB1_4_21/i0_3 ), .A2(
        \SB1_4_21/i1_7 ), .A3(\SB1_4_21/i0[8] ), .ZN(
        \SB1_4_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_31/Component_Function_1/N1  ( .A1(\SB1_4_31/i0_3 ), .A2(
        \SB1_4_31/i1[9] ), .ZN(\SB1_4_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_26/Component_Function_0/N4  ( .A1(\SB1_4_26/i0[7] ), .A2(
        \SB1_4_26/i0_3 ), .A3(\SB1_4_26/i0_0 ), .ZN(
        \SB1_4_26/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_4_0/Component_Function_0/N1  ( .A1(\SB1_4_0/i0[10] ), .A2(
        \SB1_4_0/i0[9] ), .ZN(\SB1_4_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_10/Component_Function_4/N4  ( .A1(\SB1_4_10/i1[9] ), .A2(
        \SB1_4_10/i1_5 ), .A3(\SB1_4_10/i0_4 ), .ZN(
        \SB1_4_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_31/Component_Function_1/N4  ( .A1(\SB1_4_31/i1_7 ), .A2(
        \SB1_4_31/i0[8] ), .A3(\SB1_4_31/i0_4 ), .ZN(
        \SB1_4_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_24/Component_Function_2/N4  ( .A1(\SB1_4_24/i1_5 ), .A2(
        \SB1_4_24/i0_0 ), .A3(\SB1_4_24/i0_4 ), .ZN(
        \SB1_4_24/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_22/Component_Function_4/N1  ( .A1(\SB1_4_22/i0[9] ), .A2(
        \SB1_4_22/i0_0 ), .A3(\SB1_4_22/i0[8] ), .ZN(
        \SB1_4_22/Component_Function_4/NAND4_in[0] ) );
  INV_X1 \SB2_4_0/INV_0  ( .I(\SB1_4_5/buf_output[0] ), .ZN(\SB2_4_0/i3[0] )
         );
  NAND2_X1 \SB2_4_20/Component_Function_5/N1  ( .A1(\SB2_4_20/i0_0 ), .A2(
        \SB2_4_20/i3[0] ), .ZN(\SB2_4_20/Component_Function_5/NAND4_in[0] ) );
  INV_X1 \SB2_4_23/INV_1  ( .I(\SB1_4_27/buf_output[1] ), .ZN(\SB2_4_23/i1_7 )
         );
  INV_X1 \SB2_4_1/INV_1  ( .I(\SB1_4_5/buf_output[1] ), .ZN(\SB2_4_1/i1_7 ) );
  INV_X1 \SB2_4_17/INV_1  ( .I(\SB1_4_21/buf_output[1] ), .ZN(\SB2_4_17/i1_7 )
         );
  NAND3_X1 \SB2_4_21/Component_Function_4/N2  ( .A1(\SB2_4_21/i3[0] ), .A2(
        \SB2_4_21/i0_0 ), .A3(\SB2_4_21/i1_7 ), .ZN(
        \SB2_4_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_21/Component_Function_1/N4  ( .A1(\SB2_4_21/i1_7 ), .A2(
        \SB2_4_21/i0[8] ), .A3(\SB2_4_21/i0_4 ), .ZN(
        \SB2_4_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_7/Component_Function_1/N2  ( .A1(\SB2_4_7/i0_3 ), .A2(
        \SB2_4_7/i1_7 ), .A3(\SB2_4_7/i0[8] ), .ZN(
        \SB2_4_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_0/Component_Function_3/N4  ( .A1(n3978), .A2(\SB2_4_0/i0[8] ), .A3(\SB2_4_0/i3[0] ), .ZN(\SB2_4_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_18/Component_Function_3/N4  ( .A1(\SB2_4_18/i1_5 ), .A2(
        \SB2_4_18/i0[8] ), .A3(\SB2_4_18/i3[0] ), .ZN(
        \SB2_4_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_0/Component_Function_0/N2  ( .A1(\SB2_4_0/i0[8] ), .A2(
        \SB2_4_0/i0[7] ), .A3(\SB2_4_0/i0[6] ), .ZN(
        \SB2_4_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_27/Component_Function_1/N2  ( .A1(\SB2_4_27/i0_3 ), .A2(
        \SB2_4_27/i1_7 ), .A3(\SB2_4_27/i0[8] ), .ZN(
        \SB2_4_27/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_6/Component_Function_2/N1  ( .A1(\SB2_4_6/i1_5 ), .A2(
        \SB2_4_6/i0[10] ), .A3(\SB2_4_6/i1[9] ), .ZN(
        \SB2_4_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_17/Component_Function_1/N3  ( .A1(\SB2_4_17/i1_5 ), .A2(
        \SB2_4_17/i0[6] ), .A3(\SB2_4_17/i0[9] ), .ZN(
        \SB2_4_17/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_11/Component_Function_1/N1  ( .A1(\SB2_4_11/i0_3 ), .A2(
        \SB2_4_11/i1[9] ), .ZN(\SB2_4_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_6/Component_Function_3/N1  ( .A1(\SB2_4_6/i1[9] ), .A2(
        \SB2_4_6/i0_3 ), .A3(\SB2_4_6/i0[6] ), .ZN(
        \SB2_4_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_21/Component_Function_1/N2  ( .A1(\SB2_4_21/i0_3 ), .A2(
        \SB2_4_21/i1_7 ), .A3(\SB2_4_21/i0[8] ), .ZN(
        \SB2_4_21/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_23/Component_Function_2/N1  ( .A1(\SB2_4_23/i1_5 ), .A2(
        \SB2_4_23/i0[10] ), .A3(\SB2_4_23/i1[9] ), .ZN(
        \SB2_4_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_25/Component_Function_3/N2  ( .A1(\SB2_4_25/i0_0 ), .A2(
        \SB2_4_25/i0_3 ), .A3(\SB2_4_25/i0_4 ), .ZN(
        \SB2_4_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_21/Component_Function_0/N3  ( .A1(\SB2_4_21/i0[10] ), .A2(
        \SB2_4_21/i0_4 ), .A3(\SB2_4_21/i0_3 ), .ZN(
        \SB2_4_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_27/Component_Function_3/N3  ( .A1(\SB2_4_27/i1[9] ), .A2(
        \SB2_4_27/i1_7 ), .A3(\SB2_4_27/i0[10] ), .ZN(
        \SB2_4_27/Component_Function_3/NAND4_in[2] ) );
  INV_X1 \SB3_7/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[144] ), .ZN(
        \SB3_7/i3[0] ) );
  INV_X1 \SB3_26/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[30] ), .ZN(
        \SB3_26/i3[0] ) );
  BUF_X2 \SB3_21/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[60] ), .Z(
        \SB3_21/i0[9] ) );
  BUF_X2 \SB3_4/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[162] ), .Z(
        \SB3_4/i0[9] ) );
  BUF_X2 \SB3_22/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[54] ), .Z(
        \SB3_22/i0[9] ) );
  INV_X1 \SB3_10/INV_1  ( .I(\MC_ARK_ARC_1_4/buf_output[127] ), .ZN(
        \SB3_10/i1_7 ) );
  BUF_X2 \SB3_1/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[180] ), .Z(
        \SB3_1/i0[9] ) );
  NAND3_X1 \SB3_15/Component_Function_5/N3  ( .A1(\SB3_15/i1[9] ), .A2(
        \SB3_15/i0_4 ), .A3(\SB3_15/i0_3 ), .ZN(
        \SB3_15/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB3_27/Component_Function_2/N1  ( .A1(\SB3_27/i1_5 ), .A2(
        \SB3_27/i0[10] ), .A3(\SB3_27/i1[9] ), .ZN(
        \SB3_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_4/N4  ( .A1(\SB3_14/i1[9] ), .A2(
        \SB3_14/i1_5 ), .A3(\SB3_14/i0_4 ), .ZN(
        \SB3_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_31/Component_Function_0/N4  ( .A1(\SB3_31/i0[7] ), .A2(
        \SB3_31/i0_3 ), .A3(\SB3_31/i0_0 ), .ZN(
        \SB3_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_21/Component_Function_2/N3  ( .A1(\SB3_21/i0_3 ), .A2(
        \SB3_21/i0[8] ), .A3(\SB3_21/i0[9] ), .ZN(
        \SB3_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N4  ( .A1(\SB3_26/i1[9] ), .A2(
        \SB3_26/i1_5 ), .A3(\SB3_26/i0_4 ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_19/Component_Function_4/N3  ( .A1(\SB3_19/i0[9] ), .A2(
        \SB3_19/i0[10] ), .A3(\SB3_19/i0_3 ), .ZN(
        \SB3_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_5/Component_Function_2/N3  ( .A1(\SB3_5/i0_3 ), .A2(
        \SB3_5/i0[8] ), .A3(\SB3_5/i0[9] ), .ZN(
        \SB3_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_17/Component_Function_4/N1  ( .A1(\SB3_17/i0[9] ), .A2(
        \SB3_17/i0_0 ), .A3(\SB3_17/i0[8] ), .ZN(
        \SB3_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_2/N4  ( .A1(\SB3_14/i1_5 ), .A2(
        \SB3_14/i0_0 ), .A3(\SB3_14/i0_4 ), .ZN(
        \SB3_14/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB3_30/Component_Function_3/N2  ( .A1(\SB3_30/i0_0 ), .A2(
        \SB3_30/i0_3 ), .A3(\SB3_30/i0_4 ), .ZN(
        \SB3_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_30/Component_Function_1/N4  ( .A1(\SB3_30/i1_7 ), .A2(
        \SB3_30/i0[8] ), .A3(\SB3_30/i0_4 ), .ZN(
        \SB3_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_2/Component_Function_1/N4  ( .A1(\SB3_2/i1_7 ), .A2(
        \SB3_2/i0[8] ), .A3(\SB3_2/i0_4 ), .ZN(
        \SB3_2/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB3_14/Component_Function_1/N1  ( .A1(\SB3_14/i0_3 ), .A2(
        \SB3_14/i1[9] ), .ZN(\SB3_14/Component_Function_1/NAND4_in[0] ) );
  BUF_X2 \SB4_0/BUF_0  ( .I(\SB3_5/buf_output[0] ), .Z(\SB4_0/i0[9] ) );
  INV_X1 \SB4_8/INV_3  ( .I(\SB3_10/buf_output[3] ), .ZN(\SB4_8/i0[8] ) );
  INV_X1 \SB4_11/INV_0  ( .I(\SB3_16/buf_output[0] ), .ZN(\SB4_11/i3[0] ) );
  INV_X1 \SB4_18/INV_5  ( .I(\SB3_18/buf_output[5] ), .ZN(\SB4_18/i1_5 ) );
  NAND3_X1 \SB4_18/Component_Function_2/N4  ( .A1(\SB4_18/i1_5 ), .A2(
        \SB4_18/i0_0 ), .A3(\SB4_18/i0_4 ), .ZN(
        \SB4_18/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_26/Component_Function_4/N2  ( .A1(\SB4_26/i3[0] ), .A2(
        \SB3_29/buf_output[2] ), .A3(\SB4_26/i1_7 ), .ZN(
        \SB4_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_11/Component_Function_0/N2  ( .A1(\SB4_11/i0[8] ), .A2(
        \SB4_11/i0[7] ), .A3(\SB4_11/i0[6] ), .ZN(
        \SB4_11/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_20/Component_Function_3/N1  ( .A1(\SB4_20/i1[9] ), .A2(
        \SB4_20/i0_3 ), .A3(\SB4_20/i0[6] ), .ZN(
        \SB4_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U23 ( .A1(\SB4_7/i0[6] ), .A2(\SB4_7/i0[9] ), .A3(\SB4_7/i0_4 ), 
        .ZN(\SB4_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U31 ( .A1(\SB4_14/i0_4 ), .A2(n1495), .A3(\SB4_14/i1[9] ), .ZN(
        n2490) );
  NAND3_X1 U89 ( .A1(\SB4_7/i0[6] ), .A2(\SB4_7/i1_5 ), .A3(\SB4_7/i0[9] ), 
        .ZN(n2535) );
  BUF_X2 U571 ( .I(\SB3_26/buf_output[1] ), .Z(\SB4_22/i0[6] ) );
  NAND3_X1 U575 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i0[10] ), .A3(\SB3_31/i0_4 ), 
        .ZN(\SB3_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U578 ( .A1(\SB3_2/i0[6] ), .A2(\SB3_2/i0_4 ), .A3(
        \MC_ARK_ARC_1_4/buf_output[174] ), .ZN(n2390) );
  NAND3_X1 U582 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i1[9] ), .A3(\SB3_31/i0_4 ), 
        .ZN(\SB3_31/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U592 ( .A1(\SB3_26/i0[9] ), .A2(\SB3_26/i0_4 ), .A3(\SB3_26/i0[6] ), 
        .ZN(n2879) );
  NAND3_X1 U601 ( .A1(\SB3_18/i0[10] ), .A2(\SB3_18/i0_0 ), .A3(\SB3_18/i0[6] ), .ZN(\SB3_18/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U607 ( .A1(\SB3_10/i1_5 ), .A2(\SB3_10/i0_4 ), .A3(\SB3_10/i1[9] ), 
        .ZN(\SB3_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U663 ( .A1(\SB2_4_10/i0_3 ), .A2(\SB2_4_10/i1[9] ), .A3(
        \SB1_4_11/buf_output[4] ), .ZN(
        \SB2_4_10/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U679 ( .A1(\SB2_4_20/i1_7 ), .A2(\SB2_4_20/i0[8] ), .A3(
        \SB2_4_20/i0_4 ), .ZN(\SB2_4_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U683 ( .A1(\SB2_4_15/i0_3 ), .A2(\SB2_4_15/i0_4 ), .A3(
        \SB2_4_15/i1[9] ), .ZN(n2561) );
  NAND3_X1 U714 ( .A1(\SB1_4_4/i0[10] ), .A2(\SB1_4_4/i0_3 ), .A3(
        \SB1_4_4/i0[6] ), .ZN(n1428) );
  NAND3_X1 U715 ( .A1(\SB1_4_30/i0_0 ), .A2(\SB1_4_30/i1_5 ), .A3(
        \SB1_4_30/i0_4 ), .ZN(n1344) );
  NAND3_X1 U729 ( .A1(\RI1[4][155] ), .A2(\SB1_4_6/i0[7] ), .A3(\SB1_4_6/i0_0 ), .ZN(n2583) );
  NAND3_X1 U732 ( .A1(\SB1_4_18/i1[9] ), .A2(\SB1_4_18/i1_5 ), .A3(
        \SB1_4_18/i0_4 ), .ZN(\SB1_4_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U736 ( .A1(\RI1[4][131] ), .A2(\SB1_4_10/i0[7] ), .A3(
        \SB1_4_10/i0_0 ), .ZN(n1940) );
  NAND3_X1 U751 ( .A1(\SB1_4_14/i0[6] ), .A2(\SB1_4_14/i1[9] ), .A3(
        \SB1_4_14/i0_3 ), .ZN(\SB1_4_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U753 ( .A1(\SB1_4_15/i0_0 ), .A2(\SB1_4_15/i0_4 ), .A3(
        \SB1_4_15/i1_5 ), .ZN(n1545) );
  NAND3_X1 U764 ( .A1(\SB1_4_0/i0[10] ), .A2(\SB1_4_0/i1[9] ), .A3(
        \SB1_4_0/i1_7 ), .ZN(n2967) );
  NAND3_X1 U773 ( .A1(\SB1_4_9/i0_4 ), .A2(\SB1_4_9/i1_5 ), .A3(
        \SB1_4_9/i1[9] ), .ZN(n2717) );
  NAND3_X1 U799 ( .A1(\SB2_3_27/i0[6] ), .A2(\SB2_3_27/i1_5 ), .A3(
        \SB2_3_27/i0[9] ), .ZN(\SB2_3_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U802 ( .A1(\SB2_3_16/i0_0 ), .A2(\SB1_3_16/buf_output[5] ), .A3(
        \SB2_3_16/i0[7] ), .ZN(n2870) );
  NAND3_X1 U813 ( .A1(\SB2_3_22/i0_3 ), .A2(\SB2_3_22/i0_0 ), .A3(\RI3[3][58] ), .ZN(\SB2_3_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U815 ( .A1(\SB2_3_2/i0_0 ), .A2(\SB2_3_2/i1_5 ), .A3(
        \SB1_3_3/buf_output[4] ), .ZN(n1925) );
  INV_X1 U823 ( .I(\SB1_3_3/buf_output[1] ), .ZN(\SB2_3_31/i1_7 ) );
  NAND3_X1 U834 ( .A1(\SB2_3_4/i0[9] ), .A2(\SB2_3_4/i0_4 ), .A3(
        \SB2_3_4/i0[6] ), .ZN(n1866) );
  NAND3_X1 U840 ( .A1(\SB1_3_13/i0_0 ), .A2(\SB1_3_13/i0[9] ), .A3(
        \SB1_3_13/i0[8] ), .ZN(n1591) );
  NAND3_X1 U846 ( .A1(\SB1_3_20/i0_3 ), .A2(\SB1_3_20/i0[10] ), .A3(
        \SB1_3_20/i0[6] ), .ZN(\SB1_3_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U851 ( .A1(\MC_ARK_ARC_1_2/buf_output[121] ), .A2(
        \MC_ARK_ARC_1_2/buf_output[124] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[120] ), .ZN(
        \SB1_3_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U852 ( .A1(\SB1_3_18/i0[9] ), .A2(\SB1_3_18/i0_4 ), .A3(
        \SB1_3_18/i0[6] ), .ZN(n2045) );
  NAND3_X1 U856 ( .A1(\SB1_3_29/i0_3 ), .A2(\SB1_3_29/i0[7] ), .A3(
        \SB1_3_29/i0_0 ), .ZN(n2643) );
  NAND3_X1 U865 ( .A1(n5441), .A2(\SB1_3_31/i0_4 ), .A3(\SB1_3_31/i1_7 ), .ZN(
        \SB1_3_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U882 ( .A1(\SB1_3_11/i0[10] ), .A2(\SB1_3_11/i0[6] ), .A3(
        \SB1_3_11/i0_3 ), .ZN(\SB1_3_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U884 ( .A1(\SB1_3_6/i0[9] ), .A2(\SB1_3_6/i0[8] ), .A3(
        \SB1_3_6/i0_0 ), .ZN(n874) );
  INV_X1 U894 ( .I(\MC_ARK_ARC_1_2/buf_output[168] ), .ZN(\SB1_3_3/i3[0] ) );
  NAND3_X1 U895 ( .A1(\RI1[3][167] ), .A2(\SB1_3_4/i0[7] ), .A3(\SB1_3_4/i0_0 ), .ZN(\SB1_3_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U899 ( .A1(\SB1_3_3/i0[9] ), .A2(\SB1_3_3/i0[6] ), .A3(
        \SB1_3_3/i1_5 ), .ZN(n1868) );
  NAND3_X1 U900 ( .A1(\SB1_3_10/i0_0 ), .A2(\SB1_3_10/i3[0] ), .A3(
        \SB1_3_10/i1_7 ), .ZN(\SB1_3_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U904 ( .A1(\SB1_3_0/i1_5 ), .A2(\SB1_3_0/i0_4 ), .A3(
        \SB1_3_0/i1[9] ), .ZN(\SB1_3_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U914 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0[10] ), .A3(
        \SB2_2_12/i0_4 ), .ZN(n2476) );
  NAND3_X1 U921 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i0[9] ), .A3(
        \SB2_2_11/i0[6] ), .ZN(\SB2_2_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U923 ( .A1(\SB2_2_3/i0_4 ), .A2(\SB2_2_3/i1[9] ), .A3(n3994), .ZN(
        \SB2_2_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U930 ( .A1(\SB2_2_27/i0[7] ), .A2(\SB2_2_27/i0[8] ), .A3(
        \SB2_2_27/i0[6] ), .ZN(\SB2_2_27/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U933 ( .A1(\SB2_2_6/i0_4 ), .A2(\SB2_2_6/i1_7 ), .A3(
        \SB2_2_6/i0[8] ), .ZN(\SB2_2_6/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U949 ( .I(\SB2_2_23/i0_4 ), .ZN(\SB2_2_23/i0[7] ) );
  INV_X1 U970 ( .I(\SB1_2_20/buf_output[0] ), .ZN(\SB2_2_15/i3[0] ) );
  NAND3_X1 U975 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i0[10] ), .A3(
        \SB1_2_31/i0[9] ), .ZN(n2805) );
  NAND2_X1 U980 ( .A1(n2369), .A2(\SB1_2_19/Component_Function_4/NAND4_in[0] ), 
        .ZN(n2374) );
  NAND3_X1 U982 ( .A1(\SB1_2_30/i0[6] ), .A2(\SB1_2_30/i0[10] ), .A3(
        \SB1_2_30/i0_3 ), .ZN(n936) );
  NAND3_X1 U983 ( .A1(\MC_ARK_ARC_1_1/buf_output[55] ), .A2(n6938), .A3(
        \MC_ARK_ARC_1_1/buf_output[58] ), .ZN(
        \SB1_2_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U991 ( .A1(\MC_ARK_ARC_1_1/buf_output[42] ), .A2(\SB1_2_24/i0_3 ), 
        .A3(\SB1_2_24/i0[8] ), .ZN(n1353) );
  NAND3_X1 U996 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i1_7 ), .A3(
        \SB1_2_5/i0[8] ), .ZN(\SB1_2_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U998 ( .A1(\RI1[2][149] ), .A2(\SB1_2_7/i0[7] ), .A3(\SB1_2_7/i0_0 ), .ZN(n1700) );
  NAND3_X1 U999 ( .A1(\RI1[2][59] ), .A2(\SB1_2_22/i0[7] ), .A3(
        \SB1_2_22/i0_0 ), .ZN(n1636) );
  NAND3_X1 U1005 ( .A1(\SB1_2_19/i3[0] ), .A2(\SB1_2_19/i0[8] ), .A3(
        \SB1_2_19/i1_5 ), .ZN(n2086) );
  NAND3_X1 U1014 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i1[9] ), .A3(
        \SB1_2_31/i0[6] ), .ZN(\SB1_2_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1022 ( .A1(\RI1[2][59] ), .A2(\SB1_2_22/i0[6] ), .A3(
        \SB1_2_22/i0[10] ), .ZN(\SB1_2_22/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X1 U1033 ( .A1(\SB1_2_31/i0[10] ), .A2(\SB1_2_31/i1[9] ), .A3(
        \SB1_2_31/i1_7 ), .ZN(n3127) );
  NAND3_X1 U1035 ( .A1(\SB1_2_24/i0_0 ), .A2(\SB1_2_24/i0[7] ), .A3(
        \SB1_2_24/i0_3 ), .ZN(\SB1_2_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1037 ( .A1(\SB1_2_24/i0_0 ), .A2(\SB1_2_24/i3[0] ), .A3(
        \SB1_2_24/i1_7 ), .ZN(\SB1_2_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1058 ( .A1(\SB1_1_4/buf_output[4] ), .A2(\SB2_1_3/i1_7 ), .A3(
        \SB2_1_3/i0[8] ), .ZN(n1612) );
  NAND3_X1 U1065 ( .A1(\SB2_1_7/i0_0 ), .A2(\SB2_1_7/i0[9] ), .A3(
        \SB2_1_7/i0[8] ), .ZN(n1360) );
  NAND3_X1 U1072 ( .A1(\SB2_1_17/i0_4 ), .A2(\SB2_1_17/i1[9] ), .A3(n3990), 
        .ZN(\SB2_1_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1090 ( .A1(\SB2_1_3/i3[0] ), .A2(\SB2_1_3/i1_5 ), .A3(
        \SB2_1_3/i0[8] ), .ZN(n2999) );
  INV_X2 U1096 ( .I(\SB2_1_4/i1_7 ), .ZN(\SB1_1_8/buf_output[1] ) );
  NAND3_X1 U1102 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i0[8] ), .A3(
        \SB1_1_23/i1_7 ), .ZN(\SB1_1_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1109 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i0_3 ), .A3(
        \SB1_1_2/i0_4 ), .ZN(\SB1_1_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1123 ( .A1(\SB1_1_7/i0[10] ), .A2(\SB1_1_7/i1[9] ), .A3(
        \SB1_1_7/i1_7 ), .ZN(\SB1_1_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1126 ( .A1(\SB1_1_18/i0[9] ), .A2(\SB1_1_18/i0_3 ), .A3(
        \SB1_1_18/i0[8] ), .ZN(\SB1_1_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1131 ( .A1(\SB1_1_9/i0[9] ), .A2(\SB1_1_9/i1_5 ), .A3(
        \SB1_1_9/i0[6] ), .ZN(\SB1_1_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1141 ( .A1(\SB1_1_6/i0_4 ), .A2(\SB1_1_6/i0[8] ), .A3(
        \SB1_1_6/i1_7 ), .ZN(n1918) );
  NAND3_X1 U1142 ( .A1(\SB1_1_9/i3[0] ), .A2(\SB1_1_9/i0[8] ), .A3(
        \SB1_1_9/i1_5 ), .ZN(n2157) );
  NAND3_X1 U1143 ( .A1(\SB1_1_18/i0_0 ), .A2(\SB1_1_18/i1_5 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[82] ), .ZN(n887) );
  NAND3_X1 U1149 ( .A1(\SB1_1_3/i0[9] ), .A2(\SB1_1_3/i0_3 ), .A3(
        \SB1_1_3/i0[10] ), .ZN(\SB1_1_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1155 ( .A1(\SB1_1_9/i0_0 ), .A2(\SB1_1_9/i1_5 ), .A3(
        \SB1_1_9/i0_4 ), .ZN(n3116) );
  NAND3_X1 U1162 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i3[0] ), .A3(
        \SB1_1_2/i1_7 ), .ZN(\SB1_1_2/Component_Function_4/NAND4_in[1] ) );
  BUF_X2 U1174 ( .I(Key[76]), .Z(n200) );
  NAND3_X1 U1178 ( .A1(\SB2_0_10/i0[9] ), .A2(\SB2_0_10/i0_4 ), .A3(
        \SB2_0_10/i0[6] ), .ZN(\SB2_0_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1190 ( .A1(\SB1_0_18/buf_output[0] ), .A2(\SB2_0_13/i1_5 ), .A3(
        \SB2_0_13/i0[6] ), .ZN(\SB2_0_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1194 ( .A1(\SB2_0_12/i1[9] ), .A2(\SB2_0_12/i1_7 ), .A3(
        \SB2_0_12/i0[10] ), .ZN(\SB2_0_12/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U1199 ( .A1(\SB2_0_13/i1_5 ), .A2(\SB2_0_13/i3[0] ), .A3(
        \SB2_0_13/i0[8] ), .ZN(n1835) );
  NAND3_X1 U1210 ( .A1(\RI3[0][77] ), .A2(\RI3[0][75] ), .A3(\SB2_0_19/i0[9] ), 
        .ZN(n2254) );
  NAND3_X1 U1212 ( .A1(\SB2_0_8/i0[6] ), .A2(\RI3[0][142] ), .A3(
        \SB1_0_13/buf_output[0] ), .ZN(n2097) );
  INV_X1 U1213 ( .I(\RI3[0][115] ), .ZN(\SB2_0_12/i1_7 ) );
  NAND3_X1 U1218 ( .A1(\SB2_0_27/i0[10] ), .A2(\SB2_0_27/i0_3 ), .A3(
        \SB2_0_27/i0[6] ), .ZN(\SB2_0_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1222 ( .A1(\SB2_0_7/i0[9] ), .A2(\RI3[0][148] ), .A3(
        \SB2_0_7/i0[6] ), .ZN(n2743) );
  NAND3_X1 U1224 ( .A1(\SB2_0_3/i0[6] ), .A2(\SB2_0_3/i1_5 ), .A3(
        \SB2_0_3/i0[9] ), .ZN(n1663) );
  NAND4_X2 U1231 ( .A1(\SB1_0_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_13/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][128] ) );
  NAND3_X1 U1235 ( .A1(\SB1_0_31/i0_3 ), .A2(\SB1_0_31/i0_0 ), .A3(
        \SB1_0_31/i0[7] ), .ZN(n634) );
  NAND2_X1 U1237 ( .A1(\SB1_0_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_25/Component_Function_4/NAND4_in[1] ), .ZN(n2328) );
  NAND2_X1 U1240 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i1[9] ), .ZN(n1488) );
  NAND3_X1 U1242 ( .A1(\SB1_0_17/i0[10] ), .A2(\SB1_0_17/i0_3 ), .A3(
        \SB1_0_17/i0[9] ), .ZN(n1318) );
  NAND3_X1 U1249 ( .A1(\SB1_0_0/i0_4 ), .A2(\SB1_0_0/i1[9] ), .A3(
        \SB1_0_0/i1_5 ), .ZN(n2811) );
  NAND3_X1 U1250 ( .A1(\SB1_0_9/i0[6] ), .A2(\SB1_0_9/i1_5 ), .A3(
        \SB1_0_9/i0[9] ), .ZN(\SB1_0_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1252 ( .A1(\SB1_0_19/i0_4 ), .A2(\SB1_0_19/i1_7 ), .A3(
        \SB1_0_19/i0[8] ), .ZN(\SB1_0_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1253 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i0[8] ), .A3(
        \SB1_0_16/i1_7 ), .ZN(\SB1_0_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1261 ( .A1(\SB1_0_10/i0[9] ), .A2(\SB1_0_10/i1_5 ), .A3(
        \SB1_0_10/i0[6] ), .ZN(\SB1_0_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1262 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i0_0 ), .A3(
        \SB1_0_22/i0_4 ), .ZN(\SB1_0_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1263 ( .A1(\SB1_0_23/i0[6] ), .A2(\SB1_0_23/i0[9] ), .A3(
        \SB1_0_23/i1_5 ), .ZN(n1905) );
  NAND3_X1 U1269 ( .A1(\SB1_0_26/i0[10] ), .A2(\SB1_0_26/i0_3 ), .A3(n226), 
        .ZN(\SB1_0_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1270 ( .A1(\SB1_0_24/i0[6] ), .A2(\SB1_0_24/i0_3 ), .A3(
        \SB1_0_24/i1[9] ), .ZN(\SB1_0_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1272 ( .A1(\SB1_0_26/i0_0 ), .A2(\SB1_0_26/i1_5 ), .A3(
        \SB1_0_26/i0_4 ), .ZN(\SB1_0_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1275 ( .A1(\SB1_0_11/i0_0 ), .A2(\SB1_0_11/i0[9] ), .A3(
        \SB1_0_11/i0[8] ), .ZN(n2625) );
  BUF_X4 U1278 ( .I(\SB1_0_29/buf_output[5] ), .Z(\SB2_0_29/i0_3 ) );
  INV_X2 U1283 ( .I(\MC_ARK_ARC_1_2/buf_output[59] ), .ZN(\SB1_3_22/i1_5 ) );
  NAND3_X2 U1284 ( .A1(\SB2_1_17/i0_3 ), .A2(\SB2_1_17/i0[9] ), .A3(
        \SB2_1_17/i0[8] ), .ZN(n615) );
  BUF_X2 U1285 ( .I(n238), .Z(\SB1_0_14/i0[6] ) );
  NAND3_X2 U1286 ( .A1(\RI1[5][119] ), .A2(\SB3_12/i1[9] ), .A3(\SB3_12/i0_4 ), 
        .ZN(\SB3_12/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U1288 ( .I(n339), .ZN(\SB1_0_20/i0[8] ) );
  NAND3_X2 U1289 ( .A1(\SB1_2_20/i0[10] ), .A2(\SB1_2_20/i0_0 ), .A3(
        \SB1_2_20/i0[6] ), .ZN(\SB1_2_20/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X4 U1290 ( .I(\MC_ARK_ARC_1_4/buf_output[106] ), .Z(\SB3_14/i0_4 ) );
  CLKBUF_X4 U1291 ( .I(\SB3_10/buf_output[5] ), .Z(\SB4_10/i0_3 ) );
  BUF_X2 U1292 ( .I(\SB3_12/buf_output[2] ), .Z(\SB4_9/i0_0 ) );
  BUF_X4 U1298 ( .I(\RI1[3][17] ), .Z(\SB1_3_29/i0_3 ) );
  NAND3_X1 U1307 ( .A1(\SB4_22/i1_5 ), .A2(\SB4_22/i0[6] ), .A3(\SB4_22/i0[9] ), .ZN(\SB4_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1308 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i0[6] ), .A3(
        \SB3_26/buf_output[3] ), .ZN(n897) );
  BUF_X2 U1314 ( .I(\SB3_10/buf_output[3] ), .Z(\SB4_8/i0[10] ) );
  NAND3_X1 U1316 ( .A1(\SB3_8/i1[9] ), .A2(\SB3_8/i1_5 ), .A3(\SB3_8/i0_4 ), 
        .ZN(\SB3_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1323 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i1[9] ), .A3(
        \SB2_2_29/i0[6] ), .ZN(\SB2_2_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1330 ( .A1(\SB3_9/i1[9] ), .A2(\SB3_9/i0_3 ), .A3(\SB3_9/i0[6] ), 
        .ZN(\SB3_9/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U1332 ( .A1(\SB3_17/buf_output[3] ), .A2(\SB4_15/i0[9] ), .ZN(
        \SB4_15/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U1341 ( .A1(\SB1_4_28/i0_3 ), .A2(\SB1_4_28/i1[9] ), .ZN(
        \SB1_4_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1348 ( .A1(\SB1_4_9/i1_7 ), .A2(\SB1_4_9/i0[8] ), .A3(
        \SB1_4_9/i0_4 ), .ZN(\SB1_4_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1354 ( .A1(\SB3_17/buf_output[3] ), .A2(\SB4_15/i0_3 ), .A3(
        \SB4_15/i0_4 ), .ZN(\SB4_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1357 ( .A1(\SB4_31/i0[9] ), .A2(\SB4_31/i0[6] ), .A3(\SB4_31/i0_4 ), .ZN(\SB4_31/Component_Function_5/NAND4_in[3] ) );
  INV_X1 U1358 ( .I(\SB3_4/buf_output[2] ), .ZN(\SB4_1/i1[9] ) );
  BUF_X2 U1359 ( .I(\SB3_4/buf_output[2] ), .Z(\SB4_1/i0_0 ) );
  INV_X4 U1363 ( .I(\RI1[5][119] ), .ZN(\SB3_12/i1_5 ) );
  NAND3_X1 U1379 ( .A1(\SB4_9/i0_0 ), .A2(\SB4_9/i0[9] ), .A3(n1499), .ZN(
        n2941) );
  NAND3_X1 U1380 ( .A1(\SB1_0_23/i0[8] ), .A2(\SB1_0_23/i1_7 ), .A3(
        \SB1_0_23/i0_4 ), .ZN(n1904) );
  BUF_X4 U1381 ( .I(\SB2_4_20/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[76] ) );
  CLKBUF_X4 U1382 ( .I(\SB3_19/buf_output[5] ), .Z(\SB4_19/i0_3 ) );
  INV_X1 U1384 ( .I(\MC_ARK_ARC_1_4/buf_output[165] ), .ZN(\SB3_4/i0[8] ) );
  BUF_X2 U1385 ( .I(\MC_ARK_ARC_1_4/buf_output[165] ), .Z(\SB3_4/i0[10] ) );
  INV_X1 U1395 ( .I(\SB1_4_28/buf_output[1] ), .ZN(\SB2_4_24/i1_7 ) );
  NAND3_X1 U1398 ( .A1(\SB4_8/i0[10] ), .A2(\SB4_8/i0_3 ), .A3(\SB4_8/i0[6] ), 
        .ZN(n1642) );
  NAND3_X1 U1399 ( .A1(\SB4_8/i0[10] ), .A2(n3996), .A3(\SB4_8/i1_7 ), .ZN(
        n2195) );
  NAND2_X1 U1402 ( .A1(\SB4_26/i0_3 ), .A2(n573), .ZN(
        \SB4_26/Component_Function_1/NAND4_in[0] ) );
  INV_X1 U1412 ( .I(\MC_ARK_ARC_1_2/buf_output[129] ), .ZN(\SB1_3_10/i0[8] )
         );
  BUF_X2 U1413 ( .I(\MC_ARK_ARC_1_2/buf_output[129] ), .Z(\SB1_3_10/i0[10] )
         );
  NAND3_X1 U1420 ( .A1(\SB3_9/i0_3 ), .A2(\SB3_9/i0[8] ), .A3(\SB3_9/i0[9] ), 
        .ZN(\SB3_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1428 ( .A1(\SB4_18/i0_3 ), .A2(n1496), .A3(\SB4_18/i0[6] ), .ZN(
        \SB4_18/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U1433 ( .A1(\SB3_15/i0[10] ), .A2(\SB3_15/i0[9] ), .ZN(
        \SB3_15/Component_Function_0/NAND4_in[0] ) );
  CLKBUF_X4 U1436 ( .I(\SB1_4_8/buf_output[2] ), .Z(\SB2_4_5/i0_0 ) );
  BUF_X2 U1437 ( .I(\SB3_25/buf_output[2] ), .Z(\SB4_22/i0_0 ) );
  NAND3_X1 U1439 ( .A1(\SB4_29/i0_4 ), .A2(\SB4_29/i0_0 ), .A3(\SB4_29/i1_5 ), 
        .ZN(n852) );
  INV_X1 U1440 ( .I(\MC_ARK_ARC_1_4/buf_output[108] ), .ZN(\SB3_13/i3[0] ) );
  INV_X1 U1442 ( .I(\SB1_4_28/buf_output[3] ), .ZN(\SB2_4_26/i0[8] ) );
  BUF_X2 U1443 ( .I(\SB1_4_28/buf_output[3] ), .Z(\SB2_4_26/i0[10] ) );
  NAND3_X1 U1447 ( .A1(\SB4_3/i0[6] ), .A2(\SB4_3/i0[8] ), .A3(\SB4_3/i0[7] ), 
        .ZN(\SB4_3/Component_Function_0/NAND4_in[1] ) );
  BUF_X2 U1462 ( .I(\MC_ARK_ARC_1_1/buf_output[78] ), .Z(\SB1_2_18/i0[9] ) );
  INV_X1 U1463 ( .I(\MC_ARK_ARC_1_1/buf_output[78] ), .ZN(\SB1_2_18/i3[0] ) );
  NAND3_X1 U1464 ( .A1(\SB3_10/i0_0 ), .A2(\SB3_10/i0[6] ), .A3(
        \SB3_10/i0[10] ), .ZN(\SB3_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1467 ( .A1(\SB2_4_29/i1[9] ), .A2(\SB2_4_29/i1_5 ), .A3(
        \SB2_4_29/i0_4 ), .ZN(\SB2_4_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1470 ( .A1(\SB2_4_29/i0_3 ), .A2(\SB2_4_29/i0_4 ), .A3(
        \SB2_4_29/i1[9] ), .ZN(n2349) );
  NAND3_X1 U1475 ( .A1(\SB4_26/i0[9] ), .A2(\SB3_29/buf_output[2] ), .A3(n3989), .ZN(\SB4_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1476 ( .A1(\SB4_26/i0[9] ), .A2(\SB4_26/i0_3 ), .A3(n3989), .ZN(
        n967) );
  INV_X1 U1477 ( .I(\MC_ARK_ARC_1_4/buf_output[25] ), .ZN(\SB3_27/i1_7 ) );
  BUF_X2 U1484 ( .I(\SB3_30/buf_output[2] ), .Z(\SB4_27/i0_0 ) );
  NAND2_X1 U1485 ( .A1(\SB3_26/buf_output[3] ), .A2(\SB4_24/i0[9] ), .ZN(
        \SB4_24/Component_Function_0/NAND4_in[0] ) );
  BUF_X2 U1487 ( .I(\SB3_29/buf_output[0] ), .Z(\SB4_24/i0[9] ) );
  NAND3_X1 U1491 ( .A1(\SB4_30/i0[10] ), .A2(n3973), .A3(\SB4_30/i1_7 ), .ZN(
        \SB4_30/Component_Function_3/NAND4_in[2] ) );
  NAND2_X1 U1495 ( .A1(\SB4_10/i0_3 ), .A2(\SB4_10/i1[9] ), .ZN(
        \SB4_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1496 ( .A1(\SB4_10/i0_3 ), .A2(\SB4_10/i1[9] ), .A3(\SB4_10/i0_4 ), 
        .ZN(\SB4_10/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1519 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0[10] ), .A3(
        \SB1_0_21/i0[6] ), .ZN(\SB1_0_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1525 ( .A1(\SB1_2_12/i1_5 ), .A2(\SB1_2_12/i1[9] ), .A3(
        \SB1_2_12/i0_4 ), .ZN(\SB1_2_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1530 ( .A1(\SB1_1_29/i0_0 ), .A2(\SB1_1_29/i0[6] ), .A3(
        \SB1_1_29/i0[10] ), .ZN(\SB1_1_29/Component_Function_5/NAND4_in[1] )
         );
  INV_X1 U1555 ( .I(\MC_ARK_ARC_1_4/buf_output[81] ), .ZN(\SB3_18/i0[8] ) );
  BUF_X2 U1556 ( .I(\MC_ARK_ARC_1_4/buf_output[81] ), .Z(\SB3_18/i0[10] ) );
  NAND2_X1 U1558 ( .A1(\SB1_4_8/i3[0] ), .A2(\RI1[4][140] ), .ZN(n1615) );
  NAND3_X1 U1559 ( .A1(\SB4_27/i1_5 ), .A2(\SB4_27/i0[8] ), .A3(\SB4_27/i3[0] ), .ZN(\SB4_27/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U1560 ( .I(\MC_ARK_ARC_1_0/buf_output[31] ), .ZN(\SB1_1_26/i1_7 ) );
  BUF_X4 U1569 ( .I(\SB1_2_28/buf_output[4] ), .Z(\SB2_2_27/i0_4 ) );
  NAND3_X1 U1582 ( .A1(\SB3_14/i0[8] ), .A2(\SB3_14/i0_4 ), .A3(\SB3_14/i1_7 ), 
        .ZN(n2735) );
  CLKBUF_X4 U1584 ( .I(\MC_ARK_ARC_1_1/buf_output[22] ), .Z(\SB1_2_28/i0_4 )
         );
  NAND3_X1 U1588 ( .A1(\SB3_18/i1[9] ), .A2(\SB3_18/i0_4 ), .A3(\SB3_18/i0_3 ), 
        .ZN(\SB3_18/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U1590 ( .I(\MC_ARK_ARC_1_2/buf_output[10] ), .Z(\SB1_3_30/i0_4 )
         );
  BUF_X2 U1595 ( .I(\SB3_27/buf_output[4] ), .Z(\SB4_26/i0_4 ) );
  INV_X1 U1603 ( .I(\SB3_2/buf_output[1] ), .ZN(\SB4_30/i1_7 ) );
  BUF_X2 U1616 ( .I(\SB3_28/buf_output[2] ), .Z(\SB4_25/i0_0 ) );
  INV_X1 U1620 ( .I(\MC_ARK_ARC_1_3/buf_output[96] ), .ZN(\SB1_4_15/i3[0] ) );
  NAND3_X1 U1623 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i0[10] ), .A3(
        \SB4_17/i0[6] ), .ZN(\SB4_17/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 U1625 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i1[9] ), .ZN(
        \SB4_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1627 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i1[9] ), .A3(
        \SB1_1_23/i0_4 ), .ZN(\SB1_1_23/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U1630 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i1[9] ), .ZN(
        \SB1_1_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1638 ( .A1(\SB1_4_19/i0[8] ), .A2(\SB1_4_19/i0[7] ), .A3(
        \SB1_4_19/i0[6] ), .ZN(\SB1_4_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 U1642 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i3[0] ), .ZN(
        \SB4_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1658 ( .A1(\SB4_15/i1_5 ), .A2(n1497), .A3(\SB4_15/i3[0] ), .ZN(
        \SB4_15/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U1665 ( .I(\SB3_1/buf_output[1] ), .ZN(\SB4_29/i1_7 ) );
  NAND3_X1 U1671 ( .A1(\SB1_2_30/i0_0 ), .A2(\SB1_2_30/i0_3 ), .A3(
        \SB1_2_30/i0_4 ), .ZN(\SB1_2_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1675 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB2_3_7/i0[8] ), .A3(
        \SB2_3_7/i0[9] ), .ZN(\SB2_3_7/Component_Function_2/NAND4_in[2] ) );
  INV_X1 U1676 ( .I(\MC_ARK_ARC_1_3/buf_output[48] ), .ZN(\SB1_4_23/i3[0] ) );
  CLKBUF_X4 U1690 ( .I(\SB2_3_22/buf_output[2] ), .Z(\RI5[3][74] ) );
  NAND3_X1 U1694 ( .A1(\SB1_3_3/i0_3 ), .A2(\SB1_3_3/i0[8] ), .A3(
        \SB1_3_3/i0[9] ), .ZN(\SB1_3_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1701 ( .A1(\SB1_2_15/i1[9] ), .A2(\SB1_2_15/i1_7 ), .A3(
        \SB1_2_15/i0[10] ), .ZN(\SB1_2_15/Component_Function_3/NAND4_in[2] )
         );
  BUF_X2 U1719 ( .I(\SB3_12/buf_output[3] ), .Z(\SB4_10/i0[10] ) );
  BUF_X2 U1723 ( .I(\RI1[4][140] ), .Z(\SB1_4_8/i0_0 ) );
  NAND3_X1 U1731 ( .A1(\SB4_3/i0_3 ), .A2(\SB4_3/i0[10] ), .A3(\SB4_3/i0[9] ), 
        .ZN(n2417) );
  INV_X1 U1735 ( .I(\MC_ARK_ARC_1_0/buf_output[133] ), .ZN(\SB1_1_9/i1_7 ) );
  AND4_X2 U1744 ( .A1(\SB1_3_16/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_16/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_3_16/Component_Function_5/NAND4_in[0] ), .A4(n1547), .Z(n571) );
  AND4_X2 U1748 ( .A1(\SB3_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_29/Component_Function_2/NAND4_in[3] ), .Z(n573) );
  NAND3_X1 U1749 ( .A1(\SB1_4_18/i1[9] ), .A2(\SB1_4_18/i0_4 ), .A3(
        \SB1_4_18/i0_3 ), .ZN(\SB1_4_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1761 ( .A1(\SB1_4_20/i0_3 ), .A2(\SB1_4_20/i1_7 ), .A3(
        \SB1_4_20/i0[8] ), .ZN(\SB1_4_20/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U1763 ( .I(\SB1_1_11/buf_output[5] ), .Z(\SB2_1_11/i0_3 ) );
  NAND3_X1 U1765 ( .A1(\SB1_3_17/i0[7] ), .A2(\SB1_3_17/i0_3 ), .A3(
        \SB1_3_17/i0_0 ), .ZN(\SB1_3_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1766 ( .A1(\SB1_3_17/i0_3 ), .A2(\SB1_3_17/i0[8] ), .A3(
        \SB1_3_17/i0[9] ), .ZN(\SB1_3_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1767 ( .A1(\SB1_3_17/i0[6] ), .A2(\SB1_3_17/i1[9] ), .A3(
        \SB1_3_17/i0_3 ), .ZN(n1958) );
  BUF_X4 U1776 ( .I(\MC_ARK_ARC_1_1/buf_output[23] ), .Z(\SB1_2_28/i0_3 ) );
  CLKBUF_X4 U1777 ( .I(n254), .Z(\SB1_0_31/i0_0 ) );
  INV_X1 U1796 ( .I(\MC_ARK_ARC_1_1/buf_output[79] ), .ZN(\SB1_2_18/i1_7 ) );
  INV_X1 U1797 ( .I(\SB3_30/buf_output[1] ), .ZN(\SB4_26/i1_7 ) );
  BUF_X2 U1798 ( .I(\SB3_30/buf_output[1] ), .Z(\SB4_26/i0[6] ) );
  NAND3_X1 U1799 ( .A1(\SB1_3_12/i0[6] ), .A2(\SB1_3_12/i1_5 ), .A3(
        \SB1_3_12/i0[9] ), .ZN(n1670) );
  BUF_X4 U1806 ( .I(\RI1[3][5] ), .Z(\SB1_3_31/i0_3 ) );
  NAND3_X1 U1810 ( .A1(\SB1_0_29/i1_5 ), .A2(\SB1_0_29/i1[9] ), .A3(
        \SB1_0_29/i0_4 ), .ZN(n2320) );
  CLKBUF_X4 U1819 ( .I(\MC_ARK_ARC_1_4/buf_output[86] ), .Z(\SB3_17/i0_0 ) );
  INV_X1 U1825 ( .I(n238), .ZN(\SB1_0_14/i1_7 ) );
  NAND3_X2 U1826 ( .A1(\SB2_0_21/i1[9] ), .A2(\SB2_0_21/i1_5 ), .A3(
        \SB2_0_21/i0_4 ), .ZN(\SB2_0_21/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U1830 ( .I(\MC_ARK_ARC_1_4/buf_output[115] ), .ZN(\SB3_12/i1_7 ) );
  INV_X1 U1831 ( .I(\MC_ARK_ARC_1_2/buf_output[60] ), .ZN(\SB1_3_21/i3[0] ) );
  NAND3_X1 U1833 ( .A1(\RI1[1][47] ), .A2(\SB1_1_24/i0[10] ), .A3(
        \SB1_1_24/i0[6] ), .ZN(\SB1_1_24/Component_Function_2/NAND4_in[1] ) );
  INV_X1 U1843 ( .I(n243), .ZN(\SB1_0_9/i1_7 ) );
  INV_X1 U1853 ( .I(\SB3_22/buf_output[5] ), .ZN(\SB4_22/i1_5 ) );
  INV_X1 U1856 ( .I(n295), .ZN(\SB1_0_10/i3[0] ) );
  NAND3_X1 U1873 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i0[7] ), .A3(
        \SB1_2_10/i0_3 ), .ZN(n1376) );
  NAND3_X1 U1874 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i1_5 ), .A3(
        \SB1_2_10/i0_4 ), .ZN(n2296) );
  INV_X1 U1878 ( .I(\MC_ARK_ARC_1_4/buf_output[103] ), .ZN(\SB3_14/i1_7 ) );
  NAND3_X1 U1883 ( .A1(n6290), .A2(\SB1_0_18/i0[7] ), .A3(\SB1_0_18/i0_3 ), 
        .ZN(\SB1_0_18/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U1890 ( .A1(\SB4_25/i0_3 ), .A2(\SB4_25/i1[9] ), .ZN(n946) );
  NAND3_X1 U1891 ( .A1(\SB4_25/i1[9] ), .A2(\SB4_25/i0_4 ), .A3(\SB4_25/i0_3 ), 
        .ZN(\SB4_25/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1892 ( .A1(\SB4_25/i0_3 ), .A2(\SB4_25/i0[6] ), .A3(\SB4_25/i1[9] ), .ZN(n2042) );
  BUF_X4 U1904 ( .I(\MC_ARK_ARC_1_2/buf_output[59] ), .Z(\SB1_3_22/i0_3 ) );
  OR3_X2 U1910 ( .A1(\MC_ARK_ARC_1_1/buf_output[171] ), .A2(
        \MC_ARK_ARC_1_1/buf_output[173] ), .A3(
        \MC_ARK_ARC_1_1/buf_output[168] ), .Z(
        \SB1_2_3/Component_Function_3/NAND4_in[3] ) );
  OR3_X2 U1914 ( .A1(\SB1_0_24/buf_output[3] ), .A2(\SB1_0_22/buf_output[5] ), 
        .A3(\SB1_0_27/buf_output[0] ), .Z(
        \SB2_0_22/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X4 U1915 ( .I(\MC_ARK_ARC_1_1/buf_output[74] ), .Z(\SB1_2_19/i0_0 )
         );
  OR3_X2 U1917 ( .A1(\MC_ARK_ARC_1_0/buf_output[63] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[60] ), .A3(\MC_ARK_ARC_1_0/buf_output[65] ), 
        .Z(\SB1_1_21/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U1918 ( .I(\MC_ARK_ARC_1_0/buf_output[65] ), .ZN(\SB1_1_21/i1_5 ) );
  CLKBUF_X4 U1921 ( .I(\MC_ARK_ARC_1_0/buf_output[176] ), .Z(\SB1_1_2/i0_0 )
         );
  INV_X1 U1924 ( .I(n386), .ZN(\SB1_0_26/i1_5 ) );
  CLKBUF_X4 U1939 ( .I(\RI3[5][149] ), .Z(\SB4_7/i0_3 ) );
  BUF_X2 U1954 ( .I(\MC_ARK_ARC_1_4/buf_output[67] ), .Z(\SB3_20/i0[6] ) );
  BUF_X4 U1955 ( .I(\SB2_4_18/buf_output[2] ), .Z(\RI5[4][98] ) );
  BUF_X4 U1959 ( .I(\SB2_4_8/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[148] ) );
  BUF_X4 U1961 ( .I(\SB2_4_16/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[120] ) );
  CLKBUF_X4 U1962 ( .I(\SB2_4_23/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[73] ) );
  BUF_X4 U1963 ( .I(\SB2_4_12/buf_output[4] ), .Z(\RI5[4][124] ) );
  BUF_X4 U1966 ( .I(\SB2_4_13/buf_output[5] ), .Z(\RI5[4][113] ) );
  BUF_X4 U1967 ( .I(\SB2_4_1/buf_output[5] ), .Z(\RI5[4][185] ) );
  BUF_X4 U1969 ( .I(\SB2_4_4/buf_output[0] ), .Z(\RI5[4][0] ) );
  BUF_X4 U1970 ( .I(\SB2_4_0/buf_output[1] ), .Z(\RI5[4][19] ) );
  CLKBUF_X4 U1975 ( .I(\SB1_4_14/buf_output[3] ), .Z(\SB2_4_12/i0[10] ) );
  CLKBUF_X4 U1984 ( .I(\MC_ARK_ARC_1_3/buf_output[44] ), .Z(\SB1_4_24/i0_0 )
         );
  CLKBUF_X4 U1985 ( .I(\MC_ARK_ARC_1_3/buf_output[151] ), .Z(\SB1_4_6/i0[6] )
         );
  BUF_X4 U1993 ( .I(\SB2_3_3/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[178] ) );
  CLKBUF_X4 U1995 ( .I(\SB2_3_23/buf_output[0] ), .Z(\RI5[3][78] ) );
  BUF_X4 U1996 ( .I(\SB2_3_26/buf_output[3] ), .Z(\RI5[3][45] ) );
  NAND2_X1 U2000 ( .A1(n2674), .A2(\SB1_3_22/Component_Function_4/NAND4_in[1] ), .ZN(n1775) );
  BUF_X4 U2011 ( .I(\SB2_2_5/buf_output[0] ), .Z(\RI5[2][186] ) );
  BUF_X4 U2014 ( .I(\SB2_2_1/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[3] ) );
  BUF_X4 U2017 ( .I(\SB2_2_26/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[40] ) );
  BUF_X2 U2028 ( .I(\MC_ARK_ARC_1_1/buf_output[102] ), .Z(\SB1_2_14/i0[9] ) );
  BUF_X4 U2033 ( .I(\SB2_1_19/buf_output[4] ), .Z(\RI5[1][82] ) );
  BUF_X4 U2035 ( .I(\SB2_1_13/buf_output[3] ), .Z(\RI5[1][123] ) );
  BUF_X4 U2036 ( .I(\SB2_1_15/buf_output[1] ), .Z(\RI5[1][121] ) );
  BUF_X4 U2039 ( .I(\SB2_1_28/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[48] ) );
  NAND3_X2 U2042 ( .A1(\SB2_1_4/i0_0 ), .A2(\SB2_1_4/i1_5 ), .A3(
        \SB2_1_4/i0_4 ), .ZN(n2251) );
  CLKBUF_X4 U2050 ( .I(\MC_ARK_ARC_1_0/buf_output[128] ), .Z(\SB1_1_10/i0_0 )
         );
  BUF_X4 U2057 ( .I(\SB2_0_31/buf_output[1] ), .Z(\RI5[0][25] ) );
  BUF_X4 U2058 ( .I(\SB2_0_30/buf_output[3] ), .Z(\RI5[0][21] ) );
  NAND2_X1 U2063 ( .A1(\SB1_0_27/Component_Function_4/NAND4_in[1] ), .A2(n1469), .ZN(n1468) );
  BUF_X2 U2070 ( .I(n259), .Z(\SB1_0_28/i0[9] ) );
  BUF_X2 U2071 ( .I(n255), .Z(\SB1_0_30/i0[9] ) );
  BUF_X2 U2072 ( .I(n289), .Z(\SB1_0_13/i0[9] ) );
  CLKBUF_X1 U2075 ( .I(n318), .Z(n1105) );
  NAND3_X1 U2078 ( .A1(\SB1_0_30/i0_0 ), .A2(\SB1_0_30/i3[0] ), .A3(
        \SB1_0_30/i1_7 ), .ZN(n2547) );
  INV_X2 U2079 ( .I(\SB1_0_13/i0_4 ), .ZN(\SB1_0_13/i0[7] ) );
  CLKBUF_X4 U2084 ( .I(n300), .Z(\SB1_0_8/i0_0 ) );
  BUF_X2 U2085 ( .I(n228), .Z(\SB1_0_24/i0[6] ) );
  NAND3_X1 U2089 ( .A1(\SB1_0_9/i0[9] ), .A2(\SB1_0_9/i0[10] ), .A3(
        \SB1_0_9/i0_3 ), .ZN(\SB1_0_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2090 ( .A1(\SB1_0_1/i0[9] ), .A2(\SB1_0_1/i0[10] ), .A3(
        \SB1_0_1/i0_3 ), .ZN(\SB1_0_1/Component_Function_4/NAND4_in[2] ) );
  CLKBUF_X4 U2092 ( .I(n347), .Z(\SB1_0_16/i0[10] ) );
  NAND3_X1 U2093 ( .A1(\SB1_0_8/i0_4 ), .A2(\SB1_0_8/i1[9] ), .A3(
        \SB1_0_8/i1_5 ), .ZN(\SB1_0_8/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U2094 ( .A1(\SB1_0_9/i0[10] ), .A2(\SB1_0_9/i0[9] ), .ZN(
        \SB1_0_9/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U2099 ( .A1(\SB1_0_14/i0[10] ), .A2(\SB1_0_14/i0[9] ), .ZN(n2922)
         );
  INV_X1 U2100 ( .I(n405), .ZN(\SB1_0_7/i1_5 ) );
  NAND3_X1 U2101 ( .A1(\SB1_0_3/i3[0] ), .A2(\SB1_0_3/i0_0 ), .A3(
        \SB1_0_3/i1_7 ), .ZN(\SB1_0_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2102 ( .A1(\SB1_0_19/i0_4 ), .A2(\SB1_0_19/i1_5 ), .A3(
        \SB1_0_19/i1[9] ), .ZN(n1054) );
  NAND3_X1 U2106 ( .A1(\SB1_0_24/i1_5 ), .A2(\SB1_0_24/i0[6] ), .A3(n267), 
        .ZN(\SB1_0_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2108 ( .A1(\SB1_0_25/i1_5 ), .A2(\SB1_0_25/i0[8] ), .A3(
        \SB1_0_25/i3[0] ), .ZN(\SB1_0_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2109 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0[8] ), .A3(
        \SB1_0_15/i1_7 ), .ZN(\SB1_0_15/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2110 ( .A1(\SB1_0_0/i0[9] ), .A2(\SB1_0_0/i0_0 ), .A3(
        \SB1_0_0/i0[8] ), .ZN(\SB1_0_0/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 U2111 ( .A1(\SB1_0_18/i0[10] ), .A2(\SB1_0_18/i0[9] ), .ZN(
        \SB1_0_18/Component_Function_0/NAND4_in[0] ) );
  BUF_X2 U2112 ( .I(\SB1_0_22/buf_output[0] ), .Z(\SB2_0_17/i0[9] ) );
  INV_X1 U2114 ( .I(\RI3[0][60] ), .ZN(\SB2_0_21/i3[0] ) );
  BUF_X2 U2116 ( .I(\RI3[0][121] ), .Z(\SB2_0_11/i0[6] ) );
  NAND3_X1 U2124 ( .A1(\SB2_0_10/i0[9] ), .A2(\SB2_0_10/i0[6] ), .A3(
        \SB2_0_10/i1_5 ), .ZN(\SB2_0_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2132 ( .A1(\RI3[0][49] ), .A2(\SB2_0_23/i0[9] ), .A3(\RI3[0][52] ), 
        .ZN(\SB2_0_23/Component_Function_5/NAND4_in[3] ) );
  CLKBUF_X4 U2133 ( .I(\RI3[0][111] ), .Z(\SB2_0_13/i0[10] ) );
  NAND3_X1 U2134 ( .A1(\RI3[0][77] ), .A2(\RI3[0][75] ), .A3(\RI3[0][76] ), 
        .ZN(n2736) );
  CLKBUF_X1 U2139 ( .I(n128), .Z(\MC_ARK_ARC_1_0/buf_keyinput[71] ) );
  INV_X1 U2149 ( .I(\MC_ARK_ARC_1_0/buf_output[126] ), .ZN(\SB1_1_10/i3[0] )
         );
  INV_X1 U2150 ( .I(\MC_ARK_ARC_1_0/buf_output[60] ), .ZN(\SB1_1_21/i3[0] ) );
  BUF_X2 U2152 ( .I(\MC_ARK_ARC_1_0/buf_output[73] ), .Z(\SB1_1_19/i0[6] ) );
  CLKBUF_X4 U2156 ( .I(\MC_ARK_ARC_1_0/buf_output[129] ), .Z(\SB1_1_10/i0[10] ) );
  NAND3_X1 U2158 ( .A1(\SB1_1_6/i1[9] ), .A2(\SB1_1_6/i1_5 ), .A3(
        \SB1_1_6/i0_4 ), .ZN(\SB1_1_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2161 ( .A1(\SB1_1_28/i0_3 ), .A2(\SB1_1_28/i1_7 ), .A3(
        \SB1_1_28/i0[8] ), .ZN(\SB1_1_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2166 ( .A1(\SB1_1_4/i0[10] ), .A2(\SB1_1_4/i0_4 ), .A3(
        \SB1_1_4/i0_3 ), .ZN(\SB1_1_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2167 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i0[10] ), .A3(
        \SB1_1_19/i0[6] ), .ZN(\SB1_1_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2171 ( .A1(\SB1_1_1/i1_7 ), .A2(\SB1_1_1/i0[8] ), .A3(
        \SB1_1_1/i0_4 ), .ZN(\SB1_1_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2180 ( .A1(\SB1_1_4/i0[9] ), .A2(\SB1_1_4/i0[10] ), .A3(
        \SB1_1_4/i0_3 ), .ZN(\SB1_1_4/Component_Function_4/NAND4_in[2] ) );
  BUF_X2 U2190 ( .I(\SB1_1_27/buf_output[0] ), .Z(\SB2_1_22/i0[9] ) );
  NAND3_X1 U2192 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i1_7 ), .A3(
        \SB2_1_5/i0[8] ), .ZN(\SB2_1_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2200 ( .A1(\SB2_1_22/i1_7 ), .A2(n6283), .A3(\SB2_1_22/i0_4 ), 
        .ZN(\SB2_1_22/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U2214 ( .I(\MC_ARK_ARC_1_1/buf_output[187] ), .ZN(\SB1_2_0/i1_7 ) );
  INV_X1 U2215 ( .I(\MC_ARK_ARC_1_1/buf_output[139] ), .ZN(\SB1_2_8/i1_7 ) );
  INV_X1 U2217 ( .I(\MC_ARK_ARC_1_1/buf_output[36] ), .ZN(\SB1_2_25/i3[0] ) );
  CLKBUF_X4 U2218 ( .I(\MC_ARK_ARC_1_1/buf_output[16] ), .Z(\SB1_2_29/i0_4 )
         );
  INV_X1 U2221 ( .I(\MC_ARK_ARC_1_1/buf_output[72] ), .ZN(\SB1_2_19/i3[0] ) );
  NAND3_X1 U2222 ( .A1(\SB1_2_6/i0_3 ), .A2(\SB1_2_6/i0[10] ), .A3(
        \SB1_2_6/i0[6] ), .ZN(\SB1_2_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2224 ( .A1(\SB1_2_23/i0[9] ), .A2(\SB1_2_23/i0[6] ), .A3(
        \SB1_2_23/i0_4 ), .ZN(\SB1_2_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2226 ( .A1(\SB1_2_8/i1[9] ), .A2(\SB1_2_8/i0_3 ), .A3(
        \SB1_2_8/i0[6] ), .ZN(\SB1_2_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2228 ( .A1(\SB1_2_0/i1[9] ), .A2(\SB1_2_0/i1_7 ), .A3(
        \SB1_2_0/i0[10] ), .ZN(\SB1_2_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2232 ( .A1(\SB1_2_18/i1_5 ), .A2(\SB1_2_18/i0[6] ), .A3(
        \SB1_2_18/i0[9] ), .ZN(\SB1_2_18/Component_Function_1/NAND4_in[2] ) );
  INV_X1 U2235 ( .I(\MC_ARK_ARC_1_1/buf_output[49] ), .ZN(\SB1_2_23/i1_7 ) );
  NAND3_X1 U2237 ( .A1(\SB1_2_8/i1[9] ), .A2(\SB1_2_8/i1_5 ), .A3(
        \SB1_2_8/i0_4 ), .ZN(\SB1_2_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2242 ( .A1(\SB1_2_21/i1_5 ), .A2(\SB1_2_21/i0_0 ), .A3(
        \SB1_2_21/i0_4 ), .ZN(\SB1_2_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2245 ( .A1(\RI1[2][149] ), .A2(\SB1_2_7/i0_0 ), .A3(\SB1_2_7/i0_4 ), .ZN(\SB1_2_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2248 ( .A1(\RI1[2][119] ), .A2(\SB1_2_12/i0[8] ), .A3(
        \MC_ARK_ARC_1_1/buf_output[114] ), .ZN(
        \SB1_2_12/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 U2253 ( .I(\SB1_2_31/buf_output[4] ), .Z(\SB2_2_30/i0_4 ) );
  NAND3_X1 U2270 ( .A1(\SB2_2_15/i0[10] ), .A2(\SB2_2_15/i0_4 ), .A3(
        \SB2_2_15/i0_3 ), .ZN(\SB2_2_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2277 ( .A1(\SB2_2_27/i0[7] ), .A2(\SB2_2_27/i0_3 ), .A3(
        \SB2_2_27/i0_0 ), .ZN(\SB2_2_27/Component_Function_0/NAND4_in[3] ) );
  INV_X1 U2279 ( .I(n125), .ZN(n433) );
  CLKBUF_X4 U2285 ( .I(\MC_ARK_ARC_1_2/buf_output[8] ), .Z(\SB1_3_30/i0_0 ) );
  NAND3_X1 U2292 ( .A1(\SB1_3_8/i1[9] ), .A2(\SB1_3_8/i0_3 ), .A3(
        \SB1_3_8/i0[6] ), .ZN(\SB1_3_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2293 ( .A1(\SB1_3_21/i3[0] ), .A2(\SB1_3_21/i0_0 ), .A3(
        \SB1_3_21/i1_7 ), .ZN(\SB1_3_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2297 ( .A1(\SB1_3_13/i0_3 ), .A2(\SB1_3_13/i1_7 ), .A3(
        \SB1_3_13/i0[8] ), .ZN(\SB1_3_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2301 ( .A1(\SB1_3_24/i0[10] ), .A2(\SB1_3_24/i0_3 ), .A3(
        \SB1_3_24/i0[9] ), .ZN(n2024) );
  CLKBUF_X4 U2304 ( .I(\MC_ARK_ARC_1_2/buf_output[102] ), .Z(\SB1_3_14/i0[9] )
         );
  CLKBUF_X4 U2305 ( .I(\MC_ARK_ARC_1_2/buf_output[111] ), .Z(\SB1_3_13/i0[10] ) );
  NAND3_X1 U2307 ( .A1(\SB1_3_8/i0[7] ), .A2(\SB1_3_8/i0_3 ), .A3(
        \SB1_3_8/i0_0 ), .ZN(\SB1_3_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2309 ( .A1(\SB1_3_3/i0[6] ), .A2(\SB1_3_3/i0[8] ), .A3(
        \SB1_3_3/i0[7] ), .ZN(n1870) );
  CLKBUF_X4 U2314 ( .I(\SB1_3_9/buf_output[2] ), .Z(\SB2_3_6/i0_0 ) );
  INV_X1 U2315 ( .I(\SB1_3_25/buf_output[0] ), .ZN(\SB2_3_20/i3[0] ) );
  CLKBUF_X4 U2321 ( .I(\SB1_3_1/buf_output[3] ), .Z(\SB2_3_31/i0[10] ) );
  NAND3_X1 U2333 ( .A1(\SB2_3_3/i1_5 ), .A2(\SB2_3_3/i0[6] ), .A3(
        \SB2_3_3/i0[9] ), .ZN(\SB2_3_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2334 ( .A1(\SB2_3_7/i0_0 ), .A2(\SB2_3_7/i0_4 ), .A3(
        \SB2_3_7/i1_5 ), .ZN(n2159) );
  NAND3_X1 U2347 ( .A1(\SB2_3_10/i0[7] ), .A2(\SB2_3_10/i0[8] ), .A3(
        \SB2_3_10/i0[6] ), .ZN(\SB2_3_10/Component_Function_0/NAND4_in[1] ) );
  INV_X1 U2348 ( .I(n147), .ZN(n470) );
  INV_X1 U2352 ( .I(\MC_ARK_ARC_1_3/buf_output[133] ), .ZN(\SB1_4_9/i1_7 ) );
  CLKBUF_X4 U2354 ( .I(\MC_ARK_ARC_1_3/buf_output[171] ), .Z(\SB1_4_3/i0[10] )
         );
  CLKBUF_X4 U2360 ( .I(\MC_ARK_ARC_1_3/buf_output[112] ), .Z(\SB1_4_13/i0_4 )
         );
  NAND3_X1 U2362 ( .A1(\SB1_4_8/i0[10] ), .A2(\SB1_4_8/i1_5 ), .A3(
        \SB1_4_8/i1[9] ), .ZN(n2393) );
  NAND3_X1 U2365 ( .A1(\SB1_4_14/i0[9] ), .A2(\SB1_4_14/i0_0 ), .A3(
        \SB1_4_14/i0[8] ), .ZN(\SB1_4_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2371 ( .A1(\MC_ARK_ARC_1_3/buf_output[6] ), .A2(
        \MC_ARK_ARC_1_3/buf_output[7] ), .A3(\MC_ARK_ARC_1_3/buf_output[10] ), 
        .ZN(\SB1_4_30/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2373 ( .A1(\SB1_4_20/i0[8] ), .A2(\SB1_4_20/i0[7] ), .A3(
        \SB1_4_20/i0[6] ), .ZN(\SB1_4_20/Component_Function_0/NAND4_in[1] ) );
  CLKBUF_X4 U2379 ( .I(\MC_ARK_ARC_1_3/buf_output[187] ), .Z(\SB1_4_0/i0[6] )
         );
  NAND3_X1 U2398 ( .A1(\SB2_4_15/i1_7 ), .A2(\SB2_4_15/i0[8] ), .A3(
        \SB2_4_15/i0_4 ), .ZN(\SB2_4_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2403 ( .A1(\SB2_4_11/i0[9] ), .A2(\SB2_4_11/i0[6] ), .A3(
        \SB2_4_11/i1_5 ), .ZN(n2648) );
  NAND3_X1 U2405 ( .A1(\SB2_4_18/i1[9] ), .A2(\SB2_4_18/i1_5 ), .A3(
        \SB2_4_18/i0_4 ), .ZN(\SB2_4_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2406 ( .A1(\SB1_4_1/buf_output[1] ), .A2(\SB2_4_29/i0_4 ), .A3(
        \SB2_4_29/i0[9] ), .ZN(\SB2_4_29/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2407 ( .A1(\SB2_4_15/i1[9] ), .A2(\SB2_4_15/i1_5 ), .A3(
        \SB2_4_15/i0_4 ), .ZN(\SB2_4_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2411 ( .A1(\SB2_4_23/i0_4 ), .A2(\SB2_4_23/i0[8] ), .A3(
        \SB2_4_23/i1_7 ), .ZN(n611) );
  NAND2_X1 U2416 ( .A1(\SB2_4_25/i0[10] ), .A2(\SB2_4_25/i0[9] ), .ZN(
        \SB2_4_25/Component_Function_0/NAND4_in[0] ) );
  INV_X1 U2417 ( .I(n36), .ZN(n529) );
  INV_X1 U2419 ( .I(n32), .ZN(n461) );
  CLKBUF_X4 U2425 ( .I(\MC_ARK_ARC_1_4/buf_output[8] ), .Z(\SB3_30/i0_0 ) );
  CLKBUF_X4 U2428 ( .I(\MC_ARK_ARC_1_4/buf_output[94] ), .Z(\SB3_16/i0_4 ) );
  CLKBUF_X4 U2430 ( .I(\MC_ARK_ARC_1_4/buf_output[178] ), .Z(\SB3_2/i0_4 ) );
  NAND3_X1 U2431 ( .A1(\SB3_18/i0_3 ), .A2(\SB3_18/i0[8] ), .A3(
        \MC_ARK_ARC_1_4/buf_output[78] ), .ZN(
        \SB3_18/Component_Function_2/NAND4_in[2] ) );
  INV_X1 U2436 ( .I(\MC_ARK_ARC_1_4/buf_output[121] ), .ZN(\SB3_11/i1_7 ) );
  NAND2_X1 U2437 ( .A1(\SB3_29/i0[10] ), .A2(\SB3_29/i0[9] ), .ZN(
        \SB3_29/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U2438 ( .A1(\SB3_25/i1_5 ), .A2(n774), .ZN(
        \SB3_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2439 ( .A1(\SB3_24/i0[8] ), .A2(\SB3_24/i3[0] ), .A3(\SB3_24/i1_5 ), .ZN(n1398) );
  NAND3_X1 U2447 ( .A1(\SB3_8/i1[9] ), .A2(\SB3_8/i0_4 ), .A3(\SB3_8/i0_3 ), 
        .ZN(\SB3_8/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2455 ( .A1(\SB3_17/buf_output[3] ), .A2(\SB4_15/i1[9] ), .A3(
        \SB4_15/i1_7 ), .ZN(n2027) );
  NAND3_X1 U2457 ( .A1(\SB4_8/i0[10] ), .A2(\SB4_8/i0_3 ), .A3(\SB4_8/i0_4 ), 
        .ZN(n1643) );
  NAND2_X1 U2458 ( .A1(\SB4_3/i0_3 ), .A2(\SB4_3/i1[9] ), .ZN(
        \SB4_3/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 U2460 ( .A1(\SB4_31/i0[10] ), .A2(\SB4_31/i0[9] ), .ZN(
        \SB4_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U2469 ( .A1(\SB4_24/i0_0 ), .A2(\SB4_24/i3[0] ), .A3(\SB4_24/i1_7 ), 
        .ZN(n2744) );
  CLKBUF_X2 U2473 ( .I(Key[55]), .Z(n197) );
  XNOR2_X1 U2477 ( .A1(\SB2_0_1/buf_output[5] ), .A2(n102), .ZN(n583) );
  BUF_X2 U2485 ( .I(Key[80]), .Z(n207) );
  NOR2_X1 U2486 ( .A1(\SB1_0_22/buf_output[5] ), .A2(n6288), .ZN(n593) );
  BUF_X2 U2489 ( .I(Key[101]), .Z(n212) );
  CLKBUF_X2 U2490 ( .I(Key[79]), .Z(n190) );
  BUF_X2 U2492 ( .I(Key[148]), .Z(n219) );
  XOR2_X1 U2494 ( .A1(\RI5[0][92] ), .A2(\RI5[0][86] ), .Z(n595) );
  NAND3_X1 U2497 ( .A1(\SB2_0_31/i0_0 ), .A2(\SB2_0_31/i0[9] ), .A3(
        \SB2_0_31/i0[8] ), .ZN(\SB2_0_31/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U2506 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[141] ), .A2(\RI5[2][165] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[3] ) );
  NAND3_X2 U2512 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i0_4 ), .A3(
        \SB2_3_27/i1[9] ), .ZN(n602) );
  NAND4_X2 U2513 ( .A1(\SB1_1_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_2/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_1_2/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_1_2/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_1_2/buf_output[2] ) );
  XOR2_X1 U2514 ( .A1(\RI5[4][56] ), .A2(\RI5[4][20] ), .Z(
        \MC_ARK_ARC_1_4/temp3[146] ) );
  NAND3_X1 U2527 ( .A1(\SB1_4_8/i0[9] ), .A2(\SB1_4_8/i0[6] ), .A3(
        \SB1_4_8/i1_5 ), .ZN(\SB1_4_8/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U2538 ( .A1(\RI5[1][87] ), .A2(\RI5[1][123] ), .Z(
        \MC_ARK_ARC_1_1/temp3[21] ) );
  XOR2_X1 U2543 ( .A1(\RI5[1][33] ), .A2(\RI5[1][69] ), .Z(n610) );
  NAND4_X1 U2546 ( .A1(\SB2_4_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_4_23/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_4_23/Component_Function_1/NAND4_in[2] ), .A4(n611), .ZN(
        \SB2_4_23/buf_output[1] ) );
  XOR2_X1 U2547 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[7] ), .A2(\RI5[1][13] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[13] ) );
  NAND3_X2 U2554 ( .A1(\SB1_1_21/i0_4 ), .A2(\SB1_1_21/i0[8] ), .A3(
        \SB1_1_21/i1_7 ), .ZN(n614) );
  NAND4_X2 U2556 ( .A1(\SB2_1_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_17/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_17/Component_Function_2/NAND4_in[3] ), .A4(n615), .ZN(
        \SB2_1_17/buf_output[2] ) );
  XOR2_X1 U2562 ( .A1(n617), .A2(\MC_ARK_ARC_1_2/temp5[190] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[190] ) );
  XOR2_X1 U2563 ( .A1(\MC_ARK_ARC_1_2/temp3[190] ), .A2(
        \MC_ARK_ARC_1_2/temp4[190] ), .Z(n617) );
  NAND3_X2 U2570 ( .A1(\SB1_0_9/i0_0 ), .A2(\SB1_0_9/i1_5 ), .A3(
        \SB1_0_9/i0_4 ), .ZN(n2432) );
  NAND3_X1 U2573 ( .A1(\SB2_2_3/i0[10] ), .A2(\SB2_2_3/i0_3 ), .A3(
        \SB2_2_3/i0_4 ), .ZN(n621) );
  XOR2_X1 U2578 ( .A1(\MC_ARK_ARC_1_3/temp2[160] ), .A2(
        \MC_ARK_ARC_1_3/temp1[160] ), .Z(\MC_ARK_ARC_1_3/temp5[160] ) );
  BUF_X4 U2583 ( .I(\SB2_4_1/buf_output[1] ), .Z(\RI5[4][13] ) );
  XOR2_X1 U2586 ( .A1(\MC_ARK_ARC_1_4/temp4[8] ), .A2(
        \MC_ARK_ARC_1_4/temp3[8] ), .Z(\MC_ARK_ARC_1_4/temp6[8] ) );
  INV_X2 U2595 ( .I(n630), .ZN(\SB2_0_4/i0[9] ) );
  XOR2_X1 U2599 ( .A1(n2528), .A2(\MC_ARK_ARC_1_4/temp5[25] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[25] ) );
  NAND4_X2 U2600 ( .A1(\SB1_0_3/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_3/Component_Function_5/NAND4_in[2] ), .A3(n1624), .A4(
        \SB1_0_3/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][173] ) );
  NAND3_X1 U2602 ( .A1(\SB2_3_22/i0_0 ), .A2(\SB2_3_22/i0_3 ), .A3(n1763), 
        .ZN(\SB2_3_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U2614 ( .A1(\SB1_2_17/i0_0 ), .A2(\MC_ARK_ARC_1_1/buf_output[88] ), 
        .A3(\SB1_2_17/i1_5 ), .ZN(n633) );
  NAND4_X2 U2618 ( .A1(\SB1_0_20/Component_Function_4/NAND4_in[0] ), .A2(n2482), .A3(\SB1_0_20/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_0_20/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_0_20/buf_output[4] ) );
  XOR2_X1 U2620 ( .A1(\MC_ARK_ARC_1_4/temp4[97] ), .A2(
        \MC_ARK_ARC_1_4/temp3[97] ), .Z(n635) );
  NAND4_X2 U2621 ( .A1(n1000), .A2(\SB1_0_31/Component_Function_4/NAND4_in[0] ), .A3(\SB1_0_31/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_0_31/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][10] ) );
  XOR2_X1 U2637 ( .A1(\RI5[4][69] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[75] ), 
        .Z(n642) );
  INV_X2 U2640 ( .I(\SB1_0_31/buf_output[2] ), .ZN(\SB2_0_28/i1[9] ) );
  NAND4_X2 U2641 ( .A1(\SB1_0_31/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_31/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_31/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_0_31/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_0_31/buf_output[2] ) );
  NAND4_X2 U2642 ( .A1(\SB2_4_17/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_17/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_4_17/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_4_17/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_4_17/buf_output[0] ) );
  XOR2_X1 U2643 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[94] ), .A2(\RI5[4][130] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[28] ) );
  NAND2_X1 U2647 ( .A1(\SB1_1_1/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_1_1/Component_Function_4/NAND4_in[1] ), .ZN(n648) );
  XOR2_X1 U2651 ( .A1(\MC_ARK_ARC_1_2/temp6[166] ), .A2(n650), .Z(
        \MC_ARK_ARC_1_2/buf_output[166] ) );
  XOR2_X1 U2652 ( .A1(\MC_ARK_ARC_1_2/temp1[166] ), .A2(
        \MC_ARK_ARC_1_2/temp2[166] ), .Z(n650) );
  XOR2_X1 U2655 ( .A1(\MC_ARK_ARC_1_3/temp2[169] ), .A2(
        \MC_ARK_ARC_1_3/temp1[169] ), .Z(\MC_ARK_ARC_1_3/temp5[169] ) );
  NAND2_X2 U2657 ( .A1(n2943), .A2(\SB2_1_4/Component_Function_4/NAND4_in[1] ), 
        .ZN(\MC_ARK_ARC_1_1/buf_datainput[172] ) );
  NAND3_X1 U2665 ( .A1(\SB1_4_28/i0_3 ), .A2(\SB1_4_28/i0[7] ), .A3(
        \SB1_4_28/i0_0 ), .ZN(n655) );
  XOR2_X1 U2667 ( .A1(\RI5[0][110] ), .A2(\RI5[0][86] ), .Z(n993) );
  NAND4_X2 U2668 ( .A1(\SB1_1_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_24/Component_Function_0/NAND4_in[0] ), .A4(n656), .ZN(
        \SB1_1_24/buf_output[0] ) );
  XOR2_X1 U2671 ( .A1(\RI5[2][50] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[74] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[104] ) );
  NAND4_X2 U2672 ( .A1(\SB3_27/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_27/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_27/Component_Function_0/NAND4_in[1] ), .A4(
        \SB3_27/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_27/buf_output[0] ) );
  XOR2_X1 U2678 ( .A1(\RI5[4][60] ), .A2(\RI5[4][84] ), .Z(n660) );
  NAND3_X1 U2682 ( .A1(\SB1_4_20/i0_4 ), .A2(\SB1_4_20/i1[9] ), .A3(
        \SB1_4_20/i1_5 ), .ZN(\SB1_4_20/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U2697 ( .A1(\SB2_3_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_16/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_3_16/Component_Function_3/NAND4_in[3] ), .A4(n665), .ZN(
        \SB2_3_16/buf_output[3] ) );
  XOR2_X1 U2701 ( .A1(\MC_ARK_ARC_1_1/temp4[81] ), .A2(
        \MC_ARK_ARC_1_1/temp3[81] ), .Z(n666) );
  BUF_X4 U2703 ( .I(\SB2_0_22/buf_output[1] ), .Z(\RI5[0][79] ) );
  XOR2_X1 U2706 ( .A1(n669), .A2(\MC_ARK_ARC_1_2/temp6[126] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[126] ) );
  XOR2_X1 U2707 ( .A1(\MC_ARK_ARC_1_2/temp1[126] ), .A2(
        \MC_ARK_ARC_1_2/temp2[126] ), .Z(n669) );
  NAND3_X2 U2712 ( .A1(\SB1_2_17/i0_4 ), .A2(\SB1_2_17/i1[9] ), .A3(
        \SB1_2_17/i0_3 ), .ZN(n671) );
  NAND2_X1 U2720 ( .A1(n1591), .A2(\SB1_3_13/Component_Function_4/NAND4_in[3] ), .ZN(n1590) );
  NAND4_X2 U2725 ( .A1(\SB2_1_14/Component_Function_0/NAND4_in[3] ), .A2(n1171), .A3(\SB2_1_14/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_1_14/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_14/buf_output[0] ) );
  XOR2_X1 U2728 ( .A1(\MC_ARK_ARC_1_2/temp4[111] ), .A2(n673), .Z(n940) );
  XOR2_X1 U2729 ( .A1(\RI5[2][177] ), .A2(\RI5[2][21] ), .Z(n673) );
  XOR2_X1 U2732 ( .A1(\MC_ARK_ARC_1_4/temp3[71] ), .A2(
        \MC_ARK_ARC_1_4/temp4[71] ), .Z(n674) );
  XOR2_X1 U2740 ( .A1(\MC_ARK_ARC_1_2/temp3[42] ), .A2(
        \MC_ARK_ARC_1_2/temp4[42] ), .Z(\MC_ARK_ARC_1_2/temp6[42] ) );
  BUF_X4 U2741 ( .I(\SB2_2_23/buf_output[4] ), .Z(\RI5[2][58] ) );
  NAND4_X2 U2757 ( .A1(\SB2_2_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_20/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_20/Component_Function_4/NAND4_in[1] ), .A4(n681), .ZN(
        \SB2_2_20/buf_output[4] ) );
  XOR2_X1 U2761 ( .A1(\MC_ARK_ARC_1_2/temp5[10] ), .A2(n683), .Z(
        \MC_ARK_ARC_1_2/buf_output[10] ) );
  XOR2_X1 U2762 ( .A1(\MC_ARK_ARC_1_2/temp3[10] ), .A2(
        \MC_ARK_ARC_1_2/temp4[10] ), .Z(n683) );
  XOR2_X1 U2766 ( .A1(\MC_ARK_ARC_1_3/temp1[32] ), .A2(
        \MC_ARK_ARC_1_3/temp2[32] ), .Z(n685) );
  XOR2_X1 U2767 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[24] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[60] ), .Z(\MC_ARK_ARC_1_2/temp3[150] )
         );
  NAND3_X2 U2769 ( .A1(\SB2_4_24/i0[10] ), .A2(\SB2_4_24/i0[6] ), .A3(
        \SB2_4_24/i0_0 ), .ZN(n686) );
  NAND3_X2 U2770 ( .A1(\SB1_0_19/i0_4 ), .A2(\SB1_0_19/i0[6] ), .A3(
        \SB1_0_19/i0[9] ), .ZN(\SB1_0_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2772 ( .A1(\SB2_0_6/i0_0 ), .A2(\RI3[0][154] ), .A3(\SB2_0_6/i1_5 ), .ZN(\SB2_0_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U2781 ( .A1(\SB2_1_4/i0_0 ), .A2(\SB2_1_4/i0[10] ), .A3(
        \SB1_1_8/buf_output[1] ), .ZN(n809) );
  XOR2_X1 U2787 ( .A1(\MC_ARK_ARC_1_1/temp1[139] ), .A2(
        \MC_ARK_ARC_1_1/temp2[139] ), .Z(\MC_ARK_ARC_1_1/temp5[139] ) );
  NAND3_X1 U2789 ( .A1(\SB1_4_25/i1_5 ), .A2(\SB1_4_25/i1[9] ), .A3(
        \SB1_4_25/i0_4 ), .ZN(n690) );
  BUF_X4 U2791 ( .I(\SB2_4_20/buf_output[3] ), .Z(\RI5[4][81] ) );
  INV_X2 U2792 ( .I(\SB1_3_17/buf_output[2] ), .ZN(\SB2_3_14/i1[9] ) );
  NAND3_X2 U2797 ( .A1(\SB1_1_21/i0_3 ), .A2(\SB1_1_21/i0_4 ), .A3(
        \SB1_1_21/i0_0 ), .ZN(\SB1_1_21/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U2811 ( .I(\SB3_30/buf_output[5] ), .ZN(\SB4_30/i1_5 ) );
  XOR2_X1 U2815 ( .A1(\MC_ARK_ARC_1_3/temp3[133] ), .A2(
        \MC_ARK_ARC_1_3/temp4[133] ), .Z(\MC_ARK_ARC_1_3/temp6[133] ) );
  NAND3_X1 U2827 ( .A1(\SB4_26/i0_3 ), .A2(\SB3_29/buf_output[2] ), .A3(
        \SB4_26/i0[7] ), .ZN(n702) );
  NAND3_X2 U2832 ( .A1(\SB2_2_5/i0[8] ), .A2(\SB2_2_5/i3[0] ), .A3(
        \SB2_2_5/i1_5 ), .ZN(n2226) );
  NAND3_X2 U2839 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i0[9] ), .A3(
        \SB2_3_27/i0[8] ), .ZN(n706) );
  NAND3_X1 U2840 ( .A1(n3308), .A2(\SB2_3_28/i0[6] ), .A3(\SB2_3_28/i0[8] ), 
        .ZN(\SB2_3_28/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U2846 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[79] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_2/temp3[13] )
         );
  XOR2_X1 U2848 ( .A1(\RI5[2][11] ), .A2(\RI5[2][5] ), .Z(n710) );
  XOR2_X1 U2851 ( .A1(\MC_ARK_ARC_1_4/temp4[36] ), .A2(
        \MC_ARK_ARC_1_4/temp3[36] ), .Z(\MC_ARK_ARC_1_4/temp6[36] ) );
  INV_X2 U2859 ( .I(\SB1_1_2/buf_output[3] ), .ZN(\SB2_1_0/i0[8] ) );
  INV_X2 U2867 ( .I(\SB1_4_8/buf_output[2] ), .ZN(\SB2_4_5/i1[9] ) );
  XOR2_X1 U2870 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[122] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[146] ), .Z(n1645) );
  BUF_X4 U2871 ( .I(\MC_ARK_ARC_1_3/buf_output[107] ), .Z(\SB1_4_14/i0_3 ) );
  XOR2_X1 U2872 ( .A1(n716), .A2(\MC_ARK_ARC_1_2/temp3[117] ), .Z(n1431) );
  XOR2_X1 U2873 ( .A1(\RI5[2][87] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[63] ), 
        .Z(n716) );
  INV_X2 U2885 ( .I(\SB1_1_3/buf_output[5] ), .ZN(\SB2_1_3/i1_5 ) );
  XOR2_X1 U2888 ( .A1(\RI5[4][51] ), .A2(\RI5[4][57] ), .Z(
        \MC_ARK_ARC_1_4/temp1[57] ) );
  XOR2_X1 U2892 ( .A1(\MC_ARK_ARC_1_2/temp5[154] ), .A2(n724), .Z(
        \MC_ARK_ARC_1_2/buf_output[154] ) );
  XOR2_X1 U2893 ( .A1(\MC_ARK_ARC_1_2/temp3[154] ), .A2(
        \MC_ARK_ARC_1_2/temp4[154] ), .Z(n724) );
  BUF_X4 U2894 ( .I(\SB2_2_29/buf_output[1] ), .Z(\RI5[2][37] ) );
  XOR2_X1 U2898 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[183] ), .A2(\RI5[3][27] ), 
        .Z(n727) );
  XOR2_X1 U2911 ( .A1(\MC_ARK_ARC_1_0/temp3[181] ), .A2(
        \MC_ARK_ARC_1_0/temp4[181] ), .Z(n733) );
  XOR2_X1 U2912 ( .A1(\MC_ARK_ARC_1_1/temp1[67] ), .A2(
        \MC_ARK_ARC_1_1/temp2[67] ), .Z(\MC_ARK_ARC_1_1/temp5[67] ) );
  XOR2_X1 U2930 ( .A1(n2985), .A2(\MC_ARK_ARC_1_4/temp6[188] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[188] ) );
  XOR2_X1 U2931 ( .A1(\MC_ARK_ARC_1_4/temp6[112] ), .A2(
        \MC_ARK_ARC_1_4/temp5[112] ), .Z(\MC_ARK_ARC_1_4/buf_output[112] ) );
  XOR2_X1 U2937 ( .A1(\RI5[3][137] ), .A2(n167), .Z(n741) );
  XOR2_X1 U2938 ( .A1(\RI5[3][101] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .Z(n742) );
  XOR2_X1 U2961 ( .A1(\RI5[2][116] ), .A2(\RI5[2][80] ), .Z(n753) );
  NAND3_X1 U2976 ( .A1(\SB1_3_23/i0[8] ), .A2(\SB1_3_23/i0_4 ), .A3(
        \SB1_3_23/i1_7 ), .ZN(n759) );
  XOR2_X1 U2980 ( .A1(n761), .A2(\MC_ARK_ARC_1_1/temp6[180] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[180] ) );
  XOR2_X1 U2981 ( .A1(\MC_ARK_ARC_1_1/temp1[180] ), .A2(
        \MC_ARK_ARC_1_1/temp2[180] ), .Z(n761) );
  XOR2_X1 U2982 ( .A1(\MC_ARK_ARC_1_2/temp6[156] ), .A2(
        \MC_ARK_ARC_1_2/temp5[156] ), .Z(\MC_ARK_ARC_1_2/buf_output[156] ) );
  BUF_X4 U2985 ( .I(\SB2_2_23/buf_output[1] ), .Z(\RI5[2][73] ) );
  XOR2_X1 U2987 ( .A1(\MC_ARK_ARC_1_4/temp4[31] ), .A2(
        \MC_ARK_ARC_1_4/temp3[31] ), .Z(n763) );
  NAND4_X2 U2988 ( .A1(\SB1_2_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_28/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_28/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_28/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_28/buf_output[0] ) );
  NAND3_X2 U2995 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0[9] ), .A3(
        \SB1_0_2/i0[10] ), .ZN(\SB1_0_2/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 U2996 ( .I(\SB2_4_17/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[94] ) );
  NAND3_X1 U3006 ( .A1(\SB4_18/i0[9] ), .A2(\SB4_18/i1_5 ), .A3(\SB4_18/i0[6] ), .ZN(\SB4_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3019 ( .A1(\SB1_4_8/i0[10] ), .A2(\SB1_4_8/i0_3 ), .A3(
        \SB1_4_8/i0[6] ), .ZN(\SB1_4_8/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U3024 ( .A1(\RI5[0][99] ), .A2(\RI5[0][63] ), .Z(
        \MC_ARK_ARC_1_0/temp3[189] ) );
  NAND4_X2 U3030 ( .A1(\SB1_0_16/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_16/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_16/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_16/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][120] ) );
  XOR2_X1 U3033 ( .A1(n578), .A2(\MC_ARK_ARC_1_1/buf_datainput[4] ), .Z(
        \MC_ARK_ARC_1_1/temp2[34] ) );
  XOR2_X1 U3038 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[151] ), .A2(\RI5[1][175] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[13] ) );
  XOR2_X1 U3053 ( .A1(\MC_ARK_ARC_1_3/temp3[57] ), .A2(
        \MC_ARK_ARC_1_3/temp4[57] ), .Z(\MC_ARK_ARC_1_3/temp6[57] ) );
  NAND3_X2 U3055 ( .A1(\SB1_2_13/i0[6] ), .A2(\SB1_2_13/i0_4 ), .A3(
        \SB1_2_13/i0[9] ), .ZN(n784) );
  NAND3_X2 U3066 ( .A1(\SB2_4_24/i0_4 ), .A2(\SB2_4_24/i0_0 ), .A3(n6268), 
        .ZN(\SB2_4_24/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U3073 ( .A1(\MC_ARK_ARC_1_2/temp3[85] ), .A2(
        \MC_ARK_ARC_1_2/temp4[85] ), .Z(n790) );
  NAND4_X2 U3083 ( .A1(\SB2_4_29/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_29/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_4_29/Component_Function_0/NAND4_in[0] ), .A4(n795), .ZN(
        \SB2_4_29/buf_output[0] ) );
  XOR2_X1 U3087 ( .A1(\MC_ARK_ARC_1_3/temp5[16] ), .A2(n797), .Z(
        \MC_ARK_ARC_1_3/buf_output[16] ) );
  XOR2_X1 U3088 ( .A1(\MC_ARK_ARC_1_3/temp3[16] ), .A2(
        \MC_ARK_ARC_1_3/temp4[16] ), .Z(n797) );
  XOR2_X1 U3094 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[15] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[21] ), .Z(n801) );
  XOR2_X1 U3098 ( .A1(\RI5[0][62] ), .A2(\RI5[0][68] ), .Z(n802) );
  XOR2_X1 U3107 ( .A1(\SB2_1_31/buf_output[0] ), .A2(\RI5[1][186] ), .Z(n806)
         );
  XOR2_X1 U3122 ( .A1(\MC_ARK_ARC_1_4/temp2[110] ), .A2(n813), .Z(n2980) );
  XOR2_X1 U3123 ( .A1(\RI5[4][104] ), .A2(\RI5[4][110] ), .Z(n813) );
  XOR2_X1 U3136 ( .A1(\MC_ARK_ARC_1_1/temp1[124] ), .A2(
        \MC_ARK_ARC_1_1/temp2[124] ), .Z(n817) );
  NAND3_X1 U3137 ( .A1(\SB1_0_26/i0_3 ), .A2(\SB1_0_26/i1[9] ), .A3(
        \SB1_0_26/i0_4 ), .ZN(\SB1_0_26/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U3146 ( .A1(\SB2_3_22/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_22/Component_Function_0/NAND4_in[1] ), .A3(n2033), .A4(
        \SB2_3_22/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_22/buf_output[0] ) );
  NAND3_X1 U3150 ( .A1(\RI3[0][4] ), .A2(\SB1_0_2/buf_output[2] ), .A3(
        \SB2_0_31/i1_5 ), .ZN(\SB2_0_31/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U3153 ( .A1(\SB1_2_15/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_15/Component_Function_1/NAND4_in[2] ), .A3(n2140), .A4(
        \SB1_2_15/Component_Function_1/NAND4_in[1] ), .ZN(\RI3[2][121] ) );
  XOR2_X1 U3165 ( .A1(\MC_ARK_ARC_1_0/temp1[98] ), .A2(n823), .Z(n3012) );
  XOR2_X1 U3166 ( .A1(\RI5[0][68] ), .A2(\RI5[0][44] ), .Z(n823) );
  XOR2_X1 U3169 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[73] ), .A2(\RI5[1][109] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[7] ) );
  NAND4_X2 U3173 ( .A1(\SB1_2_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_2_21/Component_Function_3/NAND4_in[3] ), .A4(n826), .ZN(
        \SB1_2_21/buf_output[3] ) );
  NAND3_X2 U3174 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i0_0 ), .A3(
        \SB1_2_21/i0_4 ), .ZN(n826) );
  NAND3_X1 U3176 ( .A1(\SB1_0_18/i0[6] ), .A2(\SB1_0_18/i0[8] ), .A3(
        \SB1_0_18/i0[7] ), .ZN(\SB1_0_18/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U3178 ( .A1(\SB1_0_3/i0[10] ), .A2(\SB1_0_3/i1[9] ), .A3(
        \SB1_0_3/i1_7 ), .ZN(n833) );
  NAND4_X2 U3184 ( .A1(\SB2_2_3/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_3/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_3/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_3/buf_output[1] ) );
  NAND4_X2 U3185 ( .A1(\SB2_2_0/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_0/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_0/Component_Function_4/NAND4_in[3] ), .A4(n829), .ZN(
        \SB2_2_0/buf_output[4] ) );
  NAND3_X2 U3186 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0[9] ), .A3(
        \SB2_2_0/i0[10] ), .ZN(n829) );
  INV_X1 U3188 ( .I(\SB3_26/buf_output[1] ), .ZN(\SB4_22/i1_7 ) );
  NAND4_X2 U3189 ( .A1(\SB3_26/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_26/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_26/buf_output[1] ) );
  NAND3_X2 U3191 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0_0 ), .A3(n5444), .ZN(
        \SB2_2_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U3194 ( .A1(\SB1_4_0/i0[10] ), .A2(\SB1_4_0/i0[6] ), .A3(
        \SB1_4_0/i0_0 ), .ZN(n830) );
  XOR2_X1 U3200 ( .A1(\RI5[3][6] ), .A2(\RI5[3][12] ), .Z(
        \MC_ARK_ARC_1_3/temp1[12] ) );
  NAND3_X2 U3206 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i0[10] ), .A3(
        \SB1_1_2/i0[6] ), .ZN(n836) );
  XOR2_X1 U3224 ( .A1(\RI5[2][95] ), .A2(\RI5[2][161] ), .Z(n845) );
  NAND3_X2 U3227 ( .A1(\SB2_1_0/i0[6] ), .A2(n590), .A3(\SB2_1_0/i0[9] ), .ZN(
        n914) );
  NAND4_X2 U3228 ( .A1(\SB2_0_9/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_9/Component_Function_3/NAND4_in[1] ), .A3(n2835), .A4(
        \SB2_0_9/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB2_0_9/buf_output[3] ) );
  XOR2_X1 U3233 ( .A1(n849), .A2(\MC_ARK_ARC_1_4/temp5[137] ), .Z(
        \RI1[5][137] ) );
  XOR2_X1 U3234 ( .A1(\MC_ARK_ARC_1_4/temp4[137] ), .A2(
        \MC_ARK_ARC_1_4/temp3[137] ), .Z(n849) );
  NAND4_X2 U3235 ( .A1(\SB1_2_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_21/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_21/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_21/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_21/buf_output[0] ) );
  XOR2_X1 U3238 ( .A1(\MC_ARK_ARC_1_0/temp6[184] ), .A2(
        \MC_ARK_ARC_1_0/temp5[184] ), .Z(\MC_ARK_ARC_1_0/buf_output[184] ) );
  BUF_X4 U3239 ( .I(\SB2_3_10/i0_4 ), .Z(n851) );
  NAND3_X2 U3241 ( .A1(\SB1_0_8/i0_4 ), .A2(\SB1_0_8/i0_3 ), .A3(
        \SB1_0_8/i1[9] ), .ZN(n2672) );
  XOR2_X1 U3243 ( .A1(\RI5[0][100] ), .A2(\RI5[0][124] ), .Z(
        \MC_ARK_ARC_1_0/temp2[154] ) );
  NAND3_X2 U3246 ( .A1(\SB2_3_3/i0_3 ), .A2(\SB2_3_3/i0[9] ), .A3(
        \SB2_3_3/i0[8] ), .ZN(n1034) );
  XOR2_X1 U3249 ( .A1(n853), .A2(\MC_ARK_ARC_1_1/temp4[101] ), .Z(n1532) );
  XOR2_X1 U3250 ( .A1(\RI5[1][167] ), .A2(\RI5[1][11] ), .Z(n853) );
  XOR2_X1 U3252 ( .A1(\RI5[3][136] ), .A2(\RI5[3][172] ), .Z(
        \MC_ARK_ARC_1_3/temp3[70] ) );
  XOR2_X1 U3253 ( .A1(n855), .A2(n854), .Z(\MC_ARK_ARC_1_0/buf_output[123] )
         );
  XOR2_X1 U3254 ( .A1(\MC_ARK_ARC_1_0/temp3[123] ), .A2(
        \MC_ARK_ARC_1_0/temp4[123] ), .Z(n854) );
  NAND3_X1 U3256 ( .A1(\SB2_0_14/i0_0 ), .A2(\SB2_0_14/i0[10] ), .A3(
        \SB2_0_14/i0[6] ), .ZN(\SB2_0_14/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U3281 ( .A1(n1095), .A2(\SB2_2_18/Component_Function_3/NAND4_in[1] ), .A3(\SB2_2_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_18/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_18/buf_output[3] ) );
  XOR2_X1 U3293 ( .A1(\MC_ARK_ARC_1_0/temp2[138] ), .A2(
        \MC_ARK_ARC_1_0/temp1[138] ), .Z(n869) );
  NAND3_X2 U3297 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i1_7 ), .A3(
        \SB2_3_19/i1[9] ), .ZN(n871) );
  XOR2_X1 U3310 ( .A1(n879), .A2(n878), .Z(Ciphertext[25]) );
  INV_X1 U3311 ( .I(n168), .ZN(n878) );
  NOR2_X1 U3312 ( .A1(n881), .A2(n880), .ZN(n879) );
  NAND2_X1 U3313 ( .A1(\SB4_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_27/Component_Function_1/NAND4_in[0] ), .ZN(n880) );
  NAND2_X1 U3314 ( .A1(\SB4_27/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_27/Component_Function_1/NAND4_in[3] ), .ZN(n881) );
  NAND4_X2 U3319 ( .A1(\SB3_17/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_17/Component_Function_1/NAND4_in[2] ), .A3(
        \SB3_17/Component_Function_1/NAND4_in[0] ), .A4(n883), .ZN(
        \SB3_17/buf_output[1] ) );
  NAND3_X2 U3320 ( .A1(\SB3_17/i0_4 ), .A2(\SB3_17/i0[8] ), .A3(\SB3_17/i1_7 ), 
        .ZN(n883) );
  XOR2_X1 U3325 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), .A2(\RI5[2][32] ), 
        .Z(n885) );
  NAND2_X1 U3335 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i0[9] ), .ZN(
        \SB4_10/Component_Function_0/NAND4_in[0] ) );
  INV_X1 U3338 ( .I(\SB3_24/buf_output[3] ), .ZN(\SB4_22/i0[8] ) );
  NAND3_X2 U3345 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0[6] ), .A3(
        \SB2_2_23/i1[9] ), .ZN(\SB2_2_23/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U3346 ( .A1(\MC_ARK_ARC_1_4/temp4[28] ), .A2(
        \MC_ARK_ARC_1_4/temp3[28] ), .Z(\MC_ARK_ARC_1_4/temp6[28] ) );
  INV_X2 U3353 ( .I(\SB1_2_31/buf_output[2] ), .ZN(\SB2_2_28/i1[9] ) );
  BUF_X4 U3355 ( .I(\MC_ARK_ARC_1_1/buf_output[26] ), .Z(\SB1_2_27/i0_0 ) );
  NAND3_X2 U3359 ( .A1(\SB1_2_27/i0_0 ), .A2(\SB1_2_27/i3[0] ), .A3(
        \SB1_2_27/i1_7 ), .ZN(\SB1_2_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3361 ( .A1(\SB3_24/i0_0 ), .A2(\SB3_24/i0[10] ), .A3(
        \SB3_24/i0[6] ), .ZN(\SB3_24/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U3362 ( .A1(\SB3_13/i0[10] ), .A2(\SB3_13/i0_0 ), .A3(
        \SB3_13/i0[6] ), .ZN(\SB3_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3376 ( .A1(\SB4_27/i0[6] ), .A2(\SB4_27/i0[7] ), .A3(
        \SB4_27/i0[8] ), .ZN(n898) );
  NAND3_X1 U3381 ( .A1(\SB1_0_18/i0_4 ), .A2(n279), .A3(n234), .ZN(n901) );
  XOR2_X1 U3388 ( .A1(n906), .A2(n905), .Z(\MC_ARK_ARC_1_4/buf_output[189] )
         );
  XOR2_X1 U3390 ( .A1(\MC_ARK_ARC_1_3/temp2[93] ), .A2(n907), .Z(
        \MC_ARK_ARC_1_3/temp5[93] ) );
  XOR2_X1 U3398 ( .A1(\MC_ARK_ARC_1_2/temp1[117] ), .A2(
        \MC_ARK_ARC_1_2/temp4[117] ), .Z(n1432) );
  NAND3_X1 U3402 ( .A1(\SB2_2_26/i0[7] ), .A2(\SB2_2_26/i0[8] ), .A3(
        \SB2_2_26/i0[6] ), .ZN(\SB2_2_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U3403 ( .A1(\SB2_0_19/i1_5 ), .A2(\RI3[0][75] ), .A3(
        \SB2_0_19/i1[9] ), .ZN(\SB2_0_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U3404 ( .A1(\SB2_1_24/i0[10] ), .A2(\SB2_1_24/i1_5 ), .A3(
        \SB2_1_24/i1[9] ), .ZN(\SB2_1_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U3415 ( .A1(\SB1_3_14/i0[10] ), .A2(\SB1_3_14/i1[9] ), .A3(
        \SB1_3_14/i1_7 ), .ZN(n913) );
  NAND4_X2 U3419 ( .A1(\SB1_1_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_1/Component_Function_3/NAND4_in[2] ), .A3(n2861), .A4(n3092), 
        .ZN(\SB1_1_1/buf_output[3] ) );
  NAND3_X1 U3420 ( .A1(\SB3_24/buf_output[2] ), .A2(\SB4_21/i0[9] ), .A3(
        \SB4_21/i0[8] ), .ZN(\SB4_21/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U3423 ( .A1(\SB3_24/Component_Function_0/NAND4_in[1] ), .A2(
        \SB3_24/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_24/Component_Function_0/NAND4_in[3] ), .A4(
        \SB3_24/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_24/buf_output[0] ) );
  NAND3_X2 U3431 ( .A1(\SB1_2_24/i0[9] ), .A2(\SB1_2_24/i0_0 ), .A3(
        \SB1_2_24/i0[8] ), .ZN(n919) );
  XOR2_X1 U3443 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[80] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[116] ), .Z(\MC_ARK_ARC_1_3/temp3[14] )
         );
  INV_X2 U3444 ( .I(\MC_ARK_ARC_1_4/buf_output[39] ), .ZN(\SB3_25/i0[8] ) );
  XOR2_X1 U3445 ( .A1(\MC_ARK_ARC_1_1/temp5[94] ), .A2(
        \MC_ARK_ARC_1_1/temp6[94] ), .Z(\MC_ARK_ARC_1_1/buf_output[94] ) );
  NAND4_X2 U3458 ( .A1(\SB3_24/Component_Function_5/NAND4_in[1] ), .A2(n966), 
        .A3(\SB3_24/Component_Function_5/NAND4_in[3] ), .A4(
        \SB3_24/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_24/buf_output[5] ) );
  INV_X2 U3459 ( .I(\SB1_1_7/buf_output[3] ), .ZN(\SB2_1_5/i0[8] ) );
  XOR2_X1 U3471 ( .A1(\MC_ARK_ARC_1_2/temp3[90] ), .A2(
        \MC_ARK_ARC_1_2/temp4[90] ), .Z(\MC_ARK_ARC_1_2/temp6[90] ) );
  XOR2_X1 U3472 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[122] ), .A2(\RI5[1][98] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[152] ) );
  XOR2_X1 U3473 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[122] ), .A2(\RI5[1][116] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[122] ) );
  NOR2_X2 U3474 ( .A1(n2328), .A2(n931), .ZN(\SB2_0_24/i0[7] ) );
  NAND3_X2 U3477 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0_0 ), .A3(
        \SB2_1_10/i0_4 ), .ZN(n932) );
  INV_X1 U3478 ( .I(\SB1_0_22/buf_output[5] ), .ZN(\SB2_0_22/i1_5 ) );
  BUF_X4 U3479 ( .I(\SB2_3_27/buf_output[0] ), .Z(\RI5[3][54] ) );
  XOR2_X1 U3481 ( .A1(\MC_ARK_ARC_1_3/temp4[18] ), .A2(
        \MC_ARK_ARC_1_3/temp3[18] ), .Z(n933) );
  NAND3_X1 U3485 ( .A1(\SB2_1_2/i0_3 ), .A2(\SB1_1_7/buf_output[0] ), .A3(
        \SB2_1_2/i0[8] ), .ZN(\SB2_1_2/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U3488 ( .A1(\RI5[0][191] ), .A2(\RI5[0][23] ), .Z(
        \MC_ARK_ARC_1_0/temp2[53] ) );
  XOR2_X1 U3494 ( .A1(\RI5[1][86] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .Z(n2951) );
  NAND3_X2 U3505 ( .A1(\SB2_2_18/i0[6] ), .A2(\SB2_2_18/i0_4 ), .A3(
        \SB2_2_18/i0[9] ), .ZN(\SB2_2_18/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U3507 ( .A1(\SB2_2_24/i0[10] ), .A2(\SB2_2_24/i0_0 ), .A3(
        \SB2_2_24/i0[6] ), .ZN(n1962) );
  NAND3_X2 U3508 ( .A1(\SB2_4_17/i0[10] ), .A2(\SB2_4_17/i1_7 ), .A3(
        \SB2_4_17/i1[9] ), .ZN(n939) );
  XOR2_X1 U3516 ( .A1(\MC_ARK_ARC_1_3/temp5[116] ), .A2(
        \MC_ARK_ARC_1_3/temp6[116] ), .Z(\MC_ARK_ARC_1_3/buf_output[116] ) );
  XOR2_X1 U3517 ( .A1(n2537), .A2(\MC_ARK_ARC_1_4/temp5[122] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[122] ) );
  NAND3_X2 U3524 ( .A1(\SB2_0_17/i0_3 ), .A2(\RI3[0][88] ), .A3(
        \SB2_0_17/i1[9] ), .ZN(\SB2_0_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3525 ( .A1(\SB2_2_4/i0_0 ), .A2(\SB2_2_4/i3[0] ), .A3(
        \SB2_2_4/i1_7 ), .ZN(\SB2_2_4/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U3527 ( .A1(\SB1_2_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_6/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_6/Component_Function_1/NAND4_in[0] ), .A4(n944), .ZN(
        \SB1_2_6/buf_output[1] ) );
  XOR2_X1 U3528 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[137] ), .A2(\RI5[0][131] ), 
        .Z(n945) );
  NAND3_X2 U3533 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0[10] ), .A3(
        \SB2_2_16/i0[9] ), .ZN(n1097) );
  INV_X2 U3536 ( .I(\SB3_18/buf_output[3] ), .ZN(\SB4_16/i0[8] ) );
  NAND3_X1 U3538 ( .A1(\SB2_3_6/i0_3 ), .A2(\SB2_3_6/i0[7] ), .A3(
        \SB2_3_6/i0_0 ), .ZN(\SB2_3_6/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U3548 ( .A1(\RI5[2][157] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[121] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[55] ) );
  INV_X2 U3551 ( .I(\SB1_1_20/buf_output[2] ), .ZN(\SB2_1_17/i1[9] ) );
  AND2_X1 U3558 ( .A1(\SB1_3_6/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_3_6/Component_Function_4/NAND4_in[1] ), .Z(n959) );
  NAND3_X2 U3560 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0_0 ), .A3(
        \SB2_2_14/i0_4 ), .ZN(\SB2_2_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U3565 ( .A1(\SB2_3_27/i0[10] ), .A2(\SB2_3_27/i1_5 ), .A3(
        \SB2_3_27/i1[9] ), .ZN(\SB2_3_27/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U3572 ( .A1(n964), .A2(n965), .Z(\MC_ARK_ARC_1_1/buf_output[103] )
         );
  XOR2_X1 U3573 ( .A1(\MC_ARK_ARC_1_1/temp3[103] ), .A2(
        \MC_ARK_ARC_1_1/temp2[103] ), .Z(n964) );
  XOR2_X1 U3574 ( .A1(\MC_ARK_ARC_1_1/temp4[103] ), .A2(
        \MC_ARK_ARC_1_1/temp1[103] ), .Z(n965) );
  NAND3_X1 U3576 ( .A1(\SB4_30/i0[6] ), .A2(\SB4_30/i0[9] ), .A3(\SB4_30/i1_5 ), .ZN(\SB4_30/Component_Function_1/NAND4_in[2] ) );
  INV_X2 U3582 ( .I(\SB1_2_6/buf_output[2] ), .ZN(\SB2_2_3/i1[9] ) );
  NAND4_X2 U3585 ( .A1(\SB2_1_17/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_17/Component_Function_4/NAND4_in[0] ), .A4(n969), .ZN(
        \SB2_1_17/buf_output[4] ) );
  NAND4_X2 U3586 ( .A1(\SB2_1_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_19/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_1_19/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_1_19/buf_output[3] ) );
  XOR2_X1 U3589 ( .A1(\RI5[1][120] ), .A2(\RI5[1][114] ), .Z(n971) );
  XOR2_X1 U3592 ( .A1(n1949), .A2(n973), .Z(\MC_ARK_ARC_1_2/buf_output[55] )
         );
  XOR2_X1 U3593 ( .A1(\MC_ARK_ARC_1_2/temp2[55] ), .A2(
        \MC_ARK_ARC_1_2/temp1[55] ), .Z(n973) );
  INV_X2 U3600 ( .I(\SB1_1_26/buf_output[5] ), .ZN(\SB2_1_26/i1_5 ) );
  XOR2_X1 U3603 ( .A1(\MC_ARK_ARC_1_3/temp1[145] ), .A2(n979), .Z(
        \MC_ARK_ARC_1_3/temp5[145] ) );
  XOR2_X1 U3604 ( .A1(\RI5[3][91] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[115] ), 
        .Z(n979) );
  XOR2_X1 U3615 ( .A1(n986), .A2(\MC_ARK_ARC_1_1/temp5[181] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[181] ) );
  XOR2_X1 U3616 ( .A1(\MC_ARK_ARC_1_1/temp4[181] ), .A2(
        \MC_ARK_ARC_1_1/temp3[181] ), .Z(n986) );
  BUF_X4 U3617 ( .I(\SB2_1_20/buf_output[1] ), .Z(\RI5[1][91] ) );
  NAND3_X1 U3630 ( .A1(\SB1_3_19/i0_0 ), .A2(\SB1_3_19/i3[0] ), .A3(
        \SB1_3_19/i1_7 ), .ZN(\SB1_3_19/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U3632 ( .A1(\MC_ARK_ARC_1_3/temp2[122] ), .A2(n994), .Z(
        \MC_ARK_ARC_1_3/temp5[122] ) );
  XOR2_X1 U3633 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), .A2(\RI5[3][122] ), 
        .Z(n994) );
  NAND4_X2 U3635 ( .A1(\SB1_3_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_0/NAND4_in[0] ), .A4(n996), .ZN(
        \SB1_3_19/buf_output[0] ) );
  NAND4_X2 U3640 ( .A1(\SB1_0_16/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_16/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_16/Component_Function_5/NAND4_in[0] ), .A4(n1862), .ZN(
        \RI3[0][95] ) );
  NAND3_X1 U3642 ( .A1(\SB4_16/i3[0] ), .A2(\SB4_16/i0[8] ), .A3(\SB4_16/i1_5 ), .ZN(\SB4_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3644 ( .A1(\SB1_4_15/i0[9] ), .A2(\SB1_4_15/i0_3 ), .A3(
        \SB1_4_15/i0[10] ), .ZN(\SB1_4_15/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U3646 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i1_5 ), .A3(n3973), .ZN(
        \SB4_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U3649 ( .A1(\SB1_0_24/i0_3 ), .A2(\SB1_0_24/i0[10] ), .A3(
        \SB1_0_24/i0_4 ), .ZN(\SB1_0_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3651 ( .A1(n1953), .A2(\SB2_3_9/i0_0 ), .A3(\SB2_3_9/i0_3 ), .ZN(
        \SB2_3_9/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U3652 ( .A1(n2584), .A2(\SB1_4_3/Component_Function_5/NAND4_in[1] ), 
        .A3(n1142), .A4(\SB1_4_3/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_4_3/buf_output[5] ) );
  XOR2_X1 U3659 ( .A1(\MC_ARK_ARC_1_3/temp6[84] ), .A2(
        \MC_ARK_ARC_1_3/temp5[84] ), .Z(\MC_ARK_ARC_1_3/buf_output[84] ) );
  XOR2_X1 U3660 ( .A1(\MC_ARK_ARC_1_1/temp6[68] ), .A2(
        \MC_ARK_ARC_1_1/temp5[68] ), .Z(\MC_ARK_ARC_1_1/buf_output[68] ) );
  NAND3_X1 U3665 ( .A1(\SB1_0_31/i0[10] ), .A2(\SB1_0_31/i0_3 ), .A3(
        \SB1_0_31/i0[9] ), .ZN(n1000) );
  XOR2_X1 U3666 ( .A1(n578), .A2(\MC_ARK_ARC_1_1/buf_datainput[178] ), .Z(
        \MC_ARK_ARC_1_1/temp1[178] ) );
  XOR2_X1 U3669 ( .A1(n1002), .A2(\MC_ARK_ARC_1_1/temp4[79] ), .Z(
        \MC_ARK_ARC_1_1/temp6[79] ) );
  XOR2_X1 U3670 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[145] ), .A2(\RI5[1][181] ), 
        .Z(n1002) );
  XOR2_X1 U3671 ( .A1(\MC_ARK_ARC_1_2/temp4[171] ), .A2(n1003), .Z(
        \MC_ARK_ARC_1_2/temp6[171] ) );
  XOR2_X1 U3672 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[45] ), .A2(\RI5[2][81] ), 
        .Z(n1003) );
  XOR2_X1 U3673 ( .A1(n1967), .A2(n1004), .Z(\MC_ARK_ARC_1_2/buf_output[78] )
         );
  XOR2_X1 U3674 ( .A1(\MC_ARK_ARC_1_2/temp3[78] ), .A2(
        \MC_ARK_ARC_1_2/temp4[78] ), .Z(n1004) );
  XOR2_X1 U3676 ( .A1(\RI5[0][26] ), .A2(\RI5[0][182] ), .Z(n1005) );
  INV_X2 U3684 ( .I(\SB1_1_25/buf_output[5] ), .ZN(\SB2_1_25/i1_5 ) );
  NAND3_X2 U3685 ( .A1(\SB2_1_25/i3[0] ), .A2(\SB2_1_25/i1_5 ), .A3(n3995), 
        .ZN(n1372) );
  XOR2_X1 U3687 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[168] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[12] ), .Z(\MC_ARK_ARC_1_4/temp3[102] )
         );
  INV_X2 U3688 ( .I(\SB1_2_24/buf_output[3] ), .ZN(\SB2_2_22/i0[8] ) );
  XOR2_X1 U3692 ( .A1(\MC_ARK_ARC_1_3/temp1[74] ), .A2(n1010), .Z(n3141) );
  XOR2_X1 U3693 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[20] ), .A2(\RI5[3][44] ), 
        .Z(n1010) );
  XOR2_X1 U3699 ( .A1(\RI5[3][9] ), .A2(\RI5[3][45] ), .Z(n1014) );
  XOR2_X1 U3712 ( .A1(\RI5[1][174] ), .A2(\RI5[1][180] ), .Z(
        \MC_ARK_ARC_1_1/temp1[180] ) );
  NAND3_X2 U3720 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i0_0 ), .A3(
        \SB4_16/i0[6] ), .ZN(n1020) );
  NAND3_X2 U3727 ( .A1(\SB2_1_31/i0_0 ), .A2(n5430), .A3(\SB2_1_31/i0_3 ), 
        .ZN(n2266) );
  XOR2_X1 U3736 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[80] ), .A2(\RI5[3][86] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[86] ) );
  NAND4_X2 U3737 ( .A1(\SB2_2_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_2/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_2/Component_Function_3/NAND4_in[2] ), .A4(n1704), .ZN(
        \SB2_2_2/buf_output[3] ) );
  NAND3_X1 U3738 ( .A1(\SB4_19/i0[10] ), .A2(n6273), .A3(\SB4_19/i1[9] ), .ZN(
        n1030) );
  NAND3_X1 U3744 ( .A1(\SB4_18/i0_3 ), .A2(n1496), .A3(\SB4_18/i0_4 ), .ZN(
        \SB4_18/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U3751 ( .I(\SB2_4_11/buf_output[5] ), .Z(\RI5[4][125] ) );
  INV_X8 U3752 ( .I(n1032), .ZN(\RI1[2][119] ) );
  INV_X2 U3753 ( .I(\MC_ARK_ARC_1_1/buf_output[119] ), .ZN(n1032) );
  XOR2_X1 U3757 ( .A1(\RI5[1][116] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .Z(n1090) );
  INV_X2 U3764 ( .I(\SB1_2_25/buf_output[2] ), .ZN(\SB2_2_22/i1[9] ) );
  XOR2_X1 U3782 ( .A1(\MC_ARK_ARC_1_3/temp2[13] ), .A2(n1046), .Z(
        \MC_ARK_ARC_1_3/temp5[13] ) );
  XOR2_X1 U3783 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[7] ), .A2(\RI5[3][13] ), 
        .Z(n1046) );
  XOR2_X1 U3785 ( .A1(\MC_ARK_ARC_1_0/temp6[171] ), .A2(n1047), .Z(
        \MC_ARK_ARC_1_0/buf_output[171] ) );
  NAND4_X2 U3788 ( .A1(\SB2_3_2/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_2/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_3_2/Component_Function_1/NAND4_in[2] ), .A4(n1048), .ZN(
        \SB2_3_2/buf_output[1] ) );
  NAND2_X2 U3789 ( .A1(\SB1_3_17/i0[9] ), .A2(n588), .ZN(
        \SB1_3_17/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U3792 ( .A1(\SB2_2_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_27/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_2_27/Component_Function_3/NAND4_in[1] ), .A4(n1923), .ZN(
        \SB2_2_27/buf_output[3] ) );
  BUF_X4 U3801 ( .I(\MC_ARK_ARC_1_2/buf_output[3] ), .Z(\SB1_3_31/i0[10] ) );
  XOR2_X1 U3817 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[182] ), .A2(n82), .Z(n1062) );
  XOR2_X1 U3818 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[182] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[188] ), .Z(\MC_ARK_ARC_1_1/temp1[188] )
         );
  XOR2_X1 U3825 ( .A1(\MC_ARK_ARC_1_3/temp3[75] ), .A2(
        \MC_ARK_ARC_1_3/temp4[75] ), .Z(n1066) );
  NAND4_X2 U3826 ( .A1(\SB2_2_16/Component_Function_0/NAND4_in[1] ), .A2(n1067), .A3(n1983), .A4(\SB2_2_16/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_16/buf_output[0] ) );
  NAND3_X1 U3829 ( .A1(\SB4_9/i0_0 ), .A2(\SB4_9/i3[0] ), .A3(\SB4_9/i1_7 ), 
        .ZN(n1068) );
  BUF_X4 U3830 ( .I(\SB2_3_2/buf_output[5] ), .Z(\RI5[3][179] ) );
  NAND3_X2 U3831 ( .A1(\SB3_12/i1_5 ), .A2(\SB3_12/i0_0 ), .A3(\SB3_12/i0_4 ), 
        .ZN(n1069) );
  NAND3_X1 U3835 ( .A1(\SB2_3_7/i0_4 ), .A2(\SB2_3_7/i1_7 ), .A3(
        \SB2_3_7/i0[8] ), .ZN(\SB2_3_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U3837 ( .A1(\SB2_3_7/i0[7] ), .A2(\SB2_3_7/i0[6] ), .A3(
        \SB2_3_7/i0[8] ), .ZN(n2274) );
  XOR2_X1 U3840 ( .A1(\MC_ARK_ARC_1_4/temp4[81] ), .A2(n1071), .Z(
        \MC_ARK_ARC_1_4/temp6[81] ) );
  XOR2_X1 U3841 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[183] ), .A2(\RI5[4][147] ), 
        .Z(n1071) );
  XOR2_X1 U3846 ( .A1(\MC_ARK_ARC_1_1/temp6[186] ), .A2(n1073), .Z(
        \MC_ARK_ARC_1_1/buf_output[186] ) );
  XOR2_X1 U3847 ( .A1(\MC_ARK_ARC_1_1/temp1[186] ), .A2(
        \MC_ARK_ARC_1_1/temp2[186] ), .Z(n1073) );
  NAND4_X2 U3853 ( .A1(\SB1_0_8/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_8/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_8/Component_Function_4/NAND4_in[3] ), .A4(n1076), .ZN(
        \SB1_0_8/buf_output[4] ) );
  XOR2_X1 U3858 ( .A1(\RI5[3][108] ), .A2(\RI5[3][114] ), .Z(n1077) );
  XOR2_X1 U3860 ( .A1(\RI5[3][51] ), .A2(\RI5[3][87] ), .Z(n1078) );
  XOR2_X1 U3862 ( .A1(\MC_ARK_ARC_1_3/temp1[115] ), .A2(n1079), .Z(
        \MC_ARK_ARC_1_3/temp5[115] ) );
  XOR2_X1 U3863 ( .A1(\RI5[3][85] ), .A2(\RI5[3][61] ), .Z(n1079) );
  NAND3_X1 U3865 ( .A1(\SB3_12/i0[8] ), .A2(\RI1[5][119] ), .A3(\SB3_12/i1_7 ), 
        .ZN(\SB3_12/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U3869 ( .A1(n1083), .A2(\MC_ARK_ARC_1_3/temp5[179] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[179] ) );
  XOR2_X1 U3870 ( .A1(\MC_ARK_ARC_1_3/temp4[179] ), .A2(
        \MC_ARK_ARC_1_3/temp3[179] ), .Z(n1083) );
  NAND3_X1 U3873 ( .A1(\SB2_4_25/i0_0 ), .A2(\SB2_4_25/i3[0] ), .A3(
        \SB2_4_25/i1_7 ), .ZN(\SB2_4_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3884 ( .A1(\SB4_10/i0[6] ), .A2(\SB4_10/i0[9] ), .A3(\SB4_10/i1_5 ), .ZN(n1087) );
  XOR2_X1 U3887 ( .A1(\MC_ARK_ARC_1_2/temp3[68] ), .A2(
        \MC_ARK_ARC_1_2/temp4[68] ), .Z(n1089) );
  XOR2_X1 U3888 ( .A1(\RI5[4][81] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[75] ), 
        .Z(n2910) );
  NAND4_X2 U3889 ( .A1(n1593), .A2(\SB1_3_17/Component_Function_5/NAND4_in[1] ), .A3(\SB1_3_17/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_3_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_17/buf_output[5] ) );
  NAND3_X2 U3897 ( .A1(\SB2_2_18/i0[6] ), .A2(\SB2_2_18/i0_3 ), .A3(
        \SB2_2_18/i1[9] ), .ZN(n1095) );
  NAND4_X2 U3902 ( .A1(\SB2_0_18/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_18/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_0_18/Component_Function_0/NAND4_in[2] ), .A4(n1096), .ZN(
        \SB2_0_18/buf_output[0] ) );
  NAND3_X1 U3903 ( .A1(\SB2_0_18/i0_3 ), .A2(\SB2_0_18/i0_0 ), .A3(
        \SB2_0_18/i0[7] ), .ZN(n1096) );
  NAND3_X1 U3905 ( .A1(n6612), .A2(\SB2_1_29/i0[8] ), .A3(\SB2_1_29/i0[6] ), 
        .ZN(\SB2_1_29/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3913 ( .A1(\SB4_25/i0_3 ), .A2(\SB4_25/i0[8] ), .A3(\SB4_25/i1_7 ), 
        .ZN(\SB4_25/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U3918 ( .A1(\SB1_3_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_7/Component_Function_3/NAND4_in[1] ), .A3(n2544), .A4(n2884), 
        .ZN(\SB1_3_7/buf_output[3] ) );
  NAND4_X2 U3919 ( .A1(\SB3_14/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_14/Component_Function_0/NAND4_in[0] ), .A4(n1103), .ZN(
        \SB3_14/buf_output[0] ) );
  NAND3_X1 U3920 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i0_3 ), .A3(\SB3_14/i0[7] ), 
        .ZN(n1103) );
  BUF_X4 U3924 ( .I(\SB2_4_13/buf_output[3] ), .Z(\RI5[4][123] ) );
  NAND3_X1 U3930 ( .A1(\SB4_13/i0[6] ), .A2(n1498), .A3(\SB4_13/i0[7] ), .ZN(
        \SB4_13/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U3931 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i0_0 ), .A3(
        \SB2_3_20/i0[6] ), .ZN(n2174) );
  NAND3_X2 U3934 ( .A1(\SB1_3_23/i0[10] ), .A2(\SB1_3_23/i1[9] ), .A3(
        \SB1_3_23/i1_7 ), .ZN(n1109) );
  XOR2_X1 U3937 ( .A1(\RI5[4][28] ), .A2(\RI5[4][52] ), .Z(n1111) );
  NAND4_X2 U3938 ( .A1(\SB3_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_0/NAND4_in[0] ), .A4(n1112), .ZN(
        \SB3_21/buf_output[0] ) );
  NAND4_X2 U3947 ( .A1(\SB1_4_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_4_2/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_4_2/Component_Function_2/NAND4_in[1] ), .A4(n1115), .ZN(
        \SB1_4_2/buf_output[2] ) );
  NAND3_X1 U3948 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i1[9] ), .A3(
        \SB1_0_8/i0[6] ), .ZN(n1116) );
  NAND3_X2 U3951 ( .A1(\SB1_1_17/i0[9] ), .A2(\SB1_1_17/i0_3 ), .A3(
        \SB1_1_17/i0[8] ), .ZN(n1192) );
  XOR2_X1 U3953 ( .A1(\RI5[4][30] ), .A2(\RI5[4][36] ), .Z(
        \MC_ARK_ARC_1_4/temp1[36] ) );
  XOR2_X1 U3954 ( .A1(n1120), .A2(n193), .Z(Ciphertext[31]) );
  XOR2_X1 U3955 ( .A1(n1121), .A2(\MC_ARK_ARC_1_4/temp6[60] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[60] ) );
  XOR2_X1 U3956 ( .A1(\MC_ARK_ARC_1_4/temp2[60] ), .A2(
        \MC_ARK_ARC_1_4/temp1[60] ), .Z(n1121) );
  XOR2_X1 U3957 ( .A1(\MC_ARK_ARC_1_0/temp1[181] ), .A2(
        \MC_ARK_ARC_1_0/temp2[181] ), .Z(\MC_ARK_ARC_1_0/temp5[181] ) );
  XOR2_X1 U3959 ( .A1(n1122), .A2(n1123), .Z(\MC_ARK_ARC_1_0/buf_output[136] )
         );
  XOR2_X1 U3960 ( .A1(\MC_ARK_ARC_1_0/temp3[136] ), .A2(
        \MC_ARK_ARC_1_0/temp1[136] ), .Z(n1122) );
  XOR2_X1 U3961 ( .A1(\MC_ARK_ARC_1_0/temp2[136] ), .A2(
        \MC_ARK_ARC_1_0/temp4[136] ), .Z(n1123) );
  NAND3_X1 U3963 ( .A1(\SB3_24/i0[10] ), .A2(\SB3_24/i1[9] ), .A3(
        \SB3_24/i1_5 ), .ZN(\SB3_24/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U3968 ( .A1(\SB2_2_27/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_27/Component_Function_0/NAND4_in[0] ), .A4(n1125), .ZN(
        \SB2_2_27/buf_output[0] ) );
  XOR2_X1 U3971 ( .A1(\RI5[1][135] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[141] ), 
        .Z(n1126) );
  NAND3_X2 U3972 ( .A1(\RI3[0][77] ), .A2(\SB2_0_19/i0_0 ), .A3(
        \SB2_0_19/i0[7] ), .ZN(n1871) );
  XOR2_X1 U3976 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[177] ), .A2(\RI5[4][153] ), 
        .Z(n1128) );
  NAND3_X2 U3998 ( .A1(\SB1_3_5/i0[9] ), .A2(\SB1_3_5/i0_4 ), .A3(
        \SB1_3_5/i0[6] ), .ZN(n2043) );
  NAND4_X1 U4000 ( .A1(\SB2_0_27/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_0_27/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_27/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_27/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_27/buf_output[4] ) );
  NAND4_X2 U4001 ( .A1(\SB2_4_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_6/Component_Function_3/NAND4_in[2] ), .A3(n1938), .A4(
        \SB2_4_6/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_4_6/buf_output[3] ) );
  NAND4_X2 U4002 ( .A1(\SB1_0_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_0/Component_Function_5/NAND4_in[1] ), .A3(n2810), .A4(
        \SB1_0_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_0/buf_output[5] ) );
  XOR2_X1 U4011 ( .A1(\RI5[2][62] ), .A2(\RI5[2][26] ), .Z(
        \MC_ARK_ARC_1_2/temp3[152] ) );
  XOR2_X1 U4013 ( .A1(n2253), .A2(\MC_ARK_ARC_1_3/temp6[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[3] ) );
  NAND4_X2 U4014 ( .A1(n2024), .A2(\SB1_3_24/Component_Function_4/NAND4_in[0] ), .A3(\SB1_3_24/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_3_24/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_24/buf_output[4] ) );
  NAND3_X1 U4015 ( .A1(\SB2_3_23/i0_4 ), .A2(\SB2_3_23/i1_7 ), .A3(
        \SB2_3_23/i0[8] ), .ZN(\SB2_3_23/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U4016 ( .A1(\SB2_1_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_27/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_1_27/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_1_27/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_1_27/buf_output[4] ) );
  NAND3_X2 U4029 ( .A1(\SB2_1_16/i0[10] ), .A2(\SB2_1_16/i0[6] ), .A3(
        \SB2_1_16/i0_0 ), .ZN(n1137) );
  XOR2_X1 U4033 ( .A1(\RI5[3][38] ), .A2(\RI5[3][74] ), .Z(
        \MC_ARK_ARC_1_3/temp3[164] ) );
  NAND3_X1 U4035 ( .A1(\SB4_24/i0_0 ), .A2(\SB4_24/i0[7] ), .A3(\SB4_24/i0_3 ), 
        .ZN(\SB4_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U4044 ( .A1(\SB1_4_3/i0_3 ), .A2(\SB1_4_3/i1[9] ), .A3(
        \SB1_4_3/i0_4 ), .ZN(n1142) );
  NAND3_X2 U4046 ( .A1(\SB2_2_2/i0_4 ), .A2(\SB2_2_2/i0_3 ), .A3(n6267), .ZN(
        n1143) );
  NAND4_X2 U4047 ( .A1(\SB2_3_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_21/Component_Function_4/NAND4_in[2] ), .A4(n1144), .ZN(
        \SB2_3_21/buf_output[4] ) );
  XOR2_X1 U4050 ( .A1(\MC_ARK_ARC_1_3/temp5[104] ), .A2(n1841), .Z(
        \MC_ARK_ARC_1_3/buf_output[104] ) );
  NAND3_X1 U4053 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i0[9] ), .A3(\SB4_10/i0[8] ), .ZN(n1146) );
  NAND4_X2 U4056 ( .A1(\SB1_0_0/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_0/Component_Function_1/NAND4_in[2] ), .A3(n2170), .A4(
        \SB1_0_0/Component_Function_1/NAND4_in[1] ), .ZN(\RI3[0][19] ) );
  XOR2_X1 U4059 ( .A1(\SB2_1_10/buf_output[4] ), .A2(\RI5[1][160] ), .Z(
        \MC_ARK_ARC_1_1/temp2[190] ) );
  NAND4_X2 U4060 ( .A1(\SB2_4_0/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_0/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_4_0/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_4_0/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_4_0/buf_output[0] ) );
  NAND4_X2 U4061 ( .A1(\SB2_1_10/Component_Function_4/NAND4_in[1] ), .A2(n2508), .A3(\SB2_1_10/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_1_10/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_10/buf_output[4] ) );
  NAND4_X2 U4066 ( .A1(\SB1_0_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_2/Component_Function_3/NAND4_in[1] ), .A3(n1920), .A4(
        \SB1_0_2/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][189] ) );
  XOR2_X1 U4082 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[129] ), .A2(\RI5[3][165] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[63] ) );
  INV_X1 U4084 ( .I(\SB1_3_17/buf_output[0] ), .ZN(\SB2_3_12/i3[0] ) );
  NAND4_X2 U4085 ( .A1(\SB1_3_17/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_17/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_3_17/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_17/buf_output[0] ) );
  XOR2_X1 U4088 ( .A1(\MC_ARK_ARC_1_1/temp5[133] ), .A2(n1155), .Z(
        \MC_ARK_ARC_1_1/buf_output[133] ) );
  XOR2_X1 U4089 ( .A1(\MC_ARK_ARC_1_1/temp3[133] ), .A2(
        \MC_ARK_ARC_1_1/temp4[133] ), .Z(n1155) );
  XOR2_X1 U4090 ( .A1(\MC_ARK_ARC_1_3/temp1[44] ), .A2(n1156), .Z(
        \MC_ARK_ARC_1_3/temp5[44] ) );
  XOR2_X1 U4091 ( .A1(\RI5[3][14] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[182] ), 
        .Z(n1156) );
  XOR2_X1 U4094 ( .A1(\MC_ARK_ARC_1_3/temp4[44] ), .A2(n1157), .Z(n2077) );
  XOR2_X1 U4095 ( .A1(\SB2_3_10/buf_output[2] ), .A2(\RI5[3][110] ), .Z(n1157)
         );
  INV_X2 U4096 ( .I(n1158), .ZN(\RI1[5][179] ) );
  XNOR2_X1 U4097 ( .A1(\MC_ARK_ARC_1_4/temp5[179] ), .A2(n3145), .ZN(n1158) );
  INV_X2 U4102 ( .I(\MC_ARK_ARC_1_3/buf_output[44] ), .ZN(\SB1_4_24/i1[9] ) );
  NAND3_X1 U4105 ( .A1(\SB2_0_28/i0[6] ), .A2(\SB2_0_28/i1_5 ), .A3(
        \SB2_0_28/i0[9] ), .ZN(\SB2_0_28/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U4110 ( .A1(\RI5[0][9] ), .A2(\RI5[0][45] ), .Z(
        \MC_ARK_ARC_1_0/temp3[135] ) );
  XOR2_X1 U4111 ( .A1(n1179), .A2(\MC_ARK_ARC_1_3/temp4[132] ), .Z(
        \MC_ARK_ARC_1_3/temp6[132] ) );
  XOR2_X1 U4112 ( .A1(\MC_ARK_ARC_1_0/temp2[145] ), .A2(
        \MC_ARK_ARC_1_0/temp1[145] ), .Z(\MC_ARK_ARC_1_0/temp5[145] ) );
  XOR2_X1 U4115 ( .A1(\RI5[2][39] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[45] ) );
  XOR2_X1 U4118 ( .A1(\RI5[2][148] ), .A2(\RI5[2][154] ), .Z(n1165) );
  NAND3_X1 U4119 ( .A1(\SB1_0_14/i0[9] ), .A2(\SB1_0_14/i0[8] ), .A3(
        \SB1_0_14/i0_3 ), .ZN(n1166) );
  XOR2_X1 U4120 ( .A1(\MC_ARK_ARC_1_1/temp6[138] ), .A2(n1167), .Z(
        \MC_ARK_ARC_1_1/buf_output[138] ) );
  XOR2_X1 U4121 ( .A1(\MC_ARK_ARC_1_1/temp1[138] ), .A2(n1369), .Z(n1167) );
  NOR2_X2 U4124 ( .A1(n2693), .A2(n1170), .ZN(\SB2_0_9/i3[0] ) );
  NAND3_X2 U4127 ( .A1(\SB2_2_20/i1[9] ), .A2(\SB2_2_20/i1_7 ), .A3(
        \SB2_2_20/i0[10] ), .ZN(\SB2_2_20/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U4128 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i0_4 ), .A3(
        \SB2_1_14/i0[10] ), .ZN(n1171) );
  NAND3_X1 U4131 ( .A1(n600), .A2(\SB2_2_23/i0[8] ), .A3(\SB2_2_23/i1_7 ), 
        .ZN(\SB2_2_23/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U4136 ( .A1(\SB2_0_24/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_0_24/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_0_24/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_0_24/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_0_24/buf_output[1] ) );
  XOR2_X1 U4145 ( .A1(\RI5[1][61] ), .A2(\RI5[1][97] ), .Z(
        \MC_ARK_ARC_1_1/temp3[187] ) );
  NAND4_X2 U4154 ( .A1(\SB1_3_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_8/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_8/Component_Function_3/NAND4_in[3] ), .A4(n1184), .ZN(
        \SB1_3_8/buf_output[3] ) );
  INV_X2 U4161 ( .I(\SB1_2_0/buf_output[5] ), .ZN(\SB2_2_0/i1_5 ) );
  XOR2_X1 U4162 ( .A1(n1189), .A2(n1188), .Z(\MC_ARK_ARC_1_3/buf_output[118] )
         );
  XOR2_X1 U4163 ( .A1(\MC_ARK_ARC_1_3/temp1[118] ), .A2(
        \MC_ARK_ARC_1_3/temp4[118] ), .Z(n1188) );
  XOR2_X1 U4168 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[43] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[19] ), .Z(n1191) );
  NAND3_X1 U4183 ( .A1(\SB4_28/i0_0 ), .A2(\SB4_28/i1_7 ), .A3(\SB4_28/i3[0] ), 
        .ZN(n1199) );
  NAND3_X1 U4187 ( .A1(n3983), .A2(\SB2_4_30/i0[8] ), .A3(\SB2_4_30/i1_5 ), 
        .ZN(\SB2_4_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U4202 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i0[8] ), .A3(
        \SB1_2_5/i0[9] ), .ZN(\SB1_2_5/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U4204 ( .A1(\RI5[0][87] ), .A2(\RI5[0][93] ), .Z(n1200) );
  XOR2_X1 U4207 ( .A1(\MC_ARK_ARC_1_4/temp4[25] ), .A2(
        \MC_ARK_ARC_1_4/temp3[25] ), .Z(n2528) );
  XOR2_X1 U4211 ( .A1(\MC_ARK_ARC_1_0/temp3[149] ), .A2(n583), .Z(n1203) );
  NAND3_X2 U4214 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i1[9] ), .A3(
        \SB1_0_22/i0_4 ), .ZN(n2074) );
  XOR2_X1 U4215 ( .A1(n1205), .A2(\MC_ARK_ARC_1_3/temp4[174] ), .Z(
        \MC_ARK_ARC_1_3/temp6[174] ) );
  NAND3_X1 U4221 ( .A1(\SB1_2_5/i0[6] ), .A2(\SB1_2_5/i0[8] ), .A3(
        \SB1_2_5/i0[7] ), .ZN(\SB1_2_5/Component_Function_0/NAND4_in[1] ) );
  BUF_X4 U4224 ( .I(\MC_ARK_ARC_1_3/buf_output[125] ), .Z(\SB1_4_11/i0_3 ) );
  NAND3_X2 U4229 ( .A1(\SB2_0_0/i0_3 ), .A2(\SB2_0_0/i1_7 ), .A3(n4003), .ZN(
        \SB2_0_0/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U4231 ( .A1(n1209), .A2(\MC_ARK_ARC_1_0/temp6[63] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[63] ) );
  BUF_X4 U4234 ( .I(\SB2_2_8/buf_output[3] ), .Z(\RI5[2][153] ) );
  NAND3_X1 U4242 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i0[9] ), .A3(n1498), .ZN(
        n1214) );
  NAND3_X2 U4246 ( .A1(\SB2_1_20/i0_3 ), .A2(\SB2_1_20/i0[9] ), .A3(
        \SB2_1_20/i0[8] ), .ZN(\SB2_1_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U4250 ( .A1(\SB2_1_2/i0[7] ), .A2(\SB2_1_2/i0[8] ), .A3(
        \SB2_1_2/i0[6] ), .ZN(\SB2_1_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U4256 ( .A1(\SB1_4_30/i1_5 ), .A2(\SB1_4_30/i0_4 ), .A3(
        \SB1_4_30/i1[9] ), .ZN(\SB1_4_30/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U4267 ( .A1(n1414), .A2(n1222), .Z(\MC_ARK_ARC_1_4/temp5[59] ) );
  XOR2_X1 U4268 ( .A1(\RI5[4][59] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[53] ), 
        .Z(n1222) );
  XOR2_X1 U4269 ( .A1(\MC_ARK_ARC_1_3/temp1[69] ), .A2(n1223), .Z(
        \MC_ARK_ARC_1_3/temp5[69] ) );
  NAND4_X2 U4279 ( .A1(\SB2_0_12/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_12/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_12/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_0_12/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_12/buf_output[3] ) );
  BUF_X4 U4282 ( .I(\SB2_4_7/buf_output[2] ), .Z(\RI5[4][164] ) );
  NAND3_X1 U4285 ( .A1(n6265), .A2(\SB2_4_30/i0[8] ), .A3(\SB2_4_30/i0[6] ), 
        .ZN(\SB2_4_30/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U4287 ( .A1(n1230), .A2(n82), .Z(Ciphertext[36]) );
  NAND4_X2 U4288 ( .A1(\SB4_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_25/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_25/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_25/Component_Function_0/NAND4_in[0] ), .ZN(n1230) );
  NAND3_X1 U4299 ( .A1(\SB1_3_6/i0_3 ), .A2(\SB1_3_6/i0[8] ), .A3(
        \SB1_3_6/i1_7 ), .ZN(\SB1_3_6/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U4302 ( .A1(\SB2_1_29/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_29/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_29/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_29/buf_output[0] ) );
  XOR2_X1 U4303 ( .A1(n1236), .A2(n1235), .Z(\MC_ARK_ARC_1_3/temp6[119] ) );
  XOR2_X1 U4304 ( .A1(\RI5[3][185] ), .A2(n87), .Z(n1235) );
  NAND3_X1 U4306 ( .A1(\SB4_26/i0[10] ), .A2(n573), .A3(\SB4_26/i1_7 ), .ZN(
        n1237) );
  XOR2_X1 U4311 ( .A1(\RI5[3][66] ), .A2(\RI5[3][90] ), .Z(
        \MC_ARK_ARC_1_3/temp2[120] ) );
  NAND3_X1 U4316 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i0[9] ), .A3(
        \SB3_23/i0[10] ), .ZN(n1242) );
  NAND4_X2 U4317 ( .A1(\SB2_0_7/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_7/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_0_7/Component_Function_0/NAND4_in[2] ), .A4(n1243), .ZN(
        \SB2_0_7/buf_output[0] ) );
  NAND3_X1 U4324 ( .A1(\SB2_4_23/i0[10] ), .A2(\SB2_4_23/i0_3 ), .A3(
        \SB2_4_23/i0[9] ), .ZN(n1246) );
  NAND4_X2 U4327 ( .A1(\SB1_0_0/Component_Function_4/NAND4_in[1] ), .A2(n2811), 
        .A3(\SB1_0_0/Component_Function_4/NAND4_in[0] ), .A4(n1248), .ZN(
        \SB1_0_0/buf_output[4] ) );
  XOR2_X1 U4335 ( .A1(\RI5[0][74] ), .A2(\RI5[0][98] ), .Z(
        \MC_ARK_ARC_1_0/temp2[128] ) );
  XOR2_X1 U4339 ( .A1(n1253), .A2(\MC_ARK_ARC_1_1/temp1[155] ), .Z(
        \MC_ARK_ARC_1_1/temp5[155] ) );
  XOR2_X1 U4340 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[125] ), .A2(\RI5[1][101] ), 
        .Z(n1253) );
  NAND3_X1 U4341 ( .A1(\SB4_21/i0[9] ), .A2(\SB4_21/i0[6] ), .A3(\SB4_21/i1_5 ), .ZN(n1254) );
  NAND4_X2 U4344 ( .A1(\SB1_4_3/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_4_3/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_4_3/Component_Function_4/NAND4_in[2] ), .A4(n1256), .ZN(
        \SB1_4_3/buf_output[4] ) );
  NAND3_X1 U4345 ( .A1(\SB1_4_3/i1[9] ), .A2(\SB1_4_3/i1_5 ), .A3(
        \SB1_4_3/i0_4 ), .ZN(n1256) );
  NAND3_X1 U4350 ( .A1(\SB4_12/i0_3 ), .A2(\SB4_12/i0[6] ), .A3(\SB4_12/i1[9] ), .ZN(\SB4_12/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U4351 ( .I(\SB2_2_28/buf_output[0] ), .Z(\RI5[2][48] ) );
  BUF_X4 U4352 ( .I(\SB2_4_5/buf_output[1] ), .Z(\RI5[4][181] ) );
  NAND3_X1 U4358 ( .A1(\SB4_27/i0[10] ), .A2(\SB4_27/i0[6] ), .A3(
        \SB4_27/i0_3 ), .ZN(n1403) );
  XOR2_X1 U4361 ( .A1(n1260), .A2(n112), .Z(Ciphertext[110]) );
  NAND3_X2 U4366 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i1[9] ), .A3(\SB3_23/i0_4 ), 
        .ZN(\SB3_23/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U4379 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[109] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_3/temp1[115] )
         );
  NAND3_X2 U4381 ( .A1(\SB2_2_12/i0_0 ), .A2(\SB2_2_12/i0_4 ), .A3(
        \SB2_2_12/i1_5 ), .ZN(n1266) );
  NAND3_X2 U4388 ( .A1(\SB2_1_27/i0_3 ), .A2(\RI3[1][26] ), .A3(
        \SB2_1_27/i0_4 ), .ZN(n1680) );
  NAND3_X2 U4391 ( .A1(\SB1_2_16/i0[10] ), .A2(\SB1_2_16/i1[9] ), .A3(
        \SB1_2_16/i1_7 ), .ZN(n1270) );
  NAND3_X2 U4393 ( .A1(\SB2_2_22/i0[10] ), .A2(\SB2_2_22/i1[9] ), .A3(
        \SB2_2_22/i1_7 ), .ZN(\SB2_2_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U4397 ( .A1(\SB1_4_6/i0[10] ), .A2(\SB1_4_6/i0_0 ), .A3(
        \SB1_4_6/i0[6] ), .ZN(\SB1_4_6/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U4402 ( .A1(n1274), .A2(\MC_ARK_ARC_1_2/temp1[34] ), .Z(
        \MC_ARK_ARC_1_2/temp5[34] ) );
  XOR2_X1 U4403 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[172] ), .A2(\RI5[2][4] ), 
        .Z(n1274) );
  XOR2_X1 U4418 ( .A1(n1282), .A2(\MC_ARK_ARC_1_0/temp5[148] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[148] ) );
  XOR2_X1 U4419 ( .A1(\MC_ARK_ARC_1_0/temp3[148] ), .A2(
        \MC_ARK_ARC_1_0/temp4[148] ), .Z(n1282) );
  INV_X1 U4420 ( .I(\SB1_4_25/buf_output[0] ), .ZN(\SB2_4_20/i3[0] ) );
  XOR2_X1 U4426 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[96] ), .A2(\RI5[3][120] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[150] ) );
  NAND3_X1 U4431 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i1_7 ), .A3(\SB4_12/i0[8] ), 
        .ZN(n1287) );
  NAND3_X2 U4434 ( .A1(\RI3[0][71] ), .A2(\SB2_0_20/i0_0 ), .A3(\RI3[0][70] ), 
        .ZN(\SB2_0_20/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 U4435 ( .I(\SB2_2_7/buf_output[1] ), .Z(\RI5[2][169] ) );
  NAND3_X1 U4436 ( .A1(\SB2_3_5/i0[7] ), .A2(\SB2_3_5/i0_0 ), .A3(
        \SB2_3_5/i0_3 ), .ZN(\SB2_3_5/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U4439 ( .A1(\SB2_3_10/Component_Function_5/NAND4_in[2] ), .A2(n2792), .A3(n1291), .A4(\SB2_3_10/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_10/buf_output[5] ) );
  INV_X2 U4442 ( .I(\RI3[0][91] ), .ZN(\SB2_0_16/i1_7 ) );
  NAND4_X2 U4443 ( .A1(\SB1_4_26/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_4_26/Component_Function_3/NAND4_in[0] ), .A3(n1795), .A4(
        \SB1_4_26/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_4_26/buf_output[3] ) );
  XOR2_X1 U4444 ( .A1(\MC_ARK_ARC_1_4/temp6[57] ), .A2(
        \MC_ARK_ARC_1_4/temp5[57] ), .Z(\MC_ARK_ARC_1_4/buf_output[57] ) );
  NAND3_X1 U4448 ( .A1(\SB1_0_8/i0_0 ), .A2(\SB1_0_8/i1_5 ), .A3(n364), .ZN(
        n1294) );
  NAND3_X1 U4450 ( .A1(\SB4_4/i0_0 ), .A2(\SB4_4/i1_5 ), .A3(\SB4_4/i0_4 ), 
        .ZN(n1295) );
  XOR2_X1 U4452 ( .A1(\RI5[2][57] ), .A2(\RI5[2][93] ), .Z(n1296) );
  NAND3_X2 U4455 ( .A1(\SB2_0_20/i0[8] ), .A2(\RI3[0][71] ), .A3(n5264), .ZN(
        \SB2_0_20/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U4465 ( .A1(\RI5[4][115] ), .A2(\RI5[4][109] ), .Z(
        \MC_ARK_ARC_1_4/temp1[115] ) );
  AND2_X1 U4467 ( .A1(\SB2_4_17/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_4_17/Component_Function_1/NAND4_in[1] ), .Z(n1303) );
  NAND4_X2 U4476 ( .A1(n1660), .A2(n1659), .A3(
        \SB2_1_18/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_1_18/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_18/buf_output[0] ) );
  BUF_X4 U4478 ( .I(\MC_ARK_ARC_1_0/buf_output[137] ), .Z(\SB1_1_9/i0_3 ) );
  XOR2_X1 U4482 ( .A1(n1312), .A2(n1313), .Z(\MC_ARK_ARC_1_0/temp5[149] ) );
  XOR2_X1 U4483 ( .A1(\RI5[0][143] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[149] ), 
        .Z(n1312) );
  XOR2_X1 U4484 ( .A1(\RI5[0][95] ), .A2(\RI5[0][119] ), .Z(n1313) );
  XOR2_X1 U4487 ( .A1(\MC_ARK_ARC_1_3/temp6[19] ), .A2(n1315), .Z(
        \MC_ARK_ARC_1_3/buf_output[19] ) );
  NAND2_X1 U4491 ( .A1(\SB1_0_17/Component_Function_4/NAND4_in[0] ), .A2(n1318), .ZN(n1317) );
  NAND2_X1 U4492 ( .A1(\SB1_0_17/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_17/Component_Function_4/NAND4_in[1] ), .ZN(n1319) );
  XOR2_X1 U4494 ( .A1(\MC_ARK_ARC_1_0/temp3[187] ), .A2(
        \MC_ARK_ARC_1_0/temp4[187] ), .Z(\MC_ARK_ARC_1_0/temp6[187] ) );
  NAND4_X2 U4496 ( .A1(\SB1_1_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_18/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_1_18/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_1_18/buf_output[4] ) );
  NAND4_X2 U4497 ( .A1(\SB1_1_15/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_15/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_15/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_1_15/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_1_15/buf_output[4] ) );
  XOR2_X1 U4498 ( .A1(\MC_ARK_ARC_1_1/temp3[16] ), .A2(
        \MC_ARK_ARC_1_1/temp4[16] ), .Z(\MC_ARK_ARC_1_1/temp6[16] ) );
  XOR2_X1 U4503 ( .A1(\RI5[3][163] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[187] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[25] ) );
  NAND4_X2 U4509 ( .A1(\SB1_0_12/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_12/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_12/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_0_12/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_0_12/buf_output[4] ) );
  INV_X2 U4512 ( .I(\SB1_3_21/buf_output[3] ), .ZN(\SB2_3_19/i0[8] ) );
  NAND3_X1 U4513 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i1[9] ), .A3(\SB4_5/i1_7 ), 
        .ZN(n1324) );
  BUF_X4 U4514 ( .I(\SB1_3_10/buf_output[5] ), .Z(\SB2_3_10/i0_3 ) );
  NAND3_X1 U4518 ( .A1(\SB2_4_3/i0_3 ), .A2(\SB2_4_3/i0[10] ), .A3(
        \SB2_4_3/i0_4 ), .ZN(\SB2_4_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4525 ( .A1(\SB3_9/i0[6] ), .A2(\MC_ARK_ARC_1_4/buf_output[132] ), 
        .A3(\SB3_9/i0_4 ), .ZN(n1327) );
  BUF_X4 U4526 ( .I(\SB2_2_8/buf_output[0] ), .Z(\RI5[2][168] ) );
  NAND3_X1 U4529 ( .A1(\SB2_2_4/i0[6] ), .A2(\SB2_2_4/i0[9] ), .A3(
        \SB2_2_4/i1_5 ), .ZN(\SB2_2_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4533 ( .A1(\SB2_4_6/i0_0 ), .A2(\SB2_4_6/i0[9] ), .A3(
        \SB2_4_6/i0[8] ), .ZN(\SB2_4_6/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U4538 ( .A1(\SB1_0_7/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_7/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_7/Component_Function_4/NAND4_in[3] ), .A4(n1333), .ZN(
        \RI3[0][154] ) );
  NAND3_X1 U4541 ( .A1(\SB1_0_31/i0_4 ), .A2(\SB1_0_31/i0_0 ), .A3(
        \SB1_0_31/i0_3 ), .ZN(\SB1_0_31/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U4542 ( .A1(\SB1_2_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_23/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_2_23/Component_Function_3/NAND4_in[1] ), .A4(n1335), .ZN(
        \SB1_2_23/buf_output[3] ) );
  NAND3_X1 U4546 ( .A1(\SB2_0_29/i0[10] ), .A2(\SB2_0_29/i0_0 ), .A3(
        \SB2_0_29/i0[6] ), .ZN(\SB2_0_29/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U4547 ( .A1(n1729), .A2(n2771), .Z(\MC_ARK_ARC_1_0/buf_output[90] )
         );
  NAND3_X1 U4559 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i0[10] ), .A3(
        \SB1_0_22/i0_4 ), .ZN(\SB1_0_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4560 ( .A1(\SB1_1_30/i1_5 ), .A2(\SB1_1_30/i1[9] ), .A3(
        \SB1_1_30/i0_4 ), .ZN(n2311) );
  XOR2_X1 U4566 ( .A1(\RI5[1][129] ), .A2(\RI5[1][105] ), .Z(
        \MC_ARK_ARC_1_1/temp2[159] ) );
  XOR2_X1 U4571 ( .A1(\MC_ARK_ARC_1_1/temp5[171] ), .A2(n1348), .Z(
        \MC_ARK_ARC_1_1/buf_output[171] ) );
  XOR2_X1 U4587 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[144] ), .A2(\RI5[3][180] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[78] ) );
  XOR2_X1 U4605 ( .A1(\MC_ARK_ARC_1_2/temp2[171] ), .A2(n1363), .Z(
        \MC_ARK_ARC_1_2/temp5[171] ) );
  XOR2_X1 U4606 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[171] ), .A2(\RI5[2][165] ), 
        .Z(n1363) );
  INV_X2 U4608 ( .I(\SB1_0_10/buf_output[2] ), .ZN(\SB2_0_7/i1[9] ) );
  AND2_X1 U4610 ( .A1(n1913), .A2(\SB1_0_10/Component_Function_2/NAND4_in[2] ), 
        .Z(n1364) );
  XOR2_X1 U4612 ( .A1(\RI5[4][65] ), .A2(\RI5[4][101] ), .Z(
        \MC_ARK_ARC_1_4/temp3[191] ) );
  XOR2_X1 U4613 ( .A1(\MC_ARK_ARC_1_0/temp6[36] ), .A2(n1366), .Z(
        \MC_ARK_ARC_1_0/buf_output[36] ) );
  XOR2_X1 U4614 ( .A1(\MC_ARK_ARC_1_0/temp2[36] ), .A2(
        \MC_ARK_ARC_1_0/temp1[36] ), .Z(n1366) );
  XOR2_X1 U4619 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[84] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[108] ), .Z(n1369) );
  XOR2_X1 U4622 ( .A1(\MC_ARK_ARC_1_0/temp1[84] ), .A2(
        \MC_ARK_ARC_1_0/temp2[84] ), .Z(\MC_ARK_ARC_1_0/temp5[84] ) );
  XOR2_X1 U4624 ( .A1(\MC_ARK_ARC_1_0/temp3[143] ), .A2(
        \MC_ARK_ARC_1_0/temp4[143] ), .Z(\MC_ARK_ARC_1_0/temp6[143] ) );
  BUF_X4 U4625 ( .I(\SB2_3_0/buf_output[4] ), .Z(\RI5[3][4] ) );
  XOR2_X1 U4626 ( .A1(\MC_ARK_ARC_1_3/temp2[188] ), .A2(
        \MC_ARK_ARC_1_3/temp1[188] ), .Z(\MC_ARK_ARC_1_3/temp5[188] ) );
  BUF_X4 U4627 ( .I(\SB2_0_7/buf_output[3] ), .Z(\RI5[0][159] ) );
  NAND4_X2 U4629 ( .A1(\SB2_1_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_25/Component_Function_3/NAND4_in[2] ), .A4(n1372), .ZN(
        \SB2_1_25/buf_output[3] ) );
  BUF_X4 U4635 ( .I(\SB2_0_10/buf_output[5] ), .Z(\RI5[0][131] ) );
  NAND3_X1 U4637 ( .A1(\SB2_0_23/i0_0 ), .A2(\SB2_0_23/i0[9] ), .A3(
        \SB2_0_23/i0[8] ), .ZN(\SB2_0_23/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U4639 ( .A1(\SB1_2_10/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_10/Component_Function_0/NAND4_in[0] ), .A4(n1376), .ZN(
        \SB1_2_10/buf_output[0] ) );
  XOR2_X1 U4644 ( .A1(n2335), .A2(n1379), .Z(\MC_ARK_ARC_1_2/temp5[5] ) );
  XOR2_X1 U4645 ( .A1(\RI5[2][167] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[143] ), 
        .Z(n1379) );
  XOR2_X1 U4653 ( .A1(\MC_ARK_ARC_1_1/temp2[161] ), .A2(n1383), .Z(
        \MC_ARK_ARC_1_1/temp5[161] ) );
  XOR2_X1 U4654 ( .A1(\RI5[1][155] ), .A2(\RI5[1][161] ), .Z(n1383) );
  XOR2_X1 U4658 ( .A1(\RI5[4][33] ), .A2(\RI5[4][57] ), .Z(n1384) );
  XOR2_X1 U4668 ( .A1(n1390), .A2(\MC_ARK_ARC_1_1/temp6[148] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[148] ) );
  XOR2_X1 U4669 ( .A1(\MC_ARK_ARC_1_3/temp1[98] ), .A2(
        \MC_ARK_ARC_1_3/temp2[98] ), .Z(\MC_ARK_ARC_1_3/temp5[98] ) );
  BUF_X4 U4671 ( .I(\SB2_2_28/buf_output[1] ), .Z(\RI5[2][43] ) );
  XOR2_X1 U4674 ( .A1(n1393), .A2(n1392), .Z(n2762) );
  XOR2_X1 U4675 ( .A1(\RI5[3][120] ), .A2(n460), .Z(n1392) );
  XOR2_X1 U4676 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[156] ), .A2(\RI5[3][90] ), 
        .Z(n1393) );
  NAND3_X1 U4682 ( .A1(\SB4_30/i0_3 ), .A2(\SB4_30/i0_4 ), .A3(n3973), .ZN(
        \SB4_30/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U4684 ( .A1(\MC_ARK_ARC_1_2/temp1[30] ), .A2(
        \MC_ARK_ARC_1_2/temp2[30] ), .Z(\MC_ARK_ARC_1_2/temp5[30] ) );
  BUF_X2 U4685 ( .I(\SB3_24/buf_output[3] ), .Z(\SB4_22/i0[10] ) );
  XOR2_X1 U4686 ( .A1(\MC_ARK_ARC_1_0/temp6[54] ), .A2(
        \MC_ARK_ARC_1_0/temp5[54] ), .Z(\MC_ARK_ARC_1_0/buf_output[54] ) );
  XOR2_X1 U4703 ( .A1(\RI5[0][185] ), .A2(\RI5[0][191] ), .Z(n1399) );
  INV_X1 U4707 ( .I(\SB3_11/buf_output[5] ), .ZN(\SB4_11/i1_5 ) );
  NAND3_X1 U4710 ( .A1(\SB3_15/i0_4 ), .A2(\SB3_15/i1[9] ), .A3(\SB3_15/i1_5 ), 
        .ZN(\SB3_15/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U4711 ( .A1(\RI5[4][51] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[75] ), 
        .Z(n1401) );
  NAND3_X2 U4714 ( .A1(\SB1_4_25/i0_0 ), .A2(\SB1_4_25/i0[10] ), .A3(
        \SB1_4_25/i0[6] ), .ZN(\SB1_4_25/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U4720 ( .A1(n1407), .A2(\MC_ARK_ARC_1_4/temp6[100] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[100] ) );
  XOR2_X1 U4721 ( .A1(\MC_ARK_ARC_1_4/temp2[100] ), .A2(
        \MC_ARK_ARC_1_4/temp1[100] ), .Z(n1407) );
  XOR2_X1 U4726 ( .A1(\RI5[1][93] ), .A2(\RI5[1][129] ), .Z(
        \MC_ARK_ARC_1_1/temp3[27] ) );
  NAND3_X2 U4733 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0_4 ), .A3(
        \SB1_3_21/i0_0 ), .ZN(n1412) );
  XOR2_X1 U4737 ( .A1(\RI5[4][29] ), .A2(\RI5[4][5] ), .Z(n1414) );
  NAND3_X2 U4740 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0_4 ), .A3(
        \SB2_2_30/i1[9] ), .ZN(n1415) );
  XOR2_X1 U4743 ( .A1(\RI5[2][54] ), .A2(\RI5[2][48] ), .Z(
        \MC_ARK_ARC_1_2/temp1[54] ) );
  BUF_X4 U4744 ( .I(\MC_ARK_ARC_1_3/buf_output[89] ), .Z(\SB1_4_17/i0_3 ) );
  NAND2_X1 U4749 ( .A1(\SB1_4_22/i0[9] ), .A2(\SB1_4_22/i0[10] ), .ZN(
        \SB1_4_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 U4750 ( .A1(\SB2_3_26/i0[10] ), .A2(\SB2_3_26/i0_0 ), .A3(
        \SB2_3_26/i0[6] ), .ZN(n2006) );
  NAND4_X2 U4751 ( .A1(\SB2_1_22/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_22/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_22/Component_Function_4/NAND4_in[3] ), .A4(n1417), .ZN(
        \SB2_1_22/buf_output[4] ) );
  NAND4_X2 U4762 ( .A1(\SB2_0_23/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_23/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_0_23/Component_Function_0/NAND4_in[2] ), .A4(n1422), .ZN(
        \SB2_0_23/buf_output[0] ) );
  NAND3_X2 U4763 ( .A1(\SB2_0_23/i0[6] ), .A2(\SB2_0_23/i0[7] ), .A3(
        \SB2_0_23/i0[8] ), .ZN(n1422) );
  XOR2_X1 U4767 ( .A1(n2334), .A2(\MC_ARK_ARC_1_0/temp4[179] ), .Z(n1423) );
  NAND4_X2 U4768 ( .A1(\SB1_1_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_2/Component_Function_1/NAND4_in[3] ), .A3(n1711), .A4(n2856), 
        .ZN(\SB1_1_2/buf_output[1] ) );
  NAND3_X1 U4772 ( .A1(\SB2_4_20/i0[9] ), .A2(\SB2_4_20/i0_0 ), .A3(
        \SB2_4_20/i0[8] ), .ZN(n1426) );
  XOR2_X1 U4781 ( .A1(n1431), .A2(n1432), .Z(\MC_ARK_ARC_1_2/buf_output[117] )
         );
  XOR2_X1 U4783 ( .A1(\RI5[3][77] ), .A2(\RI5[3][41] ), .Z(n1433) );
  XOR2_X1 U4786 ( .A1(n2552), .A2(\MC_ARK_ARC_1_1/temp2[128] ), .Z(n1436) );
  XOR2_X1 U4806 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[108] ), .A2(\RI5[0][114] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[114] ) );
  NAND3_X1 U4815 ( .A1(\SB4_9/i0[9] ), .A2(\SB4_9/i0_3 ), .A3(n1499), .ZN(
        n1447) );
  XOR2_X1 U4820 ( .A1(\RI5[2][67] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[67] ) );
  NAND3_X1 U4821 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i1[9] ), .A3(\SB4_17/i0_4 ), 
        .ZN(\SB4_17/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U4822 ( .I(\SB2_3_14/buf_output[3] ), .Z(\RI5[3][117] ) );
  NAND4_X2 U4824 ( .A1(\SB2_0_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_22/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_22/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_22/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_22/buf_output[5] ) );
  INV_X2 U4825 ( .I(\SB1_2_21/buf_output[3] ), .ZN(\SB2_2_19/i0[8] ) );
  XOR2_X1 U4827 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[179] ), .A2(n59), .Z(n1448) );
  XOR2_X1 U4828 ( .A1(\RI5[2][17] ), .A2(\RI5[2][53] ), .Z(n1449) );
  NAND3_X1 U4830 ( .A1(n221), .A2(\SB1_0_31/i0[9] ), .A3(n1105), .ZN(n1450) );
  BUF_X4 U4835 ( .I(\MC_ARK_ARC_1_3/buf_output[152] ), .Z(\SB1_4_6/i0_0 ) );
  BUF_X4 U4837 ( .I(\SB1_2_2/buf_output[5] ), .Z(\SB2_2_2/i0_3 ) );
  NAND2_X2 U4838 ( .A1(\SB3_0/i0_0 ), .A2(\SB3_0/i3[0] ), .ZN(
        \SB3_0/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U4839 ( .I(\SB1_1_24/buf_output[5] ), .Z(\SB2_1_24/i0_3 ) );
  XOR2_X1 U4842 ( .A1(\RI5[3][146] ), .A2(\RI5[3][152] ), .Z(n2241) );
  INV_X2 U4843 ( .I(\MC_ARK_ARC_1_4/buf_output[86] ), .ZN(\SB3_17/i1[9] ) );
  XOR2_X1 U4853 ( .A1(\MC_ARK_ARC_1_3/temp6[92] ), .A2(
        \MC_ARK_ARC_1_3/temp5[92] ), .Z(\MC_ARK_ARC_1_3/buf_output[92] ) );
  NAND4_X2 U4863 ( .A1(\SB3_31/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_31/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_31/Component_Function_0/NAND4_in[0] ), .A4(
        \SB3_31/Component_Function_0/NAND4_in[1] ), .ZN(\SB3_31/buf_output[0] ) );
  NAND3_X2 U4872 ( .A1(\SB1_1_14/i0[9] ), .A2(\SB1_1_14/i0[8] ), .A3(
        \SB1_1_14/i0_3 ), .ZN(\SB1_1_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4874 ( .A1(\SB4_11/i0_4 ), .A2(\SB4_11/i1[9] ), .A3(\SB4_11/i1_5 ), 
        .ZN(n1461) );
  INV_X2 U4876 ( .I(\MC_ARK_ARC_1_0/buf_output[81] ), .ZN(\SB1_1_18/i0[8] ) );
  NAND4_X2 U4885 ( .A1(\SB1_0_26/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_26/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_0_26/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_0_26/Component_Function_0/NAND4_in[1] ), .ZN(\RI3[0][60] ) );
  XOR2_X1 U4889 ( .A1(\MC_ARK_ARC_1_2/temp5[16] ), .A2(n1466), .Z(
        \MC_ARK_ARC_1_2/buf_output[16] ) );
  XOR2_X1 U4890 ( .A1(\MC_ARK_ARC_1_2/temp4[16] ), .A2(
        \MC_ARK_ARC_1_2/temp3[16] ), .Z(n1466) );
  NAND4_X2 U4893 ( .A1(\SB1_0_26/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_26/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_26/Component_Function_3/NAND4_in[2] ), .A4(n1467), .ZN(
        \SB1_0_26/buf_output[3] ) );
  NAND3_X1 U4894 ( .A1(\SB1_0_26/i3[0] ), .A2(\SB1_0_26/i1_5 ), .A3(
        \SB1_0_26/i0[8] ), .ZN(n1467) );
  NOR2_X2 U4896 ( .A1(n1470), .A2(n1468), .ZN(n2611) );
  NAND3_X1 U4897 ( .A1(n261), .A2(\SB1_0_27/i0_0 ), .A3(\SB1_0_27/i0[8] ), 
        .ZN(n1469) );
  NAND3_X2 U4899 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \SB2_3_20/i0[6] ), .ZN(\SB2_3_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U4904 ( .A1(\SB3_17/i0_3 ), .A2(\SB3_17/i1[9] ), .A3(\SB3_17/i0[6] ), .ZN(\SB3_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U4915 ( .A1(\SB2_2_28/i0_0 ), .A2(\SB2_2_28/i1_5 ), .A3(
        \SB2_2_28/i0_4 ), .ZN(n3075) );
  INV_X2 U4918 ( .I(\SB1_1_0/buf_output[5] ), .ZN(\SB2_1_0/i1_5 ) );
  XOR2_X1 U4920 ( .A1(\MC_ARK_ARC_1_2/temp4[96] ), .A2(
        \MC_ARK_ARC_1_2/temp3[96] ), .Z(n1479) );
  INV_X2 U4925 ( .I(n1482), .ZN(\RI1[1][149] ) );
  XOR2_X1 U4932 ( .A1(n1487), .A2(\MC_ARK_ARC_1_0/temp6[147] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[147] ) );
  NAND4_X2 U4934 ( .A1(\SB1_0_15/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_15/Component_Function_1/NAND4_in[3] ), .A4(n1488), .ZN(
        \RI3[0][121] ) );
  INV_X2 U4951 ( .I(\SB1_4_12/buf_output[5] ), .ZN(\SB2_4_12/i1_5 ) );
  NAND3_X1 U4964 ( .A1(\SB1_0_30/i0[7] ), .A2(\SB1_0_30/i0_3 ), .A3(
        \SB1_0_30/i0_0 ), .ZN(\SB1_0_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4965 ( .A1(\SB1_0_30/i0[9] ), .A2(\SB1_0_30/i0[10] ), .A3(
        \SB1_0_30/i0_3 ), .ZN(\SB1_0_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4969 ( .A1(\SB3_6/i1_5 ), .A2(\SB3_6/i0[6] ), .A3(\SB3_6/i0[9] ), 
        .ZN(\SB3_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4972 ( .A1(\SB2_4_8/i0_3 ), .A2(\SB2_4_8/i1_7 ), .A3(
        \SB2_4_8/i0[8] ), .ZN(\SB2_4_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4973 ( .A1(\SB2_4_8/i0[10] ), .A2(\SB2_4_8/i1[9] ), .A3(
        \SB2_4_8/i1_7 ), .ZN(\SB2_4_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4975 ( .A1(\SB4_1/i1[9] ), .A2(n5442), .A3(\SB4_1/i0_4 ), .ZN(
        \SB4_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4977 ( .A1(\SB4_3/i0[6] ), .A2(\SB4_3/i1_5 ), .A3(\SB4_3/i0[9] ), 
        .ZN(\SB4_3/Component_Function_1/NAND4_in[2] ) );
  BUF_X2 U4981 ( .I(\SB3_5/buf_output[2] ), .Z(\SB4_2/i0_0 ) );
  NAND2_X1 U4983 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i1[9] ), .ZN(
        \SB4_20/Component_Function_1/NAND4_in[0] ) );
  INV_X1 U4984 ( .I(\SB3_7/buf_output[1] ), .ZN(\SB4_3/i1_7 ) );
  NAND3_X1 U4989 ( .A1(\SB1_4_8/i0[9] ), .A2(\SB1_4_8/i0_0 ), .A3(
        \SB1_4_8/i0[8] ), .ZN(\SB1_4_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U4992 ( .A1(\SB1_4_8/i0_0 ), .A2(\SB1_4_8/i0_3 ), .A3(
        \SB1_4_8/i0_4 ), .ZN(\SB1_4_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4996 ( .A1(\SB2_0_0/i0_3 ), .A2(\SB2_0_0/i0[7] ), .A3(
        \SB2_0_0/i0_0 ), .ZN(n2207) );
  NAND3_X1 U4999 ( .A1(\SB3_6/i0_3 ), .A2(\SB3_6/i0[10] ), .A3(\SB3_6/i0[6] ), 
        .ZN(\SB3_6/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U5003 ( .I(\SB1_4_25/buf_output[5] ), .Z(\SB2_4_25/i0_3 ) );
  NAND3_X1 U5005 ( .A1(\SB4_26/i0[6] ), .A2(n3989), .A3(\SB4_26/i0[7] ), .ZN(
        \SB4_26/Component_Function_0/NAND4_in[1] ) );
  INV_X1 U5007 ( .I(\MC_ARK_ARC_1_4/buf_output[175] ), .ZN(\SB3_2/i1_7 ) );
  NAND3_X1 U5010 ( .A1(\SB4_2/i1[9] ), .A2(\SB4_2/i0_4 ), .A3(\SB4_2/i0_3 ), 
        .ZN(\SB4_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U5011 ( .A1(\SB3_23/i0[7] ), .A2(\SB3_23/i0_3 ), .A3(\SB3_23/i0_0 ), 
        .ZN(\SB3_23/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 U5013 ( .I(\SB1_4_15/buf_output[5] ), .Z(\SB2_4_15/i0_3 ) );
  NAND3_X1 U5016 ( .A1(\SB2_4_15/i0_3 ), .A2(\SB2_4_15/i1_7 ), .A3(
        \SB2_4_15/i0[8] ), .ZN(\SB2_4_15/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U5035 ( .A1(\SB3_8/i0[6] ), .A2(\SB3_8/i0_4 ), .A3(\SB3_8/i0[9] ), 
        .ZN(n2353) );
  BUF_X2 U5042 ( .I(\SB3_18/buf_output[1] ), .Z(\SB4_14/i0[6] ) );
  NAND3_X1 U5044 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0[10] ), .A3(
        \SB1_1_20/i0[6] ), .ZN(\SB1_1_20/Component_Function_2/NAND4_in[1] ) );
  INV_X1 U5047 ( .I(\SB3_28/buf_output[1] ), .ZN(\SB4_24/i1_7 ) );
  INV_X1 U5052 ( .I(\SB3_4/buf_output[3] ), .ZN(\SB4_2/i0[8] ) );
  CLKBUF_X4 U5058 ( .I(\RI3[5][171] ), .Z(\SB4_3/i0[10] ) );
  BUF_X4 U5060 ( .I(\SB2_4_30/buf_output[5] ), .Z(\RI5[4][11] ) );
  NAND3_X1 U5061 ( .A1(\SB4_10/i0_3 ), .A2(\SB3_14/buf_output[1] ), .A3(
        \SB4_10/i1[9] ), .ZN(n2921) );
  CLKBUF_X4 U5062 ( .I(\MC_ARK_ARC_1_1/buf_output[140] ), .Z(\SB1_2_8/i0_0 )
         );
  NAND3_X1 U5064 ( .A1(\SB4_2/i0[9] ), .A2(\SB4_2/i0_0 ), .A3(\SB4_2/i0[8] ), 
        .ZN(\SB4_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U5065 ( .A1(\SB4_2/i1_5 ), .A2(\SB4_2/i0_0 ), .A3(\SB4_2/i0_4 ), 
        .ZN(\SB4_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U5066 ( .A1(\SB4_2/i0[7] ), .A2(\SB4_2/i0_3 ), .A3(\SB4_2/i0_0 ), 
        .ZN(\SB4_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U5069 ( .A1(\SB2_3_18/i0_0 ), .A2(\SB2_3_18/i1_5 ), .A3(
        \SB2_3_18/i0_4 ), .ZN(n2515) );
  NAND3_X1 U5070 ( .A1(\SB3_18/i0_0 ), .A2(\SB3_18/i0_3 ), .A3(\SB3_18/i0_4 ), 
        .ZN(\SB3_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U5078 ( .A1(\SB1_4_14/i0_3 ), .A2(\SB1_4_14/i1_7 ), .A3(
        \SB1_4_14/i0[8] ), .ZN(\SB1_4_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U5079 ( .A1(\SB3_4/i1[9] ), .A2(\SB3_4/i0_3 ), .A3(\SB3_4/i0[6] ), 
        .ZN(\SB3_4/Component_Function_3/NAND4_in[0] ) );
  BUF_X2 U5080 ( .I(\MC_ARK_ARC_1_4/buf_output[85] ), .Z(\SB3_17/i0[6] ) );
  NAND3_X1 U5081 ( .A1(\SB3_17/i0_3 ), .A2(\SB3_17/i1_7 ), .A3(\SB3_17/i0[8] ), 
        .ZN(\SB3_17/Component_Function_1/NAND4_in[1] ) );
  AND4_X2 U5087 ( .A1(\SB3_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_26/Component_Function_3/NAND4_in[3] ), .Z(n1494) );
  NAND3_X1 U5088 ( .A1(\SB3_16/i1[9] ), .A2(\SB3_16/i1_5 ), .A3(\SB3_16/i0_4 ), 
        .ZN(\SB3_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U5089 ( .A1(\SB3_16/i0[9] ), .A2(\SB3_16/i0[6] ), .A3(\SB3_16/i0_4 ), .ZN(\SB3_16/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U5096 ( .A1(\SB2_4_20/i0_3 ), .A2(\SB2_4_20/i1_7 ), .A3(
        \SB2_4_20/i0[8] ), .ZN(\SB2_4_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U5097 ( .A1(\SB2_4_0/i3[0] ), .A2(\SB2_4_0/i0_0 ), .A3(
        \SB2_4_0/i1_7 ), .ZN(\SB2_4_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U5100 ( .A1(\SB3_30/i1[9] ), .A2(\SB3_30/i1_5 ), .A3(\SB3_30/i0_4 ), 
        .ZN(\SB3_30/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U5103 ( .I(\RI1[5][80] ), .Z(\SB3_18/i0_0 ) );
  BUF_X2 U5104 ( .I(n353), .Z(\SB1_0_13/i0[10] ) );
  INV_X1 U5105 ( .I(n353), .ZN(\SB1_0_13/i0[8] ) );
  NAND2_X1 U5108 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i3[0] ), .ZN(
        \SB3_14/Component_Function_5/NAND4_in[0] ) );
  AND4_X2 U5116 ( .A1(\SB3_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_21/Component_Function_2/NAND4_in[3] ), .Z(n1496) );
  NAND3_X1 U5119 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i0[10] ), .A3(
        \SB4_20/i0[9] ), .ZN(\SB4_20/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U5124 ( .A1(\SB4_28/i0_0 ), .A2(\SB4_28/i3[0] ), .ZN(
        \SB4_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U5131 ( .A1(\SB4_7/i0_3 ), .A2(\SB3_9/buf_output[3] ), .A3(
        \SB4_7/i0_4 ), .ZN(\SB4_7/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 U5132 ( .A1(\SB4_9/i0[10] ), .A2(\SB4_9/i0[9] ), .ZN(n2308) );
  NAND3_X1 U5134 ( .A1(\SB4_9/i0[10] ), .A2(\SB4_9/i1[9] ), .A3(\SB4_9/i1_7 ), 
        .ZN(n2298) );
  NAND3_X1 U5135 ( .A1(\SB4_9/i0[10] ), .A2(\SB4_9/i0[9] ), .A3(\SB4_9/i0_3 ), 
        .ZN(n2107) );
  BUF_X4 U5142 ( .I(\SB2_3_17/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[99] ) );
  CLKBUF_X4 U5147 ( .I(\SB3_6/buf_output[2] ), .Z(\SB4_3/i0_0 ) );
  NAND3_X1 U5152 ( .A1(\SB3_27/i0[8] ), .A2(\SB3_27/i0[7] ), .A3(
        \SB3_27/i0[6] ), .ZN(\SB3_27/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U5153 ( .A1(\SB3_6/i1_7 ), .A2(\SB3_6/i0[8] ), .A3(\SB3_6/i0_4 ), 
        .ZN(\SB3_6/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U5155 ( .I(\MC_ARK_ARC_1_4/buf_output[109] ), .ZN(\SB3_13/i1_7 ) );
  AND4_X2 U5157 ( .A1(\SB3_17/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_3/NAND4_in[0] ), .A4(n3020), .Z(n1497) );
  AND4_X2 U5159 ( .A1(\SB3_15/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_15/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_15/Component_Function_3/NAND4_in[3] ), .A4(n2406), .Z(n1498) );
  NAND3_X1 U5160 ( .A1(\SB3_15/i0[10] ), .A2(\SB3_15/i1_7 ), .A3(
        \SB3_15/i1[9] ), .ZN(n2406) );
  INV_X1 U5161 ( .I(\MC_ARK_ARC_1_2/buf_output[121] ), .ZN(\SB1_3_11/i1_7 ) );
  INV_X1 U5163 ( .I(\SB3_26/buf_output[5] ), .ZN(\SB4_26/i1_5 ) );
  BUF_X4 U5164 ( .I(\SB2_4_29/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[27] ) );
  CLKBUF_X4 U5167 ( .I(\SB1_4_12/buf_output[4] ), .Z(\SB2_4_11/i0_4 ) );
  NAND3_X1 U5172 ( .A1(\SB3_21/i0_3 ), .A2(\SB3_21/i0[10] ), .A3(
        \SB3_21/i0[6] ), .ZN(\SB3_21/Component_Function_2/NAND4_in[1] ) );
  INV_X1 U5176 ( .I(\SB3_25/buf_output[1] ), .ZN(\SB4_21/i1_7 ) );
  INV_X1 U5182 ( .I(\MC_ARK_ARC_1_4/buf_output[139] ), .ZN(\SB3_8/i1_7 ) );
  INV_X1 U5186 ( .I(\SB3_1/buf_output[0] ), .ZN(\SB4_28/i3[0] ) );
  NAND3_X1 U5188 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i0[10] ), .A3(\SB3_1/i0_4 ), 
        .ZN(n2409) );
  NAND3_X1 U5194 ( .A1(\SB1_4_13/i0_3 ), .A2(\SB1_4_13/i1_7 ), .A3(
        \SB1_4_13/i0[8] ), .ZN(\SB1_4_13/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X4 U5198 ( .I(\MC_ARK_ARC_1_3/buf_output[160] ), .Z(\SB1_4_5/i0_4 )
         );
  NAND3_X1 U5199 ( .A1(\SB4_2/i0_0 ), .A2(\SB4_2/i3[0] ), .A3(\SB4_2/i1_7 ), 
        .ZN(n2898) );
  NAND3_X1 U5201 ( .A1(\SB4_7/i0_4 ), .A2(\SB4_7/i1[9] ), .A3(\SB4_7/i1_5 ), 
        .ZN(n2506) );
  NAND2_X1 U5202 ( .A1(\SB4_7/i0_3 ), .A2(\SB4_7/i1[9] ), .ZN(
        \SB4_7/Component_Function_1/NAND4_in[0] ) );
  BUF_X4 U5208 ( .I(\SB2_4_6/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[170] ) );
  NAND3_X1 U5212 ( .A1(\SB4_0/i0_3 ), .A2(\SB4_0/i0_4 ), .A3(\SB4_0/i1[9] ), 
        .ZN(\SB4_0/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U5213 ( .I(\SB2_4_21/buf_output[2] ), .Z(\RI5[4][80] ) );
  CLKBUF_X4 U5214 ( .I(\SB3_27/buf_output[5] ), .Z(\SB4_27/i0_3 ) );
  BUF_X4 U5215 ( .I(\SB2_4_2/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[184] ) );
  CLKBUF_X4 U5219 ( .I(\SB1_4_4/buf_output[3] ), .Z(\SB2_4_2/i0[10] ) );
  BUF_X4 U5222 ( .I(\SB2_4_15/buf_output[4] ), .Z(\RI5[4][106] ) );
  NAND3_X1 U5223 ( .A1(\SB1_4_9/i0_3 ), .A2(\SB1_4_9/i0[7] ), .A3(
        \SB1_4_9/i0_0 ), .ZN(n2348) );
  NAND3_X1 U5224 ( .A1(\SB1_4_9/i0_3 ), .A2(\SB1_4_9/i0[10] ), .A3(
        \SB1_4_9/i0[9] ), .ZN(\SB1_4_9/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U5227 ( .I(\MC_ARK_ARC_1_0/buf_output[115] ), .ZN(\SB1_1_12/i1_7 ) );
  CLKBUF_X4 U5232 ( .I(\MC_ARK_ARC_1_2/buf_output[159] ), .Z(\SB1_3_5/i0[10] )
         );
  CLKBUF_X4 U5245 ( .I(\MC_ARK_ARC_1_0/buf_output[136] ), .Z(\SB1_1_9/i0_4 )
         );
  BUF_X4 U5254 ( .I(\SB2_2_4/buf_output[5] ), .Z(\RI5[2][167] ) );
  BUF_X4 U5255 ( .I(\SB2_4_7/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[169] ) );
  NAND3_X1 U5256 ( .A1(\SB4_1/i0_3 ), .A2(\SB4_1/i0[7] ), .A3(\SB4_1/i0_0 ), 
        .ZN(\SB4_1/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U5258 ( .A1(\SB4_1/i0_3 ), .A2(\SB4_1/i1[9] ), .ZN(
        \SB4_1/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 U5259 ( .A1(\SB4_4/i0[10] ), .A2(\SB4_4/i0[9] ), .ZN(n2684) );
  CLKBUF_X4 U5263 ( .I(\MC_ARK_ARC_1_4/buf_output[51] ), .Z(\SB3_23/i0[10] )
         );
  OR3_X2 U5269 ( .A1(\MC_ARK_ARC_1_0/buf_output[102] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[107] ), .A3(
        \MC_ARK_ARC_1_0/buf_output[105] ), .Z(n2712) );
  NAND3_X1 U5272 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i0_3 ), .A3(\SB4_8/i0_4 ), 
        .ZN(\SB4_8/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U5277 ( .I(\SB1_4_31/buf_output[1] ), .ZN(\SB2_4_27/i1_7 ) );
  NAND3_X1 U5282 ( .A1(\SB4_28/i0[9] ), .A2(\SB4_28/i0_0 ), .A3(\SB4_28/i0[8] ), .ZN(\SB4_28/Component_Function_4/NAND4_in[0] ) );
  INV_X1 U5292 ( .I(\RI1[5][167] ), .ZN(\SB3_4/i1_5 ) );
  NAND3_X1 U5297 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i1[9] ), .A3(
        \SB4_10/i1_7 ), .ZN(n2739) );
  NAND3_X1 U5298 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i0[6] ), .A3(
        \SB4_10/i0[10] ), .ZN(\SB4_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U5299 ( .A1(\SB4_10/i0_3 ), .A2(\SB4_10/i0[10] ), .A3(\SB4_10/i0_4 ), .ZN(n3157) );
  BUF_X4 U5300 ( .I(\SB2_4_14/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[132] ) );
  AND2_X2 U5301 ( .A1(\MC_ARK_ARC_1_0/buf_output[176] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[178] ), .Z(n2614) );
  NAND2_X1 U5303 ( .A1(\SB4_7/i0_0 ), .A2(\SB4_7/i3[0] ), .ZN(
        \SB4_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U5304 ( .A1(\SB4_7/i0_0 ), .A2(\SB4_7/i0[6] ), .A3(
        \SB3_9/buf_output[3] ), .ZN(\SB4_7/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U5305 ( .A1(\SB4_7/i0[7] ), .A2(\SB4_7/i0_3 ), .A3(\SB4_7/i0_0 ), 
        .ZN(\SB4_7/Component_Function_0/NAND4_in[3] ) );
  INV_X1 U5309 ( .I(\SB3_11/buf_output[1] ), .ZN(\SB4_7/i1_7 ) );
  OR3_X1 U5316 ( .A1(\RI1[2][101] ), .A2(n1509), .A3(
        \MC_ARK_ARC_1_1/buf_output[96] ), .Z(n2012) );
  INV_X1 U5317 ( .I(\MC_ARK_ARC_1_1/buf_output[96] ), .ZN(\SB1_2_15/i3[0] ) );
  CLKBUF_X4 U5318 ( .I(\MC_ARK_ARC_1_2/buf_output[171] ), .Z(\SB1_3_3/i0[10] )
         );
  NAND3_X1 U5320 ( .A1(\SB1_2_11/i0[9] ), .A2(\SB1_2_11/i0[10] ), .A3(
        \SB1_2_11/i0_3 ), .ZN(\SB1_2_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U5321 ( .A1(\SB3_3/i0_0 ), .A2(\SB3_3/i1_5 ), .A3(\SB3_3/i0_4 ), 
        .ZN(\SB3_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U5322 ( .A1(\SB3_3/i1_5 ), .A2(\SB3_3/i0[8] ), .A3(\SB3_3/i3[0] ), 
        .ZN(\SB3_3/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X4 U5323 ( .I(\RI3[0][154] ), .Z(\SB2_0_6/i0_4 ) );
  INV_X1 U5327 ( .I(\MC_ARK_ARC_1_4/buf_output[67] ), .ZN(\SB3_20/i1_7 ) );
  NAND3_X1 U5335 ( .A1(\RI1[2][101] ), .A2(\SB1_2_15/i0[9] ), .A3(
        \SB1_2_15/i0[10] ), .ZN(n2902) );
  NAND3_X1 U5336 ( .A1(\RI1[2][101] ), .A2(\SB1_2_15/i1_7 ), .A3(
        \SB1_2_15/i0[8] ), .ZN(\SB1_2_15/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X4 U5343 ( .I(n256), .Z(\SB1_0_30/i0_0 ) );
  INV_X1 U5345 ( .I(\MC_ARK_ARC_1_1/buf_output[1] ), .ZN(\SB1_2_31/i1_7 ) );
  BUF_X2 U5346 ( .I(\MC_ARK_ARC_1_1/buf_output[1] ), .Z(\SB1_2_31/i0[6] ) );
  BUF_X4 U5351 ( .I(\SB2_3_7/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[164] ) );
  NAND3_X1 U5352 ( .A1(\SB4_29/i0_4 ), .A2(\SB4_29/i1[9] ), .A3(\SB4_29/i1_5 ), 
        .ZN(n2912) );
  XOR2_X1 U5356 ( .A1(\MC_ARK_ARC_1_3/temp6[123] ), .A2(n2669), .Z(n1504) );
  INV_X1 U5359 ( .I(\SB3_8/buf_output[5] ), .ZN(\SB4_8/i1_5 ) );
  CLKBUF_X4 U5363 ( .I(\SB1_4_2/buf_output[2] ), .Z(\SB2_4_31/i0_0 ) );
  NAND2_X1 U5374 ( .A1(\SB4_21/i0_3 ), .A2(n3998), .ZN(n1699) );
  CLKBUF_X4 U5379 ( .I(\RI3[0][147] ), .Z(\SB2_0_7/i0[10] ) );
  CLKBUF_X4 U5381 ( .I(\MC_ARK_ARC_1_4/buf_output[9] ), .Z(\SB3_30/i0[10] ) );
  NAND3_X1 U5385 ( .A1(\SB1_3_5/i3[0] ), .A2(\SB1_3_5/i0_0 ), .A3(
        \SB1_3_5/i1_7 ), .ZN(\SB1_3_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U5386 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i1_7 ), .A3(
        \SB1_3_5/i0[8] ), .ZN(\SB1_3_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U5387 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i1[9] ), .A3(\SB3_7/i1_7 ), 
        .ZN(n2436) );
  CLKBUF_X4 U5394 ( .I(\MC_ARK_ARC_1_3/buf_output[122] ), .Z(\SB1_4_11/i0_0 )
         );
  NAND3_X1 U5395 ( .A1(\SB4_8/i0_4 ), .A2(n3996), .A3(\SB4_8/i1_5 ), .ZN(n2969) );
  NAND2_X1 U5396 ( .A1(\SB4_8/i0_3 ), .A2(n3996), .ZN(
        \SB4_8/Component_Function_1/NAND4_in[0] ) );
  BUF_X4 U5400 ( .I(\SB2_1_20/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[76] ) );
  BUF_X4 U5401 ( .I(\RI3[2][131] ), .Z(\SB2_2_10/i0_3 ) );
  CLKBUF_X4 U5402 ( .I(\MC_ARK_ARC_1_1/buf_output[128] ), .Z(\SB1_2_10/i0_0 )
         );
  INV_X1 U5403 ( .I(\SB3_3/buf_output[1] ), .ZN(\SB4_31/i1_7 ) );
  INV_X1 U5405 ( .I(\MC_ARK_ARC_1_3/buf_output[138] ), .ZN(\SB1_4_8/i3[0] ) );
  INV_X1 U5408 ( .I(\SB1_4_4/buf_output[1] ), .ZN(\SB2_4_0/i1_7 ) );
  NAND3_X1 U5409 ( .A1(\SB2_4_10/i0_3 ), .A2(\SB2_4_10/i1_7 ), .A3(
        \SB2_4_10/i0[8] ), .ZN(\SB2_4_10/Component_Function_1/NAND4_in[1] ) );
  INV_X1 U5416 ( .I(\SB3_14/buf_output[1] ), .ZN(\SB4_10/i1_7 ) );
  NAND3_X1 U5419 ( .A1(\SB4_28/i0_4 ), .A2(\SB4_28/i1_5 ), .A3(\SB4_28/i1[9] ), 
        .ZN(n2864) );
  NAND3_X1 U5423 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i0_4 ), .A3(\RI1[5][185] ), 
        .ZN(\SB3_1/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U5428 ( .I(\MC_ARK_ARC_1_3/buf_output[123] ), .Z(\SB1_4_11/i0[10] ) );
  CLKBUF_X4 U5432 ( .I(\MC_ARK_ARC_1_1/buf_output[2] ), .Z(\SB1_2_31/i0_0 ) );
  CLKBUF_X4 U5433 ( .I(\SB1_3_10/buf_output[2] ), .Z(\SB2_3_7/i0_0 ) );
  INV_X1 U5437 ( .I(n388), .ZN(\SB1_0_24/i1_5 ) );
  NAND3_X1 U5439 ( .A1(\SB1_4_11/i0_0 ), .A2(\SB1_4_11/i0[6] ), .A3(
        \SB1_4_11/i0[10] ), .ZN(\SB1_4_11/Component_Function_5/NAND4_in[1] )
         );
  XOR2_X1 U5440 ( .A1(Key[80]), .A2(Plaintext[80]), .Z(n1507) );
  AND4_X2 U5441 ( .A1(\SB1_0_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_18/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_18/Component_Function_2/NAND4_in[2] ), .A4(n2829), .Z(n1508) );
  XOR2_X1 U5452 ( .A1(n1546), .A2(\MC_ARK_ARC_1_2/temp6[146] ), .Z(n1510) );
  NAND3_X1 U5486 ( .A1(\SB1_0_2/i0[6] ), .A2(\SB1_0_2/i0[7] ), .A3(
        \SB1_0_2/i0[8] ), .ZN(\SB1_0_2/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U5487 ( .A1(\SB1_0_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_2/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_2/Component_Function_1/NAND4_in[0] ), .A4(n1519), .ZN(
        \SB1_0_2/buf_output[1] ) );
  XOR2_X1 U5495 ( .A1(\RI5[3][60] ), .A2(\RI5[3][84] ), .Z(
        \MC_ARK_ARC_1_3/temp2[114] ) );
  XOR2_X1 U5496 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[49] ), .A2(\RI5[2][85] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[175] ) );
  XOR2_X1 U5505 ( .A1(n1526), .A2(\MC_ARK_ARC_1_4/temp6[72] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[72] ) );
  XOR2_X1 U5506 ( .A1(\MC_ARK_ARC_1_4/temp1[72] ), .A2(
        \MC_ARK_ARC_1_4/temp2[72] ), .Z(n1526) );
  NAND4_X2 U5513 ( .A1(\SB2_2_15/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_15/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_15/Component_Function_4/NAND4_in[0] ), .A4(n1529), .ZN(
        \SB2_2_15/buf_output[4] ) );
  BUF_X4 U5516 ( .I(\SB2_1_20/buf_output[2] ), .Z(\RI5[1][86] ) );
  NAND4_X2 U5521 ( .A1(\SB2_4_28/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_4_28/Component_Function_0/NAND4_in[1] ), .A3(n2124), .A4(
        \SB2_4_28/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_4_28/buf_output[0] ) );
  NAND3_X2 U5522 ( .A1(\SB2_4_20/i0[10] ), .A2(\SB2_4_20/i1[9] ), .A3(
        \SB2_4_20/i1_7 ), .ZN(\SB2_4_20/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U5527 ( .A1(\MC_ARK_ARC_1_0/temp2[158] ), .A2(
        \MC_ARK_ARC_1_0/temp1[158] ), .Z(\MC_ARK_ARC_1_0/temp5[158] ) );
  NAND4_X2 U5534 ( .A1(\SB2_0_9/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_9/Component_Function_0/NAND4_in[0] ), .A3(n2628), .A4(
        \SB2_0_9/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_0_9/buf_output[0] ) );
  XOR2_X1 U5539 ( .A1(n1788), .A2(\MC_ARK_ARC_1_4/temp1[15] ), .Z(n1535) );
  XOR2_X1 U5546 ( .A1(\MC_ARK_ARC_1_3/temp4[103] ), .A2(n1541), .Z(
        \MC_ARK_ARC_1_3/temp6[103] ) );
  XOR2_X1 U5547 ( .A1(\RI5[3][169] ), .A2(\RI5[3][13] ), .Z(n1541) );
  XOR2_X1 U5548 ( .A1(\RI5[0][126] ), .A2(\RI5[0][162] ), .Z(
        \MC_ARK_ARC_1_0/temp3[60] ) );
  XOR2_X1 U5551 ( .A1(\MC_ARK_ARC_1_4/temp1[39] ), .A2(n1543), .Z(n2103) );
  XOR2_X1 U5552 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[9] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[177] ), .Z(n1543) );
  XOR2_X1 U5563 ( .A1(\SB2_0_16/buf_output[0] ), .A2(\RI5[0][126] ), .Z(
        \MC_ARK_ARC_1_0/temp1[126] ) );
  XOR2_X1 U5571 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[137] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[173] ), .Z(n1550) );
  NAND3_X2 U5572 ( .A1(\SB2_1_10/i0[6] ), .A2(\SB2_1_10/i0_3 ), .A3(
        \SB2_1_10/i1[9] ), .ZN(n1551) );
  NAND4_X2 U5581 ( .A1(\SB1_0_22/Component_Function_5/NAND4_in[1] ), .A2(n2074), .A3(\SB1_0_22/Component_Function_5/NAND4_in[0] ), .A4(n2400), .ZN(
        \SB1_0_22/buf_output[5] ) );
  XOR2_X1 U5584 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), .A2(\RI5[2][5] ), 
        .Z(n1557) );
  NAND3_X2 U5585 ( .A1(\SB2_1_20/i0[7] ), .A2(\SB2_1_20/i0[8] ), .A3(
        \SB2_1_20/i0[6] ), .ZN(\SB2_1_20/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U5587 ( .A1(\MC_ARK_ARC_1_3/temp4[127] ), .A2(
        \MC_ARK_ARC_1_3/temp3[127] ), .Z(n1558) );
  BUF_X4 U5588 ( .I(\SB2_1_20/buf_output[0] ), .Z(\RI5[1][96] ) );
  XOR2_X1 U5591 ( .A1(n1789), .A2(n1560), .Z(\MC_ARK_ARC_1_4/temp5[173] ) );
  XOR2_X1 U5592 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[167] ), .A2(\RI5[4][119] ), 
        .Z(n1560) );
  NAND4_X2 U5593 ( .A1(\SB2_2_1/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_2_1/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_2_1/Component_Function_2/NAND4_in[2] ), .A4(n1655), .ZN(
        \SB2_2_1/buf_output[2] ) );
  BUF_X4 U5594 ( .I(\SB2_2_1/buf_output[2] ), .Z(\RI5[2][8] ) );
  NAND3_X2 U5600 ( .A1(\SB2_4_4/i0[10] ), .A2(\SB2_4_4/i0_0 ), .A3(
        \SB2_4_4/i0[6] ), .ZN(\SB2_4_4/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U5601 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0[9] ), .A3(
        \SB2_1_10/i0[8] ), .ZN(\SB2_1_10/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U5607 ( .A1(n1566), .A2(\MC_ARK_ARC_1_0/temp4[142] ), .Z(
        \MC_ARK_ARC_1_0/temp6[142] ) );
  XOR2_X1 U5608 ( .A1(\RI5[0][16] ), .A2(\RI5[0][52] ), .Z(n1566) );
  XOR2_X1 U5614 ( .A1(n1569), .A2(\MC_ARK_ARC_1_0/temp6[47] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[47] ) );
  XOR2_X1 U5616 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[84] ), .A2(
        \SB2_2_18/buf_output[0] ), .Z(\MC_ARK_ARC_1_2/temp2[138] ) );
  BUF_X4 U5621 ( .I(\SB2_2_2/buf_output[0] ), .Z(\RI5[2][12] ) );
  XOR2_X1 U5628 ( .A1(\RI5[1][39] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[45] ), 
        .Z(n1574) );
  NAND2_X1 U5630 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i1[9] ), .ZN(n1575) );
  INV_X1 U5634 ( .I(\SB1_2_31/buf_output[0] ), .ZN(\SB2_2_26/i3[0] ) );
  NAND4_X2 U5635 ( .A1(\SB1_2_31/Component_Function_0/NAND4_in[1] ), .A2(n2642), .A3(\SB1_2_31/Component_Function_0/NAND4_in[0] ), .A4(n2641), .ZN(
        \SB1_2_31/buf_output[0] ) );
  BUF_X4 U5641 ( .I(\SB2_0_20/buf_output[4] ), .Z(\RI5[0][76] ) );
  XOR2_X1 U5642 ( .A1(\MC_ARK_ARC_1_2/temp2[95] ), .A2(n1580), .Z(
        \MC_ARK_ARC_1_2/temp5[95] ) );
  XOR2_X1 U5643 ( .A1(\RI5[2][95] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[89] ), 
        .Z(n1580) );
  NAND3_X2 U5644 ( .A1(\SB2_1_3/i0[10] ), .A2(\SB2_1_3/i1[9] ), .A3(
        \SB2_1_3/i1_7 ), .ZN(\SB2_1_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U5649 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0[8] ), .A3(
        \SB1_1_30/i1_7 ), .ZN(\SB1_1_30/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U5655 ( .A1(n2507), .A2(\SB1_1_2/Component_Function_4/NAND4_in[0] ), 
        .A3(\SB1_1_2/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_1_2/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_1_2/buf_output[4] ) );
  NAND4_X2 U5657 ( .A1(\SB2_0_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_2/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_2/Component_Function_5/NAND4_in[0] ), .A4(n1587), .ZN(
        \SB2_0_2/buf_output[5] ) );
  BUF_X4 U5658 ( .I(\SB2_1_1/buf_output[0] ), .Z(\RI5[1][18] ) );
  BUF_X4 U5661 ( .I(\SB2_3_31/buf_output[1] ), .Z(\RI5[3][25] ) );
  NAND2_X1 U5668 ( .A1(\SB1_3_13/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_3_13/Component_Function_4/NAND4_in[1] ), .ZN(n1592) );
  NAND3_X2 U5672 ( .A1(\RI1[2][149] ), .A2(\SB1_2_7/i0[10] ), .A3(
        \SB1_2_7/i0[9] ), .ZN(\SB1_2_7/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U5673 ( .A1(n1596), .A2(n2242), .Z(\MC_ARK_ARC_1_1/buf_output[149] )
         );
  XOR2_X1 U5681 ( .A1(\MC_ARK_ARC_1_4/temp1[145] ), .A2(
        \MC_ARK_ARC_1_4/temp2[145] ), .Z(\MC_ARK_ARC_1_4/temp5[145] ) );
  XOR2_X1 U5689 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[121] ), .A2(\RI5[2][145] ), 
        .Z(n1604) );
  NAND3_X2 U5698 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0_0 ), .A3(
        \SB2_2_22/i0_4 ), .ZN(\SB2_2_22/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U5699 ( .A1(n2192), .A2(\MC_ARK_ARC_1_3/temp5[80] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[80] ) );
  NAND3_X1 U5702 ( .A1(\SB2_1_7/i0_4 ), .A2(\SB2_1_7/i1_7 ), .A3(
        \SB2_1_7/i0[8] ), .ZN(\SB2_1_7/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U5706 ( .A1(\SB1_4_31/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_4_31/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_4_31/Component_Function_1/NAND4_in[1] ), .A4(n1610), .ZN(
        \SB1_4_31/buf_output[1] ) );
  NAND4_X2 U5711 ( .A1(\SB2_3_30/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_30/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_30/Component_Function_0/NAND4_in[0] ), .A4(n1613), .ZN(
        \SB2_3_30/buf_output[0] ) );
  BUF_X4 U5712 ( .I(\SB2_2_13/buf_output[5] ), .Z(\RI5[2][113] ) );
  NAND3_X2 U5716 ( .A1(\SB1_0_31/i0[10] ), .A2(\SB1_0_31/i0_0 ), .A3(
        \SB1_0_31/i0[6] ), .ZN(n1614) );
  INV_X2 U5718 ( .I(\SB1_0_2/buf_output[2] ), .ZN(\SB2_0_31/i1[9] ) );
  NAND3_X1 U5724 ( .A1(\SB1_2_31/i0_0 ), .A2(\SB1_2_31/i1_5 ), .A3(
        \SB1_2_31/i0_4 ), .ZN(n1618) );
  XOR2_X1 U5731 ( .A1(\RI5[0][189] ), .A2(\RI5[0][3] ), .Z(
        \MC_ARK_ARC_1_0/temp1[3] ) );
  NAND3_X2 U5732 ( .A1(\SB1_0_9/i0[6] ), .A2(\SB1_0_9/i0[9] ), .A3(
        \SB1_0_9/i0_4 ), .ZN(\SB1_0_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U5735 ( .A1(\SB1_1_1/i0_3 ), .A2(\SB1_1_1/i0[8] ), .A3(
        \SB1_1_1/i1_7 ), .ZN(\SB1_1_1/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U5758 ( .A1(\RI5[0][63] ), .A2(\RI5[0][27] ), .Z(
        \MC_ARK_ARC_1_0/temp3[153] ) );
  XOR2_X1 U5759 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[25] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[181] ), .Z(\MC_ARK_ARC_1_2/temp3[115] )
         );
  NAND4_X2 U5762 ( .A1(\SB1_1_31/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_31/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_1_31/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_31/buf_output[0] ) );
  NAND4_X2 U5763 ( .A1(\SB2_1_26/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_26/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_26/Component_Function_4/NAND4_in[1] ), .A4(n2047), .ZN(
        \SB2_1_26/buf_output[4] ) );
  XOR2_X1 U5765 ( .A1(\MC_ARK_ARC_1_0/temp5[115] ), .A2(
        \MC_ARK_ARC_1_0/temp6[115] ), .Z(\MC_ARK_ARC_1_0/buf_output[115] ) );
  BUF_X4 U5771 ( .I(\SB2_1_12/buf_output[0] ), .Z(\RI5[1][144] ) );
  XOR2_X1 U5772 ( .A1(\MC_ARK_ARC_1_3/temp3[68] ), .A2(
        \MC_ARK_ARC_1_3/temp4[68] ), .Z(\MC_ARK_ARC_1_3/temp6[68] ) );
  XOR2_X1 U5773 ( .A1(n1641), .A2(n1640), .Z(\MC_ARK_ARC_1_0/buf_output[172] )
         );
  XOR2_X1 U5774 ( .A1(\MC_ARK_ARC_1_0/temp4[172] ), .A2(
        \MC_ARK_ARC_1_0/temp1[172] ), .Z(n1640) );
  XOR2_X1 U5777 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[162] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[168] ), .Z(\MC_ARK_ARC_1_1/temp1[168] )
         );
  INV_X2 U5778 ( .I(\SB1_1_18/buf_output[3] ), .ZN(\SB2_1_16/i0[8] ) );
  NAND4_X2 U5779 ( .A1(\SB1_1_18/Component_Function_3/NAND4_in[1] ), .A2(n2834), .A3(n1892), .A4(\SB1_1_18/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_18/buf_output[3] ) );
  XOR2_X1 U5783 ( .A1(\MC_ARK_ARC_1_0/temp4[191] ), .A2(
        \MC_ARK_ARC_1_0/temp2[191] ), .Z(n1647) );
  NAND4_X2 U5789 ( .A1(\SB1_1_18/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_1_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_18/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_1_18/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB1_1_18/buf_output[0] ) );
  BUF_X4 U5795 ( .I(\SB2_2_6/buf_output[2] ), .Z(\RI5[2][170] ) );
  XOR2_X1 U5799 ( .A1(n1656), .A2(\MC_ARK_ARC_1_4/temp6[153] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[153] ) );
  NAND3_X1 U5805 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB2_1_18/i0[10] ), .A3(
        \SB2_1_18/i0_4 ), .ZN(n1660) );
  AND2_X1 U5807 ( .A1(\SB2_1_1/i1_7 ), .A2(\SB2_1_1/i0[8] ), .Z(n1898) );
  XOR2_X1 U5809 ( .A1(\RI5[1][65] ), .A2(\RI5[1][29] ), .Z(
        \MC_ARK_ARC_1_1/temp3[155] ) );
  XOR2_X1 U5811 ( .A1(\MC_ARK_ARC_1_1/temp6[155] ), .A2(
        \MC_ARK_ARC_1_1/temp5[155] ), .Z(\MC_ARK_ARC_1_1/buf_output[155] ) );
  XOR2_X1 U5813 ( .A1(n2304), .A2(n2305), .Z(\MC_ARK_ARC_1_2/temp6[139] ) );
  NAND4_X2 U5816 ( .A1(\SB2_2_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_1/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_1/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_1/buf_output[1] ) );
  NAND3_X1 U5821 ( .A1(\SB3_19/i0[8] ), .A2(\SB3_19/i1_5 ), .A3(\SB3_19/i3[0] ), .ZN(\SB3_19/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U5829 ( .A1(\RI5[1][55] ), .A2(\RI5[1][79] ), .Z(n1671) );
  XOR2_X1 U5831 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[117] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[93] ), .Z(n1672) );
  XOR2_X1 U5839 ( .A1(\MC_ARK_ARC_1_1/temp2[39] ), .A2(n1677), .Z(
        \MC_ARK_ARC_1_1/temp5[39] ) );
  XOR2_X1 U5840 ( .A1(\RI5[1][39] ), .A2(\RI5[1][33] ), .Z(n1677) );
  XOR2_X1 U5841 ( .A1(n1678), .A2(\MC_ARK_ARC_1_1/temp2[93] ), .Z(
        \MC_ARK_ARC_1_1/temp5[93] ) );
  NAND3_X2 U5845 ( .A1(\SB2_1_19/i0[10] ), .A2(\SB2_1_19/i1[9] ), .A3(
        \SB2_1_19/i1_7 ), .ZN(\SB2_1_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U5846 ( .A1(\SB2_4_14/i0[10] ), .A2(\SB2_4_14/i1[9] ), .A3(
        \SB2_4_14/i1_7 ), .ZN(\SB2_4_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U5850 ( .A1(\SB2_4_4/i0_4 ), .A2(\SB2_4_4/i0[6] ), .A3(
        \SB2_4_4/i0[9] ), .ZN(n1682) );
  XOR2_X1 U5852 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[167] ), .A2(\RI5[4][143] ), 
        .Z(n1683) );
  NAND3_X1 U5855 ( .A1(\SB1_3_10/i0[10] ), .A2(\SB1_3_10/i1[9] ), .A3(
        \SB1_3_10/i1_5 ), .ZN(\SB1_3_10/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U5858 ( .A1(\MC_ARK_ARC_1_3/temp6[157] ), .A2(n1685), .Z(
        \MC_ARK_ARC_1_3/buf_output[157] ) );
  XOR2_X1 U5859 ( .A1(\MC_ARK_ARC_1_3/temp1[157] ), .A2(
        \MC_ARK_ARC_1_3/temp2[157] ), .Z(n1685) );
  XOR2_X1 U5861 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[151] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[187] ), .Z(\MC_ARK_ARC_1_3/temp3[85] )
         );
  NAND2_X1 U5862 ( .A1(\SB3_12/i1[9] ), .A2(\RI1[5][119] ), .ZN(
        \SB3_12/Component_Function_1/NAND4_in[0] ) );
  XOR2_X1 U5863 ( .A1(\MC_ARK_ARC_1_3/temp5[85] ), .A2(
        \MC_ARK_ARC_1_3/temp6[85] ), .Z(\MC_ARK_ARC_1_3/buf_output[85] ) );
  NAND3_X1 U5871 ( .A1(\SB4_18/i0[8] ), .A2(\SB4_18/i3[0] ), .A3(\SB4_18/i1_5 ), .ZN(n1689) );
  NAND3_X1 U5876 ( .A1(n6716), .A2(\SB2_3_21/i0_0 ), .A3(\SB2_3_21/i0_3 ), 
        .ZN(\SB2_3_21/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U5885 ( .A1(\MC_ARK_ARC_1_0/temp6[8] ), .A2(
        \MC_ARK_ARC_1_0/temp5[8] ), .Z(\MC_ARK_ARC_1_0/buf_output[8] ) );
  BUF_X4 U5892 ( .I(\SB2_3_18/buf_output[2] ), .Z(\RI5[3][98] ) );
  INV_X2 U5895 ( .I(\SB1_3_29/buf_output[3] ), .ZN(\SB2_3_27/i0[8] ) );
  NAND3_X1 U5896 ( .A1(\SB1_1_3/buf_output[1] ), .A2(\SB2_1_31/i1_5 ), .A3(
        \SB2_1_31/i0[9] ), .ZN(\SB2_1_31/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U5898 ( .A1(n1695), .A2(\MC_ARK_ARC_1_3/temp6[101] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[101] ) );
  XOR2_X1 U5899 ( .A1(\MC_ARK_ARC_1_3/temp2[101] ), .A2(
        \MC_ARK_ARC_1_3/temp1[101] ), .Z(n1695) );
  INV_X1 U5900 ( .I(\SB3_12/buf_output[1] ), .ZN(\SB4_8/i1_7 ) );
  NAND4_X2 U5901 ( .A1(\SB3_12/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_12/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_12/buf_output[1] ) );
  NAND3_X1 U5902 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i1_5 ), .A3(
        \SB4_11/i1[9] ), .ZN(n1696) );
  XOR2_X1 U5904 ( .A1(\RI5[1][20] ), .A2(\RI5[1][56] ), .Z(
        \MC_ARK_ARC_1_1/temp3[146] ) );
  NAND3_X2 U5909 ( .A1(\SB2_2_31/i0_3 ), .A2(\SB2_2_31/i0[10] ), .A3(
        \SB2_2_31/i0[6] ), .ZN(\SB2_2_31/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U5910 ( .A1(n2243), .A2(\SB1_2_7/Component_Function_0/NAND4_in[1] ), 
        .A3(\SB1_2_7/Component_Function_0/NAND4_in[0] ), .A4(n1700), .ZN(
        \SB1_2_7/buf_output[0] ) );
  XOR2_X1 U5912 ( .A1(n2961), .A2(\MC_ARK_ARC_1_2/temp3[26] ), .Z(n1702) );
  XOR2_X1 U5916 ( .A1(\MC_ARK_ARC_1_3/temp2[1] ), .A2(
        \MC_ARK_ARC_1_3/temp1[1] ), .Z(n1705) );
  XOR2_X1 U5919 ( .A1(\MC_ARK_ARC_1_1/temp6[76] ), .A2(
        \MC_ARK_ARC_1_1/temp5[76] ), .Z(\MC_ARK_ARC_1_1/buf_output[76] ) );
  NAND3_X2 U5923 ( .A1(n2886), .A2(\SB2_0_9/i0[10] ), .A3(\SB2_0_9/i0[6] ), 
        .ZN(n1708) );
  XOR2_X1 U5925 ( .A1(n2832), .A2(n1709), .Z(\MC_ARK_ARC_1_0/buf_output[42] )
         );
  XOR2_X1 U5926 ( .A1(\MC_ARK_ARC_1_0/temp1[42] ), .A2(
        \MC_ARK_ARC_1_0/temp2[42] ), .Z(n1709) );
  NAND3_X1 U5927 ( .A1(\SB1_4_2/i0[10] ), .A2(\SB1_4_2/i1[9] ), .A3(
        \SB1_4_2/i1_5 ), .ZN(\SB1_4_2/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 U5930 ( .A1(\SB1_1_2/i1[9] ), .A2(\SB1_1_2/i0_3 ), .ZN(n1711) );
  XOR2_X1 U5936 ( .A1(\MC_ARK_ARC_1_3/temp1[80] ), .A2(n2147), .Z(
        \MC_ARK_ARC_1_3/temp5[80] ) );
  XOR2_X1 U5938 ( .A1(\RI5[0][9] ), .A2(\RI5[0][165] ), .Z(n1713) );
  NAND4_X2 U5939 ( .A1(\SB2_1_9/Component_Function_0/NAND4_in[1] ), .A2(n2270), 
        .A3(\SB2_1_9/Component_Function_0/NAND4_in[0] ), .A4(n1714), .ZN(
        \SB2_1_9/buf_output[0] ) );
  XOR2_X1 U5941 ( .A1(\RI5[0][181] ), .A2(\RI5[0][145] ), .Z(n1715) );
  NAND3_X2 U5943 ( .A1(\SB2_0_22/i0[8] ), .A2(\SB2_0_22/i0_3 ), .A3(
        \SB2_0_22/i0[9] ), .ZN(\SB2_0_22/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 U5944 ( .A1(\SB1_0_10/i0[9] ), .A2(\SB1_0_10/i0[10] ), .ZN(
        \SB1_0_10/Component_Function_0/NAND4_in[0] ) );
  NAND4_X2 U5954 ( .A1(\SB3_16/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_0/NAND4_in[0] ), .A4(n1721), .ZN(
        \SB3_16/buf_output[0] ) );
  NAND3_X1 U5959 ( .A1(\SB4_12/i0_3 ), .A2(\SB4_12/i0[10] ), .A3(
        \SB4_12/i0[9] ), .ZN(n1726) );
  XOR2_X1 U5962 ( .A1(\MC_ARK_ARC_1_1/temp5[189] ), .A2(n1728), .Z(
        \MC_ARK_ARC_1_1/buf_output[189] ) );
  XOR2_X1 U5963 ( .A1(\MC_ARK_ARC_1_1/temp3[189] ), .A2(
        \MC_ARK_ARC_1_1/temp4[189] ), .Z(n1728) );
  XOR2_X1 U5964 ( .A1(\MC_ARK_ARC_1_0/temp1[90] ), .A2(
        \MC_ARK_ARC_1_0/temp2[90] ), .Z(n1729) );
  XOR2_X1 U5967 ( .A1(\MC_ARK_ARC_1_1/temp5[1] ), .A2(
        \MC_ARK_ARC_1_1/temp6[1] ), .Z(\MC_ARK_ARC_1_1/buf_output[1] ) );
  INV_X2 U5971 ( .I(\SB1_1_29/buf_output[3] ), .ZN(\SB2_1_27/i0[8] ) );
  XOR2_X1 U5975 ( .A1(n1732), .A2(\MC_ARK_ARC_1_2/temp5[142] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[142] ) );
  XOR2_X1 U5976 ( .A1(\MC_ARK_ARC_1_2/temp3[142] ), .A2(
        \MC_ARK_ARC_1_2/temp4[142] ), .Z(n1732) );
  XOR2_X1 U5977 ( .A1(\MC_ARK_ARC_1_0/temp6[13] ), .A2(
        \MC_ARK_ARC_1_0/temp5[13] ), .Z(\MC_ARK_ARC_1_0/buf_output[13] ) );
  NAND4_X2 U5978 ( .A1(\SB2_0_18/Component_Function_5/NAND4_in[1] ), .A2(n2662), .A3(\SB2_0_18/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_18/buf_output[5] ) );
  NAND3_X2 U5985 ( .A1(\SB1_3_14/i1_5 ), .A2(\SB1_3_14/i1[9] ), .A3(
        \SB1_3_14/i0_4 ), .ZN(\SB1_3_14/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U5989 ( .A1(\SB1_2_31/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_31/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_31/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_2_31/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_31/buf_output[1] ) );
  XOR2_X1 U5994 ( .A1(\SB2_0_26/buf_output[1] ), .A2(\RI5[0][61] ), .Z(n1733)
         );
  NAND4_X2 U5995 ( .A1(\SB1_4_11/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_4_11/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_4_11/Component_Function_3/NAND4_in[2] ), .A4(n1734), .ZN(
        \SB1_4_11/buf_output[3] ) );
  NAND3_X1 U5996 ( .A1(\SB2_1_7/i0_0 ), .A2(\SB2_1_7/i3[0] ), .A3(
        \SB2_1_7/i1_7 ), .ZN(\SB2_1_7/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U5999 ( .A1(\MC_ARK_ARC_1_0/temp6[163] ), .A2(n1736), .Z(
        \MC_ARK_ARC_1_0/buf_output[163] ) );
  XOR2_X1 U6000 ( .A1(\MC_ARK_ARC_1_0/temp1[163] ), .A2(
        \MC_ARK_ARC_1_0/temp2[163] ), .Z(n1736) );
  XOR2_X1 U6008 ( .A1(n1767), .A2(n1742), .Z(\MC_ARK_ARC_1_0/buf_output[80] )
         );
  XOR2_X1 U6009 ( .A1(n2702), .A2(\MC_ARK_ARC_1_0/temp4[80] ), .Z(n1742) );
  NAND3_X2 U6010 ( .A1(\SB3_17/i0_3 ), .A2(\SB3_17/i1[9] ), .A3(\SB3_17/i0_4 ), 
        .ZN(n1743) );
  XOR2_X1 U6013 ( .A1(n1745), .A2(\MC_ARK_ARC_1_3/temp4[8] ), .Z(
        \MC_ARK_ARC_1_3/temp6[8] ) );
  XOR2_X1 U6014 ( .A1(\SB2_3_22/buf_output[2] ), .A2(\RI5[3][110] ), .Z(n1745)
         );
  NAND4_X2 U6017 ( .A1(\SB1_4_8/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_4_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_8/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_4_8/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_4_8/buf_output[1] ) );
  XOR2_X1 U6021 ( .A1(\RI5[1][31] ), .A2(\RI5[1][67] ), .Z(
        \MC_ARK_ARC_1_1/temp3[157] ) );
  NAND3_X1 U6025 ( .A1(\SB2_0_8/i0[7] ), .A2(\SB2_0_8/i0[8] ), .A3(
        \SB2_0_8/i0[6] ), .ZN(\SB2_0_8/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U6030 ( .A1(\MC_ARK_ARC_1_2/temp5[97] ), .A2(n1752), .Z(
        \MC_ARK_ARC_1_2/buf_output[97] ) );
  XOR2_X1 U6031 ( .A1(\MC_ARK_ARC_1_2/temp4[97] ), .A2(
        \MC_ARK_ARC_1_2/temp3[97] ), .Z(n1752) );
  XOR2_X1 U6032 ( .A1(\MC_ARK_ARC_1_3/temp6[13] ), .A2(
        \MC_ARK_ARC_1_3/temp5[13] ), .Z(\MC_ARK_ARC_1_3/buf_output[13] ) );
  NAND3_X2 U6033 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0[6] ), .A3(
        \SB2_0_21/i0[10] ), .ZN(\SB2_0_21/Component_Function_2/NAND4_in[1] )
         );
  NAND4_X2 U6034 ( .A1(\SB1_0_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_20/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_20/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_20/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_0_20/buf_output[5] ) );
  INV_X2 U6035 ( .I(\SB1_4_0/buf_output[2] ), .ZN(\SB2_4_29/i1[9] ) );
  XOR2_X1 U6040 ( .A1(\MC_ARK_ARC_1_1/temp1[25] ), .A2(
        \MC_ARK_ARC_1_1/temp2[25] ), .Z(n1753) );
  NAND4_X2 U6047 ( .A1(n2500), .A2(n2501), .A3(n1759), .A4(
        \SB2_1_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_31/buf_output[5] ) );
  XOR2_X1 U6050 ( .A1(\MC_ARK_ARC_1_2/temp1[143] ), .A2(
        \MC_ARK_ARC_1_2/temp2[143] ), .Z(\MC_ARK_ARC_1_2/temp5[143] ) );
  NAND3_X1 U6052 ( .A1(\SB1_2_12/i1_7 ), .A2(\RI1[2][119] ), .A3(
        \SB1_2_12/i0[8] ), .ZN(\SB1_2_12/Component_Function_1/NAND4_in[1] ) );
  NOR2_X2 U6054 ( .A1(n2521), .A2(n2255), .ZN(n1763) );
  NAND3_X1 U6058 ( .A1(\SB2_1_1/i0_0 ), .A2(\SB2_1_1/i0_3 ), .A3(
        \SB2_1_1/i0[7] ), .ZN(\SB2_1_1/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U6060 ( .A1(n2703), .A2(\MC_ARK_ARC_1_0/temp3[80] ), .Z(n1767) );
  NAND3_X2 U6062 ( .A1(\SB1_1_19/i0[10] ), .A2(\SB1_1_19/i1[9] ), .A3(
        \SB1_1_19/i1_7 ), .ZN(\SB1_1_19/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U6064 ( .A1(\MC_ARK_ARC_1_2/temp5[122] ), .A2(
        \MC_ARK_ARC_1_2/temp6[122] ), .Z(\MC_ARK_ARC_1_2/buf_output[122] ) );
  XOR2_X1 U6072 ( .A1(\MC_ARK_ARC_1_0/temp3[130] ), .A2(
        \MC_ARK_ARC_1_0/temp4[130] ), .Z(\MC_ARK_ARC_1_0/temp6[130] ) );
  NAND3_X1 U6074 ( .A1(\SB2_1_5/i0[9] ), .A2(\SB2_1_5/i1_5 ), .A3(
        \SB2_1_5/i0[6] ), .ZN(n1769) );
  XOR2_X1 U6075 ( .A1(\RI5[1][181] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[187] ) );
  XOR2_X1 U6079 ( .A1(\RI5[2][125] ), .A2(\RI5[2][149] ), .Z(
        \MC_ARK_ARC_1_2/temp2[179] ) );
  NAND4_X2 U6080 ( .A1(\SB2_1_7/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_7/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_7/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_1_7/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_1_7/buf_output[0] ) );
  NAND4_X2 U6083 ( .A1(\SB3_4/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_4/Component_Function_4/NAND4_in[3] ), .A3(
        \SB3_4/Component_Function_4/NAND4_in[1] ), .A4(
        \SB3_4/Component_Function_4/NAND4_in[0] ), .ZN(\SB3_4/buf_output[4] )
         );
  NAND4_X2 U6084 ( .A1(\SB1_1_10/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_10/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_10/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_10/buf_output[0] ) );
  XOR2_X1 U6086 ( .A1(\SB2_1_14/buf_output[2] ), .A2(n156), .Z(n1773) );
  XOR2_X1 U6091 ( .A1(\MC_ARK_ARC_1_2/temp5[129] ), .A2(n1776), .Z(
        \MC_ARK_ARC_1_2/buf_output[129] ) );
  XOR2_X1 U6093 ( .A1(\RI5[0][95] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[71] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[125] ) );
  XOR2_X1 U6094 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[124] ), .A2(\RI5[2][160] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[58] ) );
  NAND4_X2 U6096 ( .A1(\SB1_2_2/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_2/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_2/Component_Function_0/NAND4_in[0] ), .A4(n1777), .ZN(
        \SB1_2_2/buf_output[0] ) );
  NAND4_X2 U6097 ( .A1(\SB1_4_11/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_4_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_11/Component_Function_1/NAND4_in[0] ), .A4(n1778), .ZN(
        \SB1_4_11/buf_output[1] ) );
  NAND4_X2 U6102 ( .A1(\SB3_21/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_21/Component_Function_1/NAND4_in[0] ), .A4(n1780), .ZN(
        \SB3_21/buf_output[1] ) );
  NAND3_X1 U6103 ( .A1(\SB3_21/i0_4 ), .A2(\SB3_21/i1_7 ), .A3(\SB3_21/i0[8] ), 
        .ZN(n1780) );
  NOR2_X2 U6105 ( .A1(n3034), .A2(n1782), .ZN(n3033) );
  XOR2_X1 U6112 ( .A1(n1786), .A2(\MC_ARK_ARC_1_4/temp4[122] ), .Z(n2537) );
  XOR2_X1 U6113 ( .A1(\RI5[4][32] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[188] ), 
        .Z(n1786) );
  XOR2_X1 U6115 ( .A1(\RI5[4][81] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[117] ), 
        .Z(n1788) );
  XOR2_X1 U6116 ( .A1(\MC_ARK_ARC_1_2/temp1[91] ), .A2(
        \MC_ARK_ARC_1_2/temp2[91] ), .Z(\MC_ARK_ARC_1_2/temp5[91] ) );
  NAND3_X1 U6120 ( .A1(\SB4_11/i0[8] ), .A2(\SB4_11/i3[0] ), .A3(\SB4_11/i1_5 ), .ZN(n1790) );
  NAND4_X2 U6128 ( .A1(\SB2_0_24/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_24/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_24/Component_Function_3/NAND4_in[0] ), .A4(n1794), .ZN(
        \SB2_0_24/buf_output[3] ) );
  BUF_X4 U6133 ( .I(\SB2_2_15/buf_output[0] ), .Z(\RI5[2][126] ) );
  NAND3_X1 U6140 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i0[9] ), .A3(\SB3_1/i0[8] ), 
        .ZN(n1800) );
  BUF_X4 U6141 ( .I(\SB2_4_12/buf_output[0] ), .Z(\RI5[4][144] ) );
  XOR2_X1 U6143 ( .A1(n1803), .A2(\MC_ARK_ARC_1_4/temp4[108] ), .Z(
        \MC_ARK_ARC_1_4/temp6[108] ) );
  XOR2_X1 U6145 ( .A1(n1804), .A2(\MC_ARK_ARC_1_1/temp4[162] ), .Z(
        \MC_ARK_ARC_1_1/temp6[162] ) );
  XOR2_X1 U6146 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[36] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[72] ), .Z(n1804) );
  NAND4_X2 U6147 ( .A1(\SB1_2_29/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_0/NAND4_in[0] ), .A4(n1805), .ZN(
        \SB1_2_29/buf_output[0] ) );
  NAND3_X1 U6149 ( .A1(\SB2_0_5/i0_4 ), .A2(\SB2_0_5/i0[8] ), .A3(
        \SB2_0_5/i1_7 ), .ZN(\SB2_0_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U6153 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i0[10] ), .A3(
        \SB1_1_8/buf_output[1] ), .ZN(n2619) );
  XOR2_X1 U6154 ( .A1(\MC_ARK_ARC_1_3/temp4[141] ), .A2(n1807), .Z(n2394) );
  XOR2_X1 U6155 ( .A1(\RI5[3][51] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[15] ), 
        .Z(n1807) );
  XOR2_X1 U6156 ( .A1(\RI5[0][100] ), .A2(\RI5[0][76] ), .Z(
        \MC_ARK_ARC_1_0/temp2[130] ) );
  NOR2_X2 U6160 ( .A1(n1811), .A2(n1809), .ZN(n2998) );
  NAND2_X1 U6161 ( .A1(\SB1_3_20/Component_Function_4/NAND4_in[3] ), .A2(n1810), .ZN(n1809) );
  NAND3_X1 U6162 ( .A1(\SB1_3_20/i0_0 ), .A2(\SB1_3_20/i3[0] ), .A3(
        \SB1_3_20/i1_7 ), .ZN(n1810) );
  NAND2_X1 U6163 ( .A1(\SB1_3_20/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_3_20/Component_Function_4/NAND4_in[0] ), .ZN(n1811) );
  XOR2_X1 U6166 ( .A1(\MC_ARK_ARC_1_1/temp2[175] ), .A2(n1813), .Z(n1968) );
  XOR2_X1 U6167 ( .A1(\RI5[1][169] ), .A2(\RI5[1][175] ), .Z(n1813) );
  XOR2_X1 U6168 ( .A1(\MC_ARK_ARC_1_0/temp5[116] ), .A2(n1814), .Z(
        \MC_ARK_ARC_1_0/buf_output[116] ) );
  XOR2_X1 U6169 ( .A1(\MC_ARK_ARC_1_0/temp5[128] ), .A2(n1815), .Z(
        \MC_ARK_ARC_1_0/buf_output[128] ) );
  XOR2_X1 U6170 ( .A1(\MC_ARK_ARC_1_0/temp3[128] ), .A2(
        \MC_ARK_ARC_1_0/temp4[128] ), .Z(n1815) );
  NAND2_X1 U6183 ( .A1(\SB1_0_29/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_29/Component_Function_4/NAND4_in[0] ), .ZN(n2321) );
  XOR2_X1 U6185 ( .A1(\RI5[3][23] ), .A2(\RI5[3][47] ), .Z(n1819) );
  NAND4_X2 U6188 ( .A1(\SB1_0_12/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_12/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_12/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][139] ) );
  NAND3_X1 U6189 ( .A1(\SB2_3_26/i1_7 ), .A2(\SB2_3_26/i0_4 ), .A3(
        \SB2_3_26/i0[8] ), .ZN(\SB2_3_26/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 U6197 ( .I(\SB2_2_13/buf_output[4] ), .Z(\RI5[2][118] ) );
  XOR2_X1 U6199 ( .A1(\SB2_1_11/buf_output[3] ), .A2(\RI5[1][99] ), .Z(
        \MC_ARK_ARC_1_1/temp3[33] ) );
  NAND4_X2 U6200 ( .A1(\SB2_2_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_28/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_28/Component_Function_1/NAND4_in[1] ), .A4(n2237), .ZN(
        \SB2_2_28/buf_output[1] ) );
  NAND4_X2 U6205 ( .A1(\SB1_3_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_7/Component_Function_4/NAND4_in[2] ), .A4(n1825), .ZN(
        \SB1_3_7/buf_output[4] ) );
  XOR2_X1 U6206 ( .A1(\MC_ARK_ARC_1_3/temp5[131] ), .A2(n1826), .Z(
        \MC_ARK_ARC_1_3/buf_output[131] ) );
  INV_X1 U6207 ( .I(\RI3[0][151] ), .ZN(\SB2_0_6/i1_7 ) );
  NAND4_X2 U6208 ( .A1(\SB1_0_10/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_0_10/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][151] ) );
  XOR2_X1 U6209 ( .A1(n1827), .A2(\MC_ARK_ARC_1_2/temp5[102] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[102] ) );
  XOR2_X1 U6210 ( .A1(\MC_ARK_ARC_1_2/temp4[102] ), .A2(
        \MC_ARK_ARC_1_2/temp3[102] ), .Z(n1827) );
  XOR2_X1 U6216 ( .A1(n1832), .A2(\MC_ARK_ARC_1_0/temp5[167] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[167] ) );
  XOR2_X1 U6217 ( .A1(\MC_ARK_ARC_1_0/temp3[167] ), .A2(
        \MC_ARK_ARC_1_0/temp4[167] ), .Z(n1832) );
  NAND4_X2 U6220 ( .A1(\SB1_3_13/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_3_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_13/buf_output[0] ) );
  XOR2_X1 U6228 ( .A1(\MC_ARK_ARC_1_4/temp3[154] ), .A2(
        \MC_ARK_ARC_1_4/temp4[154] ), .Z(\MC_ARK_ARC_1_4/temp6[154] ) );
  NAND4_X2 U6233 ( .A1(\SB2_1_24/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_24/Component_Function_2/NAND4_in[0] ), .A4(n1844), .ZN(
        \SB2_1_24/buf_output[2] ) );
  NAND4_X2 U6242 ( .A1(\SB2_0_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_0_19/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_0_19/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_19/buf_output[5] ) );
  NAND4_X2 U6244 ( .A1(\SB2_3_12/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_12/Component_Function_1/NAND4_in[0] ), .A4(n1845), .ZN(
        \SB2_3_12/buf_output[1] ) );
  NAND4_X2 U6246 ( .A1(\SB3_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_2/NAND4_in[3] ), .A3(
        \SB3_4/Component_Function_2/NAND4_in[2] ), .A4(n1846), .ZN(
        \SB3_4/buf_output[2] ) );
  XOR2_X1 U6251 ( .A1(n2433), .A2(n1848), .Z(\MC_ARK_ARC_1_3/temp5[100] ) );
  XOR2_X1 U6252 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[94] ), .A2(\RI5[3][100] ), 
        .Z(n1848) );
  NAND4_X2 U6253 ( .A1(\SB2_4_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_4_15/Component_Function_4/NAND4_in[3] ), .A4(n1849), .ZN(
        \SB2_4_15/buf_output[4] ) );
  XOR2_X1 U6256 ( .A1(\RI5[0][100] ), .A2(\RI5[0][106] ), .Z(
        \MC_ARK_ARC_1_0/temp1[106] ) );
  XOR2_X1 U6258 ( .A1(\RI5[2][69] ), .A2(\RI5[2][75] ), .Z(n1851) );
  NAND3_X2 U6260 ( .A1(\SB2_3_17/i3[0] ), .A2(\SB2_3_17/i1_5 ), .A3(
        \SB2_3_17/i0[8] ), .ZN(n1933) );
  NAND4_X2 U6261 ( .A1(\SB2_0_20/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_20/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_20/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_0_20/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_0_20/buf_output[4] ) );
  NAND3_X1 U6267 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0[10] ), .A3(
        \SB1_1_22/i0_4 ), .ZN(\SB1_1_22/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U6270 ( .A1(\SB2_3_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_25/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_3_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_25/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_25/buf_output[1] ) );
  NAND3_X2 U6280 ( .A1(\SB2_1_20/i0[8] ), .A2(\SB2_1_20/i3[0] ), .A3(
        \SB2_1_20/i1_5 ), .ZN(n2070) );
  BUF_X4 U6282 ( .I(\SB2_2_4/buf_output[2] ), .Z(\RI5[2][182] ) );
  NAND3_X1 U6285 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i0_3 ), .A3(\SB4_14/i0[7] ), 
        .ZN(\SB4_14/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U6289 ( .A1(\MC_ARK_ARC_1_1/temp5[126] ), .A2(
        \MC_ARK_ARC_1_1/temp6[126] ), .Z(\MC_ARK_ARC_1_1/buf_output[126] ) );
  XOR2_X1 U6299 ( .A1(\MC_ARK_ARC_1_2/temp2[94] ), .A2(
        \MC_ARK_ARC_1_2/temp1[94] ), .Z(n2367) );
  NAND3_X1 U6300 ( .A1(\SB1_3_14/i0[6] ), .A2(\SB1_3_14/i0[8] ), .A3(
        \SB1_3_14/i0[7] ), .ZN(\SB1_3_14/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U6304 ( .A1(\SB1_3_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_3/Component_Function_1/NAND4_in[3] ), .A4(n1868), .ZN(
        \SB1_3_3/buf_output[1] ) );
  NAND4_X2 U6307 ( .A1(\SB1_3_3/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_3/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_3_3/Component_Function_0/NAND4_in[0] ), .A4(n1870), .ZN(
        \SB1_3_3/buf_output[0] ) );
  NAND4_X2 U6308 ( .A1(\SB2_0_19/Component_Function_0/NAND4_in[1] ), .A2(n1871), .A3(n2736), .A4(\SB2_0_19/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_19/buf_output[0] ) );
  NAND3_X2 U6310 ( .A1(\SB2_0_8/i0_3 ), .A2(\RI3[0][142] ), .A3(
        \SB2_0_8/i1[9] ), .ZN(n2096) );
  NAND3_X1 U6311 ( .A1(\SB2_2_5/i0_0 ), .A2(\SB2_2_5/i0[7] ), .A3(
        \SB2_2_5/i0_3 ), .ZN(\SB2_2_5/Component_Function_0/NAND4_in[3] ) );
  OR3_X1 U6312 ( .A1(\RI3[0][93] ), .A2(n5157), .A3(\RI3[0][95] ), .Z(
        \SB2_0_16/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U6313 ( .A1(n1873), .A2(n1874), .Z(\MC_ARK_ARC_1_0/temp6[87] ) );
  XOR2_X1 U6314 ( .A1(\RI5[0][123] ), .A2(n152), .Z(n1873) );
  XOR2_X1 U6315 ( .A1(\RI5[0][153] ), .A2(\RI5[0][189] ), .Z(n1874) );
  XOR2_X1 U6319 ( .A1(n2377), .A2(n1877), .Z(\MC_ARK_ARC_1_2/buf_output[24] )
         );
  XOR2_X1 U6321 ( .A1(\MC_ARK_ARC_1_3/temp4[125] ), .A2(
        \MC_ARK_ARC_1_3/temp3[125] ), .Z(n1879) );
  XOR2_X1 U6325 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[112] ), .A2(\RI5[2][136] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[166] ) );
  NAND4_X2 U6329 ( .A1(\SB2_2_14/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_14/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_14/Component_Function_4/NAND4_in[2] ), .A4(n1884), .ZN(
        \SB2_2_14/buf_output[4] ) );
  NAND3_X1 U6330 ( .A1(\SB2_2_14/i0_4 ), .A2(\SB2_2_14/i1[9] ), .A3(
        \SB2_2_14/i1_5 ), .ZN(n1884) );
  XOR2_X1 U6340 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[29] ), .A2(\RI5[3][59] ), 
        .Z(n1890) );
  BUF_X4 U6346 ( .I(\SB2_0_20/buf_output[0] ), .Z(\RI5[0][96] ) );
  XOR2_X1 U6347 ( .A1(n2048), .A2(n1893), .Z(\MC_ARK_ARC_1_0/buf_output[9] )
         );
  BUF_X4 U6349 ( .I(\SB2_1_24/buf_output[1] ), .Z(\RI5[1][67] ) );
  NAND4_X2 U6353 ( .A1(\SB2_1_22/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_22/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_22/Component_Function_0/NAND4_in[0] ), .A4(n1896), .ZN(
        \SB2_1_22/buf_output[0] ) );
  XOR2_X1 U6354 ( .A1(n2423), .A2(\MC_ARK_ARC_1_4/temp1[139] ), .Z(n2153) );
  OAI21_X1 U6357 ( .A1(n1898), .A2(\SB2_1_1/i1[9] ), .B(\SB2_1_1/i0_3 ), .ZN(
        n2612) );
  NAND3_X1 U6364 ( .A1(\SB4_27/i0_0 ), .A2(\SB4_27/i0[8] ), .A3(\SB4_27/i0[9] ), .ZN(n1903) );
  XOR2_X1 U6373 ( .A1(n1908), .A2(n2446), .Z(\MC_ARK_ARC_1_0/buf_output[31] )
         );
  XOR2_X1 U6374 ( .A1(\MC_ARK_ARC_1_0/temp2[31] ), .A2(
        \MC_ARK_ARC_1_0/temp1[31] ), .Z(n1908) );
  XOR2_X1 U6375 ( .A1(\RI5[2][64] ), .A2(\RI5[2][88] ), .Z(
        \MC_ARK_ARC_1_2/temp2[118] ) );
  NAND3_X1 U6379 ( .A1(\SB2_4_15/i0_3 ), .A2(\SB2_4_15/i0_0 ), .A3(
        \SB2_4_15/i0[7] ), .ZN(n2258) );
  XOR2_X1 U6381 ( .A1(\MC_ARK_ARC_1_1/temp2[51] ), .A2(
        \MC_ARK_ARC_1_1/temp1[51] ), .Z(n1910) );
  NAND4_X2 U6384 ( .A1(\SB1_0_28/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_28/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_28/Component_Function_5/NAND4_in[0] ), .A4(n1912), .ZN(
        \SB1_0_28/buf_output[5] ) );
  NAND3_X1 U6385 ( .A1(n5433), .A2(\SB1_0_28/i0[9] ), .A3(n224), .ZN(n1912) );
  NAND4_X2 U6389 ( .A1(\SB1_2_23/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_1/NAND4_in[0] ), .A4(n1915), .ZN(
        \SB1_2_23/buf_output[1] ) );
  XOR2_X1 U6395 ( .A1(n2495), .A2(\MC_ARK_ARC_1_2/temp2[7] ), .Z(n1919) );
  NAND3_X1 U6398 ( .A1(\SB4_26/i0[6] ), .A2(\SB4_26/i1_5 ), .A3(\SB4_26/i0[9] ), .ZN(\SB4_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U6407 ( .A1(\SB1_0_20/i0[10] ), .A2(\SB1_0_20/i1[9] ), .A3(
        \SB1_0_20/i1_5 ), .ZN(\SB1_0_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U6409 ( .A1(\SB2_1_0/i0_3 ), .A2(\SB2_1_0/i0[9] ), .A3(
        \SB2_1_0/i0[8] ), .ZN(\SB2_1_0/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U6418 ( .A1(n3003), .A2(n1930), .Z(\MC_ARK_ARC_1_4/buf_output[2] )
         );
  XOR2_X1 U6422 ( .A1(\MC_ARK_ARC_1_3/temp2[105] ), .A2(n1932), .Z(
        \MC_ARK_ARC_1_3/temp5[105] ) );
  XOR2_X1 U6423 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[99] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[105] ), .Z(n1932) );
  INV_X1 U6427 ( .I(\SB3_27/buf_output[5] ), .ZN(\SB4_27/i1_5 ) );
  NAND4_X2 U6433 ( .A1(\SB2_4_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_4_21/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_4_21/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_4_21/buf_output[3] ) );
  XOR2_X1 U6439 ( .A1(n1942), .A2(\MC_ARK_ARC_1_3/temp4[43] ), .Z(
        \MC_ARK_ARC_1_3/temp6[43] ) );
  XOR2_X1 U6440 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[109] ), .A2(\RI5[3][145] ), 
        .Z(n1942) );
  NAND3_X1 U6441 ( .A1(\SB2_4_20/i0_3 ), .A2(\SB2_4_20/i0[6] ), .A3(
        \SB2_4_20/i1[9] ), .ZN(\SB2_4_20/Component_Function_3/NAND4_in[0] ) );
  INV_X4 U6444 ( .I(n2998), .ZN(\SB1_3_20/buf_output[4] ) );
  XOR2_X1 U6447 ( .A1(\MC_ARK_ARC_1_1/temp5[30] ), .A2(
        \MC_ARK_ARC_1_1/temp6[30] ), .Z(\MC_ARK_ARC_1_1/buf_output[30] ) );
  XOR2_X1 U6452 ( .A1(n1946), .A2(\MC_ARK_ARC_1_2/temp5[177] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[177] ) );
  XOR2_X1 U6453 ( .A1(\MC_ARK_ARC_1_2/temp3[177] ), .A2(
        \MC_ARK_ARC_1_2/temp4[177] ), .Z(n1946) );
  XOR2_X1 U6455 ( .A1(\MC_ARK_ARC_1_2/temp3[55] ), .A2(
        \MC_ARK_ARC_1_2/temp4[55] ), .Z(n1949) );
  NAND4_X2 U6456 ( .A1(\SB2_1_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_30/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_30/Component_Function_1/NAND4_in[0] ), .A4(n1950), .ZN(
        \SB2_1_30/buf_output[1] ) );
  XOR2_X1 U6459 ( .A1(\MC_ARK_ARC_1_1/temp1[31] ), .A2(
        \MC_ARK_ARC_1_1/temp4[31] ), .Z(n1952) );
  INV_X4 U6462 ( .I(n1953), .ZN(\SB1_3_10/buf_output[4] ) );
  BUF_X4 U6464 ( .I(\SB2_2_13/buf_output[2] ), .Z(\RI5[2][128] ) );
  XOR2_X1 U6470 ( .A1(n3123), .A2(n1957), .Z(\MC_ARK_ARC_1_0/buf_output[125] )
         );
  XOR2_X1 U6472 ( .A1(\MC_ARK_ARC_1_2/temp2[85] ), .A2(n2281), .Z(
        \MC_ARK_ARC_1_2/temp5[85] ) );
  NAND4_X2 U6473 ( .A1(\SB2_2_22/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_22/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_2_22/Component_Function_1/NAND4_in[1] ), .A4(n1959), .ZN(
        \SB2_2_22/buf_output[1] ) );
  NAND3_X2 U6478 ( .A1(\SB2_1_1/i0_4 ), .A2(\SB2_1_1/i0_3 ), .A3(
        \SB2_1_1/i1[9] ), .ZN(n1963) );
  NAND4_X2 U6484 ( .A1(\SB2_2_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_25/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_25/Component_Function_2/NAND4_in[2] ), .A4(n1965), .ZN(
        \SB2_2_25/buf_output[2] ) );
  NAND3_X1 U6486 ( .A1(\SB1_3_7/i0_0 ), .A2(\SB1_3_7/i3[0] ), .A3(
        \SB1_3_7/i1_7 ), .ZN(\SB1_3_7/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U6490 ( .A1(\RI5[1][85] ), .A2(\RI5[1][121] ), .Z(
        \MC_ARK_ARC_1_1/temp3[19] ) );
  NAND3_X2 U6495 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0[9] ), .A3(
        \SB2_3_18/i0[8] ), .ZN(n1972) );
  XOR2_X1 U6497 ( .A1(\MC_ARK_ARC_1_0/temp4[120] ), .A2(
        \MC_ARK_ARC_1_0/temp3[120] ), .Z(\MC_ARK_ARC_1_0/temp6[120] ) );
  XOR2_X1 U6499 ( .A1(\MC_ARK_ARC_1_0/temp5[105] ), .A2(n1973), .Z(
        \MC_ARK_ARC_1_0/buf_output[105] ) );
  NAND3_X2 U6501 ( .A1(\RI1[4][191] ), .A2(\SB1_4_0/i1[9] ), .A3(
        \SB1_4_0/i0_4 ), .ZN(\SB1_4_0/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U6503 ( .A1(n1974), .A2(\MC_ARK_ARC_1_2/temp1[161] ), .Z(
        \MC_ARK_ARC_1_2/temp5[161] ) );
  XOR2_X1 U6504 ( .A1(\RI5[2][107] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .Z(n1974) );
  NAND3_X1 U6514 ( .A1(\SB1_1_21/i1_7 ), .A2(\SB1_1_21/i0_0 ), .A3(
        \SB1_1_21/i3[0] ), .ZN(\SB1_1_21/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U6517 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[43] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[7] ), .Z(\MC_ARK_ARC_1_3/temp3[133] ) );
  XOR2_X1 U6524 ( .A1(\RI5[3][38] ), .A2(\RI5[3][2] ), .Z(
        \MC_ARK_ARC_1_3/temp3[128] ) );
  NAND3_X1 U6527 ( .A1(\SB1_2_1/i0[6] ), .A2(\SB1_2_1/i1[9] ), .A3(
        \SB1_2_1/i0_3 ), .ZN(\SB1_2_1/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U6529 ( .A1(\RI5[2][166] ), .A2(\RI5[2][190] ), .Z(n1980) );
  XOR2_X1 U6531 ( .A1(\MC_ARK_ARC_1_4/temp6[81] ), .A2(n1982), .Z(
        \MC_ARK_ARC_1_4/buf_output[81] ) );
  XOR2_X1 U6532 ( .A1(\MC_ARK_ARC_1_4/temp2[81] ), .A2(n2910), .Z(n1982) );
  NAND2_X2 U6537 ( .A1(\SB2_1_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_4/NAND4_in[2] ), .ZN(n2945) );
  XOR2_X1 U6538 ( .A1(\MC_ARK_ARC_1_2/temp3[66] ), .A2(
        \MC_ARK_ARC_1_2/temp4[66] ), .Z(n2893) );
  NOR2_X2 U6541 ( .A1(n1986), .A2(n1984), .ZN(n2592) );
  NAND3_X2 U6542 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0[10] ), .A3(
        \SB1_0_6/i0_4 ), .ZN(n1985) );
  NAND4_X2 U6544 ( .A1(\SB2_3_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_8/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_8/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_3_8/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_3_8/buf_output[4] ) );
  BUF_X4 U6545 ( .I(\SB2_2_4/buf_output[1] ), .Z(\RI5[2][187] ) );
  XOR2_X1 U6547 ( .A1(\MC_ARK_ARC_1_3/temp5[49] ), .A2(
        \MC_ARK_ARC_1_3/temp6[49] ), .Z(\MC_ARK_ARC_1_3/buf_output[49] ) );
  NAND4_X2 U6551 ( .A1(\SB2_1_14/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_14/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_14/Component_Function_4/NAND4_in[1] ), .A4(n1991), .ZN(
        \SB2_1_14/buf_output[4] ) );
  NAND3_X1 U6554 ( .A1(\SB2_3_18/i0[6] ), .A2(\SB2_3_18/i0[9] ), .A3(
        \SB2_3_18/i1_5 ), .ZN(\SB2_3_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U6555 ( .A1(\SB2_0_8/i0[8] ), .A2(\RI3[0][142] ), .A3(
        \SB2_0_8/i1_7 ), .ZN(\SB2_0_8/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U6557 ( .A1(\RI5[0][44] ), .A2(n426), .Z(n1993) );
  XOR2_X1 U6558 ( .A1(\RI5[0][8] ), .A2(\RI5[0][170] ), .Z(n1994) );
  NAND3_X1 U6559 ( .A1(\SB1_3_22/i0_3 ), .A2(\SB1_3_22/i0[8] ), .A3(
        \SB1_3_22/i1_7 ), .ZN(\SB1_3_22/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U6561 ( .A1(\SB1_0_2/i0_0 ), .A2(\SB1_0_2/i0[10] ), .A3(
        \SB1_0_2/i0[6] ), .ZN(\SB1_0_2/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U6562 ( .A1(\SB2_3_15/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_15/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_15/Component_Function_4/NAND4_in[1] ), .A4(n1995), .ZN(
        \SB2_3_15/buf_output[4] ) );
  NAND3_X2 U6563 ( .A1(\SB2_0_20/i0_3 ), .A2(\SB2_0_20/i0[10] ), .A3(
        \RI3[0][70] ), .ZN(\SB2_0_20/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U6566 ( .A1(\MC_ARK_ARC_1_3/temp3[67] ), .A2(
        \MC_ARK_ARC_1_3/temp2[67] ), .Z(n1997) );
  NAND3_X1 U6569 ( .A1(\SB1_1_24/i0[6] ), .A2(\SB1_1_24/i1[9] ), .A3(
        \RI1[1][47] ), .ZN(\SB1_1_24/Component_Function_3/NAND4_in[0] ) );
  AND2_X1 U6572 ( .A1(\SB2_4_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_6/Component_Function_1/NAND4_in[3] ), .Z(n2001) );
  XOR2_X1 U6575 ( .A1(n2003), .A2(n2762), .Z(\MC_ARK_ARC_1_3/buf_output[54] )
         );
  NAND4_X2 U6590 ( .A1(\SB1_4_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_4_11/Component_Function_4/NAND4_in[2] ), .A4(n2009), .ZN(
        \SB1_4_11/buf_output[4] ) );
  NAND3_X2 U6593 ( .A1(\SB2_2_20/i0[6] ), .A2(\SB2_2_20/i0[9] ), .A3(
        \SB2_2_20/i0_4 ), .ZN(\SB2_2_20/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U6594 ( .A1(\RI5[3][38] ), .A2(\RI5[3][44] ), .Z(
        \MC_ARK_ARC_1_3/temp1[44] ) );
  NAND3_X2 U6596 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i0_4 ), .A3(
        \SB2_1_30/i1[9] ), .ZN(n3080) );
  NAND4_X2 U6600 ( .A1(\SB2_2_20/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_20/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_20/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_20/buf_output[1] ) );
  BUF_X4 U6604 ( .I(\SB2_2_9/buf_output[2] ), .Z(\RI5[2][152] ) );
  NAND3_X2 U6606 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i1[9] ), .A3(\SB3_2/i0_4 ), 
        .ZN(n2018) );
  NAND3_X1 U6607 ( .A1(\SB1_4_5/i0[8] ), .A2(\SB1_4_5/i1_5 ), .A3(
        \SB1_4_5/i3[0] ), .ZN(\SB1_4_5/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U6614 ( .A1(\MC_ARK_ARC_1_2/temp1[38] ), .A2(
        \MC_ARK_ARC_1_2/temp4[38] ), .Z(n2119) );
  NAND3_X1 U6615 ( .A1(\SB3_25/i0_0 ), .A2(\SB3_25/i0[9] ), .A3(\SB3_25/i0[8] ), .ZN(\SB3_25/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U6620 ( .A1(\RI5[1][181] ), .A2(\RI5[1][13] ), .Z(
        \MC_ARK_ARC_1_1/temp2[43] ) );
  XOR2_X1 U6623 ( .A1(n2976), .A2(\MC_ARK_ARC_1_4/temp6[38] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[38] ) );
  NAND3_X2 U6625 ( .A1(\SB1_1_24/i1_5 ), .A2(\SB1_1_24/i1[9] ), .A3(
        \SB1_1_24/i0_4 ), .ZN(n2022) );
  XOR2_X1 U6628 ( .A1(\MC_ARK_ARC_1_4/temp1[16] ), .A2(
        \MC_ARK_ARC_1_4/temp2[16] ), .Z(\MC_ARK_ARC_1_4/temp5[16] ) );
  XOR2_X1 U6636 ( .A1(\MC_ARK_ARC_1_4/temp2[37] ), .A2(
        \MC_ARK_ARC_1_4/temp1[37] ), .Z(\MC_ARK_ARC_1_4/temp5[37] ) );
  XOR2_X1 U6638 ( .A1(\MC_ARK_ARC_1_4/temp3[150] ), .A2(
        \MC_ARK_ARC_1_4/temp4[150] ), .Z(\MC_ARK_ARC_1_4/temp6[150] ) );
  NAND4_X2 U6645 ( .A1(\SB1_3_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_27/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_3_27/Component_Function_1/NAND4_in[0] ), .A4(n2030), .ZN(
        \SB1_3_27/buf_output[1] ) );
  XOR2_X1 U6646 ( .A1(\MC_ARK_ARC_1_1/temp2[64] ), .A2(
        \MC_ARK_ARC_1_1/temp1[64] ), .Z(\MC_ARK_ARC_1_1/temp5[64] ) );
  INV_X2 U6647 ( .I(\SB1_4_22/buf_output[3] ), .ZN(\SB2_4_20/i0[8] ) );
  XOR2_X1 U6651 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[120] ), .A2(\RI5[2][156] ), 
        .Z(n2031) );
  XOR2_X1 U6652 ( .A1(\MC_ARK_ARC_1_3/temp6[133] ), .A2(n2032), .Z(
        \MC_ARK_ARC_1_3/buf_output[133] ) );
  XOR2_X1 U6653 ( .A1(\MC_ARK_ARC_1_3/temp2[133] ), .A2(
        \MC_ARK_ARC_1_3/temp1[133] ), .Z(n2032) );
  XOR2_X1 U6654 ( .A1(\RI5[0][82] ), .A2(\RI5[0][118] ), .Z(
        \MC_ARK_ARC_1_0/temp3[16] ) );
  INV_X1 U6656 ( .I(\SB3_29/buf_output[0] ), .ZN(\SB4_24/i3[0] ) );
  NAND4_X2 U6657 ( .A1(\SB3_29/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_29/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_29/Component_Function_0/NAND4_in[1] ), .A4(
        \SB3_29/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_29/buf_output[0] ) );
  XOR2_X1 U6663 ( .A1(\RI5[4][32] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[170] ), 
        .Z(n2037) );
  XOR2_X1 U6664 ( .A1(\RI5[0][127] ), .A2(\RI5[0][163] ), .Z(
        \MC_ARK_ARC_1_0/temp3[61] ) );
  NAND4_X2 U6669 ( .A1(\SB2_4_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_6/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_4_6/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_4_6/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_4_6/buf_output[2] ) );
  XOR2_X1 U6680 ( .A1(n2206), .A2(\MC_ARK_ARC_1_0/temp4[9] ), .Z(n2048) );
  NAND3_X1 U6686 ( .A1(\SB2_1_3/i0_4 ), .A2(\SB2_1_3/i0[10] ), .A3(
        \SB2_1_3/i0_3 ), .ZN(\SB2_1_3/Component_Function_0/NAND4_in[2] ) );
  INV_X2 U6688 ( .I(\RI3[1][152] ), .ZN(\SB2_1_6/i1[9] ) );
  XOR2_X1 U6691 ( .A1(n2053), .A2(\MC_ARK_ARC_1_0/temp6[6] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[6] ) );
  XOR2_X1 U6692 ( .A1(\MC_ARK_ARC_1_0/temp2[6] ), .A2(
        \MC_ARK_ARC_1_0/temp1[6] ), .Z(n2053) );
  NAND4_X2 U6693 ( .A1(\SB1_2_12/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_12/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_12/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_2_12/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_2_12/buf_output[0] ) );
  XOR2_X1 U6696 ( .A1(\RI5[3][84] ), .A2(\RI5[3][132] ), .Z(n2054) );
  XOR2_X1 U6697 ( .A1(\RI5[3][138] ), .A2(\RI5[3][108] ), .Z(n2055) );
  NAND3_X2 U6702 ( .A1(\SB2_1_10/i0[6] ), .A2(\SB2_1_10/i0[9] ), .A3(
        \SB2_1_10/i0_4 ), .ZN(n2059) );
  NAND3_X1 U6703 ( .A1(\SB1_3_20/i0[10] ), .A2(\SB1_3_20/i0[9] ), .A3(
        \SB1_3_20/i0_3 ), .ZN(\SB1_3_20/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U6705 ( .A1(n2060), .A2(\MC_ARK_ARC_1_2/temp5[69] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[69] ) );
  XOR2_X1 U6706 ( .A1(\MC_ARK_ARC_1_2/temp3[69] ), .A2(
        \MC_ARK_ARC_1_2/temp4[69] ), .Z(n2060) );
  NAND4_X2 U6707 ( .A1(\SB2_3_18/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_18/Component_Function_0/NAND4_in[0] ), .A4(n2061), .ZN(
        \SB2_3_18/buf_output[0] ) );
  XOR2_X1 U6709 ( .A1(\MC_ARK_ARC_1_2/temp3[17] ), .A2(n2063), .Z(n2372) );
  XOR2_X1 U6710 ( .A1(\RI5[2][53] ), .A2(n436), .Z(n2063) );
  NOR2_X2 U6711 ( .A1(n2066), .A2(n2064), .ZN(n2978) );
  NAND2_X1 U6714 ( .A1(\SB1_0_26/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_26/Component_Function_4/NAND4_in[3] ), .ZN(n2066) );
  NAND4_X2 U6715 ( .A1(\SB3_8/Component_Function_5/NAND4_in[1] ), .A2(n2353), 
        .A3(\SB3_8/Component_Function_5/NAND4_in[2] ), .A4(n2067), .ZN(
        \SB3_8/buf_output[5] ) );
  NAND3_X2 U6717 ( .A1(\SB2_1_27/i0[10] ), .A2(\RI3[1][26] ), .A3(
        \SB2_1_27/i0[6] ), .ZN(\SB2_1_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U6718 ( .A1(\SB4_15/i0_4 ), .A2(\SB4_15/i1_7 ), .A3(n1497), .ZN(
        n2069) );
  NAND4_X2 U6727 ( .A1(\SB1_0_11/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_11/Component_Function_0/NAND4_in[2] ), .A4(n2076), .ZN(
        \RI3[0][150] ) );
  NAND2_X1 U6728 ( .A1(\SB1_0_11/i0[9] ), .A2(\SB1_0_11/i0[10] ), .ZN(n2076)
         );
  NAND4_X2 U6731 ( .A1(\SB1_4_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_4_5/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_4_5/Component_Function_2/NAND4_in[3] ), .A4(n2078), .ZN(
        \SB1_4_5/buf_output[2] ) );
  NAND3_X1 U6732 ( .A1(\SB1_0_6/i1[9] ), .A2(\SB1_0_6/i0[10] ), .A3(
        \SB1_0_6/i1_5 ), .ZN(n2079) );
  XOR2_X1 U6734 ( .A1(\RI5[4][8] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[2] ), 
        .Z(n2080) );
  XOR2_X1 U6736 ( .A1(\RI5[3][186] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[0] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[0] ) );
  NAND3_X1 U6737 ( .A1(\SB1_1_18/i0[6] ), .A2(\SB1_1_18/i0_3 ), .A3(
        \SB1_1_18/i0[10] ), .ZN(\SB1_1_18/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U6740 ( .A1(\MC_ARK_ARC_1_2/temp1[123] ), .A2(
        \MC_ARK_ARC_1_2/temp4[123] ), .Z(n2082) );
  XOR2_X1 U6742 ( .A1(\RI5[0][15] ), .A2(\RI5[0][183] ), .Z(
        \MC_ARK_ARC_1_0/temp2[45] ) );
  INV_X1 U6743 ( .I(\SB1_1_21/buf_output[0] ), .ZN(\SB2_1_16/i3[0] ) );
  NAND4_X2 U6744 ( .A1(\SB1_1_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_21/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_1_21/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_21/buf_output[0] ) );
  NAND3_X1 U6745 ( .A1(\SB1_1_24/i0[8] ), .A2(\SB1_1_24/i1_7 ), .A3(
        \RI1[1][47] ), .ZN(\SB1_1_24/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U6749 ( .A1(\MC_ARK_ARC_1_2/temp1[17] ), .A2(n2085), .Z(
        \MC_ARK_ARC_1_2/temp5[17] ) );
  XOR2_X1 U6750 ( .A1(\RI5[2][155] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[179] ), 
        .Z(n2085) );
  NAND4_X2 U6754 ( .A1(\SB1_0_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_25/Component_Function_5/NAND4_in[3] ), .A3(n2294), .A4(
        \SB1_0_25/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][41] ) );
  NAND3_X1 U6757 ( .A1(\SB2_3_1/i0[8] ), .A2(\SB2_3_1/i3[0] ), .A3(
        \SB2_3_1/i1_5 ), .ZN(\SB2_3_1/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U6759 ( .A1(\RI5[2][161] ), .A2(\RI5[2][155] ), .Z(
        \MC_ARK_ARC_1_2/temp1[161] ) );
  XOR2_X1 U6762 ( .A1(\MC_ARK_ARC_1_3/temp5[97] ), .A2(
        \MC_ARK_ARC_1_3/temp6[97] ), .Z(\MC_ARK_ARC_1_3/buf_output[97] ) );
  XOR2_X1 U6764 ( .A1(\MC_ARK_ARC_1_2/temp3[135] ), .A2(
        \MC_ARK_ARC_1_2/temp4[135] ), .Z(n2227) );
  NAND4_X2 U6768 ( .A1(\SB1_0_18/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_18/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_0_18/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_18/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_18/buf_output[0] ) );
  XOR2_X1 U6769 ( .A1(\RI5[3][148] ), .A2(\RI5[3][154] ), .Z(n2088) );
  XOR2_X1 U6773 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[165] ), .A2(\RI5[4][189] ), 
        .Z(n2091) );
  XOR2_X1 U6775 ( .A1(\MC_ARK_ARC_1_3/temp5[64] ), .A2(n2093), .Z(
        \MC_ARK_ARC_1_3/buf_output[64] ) );
  XOR2_X1 U6776 ( .A1(\MC_ARK_ARC_1_3/temp4[64] ), .A2(
        \MC_ARK_ARC_1_3/temp3[64] ), .Z(n2093) );
  XOR2_X1 U6777 ( .A1(\MC_ARK_ARC_1_4/temp5[63] ), .A2(n2094), .Z(
        \MC_ARK_ARC_1_4/buf_output[63] ) );
  XOR2_X1 U6778 ( .A1(\MC_ARK_ARC_1_4/temp3[63] ), .A2(
        \MC_ARK_ARC_1_4/temp4[63] ), .Z(n2094) );
  BUF_X4 U6781 ( .I(\SB2_2_12/buf_output[1] ), .Z(\RI5[2][139] ) );
  NAND4_X2 U6785 ( .A1(\SB2_1_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_2/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_1_2/Component_Function_3/NAND4_in[0] ), .A4(n2098), .ZN(
        \SB2_1_2/buf_output[3] ) );
  INV_X2 U6790 ( .I(\SB1_3_14/buf_output[3] ), .ZN(\SB2_3_12/i0[8] ) );
  NAND3_X1 U6791 ( .A1(\SB1_4_6/i0[8] ), .A2(\RI1[4][155] ), .A3(
        \SB1_4_6/i1_7 ), .ZN(\SB1_4_6/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U6795 ( .A1(\MC_ARK_ARC_1_1/temp4[175] ), .A2(
        \MC_ARK_ARC_1_1/temp3[175] ), .Z(\MC_ARK_ARC_1_1/temp6[175] ) );
  NAND4_X2 U6796 ( .A1(\SB2_2_1/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_1/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_2_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_1/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_1/buf_output[0] ) );
  XOR2_X1 U6799 ( .A1(n2103), .A2(\MC_ARK_ARC_1_4/temp6[39] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[39] ) );
  XOR2_X1 U6808 ( .A1(\MC_ARK_ARC_1_0/temp5[156] ), .A2(n2189), .Z(
        \MC_ARK_ARC_1_0/buf_output[156] ) );
  NAND3_X1 U6809 ( .A1(\SB1_3_10/i0[8] ), .A2(\SB1_3_10/i0_4 ), .A3(
        \SB1_3_10/i1_7 ), .ZN(\SB1_3_10/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U6813 ( .A1(\MC_ARK_ARC_1_0/temp6[62] ), .A2(
        \MC_ARK_ARC_1_0/temp5[62] ), .Z(\MC_ARK_ARC_1_0/buf_output[62] ) );
  XOR2_X1 U6815 ( .A1(n2110), .A2(\MC_ARK_ARC_1_0/temp4[98] ), .Z(
        \MC_ARK_ARC_1_0/temp6[98] ) );
  XOR2_X1 U6816 ( .A1(\RI5[0][8] ), .A2(\RI5[0][164] ), .Z(n2110) );
  XOR2_X1 U6817 ( .A1(\RI5[4][158] ), .A2(\RI5[4][164] ), .Z(
        \MC_ARK_ARC_1_4/temp1[164] ) );
  NOR2_X2 U6818 ( .A1(n2444), .A2(n2111), .ZN(n2748) );
  NAND3_X2 U6828 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i1[9] ), .A3(
        \SB1_1_8/buf_output[1] ), .ZN(n2815) );
  XOR2_X1 U6831 ( .A1(\RI5[2][125] ), .A2(n136), .Z(n2117) );
  XOR2_X1 U6834 ( .A1(n2120), .A2(n2119), .Z(\MC_ARK_ARC_1_2/buf_output[38] )
         );
  INV_X4 U6844 ( .I(n3104), .ZN(\SB1_2_22/buf_output[4] ) );
  NAND3_X2 U6845 ( .A1(\SB2_3_27/i0[6] ), .A2(\SB2_3_27/i0_3 ), .A3(
        \SB2_3_27/i0[10] ), .ZN(\SB2_3_27/Component_Function_2/NAND4_in[1] )
         );
  BUF_X4 U6849 ( .I(\SB2_2_24/buf_output[1] ), .Z(\RI5[2][67] ) );
  XOR2_X1 U6851 ( .A1(n2128), .A2(\MC_ARK_ARC_1_3/temp4[175] ), .Z(
        \MC_ARK_ARC_1_3/temp6[175] ) );
  INV_X2 U6853 ( .I(\SB1_2_17/buf_output[3] ), .ZN(\SB2_2_15/i0[8] ) );
  NAND3_X1 U6854 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i0[10] ), .A3(
        \SB2_0_25/i0[9] ), .ZN(\SB2_0_25/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U6855 ( .A1(n3166), .A2(\RI5[4][19] ), .Z(
        \MC_ARK_ARC_1_4/temp3[109] ) );
  NAND3_X2 U6856 ( .A1(\SB1_3_6/i0[10] ), .A2(\SB1_3_6/i0[6] ), .A3(
        \SB1_3_6/i0_0 ), .ZN(\SB1_3_6/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U6857 ( .A1(\MC_ARK_ARC_1_1/temp4[164] ), .A2(
        \MC_ARK_ARC_1_1/temp3[164] ), .Z(\MC_ARK_ARC_1_1/temp6[164] ) );
  NAND3_X2 U6864 ( .A1(\SB1_0_25/i0[10] ), .A2(\SB1_0_25/i0_3 ), .A3(
        \SB1_0_25/i0[6] ), .ZN(n2323) );
  XOR2_X1 U6867 ( .A1(\MC_ARK_ARC_1_2/temp6[140] ), .A2(
        \MC_ARK_ARC_1_2/temp5[140] ), .Z(\MC_ARK_ARC_1_2/buf_output[140] ) );
  NAND4_X2 U6871 ( .A1(\SB2_2_24/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_24/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_24/buf_output[1] ) );
  NAND4_X2 U6872 ( .A1(\SB1_2_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_28/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_28/Component_Function_1/NAND4_in[0] ), .A4(n2135), .ZN(
        \SB1_2_28/buf_output[1] ) );
  XOR2_X1 U6875 ( .A1(\RI5[2][67] ), .A2(\RI5[2][91] ), .Z(n2136) );
  NAND4_X2 U6876 ( .A1(\SB2_2_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_6/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_2_6/Component_Function_3/NAND4_in[1] ), .A4(n2983), .ZN(
        \SB2_2_6/buf_output[3] ) );
  XOR2_X1 U6877 ( .A1(\MC_ARK_ARC_1_4/temp5[167] ), .A2(
        \MC_ARK_ARC_1_4/temp6[167] ), .Z(\RI1[5][167] ) );
  NAND3_X1 U6880 ( .A1(\SB1_3_24/i0_0 ), .A2(\SB1_3_24/i3[0] ), .A3(
        \SB1_3_24/i1_7 ), .ZN(\SB1_3_24/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 U6884 ( .I(\SB2_0_20/buf_output[1] ), .Z(\RI5[0][91] ) );
  NAND2_X1 U6886 ( .A1(\SB1_2_15/i1[9] ), .A2(\RI1[2][101] ), .ZN(n2140) );
  BUF_X4 U6887 ( .I(\SB2_2_0/buf_output[1] ), .Z(\RI5[2][19] ) );
  XOR2_X1 U6892 ( .A1(n2142), .A2(\MC_ARK_ARC_1_4/temp5[27] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[27] ) );
  BUF_X4 U6896 ( .I(\SB2_1_5/buf_output[1] ), .Z(\RI5[1][181] ) );
  XOR2_X1 U6898 ( .A1(\MC_ARK_ARC_1_4/temp2[104] ), .A2(n2145), .Z(
        \MC_ARK_ARC_1_4/temp5[104] ) );
  XOR2_X1 U6899 ( .A1(\RI5[4][98] ), .A2(\RI5[4][104] ), .Z(n2145) );
  XOR2_X1 U6900 ( .A1(\RI5[3][50] ), .A2(\RI5[3][26] ), .Z(n2147) );
  XOR2_X1 U6901 ( .A1(\RI5[3][45] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[21] ), 
        .Z(n2629) );
  NAND3_X1 U6902 ( .A1(\SB2_4_8/i0_3 ), .A2(\SB2_4_8/i1[9] ), .A3(
        \SB2_4_8/i0[6] ), .ZN(\SB2_4_8/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U6904 ( .A1(n2149), .A2(\MC_ARK_ARC_1_4/temp5[184] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[184] ) );
  XOR2_X1 U6905 ( .A1(\MC_ARK_ARC_1_4/temp4[184] ), .A2(
        \MC_ARK_ARC_1_4/temp3[184] ), .Z(n2149) );
  BUF_X4 U6906 ( .I(\SB2_3_18/buf_output[3] ), .Z(\RI5[3][93] ) );
  BUF_X4 U6907 ( .I(\SB2_4_31/buf_output[2] ), .Z(\RI5[4][20] ) );
  XOR2_X1 U6908 ( .A1(\MC_ARK_ARC_1_3/temp3[93] ), .A2(
        \MC_ARK_ARC_1_3/temp4[93] ), .Z(\MC_ARK_ARC_1_3/temp6[93] ) );
  NAND3_X1 U6910 ( .A1(\SB1_0_24/i0[6] ), .A2(\SB1_0_24/i0_3 ), .A3(
        \SB1_0_24/i0[10] ), .ZN(\SB1_0_24/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U6912 ( .A1(\MC_ARK_ARC_1_3/temp5[151] ), .A2(
        \MC_ARK_ARC_1_3/temp6[151] ), .Z(\MC_ARK_ARC_1_3/buf_output[151] ) );
  XOR2_X1 U6913 ( .A1(n2153), .A2(n2503), .Z(\MC_ARK_ARC_1_4/buf_output[139] )
         );
  INV_X1 U6921 ( .I(\SB1_1_8/buf_output[0] ), .ZN(\SB2_1_3/i3[0] ) );
  NAND4_X2 U6923 ( .A1(\SB2_2_13/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_13/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_13/buf_output[1] ) );
  XOR2_X1 U6931 ( .A1(n2160), .A2(\MC_ARK_ARC_1_1/temp5[156] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[156] ) );
  XOR2_X1 U6932 ( .A1(\MC_ARK_ARC_1_1/temp3[156] ), .A2(
        \MC_ARK_ARC_1_1/temp4[156] ), .Z(n2160) );
  XOR2_X1 U6934 ( .A1(\RI5[4][59] ), .A2(n540), .Z(n2161) );
  NAND4_X2 U6940 ( .A1(\SB2_2_20/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_20/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_2_20/Component_Function_0/NAND4_in[0] ), .A4(n2165), .ZN(
        \SB2_2_20/buf_output[0] ) );
  NAND4_X2 U6943 ( .A1(\SB1_2_15/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_15/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_15/Component_Function_0/NAND4_in[1] ), .A4(n2167), .ZN(
        \SB1_2_15/buf_output[0] ) );
  XOR2_X1 U6947 ( .A1(\MC_ARK_ARC_1_2/temp4[60] ), .A2(
        \MC_ARK_ARC_1_2/temp3[60] ), .Z(n2168) );
  NAND2_X1 U6951 ( .A1(\SB1_0_0/i1[9] ), .A2(\SB1_0_0/i0_3 ), .ZN(n2170) );
  XOR2_X1 U6960 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[187] ), .A2(\RI5[1][19] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[49] ) );
  NAND4_X2 U6961 ( .A1(\SB2_2_23/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_23/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_2_23/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_23/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_23/buf_output[0] ) );
  NAND3_X2 U6962 ( .A1(\SB2_2_0/i0[7] ), .A2(\SB2_2_0/i0[6] ), .A3(
        \SB2_2_0/i0[8] ), .ZN(n2565) );
  XOR2_X1 U6963 ( .A1(n2804), .A2(n2177), .Z(\MC_ARK_ARC_1_0/buf_output[159] )
         );
  XOR2_X1 U6964 ( .A1(\MC_ARK_ARC_1_0/temp3[159] ), .A2(
        \MC_ARK_ARC_1_0/temp4[159] ), .Z(n2177) );
  XOR2_X1 U6967 ( .A1(n2179), .A2(n2178), .Z(\MC_ARK_ARC_1_1/buf_output[42] )
         );
  XOR2_X1 U6968 ( .A1(\MC_ARK_ARC_1_1/temp1[42] ), .A2(
        \MC_ARK_ARC_1_1/temp4[42] ), .Z(n2178) );
  XOR2_X1 U6969 ( .A1(n2687), .A2(\MC_ARK_ARC_1_1/temp3[42] ), .Z(n2179) );
  NAND3_X2 U6971 ( .A1(\SB2_1_27/i1[9] ), .A2(\SB2_1_27/i0[10] ), .A3(
        \SB2_1_27/i1_7 ), .ZN(\SB2_1_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U6975 ( .A1(\SB4_1/i0_3 ), .A2(\SB4_1/i0[10] ), .A3(\SB4_1/i0_4 ), 
        .ZN(\SB4_1/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U6980 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[76] ), .A2(\RI5[1][82] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[82] ) );
  NAND3_X1 U6981 ( .A1(\SB3_14/i0_3 ), .A2(\SB3_14/i0[8] ), .A3(\SB3_14/i1_7 ), 
        .ZN(\SB3_14/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U6982 ( .A1(\MC_ARK_ARC_1_4/temp3[149] ), .A2(
        \MC_ARK_ARC_1_4/temp4[149] ), .Z(n2186) );
  XOR2_X1 U6986 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[141] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[177] ), .Z(n2188) );
  XOR2_X1 U6988 ( .A1(\MC_ARK_ARC_1_0/temp3[156] ), .A2(
        \MC_ARK_ARC_1_0/temp4[156] ), .Z(n2189) );
  XOR2_X1 U6989 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[24] ), .A2(\RI5[2][48] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[78] ) );
  XOR2_X1 U6990 ( .A1(\MC_ARK_ARC_1_2/temp5[157] ), .A2(n2190), .Z(
        \MC_ARK_ARC_1_2/buf_output[157] ) );
  XOR2_X1 U6991 ( .A1(\MC_ARK_ARC_1_2/temp3[157] ), .A2(
        \MC_ARK_ARC_1_2/temp4[157] ), .Z(n2190) );
  XOR2_X1 U6994 ( .A1(\MC_ARK_ARC_1_3/temp3[80] ), .A2(
        \MC_ARK_ARC_1_3/temp4[80] ), .Z(n2192) );
  NAND4_X2 U6999 ( .A1(\SB1_1_15/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_1_15/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_1_15/Component_Function_0/NAND4_in[1] ), .A4(n2196), .ZN(
        \SB1_1_15/buf_output[0] ) );
  XOR2_X1 U7002 ( .A1(\MC_ARK_ARC_1_2/temp1[47] ), .A2(
        \MC_ARK_ARC_1_2/temp2[47] ), .Z(\MC_ARK_ARC_1_2/temp5[47] ) );
  XOR2_X1 U7003 ( .A1(\MC_ARK_ARC_1_0/temp5[40] ), .A2(
        \MC_ARK_ARC_1_0/temp6[40] ), .Z(\MC_ARK_ARC_1_0/buf_output[40] ) );
  INV_X2 U7004 ( .I(\SB1_2_10/buf_output[2] ), .ZN(\SB2_2_7/i1[9] ) );
  XOR2_X1 U7005 ( .A1(\RI5[3][113] ), .A2(\RI5[3][119] ), .Z(
        \MC_ARK_ARC_1_3/temp1[119] ) );
  NAND3_X1 U7006 ( .A1(\SB2_3_12/i0[9] ), .A2(\SB2_3_12/i1_5 ), .A3(
        \SB2_3_12/i0[6] ), .ZN(\SB2_3_12/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U7016 ( .A1(\RI5[2][105] ), .A2(\RI5[2][111] ), .Z(
        \MC_ARK_ARC_1_2/temp1[111] ) );
  XOR2_X1 U7018 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[109] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[133] ), .Z(n2204) );
  XOR2_X1 U7024 ( .A1(n2209), .A2(\MC_ARK_ARC_1_3/temp4[50] ), .Z(
        \MC_ARK_ARC_1_3/temp6[50] ) );
  NAND3_X2 U7027 ( .A1(\SB2_0_18/i0[9] ), .A2(\SB2_0_18/i0_3 ), .A3(
        \SB2_0_18/i0[8] ), .ZN(n2740) );
  NAND3_X1 U7028 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i0[10] ), .A3(
        \SB2_1_4/i0_4 ), .ZN(\SB2_1_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U7029 ( .A1(\SB2_3_3/i0[10] ), .A2(\SB2_3_3/i0_3 ), .A3(
        \SB2_3_3/i0[6] ), .ZN(\SB2_3_3/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U7030 ( .A1(n2211), .A2(n2212), .Z(\MC_ARK_ARC_1_1/temp5[0] ) );
  XOR2_X1 U7032 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[0] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[162] ), .Z(n2212) );
  NAND3_X1 U7036 ( .A1(\SB4_25/i0_4 ), .A2(n6266), .A3(\SB4_25/i0[6] ), .ZN(
        n2213) );
  BUF_X4 U7043 ( .I(\SB2_3_9/buf_output[2] ), .Z(\RI5[3][152] ) );
  NAND3_X1 U7044 ( .A1(\SB4_10/i0_4 ), .A2(\SB4_10/i1_7 ), .A3(\SB4_10/i0[8] ), 
        .ZN(\SB4_10/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U7045 ( .A1(\SB2_4_6/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_4_6/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_4_6/Component_Function_4/NAND4_in[0] ), .A4(n2216), .ZN(
        \SB2_4_6/buf_output[4] ) );
  NAND3_X1 U7048 ( .A1(\SB3_28/i0_4 ), .A2(\SB3_28/i1[9] ), .A3(\SB3_28/i1_5 ), 
        .ZN(\SB3_28/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U7054 ( .A1(n2221), .A2(\MC_ARK_ARC_1_1/temp1[74] ), .Z(
        \MC_ARK_ARC_1_1/temp5[74] ) );
  XOR2_X1 U7055 ( .A1(n2222), .A2(n2223), .Z(\MC_ARK_ARC_1_1/buf_output[69] )
         );
  XOR2_X1 U7057 ( .A1(\MC_ARK_ARC_1_1/temp1[69] ), .A2(
        \MC_ARK_ARC_1_1/temp4[69] ), .Z(n2223) );
  NAND3_X2 U7058 ( .A1(\SB2_4_3/i0[10] ), .A2(n3988), .A3(\SB2_4_3/i1[9] ), 
        .ZN(\SB2_4_3/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U7063 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[63] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[87] ), .Z(n2225) );
  NAND4_X2 U7064 ( .A1(\SB2_2_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_5/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_2_5/Component_Function_3/NAND4_in[1] ), .A4(n2226), .ZN(
        \SB2_2_5/buf_output[3] ) );
  XOR2_X1 U7066 ( .A1(\MC_ARK_ARC_1_1/temp5[100] ), .A2(
        \MC_ARK_ARC_1_1/temp6[100] ), .Z(\MC_ARK_ARC_1_1/buf_output[100] ) );
  INV_X4 U7067 ( .I(n3000), .ZN(\SB2_1_20/i0_4 ) );
  NAND3_X1 U7068 ( .A1(\SB1_4_8/i0[8] ), .A2(\SB1_4_8/i0_4 ), .A3(
        \SB1_4_8/i1_7 ), .ZN(\SB1_4_8/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U7073 ( .A1(\SB1_1_22/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_22/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_1_22/Component_Function_0/NAND4_in[1] ), .A4(n2229), .ZN(
        \SB1_1_22/buf_output[0] ) );
  XOR2_X1 U7075 ( .A1(\MC_ARK_ARC_1_0/temp2[132] ), .A2(n2230), .Z(n2767) );
  XOR2_X1 U7076 ( .A1(\RI5[0][126] ), .A2(\RI5[0][132] ), .Z(n2230) );
  NAND3_X2 U7079 ( .A1(\SB2_1_8/i0[7] ), .A2(\SB2_1_8/i0[8] ), .A3(
        \SB2_1_8/i0[6] ), .ZN(n2382) );
  NAND3_X1 U7083 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i0[8] ), .A3(\SB4_31/i0[9] ), .ZN(n2233) );
  XOR2_X1 U7086 ( .A1(\MC_ARK_ARC_1_4/temp5[175] ), .A2(
        \MC_ARK_ARC_1_4/temp6[175] ), .Z(\MC_ARK_ARC_1_4/buf_output[175] ) );
  XOR2_X1 U7088 ( .A1(\RI5[4][49] ), .A2(\RI5[4][13] ), .Z(
        \MC_ARK_ARC_1_4/temp3[139] ) );
  XOR2_X1 U7089 ( .A1(n2234), .A2(\MC_ARK_ARC_1_3/temp1[151] ), .Z(
        \MC_ARK_ARC_1_3/temp5[151] ) );
  XOR2_X1 U7090 ( .A1(\RI5[3][97] ), .A2(\RI5[3][121] ), .Z(n2234) );
  XOR2_X1 U7091 ( .A1(\MC_ARK_ARC_1_2/temp5[67] ), .A2(n2235), .Z(
        \MC_ARK_ARC_1_2/buf_output[67] ) );
  XOR2_X1 U7092 ( .A1(n2365), .A2(\MC_ARK_ARC_1_2/temp4[67] ), .Z(n2235) );
  NAND3_X1 U7099 ( .A1(\SB1_3_20/i0[6] ), .A2(\SB1_3_20/i1[9] ), .A3(
        \SB1_3_20/i0_3 ), .ZN(\SB1_3_20/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U7101 ( .I(\SB1_4_5/buf_output[2] ), .ZN(\SB2_4_2/i1[9] ) );
  NAND3_X1 U7103 ( .A1(\SB2_1_2/i0[10] ), .A2(\SB2_1_2/i0[6] ), .A3(
        \SB2_1_2/i0_0 ), .ZN(n2240) );
  XOR2_X1 U7105 ( .A1(n2241), .A2(\MC_ARK_ARC_1_3/temp2[152] ), .Z(
        \MC_ARK_ARC_1_3/temp5[152] ) );
  XOR2_X1 U7106 ( .A1(\MC_ARK_ARC_1_1/temp3[149] ), .A2(
        \MC_ARK_ARC_1_1/temp4[149] ), .Z(n2242) );
  XOR2_X1 U7109 ( .A1(n2245), .A2(\MC_ARK_ARC_1_2/temp4[8] ), .Z(n3055) );
  XOR2_X1 U7110 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[110] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[74] ), .Z(n2245) );
  XOR2_X1 U7111 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[135] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[171] ), .Z(\MC_ARK_ARC_1_4/temp3[69] )
         );
  XOR2_X1 U7114 ( .A1(\MC_ARK_ARC_1_1/temp4[53] ), .A2(
        \MC_ARK_ARC_1_1/temp3[53] ), .Z(\MC_ARK_ARC_1_1/temp6[53] ) );
  INV_X1 U7115 ( .I(\SB1_1_21/buf_output[1] ), .ZN(\SB2_1_17/i1_7 ) );
  NAND3_X2 U7116 ( .A1(\SB2_2_8/i0[10] ), .A2(\SB2_2_8/i0_0 ), .A3(
        \SB2_2_8/i0[6] ), .ZN(\SB2_2_8/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U7117 ( .A1(\SB3_4/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_4/Component_Function_0/NAND4_in[3] ), .A3(
        \SB3_4/Component_Function_0/NAND4_in[1] ), .A4(
        \SB3_4/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_4/buf_output[0] )
         );
  XOR2_X1 U7118 ( .A1(n3060), .A2(n2248), .Z(n2280) );
  XOR2_X1 U7119 ( .A1(\MC_ARK_ARC_1_3/temp3[47] ), .A2(n3179), .Z(n2248) );
  BUF_X4 U7121 ( .I(\SB2_1_0/buf_output[2] ), .Z(\RI5[1][14] ) );
  NAND4_X2 U7123 ( .A1(\SB2_1_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_2/NAND4_in[2] ), .A3(n2619), .A4(n2251), 
        .ZN(\SB2_1_4/buf_output[2] ) );
  NAND3_X1 U7124 ( .A1(\SB1_3_27/i0[8] ), .A2(\SB1_3_27/i1_7 ), .A3(
        \SB1_3_27/i0_4 ), .ZN(\SB1_3_27/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U7126 ( .A1(n3152), .A2(\SB2_1_24/Component_Function_5/NAND4_in[1] ), .A3(\SB2_1_24/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_24/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_24/buf_output[5] ) );
  NAND4_X2 U7127 ( .A1(\SB3_7/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_7/Component_Function_1/NAND4_in[2] ), .A3(
        \SB3_7/Component_Function_1/NAND4_in[0] ), .A4(
        \SB3_7/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_7/buf_output[1] )
         );
  XOR2_X1 U7131 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[80] ), .A2(\RI5[3][74] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[80] ) );
  XOR2_X1 U7132 ( .A1(\MC_ARK_ARC_1_4/temp3[24] ), .A2(
        \MC_ARK_ARC_1_4/temp4[24] ), .Z(n2256) );
  BUF_X4 U7136 ( .I(\SB2_3_27/buf_output[2] ), .Z(\RI5[3][44] ) );
  NAND3_X1 U7137 ( .A1(\SB2_2_30/i0[8] ), .A2(\SB2_2_30/i1_7 ), .A3(
        \SB1_2_31/buf_output[4] ), .ZN(
        \SB2_2_30/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U7138 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[3] ), .A2(\RI5[2][159] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[93] ) );
  XOR2_X1 U7148 ( .A1(\RI5[1][173] ), .A2(\RI5[1][137] ), .Z(n2263) );
  NAND3_X1 U7149 ( .A1(\SB1_2_23/i0[6] ), .A2(\SB1_2_23/i1[9] ), .A3(
        \SB1_2_23/i0_3 ), .ZN(\SB1_2_23/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U7150 ( .I(\SB2_2_29/buf_output[0] ), .Z(\RI5[2][42] ) );
  XOR2_X1 U7152 ( .A1(\MC_ARK_ARC_1_1/temp3[49] ), .A2(
        \MC_ARK_ARC_1_1/temp4[49] ), .Z(n2265) );
  INV_X2 U7153 ( .I(\RI3[0][39] ), .ZN(\SB2_0_25/i0[8] ) );
  NAND4_X2 U7154 ( .A1(\SB1_0_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_27/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_0_27/Component_Function_3/NAND4_in[2] ), .ZN(\RI3[0][39] ) );
  XOR2_X1 U7155 ( .A1(\MC_ARK_ARC_1_0/temp1[105] ), .A2(
        \MC_ARK_ARC_1_0/temp2[105] ), .Z(\MC_ARK_ARC_1_0/temp5[105] ) );
  NAND3_X1 U7157 ( .A1(\SB3_2/i1_5 ), .A2(\SB3_2/i1[9] ), .A3(\SB3_2/i0_4 ), 
        .ZN(\SB3_2/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U7158 ( .A1(\SB1_4_6/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_4_6/Component_Function_0/NAND4_in[0] ), .A3(n2583), .A4(n2268), 
        .ZN(\SB1_4_6/buf_output[0] ) );
  NAND4_X2 U7164 ( .A1(\SB4_2/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_2/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_2/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_2/Component_Function_1/NAND4_in[0] ), .ZN(n2457) );
  NAND4_X2 U7165 ( .A1(\SB1_3_5/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_0/NAND4_in[0] ), .A4(n2273), .ZN(
        \SB1_3_5/buf_output[0] ) );
  XOR2_X1 U7174 ( .A1(\MC_ARK_ARC_1_0/temp5[150] ), .A2(
        \MC_ARK_ARC_1_0/temp6[150] ), .Z(\MC_ARK_ARC_1_0/buf_output[150] ) );
  XOR2_X1 U7179 ( .A1(\MC_ARK_ARC_1_4/temp3[103] ), .A2(
        \MC_ARK_ARC_1_4/temp4[103] ), .Z(n2278) );
  XOR2_X1 U7180 ( .A1(\MC_ARK_ARC_1_4/temp5[106] ), .A2(n2279), .Z(
        \MC_ARK_ARC_1_4/buf_output[106] ) );
  XOR2_X1 U7181 ( .A1(\MC_ARK_ARC_1_4/temp3[106] ), .A2(
        \MC_ARK_ARC_1_4/temp4[106] ), .Z(n2279) );
  NAND3_X1 U7182 ( .A1(\SB2_4_9/i0_3 ), .A2(\SB2_4_9/i0[10] ), .A3(
        \SB2_4_9/i0_4 ), .ZN(\SB2_4_9/Component_Function_0/NAND4_in[2] ) );
  INV_X2 U7185 ( .I(n2280), .ZN(\MC_ARK_ARC_1_3/buf_output[47] ) );
  BUF_X4 U7189 ( .I(\SB2_3_15/buf_output[0] ), .Z(\RI5[3][126] ) );
  XOR2_X1 U7190 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[79] ), .A2(\RI5[2][85] ), 
        .Z(n2281) );
  NAND4_X2 U7193 ( .A1(\SB1_0_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_21/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_21/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_0_21/Component_Function_0/NAND4_in[1] ), .ZN(\RI3[0][90] ) );
  XOR2_X1 U7195 ( .A1(\RI5[4][32] ), .A2(\RI5[4][68] ), .Z(
        \MC_ARK_ARC_1_4/temp3[158] ) );
  XOR2_X1 U7196 ( .A1(n2284), .A2(\MC_ARK_ARC_1_3/temp6[89] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[89] ) );
  XOR2_X1 U7197 ( .A1(\RI5[4][152] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[188] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[86] ) );
  NAND3_X2 U7199 ( .A1(\SB2_4_18/i0_3 ), .A2(\SB2_4_18/i0_4 ), .A3(
        \SB2_4_18/i1[9] ), .ZN(n2285) );
  BUF_X4 U7201 ( .I(\SB2_2_1/buf_output[5] ), .Z(\RI5[2][185] ) );
  NAND4_X2 U7205 ( .A1(\SB2_0_29/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_0_29/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_29/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_0_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_29/buf_output[5] ) );
  NAND3_X1 U7208 ( .A1(n5429), .A2(\SB2_1_31/i1[9] ), .A3(\SB2_1_31/i1_5 ), 
        .ZN(\SB2_1_31/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U7213 ( .A1(\SB1_4_25/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_4_25/Component_Function_5/NAND4_in[3] ), .A3(n3117), .A4(
        \SB1_4_25/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_4_25/buf_output[5] ) );
  XOR2_X1 U7216 ( .A1(\MC_ARK_ARC_1_3/temp1[55] ), .A2(
        \MC_ARK_ARC_1_3/temp2[55] ), .Z(n2292) );
  NAND3_X1 U7217 ( .A1(\SB2_1_26/i0[8] ), .A2(\SB1_1_26/buf_output[5] ), .A3(
        \SB2_1_26/i0[9] ), .ZN(\SB2_1_26/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U7218 ( .A1(\MC_ARK_ARC_1_2/temp5[83] ), .A2(
        \MC_ARK_ARC_1_2/temp6[83] ), .Z(\MC_ARK_ARC_1_2/buf_output[83] ) );
  NOR2_X2 U7224 ( .A1(n2319), .A2(n2321), .ZN(\SB2_0_28/i0[7] ) );
  XOR2_X1 U7225 ( .A1(\MC_ARK_ARC_1_4/temp5[180] ), .A2(n2295), .Z(
        \MC_ARK_ARC_1_4/buf_output[180] ) );
  XOR2_X1 U7226 ( .A1(\MC_ARK_ARC_1_4/temp3[180] ), .A2(
        \MC_ARK_ARC_1_4/temp4[180] ), .Z(n2295) );
  NAND4_X2 U7231 ( .A1(\SB1_2_11/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_11/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_11/Component_Function_0/NAND4_in[1] ), .A4(n2297), .ZN(
        \SB1_2_11/buf_output[0] ) );
  XOR2_X1 U7234 ( .A1(n2300), .A2(n2299), .Z(n2987) );
  XOR2_X1 U7235 ( .A1(\RI5[0][132] ), .A2(n91), .Z(n2299) );
  XOR2_X1 U7236 ( .A1(\RI5[0][66] ), .A2(\RI5[0][96] ), .Z(n2300) );
  XOR2_X1 U7239 ( .A1(\RI5[2][13] ), .A2(n211), .Z(n2304) );
  XOR2_X1 U7243 ( .A1(\RI5[3][60] ), .A2(\RI5[3][66] ), .Z(
        \MC_ARK_ARC_1_3/temp1[66] ) );
  BUF_X4 U7244 ( .I(\SB2_4_16/buf_output[1] ), .Z(\RI5[4][115] ) );
  BUF_X4 U7250 ( .I(\SB2_4_11/buf_output[1] ), .Z(\RI5[4][145] ) );
  XOR2_X1 U7251 ( .A1(\MC_ARK_ARC_1_2/temp3[131] ), .A2(
        \MC_ARK_ARC_1_2/temp4[131] ), .Z(\MC_ARK_ARC_1_2/temp6[131] ) );
  XOR2_X1 U7253 ( .A1(\MC_ARK_ARC_1_4/temp2[119] ), .A2(n2313), .Z(
        \MC_ARK_ARC_1_4/temp5[119] ) );
  XOR2_X1 U7254 ( .A1(\RI5[4][113] ), .A2(\RI5[4][119] ), .Z(n2313) );
  NAND3_X2 U7256 ( .A1(\SB2_1_31/i0[10] ), .A2(\SB2_1_31/i1[9] ), .A3(
        \SB2_1_31/i1_7 ), .ZN(\SB2_1_31/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U7260 ( .A1(n2315), .A2(n68), .Z(Ciphertext[1]) );
  NAND4_X2 U7261 ( .A1(\SB4_31/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_31/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_31/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_31/Component_Function_1/NAND4_in[0] ), .ZN(n2315) );
  NAND3_X1 U7272 ( .A1(\SB2_4_18/i0_4 ), .A2(\SB2_4_18/i1_7 ), .A3(
        \SB2_4_18/i0[8] ), .ZN(n2316) );
  NAND3_X1 U7275 ( .A1(\SB2_2_1/i0[8] ), .A2(\SB2_2_1/i1_7 ), .A3(
        \SB1_2_2/buf_output[4] ), .ZN(
        \SB2_2_1/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U7278 ( .A1(\SB1_3_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_12/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_3_12/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_3_12/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_12/buf_output[0] ) );
  NAND3_X2 U7279 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i0_4 ), .A3(
        \SB2_1_14/i1[9] ), .ZN(\SB2_1_14/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7285 ( .A1(\MC_ARK_ARC_1_0/temp6[95] ), .A2(n2318), .Z(
        \MC_ARK_ARC_1_0/buf_output[95] ) );
  XOR2_X1 U7287 ( .A1(\RI5[1][68] ), .A2(\SB2_1_22/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/temp1[74] ) );
  XOR2_X1 U7292 ( .A1(\RI5[4][26] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[2] ), 
        .Z(n2324) );
  XOR2_X1 U7295 ( .A1(\MC_ARK_ARC_1_0/temp3[33] ), .A2(
        \MC_ARK_ARC_1_0/temp4[33] ), .Z(\MC_ARK_ARC_1_0/temp6[33] ) );
  XOR2_X1 U7297 ( .A1(\RI5[0][114] ), .A2(\RI5[0][138] ), .Z(
        \MC_ARK_ARC_1_0/temp2[168] ) );
  NAND3_X1 U7298 ( .A1(\SB2_0_17/i0_0 ), .A2(\SB2_0_17/i0_3 ), .A3(
        \SB2_0_17/i0[7] ), .ZN(\SB2_0_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U7301 ( .A1(\SB2_0_24/i0[6] ), .A2(\SB2_0_24/i0[8] ), .A3(
        \SB2_0_24/i0[7] ), .ZN(\SB2_0_24/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U7305 ( .A1(\MC_ARK_ARC_1_2/temp1[40] ), .A2(
        \MC_ARK_ARC_1_2/temp2[40] ), .Z(n2330) );
  XOR2_X1 U7309 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[73] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[97] ), .Z(n2332) );
  NAND4_X2 U7310 ( .A1(n2333), .A2(\SB2_0_18/Component_Function_3/NAND4_in[1] ), .A3(\SB2_0_18/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_0_18/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB2_0_18/buf_output[3] ) );
  XOR2_X1 U7313 ( .A1(\RI5[0][89] ), .A2(\RI5[0][53] ), .Z(n2334) );
  NAND3_X1 U7314 ( .A1(\SB1_4_13/i0_3 ), .A2(\SB1_4_13/i0[6] ), .A3(
        \SB1_4_13/i1[9] ), .ZN(\SB1_4_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U7319 ( .A1(n6277), .A2(\SB2_4_1/i0_4 ), .A3(\SB2_4_1/i0_0 ), .ZN(
        \SB2_4_1/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U7328 ( .A1(\MC_ARK_ARC_1_3/temp3[42] ), .A2(
        \MC_ARK_ARC_1_3/temp4[42] ), .Z(n2340) );
  BUF_X4 U7330 ( .I(\SB2_1_31/buf_output[5] ), .Z(\RI5[1][5] ) );
  NAND3_X1 U7337 ( .A1(\SB2_0_15/i0[10] ), .A2(n1508), .A3(\SB2_0_15/i1_7 ), 
        .ZN(\SB2_0_15/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U7338 ( .A1(n2344), .A2(\MC_ARK_ARC_1_4/temp5[0] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[0] ) );
  XOR2_X1 U7339 ( .A1(n2602), .A2(\MC_ARK_ARC_1_4/temp4[0] ), .Z(n2344) );
  NAND4_X2 U7346 ( .A1(\SB1_4_9/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_9/Component_Function_0/NAND4_in[0] ), .A4(n2348), .ZN(
        \SB1_4_9/buf_output[0] ) );
  XOR2_X1 U7347 ( .A1(\MC_ARK_ARC_1_3/temp2[178] ), .A2(
        \MC_ARK_ARC_1_3/temp1[178] ), .Z(\MC_ARK_ARC_1_3/temp5[178] ) );
  BUF_X4 U7349 ( .I(\SB2_3_12/buf_output[4] ), .Z(\RI5[3][124] ) );
  XOR2_X1 U7350 ( .A1(\MC_ARK_ARC_1_1/temp2[105] ), .A2(
        \MC_ARK_ARC_1_1/temp1[105] ), .Z(\MC_ARK_ARC_1_1/temp5[105] ) );
  NAND4_X2 U7351 ( .A1(\SB1_4_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_4_5/Component_Function_3/NAND4_in[3] ), .A4(n2350), .ZN(
        \SB1_4_5/buf_output[3] ) );
  NAND3_X1 U7352 ( .A1(\SB1_4_17/i0_0 ), .A2(\SB1_4_17/i1_7 ), .A3(
        \SB1_4_17/i3[0] ), .ZN(\SB1_4_17/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U7354 ( .A1(\MC_ARK_ARC_1_4/temp1[45] ), .A2(n2351), .Z(n2582) );
  XOR2_X1 U7355 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[183] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[15] ), .Z(n2351) );
  BUF_X4 U7356 ( .I(\SB2_3_30/buf_output[1] ), .Z(\RI5[3][31] ) );
  XOR2_X1 U7361 ( .A1(\RI5[0][115] ), .A2(\RI5[0][151] ), .Z(
        \MC_ARK_ARC_1_0/temp3[49] ) );
  NAND3_X2 U7363 ( .A1(\SB2_1_21/i0_3 ), .A2(\SB2_1_21/i0_0 ), .A3(
        \SB2_1_21/i0_4 ), .ZN(\SB2_1_21/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 U7370 ( .I(\SB2_4_24/buf_output[4] ), .Z(\RI5[4][52] ) );
  XOR2_X1 U7373 ( .A1(\RI5[3][17] ), .A2(\RI5[3][185] ), .Z(
        \MC_ARK_ARC_1_3/temp2[47] ) );
  XOR2_X1 U7375 ( .A1(n2360), .A2(n2359), .Z(\MC_ARK_ARC_1_2/buf_output[137] )
         );
  XOR2_X1 U7376 ( .A1(\MC_ARK_ARC_1_2/temp1[137] ), .A2(
        \MC_ARK_ARC_1_2/temp4[137] ), .Z(n2359) );
  XOR2_X1 U7377 ( .A1(\MC_ARK_ARC_1_1/temp1[75] ), .A2(
        \MC_ARK_ARC_1_1/temp2[75] ), .Z(n2361) );
  NAND4_X2 U7378 ( .A1(\SB2_1_31/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_1_31/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_31/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_1_31/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_1_31/buf_output[2] ) );
  NAND3_X1 U7380 ( .A1(\SB3_7/i0_3 ), .A2(\SB3_7/i0[8] ), .A3(\SB3_7/i1_7 ), 
        .ZN(\SB3_7/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U7383 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[133] ), .A2(\RI5[2][169] ), 
        .Z(n2365) );
  BUF_X4 U7384 ( .I(\SB2_0_17/buf_output[1] ), .Z(\RI5[0][109] ) );
  INV_X2 U7388 ( .I(\SB1_3_19/buf_output[5] ), .ZN(\SB2_3_19/i1_5 ) );
  XOR2_X1 U7390 ( .A1(\RI5[2][119] ), .A2(\RI5[2][83] ), .Z(
        \MC_ARK_ARC_1_2/temp3[17] ) );
  XOR2_X1 U7391 ( .A1(\MC_ARK_ARC_1_3/temp6[175] ), .A2(n2366), .Z(
        \MC_ARK_ARC_1_3/buf_output[175] ) );
  XOR2_X1 U7392 ( .A1(\MC_ARK_ARC_1_3/temp2[175] ), .A2(
        \MC_ARK_ARC_1_3/temp1[175] ), .Z(n2366) );
  NAND3_X1 U7394 ( .A1(\SB2_2_18/i1[9] ), .A2(\SB2_2_18/i0_4 ), .A3(
        \SB2_2_18/i1_5 ), .ZN(\SB2_2_18/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U7395 ( .A1(\MC_ARK_ARC_1_2/temp6[94] ), .A2(n2367), .Z(
        \MC_ARK_ARC_1_2/buf_output[94] ) );
  XOR2_X1 U7409 ( .A1(\MC_ARK_ARC_1_2/temp3[24] ), .A2(
        \MC_ARK_ARC_1_2/temp4[24] ), .Z(n2377) );
  NAND3_X1 U7412 ( .A1(\SB2_0_3/i0[7] ), .A2(\SB2_0_3/i0[8] ), .A3(
        \SB2_0_3/i0[6] ), .ZN(\SB2_0_3/Component_Function_0/NAND4_in[1] ) );
  INV_X2 U7417 ( .I(n2381), .ZN(\SB2_0_5/i0_4 ) );
  XOR2_X1 U7420 ( .A1(\MC_ARK_ARC_1_2/temp6[37] ), .A2(
        \MC_ARK_ARC_1_2/temp5[37] ), .Z(\MC_ARK_ARC_1_2/buf_output[37] ) );
  NAND3_X1 U7421 ( .A1(\SB1_1_15/i0_0 ), .A2(\SB1_1_15/i0_3 ), .A3(
        \SB1_1_15/i0[7] ), .ZN(\SB1_1_15/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U7423 ( .A1(\SB2_1_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_6/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_6/Component_Function_2/NAND4_in[1] ), .A4(n2384), .ZN(
        \SB2_1_6/buf_output[2] ) );
  NAND3_X2 U7424 ( .A1(\SB2_1_6/i0_0 ), .A2(\SB2_1_6/i1_5 ), .A3(
        \SB2_1_6/i0_4 ), .ZN(n2384) );
  AND2_X1 U7427 ( .A1(\SB2_4_6/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_4_6/Component_Function_1/NAND4_in[1] ), .Z(n2387) );
  XOR2_X1 U7428 ( .A1(n2388), .A2(\MC_ARK_ARC_1_2/temp1[101] ), .Z(
        \MC_ARK_ARC_1_2/temp5[101] ) );
  BUF_X4 U7432 ( .I(\SB2_2_20/buf_output[1] ), .Z(\RI5[2][91] ) );
  NAND3_X1 U7437 ( .A1(\SB2_4_5/i0_0 ), .A2(\SB2_4_5/i3[0] ), .A3(
        \SB2_4_5/i1_7 ), .ZN(\SB2_4_5/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U7440 ( .A1(\MC_ARK_ARC_1_1/temp5[130] ), .A2(n2395), .Z(
        \MC_ARK_ARC_1_1/buf_output[130] ) );
  XOR2_X1 U7441 ( .A1(\MC_ARK_ARC_1_1/temp3[130] ), .A2(
        \MC_ARK_ARC_1_1/temp4[130] ), .Z(n2395) );
  NAND4_X2 U7443 ( .A1(\SB1_0_24/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_24/Component_Function_4/NAND4_in[0] ), .A4(n2396), .ZN(
        \SB1_0_24/buf_output[4] ) );
  NAND3_X1 U7448 ( .A1(\SB4_9/i0[6] ), .A2(n1499), .A3(\SB4_9/i0[7] ), .ZN(
        \SB4_9/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U7449 ( .A1(\SB1_4_12/i0[8] ), .A2(\SB1_4_12/i0_4 ), .A3(
        \SB1_4_12/i1_7 ), .ZN(\SB1_4_12/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U7466 ( .A1(\SB1_3_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_3/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_3_3/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_3_3/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_3/buf_output[3] ) );
  NAND3_X1 U7467 ( .A1(\SB4_3/i0_3 ), .A2(\SB4_3/i0_0 ), .A3(\SB4_3/i0_4 ), 
        .ZN(\SB4_3/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U7472 ( .A1(\SB2_1_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_3/NAND4_in[1] ), .A3(n3101), .A4(
        \SB2_1_18/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_18/buf_output[3] ) );
  XOR2_X1 U7474 ( .A1(\RI5[4][1] ), .A2(\RI5[4][37] ), .Z(
        \MC_ARK_ARC_1_4/temp3[127] ) );
  NAND3_X2 U7480 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i0_4 ), .A3(
        \SB1_0_12/i1[9] ), .ZN(n2414) );
  XOR2_X1 U7482 ( .A1(\MC_ARK_ARC_1_3/temp2[96] ), .A2(
        \MC_ARK_ARC_1_3/temp1[96] ), .Z(\MC_ARK_ARC_1_3/temp5[96] ) );
  NAND4_X2 U7483 ( .A1(\SB2_0_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_12/Component_Function_5/NAND4_in[0] ), .A3(
        \SB2_0_12/Component_Function_5/NAND4_in[1] ), .A4(n2418), .ZN(
        \SB2_0_12/buf_output[5] ) );
  NAND4_X2 U7490 ( .A1(\SB2_1_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_4/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_1_4/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_4/buf_output[1] ) );
  XOR2_X1 U7495 ( .A1(\MC_ARK_ARC_1_3/temp6[148] ), .A2(
        \MC_ARK_ARC_1_3/temp5[148] ), .Z(\MC_ARK_ARC_1_3/buf_output[148] ) );
  XOR2_X1 U7496 ( .A1(\MC_ARK_ARC_1_0/temp1[8] ), .A2(n2421), .Z(
        \MC_ARK_ARC_1_0/temp5[8] ) );
  XOR2_X1 U7497 ( .A1(\RI5[0][146] ), .A2(\RI5[0][170] ), .Z(n2421) );
  XOR2_X1 U7499 ( .A1(\MC_ARK_ARC_1_0/temp4[23] ), .A2(
        \MC_ARK_ARC_1_0/temp3[23] ), .Z(n2422) );
  XOR2_X1 U7501 ( .A1(\RI5[4][85] ), .A2(\RI5[4][109] ), .Z(n2423) );
  XOR2_X1 U7503 ( .A1(\RI5[1][128] ), .A2(\RI5[1][134] ), .Z(n2425) );
  INV_X2 U7504 ( .I(\SB1_2_18/buf_output[5] ), .ZN(\SB2_2_18/i1_5 ) );
  NAND4_X2 U7507 ( .A1(\SB2_1_2/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_2/Component_Function_4/NAND4_in[0] ), .A4(n2427), .ZN(
        \SB2_1_2/buf_output[4] ) );
  BUF_X4 U7511 ( .I(\SB2_2_16/buf_output[3] ), .Z(\RI5[2][105] ) );
  XOR2_X1 U7514 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[46] ), .A2(\RI5[3][70] ), 
        .Z(n2433) );
  XOR2_X1 U7517 ( .A1(\RI5[0][159] ), .A2(\RI5[0][183] ), .Z(n2434) );
  NAND3_X2 U7520 ( .A1(\SB1_3_20/i0[6] ), .A2(\SB1_3_20/i0_4 ), .A3(
        \SB1_3_20/i0[9] ), .ZN(n2533) );
  XOR2_X1 U7528 ( .A1(n2439), .A2(\MC_ARK_ARC_1_2/temp6[127] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[127] ) );
  XOR2_X1 U7529 ( .A1(\MC_ARK_ARC_1_2/temp1[127] ), .A2(
        \MC_ARK_ARC_1_2/temp2[127] ), .Z(n2439) );
  BUF_X4 U7531 ( .I(\SB2_2_28/buf_output[2] ), .Z(\RI5[2][38] ) );
  XOR2_X1 U7535 ( .A1(\MC_ARK_ARC_1_4/temp2[161] ), .A2(
        \MC_ARK_ARC_1_4/temp1[161] ), .Z(n2441) );
  BUF_X4 U7536 ( .I(\SB2_2_24/buf_output[0] ), .Z(\RI5[2][72] ) );
  NAND4_X2 U7544 ( .A1(\SB1_0_20/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_20/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_20/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_20/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][96] ) );
  XOR2_X1 U7546 ( .A1(\MC_ARK_ARC_1_0/temp3[31] ), .A2(
        \MC_ARK_ARC_1_0/temp4[31] ), .Z(n2446) );
  NAND3_X1 U7547 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i0[9] ), .A3(
        \SB1_1_2/i0[8] ), .ZN(\SB1_1_2/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U7548 ( .A1(\SB1_0_24/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_24/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_24/Component_Function_1/NAND4_in[0] ), .A4(n2447), .ZN(
        \RI3[0][67] ) );
  NAND3_X1 U7555 ( .A1(\SB1_1_20/i0_0 ), .A2(\SB1_1_20/i0_4 ), .A3(
        \SB1_1_20/i1_5 ), .ZN(n2450) );
  BUF_X4 U7556 ( .I(\SB2_1_17/buf_output[0] ), .Z(\RI5[1][114] ) );
  XOR2_X1 U7558 ( .A1(n2452), .A2(\MC_ARK_ARC_1_2/temp4[127] ), .Z(
        \MC_ARK_ARC_1_2/temp6[127] ) );
  XOR2_X1 U7559 ( .A1(\RI5[2][1] ), .A2(\RI5[2][37] ), .Z(n2452) );
  XOR2_X1 U7565 ( .A1(n2457), .A2(n5), .Z(Ciphertext[175]) );
  NOR2_X2 U7567 ( .A1(n2459), .A2(n2458), .ZN(\SB2_1_19/i0[7] ) );
  XOR2_X1 U7569 ( .A1(\MC_ARK_ARC_1_4/temp5[120] ), .A2(n2460), .Z(
        \MC_ARK_ARC_1_4/buf_output[120] ) );
  XOR2_X1 U7570 ( .A1(\MC_ARK_ARC_1_4/temp3[120] ), .A2(
        \MC_ARK_ARC_1_4/temp4[120] ), .Z(n2460) );
  NAND2_X1 U7571 ( .A1(\SB1_4_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_9/Component_Function_4/NAND4_in[2] ), .ZN(n2718) );
  NAND3_X1 U7575 ( .A1(\SB4_28/i0_0 ), .A2(\SB4_28/i0[10] ), .A3(
        \SB4_28/i0[6] ), .ZN(\SB4_28/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U7582 ( .A1(\RI5[3][41] ), .A2(\RI5[3][47] ), .Z(n2462) );
  XOR2_X1 U7584 ( .A1(\MC_ARK_ARC_1_3/temp1[61] ), .A2(
        \MC_ARK_ARC_1_3/temp2[61] ), .Z(\MC_ARK_ARC_1_3/temp5[61] ) );
  XOR2_X1 U7587 ( .A1(\MC_ARK_ARC_1_4/temp1[151] ), .A2(
        \MC_ARK_ARC_1_4/temp2[151] ), .Z(\MC_ARK_ARC_1_4/temp5[151] ) );
  NAND3_X1 U7588 ( .A1(\SB4_3/i0_3 ), .A2(\SB4_3/i0_4 ), .A3(\SB4_3/i1[9] ), 
        .ZN(\SB4_3/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7589 ( .A1(\RI5[3][179] ), .A2(\RI5[3][173] ), .Z(
        \MC_ARK_ARC_1_3/temp1[179] ) );
  BUF_X4 U7598 ( .I(\SB2_1_10/buf_output[0] ), .Z(\RI5[1][156] ) );
  XOR2_X1 U7602 ( .A1(\RI5[0][115] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[139] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[169] ) );
  XOR2_X1 U7606 ( .A1(\MC_ARK_ARC_1_1/temp5[166] ), .A2(n2474), .Z(
        \MC_ARK_ARC_1_1/buf_output[166] ) );
  XOR2_X1 U7607 ( .A1(\MC_ARK_ARC_1_1/temp4[166] ), .A2(
        \MC_ARK_ARC_1_1/temp3[166] ), .Z(n2474) );
  XOR2_X1 U7619 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[184] ), .A2(\RI5[3][16] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[46] ) );
  XOR2_X1 U7620 ( .A1(n2480), .A2(\MC_ARK_ARC_1_0/temp6[26] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[26] ) );
  XOR2_X1 U7624 ( .A1(\MC_ARK_ARC_1_4/temp5[150] ), .A2(
        \MC_ARK_ARC_1_4/temp6[150] ), .Z(\MC_ARK_ARC_1_4/buf_output[150] ) );
  XOR2_X1 U7625 ( .A1(\RI5[0][120] ), .A2(\RI5[0][156] ), .Z(
        \MC_ARK_ARC_1_0/temp3[54] ) );
  XOR2_X1 U7626 ( .A1(\RI5[3][167] ), .A2(\RI5[3][131] ), .Z(
        \MC_ARK_ARC_1_3/temp3[65] ) );
  NAND3_X1 U7627 ( .A1(\SB4_31/i0[6] ), .A2(\SB4_31/i0[8] ), .A3(
        \SB4_31/i0[7] ), .ZN(\SB4_31/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U7635 ( .A1(\RI5[0][6] ), .A2(\RI5[0][42] ), .Z(n2485) );
  XOR2_X1 U7640 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[34] ), .A2(\RI5[1][70] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[160] ) );
  NAND3_X1 U7641 ( .A1(\SB4_14/i0_4 ), .A2(\SB4_14/i0[9] ), .A3(\SB4_14/i0[6] ), .ZN(\SB4_14/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 U7642 ( .I(\SB2_4_3/buf_output[0] ), .Z(\RI5[4][6] ) );
  NAND3_X2 U7648 ( .A1(\SB2_4_3/i0_0 ), .A2(\SB2_4_3/i0[10] ), .A3(
        \SB2_4_3/i0[6] ), .ZN(\SB2_4_3/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U7649 ( .A1(\RI5[2][1] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .Z(n2495) );
  NAND4_X2 U7650 ( .A1(\SB1_3_19/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_1/NAND4_in[0] ), .A4(n2497), .ZN(
        \SB1_3_19/buf_output[1] ) );
  NAND3_X2 U7656 ( .A1(\SB2_1_31/i0_3 ), .A2(\SB2_1_31/i1[9] ), .A3(n5430), 
        .ZN(n2500) );
  XOR2_X1 U7659 ( .A1(\MC_ARK_ARC_1_4/temp3[139] ), .A2(
        \MC_ARK_ARC_1_4/temp4[139] ), .Z(n2503) );
  XOR2_X1 U7660 ( .A1(\MC_ARK_ARC_1_2/temp2[77] ), .A2(
        \MC_ARK_ARC_1_2/temp1[77] ), .Z(\MC_ARK_ARC_1_2/temp5[77] ) );
  XOR2_X1 U7661 ( .A1(\MC_ARK_ARC_1_0/temp2[133] ), .A2(
        \MC_ARK_ARC_1_0/temp1[133] ), .Z(\MC_ARK_ARC_1_0/temp5[133] ) );
  XOR2_X1 U7665 ( .A1(\RI5[0][136] ), .A2(\RI5[0][142] ), .Z(
        \MC_ARK_ARC_1_0/temp1[142] ) );
  XOR2_X1 U7669 ( .A1(\MC_ARK_ARC_1_1/temp2[152] ), .A2(
        \MC_ARK_ARC_1_1/temp1[152] ), .Z(\MC_ARK_ARC_1_1/temp5[152] ) );
  XOR2_X1 U7672 ( .A1(\MC_ARK_ARC_1_0/temp2[178] ), .A2(
        \MC_ARK_ARC_1_0/temp1[178] ), .Z(\MC_ARK_ARC_1_0/temp5[178] ) );
  NAND3_X1 U7673 ( .A1(\SB1_3_25/i0_0 ), .A2(\SB1_3_25/i1_7 ), .A3(
        \SB1_3_25/i3[0] ), .ZN(\SB1_3_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U7674 ( .A1(n7587), .A2(\SB2_4_5/i0[8] ), .A3(\SB2_4_5/i0[6] ), 
        .ZN(\SB2_4_5/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U7677 ( .A1(n2511), .A2(\MC_ARK_ARC_1_4/temp5[16] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[16] ) );
  XOR2_X1 U7678 ( .A1(\MC_ARK_ARC_1_4/temp4[16] ), .A2(
        \MC_ARK_ARC_1_4/temp3[16] ), .Z(n2511) );
  NAND3_X1 U7682 ( .A1(\SB3_15/buf_output[3] ), .A2(\SB4_13/i0_3 ), .A3(
        \SB4_13/i0[9] ), .ZN(\SB4_13/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U7691 ( .A1(n2518), .A2(\MC_ARK_ARC_1_0/temp6[113] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[113] ) );
  XOR2_X1 U7695 ( .A1(\MC_ARK_ARC_1_0/temp2[1] ), .A2(
        \MC_ARK_ARC_1_0/temp1[1] ), .Z(n2520) );
  XOR2_X1 U7702 ( .A1(\MC_ARK_ARC_1_4/temp4[13] ), .A2(
        \MC_ARK_ARC_1_4/temp3[13] ), .Z(n2525) );
  NAND4_X2 U7711 ( .A1(\SB2_3_20/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_20/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_3_20/Component_Function_0/NAND4_in[3] ), .A4(n2532), .ZN(
        \SB2_3_20/buf_output[0] ) );
  NAND3_X1 U7713 ( .A1(\SB3_0/i0_4 ), .A2(\SB3_0/i0[8] ), .A3(\SB3_0/i1_7 ), 
        .ZN(n2769) );
  NAND4_X2 U7716 ( .A1(\SB1_2_31/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_31/Component_Function_5/NAND4_in[3] ), .A3(n3091), .A4(
        \SB1_2_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_31/buf_output[5] ) );
  CLKBUF_X4 U7717 ( .I(\SB2_3_22/buf_output[0] ), .Z(\RI5[3][84] ) );
  XOR2_X1 U7719 ( .A1(\RI5[0][51] ), .A2(\RI5[0][45] ), .Z(n2534) );
  NAND4_X2 U7727 ( .A1(\SB2_2_13/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_13/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_13/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_2_13/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_2_13/buf_output[4] ) );
  NAND4_X2 U7731 ( .A1(\SB2_1_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_18/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_1_18/buf_output[1] ) );
  NAND3_X1 U7734 ( .A1(\SB2_3_25/i0_3 ), .A2(\SB2_3_25/i0[10] ), .A3(
        \SB2_3_25/i0_4 ), .ZN(\SB2_3_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U7735 ( .A1(\SB1_4_13/i0_3 ), .A2(\SB1_4_13/i0_0 ), .A3(
        \SB1_4_13/i0_4 ), .ZN(\SB1_4_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U7736 ( .A1(\SB2_4_12/i0[6] ), .A2(\SB2_4_12/i1_5 ), .A3(
        \SB2_4_12/i0[9] ), .ZN(\SB2_4_12/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U7740 ( .A1(\SB1_0_17/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_17/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_17/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_0_17/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][89] ) );
  BUF_X4 U7743 ( .I(\SB2_1_12/buf_output[3] ), .Z(\RI5[1][129] ) );
  XOR2_X1 U7753 ( .A1(\MC_ARK_ARC_1_4/temp6[187] ), .A2(
        \MC_ARK_ARC_1_4/temp5[187] ), .Z(\MC_ARK_ARC_1_4/buf_output[187] ) );
  NAND4_X2 U7754 ( .A1(\SB1_0_17/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_17/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][109] ) );
  XOR2_X1 U7755 ( .A1(\RI5[2][32] ), .A2(\RI5[2][38] ), .Z(
        \MC_ARK_ARC_1_2/temp1[38] ) );
  NAND3_X1 U7756 ( .A1(\SB1_1_18/i0[10] ), .A2(\SB1_1_18/i1[9] ), .A3(
        \SB1_1_18/i1_5 ), .ZN(\SB1_1_18/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U7760 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[122] ), .A2(\RI5[1][128] ), 
        .Z(n2552) );
  XOR2_X1 U7761 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[74] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[98] ), .Z(\MC_ARK_ARC_1_2/temp2[128] )
         );
  XOR2_X1 U7762 ( .A1(\MC_ARK_ARC_1_1/temp3[191] ), .A2(
        \MC_ARK_ARC_1_1/temp4[191] ), .Z(n2553) );
  NAND4_X2 U7763 ( .A1(\SB2_3_25/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_25/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_25/Component_Function_3/NAND4_in[3] ), .A4(n3106), .ZN(
        \SB2_3_25/buf_output[3] ) );
  XOR2_X1 U7765 ( .A1(\SB2_4_6/buf_output[3] ), .A2(\SB2_4_10/buf_output[3] ), 
        .Z(n3070) );
  BUF_X4 U7766 ( .I(\SB2_3_25/buf_output[3] ), .Z(\RI5[3][51] ) );
  XOR2_X1 U7774 ( .A1(\MC_ARK_ARC_1_3/temp4[2] ), .A2(n2563), .Z(
        \MC_ARK_ARC_1_3/temp6[2] ) );
  XOR2_X1 U7775 ( .A1(\RI5[3][68] ), .A2(\RI5[3][104] ), .Z(n2563) );
  INV_X2 U7777 ( .I(\SB1_1_15/buf_output[5] ), .ZN(\SB2_1_15/i1_5 ) );
  XOR2_X1 U7779 ( .A1(\MC_ARK_ARC_1_4/temp2[128] ), .A2(
        \MC_ARK_ARC_1_4/temp1[128] ), .Z(\MC_ARK_ARC_1_4/temp5[128] ) );
  XOR2_X1 U7780 ( .A1(\MC_ARK_ARC_1_2/temp5[176] ), .A2(
        \MC_ARK_ARC_1_2/temp6[176] ), .Z(\MC_ARK_ARC_1_2/buf_output[176] ) );
  INV_X2 U7782 ( .I(\SB1_3_12/buf_output[3] ), .ZN(\SB2_3_10/i0[8] ) );
  NAND4_X2 U7784 ( .A1(\SB2_2_0/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_0/Component_Function_0/NAND4_in[0] ), .A3(n2566), .A4(n2565), 
        .ZN(\SB2_2_0/buf_output[0] ) );
  NAND3_X1 U7790 ( .A1(\SB1_0_17/i0_0 ), .A2(\SB1_0_17/i1_5 ), .A3(
        \SB1_0_17/i0_4 ), .ZN(n2569) );
  INV_X2 U7796 ( .I(n2572), .ZN(\RI1[4][5] ) );
  XNOR2_X1 U7797 ( .A1(\MC_ARK_ARC_1_3/temp5[5] ), .A2(
        \MC_ARK_ARC_1_3/temp6[5] ), .ZN(n2572) );
  XOR2_X1 U7807 ( .A1(\RI5[2][108] ), .A2(\RI5[2][114] ), .Z(
        \MC_ARK_ARC_1_2/temp1[114] ) );
  NAND4_X2 U7810 ( .A1(\SB3_12/Component_Function_0/NAND4_in[1] ), .A2(
        \SB3_12/Component_Function_0/NAND4_in[0] ), .A3(n2581), .A4(n2580), 
        .ZN(\SB3_12/buf_output[0] ) );
  XOR2_X1 U7812 ( .A1(n2582), .A2(\MC_ARK_ARC_1_4/temp6[45] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[45] ) );
  BUF_X4 U7814 ( .I(\SB2_1_26/buf_output[0] ), .Z(\RI5[1][60] ) );
  NAND3_X2 U7818 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i1[9] ), .A3(\SB3_30/i0_4 ), 
        .ZN(n2585) );
  XOR2_X1 U7821 ( .A1(\MC_ARK_ARC_1_1/temp6[3] ), .A2(n2590), .Z(
        \MC_ARK_ARC_1_1/buf_output[3] ) );
  XOR2_X1 U7822 ( .A1(\MC_ARK_ARC_1_1/temp2[3] ), .A2(
        \MC_ARK_ARC_1_1/temp1[3] ), .Z(n2590) );
  NAND4_X2 U7823 ( .A1(\SB2_2_29/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_29/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_2_29/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_2_29/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_29/buf_output[0] ) );
  NAND4_X2 U7826 ( .A1(\SB1_4_16/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_4_16/Component_Function_4/NAND4_in[0] ), .A3(n2905), .A4(
        \SB1_4_16/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_4_16/buf_output[4] ) );
  BUF_X4 U7828 ( .I(\SB2_1_5/buf_output[2] ), .Z(\RI5[1][176] ) );
  BUF_X4 U7834 ( .I(\SB2_2_3/buf_output[1] ), .Z(\RI5[2][1] ) );
  NAND3_X1 U7835 ( .A1(\SB2_3_4/i0[6] ), .A2(\SB2_3_4/i0[8] ), .A3(n5683), 
        .ZN(\SB2_3_4/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U7838 ( .A1(\SB2_0_12/i1_5 ), .A2(\SB2_0_12/i3[0] ), .A3(
        \SB2_0_12/i0[8] ), .ZN(\SB2_0_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U7843 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i0[8] ), .A3(\SB3_2/i1_7 ), 
        .ZN(\SB3_2/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U7845 ( .A1(\RI5[4][66] ), .A2(\RI5[4][102] ), .Z(n2602) );
  XOR2_X1 U7846 ( .A1(\RI5[4][17] ), .A2(\RI5[4][11] ), .Z(
        \MC_ARK_ARC_1_4/temp1[17] ) );
  NAND3_X1 U7851 ( .A1(\SB4_31/i0[10] ), .A2(\SB4_31/i1_5 ), .A3(
        \SB4_31/i1[9] ), .ZN(\SB4_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U7852 ( .A1(\SB2_2_10/i0[10] ), .A2(\SB2_2_10/i0_0 ), .A3(
        \SB2_2_10/i0[6] ), .ZN(\SB2_2_10/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U7860 ( .A1(\RI5[1][191] ), .A2(\RI5[1][5] ), .Z(
        \MC_ARK_ARC_1_1/temp1[5] ) );
  XOR2_X1 U7862 ( .A1(\RI5[1][169] ), .A2(\RI5[1][13] ), .Z(
        \MC_ARK_ARC_1_1/temp3[103] ) );
  AND2_X1 U7863 ( .A1(\SB2_1_1/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_1/Component_Function_1/NAND4_in[2] ), .Z(n2613) );
  NAND2_X1 U7864 ( .A1(\SB3_15/i1[9] ), .A2(\SB3_15/i0_3 ), .ZN(
        \SB3_15/Component_Function_1/NAND4_in[0] ) );
  NAND4_X2 U7865 ( .A1(n2738), .A2(\SB1_0_6/Component_Function_1/NAND4_in[1] ), 
        .A3(\SB1_0_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_6/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][175] ) );
  NAND2_X1 U7867 ( .A1(\SB1_1_2/i1_5 ), .A2(n2614), .ZN(
        \SB1_1_2/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U7870 ( .A1(\SB1_2_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_3/NAND4_in[3] ), .A4(n2616), .ZN(
        \SB1_2_6/buf_output[3] ) );
  NAND3_X2 U7874 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i1[9] ), .A3(
        \SB2_1_22/i0_4 ), .ZN(\SB2_1_22/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7876 ( .A1(\MC_ARK_ARC_1_0/temp1[46] ), .A2(n2618), .Z(
        \MC_ARK_ARC_1_0/temp5[46] ) );
  NAND3_X1 U7885 ( .A1(\SB4_1/i0_3 ), .A2(\SB4_1/i1[9] ), .A3(
        \SB3_5/buf_output[1] ), .ZN(\SB4_1/Component_Function_3/NAND4_in[0] )
         );
  NOR2_X2 U7886 ( .A1(n2626), .A2(n2624), .ZN(n2965) );
  NAND3_X1 U7891 ( .A1(\SB2_2_0/i1[9] ), .A2(n5444), .A3(\SB2_2_0/i1_5 ), .ZN(
        \SB2_2_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U7894 ( .A1(\SB4_15/i0_4 ), .A2(\SB4_15/i1[9] ), .A3(\SB4_15/i1_5 ), 
        .ZN(\SB4_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U7895 ( .A1(\SB2_1_21/i0_3 ), .A2(\SB2_1_21/i0_4 ), .A3(
        \SB2_1_21/i1[9] ), .ZN(n2630) );
  NAND3_X1 U7896 ( .A1(\SB1_2_20/i0[10] ), .A2(\SB1_2_20/i0_3 ), .A3(
        \SB1_2_20/i0[6] ), .ZN(\SB1_2_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U7900 ( .A1(\SB2_2_18/i0_0 ), .A2(\SB2_2_18/i1_5 ), .A3(
        \SB2_2_18/i0_4 ), .ZN(\SB2_2_18/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U7902 ( .A1(\SB1_4_4/i0[10] ), .A2(\SB1_4_4/i0_0 ), .A3(
        \SB1_4_4/i0[6] ), .ZN(\SB1_4_4/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U7903 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[41] ), .A2(\RI5[2][77] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[167] ) );
  NAND3_X2 U7904 ( .A1(\SB1_4_10/i0[10] ), .A2(\RI1[4][131] ), .A3(
        \SB1_4_10/i0[6] ), .ZN(\SB1_4_10/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U7914 ( .A1(\MC_ARK_ARC_1_3/temp2[110] ), .A2(n2632), .Z(
        \MC_ARK_ARC_1_3/temp5[110] ) );
  XOR2_X1 U7915 ( .A1(\RI5[3][104] ), .A2(\RI5[3][110] ), .Z(n2632) );
  XOR2_X1 U7916 ( .A1(\RI5[1][165] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[189] ), 
        .Z(n2633) );
  NAND4_X2 U7918 ( .A1(\SB2_3_6/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_6/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_6/Component_Function_4/NAND4_in[1] ), .A4(n2634), .ZN(
        \SB2_3_6/buf_output[4] ) );
  XOR2_X1 U7920 ( .A1(n2635), .A2(n2636), .Z(\MC_ARK_ARC_1_3/buf_output[90] )
         );
  XOR2_X1 U7921 ( .A1(\MC_ARK_ARC_1_3/temp2[90] ), .A2(
        \MC_ARK_ARC_1_3/temp3[90] ), .Z(n2635) );
  XOR2_X1 U7922 ( .A1(\MC_ARK_ARC_1_3/temp1[90] ), .A2(
        \MC_ARK_ARC_1_3/temp4[90] ), .Z(n2636) );
  NAND3_X2 U7923 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i1[9] ), .A3(
        \SB2_2_24/i0_4 ), .ZN(\SB2_2_24/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7924 ( .A1(\RI5[3][160] ), .A2(\RI5[3][4] ), .Z(
        \MC_ARK_ARC_1_3/temp3[94] ) );
  XOR2_X1 U7935 ( .A1(\MC_ARK_ARC_1_1/temp4[87] ), .A2(
        \MC_ARK_ARC_1_1/temp3[87] ), .Z(\MC_ARK_ARC_1_1/temp6[87] ) );
  NAND3_X1 U7939 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i0[10] ), .A3(
        \SB1_2_31/i0_4 ), .ZN(n2642) );
  NAND4_X2 U7950 ( .A1(\SB1_0_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_12/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_12/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_12/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][144] ) );
  NAND3_X1 U7954 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i0_4 ), .A3(\SB4_31/i1_5 ), 
        .ZN(n2649) );
  XOR2_X1 U7957 ( .A1(\RI5[4][136] ), .A2(\RI5[4][142] ), .Z(
        \MC_ARK_ARC_1_4/temp1[142] ) );
  XOR2_X1 U7959 ( .A1(\RI5[2][169] ), .A2(\RI5[2][13] ), .Z(n2651) );
  NAND3_X1 U7960 ( .A1(\SB2_4_1/i0[9] ), .A2(n6277), .A3(\SB2_4_1/i0[6] ), 
        .ZN(\SB2_4_1/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U7962 ( .A1(\MC_ARK_ARC_1_3/temp3[73] ), .A2(
        \MC_ARK_ARC_1_3/temp4[73] ), .Z(n2652) );
  INV_X2 U7964 ( .I(\SB1_1_21/buf_output[5] ), .ZN(\SB2_1_21/i1_5 ) );
  XOR2_X1 U7965 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[102] ), .A2(\RI5[3][108] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[108] ) );
  NAND3_X2 U7967 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i1[9] ), .A3(
        \SB2_2_22/i0_4 ), .ZN(\SB2_2_22/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7968 ( .A1(\MC_ARK_ARC_1_1/temp6[72] ), .A2(
        \MC_ARK_ARC_1_1/temp5[72] ), .Z(\MC_ARK_ARC_1_1/buf_output[72] ) );
  BUF_X4 U7969 ( .I(\SB2_2_27/buf_output[2] ), .Z(\RI5[2][44] ) );
  NAND3_X1 U7970 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i1_5 ), .A3(
        \SB2_0_4/i1[9] ), .ZN(\SB2_0_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U7973 ( .A1(\SB2_4_8/i0_3 ), .A2(\SB2_4_8/i0[10] ), .A3(
        \SB2_4_8/i0[9] ), .ZN(n2655) );
  XOR2_X1 U7974 ( .A1(\MC_ARK_ARC_1_4/temp4[127] ), .A2(
        \MC_ARK_ARC_1_4/temp3[127] ), .Z(\MC_ARK_ARC_1_4/temp6[127] ) );
  XOR2_X1 U7975 ( .A1(\MC_ARK_ARC_1_1/temp6[70] ), .A2(
        \MC_ARK_ARC_1_1/temp5[70] ), .Z(\MC_ARK_ARC_1_1/buf_output[70] ) );
  INV_X4 U7978 ( .I(n2657), .ZN(\SB2_0_29/i0_4 ) );
  BUF_X4 U7983 ( .I(\SB2_2_20/buf_output[3] ), .Z(\RI5[2][81] ) );
  NAND3_X1 U7985 ( .A1(\SB1_0_7/i0_0 ), .A2(\SB1_0_7/i0[9] ), .A3(
        \SB1_0_7/i0[8] ), .ZN(\SB1_0_7/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U7986 ( .A1(\MC_ARK_ARC_1_1/temp5[78] ), .A2(n2661), .Z(
        \MC_ARK_ARC_1_1/buf_output[78] ) );
  XOR2_X1 U7987 ( .A1(\MC_ARK_ARC_1_1/temp3[78] ), .A2(
        \MC_ARK_ARC_1_1/temp4[78] ), .Z(n2661) );
  NAND3_X2 U7990 ( .A1(\SB2_0_18/i0_3 ), .A2(\RI3[0][82] ), .A3(
        \SB2_0_18/i1[9] ), .ZN(n2662) );
  BUF_X4 U7992 ( .I(\SB2_2_4/buf_output[3] ), .Z(\RI5[2][177] ) );
  NAND3_X1 U7994 ( .A1(\SB4_15/i0_3 ), .A2(\SB4_15/i0_4 ), .A3(\SB4_15/i1[9] ), 
        .ZN(n2664) );
  BUF_X4 U7996 ( .I(\SB2_3_30/buf_output[0] ), .Z(\RI5[3][36] ) );
  XOR2_X1 U7997 ( .A1(\RI5[2][108] ), .A2(\RI5[2][132] ), .Z(
        \MC_ARK_ARC_1_2/temp2[162] ) );
  XOR2_X1 U7998 ( .A1(n2668), .A2(\MC_ARK_ARC_1_2/temp5[6] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[6] ) );
  XOR2_X1 U7999 ( .A1(\MC_ARK_ARC_1_2/temp3[6] ), .A2(
        \MC_ARK_ARC_1_2/temp4[6] ), .Z(n2668) );
  XOR2_X1 U8005 ( .A1(\RI5[0][21] ), .A2(\RI5[0][57] ), .Z(
        \MC_ARK_ARC_1_0/temp3[147] ) );
  NAND3_X1 U8007 ( .A1(\SB4_7/i0_3 ), .A2(\SB4_7/i0[9] ), .A3(
        \SB3_9/buf_output[3] ), .ZN(n2673) );
  NAND3_X1 U8008 ( .A1(\SB4_7/i0_3 ), .A2(\SB4_7/i0_4 ), .A3(\SB4_7/i1[9] ), 
        .ZN(\SB4_7/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U8009 ( .I(\RI3[0][117] ), .ZN(\SB2_0_12/i0[8] ) );
  NAND3_X1 U8012 ( .A1(\SB4_30/i0[6] ), .A2(\SB4_30/i0[8] ), .A3(
        \SB4_30/i0[7] ), .ZN(\SB4_30/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U8016 ( .A1(\MC_ARK_ARC_1_0/temp2[150] ), .A2(n2680), .Z(
        \MC_ARK_ARC_1_0/temp5[150] ) );
  XOR2_X1 U8017 ( .A1(\RI5[0][144] ), .A2(\RI5[0][150] ), .Z(n2680) );
  NAND4_X1 U8019 ( .A1(\SB2_0_12/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_12/Component_Function_0/NAND4_in[0] ), .A3(n2682), .A4(
        \SB2_0_12/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_0_12/buf_output[0] ) );
  XOR2_X1 U8033 ( .A1(\MC_ARK_ARC_1_2/temp1[61] ), .A2(
        \MC_ARK_ARC_1_2/temp2[61] ), .Z(\MC_ARK_ARC_1_2/temp5[61] ) );
  NAND4_X2 U8039 ( .A1(\SB1_0_14/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_14/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][127] ) );
  NAND3_X1 U8042 ( .A1(n3966), .A2(\SB4_23/i0_3 ), .A3(\SB4_23/i0[9] ), .ZN(
        n2695) );
  NAND4_X2 U8045 ( .A1(\SB2_3_22/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_22/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_22/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_22/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB2_3_22/buf_output[4] ) );
  NAND3_X1 U8047 ( .A1(\SB4_20/i0_0 ), .A2(\SB4_20/i0[10] ), .A3(
        \SB4_20/i0[6] ), .ZN(n2700) );
  XOR2_X1 U8051 ( .A1(\RI5[0][74] ), .A2(\RI5[0][80] ), .Z(n2703) );
  NAND4_X2 U8058 ( .A1(\SB1_3_22/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_22/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_22/Component_Function_1/NAND4_in[0] ), .A4(n2713), .ZN(
        \SB1_3_22/buf_output[1] ) );
  NAND3_X2 U8060 ( .A1(\SB1_2_3/i0[10] ), .A2(\SB1_2_3/i1[9] ), .A3(
        \SB1_2_3/i1_7 ), .ZN(\SB1_2_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U8067 ( .A1(n232), .A2(n340), .A3(n275), .ZN(
        \SB1_0_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U8071 ( .A1(\SB2_0_29/i0[9] ), .A2(\SB2_0_29/i0_4 ), .A3(
        \SB2_0_29/i0[6] ), .ZN(\SB2_0_29/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U8075 ( .A1(\SB1_0_11/i0_0 ), .A2(\SB1_0_11/i3[0] ), .A3(
        \SB1_0_11/i1_7 ), .ZN(\SB1_0_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U8077 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i0_0 ), .A3(\SB4_5/i0[6] ), 
        .ZN(\SB4_5/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U8078 ( .I(\SB2_4_9/buf_output[0] ), .Z(\RI5[4][162] ) );
  XOR2_X1 U8081 ( .A1(\MC_ARK_ARC_1_4/temp5[126] ), .A2(n2730), .Z(
        \MC_ARK_ARC_1_4/buf_output[126] ) );
  XOR2_X1 U8082 ( .A1(\MC_ARK_ARC_1_4/temp3[126] ), .A2(
        \MC_ARK_ARC_1_4/temp4[126] ), .Z(n2730) );
  NAND4_X2 U8083 ( .A1(\SB2_4_10/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_4_10/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_4_10/Component_Function_3/NAND4_in[1] ), .A4(n2731), .ZN(
        \SB2_4_10/buf_output[3] ) );
  NAND4_X2 U8089 ( .A1(\SB3_14/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_14/Component_Function_1/NAND4_in[0] ), .A4(n2735), .ZN(
        \SB3_14/buf_output[1] ) );
  NAND3_X1 U8092 ( .A1(\SB1_0_6/i0_4 ), .A2(\SB1_0_6/i1_7 ), .A3(
        \SB1_0_6/i0[8] ), .ZN(n2738) );
  BUF_X4 U8093 ( .I(\SB2_2_8/buf_output[1] ), .Z(\RI5[2][163] ) );
  NAND3_X1 U8098 ( .A1(\SB1_3_3/i0[6] ), .A2(\SB1_3_3/i1[9] ), .A3(
        \SB1_3_3/i0_3 ), .ZN(\SB1_3_3/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U8100 ( .A1(\SB1_0_23/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_23/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_0_23/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_23/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][78] ) );
  XOR2_X1 U8102 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[25] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[61] ), .Z(\MC_ARK_ARC_1_2/temp3[151] )
         );
  XOR2_X1 U8106 ( .A1(n2746), .A2(\MC_ARK_ARC_1_4/temp2[26] ), .Z(
        \MC_ARK_ARC_1_4/temp5[26] ) );
  XOR2_X1 U8107 ( .A1(\RI5[4][20] ), .A2(\RI5[4][26] ), .Z(n2746) );
  XOR2_X1 U8108 ( .A1(n2747), .A2(\MC_ARK_ARC_1_3/temp5[99] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[99] ) );
  BUF_X4 U8117 ( .I(\SB2_2_30/buf_output[2] ), .Z(\RI5[2][26] ) );
  NAND3_X1 U8119 ( .A1(\SB1_1_20/i0[6] ), .A2(\SB1_1_20/i1[9] ), .A3(
        \SB1_1_20/i0_3 ), .ZN(\SB1_1_20/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U8123 ( .A1(n2753), .A2(\MC_ARK_ARC_1_4/temp5[119] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[119] ) );
  XOR2_X1 U8124 ( .A1(\MC_ARK_ARC_1_4/temp3[119] ), .A2(
        \MC_ARK_ARC_1_4/temp4[119] ), .Z(n2753) );
  XOR2_X1 U8125 ( .A1(\RI5[2][8] ), .A2(\RI5[2][44] ), .Z(
        \MC_ARK_ARC_1_2/temp3[134] ) );
  NOR2_X2 U8135 ( .A1(n2756), .A2(n2755), .ZN(\SB2_1_4/i1_7 ) );
  XOR2_X1 U8140 ( .A1(\MC_ARK_ARC_1_1/temp6[150] ), .A2(
        \MC_ARK_ARC_1_1/temp5[150] ), .Z(\MC_ARK_ARC_1_1/buf_output[150] ) );
  XOR2_X1 U8142 ( .A1(\RI5[3][47] ), .A2(n27), .Z(n2759) );
  XOR2_X1 U8143 ( .A1(n2761), .A2(\MC_ARK_ARC_1_1/temp6[15] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[15] ) );
  NAND3_X2 U8145 ( .A1(\SB2_2_13/i0_3 ), .A2(\SB2_2_13/i1[9] ), .A3(
        \SB2_2_13/i0_4 ), .ZN(\SB2_2_13/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8146 ( .A1(\RI5[1][63] ), .A2(\RI5[1][69] ), .Z(
        \MC_ARK_ARC_1_1/temp1[69] ) );
  XOR2_X1 U8150 ( .A1(n2768), .A2(\MC_ARK_ARC_1_0/temp1[146] ), .Z(
        \MC_ARK_ARC_1_0/temp5[146] ) );
  XOR2_X1 U8151 ( .A1(\RI5[0][116] ), .A2(\RI5[0][92] ), .Z(n2768) );
  BUF_X4 U8152 ( .I(\SB2_0_20/buf_output[3] ), .Z(\RI5[0][81] ) );
  XOR2_X1 U8154 ( .A1(\MC_ARK_ARC_1_0/temp3[90] ), .A2(
        \MC_ARK_ARC_1_0/temp4[90] ), .Z(n2771) );
  XOR2_X1 U8155 ( .A1(\MC_ARK_ARC_1_4/temp3[30] ), .A2(
        \MC_ARK_ARC_1_4/temp4[30] ), .Z(\MC_ARK_ARC_1_4/temp6[30] ) );
  NAND4_X2 U8156 ( .A1(\SB1_0_8/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_8/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][163] ) );
  BUF_X4 U8157 ( .I(\SB2_3_14/buf_output[2] ), .Z(\RI5[3][122] ) );
  NAND3_X1 U8158 ( .A1(\SB1_0_27/i0_0 ), .A2(\SB1_0_27/i3[0] ), .A3(
        \SB1_0_27/i1_7 ), .ZN(\SB1_0_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U8159 ( .A1(\SB1_0_0/i0_4 ), .A2(\SB1_0_0/i0_0 ), .A3(
        \SB1_0_0/i1_5 ), .ZN(n2772) );
  XOR2_X1 U8161 ( .A1(\MC_ARK_ARC_1_2/temp3[160] ), .A2(
        \MC_ARK_ARC_1_2/temp4[160] ), .Z(\MC_ARK_ARC_1_2/temp6[160] ) );
  XOR2_X1 U8162 ( .A1(n2779), .A2(\MC_ARK_ARC_1_4/temp6[33] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[33] ) );
  XOR2_X1 U8164 ( .A1(\MC_ARK_ARC_1_4/temp6[99] ), .A2(n2780), .Z(
        \MC_ARK_ARC_1_4/buf_output[99] ) );
  XOR2_X1 U8165 ( .A1(n2781), .A2(n56), .Z(Ciphertext[186]) );
  XOR2_X1 U8172 ( .A1(\RI5[0][135] ), .A2(\RI5[0][141] ), .Z(
        \MC_ARK_ARC_1_0/temp1[141] ) );
  NAND3_X1 U8178 ( .A1(\SB4_3/i0_4 ), .A2(\SB4_3/i1[9] ), .A3(\SB4_3/i1_5 ), 
        .ZN(n2789) );
  NAND4_X2 U8181 ( .A1(\SB1_0_7/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_7/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_7/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_0_7/Component_Function_1/NAND4_in[2] ), .ZN(\RI3[0][169] ) );
  NAND4_X2 U8182 ( .A1(\SB1_0_17/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_17/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_0_17/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_17/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][114] ) );
  NAND3_X1 U8186 ( .A1(\SB4_12/i0[10] ), .A2(\SB4_12/i1[9] ), .A3(
        \SB4_12/i1_7 ), .ZN(n2791) );
  NAND3_X1 U8187 ( .A1(\SB2_4_23/i0[9] ), .A2(\SB2_4_23/i1_5 ), .A3(
        \SB2_4_23/i0[6] ), .ZN(\SB2_4_23/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U8191 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[43] ), .A2(\RI5[4][67] ), 
        .Z(n2795) );
  XOR2_X1 U8196 ( .A1(\MC_ARK_ARC_1_2/temp3[89] ), .A2(
        \MC_ARK_ARC_1_2/temp4[89] ), .Z(n2803) );
  NAND4_X2 U8200 ( .A1(\SB1_2_31/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_31/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_31/Component_Function_4/NAND4_in[3] ), .A4(n2805), .ZN(
        \SB1_2_31/buf_output[4] ) );
  XOR2_X1 U8201 ( .A1(\MC_ARK_ARC_1_3/temp4[109] ), .A2(
        \MC_ARK_ARC_1_3/temp3[109] ), .Z(n2806) );
  XOR2_X1 U8202 ( .A1(\MC_ARK_ARC_1_0/temp1[169] ), .A2(
        \MC_ARK_ARC_1_0/temp2[169] ), .Z(\MC_ARK_ARC_1_0/temp5[169] ) );
  INV_X2 U8209 ( .I(\SB1_1_14/buf_output[2] ), .ZN(\SB2_1_11/i1[9] ) );
  NAND4_X2 U8210 ( .A1(\SB1_1_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_14/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_14/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_1_14/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_1_14/buf_output[2] ) );
  NAND3_X1 U8212 ( .A1(\SB4_10/i0[8] ), .A2(\SB4_10/i1_5 ), .A3(\SB4_10/i3[0] ), .ZN(\SB4_10/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U8213 ( .A1(\MC_ARK_ARC_1_3/temp6[66] ), .A2(
        \MC_ARK_ARC_1_3/temp5[66] ), .Z(\MC_ARK_ARC_1_3/buf_output[66] ) );
  XOR2_X1 U8216 ( .A1(\MC_ARK_ARC_1_4/temp4[5] ), .A2(n3007), .Z(
        \MC_ARK_ARC_1_4/temp6[5] ) );
  NAND3_X2 U8218 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i0[10] ), .A3(
        \SB2_1_4/i0[9] ), .ZN(\SB2_1_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U8219 ( .A1(\SB1_4_0/i0_3 ), .A2(\SB1_4_0/i0[9] ), .A3(
        \SB1_4_0/i0[10] ), .ZN(\SB1_4_0/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U8221 ( .A1(\MC_ARK_ARC_1_4/temp1[67] ), .A2(
        \MC_ARK_ARC_1_4/temp2[67] ), .Z(\MC_ARK_ARC_1_4/temp5[67] ) );
  BUF_X4 U8222 ( .I(\SB2_4_29/buf_output[1] ), .Z(\RI5[4][37] ) );
  XOR2_X1 U8223 ( .A1(\RI5[1][148] ), .A2(\RI5[1][184] ), .Z(
        \MC_ARK_ARC_1_1/temp3[82] ) );
  XOR2_X1 U8229 ( .A1(\MC_ARK_ARC_1_2/temp5[100] ), .A2(n2814), .Z(
        \MC_ARK_ARC_1_2/buf_output[100] ) );
  NAND4_X2 U8230 ( .A1(n2986), .A2(\SB2_1_4/Component_Function_3/NAND4_in[1] ), 
        .A3(\SB2_1_4/Component_Function_3/NAND4_in[3] ), .A4(n2815), .ZN(
        \SB2_1_4/buf_output[3] ) );
  NAND3_X1 U8231 ( .A1(\SB1_0_8/i0_4 ), .A2(\SB1_0_8/i0[9] ), .A3(
        \SB1_0_8/i0[6] ), .ZN(n2816) );
  XOR2_X1 U8234 ( .A1(\MC_ARK_ARC_1_2/temp4[2] ), .A2(
        \MC_ARK_ARC_1_2/temp3[2] ), .Z(n2819) );
  NAND4_X2 U8239 ( .A1(\SB2_3_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_19/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_19/Component_Function_4/NAND4_in[1] ), .A4(n2823), .ZN(
        \SB2_3_19/buf_output[4] ) );
  XOR2_X1 U8245 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[83] ), .A2(\RI5[1][119] ), 
        .Z(n2827) );
  NAND3_X1 U8246 ( .A1(\SB4_17/i0_0 ), .A2(\SB4_17/i3[0] ), .A3(\SB4_17/i1_7 ), 
        .ZN(n2828) );
  BUF_X4 U8248 ( .I(\SB2_2_10/buf_output[0] ), .Z(\RI5[2][156] ) );
  NAND4_X2 U8251 ( .A1(\SB1_1_4/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_4/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_1_4/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_1_4/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_4/buf_output[0] ) );
  XOR2_X1 U8253 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[100] ), .A2(\RI5[2][136] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[34] ) );
  BUF_X4 U8254 ( .I(\SB2_2_30/buf_output[3] ), .Z(\RI5[2][21] ) );
  XOR2_X1 U8255 ( .A1(\MC_ARK_ARC_1_0/temp3[42] ), .A2(
        \MC_ARK_ARC_1_0/temp4[42] ), .Z(n2832) );
  NAND3_X1 U8256 ( .A1(\SB2_0_9/i0[10] ), .A2(\SB2_0_9/i1[9] ), .A3(
        \SB2_0_9/i1_7 ), .ZN(n2835) );
  XOR2_X1 U8259 ( .A1(n2837), .A2(\MC_ARK_ARC_1_3/temp1[92] ), .Z(
        \MC_ARK_ARC_1_3/temp5[92] ) );
  NAND3_X1 U8261 ( .A1(\SB1_0_5/i1[9] ), .A2(\SB1_0_5/i0[10] ), .A3(
        \SB1_0_5/i1_5 ), .ZN(\SB1_0_5/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U8262 ( .A1(\RI5[0][179] ), .A2(\RI5[0][23] ), .Z(
        \MC_ARK_ARC_1_0/temp3[113] ) );
  XOR2_X1 U8265 ( .A1(\MC_ARK_ARC_1_0/temp2[128] ), .A2(
        \MC_ARK_ARC_1_0/temp1[128] ), .Z(\MC_ARK_ARC_1_0/temp5[128] ) );
  XOR2_X1 U8266 ( .A1(\MC_ARK_ARC_1_3/temp5[12] ), .A2(n2838), .Z(
        \MC_ARK_ARC_1_3/buf_output[12] ) );
  XOR2_X1 U8267 ( .A1(\MC_ARK_ARC_1_3/temp4[12] ), .A2(
        \MC_ARK_ARC_1_3/temp3[12] ), .Z(n2838) );
  NAND3_X2 U8270 ( .A1(\SB1_0_20/i0[10] ), .A2(\SB1_0_20/i1[9] ), .A3(
        \SB1_0_20/i1_7 ), .ZN(\SB1_0_20/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U8272 ( .A1(\MC_ARK_ARC_1_2/temp5[58] ), .A2(n2841), .Z(
        \MC_ARK_ARC_1_2/buf_output[58] ) );
  XOR2_X1 U8273 ( .A1(\MC_ARK_ARC_1_2/temp3[58] ), .A2(
        \MC_ARK_ARC_1_2/temp4[58] ), .Z(n2841) );
  BUF_X4 U8274 ( .I(\SB2_3_18/buf_output[1] ), .Z(\RI5[3][103] ) );
  NAND2_X2 U8276 ( .A1(n2843), .A2(n2842), .ZN(\SB2_0_14/i0[6] ) );
  XOR2_X1 U8278 ( .A1(n2845), .A2(n2846), .Z(\MC_ARK_ARC_1_3/buf_output[95] )
         );
  XOR2_X1 U8281 ( .A1(\RI5[4][83] ), .A2(\RI5[4][119] ), .Z(n2847) );
  NAND3_X2 U8286 ( .A1(\SB2_3_21/i0[6] ), .A2(\RI3[3][64] ), .A3(
        \SB2_3_21/i0[9] ), .ZN(n2848) );
  NAND3_X2 U8288 ( .A1(\SB2_3_18/i0_0 ), .A2(\SB2_3_18/i0[10] ), .A3(
        \SB2_3_18/i0[6] ), .ZN(n2932) );
  NAND3_X2 U8290 ( .A1(\SB2_2_13/i0_3 ), .A2(\SB2_2_13/i0_0 ), .A3(
        \SB2_2_13/i0_4 ), .ZN(\SB2_2_13/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U8291 ( .A1(\MC_ARK_ARC_1_0/temp3[67] ), .A2(
        \MC_ARK_ARC_1_0/temp4[67] ), .Z(\MC_ARK_ARC_1_0/temp6[67] ) );
  XOR2_X1 U8295 ( .A1(\MC_ARK_ARC_1_2/temp2[168] ), .A2(
        \MC_ARK_ARC_1_2/temp1[168] ), .Z(n2852) );
  INV_X2 U8296 ( .I(n2854), .ZN(\RI1[5][185] ) );
  XNOR2_X1 U8297 ( .A1(\MC_ARK_ARC_1_4/temp6[185] ), .A2(
        \MC_ARK_ARC_1_4/temp5[185] ), .ZN(n2854) );
  XOR2_X1 U8298 ( .A1(\MC_ARK_ARC_1_4/temp3[115] ), .A2(
        \MC_ARK_ARC_1_4/temp4[115] ), .Z(n2855) );
  NAND3_X1 U8299 ( .A1(\SB2_3_22/i0[8] ), .A2(\RI3[3][58] ), .A3(
        \SB2_3_22/i1_7 ), .ZN(\SB2_3_22/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U8304 ( .A1(n2858), .A2(\MC_ARK_ARC_1_0/temp5[166] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[166] ) );
  NAND3_X1 U8306 ( .A1(\SB4_21/i0_3 ), .A2(\SB4_21/i0_4 ), .A3(n3998), .ZN(
        n2860) );
  NAND3_X1 U8317 ( .A1(\SB4_18/i0_3 ), .A2(\SB4_18/i0_0 ), .A3(\SB4_18/i0_4 ), 
        .ZN(\SB4_18/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U8320 ( .A1(\SB2_3_16/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_16/Component_Function_0/NAND4_in[0] ), .A3(n2870), .A4(n2869), 
        .ZN(\SB2_3_16/buf_output[0] ) );
  XOR2_X1 U8326 ( .A1(n2872), .A2(n121), .Z(Ciphertext[42]) );
  XOR2_X1 U8328 ( .A1(\RI5[0][120] ), .A2(\RI5[0][144] ), .Z(
        \MC_ARK_ARC_1_0/temp2[174] ) );
  BUF_X4 U8329 ( .I(\SB2_2_31/buf_output[3] ), .Z(\RI5[2][15] ) );
  BUF_X4 U8333 ( .I(\SB2_1_9/buf_output[1] ), .Z(\RI5[1][157] ) );
  NAND3_X1 U8336 ( .A1(\SB1_4_28/i0_3 ), .A2(\SB1_4_28/i0[10] ), .A3(
        \SB1_4_28/i0_4 ), .ZN(\SB1_4_28/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U8337 ( .A1(\SB1_3_21/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_21/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_21/Component_Function_1/NAND4_in[0] ), .A4(n2880), .ZN(
        \SB1_3_21/buf_output[1] ) );
  NAND3_X1 U8338 ( .A1(\SB4_31/i0_3 ), .A2(\SB4_31/i0_4 ), .A3(\SB4_31/i1[9] ), 
        .ZN(n2881) );
  XOR2_X1 U8339 ( .A1(\RI5[4][136] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[160] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[190] ) );
  NAND3_X1 U8340 ( .A1(\SB4_26/i0_3 ), .A2(\SB4_26/i0[10] ), .A3(
        \SB4_26/i0[9] ), .ZN(n2882) );
  XOR2_X1 U8345 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[156] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[0] ), .Z(\MC_ARK_ARC_1_3/temp3[90] ) );
  NAND3_X1 U8347 ( .A1(\SB1_3_13/i0[10] ), .A2(\SB1_3_13/i0[6] ), .A3(
        \SB1_3_13/i0_3 ), .ZN(\SB1_3_13/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U8348 ( .I(\SB1_1_6/buf_output[5] ), .ZN(\SB2_1_6/i1_5 ) );
  BUF_X4 U8349 ( .I(\SB2_1_6/buf_output[1] ), .Z(\RI5[1][175] ) );
  INV_X2 U8352 ( .I(n2887), .ZN(\RI1[5][89] ) );
  XNOR2_X1 U8353 ( .A1(\MC_ARK_ARC_1_4/temp5[89] ), .A2(n3001), .ZN(n2887) );
  XOR2_X1 U8357 ( .A1(\MC_ARK_ARC_1_1/temp1[112] ), .A2(
        \MC_ARK_ARC_1_1/temp2[112] ), .Z(n2891) );
  XOR2_X1 U8358 ( .A1(\RI5[0][93] ), .A2(\RI5[0][57] ), .Z(
        \MC_ARK_ARC_1_0/temp3[183] ) );
  NAND4_X2 U8360 ( .A1(\SB2_1_30/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_1_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_30/Component_Function_4/NAND4_in[0] ), .A4(n3086), .ZN(
        \SB2_1_30/buf_output[4] ) );
  NAND3_X2 U8361 ( .A1(\SB1_4_10/i0[10] ), .A2(\SB1_4_10/i0_0 ), .A3(
        \SB1_4_10/i0[6] ), .ZN(\SB1_4_10/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U8363 ( .A1(\SB3_11/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_1/NAND4_in[3] ), .A4(
        \SB3_11/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_11/buf_output[1] ) );
  INV_X2 U8368 ( .I(\RI3[0][147] ), .ZN(\SB2_0_7/i0[8] ) );
  XOR2_X1 U8369 ( .A1(\MC_ARK_ARC_1_2/temp5[66] ), .A2(n2893), .Z(
        \MC_ARK_ARC_1_2/buf_output[66] ) );
  NAND3_X2 U8377 ( .A1(\SB1_4_9/i0_3 ), .A2(\SB1_4_9/i1[9] ), .A3(
        \SB1_4_9/i0_4 ), .ZN(n2897) );
  INV_X2 U8381 ( .I(\SB1_1_28/buf_output[2] ), .ZN(\SB2_1_25/i1[9] ) );
  NAND3_X2 U8383 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i0_4 ), .A3(
        \SB1_1_15/i1[9] ), .ZN(n2903) );
  NAND3_X1 U8386 ( .A1(\SB1_4_16/i0_4 ), .A2(\SB1_4_16/i1_5 ), .A3(
        \SB1_4_16/i1[9] ), .ZN(n2905) );
  XOR2_X1 U8388 ( .A1(n2907), .A2(n144), .Z(Ciphertext[83]) );
  NAND4_X2 U8389 ( .A1(\SB4_18/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_18/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_18/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_18/Component_Function_5/NAND4_in[0] ), .ZN(n2907) );
  NAND4_X2 U8392 ( .A1(\SB2_1_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_27/Component_Function_0/NAND4_in[1] ), .A3(n2909), .A4(
        \SB2_1_27/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_27/buf_output[0] ) );
  XOR2_X1 U8397 ( .A1(\RI5[4][136] ), .A2(\RI5[4][172] ), .Z(
        \MC_ARK_ARC_1_4/temp3[70] ) );
  XOR2_X1 U8402 ( .A1(\MC_ARK_ARC_1_0/temp3[4] ), .A2(
        \MC_ARK_ARC_1_0/temp4[4] ), .Z(n2914) );
  NAND3_X1 U8405 ( .A1(\SB3_11/i0[9] ), .A2(\SB3_11/i0[6] ), .A3(\SB3_11/i1_5 ), .ZN(\SB3_11/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U8408 ( .A1(\RI5[3][25] ), .A2(\RI5[3][73] ), .Z(n2916) );
  XOR2_X1 U8409 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), .A2(\RI5[3][79] ), 
        .Z(n2917) );
  BUF_X4 U8410 ( .I(\SB2_1_2/buf_output[0] ), .Z(\RI5[1][12] ) );
  XOR2_X1 U8413 ( .A1(\MC_ARK_ARC_1_1/temp3[119] ), .A2(
        \MC_ARK_ARC_1_1/temp4[119] ), .Z(\MC_ARK_ARC_1_1/temp6[119] ) );
  BUF_X4 U8415 ( .I(\SB2_1_14/buf_output[1] ), .Z(\RI5[1][127] ) );
  XOR2_X1 U8419 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[20] ), .A2(\RI5[3][26] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[26] ) );
  XOR2_X1 U8420 ( .A1(\MC_ARK_ARC_1_4/temp2[98] ), .A2(
        \MC_ARK_ARC_1_4/temp1[98] ), .Z(\MC_ARK_ARC_1_4/temp5[98] ) );
  XOR2_X1 U8421 ( .A1(\MC_ARK_ARC_1_4/temp5[85] ), .A2(
        \MC_ARK_ARC_1_4/temp6[85] ), .Z(\MC_ARK_ARC_1_4/buf_output[85] ) );
  NAND3_X2 U8423 ( .A1(\SB1_4_8/i0_3 ), .A2(\SB1_4_8/i1[9] ), .A3(
        \SB1_4_8/i0_4 ), .ZN(n2927) );
  NAND4_X2 U8427 ( .A1(\SB1_1_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_2/Component_Function_0/NAND4_in[0] ), .A4(n2928), .ZN(
        \SB1_1_2/buf_output[0] ) );
  NAND3_X1 U8429 ( .A1(\SB3_25/i0_0 ), .A2(\SB3_25/i0_3 ), .A3(\SB3_25/i0[7] ), 
        .ZN(n2929) );
  XOR2_X1 U8430 ( .A1(\MC_ARK_ARC_1_4/temp4[87] ), .A2(n2930), .Z(n2933) );
  XOR2_X1 U8431 ( .A1(\RI5[4][153] ), .A2(\RI5[4][189] ), .Z(n2930) );
  NAND3_X1 U8432 ( .A1(\SB1_1_6/i0_0 ), .A2(\SB1_1_6/i1_7 ), .A3(
        \SB1_1_6/i3[0] ), .ZN(\SB1_1_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U8433 ( .A1(\SB2_1_21/i0_0 ), .A2(\SB2_1_21/i0_4 ), .A3(
        \SB2_1_21/i1_5 ), .ZN(n2931) );
  NAND3_X1 U8444 ( .A1(\SB4_26/i0_4 ), .A2(n573), .A3(\SB4_26/i1_5 ), .ZN(
        n2938) );
  XOR2_X1 U8446 ( .A1(\MC_ARK_ARC_1_0/temp1[74] ), .A2(n2939), .Z(
        \MC_ARK_ARC_1_0/temp5[74] ) );
  XOR2_X1 U8447 ( .A1(\RI5[0][20] ), .A2(\RI5[0][44] ), .Z(n2939) );
  XOR2_X1 U8453 ( .A1(\MC_ARK_ARC_1_1/temp2[10] ), .A2(
        \MC_ARK_ARC_1_1/temp1[10] ), .Z(\MC_ARK_ARC_1_1/temp5[10] ) );
  XOR2_X1 U8454 ( .A1(\MC_ARK_ARC_1_1/temp1[178] ), .A2(
        \MC_ARK_ARC_1_1/temp2[178] ), .Z(\MC_ARK_ARC_1_1/temp5[178] ) );
  XOR2_X1 U8455 ( .A1(\MC_ARK_ARC_1_4/temp3[26] ), .A2(
        \MC_ARK_ARC_1_4/temp4[26] ), .Z(n3139) );
  NOR2_X2 U8457 ( .A1(n2945), .A2(n3180), .ZN(n2943) );
  AND2_X1 U8459 ( .A1(\SB1_0_20/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_0_20/Component_Function_3/NAND4_in[3] ), .Z(n2946) );
  XOR2_X1 U8460 ( .A1(\MC_ARK_ARC_1_1/temp6[136] ), .A2(
        \MC_ARK_ARC_1_1/temp5[136] ), .Z(\MC_ARK_ARC_1_1/buf_output[136] ) );
  XOR2_X1 U8464 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[14] ), .A2(\RI5[2][38] ), 
        .Z(n2948) );
  XOR2_X1 U8465 ( .A1(\MC_ARK_ARC_1_1/temp5[125] ), .A2(
        \MC_ARK_ARC_1_1/temp6[125] ), .Z(\RI1[2][125] ) );
  XOR2_X1 U8470 ( .A1(\MC_ARK_ARC_1_0/temp3[44] ), .A2(
        \MC_ARK_ARC_1_0/temp4[44] ), .Z(n2952) );
  XOR2_X1 U8477 ( .A1(\SB2_3_29/buf_output[5] ), .A2(\RI5[3][41] ), .Z(
        \MC_ARK_ARC_1_3/temp2[71] ) );
  BUF_X4 U8485 ( .I(\SB2_1_25/buf_output[2] ), .Z(\RI5[1][56] ) );
  XOR2_X1 U8487 ( .A1(n2962), .A2(\MC_ARK_ARC_1_0/temp5[18] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[18] ) );
  XOR2_X1 U8488 ( .A1(\MC_ARK_ARC_1_0/temp3[18] ), .A2(
        \MC_ARK_ARC_1_0/temp4[18] ), .Z(n2962) );
  NAND3_X2 U8489 ( .A1(\SB2_1_19/i0_3 ), .A2(\SB2_1_19/i1[9] ), .A3(
        \SB2_1_19/i0_4 ), .ZN(n2963) );
  NAND3_X1 U8491 ( .A1(\SB4_0/i0_3 ), .A2(\SB4_0/i0_0 ), .A3(\SB4_0/i0[7] ), 
        .ZN(n2966) );
  NAND3_X1 U8492 ( .A1(\SB1_3_1/i0_0 ), .A2(\SB1_3_1/i3[0] ), .A3(
        \SB1_3_1/i1_7 ), .ZN(\SB1_3_1/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U8494 ( .A1(\SB1_3_1/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_1/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_3_1/Component_Function_0/NAND4_in[1] ), .A4(n2971), .ZN(
        \SB1_3_1/buf_output[0] ) );
  XOR2_X1 U8499 ( .A1(\MC_ARK_ARC_1_3/temp3[164] ), .A2(
        \MC_ARK_ARC_1_3/temp4[164] ), .Z(\MC_ARK_ARC_1_3/temp6[164] ) );
  NAND3_X1 U8502 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i0_3 ), .A3(\SB4_11/i0_4 ), .ZN(\SB4_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U8503 ( .A1(n1763), .A2(\SB2_3_22/i0[8] ), .A3(\SB2_3_22/i0[6] ), 
        .ZN(\SB2_3_22/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U8512 ( .A1(n2982), .A2(\MC_ARK_ARC_1_4/temp6[190] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[190] ) );
  XOR2_X1 U8513 ( .A1(\MC_ARK_ARC_1_4/temp1[190] ), .A2(
        \MC_ARK_ARC_1_4/temp2[190] ), .Z(n2982) );
  NAND3_X1 U8515 ( .A1(\SB2_4_12/i0[10] ), .A2(\SB2_4_12/i0_3 ), .A3(
        \SB2_4_12/i0[9] ), .ZN(\SB2_4_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U8516 ( .A1(\RI1[1][149] ), .A2(\SB1_1_7/i1[9] ), .A3(
        \SB1_1_7/i0_4 ), .ZN(\SB1_1_7/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8517 ( .A1(\MC_ARK_ARC_1_0/temp5[30] ), .A2(n2987), .Z(
        \MC_ARK_ARC_1_0/buf_output[30] ) );
  XOR2_X1 U8518 ( .A1(\MC_ARK_ARC_1_1/temp5[10] ), .A2(n2988), .Z(
        \MC_ARK_ARC_1_1/buf_output[10] ) );
  XOR2_X1 U8519 ( .A1(\MC_ARK_ARC_1_1/temp3[10] ), .A2(
        \MC_ARK_ARC_1_1/temp4[10] ), .Z(n2988) );
  XOR2_X1 U8520 ( .A1(\RI5[2][71] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[35] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[161] ) );
  NAND4_X2 U8521 ( .A1(\SB1_1_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_7/Component_Function_0/NAND4_in[0] ), .A4(n2989), .ZN(
        \SB1_1_7/buf_output[0] ) );
  NAND3_X1 U8527 ( .A1(\SB4_19/i0_0 ), .A2(\SB4_19/i3[0] ), .A3(\SB4_19/i1_7 ), 
        .ZN(\SB4_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U8528 ( .A1(\SB2_3_6/i0_3 ), .A2(\SB2_3_6/i1[9] ), .A3(
        \SB2_3_6/i0_4 ), .ZN(\SB2_3_6/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8531 ( .A1(\SB2_2_22/buf_output[3] ), .A2(\RI5[2][105] ), .Z(
        \MC_ARK_ARC_1_2/temp3[3] ) );
  XOR2_X1 U8533 ( .A1(n3078), .A2(\MC_ARK_ARC_1_0/temp1[23] ), .Z(
        \MC_ARK_ARC_1_0/temp5[23] ) );
  NAND3_X2 U8534 ( .A1(\RI1[4][155] ), .A2(\SB1_4_6/i1[9] ), .A3(
        \SB1_4_6/i0_4 ), .ZN(n2997) );
  NAND3_X1 U8543 ( .A1(\SB1_0_29/i0_0 ), .A2(\SB1_0_29/i0[9] ), .A3(
        \SB1_0_29/i0[8] ), .ZN(\SB1_0_29/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U8545 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[171] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[3] ), .Z(n3004) );
  NAND3_X1 U8547 ( .A1(\SB3_9/buf_output[3] ), .A2(\SB4_7/i1[9] ), .A3(
        \SB4_7/i1_7 ), .ZN(n3006) );
  XOR2_X1 U8548 ( .A1(\RI5[4][107] ), .A2(\RI5[4][71] ), .Z(n3007) );
  XOR2_X1 U8555 ( .A1(\MC_ARK_ARC_1_2/temp3[39] ), .A2(
        \MC_ARK_ARC_1_2/temp4[39] ), .Z(n3011) );
  XOR2_X1 U8556 ( .A1(\RI5[3][65] ), .A2(\RI5[3][59] ), .Z(
        \MC_ARK_ARC_1_3/temp1[65] ) );
  XOR2_X1 U8557 ( .A1(\RI5[3][48] ), .A2(\RI5[3][72] ), .Z(
        \MC_ARK_ARC_1_3/temp2[102] ) );
  XOR2_X1 U8558 ( .A1(n3012), .A2(\MC_ARK_ARC_1_0/temp6[98] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[98] ) );
  NAND3_X1 U8559 ( .A1(\SB2_4_12/i0[10] ), .A2(\SB2_4_12/i1[9] ), .A3(
        \SB2_4_12/i1_7 ), .ZN(\SB2_4_12/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U8561 ( .I(\SB2_2_3/buf_output[2] ), .Z(\RI5[2][188] ) );
  BUF_X4 U8566 ( .I(\SB2_4_24/buf_output[5] ), .Z(\RI5[4][47] ) );
  NAND3_X1 U8568 ( .A1(\SB1_2_19/i0_0 ), .A2(\SB1_2_19/i1_5 ), .A3(
        \SB1_2_19/i0_4 ), .ZN(n3016) );
  BUF_X4 U8570 ( .I(\SB2_2_1/buf_output[4] ), .Z(\RI5[2][190] ) );
  XOR2_X1 U8573 ( .A1(n3018), .A2(n97), .Z(Ciphertext[89]) );
  NAND4_X2 U8574 ( .A1(\SB4_17/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_17/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_17/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_17/Component_Function_5/NAND4_in[0] ), .ZN(n3018) );
  NAND4_X2 U8576 ( .A1(\SB1_0_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_7/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_7/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_7/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][174] ) );
  NAND4_X2 U8577 ( .A1(\SB3_17/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_3/NAND4_in[0] ), .A4(n3020), .ZN(
        \SB3_17/buf_output[3] ) );
  XOR2_X1 U8580 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[143] ), .A2(\RI5[3][119] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[173] ) );
  NAND3_X1 U8582 ( .A1(\SB3_25/i0_0 ), .A2(\SB3_25/i3[0] ), .A3(\SB3_25/i1_7 ), 
        .ZN(\SB3_25/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U8583 ( .A1(\RI5[1][107] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[71] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[5] ) );
  XOR2_X1 U8585 ( .A1(\MC_ARK_ARC_1_4/temp3[128] ), .A2(
        \MC_ARK_ARC_1_4/temp4[128] ), .Z(\MC_ARK_ARC_1_4/temp6[128] ) );
  NAND4_X2 U8587 ( .A1(\SB3_29/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_29/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_29/Component_Function_4/NAND4_in[2] ), .A4(n3027), .ZN(
        \SB3_29/buf_output[4] ) );
  NAND3_X2 U8588 ( .A1(\SB2_2_18/i0_3 ), .A2(\SB2_2_18/i0_0 ), .A3(
        \SB2_2_18/i0_4 ), .ZN(\SB2_2_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U8592 ( .A1(\SB2_4_5/i1[9] ), .A2(\SB1_4_6/buf_output[4] ), .A3(
        \SB2_4_5/i1_5 ), .ZN(n3029) );
  XOR2_X1 U8593 ( .A1(\MC_ARK_ARC_1_1/temp6[160] ), .A2(n3030), .Z(
        \MC_ARK_ARC_1_1/buf_output[160] ) );
  XOR2_X1 U8594 ( .A1(\MC_ARK_ARC_1_1/temp2[160] ), .A2(
        \MC_ARK_ARC_1_1/temp1[160] ), .Z(n3030) );
  BUF_X4 U8600 ( .I(\SB2_2_30/buf_output[0] ), .Z(\RI5[2][36] ) );
  BUF_X4 U8602 ( .I(\SB2_4_18/buf_output[4] ), .Z(\RI5[4][88] ) );
  XOR2_X1 U8607 ( .A1(\RI5[4][137] ), .A2(\RI5[4][131] ), .Z(
        \MC_ARK_ARC_1_4/temp1[137] ) );
  NAND4_X2 U8609 ( .A1(\SB3_9/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_9/Component_Function_0/NAND4_in[3] ), .A3(
        \SB3_9/Component_Function_0/NAND4_in[1] ), .A4(
        \SB3_9/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_9/buf_output[0] )
         );
  NAND4_X2 U8610 ( .A1(\SB2_4_25/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_4_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_4_25/Component_Function_3/NAND4_in[0] ), .A4(n3039), .ZN(
        \SB2_4_25/buf_output[3] ) );
  NAND3_X1 U8614 ( .A1(\SB4_4/i0_4 ), .A2(\SB4_4/i1_7 ), .A3(\SB4_4/i0[8] ), 
        .ZN(\SB4_4/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U8621 ( .A1(\SB1_0_15/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_15/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_15/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_15/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][126] ) );
  XOR2_X1 U8626 ( .A1(\RI5[3][167] ), .A2(\RI5[3][173] ), .Z(
        \MC_ARK_ARC_1_3/temp1[173] ) );
  BUF_X4 U8628 ( .I(\SB2_4_22/buf_output[5] ), .Z(\RI5[4][59] ) );
  NAND3_X1 U8629 ( .A1(\SB3_1/i1_5 ), .A2(\SB3_1/i1[9] ), .A3(\SB3_1/i0_4 ), 
        .ZN(\SB3_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U8630 ( .A1(\SB4_0/i0_4 ), .A2(\SB4_0/i1_7 ), .A3(\SB4_0/i0[8] ), 
        .ZN(n3046) );
  XOR2_X1 U8635 ( .A1(\MC_ARK_ARC_1_2/temp2[32] ), .A2(
        \MC_ARK_ARC_1_2/temp3[32] ), .Z(n3049) );
  XOR2_X1 U8641 ( .A1(\MC_ARK_ARC_1_2/temp5[8] ), .A2(n3055), .Z(
        \MC_ARK_ARC_1_2/buf_output[8] ) );
  NAND3_X2 U8643 ( .A1(\SB2_0_16/i0_3 ), .A2(n594), .A3(\SB2_0_16/i1[9] ), 
        .ZN(\SB2_0_16/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8646 ( .A1(n3056), .A2(\MC_ARK_ARC_1_3/temp5[172] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[172] ) );
  XOR2_X1 U8647 ( .A1(\MC_ARK_ARC_1_3/temp3[172] ), .A2(
        \MC_ARK_ARC_1_3/temp4[172] ), .Z(n3056) );
  XOR2_X1 U8651 ( .A1(\MC_ARK_ARC_1_1/temp1[150] ), .A2(
        \MC_ARK_ARC_1_1/temp2[150] ), .Z(\MC_ARK_ARC_1_1/temp5[150] ) );
  NAND3_X1 U8654 ( .A1(\SB3_24/i0_3 ), .A2(\SB3_24/i0[10] ), .A3(\SB3_24/i0_4 ), .ZN(\SB3_24/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U8656 ( .A1(\SB1_0_1/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_1/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_1/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_1/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][18] ) );
  NAND3_X1 U8663 ( .A1(\SB3_5/i0[10] ), .A2(\SB3_5/i1[9] ), .A3(\SB3_5/i1_5 ), 
        .ZN(\SB3_5/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U8669 ( .A1(\SB1_4_31/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_4_31/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_4_31/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_4_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_4_31/buf_output[5] ) );
  XOR2_X1 U8670 ( .A1(\MC_ARK_ARC_1_4/temp5[59] ), .A2(
        \MC_ARK_ARC_1_4/temp6[59] ), .Z(\RI1[5][59] ) );
  NAND3_X1 U8674 ( .A1(\SB2_0_7/i0[8] ), .A2(\SB2_0_7/i1_7 ), .A3(
        \RI3[0][148] ), .ZN(\SB2_0_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U8675 ( .A1(\SB4_3/i0_4 ), .A2(\SB4_3/i1_7 ), .A3(\SB4_3/i0[8] ), 
        .ZN(\SB4_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U8683 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0[7] ), .A3(
        \SB2_1_23/i0_0 ), .ZN(\SB2_1_23/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U8685 ( .A1(\RI5[4][158] ), .A2(\RI5[4][182] ), .Z(n3079) );
  BUF_X4 U8688 ( .I(\SB2_4_25/buf_output[0] ), .Z(\RI5[4][66] ) );
  NAND3_X1 U8689 ( .A1(\SB1_1_21/i0_4 ), .A2(\SB1_1_21/i1_5 ), .A3(
        \SB1_1_21/i0_0 ), .ZN(n3083) );
  XOR2_X1 U8690 ( .A1(\MC_ARK_ARC_1_3/temp1[177] ), .A2(
        \MC_ARK_ARC_1_3/temp2[177] ), .Z(n3085) );
  NAND4_X2 U8691 ( .A1(\SB2_4_5/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_4_5/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_4_5/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_4_5/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_4_5/buf_output[2] ) );
  XOR2_X1 U8694 ( .A1(\MC_ARK_ARC_1_1/temp3[170] ), .A2(
        \MC_ARK_ARC_1_1/temp4[170] ), .Z(n3087) );
  XOR2_X1 U8695 ( .A1(\RI5[4][125] ), .A2(\RI5[4][149] ), .Z(n3088) );
  BUF_X4 U8696 ( .I(\SB2_2_31/buf_output[2] ), .Z(\RI5[2][20] ) );
  XOR2_X1 U8697 ( .A1(\MC_ARK_ARC_1_4/temp3[177] ), .A2(
        \MC_ARK_ARC_1_4/temp1[177] ), .Z(n3089) );
  XOR2_X1 U8698 ( .A1(\MC_ARK_ARC_1_4/temp2[177] ), .A2(
        \MC_ARK_ARC_1_4/temp4[177] ), .Z(n3090) );
  NAND3_X1 U8700 ( .A1(\SB1_1_1/i0[8] ), .A2(\SB1_1_1/i3[0] ), .A3(
        \SB1_1_1/i1_5 ), .ZN(n3092) );
  NAND3_X1 U8704 ( .A1(\SB3_17/buf_output[3] ), .A2(\SB4_15/i0_0 ), .A3(
        \SB4_15/i0[6] ), .ZN(\SB4_15/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U8705 ( .A1(\MC_ARK_ARC_1_2/temp5[77] ), .A2(n3094), .Z(
        \MC_ARK_ARC_1_2/buf_output[77] ) );
  XOR2_X1 U8706 ( .A1(\MC_ARK_ARC_1_2/temp3[77] ), .A2(
        \MC_ARK_ARC_1_2/temp4[77] ), .Z(n3094) );
  NAND3_X2 U8708 ( .A1(\SB2_4_4/i0_3 ), .A2(\SB2_4_4/i1[9] ), .A3(
        \SB2_4_4/i0_4 ), .ZN(n3097) );
  XNOR2_X1 U8714 ( .A1(\MC_ARK_ARC_1_2/temp6[28] ), .A2(
        \MC_ARK_ARC_1_2/temp5[28] ), .ZN(n3100) );
  NAND3_X1 U8716 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i0[8] ), .A3(\SB3_31/i1_7 ), 
        .ZN(\SB3_31/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U8717 ( .A1(\MC_ARK_ARC_1_4/temp1[70] ), .A2(
        \MC_ARK_ARC_1_4/temp2[70] ), .Z(\MC_ARK_ARC_1_4/temp5[70] ) );
  BUF_X4 U8720 ( .I(\SB2_3_19/buf_output[4] ), .Z(\RI5[3][82] ) );
  XOR2_X1 U8721 ( .A1(\MC_ARK_ARC_1_1/temp5[151] ), .A2(
        \MC_ARK_ARC_1_1/temp6[151] ), .Z(\MC_ARK_ARC_1_1/buf_output[151] ) );
  NAND4_X2 U8722 ( .A1(\SB1_0_23/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_23/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_23/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_0_23/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][53] ) );
  BUF_X4 U8725 ( .I(\SB2_1_16/buf_output[1] ), .Z(\RI5[1][115] ) );
  BUF_X4 U8728 ( .I(\SB2_1_27/buf_output[3] ), .Z(\RI5[1][39] ) );
  BUF_X4 U8729 ( .I(\SB2_3_13/buf_output[5] ), .Z(\RI5[3][113] ) );
  NAND3_X2 U8731 ( .A1(\SB1_1_28/i0_3 ), .A2(\SB1_1_28/i1[9] ), .A3(
        \SB1_1_28/i0_4 ), .ZN(n3107) );
  XOR2_X1 U8732 ( .A1(\RI5[1][68] ), .A2(\RI5[1][104] ), .Z(
        \MC_ARK_ARC_1_1/temp3[2] ) );
  NAND3_X2 U8734 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i1[9] ), .A3(
        \SB2_1_28/i0_4 ), .ZN(\SB2_1_28/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U8736 ( .I(\SB2_4_10/buf_output[0] ), .Z(\RI5[4][156] ) );
  NAND3_X1 U8737 ( .A1(\SB1_1_14/i0[10] ), .A2(\SB1_1_14/i0_3 ), .A3(
        \SB1_1_14/i0_4 ), .ZN(\SB1_1_14/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 U8740 ( .I(\SB2_4_21/buf_output[0] ), .Z(\RI5[4][90] ) );
  NAND3_X1 U8742 ( .A1(\SB3_14/i0_3 ), .A2(\SB3_14/i0[9] ), .A3(
        \SB3_14/i0[10] ), .ZN(\SB3_14/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U8749 ( .A1(\SB3_4/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_4/Component_Function_5/NAND4_in[0] ), .A3(
        \SB3_4/Component_Function_5/NAND4_in[3] ), .A4(n3118), .ZN(
        \SB3_4/buf_output[5] ) );
  BUF_X4 U8755 ( .I(\SB2_4_0/buf_output[5] ), .Z(\RI5[4][191] ) );
  NAND4_X2 U8758 ( .A1(\SB3_23/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_23/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[5][73] ) );
  INV_X2 U8763 ( .I(n3125), .ZN(\RI1[3][17] ) );
  BUF_X4 U8765 ( .I(\SB2_3_6/buf_output[0] ), .Z(\RI5[3][180] ) );
  INV_X1 U8769 ( .I(\SB3_31/buf_output[1] ), .ZN(\SB4_27/i1_7 ) );
  NAND4_X2 U8770 ( .A1(\SB3_31/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_31/buf_output[1] ) );
  XOR2_X1 U8778 ( .A1(\MC_ARK_ARC_1_1/temp3[190] ), .A2(
        \MC_ARK_ARC_1_1/temp4[190] ), .Z(n3133) );
  XOR2_X1 U8779 ( .A1(\MC_ARK_ARC_1_4/temp5[152] ), .A2(n3134), .Z(
        \MC_ARK_ARC_1_4/buf_output[152] ) );
  NAND3_X2 U8781 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i1[9] ), .A3(
        \SB2_2_28/i0_4 ), .ZN(\SB2_2_28/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8784 ( .A1(\MC_ARK_ARC_1_4/temp5[26] ), .A2(n3139), .Z(
        \MC_ARK_ARC_1_4/buf_output[26] ) );
  XOR2_X1 U8785 ( .A1(\MC_ARK_ARC_1_3/temp5[105] ), .A2(
        \MC_ARK_ARC_1_3/temp6[105] ), .Z(\RI1[4][105] ) );
  XOR2_X1 U8786 ( .A1(\MC_ARK_ARC_1_1/temp6[9] ), .A2(
        \MC_ARK_ARC_1_1/temp5[9] ), .Z(\RI1[2][9] ) );
  NAND3_X1 U8788 ( .A1(\SB1_4_16/i0_3 ), .A2(\SB1_4_16/i0_0 ), .A3(
        \SB1_4_16/i0_4 ), .ZN(\SB1_4_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U8789 ( .A1(n1499), .A2(\SB4_9/i3[0] ), .A3(\SB4_9/i1_5 ), .ZN(
        n3140) );
  BUF_X4 U8796 ( .I(\SB2_3_2/buf_output[0] ), .Z(\RI5[3][12] ) );
  XOR2_X1 U8800 ( .A1(\MC_ARK_ARC_1_4/temp3[159] ), .A2(
        \MC_ARK_ARC_1_4/temp4[159] ), .Z(n3148) );
  XOR2_X1 U8804 ( .A1(\RI5[1][77] ), .A2(\RI5[1][101] ), .Z(n3150) );
  NAND3_X2 U8809 ( .A1(\SB3_14/i0_3 ), .A2(\SB3_14/i1[9] ), .A3(\SB3_14/i0_4 ), 
        .ZN(\SB3_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U8810 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i1[9] ), .A3(
        \SB1_3_21/i0_4 ), .ZN(\SB1_3_21/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8819 ( .A1(\MC_ARK_ARC_1_4/temp3[170] ), .A2(
        \MC_ARK_ARC_1_4/temp4[170] ), .Z(n3159) );
  NAND3_X2 U8823 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i1[9] ), .A3(
        \SB2_1_23/i0_4 ), .ZN(n3161) );
  XOR2_X1 U8826 ( .A1(\MC_ARK_ARC_1_2/temp5[165] ), .A2(
        \MC_ARK_ARC_1_2/temp6[165] ), .Z(\RI1[3][165] ) );
  BUF_X4 U8829 ( .I(\SB2_3_16/buf_output[2] ), .Z(\RI5[3][110] ) );
  BUF_X4 U8830 ( .I(\SB2_2_7/buf_output[0] ), .Z(\RI5[2][174] ) );
  BUF_X4 U8831 ( .I(\SB2_3_12/buf_output[2] ), .Z(\RI5[3][134] ) );
  BUF_X4 U8832 ( .I(\SB2_4_5/buf_output[5] ), .Z(\RI5[4][161] ) );
  BUF_X4 U8833 ( .I(\SB2_4_6/buf_output[5] ), .Z(\RI5[4][155] ) );
  BUF_X4 U8835 ( .I(\SB2_1_2/buf_output[5] ), .Z(\RI5[1][179] ) );
  BUF_X4 U8836 ( .I(\SB2_2_29/buf_output[2] ), .Z(\RI5[2][32] ) );
  BUF_X4 U8837 ( .I(\SB2_1_6/buf_output[3] ), .Z(\RI5[1][165] ) );
  BUF_X4 U8839 ( .I(\SB2_4_4/buf_output[2] ), .Z(\RI5[4][182] ) );
  BUF_X4 U8840 ( .I(\SB2_2_3/buf_output[5] ), .Z(\RI5[2][173] ) );
  BUF_X4 U8841 ( .I(\SB2_3_2/buf_output[3] ), .Z(\RI5[3][189] ) );
  BUF_X4 U8842 ( .I(\SB2_3_7/buf_output[5] ), .Z(\RI5[3][149] ) );
  BUF_X4 U8843 ( .I(\SB2_0_19/buf_output[4] ), .Z(\RI5[0][82] ) );
  BUF_X4 U8846 ( .I(\SB2_0_17/buf_output[0] ), .Z(\RI5[0][114] ) );
  BUF_X4 U8847 ( .I(\SB2_0_17/buf_output[4] ), .Z(\RI5[0][94] ) );
  BUF_X4 U8848 ( .I(\SB2_0_17/buf_output[5] ), .Z(\RI5[0][89] ) );
  BUF_X4 U8850 ( .I(\SB2_0_18/buf_output[2] ), .Z(\RI5[0][98] ) );
  NAND4_X2 U8853 ( .A1(\SB1_1_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_1/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_1/buf_output[0] ) );
  BUF_X4 U8856 ( .I(\SB2_0_21/buf_output[0] ), .Z(\RI5[0][90] ) );
  BUF_X4 U8861 ( .I(\SB2_0_21/buf_output[1] ), .Z(\RI5[0][85] ) );
  NAND4_X2 U8862 ( .A1(\SB1_1_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_3/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_3/buf_output[0] ) );
  NAND4_X2 U8866 ( .A1(\SB1_1_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_13/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_13/buf_output[1] ) );
  NAND4_X2 U8867 ( .A1(\SB1_1_17/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_17/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_17/buf_output[0] ) );
  NAND4_X2 U8870 ( .A1(\SB1_1_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_29/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_29/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_1_29/buf_output[2] ) );
  NAND4_X2 U8876 ( .A1(\SB1_1_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_12/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_12/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_12/buf_output[4] ) );
  BUF_X4 U8882 ( .I(\SB2_0_21/buf_output[5] ), .Z(\RI5[0][65] ) );
  NAND4_X2 U8886 ( .A1(\SB1_1_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_10/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_10/buf_output[4] ) );
  NAND4_X2 U8888 ( .A1(\SB1_1_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_18/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_18/buf_output[1] ) );
  NAND4_X2 U8889 ( .A1(\SB1_1_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_25/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_25/buf_output[1] ) );
  NAND4_X2 U8891 ( .A1(\SB1_1_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_30/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_30/buf_output[0] ) );
  BUF_X4 U8895 ( .I(\SB2_1_3/buf_output[5] ), .Z(\RI5[1][173] ) );
  NAND4_X2 U8896 ( .A1(\SB2_1_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_0/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_0/buf_output[4] ) );
  NAND4_X2 U8897 ( .A1(\SB1_1_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_5/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_5/buf_output[0] ) );
  BUF_X4 U8899 ( .I(\SB2_1_1/buf_output[5] ), .Z(\RI5[1][185] ) );
  BUF_X4 U8901 ( .I(\SB2_1_4/buf_output[5] ), .Z(\RI5[1][167] ) );
  NAND4_X2 U8902 ( .A1(\SB1_1_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_5/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_5/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_5/buf_output[4] ) );
  BUF_X4 U8904 ( .I(\SB2_1_8/buf_output[5] ), .Z(\RI5[1][143] ) );
  BUF_X4 U8906 ( .I(\SB2_1_9/buf_output[5] ), .Z(\RI5[1][137] ) );
  BUF_X4 U8907 ( .I(\SB2_1_6/buf_output[5] ), .Z(\RI5[1][155] ) );
  BUF_X4 U8910 ( .I(\SB2_1_10/buf_output[5] ), .Z(\RI5[1][131] ) );
  BUF_X4 U8911 ( .I(\SB2_1_11/buf_output[2] ), .Z(\RI5[1][140] ) );
  BUF_X4 U8913 ( .I(\SB2_1_11/buf_output[4] ), .Z(\RI5[1][130] ) );
  BUF_X4 U8915 ( .I(\SB2_1_13/buf_output[1] ), .Z(\RI5[1][133] ) );
  BUF_X4 U8916 ( .I(\SB2_1_13/buf_output[2] ), .Z(\RI5[1][128] ) );
  BUF_X4 U8917 ( .I(\SB2_1_13/buf_output[0] ), .Z(\RI5[1][138] ) );
  BUF_X4 U8918 ( .I(\SB2_1_13/buf_output[5] ), .Z(\RI5[1][113] ) );
  BUF_X4 U8919 ( .I(\SB2_1_12/buf_output[5] ), .Z(\RI5[1][119] ) );
  NAND4_X2 U8921 ( .A1(\SB1_1_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_19/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_1_19/buf_output[2] ) );
  NAND4_X2 U8923 ( .A1(\SB1_1_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_19/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_19/buf_output[4] ) );
  BUF_X4 U8924 ( .I(\SB2_1_14/buf_output[4] ), .Z(\RI5[1][112] ) );
  BUF_X4 U8925 ( .I(\SB2_1_14/buf_output[5] ), .Z(\RI5[1][107] ) );
  NAND4_X2 U8926 ( .A1(\SB1_1_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_19/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_19/buf_output[0] ) );
  BUF_X4 U8928 ( .I(\SB2_1_17/buf_output[2] ), .Z(\RI5[1][104] ) );
  BUF_X4 U8929 ( .I(\SB2_1_17/buf_output[3] ), .Z(\RI5[1][99] ) );
  BUF_X4 U8931 ( .I(\SB2_1_18/buf_output[4] ), .Z(\RI5[1][88] ) );
  NAND4_X2 U8932 ( .A1(\SB1_1_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_20/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_20/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_20/buf_output[3] ) );
  BUF_X4 U8934 ( .I(\SB2_1_15/buf_output[2] ), .Z(\RI5[1][116] ) );
  BUF_X4 U8935 ( .I(\SB2_1_15/buf_output[0] ), .Z(\RI5[1][126] ) );
  NAND4_X2 U8936 ( .A1(\SB1_1_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_20/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_20/buf_output[0] ) );
  BUF_X4 U8937 ( .I(\SB2_1_16/buf_output[4] ), .Z(\RI5[1][100] ) );
  BUF_X4 U8938 ( .I(\SB2_1_16/buf_output[5] ), .Z(\RI5[1][95] ) );
  BUF_X4 U8941 ( .I(\SB2_1_28/buf_output[5] ), .Z(\RI5[1][23] ) );
  BUF_X4 U8942 ( .I(\SB2_1_28/buf_output[4] ), .Z(\RI5[1][28] ) );
  BUF_X4 U8946 ( .I(\SB2_1_30/buf_output[2] ), .Z(\RI5[1][26] ) );
  BUF_X4 U8947 ( .I(\SB2_1_30/buf_output[4] ), .Z(\RI5[1][16] ) );
  BUF_X4 U8949 ( .I(\SB2_1_30/buf_output[5] ), .Z(\RI5[1][11] ) );
  BUF_X4 U8952 ( .I(\SB2_1_27/buf_output[5] ), .Z(\RI5[1][29] ) );
  NAND4_X2 U8954 ( .A1(\SB1_0_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_22/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_22/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_0_22/buf_output[4] ) );
  BUF_X4 U8957 ( .I(\SB2_1_24/buf_output[5] ), .Z(\RI5[1][47] ) );
  BUF_X4 U8958 ( .I(\SB2_1_21/buf_output[0] ), .Z(\RI5[1][90] ) );
  BUF_X4 U8959 ( .I(\SB2_1_21/buf_output[5] ), .Z(\RI5[1][65] ) );
  BUF_X4 U8960 ( .I(\SB2_1_21/buf_output[2] ), .Z(\RI5[1][80] ) );
  BUF_X4 U8961 ( .I(\SB2_1_21/buf_output[4] ), .Z(\RI5[1][70] ) );
  NAND4_X2 U8962 ( .A1(\SB1_1_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_26/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_26/buf_output[0] ) );
  BUF_X4 U8963 ( .I(\SB2_1_26/buf_output[5] ), .Z(\RI5[1][35] ) );
  BUF_X4 U8965 ( .I(\SB2_1_26/buf_output[4] ), .Z(\RI5[1][40] ) );
  BUF_X4 U8966 ( .I(\SB2_1_26/buf_output[1] ), .Z(\RI5[1][55] ) );
  NAND4_X2 U8973 ( .A1(\SB1_2_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_13/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_13/buf_output[1] ) );
  NAND4_X2 U8977 ( .A1(\SB1_2_2/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_2/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_2/buf_output[1] ) );
  NAND4_X2 U8978 ( .A1(\SB1_2_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_8/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_8/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_8/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_2_8/buf_output[4] ) );
  NAND4_X2 U8980 ( .A1(\SB1_2_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_8/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_8/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_8/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_8/buf_output[3] ) );
  NAND4_X2 U8982 ( .A1(\SB1_2_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_18/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_18/buf_output[1] ) );
  NAND4_X2 U8985 ( .A1(\SB1_2_22/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_2_22/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_22/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_2_22/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_2_22/buf_output[5] ) );
  NAND4_X2 U8990 ( .A1(\SB1_2_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_9/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_9/buf_output[0] ) );
  NAND4_X2 U8991 ( .A1(\SB1_2_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_23/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_2_23/buf_output[4] ) );
  NAND4_X2 U8994 ( .A1(\SB1_2_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_30/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_30/buf_output[1] ) );
  NAND4_X2 U8998 ( .A1(\SB1_2_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_19/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_19/buf_output[0] ) );
  NAND4_X2 U9004 ( .A1(\SB1_2_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_21/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_21/buf_output[1] ) );
  NAND4_X2 U9007 ( .A1(\SB1_2_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_4/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_4/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_4/buf_output[2] ) );
  BUF_X4 U9011 ( .I(\SB2_2_5/buf_output[4] ), .Z(\RI5[2][166] ) );
  BUF_X4 U9012 ( .I(\SB2_2_5/buf_output[5] ), .Z(\RI5[2][161] ) );
  BUF_X4 U9013 ( .I(\SB2_2_6/buf_output[4] ), .Z(\RI5[2][160] ) );
  BUF_X4 U9014 ( .I(\SB2_2_6/buf_output[0] ), .Z(\RI5[2][180] ) );
  BUF_X4 U9015 ( .I(\SB2_2_6/buf_output[5] ), .Z(\RI5[2][155] ) );
  BUF_X4 U9019 ( .I(\SB2_2_14/buf_output[5] ), .Z(\RI5[2][107] ) );
  BUF_X4 U9023 ( .I(\SB2_2_15/buf_output[5] ), .Z(\RI5[2][101] ) );
  BUF_X4 U9024 ( .I(\SB2_2_17/buf_output[1] ), .Z(\RI5[2][109] ) );
  BUF_X4 U9027 ( .I(\SB2_2_18/buf_output[5] ), .Z(\RI5[2][83] ) );
  BUF_X4 U9028 ( .I(\SB2_2_18/buf_output[4] ), .Z(\RI5[2][88] ) );
  NAND4_X2 U9029 ( .A1(\SB1_2_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_20/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_2_20/buf_output[4] ) );
  BUF_X4 U9030 ( .I(\SB2_2_16/buf_output[5] ), .Z(\RI5[2][95] ) );
  NAND4_X2 U9031 ( .A1(\SB1_2_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_20/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_20/buf_output[1] ) );
  BUF_X4 U9033 ( .I(\SB2_2_19/buf_output[4] ), .Z(\RI5[2][82] ) );
  BUF_X4 U9034 ( .I(\SB2_2_19/buf_output[5] ), .Z(\RI5[2][77] ) );
  BUF_X4 U9040 ( .I(\SB2_2_24/buf_output[2] ), .Z(\RI5[2][62] ) );
  BUF_X4 U9041 ( .I(\SB2_2_24/buf_output[3] ), .Z(\RI5[2][57] ) );
  BUF_X4 U9044 ( .I(\SB2_2_22/buf_output[5] ), .Z(\RI5[2][59] ) );
  BUF_X4 U9045 ( .I(\SB2_2_29/buf_output[5] ), .Z(\RI5[2][17] ) );
  BUF_X4 U9048 ( .I(\SB2_2_31/buf_output[5] ), .Z(\RI5[2][5] ) );
  BUF_X4 U9050 ( .I(\SB2_1_25/buf_output[5] ), .Z(\RI5[1][41] ) );
  BUF_X4 U9053 ( .I(\SB2_2_7/buf_output[4] ), .Z(\RI5[2][154] ) );
  BUF_X4 U9054 ( .I(\SB2_2_12/buf_output[5] ), .Z(\RI5[2][119] ) );
  BUF_X4 U9055 ( .I(\SB2_2_9/buf_output[5] ), .Z(\RI5[2][137] ) );
  NAND4_X2 U9056 ( .A1(\SB2_2_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_9/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_9/buf_output[3] ) );
  NAND4_X2 U9059 ( .A1(\SB1_3_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_15/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_15/buf_output[1] ) );
  NAND4_X2 U9061 ( .A1(\SB1_3_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_15/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_15/buf_output[0] ) );
  NAND4_X2 U9071 ( .A1(\SB1_3_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_13/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_13/buf_output[1] ) );
  NAND4_X2 U9074 ( .A1(\SB1_3_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_18/buf_output[1] ) );
  NAND4_X2 U9081 ( .A1(\SB1_3_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_1/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_1/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_1/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_1/buf_output[3] ) );
  NAND4_X2 U9083 ( .A1(\SB1_3_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_5/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_5/buf_output[1] ) );
  NAND4_X2 U9087 ( .A1(\SB1_3_16/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_16/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_16/buf_output[0] ) );
  NAND4_X2 U9098 ( .A1(\SB1_3_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_22/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_22/buf_output[0] ) );
  BUF_X4 U9105 ( .I(\SB2_3_3/buf_output[5] ), .Z(\RI5[3][173] ) );
  BUF_X4 U9106 ( .I(\SB2_3_5/buf_output[5] ), .Z(\RI5[3][161] ) );
  NAND4_X2 U9110 ( .A1(\SB1_3_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_8/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_8/buf_output[1] ) );
  BUF_X4 U9113 ( .I(\SB2_3_9/buf_output[5] ), .Z(\RI5[3][137] ) );
  NAND4_X2 U9114 ( .A1(\SB2_3_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_13/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_3_13/buf_output[4] ) );
  BUF_X4 U9116 ( .I(\SB2_3_17/buf_output[0] ), .Z(\RI5[3][114] ) );
  BUF_X4 U9117 ( .I(\SB2_3_17/buf_output[5] ), .Z(\RI5[3][89] ) );
  BUF_X4 U9118 ( .I(\SB2_3_17/buf_output[2] ), .Z(\RI5[3][104] ) );
  BUF_X4 U9120 ( .I(\SB2_3_22/buf_output[5] ), .Z(\RI5[3][59] ) );
  BUF_X4 U9123 ( .I(\SB2_3_21/buf_output[4] ), .Z(\RI5[3][70] ) );
  BUF_X4 U9124 ( .I(\SB2_3_21/buf_output[5] ), .Z(\RI5[3][65] ) );
  NAND4_X2 U9125 ( .A1(\SB1_3_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_25/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_25/buf_output[1] ) );
  BUF_X4 U9127 ( .I(\SB2_3_24/buf_output[5] ), .Z(\RI5[3][47] ) );
  BUF_X4 U9130 ( .I(\SB2_3_28/buf_output[4] ), .Z(\RI5[3][28] ) );
  BUF_X4 U9131 ( .I(\SB2_3_28/buf_output[5] ), .Z(\RI5[3][23] ) );
  BUF_X4 U9133 ( .I(\SB2_3_29/buf_output[4] ), .Z(\RI5[3][22] ) );
  BUF_X4 U9135 ( .I(\SB2_3_27/buf_output[4] ), .Z(\RI5[3][34] ) );
  NAND4_X2 U9137 ( .A1(\SB2_3_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_31/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_31/buf_output[3] ) );
  NAND4_X2 U9139 ( .A1(\SB1_4_2/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_4_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_2/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_4_2/buf_output[0] ) );
  NAND4_X2 U9141 ( .A1(\SB1_4_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_4_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_4_7/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_4_7/buf_output[1] ) );
  NAND4_X2 U9150 ( .A1(\SB1_4_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_4_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_4_31/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_4_31/buf_output[3] ) );
  NAND4_X2 U9153 ( .A1(\SB1_4_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_4_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_4_0/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_4_0/buf_output[1] ) );
  NAND4_X2 U9154 ( .A1(\SB1_4_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_4_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_4_5/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_4_5/buf_output[1] ) );
  NAND4_X2 U9155 ( .A1(\SB1_4_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_4_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_11/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_4_11/buf_output[0] ) );
  NAND4_X2 U9156 ( .A1(\SB1_4_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_4_17/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_4_17/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_4_17/buf_output[4] ) );
  NAND4_X2 U9165 ( .A1(\SB1_4_21/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_4_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_21/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_21/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_4_21/buf_output[0] ) );
  NAND4_X2 U9170 ( .A1(\SB1_4_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_4_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_4_30/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_4_30/buf_output[1] ) );
  BUF_X4 U9171 ( .I(\SB2_3_30/buf_output[5] ), .Z(\RI5[3][11] ) );
  NAND4_X2 U9179 ( .A1(\SB1_4_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_4_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_4_22/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_4_22/buf_output[1] ) );
  NAND4_X2 U9180 ( .A1(\SB1_4_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_4_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_4_26/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_4_26/buf_output[4] ) );
  BUF_X4 U9186 ( .I(\SB2_4_2/buf_output[5] ), .Z(\RI5[4][179] ) );
  BUF_X4 U9187 ( .I(\SB2_4_30/buf_output[2] ), .Z(\RI5[4][26] ) );
  BUF_X4 U9190 ( .I(\SB2_4_30/buf_output[4] ), .Z(\RI5[4][16] ) );
  BUF_X4 U9198 ( .I(\SB2_4_7/buf_output[5] ), .Z(\RI5[4][149] ) );
  BUF_X4 U9201 ( .I(\SB2_4_11/buf_output[0] ), .Z(\RI5[4][150] ) );
  BUF_X4 U9202 ( .I(\SB2_4_11/buf_output[2] ), .Z(\RI5[4][140] ) );
  BUF_X4 U9203 ( .I(\SB2_4_11/buf_output[4] ), .Z(\RI5[4][130] ) );
  BUF_X4 U9206 ( .I(\SB2_4_9/buf_output[4] ), .Z(\RI5[4][142] ) );
  BUF_X4 U9209 ( .I(\SB2_4_10/buf_output[2] ), .Z(\RI5[4][146] ) );
  BUF_X4 U9210 ( .I(\SB2_4_14/buf_output[5] ), .Z(\RI5[4][107] ) );
  NAND4_X2 U9211 ( .A1(\SB2_4_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_4_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_4_14/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_4_14/buf_output[3] ) );
  BUF_X4 U9212 ( .I(\SB2_4_14/buf_output[4] ), .Z(\RI5[4][112] ) );
  BUF_X4 U9214 ( .I(\SB2_4_14/buf_output[2] ), .Z(\RI5[4][122] ) );
  BUF_X4 U9215 ( .I(\SB2_4_13/buf_output[2] ), .Z(\RI5[4][128] ) );
  BUF_X4 U9216 ( .I(\SB2_4_17/buf_output[2] ), .Z(\RI5[4][104] ) );
  BUF_X4 U9217 ( .I(\SB2_4_17/buf_output[0] ), .Z(\RI5[4][114] ) );
  BUF_X4 U9218 ( .I(\SB2_4_17/buf_output[5] ), .Z(\RI5[4][89] ) );
  BUF_X4 U9219 ( .I(\SB2_4_18/buf_output[5] ), .Z(\RI5[4][83] ) );
  BUF_X4 U9221 ( .I(\SB2_4_15/buf_output[5] ), .Z(\RI5[4][101] ) );
  BUF_X4 U9223 ( .I(\SB2_4_16/buf_output[4] ), .Z(\RI5[4][100] ) );
  BUF_X4 U9224 ( .I(\SB2_4_16/buf_output[2] ), .Z(\RI5[4][110] ) );
  BUF_X4 U9225 ( .I(\SB2_4_16/buf_output[5] ), .Z(\RI5[4][95] ) );
  BUF_X4 U9229 ( .I(\SB2_4_19/buf_output[4] ), .Z(\RI5[4][82] ) );
  BUF_X4 U9231 ( .I(\SB2_4_20/buf_output[0] ), .Z(\RI5[4][96] ) );
  BUF_X4 U9232 ( .I(\SB2_4_20/buf_output[5] ), .Z(\RI5[4][71] ) );
  BUF_X4 U9235 ( .I(\SB2_4_21/buf_output[5] ), .Z(\RI5[4][65] ) );
  BUF_X4 U9236 ( .I(\SB2_4_21/buf_output[4] ), .Z(\RI5[4][70] ) );
  NAND4_X2 U9237 ( .A1(\SB2_4_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_4_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_4_23/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_4_23/buf_output[3] ) );
  BUF_X4 U9239 ( .I(\SB2_4_23/buf_output[0] ), .Z(\RI5[4][78] ) );
  BUF_X4 U9240 ( .I(\SB2_4_23/buf_output[4] ), .Z(\RI5[4][58] ) );
  BUF_X4 U9241 ( .I(\SB2_4_26/buf_output[2] ), .Z(\RI5[4][50] ) );
  BUF_X4 U9243 ( .I(\SB2_4_26/buf_output[5] ), .Z(\RI5[4][35] ) );
  BUF_X4 U9247 ( .I(\SB2_4_28/buf_output[4] ), .Z(\RI5[4][28] ) );
  BUF_X4 U9248 ( .I(\SB2_4_28/buf_output[0] ), .Z(\RI5[4][48] ) );
  NAND4_X2 U9249 ( .A1(\SB2_4_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_28/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_4_28/buf_output[1] ) );
  BUF_X4 U9254 ( .I(\SB2_4_25/buf_output[4] ), .Z(\RI5[4][46] ) );
  BUF_X4 U9256 ( .I(\SB2_4_25/buf_output[3] ), .Z(\RI5[4][51] ) );
  BUF_X4 U9257 ( .I(\SB2_4_25/buf_output[5] ), .Z(\RI5[4][41] ) );
  NAND4_X2 U9261 ( .A1(\SB3_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_9/buf_output[4] )
         );
  NAND4_X2 U9263 ( .A1(\SB3_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_3/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_3/buf_output[1] )
         );
  NAND4_X2 U9264 ( .A1(\SB3_8/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_8/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_8/buf_output[0] )
         );
  NAND4_X2 U9266 ( .A1(\SB3_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_8/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_8/Component_Function_3/NAND4_in[3] ), .ZN(\SB3_8/buf_output[3] )
         );
  NAND4_X2 U9268 ( .A1(\SB3_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_29/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_29/buf_output[1] ) );
  BUF_X4 U9269 ( .I(\SB2_4_29/buf_output[5] ), .Z(\RI5[4][17] ) );
  NAND4_X2 U9271 ( .A1(\SB3_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_5/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_5/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_5/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_5/buf_output[4] )
         );
  NAND4_X2 U9278 ( .A1(\SB3_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_6/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_6/buf_output[0] )
         );
  NAND4_X2 U9280 ( .A1(\SB3_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_18/buf_output[1] ) );
  NAND4_X2 U9282 ( .A1(\SB3_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_18/buf_output[4] ) );
  NAND4_X2 U9283 ( .A1(\SB3_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_18/buf_output[0] ) );
  NAND4_X2 U9284 ( .A1(\SB3_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_22/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_22/buf_output[1] ) );
  NAND4_X2 U9286 ( .A1(\SB3_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_22/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_22/buf_output[4] ) );
  NAND4_X2 U9288 ( .A1(\SB3_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_26/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_26/buf_output[4] ) );
  NAND4_X2 U9293 ( .A1(\SB3_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_10/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_10/buf_output[1] ) );
  NAND4_X2 U9294 ( .A1(\SB3_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_16/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_16/buf_output[1] ) );
  NAND4_X2 U9296 ( .A1(\SB3_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_20/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_20/buf_output[0] ) );
  NAND4_X2 U9299 ( .A1(\SB3_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_25/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_25/buf_output[1] ) );
  NAND4_X2 U9301 ( .A1(\SB3_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_2/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_2/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_2/buf_output[4] )
         );
  INV_X2 \SB1_2_22/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[57] ), .ZN(
        \SB1_2_22/i0[8] ) );
  NAND3_X2 \SB1_1_30/Component_Function_5/N2  ( .A1(\SB1_1_30/i0_0 ), .A2(
        \SB1_1_30/i0[6] ), .A3(\SB1_1_30/i0[10] ), .ZN(
        \SB1_1_30/Component_Function_5/NAND4_in[1] ) );
  AND2_X1 U1838 ( .A1(\SB1_4_27/buf_output[3] ), .A2(\SB1_4_28/buf_output[2] ), 
        .Z(n1026) );
  NAND2_X2 \SB1_1_7/Component_Function_5/N1  ( .A1(\SB1_1_7/i0_0 ), .A2(
        \SB1_1_7/i3[0] ), .ZN(\SB1_1_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U1740 ( .A1(\SB2_2_9/i0_0 ), .A2(\SB2_2_9/i0_4 ), .A3(
        \SB2_2_9/i1_5 ), .ZN(n2844) );
  INV_X4 U8110 ( .I(n2748), .ZN(\SB1_2_2/buf_output[4] ) );
  NAND3_X2 \SB3_30/Component_Function_2/N1  ( .A1(\SB3_30/i1_5 ), .A2(
        \SB3_30/i0[10] ), .A3(\SB3_30/i1[9] ), .ZN(
        \SB3_30/Component_Function_2/NAND4_in[0] ) );
  BUF_X2 U2045 ( .I(\SB1_1_14/buf_output[4] ), .Z(n2156) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_34  ( .I(\SB2_1_27/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[34] ) );
  NAND3_X2 \SB2_1_6/Component_Function_5/N2  ( .A1(\SB2_1_6/i0_0 ), .A2(
        \SB2_1_6/i0[6] ), .A3(\SB2_1_6/i0[10] ), .ZN(
        \SB2_1_6/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB2_1_28/INV_5  ( .I(\SB1_1_28/buf_output[5] ), .ZN(\SB2_1_28/i1_5 )
         );
  NAND3_X2 U5461 ( .A1(\SB2_3_26/i0[9] ), .A2(\SB2_3_26/i0_4 ), .A3(
        \SB2_3_26/i0[6] ), .ZN(\SB2_3_26/Component_Function_5/NAND4_in[3] ) );
  BUF_X2 \SB3_10/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[126] ), .Z(
        \SB3_10/i0[9] ) );
  INV_X2 U2356 ( .I(\RI1[4][65] ), .ZN(\SB1_4_21/i1_5 ) );
  NAND3_X2 U1148 ( .A1(\SB1_1_17/i0_3 ), .A2(\SB1_1_17/i0_4 ), .A3(
        \SB1_1_17/i1[9] ), .ZN(n1187) );
  NAND3_X2 U588 ( .A1(\SB3_29/i0_4 ), .A2(\SB3_29/i0[6] ), .A3(\SB3_29/i0[9] ), 
        .ZN(\SB3_29/Component_Function_5/NAND4_in[3] ) );
  INV_X2 \SB1_2_22/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[56] ), .ZN(
        \SB1_2_22/i1[9] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_144  ( .I(\SB2_3_12/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[144] ) );
  INV_X2 \SB2_4_21/INV_5  ( .I(\SB1_4_21/buf_output[5] ), .ZN(\SB2_4_21/i1_5 )
         );
  NAND3_X2 \SB2_2_19/Component_Function_5/N4  ( .A1(\SB2_2_19/i0[9] ), .A2(
        \SB2_2_19/i0[6] ), .A3(\SB2_2_19/i0_4 ), .ZN(
        \SB2_2_19/Component_Function_5/NAND4_in[3] ) );
  INV_X2 \SB2_3_9/INV_5  ( .I(\SB1_3_9/buf_output[5] ), .ZN(\SB2_3_9/i1_5 ) );
  INV_X2 \SB2_4_2/INV_5  ( .I(\SB1_4_2/buf_output[5] ), .ZN(\SB2_4_2/i1_5 ) );
  INV_X2 \SB1_0_29/INV_3  ( .I(n321), .ZN(\SB1_0_29/i0[8] ) );
  NAND3_X2 \SB2_1_28/Component_Function_5/N2  ( .A1(\SB2_1_28/i0_0 ), .A2(
        \SB2_1_28/i0[6] ), .A3(\SB2_1_28/i0[10] ), .ZN(
        \SB2_1_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X2 \SB1_0_17/Component_Function_5/N1  ( .A1(\SB1_0_17/i0_0 ), .A2(
        \SB1_0_17/i3[0] ), .ZN(\SB1_0_17/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U1860 ( .I(\SB1_3_3/buf_output[5] ), .Z(\SB2_3_3/i0_3 ) );
  INV_X2 \SB2_1_31/INV_4  ( .I(n5429), .ZN(\SB2_1_31/i0[7] ) );
  NAND3_X2 U922 ( .A1(\SB2_2_7/i0[10] ), .A2(\SB2_2_7/i0_0 ), .A3(
        \SB2_2_7/i0[6] ), .ZN(\SB2_2_7/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB1_3_2/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[179] ), .ZN(
        \SB1_3_2/i1_5 ) );
  INV_X2 U4398 ( .I(\SB1_2_4/buf_output[5] ), .ZN(\SB2_2_4/i1_5 ) );
  NAND3_X2 \SB2_3_27/Component_Function_4/N4  ( .A1(\SB2_3_27/i1[9] ), .A2(
        \SB2_3_27/i1_5 ), .A3(\SB2_3_27/i0_4 ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 U2016 ( .I(\SB2_2_4/buf_output[0] ), .Z(\RI5[2][0] ) );
  NAND4_X2 U4695 ( .A1(\SB2_2_4/Component_Function_0/NAND4_in[1] ), .A2(n1600), 
        .A3(\SB2_2_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_4/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_4/buf_output[0] ) );
  NAND3_X2 \SB1_2_28/Component_Function_2/N2  ( .A1(\SB1_2_28/i0_3 ), .A2(
        \SB1_2_28/i0[10] ), .A3(\SB1_2_28/i0[6] ), .ZN(
        \SB1_2_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U1086 ( .A1(\SB2_1_31/i0[6] ), .A2(\SB2_1_31/i0[9] ), .A3(n5430), 
        .ZN(n1759) );
  NAND3_X2 \SB2_1_8/Component_Function_3/N3  ( .A1(\SB2_1_8/i1[9] ), .A2(
        \SB2_1_8/i1_7 ), .A3(\SB2_1_8/i0[10] ), .ZN(
        \SB2_1_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_23/Component_Function_3/N1  ( .A1(\SB2_0_23/i1[9] ), .A2(
        \SB2_0_23/i0_3 ), .A3(\SB2_0_23/i0[6] ), .ZN(
        \SB2_0_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U818 ( .A1(\SB2_3_3/i0[10] ), .A2(\SB2_3_3/i0_0 ), .A3(
        \SB2_3_3/i0[6] ), .ZN(\SB2_3_3/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U3111 ( .A1(\SB2_1_31/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_31/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_31/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_31/buf_output[0] ) );
  NAND3_X2 U820 ( .A1(\SB2_3_3/i0_3 ), .A2(\SB2_3_3/i0_4 ), .A3(
        \SB2_3_3/i1[9] ), .ZN(n916) );
  BUF_X4 \SB2_3_8/BUF_3_0  ( .I(\SB2_3_8/buf_output[3] ), .Z(\RI5[3][153] ) );
  NAND3_X2 U956 ( .A1(\SB2_2_7/i0[10] ), .A2(\SB2_2_7/i0_3 ), .A3(
        \SB2_2_7/i0[9] ), .ZN(\SB2_2_7/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_15/Component_Function_2/N3  ( .A1(\SB2_3_15/i0_3 ), .A2(
        \SB2_3_15/i0[8] ), .A3(\SB2_3_15/i0[9] ), .ZN(
        \SB2_3_15/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB1_2_15/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[98] ), .ZN(
        \SB1_2_15/i1[9] ) );
  INV_X2 \SB2_2_2/INV_5  ( .I(\SB1_2_2/buf_output[5] ), .ZN(\SB2_2_2/i1_5 ) );
  NAND4_X2 U6316 ( .A1(\SB2_3_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_4/Component_Function_2/NAND4_in[2] ), .A4(n1875), .ZN(
        \SB2_3_4/buf_output[2] ) );
  INV_X2 U2588 ( .I(\SB1_2_12/buf_output[5] ), .ZN(\SB2_2_12/i1_5 ) );
  NAND4_X2 U4600 ( .A1(\SB2_1_10/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_1_10/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_10/Component_Function_1/NAND4_in[0] ), .A4(n1359), .ZN(
        \SB2_1_10/buf_output[1] ) );
  BUF_X4 U644 ( .I(\SB2_4_8/buf_output[1] ), .Z(\RI5[4][163] ) );
  BUF_X4 U1859 ( .I(\RI5[3][123] ), .Z(n575) );
  NAND3_X2 U1080 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i0[6] ), .A3(
        \SB2_1_20/i0_3 ), .ZN(\SB2_1_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_3_16/Component_Function_2/N2  ( .A1(\SB2_3_16/i0_3 ), .A2(
        \SB2_3_16/i0[10] ), .A3(\SB2_3_16/i0[6] ), .ZN(
        \SB2_3_16/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U1823 ( .I(\SB1_1_9/buf_output[5] ), .ZN(\SB2_1_9/i1_5 ) );
  NAND3_X2 U4789 ( .A1(\SB2_0_23/i0[6] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i0[10] ), .ZN(\SB2_0_23/Component_Function_2/NAND4_in[1] )
         );
  INV_X2 U1711 ( .I(\MC_ARK_ARC_1_0/buf_output[32] ), .ZN(\SB1_1_26/i1[9] ) );
  BUF_X4 \SB2_3_26/BUF_4_0  ( .I(\SB2_3_26/buf_output[4] ), .Z(\RI5[3][40] )
         );
  INV_X2 \SB2_4_25/INV_5  ( .I(\SB1_4_25/buf_output[5] ), .ZN(\SB2_4_25/i1_5 )
         );
  BUF_X4 \SB2_2_2/BUF_2_0  ( .I(\SB2_2_2/buf_output[2] ), .Z(\RI5[2][2] ) );
  NAND3_X2 U668 ( .A1(\SB2_4_2/i0[10] ), .A2(\SB2_4_2/i1[9] ), .A3(
        \SB2_4_2/i1_7 ), .ZN(\SB2_4_2/Component_Function_3/NAND4_in[2] ) );
  INV_X2 U5333 ( .I(\SB1_4_24/buf_output[3] ), .ZN(\SB2_4_22/i0[8] ) );
  BUF_X2 \SB2_4_15/BUF_0  ( .I(\SB1_4_20/buf_output[0] ), .Z(\SB2_4_15/i0[9] )
         );
  BUF_X2 U5128 ( .I(\SB3_22/buf_output[3] ), .Z(\SB4_20/i0[10] ) );
  INV_X2 U1871 ( .I(\SB1_2_22/buf_output[5] ), .ZN(\SB2_2_22/i1_5 ) );
  NAND3_X2 U898 ( .A1(\SB1_3_2/i0_3 ), .A2(\SB1_3_2/i0[8] ), .A3(
        \SB1_3_2/i0[9] ), .ZN(\SB1_3_2/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U1870 ( .I(\SB1_2_22/buf_output[5] ), .Z(\SB2_2_22/i0_3 ) );
  INV_X2 U1514 ( .I(\MC_ARK_ARC_1_2/buf_output[177] ), .ZN(\SB1_3_2/i0[8] ) );
  NAND3_X2 \SB1_3_14/Component_Function_5/N3  ( .A1(\SB1_3_14/i1[9] ), .A2(
        \SB1_3_14/i0_4 ), .A3(\RI1[3][107] ), .ZN(
        \SB1_3_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U7345 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0[10] ), .A3(
        \SB2_2_24/i0[6] ), .ZN(\SB2_2_24/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U6729 ( .I(\SB1_1_7/buf_output[5] ), .ZN(\SB2_1_7/i1_5 ) );
  NAND3_X2 \SB2_3_15/Component_Function_1/N2  ( .A1(\SB2_3_15/i0_3 ), .A2(
        \SB2_3_15/i1_7 ), .A3(\SB2_3_15/i0[8] ), .ZN(
        \SB2_3_15/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \SB2_1_7/BUF_4_0  ( .I(\SB2_1_7/buf_output[4] ), .Z(\RI5[1][154] ) );
  NAND4_X2 U4601 ( .A1(\SB2_1_7/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_7/Component_Function_4/NAND4_in[1] ), .A3(n1360), .A4(
        \SB2_1_7/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_1_7/buf_output[4] ) );
  NAND4_X2 \SB2_3_21/Component_Function_1/N5  ( .A1(
        \SB2_3_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_21/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_21/buf_output[1] ) );
  NAND3_X2 \SB2_2_23/Component_Function_2/N3  ( .A1(\SB2_2_23/i0_3 ), .A2(
        \SB2_2_23/i0[8] ), .A3(\SB2_2_23/i0[9] ), .ZN(
        \SB2_2_23/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB2_0_27/BUF_0_0  ( .I(\SB2_0_27/buf_output[0] ), .Z(\RI5[0][54] )
         );
  NAND2_X2 \SB2_1_20/Component_Function_5/N1  ( .A1(\SB2_1_20/i0_0 ), .A2(
        \SB2_1_20/i3[0] ), .ZN(\SB2_1_20/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U9253 ( .I(\SB2_4_24/buf_output[0] ), .Z(\RI5[4][72] ) );
  NAND3_X2 \SB2_1_25/Component_Function_1/N4  ( .A1(\SB2_1_25/i1_7 ), .A2(
        n3995), .A3(\SB2_1_25/i0_4 ), .ZN(
        \SB2_1_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U976 ( .A1(\SB1_2_27/i1[9] ), .A2(\SB1_2_27/i0_4 ), .A3(
        \SB1_2_27/i0_3 ), .ZN(n2151) );
  BUF_X4 U961 ( .I(\SB1_2_8/buf_output[4] ), .Z(\SB2_2_7/i0_4 ) );
  NAND2_X2 U1089 ( .A1(\SB2_1_4/i0_0 ), .A2(\SB2_1_4/i3[0] ), .ZN(n2104) );
  INV_X2 \SB1_1_22/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[56] ), .ZN(
        \SB1_1_22/i1[9] ) );
  CLKBUF_X4 \SB2_0_15/BUF_3  ( .I(\RI3[0][99] ), .Z(\SB2_0_15/i0[10] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_188  ( .I(\SB2_1_3/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[188] ) );
  NAND4_X2 U8268 ( .A1(\SB2_1_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_3/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_3/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_1_3/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_1_3/buf_output[2] ) );
  BUF_X4 U9252 ( .I(\SB2_4_24/buf_output[2] ), .Z(\RI5[4][62] ) );
  NAND3_X2 \SB2_2_0/Component_Function_2/N2  ( .A1(\SB2_2_0/i0_3 ), .A2(
        \SB2_2_0/i0[10] ), .A3(\SB2_2_0/i0[6] ), .ZN(
        \SB2_2_0/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U1375 ( .I(\MC_ARK_ARC_1_2/buf_output[117] ), .ZN(\SB1_3_12/i0[8] )
         );
  NAND3_X2 \SB1_2_4/Component_Function_1/N4  ( .A1(\SB1_2_4/i1_7 ), .A2(
        \SB1_2_4/i0[8] ), .A3(\SB1_2_4/i0_4 ), .ZN(
        \SB1_2_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U1800 ( .A1(\SB2_4_26/i1[9] ), .A2(\SB2_4_26/i0_3 ), .A3(
        \SB2_4_26/i0[6] ), .ZN(\SB2_4_26/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_0_6/BUF_1_0  ( .I(\SB2_0_6/buf_output[1] ), .Z(\RI5[0][175] ) );
  NAND3_X2 \SB2_2_23/Component_Function_3/N2  ( .A1(\SB2_2_23/i0_0 ), .A2(
        \SB2_2_23/i0_3 ), .A3(n600), .ZN(
        \SB2_2_23/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB2_0_23/BUF_1  ( .I(\RI3[0][49] ), .Z(\SB2_0_23/i0[6] ) );
  BUF_X2 U1097 ( .I(\SB1_1_12/buf_output[1] ), .Z(\SB2_1_8/i0[6] ) );
  NAND3_X2 U4696 ( .A1(\SB2_2_2/i0_3 ), .A2(\SB2_2_2/i0[9] ), .A3(
        \SB2_2_2/i0[8] ), .ZN(\SB2_2_2/Component_Function_2/NAND4_in[2] ) );
  AND4_X2 U236 ( .A1(\SB3_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_11/Component_Function_3/NAND4_in[3] ), .Z(n1499) );
  NAND3_X2 \SB1_3_25/Component_Function_2/N2  ( .A1(\SB1_3_25/i0_3 ), .A2(
        \SB1_3_25/i0[10] ), .A3(\SB1_3_25/i0[6] ), .ZN(
        \SB1_3_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB1_3_7/Component_Function_2/N2  ( .A1(\SB1_3_7/i0_3 ), .A2(
        \SB1_3_7/i0[10] ), .A3(\SB1_3_7/i0[6] ), .ZN(
        \SB1_3_7/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U1912 ( .I(\MC_ARK_ARC_1_2/buf_output[131] ), .Z(\SB1_3_10/i0_3 ) );
  INV_X2 U1499 ( .I(\MC_ARK_ARC_1_3/buf_output[170] ), .ZN(\SB1_4_3/i1[9] ) );
  BUF_X4 \SB1_3_7/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[148] ), .Z(
        \SB1_3_7/i0_4 ) );
  NAND3_X2 U667 ( .A1(\SB2_4_1/i0[10] ), .A2(\SB2_4_1/i0_0 ), .A3(
        \SB2_4_1/i0[6] ), .ZN(\SB2_4_1/Component_Function_5/NAND4_in[1] ) );
  NAND2_X2 U2091 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i1[9] ), .ZN(
        \SB1_0_20/Component_Function_1/NAND4_in[0] ) );
  NAND4_X2 \SB2_1_12/Component_Function_1/N5  ( .A1(
        \SB2_1_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_12/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_1_12/buf_output[1] ) );
  INV_X2 \SB1_0_18/INV_2  ( .I(n1507), .ZN(\SB1_0_18/i1[9] ) );
  NAND3_X2 \SB2_0_16/Component_Function_5/N2  ( .A1(\SB2_0_16/i0_0 ), .A2(
        \SB2_0_16/i0[6] ), .A3(\RI3[0][93] ), .ZN(
        \SB2_0_16/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_0_2/BUF_4_0  ( .I(\SB2_0_2/buf_output[4] ), .Z(\RI5[0][184] ) );
  NAND3_X2 U1092 ( .A1(\SB2_1_31/i0_0 ), .A2(\SB2_1_31/i0[10] ), .A3(
        \SB2_1_31/i0[6] ), .ZN(n2501) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_187  ( .I(\SB2_3_4/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[187] ) );
  NAND4_X2 \SB2_3_4/Component_Function_1/N5  ( .A1(
        \SB2_3_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_4/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_3_4/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_4/buf_output[1] ) );
  NAND3_X2 \SB2_3_16/Component_Function_1/N4  ( .A1(\SB2_3_16/i1_7 ), .A2(
        \SB2_3_16/i0[8] ), .A3(\SB2_3_16/i0_4 ), .ZN(
        \SB2_3_16/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 \SB2_0_16/BUF_1_0  ( .I(\SB2_0_16/buf_output[1] ), .Z(\RI5[0][115] )
         );
  AND4_X2 U959 ( .A1(\SB1_2_10/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_2_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_10/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_2_10/Component_Function_5/NAND4_in[2] ), .Z(n589) );
  NAND2_X2 \SB2_3_3/Component_Function_5/N1  ( .A1(\SB2_3_3/i0_0 ), .A2(
        \SB2_3_3/i3[0] ), .ZN(\SB2_3_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_21/Component_Function_2/N2  ( .A1(\SB2_1_21/i0_3 ), .A2(
        \SB2_1_21/i0[10] ), .A3(\SB2_1_21/i0[6] ), .ZN(
        \SB2_1_21/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U1585 ( .I(\MC_ARK_ARC_1_2/buf_output[45] ), .ZN(\SB1_3_24/i0[8] ) );
  NAND3_X2 U2207 ( .A1(\SB2_1_27/i0_3 ), .A2(\SB2_1_27/i0[9] ), .A3(
        \SB2_1_27/i0[10] ), .ZN(\SB2_1_27/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X2 \SB2_1_19/Component_Function_3/N2  ( .A1(\SB2_1_19/i0_0 ), .A2(
        \SB2_1_19/i0_3 ), .A3(\SB2_1_19/i0_4 ), .ZN(
        \SB2_1_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_3_16/Component_Function_3/N3  ( .A1(\SB2_3_16/i1[9] ), .A2(
        \SB2_3_16/i1_7 ), .A3(\SB2_3_16/i0[10] ), .ZN(
        \SB2_3_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U1517 ( .A1(\SB1_0_21/i0[10] ), .A2(\SB1_0_21/i0_0 ), .A3(
        \SB1_0_21/i0[6] ), .ZN(\SB1_0_21/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U2331 ( .A1(\SB2_3_27/i1_5 ), .A2(\SB2_3_27/i0_0 ), .A3(
        \SB2_3_27/i0_4 ), .ZN(\SB2_3_27/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U886 ( .A1(\SB1_3_31/i0[10] ), .A2(\SB1_3_31/i0_0 ), .A3(
        \SB1_3_31/i0[6] ), .ZN(\SB1_3_31/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U7485 ( .I(\SB2_3_21/buf_output[0] ), .Z(\RI5[3][90] ) );
  NAND3_X2 \SB1_0_12/Component_Function_5/N2  ( .A1(\SB1_0_12/i0_0 ), .A2(
        \SB1_0_12/i0[6] ), .A3(\SB1_0_12/i0[10] ), .ZN(
        \SB1_0_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_20/Component_Function_2/N2  ( .A1(\SB1_0_20/i0_3 ), .A2(
        \SB1_0_20/i0[10] ), .A3(\SB1_0_20/i0[6] ), .ZN(
        \SB1_0_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_3_15/Component_Function_3/N4  ( .A1(\SB2_3_15/i1_5 ), .A2(
        \SB2_3_15/i0[8] ), .A3(\SB2_3_15/i3[0] ), .ZN(
        \SB2_3_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U660 ( .A1(\SB2_4_24/i0_4 ), .A2(\SB2_4_24/i0_3 ), .A3(
        \SB2_4_24/i0_0 ), .ZN(\SB2_4_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U2409 ( .A1(\SB2_4_4/i0[10] ), .A2(\SB2_4_4/i1[9] ), .A3(
        \SB2_4_4/i1_7 ), .ZN(\SB2_4_4/Component_Function_3/NAND4_in[2] ) );
  BUF_X2 U1597 ( .I(\SB3_7/buf_output[3] ), .Z(\SB4_5/i0[10] ) );
  NAND3_X2 U1674 ( .A1(\SB2_3_7/i0[7] ), .A2(\SB2_3_7/i0_3 ), .A3(
        \SB2_3_7/i0_0 ), .ZN(\SB2_3_7/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 U5469 ( .I(\MC_ARK_ARC_1_1/buf_output[120] ), .Z(\SB1_2_11/i0[9] )
         );
  BUF_X4 U5196 ( .I(\SB1_2_10/buf_output[2] ), .Z(\SB2_2_7/i0_0 ) );
  BUF_X4 U2056 ( .I(\SB2_0_18/buf_output[3] ), .Z(\RI5[0][93] ) );
  NAND2_X2 \SB2_2_0/Component_Function_1/N1  ( .A1(\SB2_2_0/i0_3 ), .A2(
        \SB2_2_0/i1[9] ), .ZN(\SB2_2_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_7/Component_Function_2/N2  ( .A1(\SB1_1_7/i0_3 ), .A2(
        \SB1_1_7/i0[10] ), .A3(\SB1_1_7/i0[6] ), .ZN(
        \SB1_1_7/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB1_2_10/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[130] ), .Z(
        \SB1_2_10/i0_4 ) );
  NAND3_X2 \SB1_3_25/Component_Function_3/N2  ( .A1(\SB1_3_25/i0_0 ), .A2(
        \SB1_3_25/i0_3 ), .A3(\SB1_3_25/i0_4 ), .ZN(
        \SB1_3_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U2402 ( .A1(\SB2_4_3/i0_0 ), .A2(\SB2_4_3/i0_3 ), .A3(
        \SB2_4_3/i0_4 ), .ZN(\SB2_4_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U658 ( .A1(\SB2_4_3/i0_0 ), .A2(n3988), .A3(\SB2_4_3/i0_4 ), .ZN(
        \SB2_4_3/Component_Function_2/NAND4_in[3] ) );
  INV_X2 \SB2_4_4/INV_5  ( .I(\SB1_4_4/buf_output[5] ), .ZN(\SB2_4_4/i1_5 ) );
  NAND2_X2 \SB2_1_29/Component_Function_5/N1  ( .A1(\SB2_1_29/i0_0 ), .A2(
        \SB2_1_29/i3[0] ), .ZN(\SB2_1_29/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 \SB2_0_6/Component_Function_2/N5  ( .A1(
        \SB2_0_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_6/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_6/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_6/buf_output[2] ) );
  NAND3_X2 \SB1_1_12/Component_Function_2/N1  ( .A1(\SB1_1_12/i1_5 ), .A2(
        \SB1_1_12/i0[10] ), .A3(\SB1_1_12/i1[9] ), .ZN(
        \SB1_1_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_4/Component_Function_2/N3  ( .A1(\SB2_1_4/i0_3 ), .A2(
        \SB2_1_4/i0[8] ), .A3(\SB2_1_4/i0[9] ), .ZN(
        \SB2_1_4/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 \SB1_0_11/Component_Function_1/N5  ( .A1(
        \SB1_0_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_11/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_11/buf_output[1] ) );
  NAND3_X2 \SB2_2_16/Component_Function_3/N3  ( .A1(\SB2_2_16/i1[9] ), .A2(
        \SB2_2_16/i1_7 ), .A3(\SB2_2_16/i0[10] ), .ZN(
        \SB2_2_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U1100 ( .A1(\SB1_1_15/i0[10] ), .A2(\SB1_1_15/i0[9] ), .A3(
        \SB1_1_15/i0_3 ), .ZN(\SB1_1_15/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 U1866 ( .I(\MC_ARK_ARC_1_1/buf_datainput[172] ), .Z(n578) );
  INV_X2 U1732 ( .I(\MC_ARK_ARC_1_3/buf_output[164] ), .ZN(\SB1_4_4/i1[9] ) );
  BUF_X4 U1168 ( .I(\MC_ARK_ARC_1_0/buf_output[124] ), .Z(\SB1_1_11/i0_4 ) );
  BUF_X4 U7393 ( .I(\SB2_3_15/buf_output[1] ), .Z(\RI5[3][121] ) );
  NAND2_X2 \SB2_1_5/Component_Function_1/N1  ( .A1(\SB2_1_5/i0_3 ), .A2(
        \SB2_1_5/i1[9] ), .ZN(\SB2_1_5/Component_Function_1/NAND4_in[0] ) );
  INV_X2 U2449 ( .I(\RI1[5][77] ), .ZN(\SB3_19/i1_5 ) );
  BUF_X4 U1854 ( .I(\MC_ARK_ARC_1_0/buf_output[99] ), .Z(\SB1_1_15/i0[10] ) );
  INV_X2 U1862 ( .I(\MC_ARK_ARC_1_3/buf_output[159] ), .ZN(\SB1_4_5/i0[8] ) );
  INV_X2 \SB1_1_12/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[119] ), .ZN(
        \SB1_1_12/i1_5 ) );
  INV_X2 U5123 ( .I(\MC_ARK_ARC_1_2/buf_output[23] ), .ZN(\SB1_3_28/i1_5 ) );
  NAND3_X2 U1041 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0[10] ), .A3(
        \SB2_1_10/i0_4 ), .ZN(n775) );
  CLKBUF_X4 \SB1_1_21/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[61] ), .Z(
        \SB1_1_21/i0[6] ) );
  BUF_X4 U5122 ( .I(\MC_ARK_ARC_1_2/buf_output[23] ), .Z(\SB1_3_28/i0_3 ) );
  NAND3_X2 \SB2_3_16/Component_Function_1/N2  ( .A1(\SB2_3_16/i0_3 ), .A2(
        \SB2_3_16/i1_7 ), .A3(\SB2_3_16/i0[8] ), .ZN(
        \SB2_3_16/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U2022 ( .I(\SB1_2_0/buf_output[5] ), .Z(\SB2_2_0/i0_3 ) );
  NAND2_X2 U741 ( .A1(\SB1_4_22/i0_0 ), .A2(\SB1_4_22/i3[0] ), .ZN(n1091) );
  NAND3_X2 \SB2_1_13/Component_Function_1/N4  ( .A1(\SB2_1_13/i1_7 ), .A2(
        \SB2_1_13/i0[8] ), .A3(\SB2_1_13/i0_4 ), .ZN(
        \SB2_1_13/Component_Function_1/NAND4_in[3] ) );
  INV_X2 \SB1_3_13/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[109] ), .ZN(
        \SB1_3_13/i1_7 ) );
  NAND3_X2 \SB1_1_12/Component_Function_1/N2  ( .A1(\SB1_1_12/i0_3 ), .A2(
        \SB1_1_12/i1_7 ), .A3(\SB1_1_12/i0[8] ), .ZN(
        \SB1_1_12/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \SB2_2_14/BUF_4  ( .I(\SB1_2_15/buf_output[4] ), .Z(\SB2_2_14/i0_4 )
         );
  NAND3_X2 U5431 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0[8] ), .A3(
        \SB1_0_2/i0[9] ), .ZN(\SB1_0_2/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB1_3_1/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[185] ), .ZN(
        \SB1_3_1/i1_5 ) );
  INV_X2 \SB2_0_30/INV_1  ( .I(\SB1_0_2/buf_output[1] ), .ZN(\SB2_0_30/i1_7 )
         );
  NAND3_X2 \SB2_2_21/Component_Function_5/N2  ( .A1(\SB2_2_21/i0_0 ), .A2(
        \SB2_2_21/i0[6] ), .A3(\SB2_2_21/i0[10] ), .ZN(
        \SB2_2_21/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB1_1_29/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[17] ), .Z(
        \SB1_1_29/i0_3 ) );
  NAND3_X2 U1608 ( .A1(\SB1_0_0/i0[10] ), .A2(\SB1_0_0/i1[9] ), .A3(
        \SB1_0_0/i1_7 ), .ZN(n1169) );
  NAND3_X2 U888 ( .A1(\SB1_3_4/i0_4 ), .A2(\SB1_3_4/i1[9] ), .A3(\RI1[3][167] ), .ZN(n643) );
  NAND4_X2 U9196 ( .A1(\SB2_4_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_7/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_4_7/buf_output[1] ) );
  BUF_X4 U9220 ( .I(\SB2_4_15/buf_output[0] ), .Z(\RI5[4][126] ) );
  NAND4_X2 U7133 ( .A1(\SB2_4_15/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_15/Component_Function_0/NAND4_in[2] ), .A3(n2258), .A4(
        \SB2_4_15/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_4_15/buf_output[0] ) );
  BUF_X2 U5053 ( .I(\SB3_4/buf_output[3] ), .Z(\SB4_2/i0[10] ) );
  NAND3_X2 U1610 ( .A1(\SB1_0_0/i0[10] ), .A2(\SB1_0_0/i0_3 ), .A3(
        \SB1_0_0/i0[6] ), .ZN(n1552) );
  INV_X2 U1885 ( .I(\RI1[4][105] ), .ZN(\SB1_4_14/i0[8] ) );
  INV_X2 \SB1_1_8/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[143] ), .ZN(
        \SB1_1_8/i1_5 ) );
  NAND3_X2 U610 ( .A1(\SB3_17/i0[8] ), .A2(\SB3_17/i1_5 ), .A3(\SB3_17/i3[0] ), 
        .ZN(n3020) );
  NAND3_X2 U1095 ( .A1(\SB2_1_4/i0_0 ), .A2(\SB2_1_4/i0[8] ), .A3(
        \SB2_1_4/i0[9] ), .ZN(\SB2_1_4/Component_Function_4/NAND4_in[0] ) );
  BUF_X4 U3648 ( .I(\SB2_3_9/buf_output[0] ), .Z(\RI5[3][162] ) );
  NAND2_X2 \SB1_1_10/Component_Function_5/N1  ( .A1(\SB1_1_10/i0_0 ), .A2(
        \SB1_1_10/i3[0] ), .ZN(\SB1_1_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_8/Component_Function_0/N4  ( .A1(\SB2_1_8/i0[7] ), .A2(
        \SB2_1_8/i0_3 ), .A3(\SB2_1_8/i0_0 ), .ZN(
        \SB2_1_8/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 U5434 ( .I(\SB1_2_12/buf_output[5] ), .Z(\SB2_2_12/i0_3 ) );
  BUF_X4 \SB1_3_28/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[22] ), .Z(
        \SB1_3_28/i0_4 ) );
  NAND4_X2 \SB2_0_4/Component_Function_1/N5  ( .A1(
        \SB2_0_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_4/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_4/buf_output[1] ) );
  NAND3_X2 U816 ( .A1(\SB2_3_2/i0[9] ), .A2(\SB2_3_2/i0_3 ), .A3(
        \SB2_3_2/i0[8] ), .ZN(n1092) );
  NAND3_X2 \SB1_0_6/Component_Function_2/N3  ( .A1(\SB1_0_6/i0_3 ), .A2(
        \SB1_0_6/i0[8] ), .A3(\SB1_0_6/i0[9] ), .ZN(
        \SB1_0_6/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U70 ( .I(Key[30]), .Z(n30) );
  NAND2_X2 \SB1_1_29/Component_Function_5/N1  ( .A1(\SB1_1_29/i0_0 ), .A2(
        \SB1_1_29/i3[0] ), .ZN(\SB1_1_29/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_0_6/BUF_2_0  ( .I(\SB2_0_6/buf_output[2] ), .Z(\RI5[0][170] ) );
  NAND2_X2 \SB1_4_9/Component_Function_5/N1  ( .A1(\SB1_4_9/i0_0 ), .A2(
        \SB1_4_9/i3[0] ), .ZN(\SB1_4_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U953 ( .A1(\SB2_2_27/i3[0] ), .A2(\SB2_2_27/i0[8] ), .A3(
        \SB2_2_27/i1_5 ), .ZN(n1923) );
  NAND2_X2 \SB2_0_31/Component_Function_5/N1  ( .A1(\SB2_0_31/i0_0 ), .A2(
        n5450), .ZN(\SB2_0_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_4_0/Component_Function_5/N4  ( .A1(\SB1_4_0/i0[9] ), .A2(
        \SB1_4_0/i0[6] ), .A3(\SB1_4_0/i0_4 ), .ZN(
        \SB1_4_0/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \SB2_3_9/BUF_1  ( .I(\SB1_3_13/buf_output[1] ), .Z(\SB2_3_9/i0[6] )
         );
  BUF_X2 \SB1_1_6/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[151] ), .Z(
        \SB1_1_6/i0[6] ) );
  NAND3_X2 U1145 ( .A1(\SB1_1_14/i0[10] ), .A2(\SB1_1_14/i1[9] ), .A3(
        \SB1_1_14/i1_7 ), .ZN(\SB1_1_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_6/Component_Function_3/N4  ( .A1(\SB2_0_6/i1_5 ), .A2(
        \SB2_0_6/i0[8] ), .A3(\SB2_0_6/i3[0] ), .ZN(
        \SB2_0_6/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_0_9/BUF_0_0  ( .I(\SB2_0_9/buf_output[0] ), .Z(\RI5[0][162] ) );
  NAND2_X2 \SB4_16/Component_Function_0/N1  ( .A1(\SB4_16/i0[10] ), .A2(
        \SB4_16/i0[9] ), .ZN(\SB4_16/Component_Function_0/NAND4_in[0] ) );
  BUF_X4 \SB1_3_30/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[11] ), .Z(
        \SB1_3_30/i0_3 ) );
  BUF_X4 U7599 ( .I(\SB2_3_1/buf_output[1] ), .Z(\RI5[3][13] ) );
  NAND3_X2 \SB1_3_28/Component_Function_1/N4  ( .A1(\SB1_3_28/i1_7 ), .A2(
        \SB1_3_28/i0[8] ), .A3(\SB1_3_28/i0_4 ), .ZN(
        \SB1_3_28/Component_Function_1/NAND4_in[3] ) );
  INV_X2 \SB1_0_25/INV_2  ( .I(n266), .ZN(\SB1_0_25/i1[9] ) );
  INV_X4 U1229 ( .I(\SB2_0_24/i0[7] ), .ZN(\RI3[0][46] ) );
  INV_X2 \SB1_2_30/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[11] ), .ZN(
        \SB1_2_30/i1_5 ) );
  NAND2_X2 U1266 ( .A1(\SB1_0_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_0/Component_Function_0/NAND4_in[1] ), .ZN(n3034) );
  BUF_X2 U1301 ( .I(\SB3_2/buf_output[3] ), .Z(\SB4_0/i0[10] ) );
  NAND3_X2 \SB3_25/Component_Function_1/N3  ( .A1(\SB3_25/i1_5 ), .A2(
        \SB3_25/i0[6] ), .A3(\SB3_25/i0[9] ), .ZN(
        \SB3_25/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 U1968 ( .I(\SB2_4_27/buf_output[1] ), .Z(\RI5[4][49] ) );
  NAND3_X2 U1459 ( .A1(\SB2_4_0/i0_3 ), .A2(\SB2_4_0/i0_4 ), .A3(
        \SB2_4_0/i1[9] ), .ZN(\SB2_4_0/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB1_4_22/Component_Function_1/N4  ( .A1(\SB1_4_22/i1_7 ), .A2(
        \SB1_4_22/i0[8] ), .A3(\SB1_4_22/i0_4 ), .ZN(
        \SB1_4_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_10/Component_Function_0/N3  ( .A1(\SB2_2_10/i0[10] ), .A2(
        \SB2_2_10/i0_4 ), .A3(\SB2_2_10/i0_3 ), .ZN(
        \SB2_2_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB1_4_27/Component_Function_2/N2  ( .A1(\SB1_4_27/i0_3 ), .A2(
        \SB1_4_27/i0[10] ), .A3(\SB1_4_27/i0[6] ), .ZN(
        \SB1_4_27/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U1889 ( .I(\MC_ARK_ARC_1_4/buf_output[38] ), .ZN(\SB3_25/i1[9] ) );
  NAND3_X2 \SB2_4_29/Component_Function_2/N3  ( .A1(\SB2_4_29/i0_3 ), .A2(
        \SB2_4_29/i0[8] ), .A3(\SB2_4_29/i0[9] ), .ZN(
        \SB2_4_29/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U908 ( .I(\RI1[3][17] ), .ZN(\SB1_3_29/i1_5 ) );
  INV_X2 \SB1_0_21/INV_2  ( .I(n274), .ZN(\SB1_0_21/i1[9] ) );
  BUF_X2 U574 ( .I(\SB3_10/buf_output[1] ), .Z(\SB4_6/i0[6] ) );
  INV_X2 \SB2_1_14/INV_1  ( .I(\SB1_1_18/buf_output[1] ), .ZN(\SB2_1_14/i1_7 )
         );
  NAND3_X2 \SB2_4_12/Component_Function_0/N4  ( .A1(\SB2_4_12/i0[7] ), .A2(
        \SB2_4_12/i0_3 ), .A3(\SB2_4_12/i0_0 ), .ZN(
        \SB2_4_12/Component_Function_0/NAND4_in[3] ) );
  INV_X4 U1571 ( .I(n2554), .ZN(\SB1_4_31/buf_output[4] ) );
  NAND3_X2 U3985 ( .A1(\SB2_3_6/i0_3 ), .A2(\SB2_3_6/i0[6] ), .A3(
        \SB2_3_6/i1[9] ), .ZN(\SB2_3_6/Component_Function_3/NAND4_in[0] ) );
  INV_X2 \SB1_1_17/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[89] ), .ZN(
        \SB1_1_17/i1_5 ) );
  BUF_X4 \SB2_3_9/BUF_5  ( .I(\SB1_3_9/buf_output[5] ), .Z(\SB2_3_9/i0_3 ) );
  NAND3_X2 U1122 ( .A1(\SB1_1_3/i0[9] ), .A2(\SB1_1_3/i0_3 ), .A3(
        \SB1_1_3/i0[8] ), .ZN(n2021) );
  NAND2_X2 \SB1_1_0/Component_Function_5/N1  ( .A1(\SB1_1_0/i0_0 ), .A2(
        \SB1_1_0/i3[0] ), .ZN(\SB1_1_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_17/Component_Function_2/N1  ( .A1(\SB2_3_17/i1_5 ), .A2(
        \SB2_3_17/i0[10] ), .A3(\SB2_3_17/i1[9] ), .ZN(
        \SB2_3_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4912 ( .A1(\SB2_2_11/i0[8] ), .A2(\SB2_2_11/i3[0] ), .A3(
        \SB2_2_11/i1_5 ), .ZN(\SB2_2_11/Component_Function_3/NAND4_in[3] ) );
  NAND2_X2 \SB1_0_21/Component_Function_5/N1  ( .A1(\SB1_0_21/i0_0 ), .A2(
        \SB1_0_21/i3[0] ), .ZN(\SB1_0_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_14/Component_Function_3/N4  ( .A1(\SB2_1_14/i1_5 ), .A2(
        \SB2_1_14/i0[8] ), .A3(\SB2_1_14/i3[0] ), .ZN(
        \SB2_1_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U1570 ( .A1(\SB2_4_30/i0_3 ), .A2(\SB2_4_30/i0[8] ), .A3(
        \SB2_4_30/i0[9] ), .ZN(\SB2_4_30/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB2_1_16/BUF_3_0  ( .I(\SB2_1_16/buf_output[3] ), .Z(\RI5[1][105] )
         );
  NAND4_X2 U4235 ( .A1(\SB2_1_16/Component_Function_3/NAND4_in[0] ), .A2(n1212), .A3(n1211), .A4(n1210), .ZN(\SB2_1_16/buf_output[3] ) );
  NAND4_X2 \SB2_3_0/Component_Function_3/N5  ( .A1(
        \SB2_3_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_0/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_0/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_0/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_0/buf_output[3] ) );
  BUF_X2 U1079 ( .I(\SB1_1_8/buf_output[0] ), .Z(\SB2_1_3/i0[9] ) );
  BUF_X4 \SB1_0_21/BUF_2  ( .I(n274), .Z(\SB1_0_21/i0_0 ) );
  INV_X2 U4661 ( .I(\SB1_4_16/buf_output[5] ), .ZN(\SB2_4_16/i1_5 ) );
  NAND3_X2 U1516 ( .A1(\SB1_0_21/i0[10] ), .A2(\SB1_0_21/i1[9] ), .A3(
        \SB1_0_21/i1_7 ), .ZN(\SB1_0_21/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U2055 ( .I(\SB2_0_18/buf_output[4] ), .Z(\RI5[0][88] ) );
  NAND3_X2 \SB2_3_9/Component_Function_5/N3  ( .A1(\SB2_3_9/i1[9] ), .A2(
        \SB1_3_10/buf_output[4] ), .A3(\SB2_3_9/i0_3 ), .ZN(
        \SB2_3_9/Component_Function_5/NAND4_in[2] ) );
  INV_X4 U960 ( .I(n1102), .ZN(\SB2_2_18/i0_4 ) );
  NAND3_X2 \SB2_4_1/Component_Function_3/N4  ( .A1(n6277), .A2(\SB2_4_1/i0[8] ), .A3(\SB2_4_1/i3[0] ), .ZN(\SB2_4_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB3_13/Component_Function_0/N3  ( .A1(\SB3_13/i0[10] ), .A2(
        \SB3_13/i0_4 ), .A3(\SB3_13/i0_3 ), .ZN(
        \SB3_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_6/Component_Function_2/N1  ( .A1(\SB2_3_6/i1_5 ), .A2(
        \SB2_3_6/i0[10] ), .A3(\SB2_3_6/i1[9] ), .ZN(
        \SB2_3_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_4_16/Component_Function_3/N1  ( .A1(\SB2_4_16/i1[9] ), .A2(
        \SB2_4_16/i0_3 ), .A3(\SB2_4_16/i0[6] ), .ZN(
        \SB2_4_16/Component_Function_3/NAND4_in[0] ) );
  INV_X2 \SB2_3_28/INV_5  ( .I(\SB1_3_28/buf_output[5] ), .ZN(\SB2_3_28/i1_5 )
         );
  NAND2_X2 \SB1_3_28/Component_Function_5/N1  ( .A1(\SB1_3_28/i0_0 ), .A2(
        \SB1_3_28/i3[0] ), .ZN(\SB1_3_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U8425 ( .A1(\SB1_4_0/i0[8] ), .A2(\SB1_4_0/i1_5 ), .A3(
        \SB1_4_0/i3[0] ), .ZN(\SB1_4_0/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 U9122 ( .I(\SB2_3_23/buf_output[1] ), .Z(\RI5[3][73] ) );
  NAND3_X2 U924 ( .A1(\SB2_2_10/i0_3 ), .A2(\SB2_2_10/i0_0 ), .A3(
        \SB2_2_10/i0_4 ), .ZN(\SB2_2_10/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 U2024 ( .I(\SB1_2_11/buf_output[4] ), .Z(\SB2_2_10/i0_4 ) );
  BUF_X4 \SB2_4_1/BUF_4_0  ( .I(\SB2_4_1/buf_output[4] ), .Z(\RI5[4][190] ) );
  BUF_X4 U1980 ( .I(\SB1_4_12/buf_output[5] ), .Z(\SB2_4_12/i0_3 ) );
  INV_X2 U1801 ( .I(\MC_ARK_ARC_1_4/buf_output[176] ), .ZN(\SB3_2/i1[9] ) );
  BUF_X4 \SB2_0_21/BUF_5  ( .I(\RI3[0][65] ), .Z(\SB2_0_21/i0_3 ) );
  INV_X2 U1708 ( .I(\MC_ARK_ARC_1_1/buf_output[63] ), .ZN(\SB1_2_21/i0[8] ) );
  NAND3_X2 \SB3_2/Component_Function_2/N4  ( .A1(\SB3_2/i1_5 ), .A2(
        \SB3_2/i0_0 ), .A3(\SB3_2/i0_4 ), .ZN(
        \SB3_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U1884 ( .A1(\SB1_0_18/i0[6] ), .A2(\SB1_0_18/i0_3 ), .A3(
        \SB1_0_18/i1[9] ), .ZN(\SB1_0_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_28/Component_Function_5/N2  ( .A1(\SB1_2_28/i0_0 ), .A2(
        \SB1_2_28/i0[6] ), .A3(\SB1_2_28/i0[10] ), .ZN(
        \SB1_2_28/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U1827 ( .I(\SB2_1_19/buf_output[2] ), .Z(\RI5[1][92] ) );
  INV_X2 \SB1_4_18/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[83] ), .ZN(
        \SB1_4_18/i1_5 ) );
  NAND3_X2 U2189 ( .A1(\SB2_1_30/i1_5 ), .A2(\SB2_1_30/i0[10] ), .A3(
        \SB2_1_30/i1[9] ), .ZN(\SB2_1_30/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U7262 ( .I(\SB2_3_7/buf_output[1] ), .Z(\RI5[3][169] ) );
  BUF_X4 \SB1_2_29/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[14] ), .Z(
        \SB1_2_29/i0_0 ) );
  BUF_X4 \SB2_0_13/BUF_5  ( .I(\RI3[0][113] ), .Z(\SB2_0_13/i0_3 ) );
  NAND3_X2 U1321 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i1[9] ), .A3(
        \SB2_2_29/i0_4 ), .ZN(\SB2_2_29/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB2_4_20/INV_4  ( .I(\SB2_4_20/i0_4 ), .ZN(\SB2_4_20/i0[7] ) );
  NAND3_X2 \SB2_4_13/Component_Function_2/N3  ( .A1(\SB2_4_13/i0_3 ), .A2(
        \SB2_4_13/i0[8] ), .A3(\SB2_4_13/i0[9] ), .ZN(
        \SB2_4_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_26/Component_Function_3/N1  ( .A1(\SB2_2_26/i1[9] ), .A2(
        \SB2_2_26/i0_3 ), .A3(\SB2_2_26/i0[6] ), .ZN(
        \SB2_2_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U1602 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i0[10] ), .A3(\SB3_1/i0[6] ), 
        .ZN(\SB3_1/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U1686 ( .I(\MC_ARK_ARC_1_3/buf_output[113] ), .Z(\SB1_4_13/i0_3 ) );
  NAND3_X2 \SB2_1_23/Component_Function_2/N2  ( .A1(\SB2_1_23/i0_3 ), .A2(
        \SB2_1_23/i0[10] ), .A3(\SB2_1_23/i0[6] ), .ZN(
        \SB2_1_23/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U1685 ( .I(\MC_ARK_ARC_1_3/buf_output[113] ), .ZN(\SB1_4_13/i1_5 ) );
  NAND3_X2 \SB2_0_13/Component_Function_1/N2  ( .A1(\SB2_0_13/i0_3 ), .A2(
        \SB2_0_13/i1_7 ), .A3(\SB2_0_13/i0[8] ), .ZN(
        \SB2_0_13/Component_Function_1/NAND4_in[1] ) );
  INV_X2 U1410 ( .I(\MC_ARK_ARC_1_4/buf_output[171] ), .ZN(\SB3_3/i0[8] ) );
  BUF_X4 U5376 ( .I(\SB1_4_16/buf_output[5] ), .Z(\SB2_4_16/i0_3 ) );
  INV_X2 U5449 ( .I(\RI3[0][21] ), .ZN(\SB2_0_28/i0[8] ) );
  BUF_X4 \SB2_0_21/BUF_4  ( .I(\SB1_0_22/buf_output[4] ), .Z(\SB2_0_21/i0_4 )
         );
  NAND3_X2 \SB1_3_20/Component_Function_0/N4  ( .A1(\SB1_3_20/i0[7] ), .A2(
        \SB1_3_20/i0_3 ), .A3(\SB1_3_20/i0_0 ), .ZN(
        \SB1_3_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 \SB1_0_19/Component_Function_5/N2  ( .A1(\SB1_0_19/i0_0 ), .A2(
        \SB1_0_19/i0[6] ), .A3(\SB1_0_19/i0[10] ), .ZN(
        \SB1_0_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_7/Component_Function_1/N3  ( .A1(\SB2_2_7/i1_5 ), .A2(
        \SB2_2_7/i0[6] ), .A3(\SB2_2_7/i0[9] ), .ZN(
        \SB2_2_7/Component_Function_1/NAND4_in[2] ) );
  INV_X2 U1404 ( .I(\MC_ARK_ARC_1_4/buf_output[170] ), .ZN(\SB3_3/i1[9] ) );
  NAND3_X2 U810 ( .A1(\SB2_3_12/i0_3 ), .A2(\SB2_3_12/i0[9] ), .A3(
        \SB2_3_12/i0[10] ), .ZN(\SB2_3_12/Component_Function_4/NAND4_in[2] )
         );
  BUF_X4 \SB2_3_14/BUF_5  ( .I(\SB1_3_14/buf_output[5] ), .Z(\SB2_3_14/i0_3 )
         );
  NAND3_X2 \SB2_1_12/Component_Function_3/N1  ( .A1(\SB2_1_12/i1[9] ), .A2(
        \SB2_1_12/i0_3 ), .A3(\SB2_1_12/i0[6] ), .ZN(
        \SB2_1_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB1_0_6/Component_Function_3/N1  ( .A1(\SB1_0_6/i1[9] ), .A2(
        \SB1_0_6/i0_3 ), .A3(\SB1_0_6/i0[6] ), .ZN(
        \SB1_0_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U2296 ( .A1(\SB1_3_13/i3[0] ), .A2(\SB1_3_13/i0[8] ), .A3(
        \SB1_3_13/i1_5 ), .ZN(n715) );
  NAND3_X2 \SB2_2_5/Component_Function_3/N3  ( .A1(\SB2_2_5/i1[9] ), .A2(
        \SB2_2_5/i1_7 ), .A3(\SB2_2_5/i0[10] ), .ZN(
        \SB2_2_5/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U4991 ( .I(\MC_ARK_ARC_1_3/buf_output[143] ), .Z(\SB1_4_8/i0_3 ) );
  NAND3_X2 \SB2_0_26/Component_Function_5/N4  ( .A1(\SB2_0_26/i0[9] ), .A2(
        \SB2_0_26/i0[6] ), .A3(\SB2_0_26/i0_4 ), .ZN(
        \SB2_0_26/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \SB2_0_4/BUF_1_0  ( .I(\SB2_0_4/buf_output[1] ), .Z(\RI5[0][187] ) );
  INV_X2 \SB1_0_19/INV_2  ( .I(n278), .ZN(\SB1_0_19/i1[9] ) );
  NAND2_X2 \SB2_2_24/Component_Function_1/N1  ( .A1(\SB2_2_24/i0_3 ), .A2(
        \SB2_2_24/i1[9] ), .ZN(\SB2_2_24/Component_Function_1/NAND4_in[0] ) );
  INV_X2 U1577 ( .I(\MC_ARK_ARC_1_3/buf_output[165] ), .ZN(\SB1_4_4/i0[8] ) );
  NAND3_X2 U3828 ( .A1(\SB2_3_19/i0[9] ), .A2(\SB2_3_19/i0[6] ), .A3(
        \SB1_3_20/buf_output[4] ), .ZN(
        \SB2_3_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U7479 ( .A1(\SB1_0_12/i0_4 ), .A2(\SB1_0_12/i0[9] ), .A3(
        \SB1_0_12/i0[6] ), .ZN(n2413) );
  NAND3_X2 U2308 ( .A1(\SB1_3_15/i0_3 ), .A2(\SB1_3_15/i0[8] ), .A3(
        \SB1_3_15/i0[9] ), .ZN(\SB1_3_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_23/Component_Function_2/N1  ( .A1(\SB2_2_23/i1_5 ), .A2(
        \SB2_2_23/i0[10] ), .A3(\SB2_2_23/i1[9] ), .ZN(
        \SB2_2_23/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 \SB1_1_2/Component_Function_5/N1  ( .A1(\SB1_1_2/i0_0 ), .A2(
        \SB1_1_2/i3[0] ), .ZN(\SB1_1_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_23/Component_Function_0/N3  ( .A1(\SB2_2_23/i0[10] ), .A2(
        n600), .A3(\SB2_2_23/i0_3 ), .ZN(
        \SB2_2_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_21/Component_Function_3/N1  ( .A1(\SB2_0_21/i1[9] ), .A2(
        \SB2_0_21/i0_3 ), .A3(\SB2_0_21/i0[6] ), .ZN(
        \SB2_0_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_21/Component_Function_3/N4  ( .A1(\SB2_0_21/i1_5 ), .A2(
        \SB2_0_21/i0[8] ), .A3(\SB2_0_21/i3[0] ), .ZN(
        \SB2_0_21/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 U1916 ( .I(\MC_ARK_ARC_1_0/buf_output[65] ), .Z(\SB1_1_21/i0_3 ) );
  NAND2_X2 U1875 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i3[0] ), .ZN(
        \SB1_2_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_21/Component_Function_1/N4  ( .A1(\SB2_0_21/i1_7 ), .A2(
        \SB2_0_21/i0[8] ), .A3(\SB2_0_21/i0_4 ), .ZN(
        \SB2_0_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U1044 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0[8] ), .A3(
        \SB2_1_9/i1_7 ), .ZN(n2378) );
  NAND3_X2 U710 ( .A1(\SB1_4_28/i0[10] ), .A2(\SB1_4_28/i0_0 ), .A3(
        \SB1_4_28/i0[6] ), .ZN(\SB1_4_28/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_37  ( .I(\SB2_1_29/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[37] ) );
  BUF_X4 U5340 ( .I(\SB1_0_30/buf_output[5] ), .Z(\SB2_0_30/i0_3 ) );
  BUF_X4 U1824 ( .I(\SB1_1_9/buf_output[5] ), .Z(\SB2_1_9/i0_3 ) );
  NAND3_X2 \SB1_0_21/Component_Function_3/N2  ( .A1(\SB1_0_21/i0_0 ), .A2(
        \SB1_0_21/i0_3 ), .A3(\SB1_0_21/i0_4 ), .ZN(
        \SB1_0_21/Component_Function_3/NAND4_in[1] ) );
  NAND2_X2 U720 ( .A1(\SB1_4_28/i0_0 ), .A2(\SB1_4_28/i3[0] ), .ZN(n1311) );
  NAND3_X2 U7203 ( .A1(\SB1_0_29/i0[10] ), .A2(\SB1_0_29/i1[9] ), .A3(
        \SB1_0_29/i1_7 ), .ZN(\SB1_0_29/Component_Function_3/NAND4_in[2] ) );
  INV_X2 \SB1_0_29/INV_2  ( .I(n258), .ZN(\SB1_0_29/i1[9] ) );
  NAND3_X2 \SB1_4_4/Component_Function_2/N3  ( .A1(\SB1_4_4/i0_3 ), .A2(
        \SB1_4_4/i0[8] ), .A3(\SB1_4_4/i0[9] ), .ZN(
        \SB1_4_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U936 ( .A1(\SB2_2_5/i0_0 ), .A2(\SB2_2_5/i1_5 ), .A3(\SB2_2_5/i0_4 ), .ZN(\SB2_2_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_1_20/Component_Function_2/N1  ( .A1(\SB2_1_20/i1_5 ), .A2(
        \SB2_1_20/i0[10] ), .A3(\SB2_1_20/i1[9] ), .ZN(
        \SB2_1_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_4/Component_Function_3/N4  ( .A1(\SB2_1_4/i1_5 ), .A2(
        \SB2_1_4/i0[8] ), .A3(\SB2_1_4/i3[0] ), .ZN(
        \SB2_1_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_1_24/Component_Function_3/N4  ( .A1(\SB1_1_24/i1_5 ), .A2(
        \SB1_1_24/i0[8] ), .A3(\SB1_1_24/i3[0] ), .ZN(
        \SB1_1_24/Component_Function_3/NAND4_in[3] ) );
  INV_X2 U1807 ( .I(\RI1[3][5] ), .ZN(\SB1_3_31/i1_5 ) );
  BUF_X4 \SB2_1_26/BUF_5  ( .I(\SB1_1_26/buf_output[5] ), .Z(\SB2_1_26/i0_3 )
         );
  NAND3_X2 U937 ( .A1(\SB2_2_10/i0[10] ), .A2(\SB2_2_10/i0_3 ), .A3(
        \SB2_2_10/i0[6] ), .ZN(\SB2_2_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U2396 ( .A1(\SB2_4_13/i1_5 ), .A2(\SB2_4_13/i0[8] ), .A3(
        \SB2_4_13/i3[0] ), .ZN(\SB2_4_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U2262 ( .A1(\SB2_2_31/i1[9] ), .A2(\SB2_2_31/i1_7 ), .A3(
        \SB2_2_31/i0[10] ), .ZN(\SB2_2_31/Component_Function_3/NAND4_in[2] )
         );
  NAND2_X2 U2103 ( .A1(\SB1_0_19/i0_0 ), .A2(\SB1_0_19/i3[0] ), .ZN(
        \SB1_0_19/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_0_2/BUF_5  ( .I(\RI3[0][179] ), .Z(\SB2_0_2/i0_3 ) );
  NAND3_X2 \SB2_1_4/Component_Function_1/N4  ( .A1(n2656), .A2(\SB2_1_4/i0[8] ), .A3(\SB2_1_4/i0_4 ), .ZN(\SB2_1_4/Component_Function_1/NAND4_in[3] ) );
  NAND2_X2 \SB1_0_4/Component_Function_5/N1  ( .A1(\SB1_0_4/i0_0 ), .A2(
        \SB1_0_4/i3[0] ), .ZN(\SB1_0_4/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_1/Component_Function_1/N1  ( .A1(\SB2_2_1/i0_3 ), .A2(
        \SB2_2_1/i1[9] ), .ZN(\SB2_2_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U804 ( .A1(\SB2_3_25/i0[10] ), .A2(\SB2_3_25/i1_7 ), .A3(
        \SB2_3_25/i1[9] ), .ZN(n3106) );
  NAND3_X2 \SB1_4_27/Component_Function_3/N2  ( .A1(\RI1[4][26] ), .A2(
        \SB1_4_27/i0_3 ), .A3(\SB1_4_27/i0_4 ), .ZN(
        \SB1_4_27/Component_Function_3/NAND4_in[1] ) );
  INV_X2 \SB1_4_27/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[29] ), .ZN(
        \SB1_4_27/i1_5 ) );
  NAND3_X2 \SB2_1_20/Component_Function_1/N3  ( .A1(\SB2_1_20/i1_5 ), .A2(
        \SB2_1_20/i0[6] ), .A3(\SB2_1_20/i0[9] ), .ZN(
        \SB2_1_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_8/Component_Function_2/N3  ( .A1(\SB1_1_8/i0_3 ), .A2(
        \SB1_1_8/i0[8] ), .A3(\SB1_1_8/i0[9] ), .ZN(
        \SB1_1_8/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 \SB1_2_16/Component_Function_5/N1  ( .A1(\SB1_2_16/i0_0 ), .A2(
        \SB1_2_16/i3[0] ), .ZN(\SB1_2_16/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB2_3_26/INV_5  ( .I(\SB1_3_26/buf_output[5] ), .ZN(\SB2_3_26/i1_5 )
         );
  NAND3_X2 U1600 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i1[9] ), .A3(\SB3_1/i0_4 ), 
        .ZN(\SB3_1/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U2034 ( .I(\SB2_1_7/buf_output[0] ), .Z(\RI5[1][174] ) );
  NAND3_X2 U94 ( .A1(\SB4_0/i0_4 ), .A2(\SB4_0/i1[9] ), .A3(\SB4_0/i1_5 ), 
        .ZN(n1801) );
  BUF_X2 U1082 ( .I(\SB2_1_4/i1_7 ), .Z(n2656) );
  BUF_X4 \SB3_8/BUF_5  ( .I(\MC_ARK_ARC_1_4/buf_output[143] ), .Z(\SB3_8/i0_3 ) );
  NAND3_X2 \SB1_4_27/Component_Function_1/N4  ( .A1(\SB1_4_27/i1_7 ), .A2(
        \SB1_4_27/i0[8] ), .A3(\SB1_4_27/i0_4 ), .ZN(
        \SB1_4_27/Component_Function_1/NAND4_in[3] ) );
  INV_X2 \SB1_0_21/INV_5  ( .I(n3985), .ZN(\SB1_0_21/i1_5 ) );
  NAND3_X2 \SB1_0_21/Component_Function_3/N1  ( .A1(\SB1_0_21/i1[9] ), .A2(
        \SB1_0_21/i0_3 ), .A3(\SB1_0_21/i0[6] ), .ZN(
        \SB1_0_21/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U7631 ( .I(\SB1_2_6/buf_output[5] ), .ZN(\SB2_2_6/i1_5 ) );
  INV_X8 \SB2_0_19/INV_3  ( .I(\RI3[0][75] ), .ZN(\SB2_0_19/i0[8] ) );
  NAND3_X2 U1633 ( .A1(\SB2_0_0/i1_5 ), .A2(\SB2_0_0/i0[10] ), .A3(
        \SB2_0_0/i1[9] ), .ZN(\SB2_0_0/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_4_16/BUF_4  ( .I(\SB1_4_17/buf_output[4] ), .Z(\SB2_4_16/i0_4 )
         );
  NAND3_X2 \SB2_1_24/Component_Function_2/N2  ( .A1(\SB2_1_24/i0_3 ), .A2(
        \SB2_1_24/i0[10] ), .A3(\SB2_1_24/i0[6] ), .ZN(
        \SB2_1_24/Component_Function_2/NAND4_in[1] ) );
  BUF_X2 \SB1_2_18/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[79] ), .Z(
        \SB1_2_18/i0[6] ) );
  NAND3_X2 \SB1_1_2/Component_Function_2/N3  ( .A1(\SB1_1_2/i0_3 ), .A2(
        \SB1_1_2/i0[8] ), .A3(\SB1_1_2/i0[9] ), .ZN(
        \SB1_1_2/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U2254 ( .I(\SB1_2_21/buf_output[4] ), .Z(\SB2_2_20/i0_4 ) );
  NAND3_X2 \SB1_0_20/Component_Function_0/N2  ( .A1(\SB1_0_20/i0[8] ), .A2(
        \SB1_0_20/i0[7] ), .A3(\SB1_0_20/i0[6] ), .ZN(
        \SB1_0_20/Component_Function_0/NAND4_in[1] ) );
  BUF_X4 U2122 ( .I(\SB1_0_4/buf_output[4] ), .Z(\RI3[0][172] ) );
  INV_X2 \SB2_0_7/INV_5  ( .I(\RI3[0][149] ), .ZN(\SB2_0_7/i1_5 ) );
  BUF_X4 U1907 ( .I(n390), .Z(\SB1_0_22/i0_3 ) );
  BUF_X4 U1771 ( .I(\MC_ARK_ARC_1_1/buf_output[109] ), .Z(\SB1_2_13/i0[6] ) );
  NAND3_X2 \SB1_4_3/Component_Function_5/N2  ( .A1(\SB1_4_3/i0_0 ), .A2(
        \SB1_4_3/i0[6] ), .A3(\SB1_4_3/i0[10] ), .ZN(
        \SB1_4_3/Component_Function_5/NAND4_in[1] ) );
  NAND2_X2 \SB2_2_7/Component_Function_5/N1  ( .A1(\SB2_2_7/i0_0 ), .A2(
        \SB2_2_7/i3[0] ), .ZN(\SB2_2_7/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U1974 ( .I(\SB1_4_30/buf_output[5] ), .Z(\SB2_4_30/i0_3 ) );
  NAND3_X2 \SB2_0_21/Component_Function_1/N2  ( .A1(\SB2_0_21/i0_3 ), .A2(
        \SB2_0_21/i1_7 ), .A3(\SB2_0_21/i0[8] ), .ZN(
        \SB2_0_21/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U8930 ( .I(\SB2_1_17/buf_output[1] ), .Z(\RI5[1][109] ) );
  NAND4_X2 U6027 ( .A1(\SB2_1_17/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_17/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_17/buf_output[1] ) );
  NAND4_X2 \SB2_1_7/Component_Function_1/N5  ( .A1(
        \SB2_1_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_7/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_1_7/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_7/buf_output[1] ) );
  CLKBUF_X2 U15 ( .I(Key[116]), .Z(n205) );
  NAND3_X2 U807 ( .A1(\SB2_3_2/i0_3 ), .A2(\SB2_3_2/i1_7 ), .A3(
        \SB2_3_2/i0[8] ), .ZN(n1048) );
  BUF_X4 U2155 ( .I(\MC_ARK_ARC_1_0/buf_output[119] ), .Z(\SB1_1_12/i0_3 ) );
  INV_X2 U1779 ( .I(\MC_ARK_ARC_1_0/buf_output[95] ), .ZN(\SB1_1_16/i1_5 ) );
  NAND3_X2 U8733 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i0[9] ), .A3(\SB3_1/i0[10] ), 
        .ZN(\SB3_1/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 \SB1_3_2/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[176] ), .Z(
        \SB1_3_2/i0_0 ) );
  BUF_X4 U9199 ( .I(\SB2_4_4/buf_output[1] ), .Z(\RI5[4][187] ) );
  NAND4_X2 \SB2_4_4/Component_Function_1/N5  ( .A1(
        \SB2_4_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_4/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_4_4/buf_output[1] ) );
  NAND3_X2 U1234 ( .A1(\SB1_0_25/i0[10] ), .A2(\SB1_0_25/i0_0 ), .A3(
        \SB1_0_25/i0[6] ), .ZN(n2294) );
  BUF_X4 \SB2_0_11/BUF_1_0  ( .I(\SB2_0_11/buf_output[1] ), .Z(\RI5[0][145] )
         );
  NAND4_X2 \SB2_0_11/Component_Function_1/N5  ( .A1(
        \SB2_0_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_11/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_11/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_11/buf_output[1] ) );
  INV_X2 \SB2_0_25/INV_5  ( .I(\RI3[0][41] ), .ZN(\SB2_0_25/i1_5 ) );
  BUF_X4 \SB2_1_25/BUF_3_0  ( .I(\SB2_1_25/buf_output[3] ), .Z(\RI5[1][51] )
         );
  NAND3_X2 U809 ( .A1(\SB2_3_3/i0[10] ), .A2(\SB2_3_3/i1_7 ), .A3(
        \SB2_3_3/i1[9] ), .ZN(\SB2_3_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U1191 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0_4 ), .A3(
        \SB2_0_5/i1[9] ), .ZN(n1771) );
  NAND3_X2 \SB2_4_17/Component_Function_2/N4  ( .A1(\SB2_4_17/i1_5 ), .A2(
        \SB2_4_17/i0_0 ), .A3(\SB2_4_17/i0_4 ), .ZN(
        \SB2_4_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U1507 ( .A1(\RI1[4][119] ), .A2(\SB1_4_12/i1[9] ), .A3(
        \SB1_4_12/i0_4 ), .ZN(\SB1_4_12/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_1_23/BUF_5  ( .I(\SB1_1_23/buf_output[5] ), .Z(\SB2_1_23/i0_3 )
         );
  NAND3_X2 U2368 ( .A1(\SB1_4_3/i0[10] ), .A2(\SB1_4_3/i1[9] ), .A3(
        \SB1_4_3/i1_7 ), .ZN(n1101) );
  BUF_X4 U8844 ( .I(\SB2_0_20/buf_output[2] ), .Z(\RI5[0][86] ) );
  NAND4_X2 \SB2_0_20/Component_Function_2/N5  ( .A1(
        \SB2_0_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_20/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_20/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_20/buf_output[2] ) );
  NAND3_X2 \SB3_17/Component_Function_5/N2  ( .A1(\SB3_17/i0_0 ), .A2(
        \SB3_17/i0[6] ), .A3(\SB3_17/i0[10] ), .ZN(
        \SB3_17/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB1_3_5/BUF_5  ( .I(\RI1[3][161] ), .Z(\SB1_3_5/i0_3 ) );
  NAND4_X2 U2752 ( .A1(\SB1_4_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_4_27/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_4_27/Component_Function_2/NAND4_in[1] ), .A4(n3069), .ZN(
        \SB1_4_27/buf_output[2] ) );
  INV_X2 U1631 ( .I(\MC_ARK_ARC_1_0/buf_output[50] ), .ZN(\SB1_1_23/i1[9] ) );
  NAND4_X2 \SB2_0_7/Component_Function_3/N5  ( .A1(
        \SB2_0_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_7/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_7/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_7/buf_output[3] ) );
  NAND3_X2 U5041 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i0[10] ), .A3(\SB3_2/i0[6] ), 
        .ZN(\SB3_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB1_1_0/Component_Function_0/N4  ( .A1(\SB1_1_0/i0[7] ), .A2(
        \SB1_1_0/i0_3 ), .A3(\SB1_1_0/i0_0 ), .ZN(
        \SB1_1_0/Component_Function_0/NAND4_in[3] ) );
  BUF_X2 \SB3_17/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[84] ), .Z(
        \SB3_17/i0[9] ) );
  INV_X2 U1795 ( .I(\MC_ARK_ARC_1_2/buf_output[29] ), .ZN(\SB1_3_27/i1_5 ) );
  INV_X2 U1895 ( .I(\MC_ARK_ARC_1_0/buf_output[53] ), .ZN(\SB1_1_23/i1_5 ) );
  BUF_X4 U1794 ( .I(\MC_ARK_ARC_1_2/buf_output[29] ), .Z(\SB1_3_27/i0_3 ) );
  INV_X2 U1230 ( .I(\RI3[0][179] ), .ZN(\SB2_0_2/i1_5 ) );
  CLKBUF_X2 U175 ( .I(Key[181]), .Z(n118) );
  NAND2_X2 \SB2_4_31/Component_Function_5/N1  ( .A1(\SB2_4_31/i0_0 ), .A2(
        \SB2_4_31/i3[0] ), .ZN(\SB2_4_31/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U790 ( .I(\SB2_3_14/buf_output[1] ), .Z(\RI5[3][127] ) );
  NAND2_X2 \SB1_2_30/Component_Function_5/N1  ( .A1(\SB1_2_30/i0_0 ), .A2(
        \SB1_2_30/i3[0] ), .ZN(\SB1_2_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U985 ( .A1(\SB1_2_30/i0[10] ), .A2(\SB1_2_30/i0_0 ), .A3(
        \SB1_2_30/i0[6] ), .ZN(\SB1_2_30/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U1758 ( .A1(\SB2_2_30/i0_0 ), .A2(\SB2_2_30/i0_3 ), .A3(
        \SB2_2_30/i0_4 ), .ZN(\SB2_2_30/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB2_0_10/BUF_5  ( .I(\RI3[0][131] ), .Z(\SB2_0_10/i0_3 ) );
  NAND4_X2 U1175 ( .A1(\SB2_0_2/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_2/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_2/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_2/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_2/buf_output[0] ) );
  INV_X2 U1344 ( .I(\MC_ARK_ARC_1_0/buf_output[75] ), .ZN(\SB1_1_19/i0[8] ) );
  INV_X2 U5468 ( .I(n343), .ZN(\SB1_0_18/i0[8] ) );
  BUF_X4 U5267 ( .I(\SB1_3_20/buf_output[5] ), .Z(\SB2_3_20/i0_3 ) );
  BUF_X4 \SB1_3_31/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[2] ), .Z(
        \SB1_3_31/i0_0 ) );
  NAND2_X2 \SB1_2_8/Component_Function_5/N1  ( .A1(\SB1_2_8/i0_0 ), .A2(
        \SB1_2_8/i3[0] ), .ZN(\SB1_2_8/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB1_4_24/BUF_5  ( .I(\MC_ARK_ARC_1_3/buf_output[47] ), .Z(
        \SB1_4_24/i0_3 ) );
  NAND3_X2 \SB1_0_23/Component_Function_3/N3  ( .A1(\SB1_0_23/i1[9] ), .A2(
        \SB1_0_23/i1_7 ), .A3(\SB1_0_23/i0[10] ), .ZN(
        \SB1_0_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_23/Component_Function_2/N3  ( .A1(\SB2_0_23/i0_3 ), .A2(
        \SB2_0_23/i0[8] ), .A3(\SB2_0_23/i0[9] ), .ZN(
        \SB2_0_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U1762 ( .A1(\SB1_4_20/i0[10] ), .A2(\SB1_4_20/i1[9] ), .A3(
        \SB1_4_20/i1_7 ), .ZN(n1793) );
  NAND3_X2 \SB1_1_30/Component_Function_0/N4  ( .A1(\SB1_1_30/i0[7] ), .A2(
        \SB1_1_30/i0_3 ), .A3(\SB1_1_30/i0_0 ), .ZN(
        \SB1_1_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U821 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i1[9] ), .A3(
        \SB2_3_16/i0_4 ), .ZN(\SB2_3_16/Component_Function_5/NAND4_in[2] ) );
  NAND2_X2 U1506 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i1[9] ), .ZN(
        \SB2_1_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_4/Component_Function_2/N2  ( .A1(\SB2_2_4/i0_3 ), .A2(
        \SB2_2_4/i0[10] ), .A3(\SB2_2_4/i0[6] ), .ZN(
        \SB2_2_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_15/Component_Function_2/N2  ( .A1(\SB2_1_15/i0_3 ), .A2(
        \SB2_1_15/i0[10] ), .A3(\SB2_1_15/i0[6] ), .ZN(
        \SB2_1_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U4804 ( .A1(\SB2_2_2/i0[10] ), .A2(\SB2_2_2/i1_5 ), .A3(n6267), 
        .ZN(\SB2_2_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_8/Component_Function_3/N3  ( .A1(\SB2_0_8/i1[9] ), .A2(
        \SB2_0_8/i1_7 ), .A3(\SB2_0_8/i0[10] ), .ZN(
        \SB2_0_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_23/Component_Function_3/N2  ( .A1(\SB1_1_23/i0_0 ), .A2(
        \SB1_1_23/i0_3 ), .A3(\SB1_1_23/i0_4 ), .ZN(
        \SB1_1_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_8/Component_Function_2/N1  ( .A1(\SB2_0_8/i1_5 ), .A2(
        \SB2_0_8/i0[10] ), .A3(\SB2_0_8/i1[9] ), .ZN(
        \SB2_0_8/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 \SB2_0_14/Component_Function_0/N5  ( .A1(
        \SB2_0_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_14/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_0_14/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_0_14/buf_output[0] ) );
  BUF_X4 \SB2_0_8/BUF_3  ( .I(\RI3[0][141] ), .Z(\SB2_0_8/i0[10] ) );
  BUF_X4 U8644 ( .I(\SB2_1_8/buf_output[2] ), .Z(\RI5[1][158] ) );
  BUF_X4 U8944 ( .I(\SB2_1_29/buf_output[3] ), .Z(\RI5[1][27] ) );
  BUF_X4 \SB2_0_14/BUF_0_0  ( .I(\SB2_0_14/buf_output[0] ), .Z(\RI5[0][132] )
         );
  NAND2_X2 \SB1_2_23/Component_Function_5/N1  ( .A1(\SB1_2_23/i0_0 ), .A2(
        \SB1_2_23/i3[0] ), .ZN(\SB1_2_23/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_3_28/BUF_5  ( .I(\SB1_3_28/buf_output[5] ), .Z(\SB2_3_28/i0_3 )
         );
  NAND3_X1 \SB3_23/Component_Function_3/N3  ( .A1(\SB3_23/i1[9] ), .A2(
        \SB3_23/i1_7 ), .A3(\SB3_23/i0[10] ), .ZN(
        \SB3_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U1201 ( .A1(\SB2_0_2/i0[10] ), .A2(\SB2_0_2/i0_0 ), .A3(
        \SB2_0_2/i0[6] ), .ZN(n1587) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_3  ( .I(\SB2_1_1/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[3] ) );
  NAND3_X2 U4773 ( .A1(\SB3_1/i0[6] ), .A2(\SB3_1/i0_0 ), .A3(\SB3_1/i0[10] ), 
        .ZN(\SB3_1/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U1822 ( .I(n6278), .ZN(\SB1_1_31/i1_5 ) );
  NAND3_X2 \SB2_1_14/Component_Function_3/N3  ( .A1(\SB2_1_14/i1[9] ), .A2(
        \SB2_1_14/i1_7 ), .A3(\SB2_1_14/i0[10] ), .ZN(
        \SB2_1_14/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB1_1_29/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[14] ), .Z(
        \SB1_1_29/i0_0 ) );
  BUF_X4 \SB3_28/BUF_5  ( .I(\MC_ARK_ARC_1_4/buf_output[23] ), .Z(
        \SB3_28/i0_3 ) );
  NAND3_X2 \SB2_0_8/Component_Function_2/N3  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \SB2_0_8/i0[8] ), .A3(\SB2_0_8/i0[9] ), .ZN(
        \SB2_0_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_28/Component_Function_3/N1  ( .A1(\SB2_1_28/i1[9] ), .A2(
        \SB2_1_28/i0_3 ), .A3(\SB2_1_28/i0[6] ), .ZN(
        \SB2_1_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_19/Component_Function_2/N4  ( .A1(\SB2_2_19/i1_5 ), .A2(
        \SB2_2_19/i0_0 ), .A3(\SB2_2_19/i0_4 ), .ZN(
        \SB2_2_19/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 U1983 ( .I(n5424), .Z(\SB1_4_9/i0_3 ) );
  NAND3_X2 U890 ( .A1(\SB1_3_27/i0[10] ), .A2(\SB1_3_27/i1[9] ), .A3(
        \SB1_3_27/i1_7 ), .ZN(n2763) );
  BUF_X2 U73 ( .I(Key[120]), .Z(n29) );
  BUF_X4 \SB2_0_4/BUF_2_0  ( .I(\SB2_0_4/buf_output[2] ), .Z(\RI5[0][182] ) );
  NAND3_X2 \SB2_4_17/Component_Function_3/N1  ( .A1(\SB2_4_17/i1[9] ), .A2(
        \SB2_4_17/i0_3 ), .A3(\SB2_4_17/i0[6] ), .ZN(
        \SB2_4_17/Component_Function_3/NAND4_in[0] ) );
  INV_X4 U910 ( .I(n3100), .ZN(\SB1_3_27/i0_4 ) );
  NAND3_X2 \SB2_4_26/Component_Function_3/N2  ( .A1(\SB2_4_26/i0_0 ), .A2(
        \SB2_4_26/i0_3 ), .A3(\SB2_4_26/i0_4 ), .ZN(
        \SB2_4_26/Component_Function_3/NAND4_in[1] ) );
  NAND2_X2 \SB1_1_24/Component_Function_5/N1  ( .A1(\SB1_1_24/i0_0 ), .A2(
        \SB1_1_24/i3[0] ), .ZN(\SB1_1_24/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U5266 ( .I(\SB1_2_4/buf_output[5] ), .Z(\SB2_2_4/i0_3 ) );
  BUF_X4 U1751 ( .I(\SB1_1_10/buf_output[5] ), .Z(\SB2_1_10/i0_3 ) );
  INV_X2 U1376 ( .I(\MC_ARK_ARC_1_4/buf_output[182] ), .ZN(\SB3_1/i1[9] ) );
  BUF_X4 \SB1_0_28/BUF_4_0  ( .I(\SB1_0_28/buf_output[4] ), .Z(\RI3[0][28] )
         );
  BUF_X4 \SB2_0_27/BUF_1_0  ( .I(\SB2_0_27/buf_output[1] ), .Z(\RI5[0][49] )
         );
  NAND3_X2 \SB2_2_12/Component_Function_3/N3  ( .A1(\SB2_2_12/i1[9] ), .A2(
        \SB2_2_12/i1_7 ), .A3(\SB2_2_12/i0[10] ), .ZN(
        \SB2_2_12/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB1_4_29/BUF_2  ( .I(\MC_ARK_ARC_1_3/buf_output[14] ), .Z(
        \SB1_4_29/i0_0 ) );
  INV_X2 \SB2_1_8/INV_5  ( .I(\SB1_1_8/buf_output[5] ), .ZN(\SB2_1_8/i1_5 ) );
  NAND3_X2 \SB1_1_7/Component_Function_3/N4  ( .A1(\SB1_1_7/i1_5 ), .A2(
        \SB1_1_7/i0[8] ), .A3(\SB1_1_7/i3[0] ), .ZN(
        \SB1_1_7/Component_Function_3/NAND4_in[3] ) );
  INV_X2 U5190 ( .I(\MC_ARK_ARC_1_3/buf_output[50] ), .ZN(\SB1_4_23/i1[9] ) );
  BUF_X4 \SB1_1_14/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[103] ), .Z(
        \SB1_1_14/i0[6] ) );
  BUF_X4 \SB2_2_16/BUF_1  ( .I(\SB1_2_20/buf_output[1] ), .Z(\SB2_2_16/i0[6] )
         );
  CLKBUF_X2 U18 ( .I(Key[154]), .Z(n211) );
  CLKBUF_X2 U225 ( .I(Key[104]), .Z(n175) );
  INV_X4 U4776 ( .I(n1427), .ZN(\RI3[3][64] ) );
  NAND3_X2 \SB2_1_8/Component_Function_2/N1  ( .A1(\SB2_1_8/i1_5 ), .A2(
        \SB2_1_8/i0[10] ), .A3(\SB2_1_8/i1[9] ), .ZN(
        \SB2_1_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_13/Component_Function_1/N2  ( .A1(\SB1_1_13/i0_3 ), .A2(
        \SB1_1_13/i1_7 ), .A3(\SB1_1_13/i0[8] ), .ZN(
        \SB1_1_13/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \SB2_3_16/BUF_4  ( .I(\SB1_3_17/buf_output[4] ), .Z(\SB2_3_16/i0_4 )
         );
  BUF_X4 \SB2_0_30/BUF_4_0  ( .I(\SB2_0_30/buf_output[4] ), .Z(\RI5[0][16] )
         );
  NAND3_X2 \SB2_2_20/Component_Function_3/N1  ( .A1(\SB2_2_20/i1[9] ), .A2(
        \SB2_2_20/i0_3 ), .A3(\SB2_2_20/i0[6] ), .ZN(
        \SB2_2_20/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_0_30/BUF_3  ( .I(\RI3[0][9] ), .Z(\SB2_0_30/i0[10] ) );
  BUF_X4 U2023 ( .I(\SB1_2_29/buf_output[4] ), .Z(\SB2_2_28/i0_4 ) );
  NAND2_X2 \SB1_1_30/Component_Function_5/N1  ( .A1(\SB1_1_30/i0_0 ), .A2(
        \SB1_1_30/i3[0] ), .ZN(\SB1_1_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_13/Component_Function_1/N4  ( .A1(\SB1_1_13/i1_7 ), .A2(
        \SB1_1_13/i0[8] ), .A3(\SB1_1_13/i0_4 ), .ZN(
        \SB1_1_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U2138 ( .A1(\SB2_0_26/i0[9] ), .A2(\SB2_0_26/i0_0 ), .A3(
        \SB2_0_26/i0[8] ), .ZN(\SB2_0_26/Component_Function_4/NAND4_in[0] ) );
  INV_X2 \SB2_1_26/INV_1  ( .I(\SB1_1_30/buf_output[1] ), .ZN(\SB2_1_26/i1_7 )
         );
  BUF_X4 U1846 ( .I(\MC_ARK_ARC_1_0/buf_output[185] ), .Z(\SB1_1_1/i0_3 ) );
  NAND3_X2 \SB1_1_19/Component_Function_3/N2  ( .A1(\SB1_1_19/i0_0 ), .A2(
        \SB1_1_19/i0_3 ), .A3(\SB1_1_19/i0_4 ), .ZN(
        \SB1_1_19/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB2_0_28/BUF_2_0  ( .I(\SB2_0_28/buf_output[2] ), .Z(\RI5[0][38] )
         );
  BUF_X4 U8933 ( .I(\SB2_1_19/buf_output[1] ), .Z(\RI5[1][97] ) );
  CLKBUF_X4 U1872 ( .I(\MC_ARK_ARC_1_0/buf_output[189] ), .Z(\SB1_1_0/i0[10] )
         );
  CLKBUF_X2 U120 ( .I(Key[61]), .Z(n48) );
  NAND3_X2 \SB2_2_14/Component_Function_2/N3  ( .A1(\SB2_2_14/i0_3 ), .A2(
        \SB2_2_14/i0[8] ), .A3(\SB2_2_14/i0[9] ), .ZN(
        \SB2_2_14/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB2_4_31/BUF_4_0  ( .I(\SB2_4_31/buf_output[4] ), .Z(\RI5[4][10] )
         );
  NAND3_X2 U6485 ( .A1(\SB2_2_25/i0_0 ), .A2(\SB2_2_25/i0_4 ), .A3(
        \SB2_2_25/i1_5 ), .ZN(n1965) );
  BUF_X4 U9038 ( .I(\SB2_2_21/buf_output[3] ), .Z(\RI5[2][75] ) );
  NAND4_X2 U5793 ( .A1(\SB2_2_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_21/Component_Function_3/NAND4_in[1] ), .A3(n1654), .A4(
        \SB2_2_21/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_21/buf_output[3] ) );
  INV_X2 U1083 ( .I(\SB1_1_12/buf_output[5] ), .ZN(\SB2_1_12/i1_5 ) );
  BUF_X4 U9022 ( .I(\SB2_2_15/buf_output[3] ), .Z(\RI5[2][111] ) );
  NAND3_X2 U1725 ( .A1(\SB2_4_1/i0[9] ), .A2(\SB2_4_1/i0_4 ), .A3(
        \SB2_4_1/i0[6] ), .ZN(\SB2_4_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB1_1_16/Component_Function_0/N4  ( .A1(\SB1_1_16/i0[7] ), .A2(
        \SB1_1_16/i0_3 ), .A3(\SB1_1_16/i0_0 ), .ZN(
        \SB1_1_16/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 U1172 ( .I(\SB2_0_9/buf_output[2] ), .Z(\RI5[0][152] ) );
  BUF_X4 U5228 ( .I(\SB1_1_12/buf_output[5] ), .Z(\SB2_1_12/i0_3 ) );
  NAND4_X2 \SB2_3_14/Component_Function_1/N5  ( .A1(
        \SB2_3_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_14/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_3_14/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_14/buf_output[1] ) );
  NAND3_X2 \SB1_2_0/Component_Function_3/N1  ( .A1(\SB1_2_0/i1[9] ), .A2(
        \RI1[2][191] ), .A3(\SB1_2_0/i0[6] ), .ZN(
        \SB1_2_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U6608 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0_4 ), .A3(
        \SB1_0_2/i1[9] ), .ZN(\SB1_0_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB2_4_12/Component_Function_3/N2  ( .A1(\SB2_4_12/i0_0 ), .A2(
        \SB2_4_12/i0_3 ), .A3(\SB2_4_12/i0_4 ), .ZN(
        \SB2_4_12/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB1_1_12/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[118] ), .Z(
        \SB1_1_12/i0_4 ) );
  NAND3_X2 \SB1_4_27/Component_Function_0/N3  ( .A1(\SB1_4_27/i0[10] ), .A2(
        \SB1_4_27/i0_4 ), .A3(\SB1_4_27/i0_3 ), .ZN(
        \SB1_4_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U837 ( .A1(\SB1_3_31/i0[10] ), .A2(\SB1_3_31/i1[9] ), .A3(
        \SB1_3_31/i1_7 ), .ZN(\SB1_3_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U3735 ( .A1(\SB1_1_17/i0[10] ), .A2(\SB1_1_17/i0_3 ), .A3(
        \SB1_1_17/i0_4 ), .ZN(\SB1_1_17/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 U9037 ( .I(\SB2_2_21/buf_output[2] ), .Z(\RI5[2][80] ) );
  INV_X2 \SB1_1_5/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[161] ), .ZN(
        \SB1_1_5/i1_5 ) );
  INV_X2 U1369 ( .I(\MC_ARK_ARC_1_2/buf_output[115] ), .ZN(\SB1_3_12/i1_7 ) );
  NAND3_X2 \SB2_2_10/Component_Function_1/N3  ( .A1(n589), .A2(
        \SB2_2_10/i0[6] ), .A3(\SB2_2_10/i0[9] ), .ZN(
        \SB2_2_10/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 \SB1_0_21/BUF_3_0  ( .I(\SB1_0_21/buf_output[3] ), .Z(\RI3[0][75] )
         );
  NAND3_X2 U1160 ( .A1(\SB1_1_21/i0_3 ), .A2(\SB1_1_21/i0[9] ), .A3(
        \SB1_1_21/i0[10] ), .ZN(n2801) );
  BUF_X4 \SB2_1_31/BUF_4_0  ( .I(\SB2_1_31/buf_output[4] ), .Z(\RI5[1][10] )
         );
  NAND3_X2 U2376 ( .A1(\SB1_4_12/i1_5 ), .A2(\SB1_4_12/i0_4 ), .A3(
        \SB1_4_12/i0_0 ), .ZN(n1483) );
  NAND3_X2 \SB2_0_14/Component_Function_4/N2  ( .A1(\SB2_0_14/i3[0] ), .A2(
        \SB2_0_14/i0_0 ), .A3(\SB2_0_14/i1_7 ), .ZN(
        \SB2_0_14/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 \SB2_0_11/BUF_4_0  ( .I(\SB2_0_11/buf_output[4] ), .Z(\RI5[0][130] )
         );
  BUF_X4 \SB2_0_11/BUF_5  ( .I(\RI3[0][125] ), .Z(\SB2_0_11/i0_3 ) );
  BUF_X4 \SB2_0_12/BUF_2_0  ( .I(\SB2_0_12/buf_output[2] ), .Z(\RI5[0][134] )
         );
  BUF_X4 \SB2_1_8/BUF_4  ( .I(\SB1_1_9/buf_output[4] ), .Z(\SB2_1_8/i0_4 ) );
  NAND3_X2 \SB1_3_5/Component_Function_2/N4  ( .A1(\SB1_3_5/i1_5 ), .A2(
        \SB1_3_5/i0_0 ), .A3(\SB1_3_5/i0_4 ), .ZN(
        \SB1_3_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U1189 ( .A1(\SB2_0_20/i0_3 ), .A2(\SB2_0_20/i1[9] ), .A3(
        \SB2_0_20/i0[6] ), .ZN(\SB2_0_20/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U1400 ( .I(\SB2_0_17/buf_output[3] ), .Z(\RI5[0][99] ) );
  NAND3_X2 \SB2_1_8/Component_Function_3/N2  ( .A1(\SB2_1_8/i0_0 ), .A2(
        \SB2_1_8/i0_3 ), .A3(\SB2_1_8/i0_4 ), .ZN(
        \SB2_1_8/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U4309 ( .A1(\SB2_0_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_4/NAND4_in[1] ), .A3(n1239), .A4(
        \SB2_0_5/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_5/buf_output[4] ) );
  NAND3_X2 U5931 ( .A1(\SB2_1_3/i0[10] ), .A2(\SB2_1_3/i1_5 ), .A3(
        \SB2_1_3/i1[9] ), .ZN(\SB2_1_3/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_0_31/BUF_4_0  ( .I(\SB2_0_31/buf_output[4] ), .Z(\RI5[0][10] )
         );
  NAND3_X2 U931 ( .A1(\SB2_2_15/i0[10] ), .A2(\SB2_2_15/i1_7 ), .A3(
        \SB2_2_15/i1[9] ), .ZN(n1802) );
  CLKBUF_X4 \SB2_0_19/BUF_1  ( .I(\SB1_0_23/buf_output[1] ), .Z(
        \SB2_0_19/i0[6] ) );
  NAND3_X1 U6789 ( .A1(\SB1_1_6/i0_0 ), .A2(\SB1_1_6/i0_4 ), .A3(
        \SB1_1_6/i1_5 ), .ZN(n2100) );
  BUF_X4 \SB2_4_12/BUF_1_0  ( .I(\SB2_4_12/buf_output[1] ), .Z(\RI5[4][139] )
         );
  INV_X2 \SB2_3_6/INV_4  ( .I(\SB2_3_6/i0_4 ), .ZN(\SB2_3_6/i0[7] ) );
  BUF_X4 \SB2_3_16/BUF_5  ( .I(\SB1_3_16/buf_output[5] ), .Z(\SB2_3_16/i0_3 )
         );
  NAND3_X2 U948 ( .A1(\SB2_2_31/i0_3 ), .A2(\SB2_2_31/i0_0 ), .A3(
        \SB2_2_31/i0_4 ), .ZN(\SB2_2_31/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 U85 ( .I(Key[18]), .Z(n56) );
  BUF_X4 U2053 ( .I(\SB2_0_17/buf_output[2] ), .Z(\RI5[0][104] ) );
  CLKBUF_X2 U153 ( .I(Key[12]), .Z(n95) );
  NAND4_X2 \SB2_0_31/Component_Function_1/N5  ( .A1(
        \SB2_0_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_31/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_31/buf_output[1] ) );
  INV_X4 \SB2_0_22/INV_3  ( .I(\RI3[0][57] ), .ZN(\SB2_0_22/i0[8] ) );
  BUF_X4 U1821 ( .I(\MC_ARK_ARC_1_0/buf_output[5] ), .Z(\SB1_1_31/i0_3 ) );
  BUF_X4 U9046 ( .I(\SB2_2_26/buf_output[2] ), .Z(\RI5[2][50] ) );
  NAND2_X2 U1601 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i1[9] ), .ZN(
        \SB3_1/Component_Function_1/NAND4_in[0] ) );
  INV_X1 \SB1_4_29/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[12] ), .ZN(
        \SB1_4_29/i3[0] ) );
  BUF_X2 \SB2_0_22/BUF_3  ( .I(\SB1_0_24/buf_output[3] ), .Z(\SB2_0_22/i0[10] ) );
  INV_X2 \SB1_0_24/INV_0  ( .I(n267), .ZN(\SB1_0_24/i3[0] ) );
  NAND3_X2 U590 ( .A1(\SB3_14/i0[6] ), .A2(\SB3_14/i0[9] ), .A3(\SB3_14/i0_4 ), 
        .ZN(n1628) );
  NAND3_X2 U2216 ( .A1(\SB1_2_22/i0[9] ), .A2(\SB1_2_22/i0_0 ), .A3(
        \SB1_2_22/i0[8] ), .ZN(\SB1_2_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_7/Component_Function_4/N4  ( .A1(\SB2_2_7/i1[9] ), .A2(
        \SB2_2_7/i1_5 ), .A3(\SB2_2_7/i0_4 ), .ZN(
        \SB2_2_7/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \SB2_0_31/BUF_3_0  ( .I(\SB2_0_31/buf_output[3] ), .Z(\RI5[0][15] )
         );
  BUF_X2 \SB2_0_27/BUF_4_0  ( .I(\SB2_0_27/buf_output[4] ), .Z(\RI5[0][34] )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_45  ( .I(\SB2_2_26/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[45] ) );
  NAND3_X1 \SB4_4/Component_Function_0/N3  ( .A1(\SB4_4/i0[10] ), .A2(
        \SB4_4/i0_4 ), .A3(\SB4_4/i0_3 ), .ZN(
        \SB4_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB1_0_19/Component_Function_3/N2  ( .A1(\SB1_0_19/i0_0 ), .A2(
        \SB1_0_19/i0_3 ), .A3(\SB1_0_19/i0_4 ), .ZN(
        \SB1_0_19/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U5055 ( .I(\SB2_3_29/buf_output[5] ), .Z(\RI5[3][17] ) );
  NAND3_X2 U1206 ( .A1(\SB2_0_22/i0[8] ), .A2(\SB2_0_22/i0_0 ), .A3(
        \SB2_0_22/i0[9] ), .ZN(\SB2_0_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_20/Component_Function_4/N2  ( .A1(\SB2_0_20/i3[0] ), .A2(
        \SB2_0_20/i0_0 ), .A3(\SB2_0_20/i1_7 ), .ZN(
        \SB2_0_20/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 U2154 ( .I(\MC_ARK_ARC_1_0/buf_output[112] ), .Z(\SB1_1_13/i0_4 ) );
  NAND3_X2 \SB1_0_27/Component_Function_2/N2  ( .A1(\SB1_0_27/i0_3 ), .A2(
        \SB1_0_27/i0[10] ), .A3(\SB1_0_27/i0[6] ), .ZN(
        \SB1_0_27/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB1_0_27/BUF_5  ( .I(n385), .Z(\SB1_0_27/i0_3 ) );
  CLKBUF_X4 \SB2_3_1/BUF_0  ( .I(\SB1_3_6/buf_output[0] ), .Z(\SB2_3_1/i0[9] )
         );
  BUF_X4 \SB2_0_5/BUF_4_0  ( .I(\SB2_0_5/buf_output[4] ), .Z(\RI5[0][166] ) );
  NAND3_X2 U762 ( .A1(\SB1_4_3/i0_0 ), .A2(\SB1_4_3/i0_4 ), .A3(\SB1_4_3/i1_5 ), .ZN(\SB1_4_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB1_1_16/Component_Function_2/N3  ( .A1(\SB1_1_16/i0_3 ), .A2(
        \SB1_1_16/i0[8] ), .A3(\SB1_1_16/i0[9] ), .ZN(
        \SB1_1_16/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB1_4_15/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[100] ), .Z(
        \SB1_4_15/i0_4 ) );
  NAND3_X2 \SB2_0_18/Component_Function_0/N2  ( .A1(\SB2_0_18/i0[8] ), .A2(
        \SB2_0_18/i0[7] ), .A3(\SB2_0_18/i0[6] ), .ZN(
        \SB2_0_18/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 \SB2_4_24/Component_Function_3/N1  ( .A1(n5443), .A2(
        \SB2_4_24/i0_3 ), .A3(\SB2_4_24/i0[6] ), .ZN(
        \SB2_4_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_13/Component_Function_2/N3  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i0[8] ), .A3(\SB2_3_13/i0[9] ), .ZN(
        \SB2_3_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U5197 ( .A1(\SB2_0_3/i1_5 ), .A2(\SB2_0_3/i0[10] ), .A3(
        \SB2_0_3/i1[9] ), .ZN(\SB2_0_3/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U5470 ( .I(\MC_ARK_ARC_1_1/buf_output[120] ), .ZN(\SB1_2_11/i3[0] )
         );
  NAND3_X1 U8667 ( .A1(\SB1_3_26/i0[10] ), .A2(\SB1_3_26/i1[9] ), .A3(
        \SB1_3_26/i1_7 ), .ZN(\SB1_3_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U678 ( .A1(\SB2_4_4/i0_3 ), .A2(\SB2_4_4/i1_7 ), .A3(
        \SB2_4_4/i0[8] ), .ZN(\SB2_4_4/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U847 ( .A1(\SB1_3_11/i0_3 ), .A2(\SB1_3_11/i1[9] ), .A3(
        \SB1_3_11/i0_4 ), .ZN(\SB1_3_11/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB1_3_2/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[178] ), .Z(
        \SB1_3_2/i0_4 ) );
  BUF_X4 \SB2_3_8/BUF_4  ( .I(\SB1_3_9/buf_output[4] ), .Z(\SB2_3_8/i0_4 ) );
  INV_X8 \SB1_3_4/INV_5  ( .I(\RI1[3][167] ), .ZN(\SB1_3_4/i1_5 ) );
  NAND3_X2 U978 ( .A1(\SB1_2_24/i0[6] ), .A2(\SB1_2_24/i0[9] ), .A3(
        \SB1_2_24/i0_4 ), .ZN(n2454) );
  NAND3_X2 \SB2_3_12/Component_Function_1/N2  ( .A1(\SB2_3_12/i0_3 ), .A2(
        \SB2_3_12/i1_7 ), .A3(\SB2_3_12/i0[8] ), .ZN(
        \SB2_3_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X2 U1245 ( .A1(\SB1_0_3/i0_0 ), .A2(\SB1_0_3/i3[0] ), .ZN(n1624) );
  BUF_X4 U8920 ( .I(\SB2_1_12/buf_output[2] ), .Z(\RI5[1][134] ) );
  INV_X4 \SB2_0_14/INV_1  ( .I(\SB2_0_14/i0[6] ), .ZN(\SB2_0_14/i1_7 ) );
  NAND3_X2 \SB1_2_4/Component_Function_2/N3  ( .A1(\SB1_2_4/i0_3 ), .A2(
        \SB1_2_4/i0[8] ), .A3(\SB1_2_4/i0[9] ), .ZN(
        \SB1_2_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U853 ( .A1(n3757), .A2(\SB1_3_29/i1[9] ), .A3(\SB1_3_29/i0_4 ), 
        .ZN(\SB1_3_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_25/Component_Function_2/N2  ( .A1(\SB1_1_25/i0_3 ), .A2(
        \SB1_1_25/i0[10] ), .A3(\SB1_1_25/i0[6] ), .ZN(
        \SB1_1_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB4_0/Component_Function_2/N2  ( .A1(\SB4_0/i0_3 ), .A2(
        \SB4_0/i0[10] ), .A3(\SB4_0/i0[6] ), .ZN(
        \SB4_0/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_2_3/BUF_3  ( .I(\SB1_2_5/buf_output[3] ), .Z(\SB2_2_3/i0[10] )
         );
  NAND3_X2 U5529 ( .A1(\SB1_1_25/i0_3 ), .A2(\SB1_1_25/i1[9] ), .A3(
        \SB1_1_25/i0[6] ), .ZN(\SB1_1_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_4_25/Component_Function_1/N3  ( .A1(\SB2_4_25/i1_5 ), .A2(
        \SB2_4_25/i0[6] ), .A3(\SB2_4_25/i0[9] ), .ZN(
        \SB2_4_25/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X2 U227 ( .I(Key[44]), .Z(n177) );
  NAND3_X2 U1196 ( .A1(\SB2_0_6/i0_4 ), .A2(\SB2_0_6/i0[9] ), .A3(
        \SB2_0_6/i0[6] ), .ZN(n2437) );
  INV_X2 U1908 ( .I(n390), .ZN(\SB1_0_22/i1_5 ) );
  INV_X2 U1471 ( .I(\MC_ARK_ARC_1_1/buf_output[105] ), .ZN(\SB1_2_14/i0[8] )
         );
  NAND3_X2 \SB2_0_20/Component_Function_5/N2  ( .A1(\SB2_0_20/i0_0 ), .A2(
        \SB2_0_20/i0[6] ), .A3(\SB2_0_20/i0[10] ), .ZN(
        \SB2_0_20/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB1_4_27/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[27] ), .Z(
        \SB1_4_27/i0[10] ) );
  NAND2_X2 \SB2_0_20/Component_Function_5/N1  ( .A1(\SB2_0_20/i0_0 ), .A2(
        \SB2_0_20/i3[0] ), .ZN(\SB2_0_20/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_4_23/BUF_5  ( .I(\SB1_4_23/buf_output[5] ), .Z(\SB2_4_23/i0_3 )
         );
  NAND2_X2 \SB1_4_29/Component_Function_5/N1  ( .A1(\SB1_4_29/i0_0 ), .A2(
        \SB1_4_29/i3[0] ), .ZN(\SB1_4_29/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U2038 ( .I(\SB2_1_12/buf_output[1] ), .Z(\RI5[1][139] ) );
  BUF_X4 \SB2_0_7/BUF_2_0  ( .I(\SB2_0_7/buf_output[2] ), .Z(\RI5[0][164] ) );
  BUF_X4 \SB1_0_11/BUF_5  ( .I(n401), .Z(\SB1_0_11/i0_3 ) );
  NAND3_X2 \SB2_0_31/Component_Function_5/N3  ( .A1(\SB2_0_31/i1[9] ), .A2(
        \RI3[0][4] ), .A3(\SB2_0_31/i0_3 ), .ZN(
        \SB2_0_31/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X2 U217 ( .I(Key[173]), .Z(n165) );
  INV_X2 \SB1_2_9/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[132] ), .ZN(
        \SB1_2_9/i3[0] ) );
  NAND3_X2 \SB1_2_24/Component_Function_3/N2  ( .A1(\SB1_2_24/i0_0 ), .A2(
        \SB1_2_24/i0_3 ), .A3(\SB1_2_24/i0_4 ), .ZN(
        \SB1_2_24/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB1_0_5/BUF_3  ( .I(n369), .Z(\SB1_0_5/i0[10] ) );
  INV_X2 \SB1_0_5/INV_3  ( .I(n369), .ZN(\SB1_0_5/i0[8] ) );
  BUF_X4 \SB1_3_6/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[154] ), .Z(
        \SB1_3_6/i0_4 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_107_1  ( .I(\MC_ARK_ARC_1_1/buf_output[107] ), 
        .Z(\RI1[2][107] ) );
  NAND2_X2 \SB2_1_11/Component_Function_5/N1  ( .A1(\SB2_1_11/i0_0 ), .A2(
        \SB2_1_11/i3[0] ), .ZN(\SB2_1_11/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U1663 ( .I(\SB3_27/buf_output[3] ), .ZN(\SB4_25/i0[8] ) );
  NAND3_X2 U1103 ( .A1(\SB1_1_25/i0_3 ), .A2(\SB1_1_25/i0_4 ), .A3(
        \SB1_1_25/i1[9] ), .ZN(\SB1_1_25/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_0_0/BUF_1_0  ( .I(\SB2_0_0/buf_output[1] ), .Z(\RI5[0][19] ) );
  NAND2_X2 U2440 ( .A1(\SB3_25/i0_0 ), .A2(\SB3_25/i3[0] ), .ZN(
        \SB3_25/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB1_1_11/Component_Function_5/N1  ( .A1(\SB1_1_11/i0_0 ), .A2(
        \SB1_1_11/i3[0] ), .ZN(\SB1_1_11/Component_Function_5/NAND4_in[0] ) );
  INV_X8 \SB1_4_27/INV_2  ( .I(\RI1[4][26] ), .ZN(\SB1_4_27/i1[9] ) );
  NAND3_X2 U4956 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i0[7] ), .A3(\SB3_1/i0_0 ), 
        .ZN(n2408) );
  CLKBUF_X4 \SB1_0_24/BUF_0  ( .I(n267), .Z(\SB1_0_24/i0[9] ) );
  BUF_X4 U9185 ( .I(\SB2_4_2/buf_output[1] ), .Z(\RI5[4][7] ) );
  NAND3_X2 \SB2_4_20/Component_Function_2/N1  ( .A1(\SB2_4_20/i1_5 ), .A2(
        \SB2_4_20/i0[10] ), .A3(\SB2_4_20/i1[9] ), .ZN(
        \SB2_4_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB3_25/Component_Function_5/N2  ( .A1(\SB3_25/i0_0 ), .A2(
        \SB3_25/i0[6] ), .A3(\SB3_25/i0[10] ), .ZN(
        \SB3_25/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X2 U173 ( .I(Key[85]), .Z(n116) );
  NAND3_X2 \SB1_0_22/Component_Function_2/N2  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i0[10] ), .A3(\SB1_0_22/i0[6] ), .ZN(
        \SB1_0_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_22/Component_Function_2/N1  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0[10] ), .A3(\SB1_0_22/i1[9] ), .ZN(
        \SB1_0_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_14/Component_Function_2/N2  ( .A1(\SB2_2_14/i0_3 ), .A2(
        \SB2_2_14/i0[10] ), .A3(\SB2_2_14/i0[6] ), .ZN(
        \SB2_2_14/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 U1247 ( .A1(\SB1_0_29/Component_Function_4/NAND4_in[2] ), .A2(n2320), .ZN(n2319) );
  NAND3_X2 \SB2_2_25/Component_Function_2/N3  ( .A1(\SB2_2_25/i0_3 ), .A2(
        \SB2_2_25/i0[8] ), .A3(\SB2_2_25/i0[9] ), .ZN(
        \SB2_2_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U1575 ( .A1(\SB2_0_6/i0[10] ), .A2(\SB2_0_6/i0_3 ), .A3(
        \SB2_0_6/i0[6] ), .ZN(\SB2_0_6/Component_Function_2/NAND4_in[1] ) );
  INV_X2 \SB1_2_4/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[163] ), .ZN(
        \SB1_2_4/i1_7 ) );
  INV_X2 \SB2_2_28/INV_1  ( .I(\SB1_2_0/buf_output[1] ), .ZN(\SB2_2_28/i1_7 )
         );
  BUF_X4 U1408 ( .I(\RI1[4][53] ), .Z(\SB1_4_23/i0_3 ) );
  NAND2_X2 U1265 ( .A1(\SB1_0_6/Component_Function_0/NAND4_in[0] ), .A2(n1985), 
        .ZN(n1984) );
  NAND3_X2 \SB2_3_2/Component_Function_3/N3  ( .A1(\SB2_3_2/i1[9] ), .A2(
        \SB2_3_2/i1_7 ), .A3(\SB2_3_2/i0[10] ), .ZN(
        \SB2_3_2/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 \SB2_0_5/Component_Function_1/N5  ( .A1(
        \SB2_0_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_5/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_5/buf_output[1] ) );
  NAND3_X2 \SB1_0_13/Component_Function_2/N3  ( .A1(\SB1_0_13/i0_3 ), .A2(
        n5428), .A3(\SB1_0_13/i0[9] ), .ZN(
        \SB1_0_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U7808 ( .A1(\SB2_2_18/i0_3 ), .A2(\SB2_2_18/i0[10] ), .A3(
        \SB2_2_18/i0_4 ), .ZN(\SB2_2_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_23/Component_Function_0/N2  ( .A1(\SB1_1_23/i0[8] ), .A2(
        \SB1_1_23/i0[7] ), .A3(\SB1_1_23/i0[6] ), .ZN(
        \SB1_1_23/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_14/Component_Function_5/N2  ( .A1(\SB2_1_14/i0_0 ), .A2(
        \SB2_1_14/i0[6] ), .A3(\SB2_1_14/i0[10] ), .ZN(
        \SB2_1_14/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X4 \SB2_0_1/BUF_3  ( .I(\RI3[0][183] ), .Z(\SB2_0_1/i0[10] ) );
  BUF_X2 U82 ( .I(Key[1]), .Z(n78) );
  CLKBUF_X4 U2087 ( .I(n340), .Z(\SB1_0_20/i0_4 ) );
  NAND3_X1 U170 ( .A1(\SB4_29/i0[6] ), .A2(\SB4_29/i0[9] ), .A3(
        \SB3_30/buf_output[4] ), .ZN(n2200) );
  CLKBUF_X2 U219 ( .I(Key[97]), .Z(n168) );
  NAND3_X2 \SB2_1_23/Component_Function_2/N1  ( .A1(\SB2_1_23/i1_5 ), .A2(
        \SB2_1_23/i0[10] ), .A3(\SB2_1_23/i1[9] ), .ZN(
        \SB2_1_23/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U9193 ( .I(\SB2_4_31/buf_output[0] ), .Z(\RI5[4][30] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_73  ( .I(\SB2_1_23/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[73] ) );
  BUF_X8 U1388 ( .I(\RI3[2][95] ), .Z(\SB2_2_16/i0_3 ) );
  NAND3_X2 \SB1_0_5/Component_Function_5/N2  ( .A1(\SB1_0_5/i0_0 ), .A2(
        \SB1_0_5/i0[6] ), .A3(\SB1_0_5/i0[10] ), .ZN(
        \SB1_0_5/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_0_25/BUF_5  ( .I(\RI3[0][41] ), .Z(\SB2_0_25/i0_3 ) );
  NAND3_X2 \SB1_0_25/Component_Function_2/N4  ( .A1(\SB1_0_25/i1_5 ), .A2(
        \SB1_0_25/i0_0 ), .A3(\SB1_0_25/i0_4 ), .ZN(
        \SB1_0_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_24/Component_Function_2/N1  ( .A1(\SB1_3_24/i1_5 ), .A2(
        \SB1_3_24/i0[10] ), .A3(\SB1_3_24/i1[9] ), .ZN(
        \SB1_3_24/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 U9020 ( .I(\SB2_2_14/buf_output[0] ), .Z(\RI5[2][132] ) );
  CLKBUF_X4 \SB2_0_2/BUF_3_0  ( .I(\SB2_0_2/buf_output[3] ), .Z(\RI5[0][189] )
         );
  NAND3_X1 U6748 ( .A1(\SB2_3_27/i0[8] ), .A2(\SB2_3_27/i3[0] ), .A3(
        \SB2_3_27/i1_5 ), .ZN(\SB2_3_27/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X2 U198 ( .I(Key[75]), .Z(n141) );
  NAND3_X2 \SB1_1_13/Component_Function_3/N2  ( .A1(\SB1_1_13/i0_0 ), .A2(
        \SB1_1_13/i0_3 ), .A3(\SB1_1_13/i0_4 ), .ZN(
        \SB1_1_13/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 U2086 ( .I(n305), .Z(\SB1_0_5/i0[9] ) );
  NAND3_X2 U1207 ( .A1(\SB2_0_26/i0_0 ), .A2(\SB2_0_26/i0_4 ), .A3(
        \SB2_0_26/i0_3 ), .ZN(\SB2_0_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U4328 ( .A1(\SB1_0_0/i0[10] ), .A2(\SB1_0_0/i0[9] ), .A3(
        \SB1_0_0/i0_3 ), .ZN(n1248) );
  NAND3_X2 \SB1_2_6/Component_Function_2/N1  ( .A1(\SB1_2_6/i1_5 ), .A2(
        \SB1_2_6/i0[10] ), .A3(\SB1_2_6/i1[9] ), .ZN(
        \SB1_2_6/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U8194 ( .A1(\SB1_1_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_21/Component_Function_4/NAND4_in[1] ), .ZN(n2802) );
  NAND2_X2 \SB1_2_4/Component_Function_5/N1  ( .A1(\SB1_2_4/i0_0 ), .A2(
        \SB1_2_4/i3[0] ), .ZN(\SB1_2_4/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_3_19/Component_Function_5/N1  ( .A1(\SB2_3_19/i0_0 ), .A2(
        \SB2_3_19/i3[0] ), .ZN(\SB2_3_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_31/Component_Function_3/N1  ( .A1(\SB1_1_31/i1[9] ), .A2(
        \SB1_1_31/i0_3 ), .A3(\SB1_1_31/i0[6] ), .ZN(
        \SB1_1_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_9/Component_Function_2/N1  ( .A1(\SB2_1_9/i1_5 ), .A2(
        \SB2_1_9/i0[10] ), .A3(\SB2_1_9/i1[9] ), .ZN(
        \SB2_1_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_29/Component_Function_2/N3  ( .A1(\SB1_1_29/i0_3 ), .A2(
        \SB1_1_29/i0[8] ), .A3(\SB1_1_29/i0[9] ), .ZN(
        \SB1_1_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_28/Component_Function_3/N1  ( .A1(\SB2_3_28/i1[9] ), .A2(
        \SB2_3_28/i0_3 ), .A3(\SB2_3_28/i0[6] ), .ZN(
        \SB2_3_28/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_0_29/BUF_0_0  ( .I(\SB2_0_29/buf_output[0] ), .Z(\RI5[0][42] )
         );
  NAND3_X2 U4068 ( .A1(\SB2_4_31/i0[7] ), .A2(\SB2_4_31/i0[8] ), .A3(
        \SB2_4_31/i0[6] ), .ZN(\SB2_4_31/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_4/Component_Function_3/N3  ( .A1(\SB2_2_4/i1[9] ), .A2(
        \SB2_2_4/i1_7 ), .A3(\SB2_2_4/i0[10] ), .ZN(
        \SB2_2_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB1_0_9/Component_Function_2/N3  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i0[8] ), .A3(\SB1_0_9/i0[9] ), .ZN(
        \SB1_0_9/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_41_1  ( .I(\MC_ARK_ARC_1_3/buf_output[41] ), .Z(
        \RI1[4][41] ) );
  CLKBUF_X4 \SB2_4_9/BUF_0  ( .I(\SB1_4_14/buf_output[0] ), .Z(\SB2_4_9/i0[9] ) );
  CLKBUF_X4 \SB2_0_11/BUF_2  ( .I(\RI3[0][122] ), .Z(\SB2_0_11/i0_0 ) );
  BUF_X4 \SB1_1_13/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[110] ), .Z(
        \SB1_1_13/i0_0 ) );
  NAND3_X2 U5430 ( .A1(\SB1_0_2/i1_5 ), .A2(\SB1_0_2/i0[8] ), .A3(
        \SB1_0_2/i3[0] ), .ZN(\SB1_0_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB2_1_29/Component_Function_2/N1  ( .A1(\SB2_1_29/i1_5 ), .A2(
        \SB2_1_29/i0[10] ), .A3(\SB2_1_29/i1[9] ), .ZN(
        \SB2_1_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_16/Component_Function_3/N1  ( .A1(\SB2_3_16/i1[9] ), .A2(
        \SB2_3_16/i0_3 ), .A3(\SB2_3_16/i0[6] ), .ZN(
        \SB2_3_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_4_0/Component_Function_1/N4  ( .A1(\SB2_4_0/i1_7 ), .A2(
        \SB2_4_0/i0[8] ), .A3(\SB2_4_0/i0_4 ), .ZN(
        \SB2_4_0/Component_Function_1/NAND4_in[3] ) );
  INV_X4 U1919 ( .I(n4734), .ZN(\SB2_2_31/i1_5 ) );
  NAND3_X2 \SB2_3_16/Component_Function_2/N1  ( .A1(n571), .A2(
        \SB2_3_16/i0[10] ), .A3(\SB2_3_16/i1[9] ), .ZN(
        \SB2_3_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_16/Component_Function_1/N3  ( .A1(n571), .A2(
        \SB2_3_16/i0[6] ), .A3(\SB2_3_16/i0[9] ), .ZN(
        \SB2_3_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U1226 ( .A1(\SB2_0_5/i0[10] ), .A2(\SB2_0_5/i1[9] ), .A3(
        \SB2_0_5/i1_7 ), .ZN(\SB2_0_5/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_7  ( .I(\SB2_1_2/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[7] ) );
  NAND3_X2 \SB1_3_12/Component_Function_4/N2  ( .A1(\SB1_3_12/i3[0] ), .A2(
        \SB1_3_12/i0_0 ), .A3(\SB1_3_12/i1_7 ), .ZN(
        \SB1_3_12/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 U1391 ( .I(\SB1_2_16/buf_output[5] ), .Z(\RI3[2][95] ) );
  NAND3_X2 \SB2_3_2/Component_Function_2/N1  ( .A1(\SB2_3_2/i1_5 ), .A2(
        \SB2_3_2/i0[10] ), .A3(\SB2_3_2/i1[9] ), .ZN(
        \SB2_3_2/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_3_7/BUF_5  ( .I(\SB1_3_7/buf_output[5] ), .Z(\SB2_3_7/i0_3 ) );
  CLKBUF_X4 \SB2_4_1/BUF_2  ( .I(\SB1_4_4/buf_output[2] ), .Z(\SB2_4_1/i0_0 )
         );
  INV_X4 \SB1_4_25/INV_5  ( .I(\RI1[4][41] ), .ZN(\SB1_4_25/i1_5 ) );
  BUF_X4 \SB2_0_20/BUF_2  ( .I(\RI3[0][68] ), .Z(\SB2_0_20/i0_0 ) );
  NAND3_X2 U8090 ( .A1(\SB2_1_8/i0_4 ), .A2(\SB2_1_8/i0[9] ), .A3(
        \SB2_1_8/i0[6] ), .ZN(\SB2_1_8/Component_Function_5/NAND4_in[3] ) );
  BUF_X2 U19 ( .I(Key[147]), .Z(n206) );
  BUF_X2 U609 ( .I(Key[62]), .Z(n182) );
  NAND3_X2 U2256 ( .A1(\SB2_2_5/i0_3 ), .A2(\SB2_2_5/i1[9] ), .A3(
        \SB2_2_5/i0_4 ), .ZN(n3031) );
  CLKBUF_X2 U4968 ( .I(Key[43]), .Z(n214) );
  CLKBUF_X2 U124 ( .I(Key[102]), .Z(n54) );
  CLKBUF_X4 \SB1_0_17/BUF_4  ( .I(n346), .Z(\SB1_0_17/i0_4 ) );
  INV_X1 U2278 ( .I(n28), .ZN(n457) );
  INV_X1 U289 ( .I(n101), .ZN(n431) );
  BUF_X2 \SB1_0_8/BUF_4  ( .I(n364), .Z(\SB1_0_8/i0_4 ) );
  CLKBUF_X4 \SB1_0_10/BUF_2  ( .I(n296), .Z(\SB1_0_10/i0_0 ) );
  INV_X1 U56 ( .I(n62), .ZN(n465) );
  CLKBUF_X4 \SB1_0_0/BUF_2  ( .I(n316), .Z(\SB1_0_0/i0_0 ) );
  INV_X1 U30 ( .I(n23), .ZN(n440) );
  CLKBUF_X4 U2088 ( .I(n329), .Z(\SB1_0_25/i0[10] ) );
  CLKBUF_X4 \SB1_0_23/BUF_4  ( .I(n334), .Z(\SB1_0_23/i0_4 ) );
  INV_X1 U37 ( .I(n55), .ZN(n462) );
  CLKBUF_X4 \SB1_0_29/BUF_1  ( .I(n223), .Z(\SB1_0_29/i0[6] ) );
  INV_X1 U34 ( .I(n81), .ZN(n477) );
  CLKBUF_X4 \SB1_0_21/BUF_4  ( .I(n338), .Z(\SB1_0_21/i0_4 ) );
  INV_X1 U55 ( .I(n66), .ZN(n546) );
  CLKBUF_X4 \SB1_0_29/BUF_3  ( .I(n321), .Z(\SB1_0_29/i0[10] ) );
  INV_X1 U40 ( .I(n7), .ZN(n540) );
  CLKBUF_X4 U2074 ( .I(n343), .Z(\SB1_0_18/i0[10] ) );
  CLKBUF_X4 \SB1_0_4/BUF_2  ( .I(n308), .Z(\SB1_0_4/i0_0 ) );
  CLKBUF_X4 \SB1_0_6/BUF_4  ( .I(n368), .Z(\SB1_0_6/i0_4 ) );
  NAND2_X1 U8041 ( .A1(\SB1_0_14/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_14/Component_Function_0/NAND4_in[1] ), .ZN(n2693) );
  CLKBUF_X4 U5274 ( .I(\SB1_0_16/buf_output[3] ), .Z(\SB2_0_14/i0[10] ) );
  CLKBUF_X4 \SB1_0_8/BUF_4_0  ( .I(\SB1_0_8/buf_output[4] ), .Z(\RI3[0][148] )
         );
  BUF_X2 \SB2_0_7/BUF_0  ( .I(\RI3[0][144] ), .Z(\SB2_0_7/i0[9] ) );
  CLKBUF_X4 \SB2_0_26/BUF_1  ( .I(\SB1_0_30/buf_output[1] ), .Z(
        \SB2_0_26/i0[6] ) );
  CLKBUF_X4 U2060 ( .I(\RI3[0][21] ), .Z(\SB2_0_28/i0[10] ) );
  CLKBUF_X4 \SB2_0_9/BUF_5  ( .I(\SB1_0_9/buf_output[5] ), .Z(\SB2_0_9/i0_3 )
         );
  CLKBUF_X4 \SB2_0_1/BUF_4  ( .I(\RI3[0][184] ), .Z(\SB2_0_1/i0_4 ) );
  CLKBUF_X4 \SB2_0_27/BUF_1  ( .I(\SB1_0_31/buf_output[1] ), .Z(
        \SB2_0_27/i0[6] ) );
  CLKBUF_X4 \SB2_0_21/BUF_0  ( .I(\RI3[0][60] ), .Z(\SB2_0_21/i0[9] ) );
  BUF_X2 \SB2_0_8/BUF_1  ( .I(\RI3[0][139] ), .Z(\SB2_0_8/i0[6] ) );
  CLKBUF_X4 \SB2_0_18/BUF_0  ( .I(\RI3[0][78] ), .Z(\SB2_0_18/i0[9] ) );
  CLKBUF_X4 U2118 ( .I(\RI3[0][115] ), .Z(\SB2_0_12/i0[6] ) );
  CLKBUF_X4 \SB2_0_24/BUF_2  ( .I(\RI3[0][44] ), .Z(\SB2_0_24/i0_0 ) );
  CLKBUF_X4 U5289 ( .I(\RI3[0][117] ), .Z(\SB2_0_12/i0[10] ) );
  CLKBUF_X4 \SB1_0_24/BUF_4_0  ( .I(\SB1_0_24/buf_output[4] ), .Z(\RI3[0][52] ) );
  CLKBUF_X4 \SB2_0_25/BUF_1  ( .I(\SB1_0_29/buf_output[1] ), .Z(
        \SB2_0_25/i0[6] ) );
  CLKBUF_X8 \SB2_0_20/BUF_5  ( .I(\RI3[0][71] ), .Z(\SB2_0_20/i0_3 ) );
  CLKBUF_X4 \SB2_0_19/BUF_0  ( .I(\RI3[0][72] ), .Z(\SB2_0_19/i0[9] ) );
  CLKBUF_X4 \SB2_0_13/BUF_3_0  ( .I(\SB2_0_13/buf_output[3] ), .Z(
        \RI5[0][123] ) );
  BUF_X4 \SB2_0_3/BUF_3_0  ( .I(\SB2_0_3/buf_output[3] ), .Z(\RI5[0][183] ) );
  BUF_X4 \SB2_0_15/BUF_0_0  ( .I(\SB2_0_15/buf_output[0] ), .Z(\RI5[0][126] )
         );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_67  ( .I(\SB2_0_24/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[67] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_0/BUF_77  ( .I(\SB2_0_19/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[77] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_0/BUF_35  ( .I(\SB2_0_26/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[35] ) );
  CLKBUF_X4 \SB2_0_1/BUF_5_0  ( .I(\SB2_0_1/buf_output[5] ), .Z(\RI5[0][185] )
         );
  CLKBUF_X4 \SB2_0_27/BUF_3_0  ( .I(\SB2_0_27/buf_output[3] ), .Z(\RI5[0][39] ) );
  BUF_X4 \SB2_0_14/BUF_4_0  ( .I(\SB2_0_14/buf_output[4] ), .Z(\RI5[0][112] )
         );
  CLKBUF_X4 \SB1_1_6/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[154] ), .Z(
        \SB1_1_6/i0_4 ) );
  CLKBUF_X4 \SB1_1_30/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[7] ), .Z(
        \SB1_1_30/i0[6] ) );
  CLKBUF_X4 \SB1_1_28/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[18] ), .Z(
        \SB1_1_28/i0[9] ) );
  CLKBUF_X4 \SB1_1_20/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[70] ), .Z(
        \SB1_1_20/i0_4 ) );
  CLKBUF_X4 U2153 ( .I(\MC_ARK_ARC_1_0/buf_output[68] ), .Z(\SB1_1_20/i0_0 )
         );
  CLKBUF_X4 \SB1_1_20/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[67] ), .Z(
        \SB1_1_20/i0[6] ) );
  CLKBUF_X4 \SB1_1_27/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[28] ), .Z(
        \SB1_1_27/i0_4 ) );
  CLKBUF_X4 \SB1_1_4/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[162] ), .Z(
        \SB1_1_4/i0[9] ) );
  CLKBUF_X4 \SB1_1_1/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[181] ), .Z(
        \SB1_1_1/i0[6] ) );
  CLKBUF_X4 U1343 ( .I(\MC_ARK_ARC_1_0/buf_output[75] ), .Z(\SB1_1_19/i0[10] )
         );
  CLKBUF_X4 \SB1_1_18/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[78] ), .Z(
        \SB1_1_18/i0[9] ) );
  CLKBUF_X4 \SB1_1_20/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[69] ), .Z(
        \SB1_1_20/i0[10] ) );
  CLKBUF_X4 \SB1_1_5/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[160] ), .Z(
        \SB1_1_5/i0_4 ) );
  CLKBUF_X4 \SB1_1_24/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[46] ), .Z(
        \SB1_1_24/i0_4 ) );
  CLKBUF_X4 \SB1_1_25/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[39] ), .Z(
        \SB1_1_25/i0[10] ) );
  CLKBUF_X4 \SB2_1_13/BUF_3  ( .I(\RI3[1][111] ), .Z(\SB2_1_13/i0[10] ) );
  CLKBUF_X4 \SB2_1_24/BUF_3  ( .I(\SB1_1_26/buf_output[3] ), .Z(
        \SB2_1_24/i0[10] ) );
  CLKBUF_X4 \SB2_1_23/BUF_1  ( .I(\SB1_1_27/buf_output[1] ), .Z(
        \SB2_1_23/i0[6] ) );
  CLKBUF_X4 \SB2_1_3/BUF_1  ( .I(\SB1_1_7/buf_output[1] ), .Z(\SB2_1_3/i0[6] )
         );
  CLKBUF_X4 \SB2_1_19/BUF_1  ( .I(\SB1_1_23/buf_output[1] ), .Z(
        \SB2_1_19/i0[6] ) );
  CLKBUF_X4 \SB2_1_14/BUF_3  ( .I(\SB1_1_16/buf_output[3] ), .Z(
        \SB2_1_14/i0[10] ) );
  CLKBUF_X4 \SB2_1_13/BUF_0  ( .I(\SB1_1_18/buf_output[0] ), .Z(
        \SB2_1_13/i0[9] ) );
  CLKBUF_X4 \SB2_1_13/BUF_1  ( .I(\SB1_1_17/buf_output[1] ), .Z(
        \SB2_1_13/i0[6] ) );
  CLKBUF_X4 \SB2_1_4/BUF_2  ( .I(\SB1_1_7/buf_output[2] ), .Z(\SB2_1_4/i0_0 )
         );
  CLKBUF_X4 \SB2_1_2/BUF_3  ( .I(\SB1_1_4/buf_output[3] ), .Z(\SB2_1_2/i0[10] ) );
  CLKBUF_X4 \SB2_1_8/BUF_3  ( .I(\SB1_1_10/buf_output[3] ), .Z(
        \SB2_1_8/i0[10] ) );
  CLKBUF_X4 \SB2_1_8/BUF_0  ( .I(\SB1_1_13/buf_output[0] ), .Z(\SB2_1_8/i0[9] ) );
  CLKBUF_X4 \SB2_1_12/BUF_0  ( .I(\SB1_1_17/buf_output[0] ), .Z(
        \SB2_1_12/i0[9] ) );
  CLKBUF_X4 \SB2_1_17/BUF_2  ( .I(\SB1_1_20/buf_output[2] ), .Z(
        \SB2_1_17/i0_0 ) );
  CLKBUF_X4 \SB2_1_22/BUF_3  ( .I(\SB1_1_24/buf_output[3] ), .Z(
        \SB2_1_22/i0[10] ) );
  CLKBUF_X4 \SB2_1_25/BUF_0  ( .I(\SB1_1_30/buf_output[0] ), .Z(
        \SB2_1_25/i0[9] ) );
  CLKBUF_X4 \SB2_1_31/BUF_0  ( .I(\SB1_1_4/buf_output[0] ), .Z(
        \SB2_1_31/i0[9] ) );
  CLKBUF_X4 U7815 ( .I(\SB2_1_28/buf_output[1] ), .Z(\RI5[1][43] ) );
  CLKBUF_X4 \SB2_1_5/BUF_0_0  ( .I(\SB2_1_5/buf_output[0] ), .Z(\RI5[1][186] )
         );
  BUF_X4 U2037 ( .I(\SB2_1_7/buf_output[1] ), .Z(\RI5[1][169] ) );
  CLKBUF_X4 \SB1_2_6/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[152] ), .Z(
        \SB1_2_6/i0_0 ) );
  CLKBUF_X4 \SB1_2_25/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[37] ), .Z(
        \SB1_2_25/i0[6] ) );
  CLKBUF_X4 U5371 ( .I(\MC_ARK_ARC_1_1/buf_output[111] ), .Z(\SB1_2_13/i0[10] ) );
  CLKBUF_X4 \SB1_2_19/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[76] ), .Z(
        \SB1_2_19/i0_4 ) );
  CLKBUF_X4 \SB1_2_19/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[73] ), .Z(
        \SB1_2_19/i0[6] ) );
  CLKBUF_X4 \SB1_2_19/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[75] ), .Z(
        \SB1_2_19/i0[10] ) );
  CLKBUF_X4 \SB1_2_2/BUF_2  ( .I(n6279), .Z(\SB1_2_2/i0_0 ) );
  CLKBUF_X4 U1287 ( .I(\MC_ARK_ARC_1_1/buf_output[68] ), .Z(\SB1_2_20/i0_0 )
         );
  CLKBUF_X4 \SB1_2_12/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[115] ), .Z(
        \SB1_2_12/i0[6] ) );
  CLKBUF_X4 \SB1_2_25/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[40] ), .Z(
        \SB1_2_25/i0_4 ) );
  CLKBUF_X4 \SB1_2_4/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[163] ), .Z(
        \SB1_2_4/i0[6] ) );
  CLKBUF_X4 U5447 ( .I(\MC_ARK_ARC_1_1/buf_output[13] ), .Z(\SB1_2_29/i0[6] )
         );
  CLKBUF_X4 \SB1_2_29/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[12] ), .Z(
        \SB1_2_29/i0[9] ) );
  CLKBUF_X4 \SB1_2_8/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[142] ), .Z(
        \SB1_2_8/i0_4 ) );
  CLKBUF_X4 \SB2_2_11/BUF_3  ( .I(\SB1_2_13/buf_output[3] ), .Z(
        \SB2_2_11/i0[10] ) );
  CLKBUF_X4 \SB2_2_6/BUF_3  ( .I(\SB1_2_8/buf_output[3] ), .Z(\SB2_2_6/i0[10] ) );
  CLKBUF_X4 \SB2_2_15/BUF_4  ( .I(\SB1_2_16/buf_output[4] ), .Z(
        \SB2_2_15/i0_4 ) );
  CLKBUF_X4 \SB2_2_15/BUF_2  ( .I(\SB1_2_18/buf_output[2] ), .Z(
        \SB2_2_15/i0_0 ) );
  CLKBUF_X4 \SB2_2_1/BUF_2  ( .I(\SB1_2_4/buf_output[2] ), .Z(\SB2_2_1/i0_0 )
         );
  CLKBUF_X4 \SB2_2_4/BUF_1  ( .I(\SB1_2_8/buf_output[1] ), .Z(\SB2_2_4/i0[6] )
         );
  CLKBUF_X4 \SB2_2_30/BUF_3  ( .I(\SB1_2_0/buf_output[3] ), .Z(
        \SB2_2_30/i0[10] ) );
  CLKBUF_X4 \SB2_2_16/BUF_0  ( .I(\SB1_2_21/buf_output[0] ), .Z(
        \SB2_2_16/i0[9] ) );
  CLKBUF_X4 \SB2_2_29/BUF_4  ( .I(\SB1_2_30/buf_output[4] ), .Z(
        \SB2_2_29/i0_4 ) );
  CLKBUF_X4 \SB2_2_27/BUF_2  ( .I(\SB1_2_30/buf_output[2] ), .Z(
        \SB2_2_27/i0_0 ) );
  CLKBUF_X4 \SB2_2_21/BUF_0  ( .I(\SB1_2_26/buf_output[0] ), .Z(
        \SB2_2_21/i0[9] ) );
  CLKBUF_X4 \SB2_2_19/BUF_0  ( .I(\SB1_2_24/buf_output[0] ), .Z(
        \SB2_2_19/i0[9] ) );
  CLKBUF_X4 \SB2_2_20/BUF_2  ( .I(\SB1_2_23/buf_output[2] ), .Z(
        \SB2_2_20/i0_0 ) );
  CLKBUF_X4 \SB2_2_20/BUF_1  ( .I(\SB1_2_24/buf_output[1] ), .Z(
        \SB2_2_20/i0[6] ) );
  CLKBUF_X4 \SB2_2_3/BUF_1  ( .I(\SB1_2_7/buf_output[1] ), .Z(\SB2_2_3/i0[6] )
         );
  CLKBUF_X4 \SB2_2_31/BUF_2  ( .I(\SB1_2_2/buf_output[2] ), .Z(\SB2_2_31/i0_0 ) );
  CLKBUF_X4 \SB2_2_4/BUF_3  ( .I(\SB1_2_6/buf_output[3] ), .Z(\SB2_2_4/i0[10] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_133  ( .I(\SB2_2_13/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[133] ) );
  CLKBUF_X4 U2013 ( .I(\SB2_2_24/buf_output[5] ), .Z(\RI5[2][47] ) );
  CLKBUF_X4 U5252 ( .I(\SB2_2_27/buf_output[0] ), .Z(\RI5[2][54] ) );
  CLKBUF_X4 \SB1_3_16/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[94] ), .Z(
        \SB1_3_16/i0_4 ) );
  CLKBUF_X4 \SB1_3_7/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[144] ), .Z(
        \SB1_3_7/i0[9] ) );
  CLKBUF_X4 \SB1_3_15/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[96] ), .Z(
        \SB1_3_15/i0[9] ) );
  CLKBUF_X4 \SB1_3_26/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[34] ), .Z(
        \SB1_3_26/i0_4 ) );
  CLKBUF_X4 \SB1_3_22/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[54] ), .Z(
        \SB1_3_22/i0[9] ) );
  CLKBUF_X4 \SB1_3_22/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[57] ), .Z(
        \SB1_3_22/i0[10] ) );
  CLKBUF_X4 U1356 ( .I(\MC_ARK_ARC_1_2/buf_output[66] ), .Z(\SB1_3_20/i0[9] )
         );
  CLKBUF_X4 \SB1_3_8/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[140] ), .Z(
        \SB1_3_8/i0_0 ) );
  BUF_X4 \SB1_3_6/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[155] ), .Z(
        \SB1_3_6/i0_3 ) );
  CLKBUF_X4 \SB1_3_8/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[142] ), .Z(
        \SB1_3_8/i0_4 ) );
  CLKBUF_X4 \SB1_3_6/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[151] ), .Z(
        \SB1_3_6/i0[6] ) );
  CLKBUF_X4 U1586 ( .I(\MC_ARK_ARC_1_2/buf_output[45] ), .Z(\SB1_3_24/i0[10] )
         );
  CLKBUF_X4 \SB1_3_14/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[105] ), .Z(
        \SB1_3_14/i0[10] ) );
  CLKBUF_X4 \SB2_3_1/BUF_4  ( .I(\SB1_3_2/buf_output[4] ), .Z(\SB2_3_1/i0_4 )
         );
  CLKBUF_X4 \SB2_3_21/BUF_2  ( .I(\SB1_3_24/buf_output[2] ), .Z(
        \SB2_3_21/i0_0 ) );
  CLKBUF_X4 \SB2_3_7/BUF_3  ( .I(\SB1_3_9/buf_output[3] ), .Z(\SB2_3_7/i0[10] ) );
  CLKBUF_X4 U2316 ( .I(\SB1_3_1/buf_output[2] ), .Z(\SB2_3_30/i0_0 ) );
  CLKBUF_X4 \SB2_3_0/BUF_4  ( .I(\SB1_3_1/buf_output[4] ), .Z(\SB2_3_0/i0_4 )
         );
  CLKBUF_X4 \SB2_3_15/BUF_2  ( .I(\SB1_3_18/buf_output[2] ), .Z(
        \SB2_3_15/i0_0 ) );
  CLKBUF_X4 \SB2_3_11/BUF_3  ( .I(\SB1_3_13/buf_output[3] ), .Z(
        \SB2_3_11/i0[10] ) );
  CLKBUF_X4 U2318 ( .I(\SB1_3_19/buf_output[4] ), .Z(\SB2_3_18/i0_4 ) );
  CLKBUF_X4 \SB2_3_22/BUF_2  ( .I(\SB1_3_25/buf_output[2] ), .Z(
        \SB2_3_22/i0_0 ) );
  CLKBUF_X4 U5310 ( .I(\SB1_3_24/buf_output[3] ), .Z(\SB2_3_22/i0[10] ) );
  CLKBUF_X4 U2323 ( .I(\SB1_3_21/buf_output[1] ), .Z(\SB2_3_17/i0[6] ) );
  CLKBUF_X4 U5102 ( .I(\SB1_3_21/buf_output[2] ), .Z(\SB2_3_18/i0_0 ) );
  CLKBUF_X4 U2320 ( .I(\SB1_3_20/buf_output[2] ), .Z(\SB2_3_17/i0_0 ) );
  CLKBUF_X4 U2317 ( .I(\SB1_3_19/buf_output[1] ), .Z(\SB2_3_15/i0[6] ) );
  CLKBUF_X4 \SB2_3_20/BUF_1  ( .I(\SB1_3_24/buf_output[1] ), .Z(
        \SB2_3_20/i0[6] ) );
  CLKBUF_X4 \SB2_3_15/BUF_0  ( .I(\SB1_3_20/buf_output[0] ), .Z(
        \SB2_3_15/i0[9] ) );
  NAND3_X2 U8481 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i0[9] ), .A3(
        \SB2_3_16/i0[10] ), .ZN(\SB2_3_16/Component_Function_4/NAND4_in[2] )
         );
  CLKBUF_X4 \SB2_3_0/BUF_1  ( .I(\SB1_3_4/buf_output[1] ), .Z(\SB2_3_0/i0[6] )
         );
  CLKBUF_X4 U1994 ( .I(\SB2_3_18/buf_output[5] ), .Z(\RI5[3][83] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_3/BUF_24  ( .I(\SB2_3_0/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[24] ) );
  CLKBUF_X4 \SB1_4_22/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[55] ), .Z(
        \SB1_4_22/i0[6] ) );
  CLKBUF_X4 \SB1_4_13/BUF_2  ( .I(\MC_ARK_ARC_1_3/buf_output[110] ), .Z(
        \SB1_4_13/i0_0 ) );
  CLKBUF_X4 \SB1_4_14/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[106] ), .Z(
        \SB1_4_14/i0_4 ) );
  CLKBUF_X4 U3838 ( .I(\MC_ARK_ARC_1_3/buf_output[133] ), .Z(\SB1_4_9/i0[6] )
         );
  CLKBUF_X4 U4987 ( .I(\MC_ARK_ARC_1_3/buf_output[172] ), .Z(\SB1_4_3/i0_4 )
         );
  CLKBUF_X4 \SB1_4_17/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[88] ), .Z(
        \SB1_4_17/i0_4 ) );
  CLKBUF_X4 U1578 ( .I(\MC_ARK_ARC_1_3/buf_output[165] ), .Z(\SB1_4_4/i0[10] )
         );
  CLKBUF_X4 U1733 ( .I(\MC_ARK_ARC_1_3/buf_output[164] ), .Z(\SB1_4_4/i0_0 )
         );
  CLKBUF_X4 U788 ( .I(\MC_ARK_ARC_1_3/buf_output[0] ), .Z(\SB1_4_31/i0[9] ) );
  CLKBUF_X4 U1979 ( .I(\SB1_4_17/buf_output[3] ), .Z(\SB2_4_15/i0[10] ) );
  CLKBUF_X4 \SB2_4_30/BUF_1  ( .I(\SB1_4_2/buf_output[1] ), .Z(
        \SB2_4_30/i0[6] ) );
  CLKBUF_X4 \SB2_4_17/BUF_4  ( .I(\SB1_4_18/buf_output[4] ), .Z(
        \SB2_4_17/i0_4 ) );
  CLKBUF_X4 \SB2_4_0/BUF_3  ( .I(\SB1_4_2/buf_output[3] ), .Z(\SB2_4_0/i0[10] ) );
  CLKBUF_X4 \SB2_4_0/BUF_4  ( .I(\SB1_4_1/buf_output[4] ), .Z(\SB2_4_0/i0_4 )
         );
  CLKBUF_X4 \SB2_4_13/BUF_4  ( .I(\SB1_4_14/buf_output[4] ), .Z(
        \SB2_4_13/i0_4 ) );
  CLKBUF_X4 \MC_ARK_ARC_1_4/BUF_141  ( .I(\SB2_4_10/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[141] ) );
  BUF_X4 U1956 ( .I(\SB2_4_22/buf_output[1] ), .Z(\RI5[4][79] ) );
  BUF_X2 \SB3_7/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[144] ), .Z(
        \SB3_7/i0[9] ) );
  CLKBUF_X4 U1812 ( .I(\MC_ARK_ARC_1_4/buf_output[26] ), .Z(\SB3_27/i0_0 ) );
  CLKBUF_X4 \SB3_11/BUF_1  ( .I(\MC_ARK_ARC_1_4/buf_output[121] ), .Z(
        \SB3_11/i0[6] ) );
  CLKBUF_X4 U2429 ( .I(\MC_ARK_ARC_1_4/buf_output[70] ), .Z(\SB3_20/i0_4 ) );
  CLKBUF_X4 U1377 ( .I(\MC_ARK_ARC_1_4/buf_output[182] ), .Z(\SB3_1/i0_0 ) );
  CLKBUF_X4 \SB3_24/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[42] ), .Z(
        \SB3_24/i0[9] ) );
  CLKBUF_X4 \SB4_17/BUF_4  ( .I(\SB3_18/buf_output[4] ), .Z(\SB4_17/i0_4 ) );
  CLKBUF_X4 U1662 ( .I(\SB3_27/buf_output[3] ), .Z(\SB4_25/i0[10] ) );
  BUF_X4 \SB2_2_6/BUF_2  ( .I(\SB1_2_9/buf_output[2] ), .Z(\SB2_2_6/i0_0 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_149_1  ( .I(\MC_ARK_ARC_1_1/buf_output[149] ), 
        .Z(\RI1[2][149] ) );
  BUF_X4 U9195 ( .I(\SB2_4_5/buf_output[0] ), .Z(\RI5[4][186] ) );
  INV_X2 \SB1_3_9/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[132] ), .ZN(
        \SB1_3_9/i3[0] ) );
  INV_X1 \SB1_0_20/INV_0  ( .I(n275), .ZN(\SB1_0_20/i3[0] ) );
  BUF_X2 \SB1_0_21/BUF_1  ( .I(n231), .Z(\SB1_0_21/i0[6] ) );
  NAND3_X1 U2081 ( .A1(\SB1_0_19/i0[8] ), .A2(\SB1_0_19/i0[7] ), .A3(n233), 
        .ZN(\SB1_0_19/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_18/Component_Function_1/N4  ( .A1(\SB1_0_18/i1_7 ), .A2(
        \SB1_0_18/i0[8] ), .A3(\SB1_0_18/i0_4 ), .ZN(
        \SB1_0_18/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_18/Component_Function_1/N1  ( .A1(\SB1_0_18/i0_3 ), .A2(
        \SB1_0_18/i1[9] ), .ZN(\SB1_0_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1273 ( .A1(\SB1_0_12/i0[10] ), .A2(\SB1_0_12/i1[9] ), .A3(
        \SB1_0_12/i1_5 ), .ZN(n1836) );
  NAND3_X1 U3203 ( .A1(\SB1_0_12/i0[10] ), .A2(\SB1_0_12/i0_3 ), .A3(
        \SB1_0_12/i0[6] ), .ZN(n835) );
  BUF_X2 \SB1_0_7/BUF_3  ( .I(n365), .Z(\SB1_0_7/i0[10] ) );
  INV_X1 \SB1_0_31/INV_5  ( .I(n381), .ZN(\SB1_0_31/i1_5 ) );
  INV_X1 \SB1_0_23/INV_1  ( .I(n229), .ZN(\SB1_0_23/i1_7 ) );
  BUF_X2 \SB1_0_21/BUF_0  ( .I(n273), .Z(\SB1_0_21/i0[9] ) );
  INV_X1 \SB1_0_17/INV_4  ( .I(\SB1_0_17/i0_4 ), .ZN(\SB1_0_17/i0[7] ) );
  NAND3_X1 \SB1_0_7/Component_Function_4/N4  ( .A1(\SB1_0_7/i1[9] ), .A2(
        \SB1_0_7/i1_5 ), .A3(\SB1_0_7/i0_4 ), .ZN(
        \SB1_0_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_1/N4  ( .A1(\SB1_0_10/i1_7 ), .A2(
        \SB1_0_10/i0[8] ), .A3(\SB1_0_10/i0_4 ), .ZN(
        \SB1_0_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4966 ( .A1(\SB1_0_30/i0_3 ), .A2(\SB1_0_30/i0[8] ), .A3(
        \SB1_0_30/i0[9] ), .ZN(\SB1_0_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_3/Component_Function_0/N4  ( .A1(\SB1_0_3/i0[7] ), .A2(
        \SB1_0_3/i0_3 ), .A3(\SB1_0_3/i0_0 ), .ZN(
        \SB1_0_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_5/N3  ( .A1(\SB1_0_7/i1[9] ), .A2(
        \SB1_0_7/i0_4 ), .A3(\SB1_0_7/i0_3 ), .ZN(
        \SB1_0_7/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_14/Component_Function_3/N4  ( .A1(\SB1_0_14/i1_5 ), .A2(
        \SB1_0_14/i0[8] ), .A3(\SB1_0_14/i3[0] ), .ZN(
        \SB1_0_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_18/Component_Function_2/N3  ( .A1(\SB1_0_18/i0_3 ), .A2(
        \SB1_0_18/i0[8] ), .A3(\SB1_0_18/i0[9] ), .ZN(
        \SB1_0_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_1/Component_Function_3/N4  ( .A1(\SB1_0_1/i1_5 ), .A2(
        \SB1_0_1/i0[8] ), .A3(\SB1_0_1/i3[0] ), .ZN(
        \SB1_0_1/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_7/Component_Function_5/N1  ( .A1(\SB1_0_7/i0_0 ), .A2(
        \SB1_0_7/i3[0] ), .ZN(\SB1_0_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_1/N4  ( .A1(\SB1_0_31/i1_7 ), .A2(
        \SB1_0_31/i0[8] ), .A3(\SB1_0_31/i0_4 ), .ZN(
        \SB1_0_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_1/N2  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i1_7 ), .A3(\SB1_0_31/i0[8] ), .ZN(
        \SB1_0_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_29/Component_Function_0/N1  ( .A1(\SB1_0_29/i0[10] ), .A2(
        \SB1_0_29/i0[9] ), .ZN(\SB1_0_29/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_22/Component_Function_5/N1  ( .A1(\SB1_0_22/i0_0 ), .A2(
        \SB1_0_22/i3[0] ), .ZN(\SB1_0_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_3/N3  ( .A1(\SB1_0_6/i1[9] ), .A2(
        \SB1_0_6/i1_7 ), .A3(\SB1_0_6/i0[10] ), .ZN(
        \SB1_0_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2067 ( .A1(n230), .A2(\SB1_0_22/i0[9] ), .A3(n336), .ZN(n2400) );
  NAND2_X1 U4125 ( .A1(n1460), .A2(n2922), .ZN(n1170) );
  NAND3_X1 \SB1_0_10/Component_Function_0/N4  ( .A1(\SB1_0_10/i0[7] ), .A2(
        \SB1_0_10/i0_3 ), .A3(\SB1_0_10/i0_0 ), .ZN(
        \SB1_0_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_3/N2  ( .A1(\SB1_0_9/i0_0 ), .A2(
        \SB1_0_9/i0_3 ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U5473 ( .A1(\SB1_0_0/i0_0 ), .A2(\SB1_0_0/i0_3 ), .A3(
        \SB1_0_0/i0_4 ), .ZN(n1512) );
  NAND3_X1 U6022 ( .A1(\SB1_0_6/i0[10] ), .A2(\SB1_0_6/i0_3 ), .A3(
        \SB1_0_6/i0[6] ), .ZN(n1749) );
  NAND3_X1 \SB1_0_8/Component_Function_5/N2  ( .A1(\SB1_0_8/i0_0 ), .A2(
        \SB1_0_8/i0[6] ), .A3(\SB1_0_8/i0[10] ), .ZN(
        \SB1_0_8/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U7135 ( .A1(\SB1_0_14/i0[6] ), .A2(n352), .A3(\SB1_0_14/i0[9] ), 
        .ZN(n2483) );
  NAND3_X1 \SB1_0_30/Component_Function_5/N2  ( .A1(\SB1_0_30/i0_0 ), .A2(
        \SB1_0_30/i0[6] ), .A3(\SB1_0_30/i0[10] ), .ZN(
        \SB1_0_30/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U7188 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i1[9] ), .A3(
        \SB1_0_29/i0[6] ), .ZN(\SB1_0_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_0/N4  ( .A1(\SB1_0_5/i0[7] ), .A2(
        \SB1_0_5/i0_3 ), .A3(\SB1_0_5/i0_0 ), .ZN(
        \SB1_0_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_5/N3  ( .A1(\SB1_0_31/i1[9] ), .A2(
        \SB1_0_31/i0_4 ), .A3(\SB1_0_31/i0_3 ), .ZN(
        \SB1_0_31/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_8/Component_Function_1/N1  ( .A1(\SB1_0_8/i0_3 ), .A2(
        \SB1_0_8/i1[9] ), .ZN(\SB1_0_8/Component_Function_1/NAND4_in[0] ) );
  INV_X2 U1204 ( .I(\SB2_0_9/i3[0] ), .ZN(\SB2_0_9/i0[9] ) );
  INV_X1 U2117 ( .I(\SB1_0_26/buf_output[1] ), .ZN(\SB2_0_22/i1_7 ) );
  BUF_X2 \SB2_0_3/BUF_1  ( .I(\RI3[0][169] ), .Z(\SB2_0_3/i0[6] ) );
  INV_X1 U3029 ( .I(\RI3[0][120] ), .ZN(\SB2_0_11/i3[0] ) );
  INV_X4 \SB2_0_16/INV_3  ( .I(\RI3[0][93] ), .ZN(\SB2_0_16/i0[8] ) );
  BUF_X2 \SB2_0_13/BUF_1  ( .I(\RI3[0][109] ), .Z(\SB2_0_13/i0[6] ) );
  INV_X4 \SB2_0_26/INV_3  ( .I(\RI3[0][33] ), .ZN(\SB2_0_26/i0[8] ) );
  INV_X2 U7859 ( .I(n2611), .ZN(\SB2_0_26/i0_4 ) );
  INV_X1 \SB2_0_25/INV_1  ( .I(\SB1_0_29/buf_output[1] ), .ZN(\SB2_0_25/i1_7 )
         );
  INV_X1 \SB2_0_2/INV_4  ( .I(\SB1_0_3/buf_output[4] ), .ZN(\SB2_0_2/i0[7] )
         );
  NAND3_X1 \SB2_0_3/Component_Function_5/N3  ( .A1(\SB2_0_3/i1[9] ), .A2(
        \RI3[0][172] ), .A3(\SB2_0_3/i0_3 ), .ZN(
        \SB2_0_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_2/Component_Function_4/N3  ( .A1(\SB2_0_2/i0[9] ), .A2(
        \SB2_0_2/i0[10] ), .A3(\SB2_0_2/i0_3 ), .ZN(
        \SB2_0_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_30/Component_Function_4/N2  ( .A1(\SB2_0_30/i3[0] ), .A2(
        \SB2_0_30/i0_0 ), .A3(\SB2_0_30/i1_7 ), .ZN(
        \SB2_0_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_4/Component_Function_4/N2  ( .A1(n630), .A2(\SB2_0_4/i0_0 ), 
        .A3(\SB2_0_4/i1_7 ), .ZN(\SB2_0_4/Component_Function_4/NAND4_in[1] )
         );
  NAND3_X1 U4651 ( .A1(\SB2_0_4/i1[9] ), .A2(\RI3[0][166] ), .A3(
        \SB2_0_4/i1_5 ), .ZN(n1381) );
  NAND3_X1 U1219 ( .A1(\SB2_0_10/i0_3 ), .A2(\RI3[0][126] ), .A3(
        \SB2_0_10/i0[8] ), .ZN(\SB2_0_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_9/Component_Function_3/N4  ( .A1(\SB2_0_9/i1_5 ), .A2(
        \SB2_0_9/i0[8] ), .A3(n4847), .ZN(
        \SB2_0_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_26/Component_Function_0/N4  ( .A1(n3510), .A2(
        \SB2_0_26/i0_3 ), .A3(\SB2_0_26/i0_0 ), .ZN(
        \SB2_0_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_11/Component_Function_4/N4  ( .A1(\SB2_0_11/i1[9] ), .A2(
        \SB2_0_11/i1_5 ), .A3(\SB2_0_11/i0_4 ), .ZN(
        \SB2_0_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U5786 ( .A1(n2965), .A2(\RI3[0][128] ), .A3(\SB2_0_10/i0_3 ), .ZN(
        n1651) );
  NAND2_X1 \SB2_0_11/Component_Function_5/N1  ( .A1(\SB2_0_11/i0_0 ), .A2(
        \SB2_0_11/i3[0] ), .ZN(\SB2_0_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U6798 ( .A1(\SB2_0_3/i0_0 ), .A2(\SB2_0_3/i0[7] ), .A3(
        \SB2_0_3/i0_3 ), .ZN(\SB2_0_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1186 ( .A1(\SB2_0_11/i0[6] ), .A2(\SB2_0_11/i0_4 ), .A3(
        \SB2_0_11/i0[9] ), .ZN(n1854) );
  NAND3_X1 \SB2_0_17/Component_Function_0/N3  ( .A1(\SB2_0_17/i0[10] ), .A2(
        \RI3[0][88] ), .A3(\SB2_0_17/i0_3 ), .ZN(
        \SB2_0_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_13/Component_Function_4/N4  ( .A1(\SB2_0_13/i1[9] ), .A2(
        \SB2_0_13/i1_5 ), .A3(\RI3[0][112] ), .ZN(
        \SB2_0_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3702 ( .A1(\SB2_0_30/i0_4 ), .A2(\SB2_0_30/i1_5 ), .A3(
        \SB2_0_30/i0_0 ), .ZN(\SB2_0_30/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_12/Component_Function_0/N3  ( .A1(\SB2_0_12/i0[10] ), .A2(
        \RI3[0][118] ), .A3(\RI3[0][119] ), .ZN(
        \SB2_0_12/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 U5866 ( .A1(\RI3[0][57] ), .A2(n593), .ZN(
        \SB2_0_22/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_1/Component_Function_5/N1  ( .A1(\SB2_0_1/i0_0 ), .A2(n2592), 
        .ZN(\SB2_0_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_1/N2  ( .A1(\SB2_0_1/i0_3 ), .A2(
        \SB2_0_1/i1_7 ), .A3(\SB2_0_1/i0[8] ), .ZN(
        \SB2_0_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U5288 ( .A1(\SB2_0_12/i0[9] ), .A2(\SB2_0_12/i0[10] ), .A3(
        \RI3[0][119] ), .ZN(\SB2_0_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U5612 ( .A1(\SB2_0_30/i0_3 ), .A2(\SB2_0_30/i0_0 ), .A3(
        \SB2_0_30/i0[7] ), .ZN(n1568) );
  NAND3_X1 U2717 ( .A1(\SB2_0_28/i0_0 ), .A2(\SB2_0_28/i1_5 ), .A3(
        \SB2_0_28/i0_4 ), .ZN(\SB2_0_28/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4870 ( .A1(\SB2_0_23/i0_0 ), .A2(\SB2_0_23/i3[0] ), .A3(
        \SB2_0_23/i1_7 ), .ZN(\SB2_0_23/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_23/Component_Function_5/N1  ( .A1(\SB2_0_23/i0_0 ), .A2(
        \SB2_0_23/i3[0] ), .ZN(\SB2_0_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_3/Component_Function_3/N1  ( .A1(\SB2_0_3/i1[9] ), .A2(
        \SB2_0_3/i0_3 ), .A3(\SB2_0_3/i0[6] ), .ZN(
        \SB2_0_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1183 ( .A1(\SB2_0_31/i0_3 ), .A2(\SB2_0_31/i0[9] ), .A3(
        \SB2_0_31/i0[8] ), .ZN(\SB2_0_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_20/Component_Function_1/N3  ( .A1(\SB2_0_20/i1_5 ), .A2(
        \SB2_0_20/i0[6] ), .A3(n5264), .ZN(
        \SB2_0_20/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_22/Component_Function_0/N1  ( .A1(\SB2_0_22/i0[10] ), .A2(
        \SB2_0_22/i0[9] ), .ZN(\SB2_0_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_21/Component_Function_0/N2  ( .A1(\SB2_0_21/i0[8] ), .A2(
        \SB2_0_21/i0[7] ), .A3(\SB2_0_21/i0[6] ), .ZN(
        \SB2_0_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_23/Component_Function_4/N4  ( .A1(\SB2_0_23/i1[9] ), .A2(
        \SB2_0_23/i1_5 ), .A3(\SB1_0_24/buf_output[4] ), .ZN(
        \SB2_0_23/Component_Function_4/NAND4_in[3] ) );
  BUF_X2 U191 ( .I(Key[130]), .Z(n134) );
  INV_X1 U44 ( .I(n40), .ZN(n517) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_43  ( .I(\SB2_0_28/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[43] ) );
  INV_X1 U2420 ( .I(n76), .ZN(n450) );
  BUF_X2 \SB2_0_29/BUF_1_0  ( .I(\SB2_0_29/buf_output[1] ), .Z(\RI5[0][37] )
         );
  INV_X1 U385 ( .I(Key[145]), .ZN(n452) );
  BUF_X2 \SB1_1_5/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[157] ), .Z(
        \SB1_1_5/i0[6] ) );
  INV_X1 \SB1_1_1/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[181] ), .ZN(
        \SB1_1_1/i1_7 ) );
  INV_X1 \SB1_1_24/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[42] ), .ZN(
        \SB1_1_24/i3[0] ) );
  INV_X1 \SB1_1_2/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[175] ), .ZN(
        \SB1_1_2/i1_7 ) );
  INV_X1 \SB1_1_28/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[18] ), .ZN(
        \SB1_1_28/i3[0] ) );
  INV_X1 \SB1_1_19/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[72] ), .ZN(
        \SB1_1_19/i3[0] ) );
  INV_X1 \SB1_1_7/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[144] ), .ZN(
        \SB1_1_7/i3[0] ) );
  INV_X1 \SB1_1_22/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[54] ), .ZN(
        \SB1_1_22/i3[0] ) );
  BUF_X2 \SB1_1_25/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[36] ), .Z(
        \SB1_1_25/i0[9] ) );
  INV_X1 \SB1_1_28/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[19] ), .ZN(
        \SB1_1_28/i1_7 ) );
  INV_X1 \SB1_1_23/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[49] ), .ZN(
        \SB1_1_23/i1_7 ) );
  BUF_X2 \SB1_1_17/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[85] ), .Z(
        \SB1_1_17/i0[6] ) );
  BUF_X2 \SB1_1_26/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[30] ), .Z(
        \SB1_1_26/i0[9] ) );
  BUF_X2 \SB1_1_31/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[3] ), .Z(
        \SB1_1_31/i0[10] ) );
  INV_X1 \SB1_1_20/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[67] ), .ZN(
        \SB1_1_20/i1_7 ) );
  BUF_X2 \SB1_1_8/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[139] ), .Z(
        \SB1_1_8/i0[6] ) );
  NAND3_X1 \SB1_1_19/Component_Function_4/N3  ( .A1(\SB1_1_19/i0[9] ), .A2(
        \SB1_1_19/i0[10] ), .A3(\SB1_1_19/i0_3 ), .ZN(
        \SB1_1_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_3/Component_Function_0/N3  ( .A1(\SB1_1_3/i0[10] ), .A2(
        \SB1_1_3/i0_4 ), .A3(\SB1_1_3/i0_3 ), .ZN(
        \SB1_1_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_27/Component_Function_1/N3  ( .A1(\SB1_1_27/i1_5 ), .A2(
        \SB1_1_27/i0[6] ), .A3(\SB1_1_27/i0[9] ), .ZN(
        \SB1_1_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1140 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i0_0 ), .A3(
        \SB1_1_7/i0[7] ), .ZN(n2989) );
  NAND3_X1 \SB1_1_9/Component_Function_0/N4  ( .A1(\SB1_1_9/i0[7] ), .A2(
        \SB1_1_9/i0_3 ), .A3(\SB1_1_9/i0_0 ), .ZN(
        \SB1_1_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U7542 ( .A1(\SB1_1_18/i0_0 ), .A2(\SB1_1_18/i3[0] ), .A3(
        \SB1_1_18/i1_7 ), .ZN(\SB1_1_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_10/Component_Function_1/N2  ( .A1(\SB1_1_10/i0_3 ), .A2(
        \SB1_1_10/i1_7 ), .A3(\SB1_1_10/i0[8] ), .ZN(
        \SB1_1_10/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_18/Component_Function_4/N3  ( .A1(\SB1_1_18/i0[9] ), .A2(
        \SB1_1_18/i0[10] ), .A3(\SB1_1_18/i0_3 ), .ZN(
        \SB1_1_18/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U2164 ( .A1(\SB1_1_8/i0_3 ), .A2(\SB1_1_8/i1[9] ), .ZN(
        \SB1_1_8/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_7/Component_Function_0/N1  ( .A1(\SB1_1_7/i0[10] ), .A2(
        \SB1_1_7/i0[9] ), .ZN(\SB1_1_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_2/N2  ( .A1(\SB1_1_15/i0_3 ), .A2(
        \SB1_1_15/i0[10] ), .A3(\SB1_1_15/i0[6] ), .ZN(
        \SB1_1_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U7737 ( .A1(\SB1_1_16/i0[9] ), .A2(\SB1_1_16/i0[6] ), .A3(
        \SB1_1_16/i1_5 ), .ZN(\SB1_1_16/Component_Function_1/NAND4_in[2] ) );
  INV_X2 \SB1_1_16/INV_4  ( .I(\SB1_1_16/i0_4 ), .ZN(\SB1_1_16/i0[7] ) );
  NAND3_X1 \SB1_1_10/Component_Function_3/N2  ( .A1(\SB1_1_10/i0_0 ), .A2(
        \SB1_1_10/i0_3 ), .A3(\SB1_1_10/i0_4 ), .ZN(
        \SB1_1_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U6292 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0_0 ), .A3(
        \SB1_1_22/i0_4 ), .ZN(n1863) );
  NAND3_X1 \SB1_1_12/Component_Function_0/N4  ( .A1(\SB1_1_12/i0[7] ), .A2(
        \SB1_1_12/i0_3 ), .A3(\SB1_1_12/i0_0 ), .ZN(
        \SB1_1_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1121 ( .A1(\SB1_1_3/i0[9] ), .A2(\SB1_1_3/i0[6] ), .A3(
        \SB1_1_3/i1_5 ), .ZN(n1662) );
  NAND3_X1 \SB1_1_19/Component_Function_1/N4  ( .A1(\SB1_1_19/i1_7 ), .A2(
        \SB1_1_19/i0[8] ), .A3(\SB1_1_19/i0_4 ), .ZN(
        \SB1_1_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_19/Component_Function_0/N4  ( .A1(\SB1_1_19/i0[7] ), .A2(
        \SB1_1_19/i0_3 ), .A3(\SB1_1_19/i0_0 ), .ZN(
        \SB1_1_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3761 ( .A1(\SB1_1_8/i0[7] ), .A2(\SB1_1_8/i0[8] ), .A3(
        \SB1_1_8/i0[6] ), .ZN(\SB1_1_8/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_5/Component_Function_4/N4  ( .A1(\SB1_1_5/i1[9] ), .A2(
        \SB1_1_5/i1_5 ), .A3(\SB1_1_5/i0_4 ), .ZN(
        \SB1_1_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1144 ( .A1(\SB1_1_18/i0[10] ), .A2(\SB1_1_18/i1[9] ), .A3(
        \SB1_1_18/i1_7 ), .ZN(n2834) );
  NAND3_X1 U2162 ( .A1(\SB1_1_16/i1[9] ), .A2(\SB1_1_16/i1_5 ), .A3(
        \SB1_1_16/i0_4 ), .ZN(\SB1_1_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_29/Component_Function_1/N3  ( .A1(\SB1_1_29/i1_5 ), .A2(
        \SB1_1_29/i0[6] ), .A3(\SB1_1_29/i0[9] ), .ZN(
        \SB1_1_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_26/Component_Function_1/N3  ( .A1(\SB1_1_26/i1_5 ), .A2(
        \SB1_1_26/i0[6] ), .A3(\SB1_1_26/i0[9] ), .ZN(
        \SB1_1_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_19/Component_Function_1/N3  ( .A1(\SB1_1_19/i1_5 ), .A2(
        \SB1_1_19/i0[6] ), .A3(\SB1_1_19/i0[9] ), .ZN(
        \SB1_1_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_23/Component_Function_1/N3  ( .A1(\SB1_1_23/i1_5 ), .A2(
        \SB1_1_23/i0[6] ), .A3(\SB1_1_23/i0[9] ), .ZN(
        \SB1_1_23/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_29/Component_Function_1/N1  ( .A1(\SB1_1_29/i0_3 ), .A2(
        \SB1_1_29/i1[9] ), .ZN(\SB1_1_29/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_27/Component_Function_0/N1  ( .A1(\SB1_1_27/i0[10] ), .A2(
        \SB1_1_27/i0[9] ), .ZN(\SB1_1_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_1/Component_Function_0/N4  ( .A1(\SB1_1_1/i0[7] ), .A2(
        \SB1_1_1/i0_3 ), .A3(\SB1_1_1/i0_0 ), .ZN(
        \SB1_1_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_0/Component_Function_5/N4  ( .A1(\SB1_1_0/i0[9] ), .A2(
        \SB1_1_0/i0[6] ), .A3(\MC_ARK_ARC_1_0/buf_output[190] ), .ZN(
        \SB1_1_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2693 ( .A1(\SB1_1_19/i0_0 ), .A2(\SB1_1_19/i0[10] ), .A3(
        \SB1_1_19/i0[6] ), .ZN(\SB1_1_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_12/Component_Function_0/N3  ( .A1(\SB1_1_12/i0[10] ), .A2(
        \SB1_1_12/i0_4 ), .A3(\SB1_1_12/i0_3 ), .ZN(
        \SB1_1_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_28/Component_Function_3/N1  ( .A1(\SB1_1_28/i1[9] ), .A2(
        \SB1_1_28/i0_3 ), .A3(\SB1_1_28/i0[6] ), .ZN(
        \SB1_1_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_0/N2  ( .A1(\SB1_1_13/i0[8] ), .A2(
        \SB1_1_13/i0[7] ), .A3(\SB1_1_13/i0[6] ), .ZN(
        \SB1_1_13/Component_Function_0/NAND4_in[1] ) );
  INV_X1 \SB2_1_5/INV_0  ( .I(\SB1_1_10/buf_output[0] ), .ZN(\SB2_1_5/i3[0] )
         );
  INV_X1 \SB2_1_25/INV_1  ( .I(\SB1_1_29/buf_output[1] ), .ZN(\SB2_1_25/i1_7 )
         );
  NAND2_X1 \SB2_1_17/Component_Function_1/N1  ( .A1(\SB2_1_17/i0_3 ), .A2(
        \SB2_1_17/i1[9] ), .ZN(\SB2_1_17/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_5/Component_Function_5/N1  ( .A1(\SB2_1_5/i0_0 ), .A2(
        \SB2_1_5/i3[0] ), .ZN(\SB2_1_5/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_7/Component_Function_5/N1  ( .A1(\SB2_1_7/i0_0 ), .A2(
        \SB2_1_7/i3[0] ), .ZN(\SB2_1_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_2/N4  ( .A1(\SB2_1_5/i1_5 ), .A2(
        \SB2_1_5/i0_0 ), .A3(\SB2_1_5/i0_4 ), .ZN(
        \SB2_1_5/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_5/Component_Function_0/N1  ( .A1(\SB2_1_5/i0[10] ), .A2(
        \SB2_1_5/i0[9] ), .ZN(\SB2_1_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_1/Component_Function_1/N3  ( .A1(\SB2_1_1/i1_5 ), .A2(
        \SB2_1_1/i0[6] ), .A3(\SB2_1_1/i0[9] ), .ZN(
        \SB2_1_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_4/Component_Function_1/N3  ( .A1(\SB2_1_4/i1_5 ), .A2(
        \SB1_1_8/buf_output[1] ), .A3(\SB2_1_4/i0[9] ), .ZN(
        \SB2_1_4/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_10/Component_Function_5/N1  ( .A1(\SB2_1_10/i0_0 ), .A2(
        \SB2_1_10/i3[0] ), .ZN(\SB2_1_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_21/Component_Function_4/N2  ( .A1(\SB2_1_21/i3[0] ), .A2(
        \SB2_1_21/i0_0 ), .A3(\SB2_1_21/i1_7 ), .ZN(
        \SB2_1_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N2  ( .A1(\SB2_1_26/i3[0] ), .A2(
        \SB2_1_26/i0_0 ), .A3(\SB2_1_26/i1_7 ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1067 ( .A1(\SB2_1_24/i0_4 ), .A2(\SB2_1_24/i1_7 ), .A3(
        \SB2_1_24/i0[8] ), .ZN(n1936) );
  NAND3_X1 U4236 ( .A1(\SB2_1_16/i0[10] ), .A2(\SB2_1_16/i1_7 ), .A3(
        \SB2_1_16/i1[9] ), .ZN(n1212) );
  NAND3_X1 U7945 ( .A1(\SB2_1_16/i0[9] ), .A2(\SB2_1_16/i1_5 ), .A3(
        \SB2_1_16/i0[6] ), .ZN(\SB2_1_16/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_2/Component_Function_1/N1  ( .A1(\SB2_1_2/i0_3 ), .A2(
        \SB2_1_2/i1[9] ), .ZN(\SB2_1_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U4093 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB2_1_18/i0[10] ), .A3(
        \SB2_1_18/i0[9] ), .ZN(\SB2_1_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_31/Component_Function_0/N3  ( .A1(\SB2_1_31/i0[10] ), .A2(
        n5429), .A3(\SB2_1_31/i0_3 ), .ZN(
        \SB2_1_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_25/Component_Function_0/N4  ( .A1(\SB2_1_25/i0[7] ), .A2(
        \SB2_1_25/i0_3 ), .A3(\SB2_1_25/i0_0 ), .ZN(
        \SB2_1_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_12/Component_Function_4/N4  ( .A1(\SB2_1_12/i1[9] ), .A2(
        \SB2_1_12/i1_5 ), .A3(\SB2_1_12/i0_4 ), .ZN(
        \SB2_1_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1073 ( .A1(\SB2_1_17/i0_3 ), .A2(\SB2_1_17/i0[10] ), .A3(
        \SB2_1_17/i0[9] ), .ZN(n969) );
  NAND3_X1 \SB2_1_25/Component_Function_2/N2  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB1_1_27/buf_output[3] ), .A3(\SB2_1_25/i0[6] ), .ZN(
        \SB2_1_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_25/Component_Function_4/N3  ( .A1(\SB2_1_25/i0[9] ), .A2(
        \SB1_1_27/buf_output[3] ), .A3(\SB2_1_25/i0_3 ), .ZN(
        \SB2_1_25/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_31/Component_Function_0/N1  ( .A1(\SB2_1_31/i0[10] ), .A2(
        \SB2_1_31/i0[9] ), .ZN(\SB2_1_31/Component_Function_0/NAND4_in[0] ) );
  BUF_X2 \SB1_2_24/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[42] ), .Z(
        \SB1_2_24/i0[9] ) );
  BUF_X2 \SB1_2_19/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[72] ), .Z(
        \SB1_2_19/i0[9] ) );
  BUF_X2 \SB1_2_30/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[6] ), .Z(
        \SB1_2_30/i0[9] ) );
  INV_X1 \SB1_2_10/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[126] ), .ZN(
        \SB1_2_10/i3[0] ) );
  BUF_X2 \SB1_2_25/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[36] ), .Z(
        \SB1_2_25/i0[9] ) );
  INV_X1 \SB1_2_20/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[67] ), .ZN(
        \SB1_2_20/i1_7 ) );
  INV_X1 \SB1_2_6/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[151] ), .ZN(
        \SB1_2_6/i1_7 ) );
  NAND3_X1 \SB1_2_17/Component_Function_3/N1  ( .A1(\SB1_2_17/i1[9] ), .A2(
        \SB1_2_17/i0_3 ), .A3(\SB1_2_17/i0[6] ), .ZN(
        \SB1_2_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U7543 ( .A1(\SB1_2_2/i0[10] ), .A2(\SB1_2_2/i0[9] ), .A3(
        \SB1_2_2/i0_3 ), .ZN(n2445) );
  NAND3_X1 \SB1_2_2/Component_Function_4/N4  ( .A1(\SB1_2_2/i1[9] ), .A2(
        \SB1_2_2/i1_5 ), .A3(\SB1_2_2/i0_4 ), .ZN(
        \SB1_2_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_4/N2  ( .A1(\SB1_2_2/i3[0] ), .A2(
        \SB1_2_2/i0_0 ), .A3(\SB1_2_2/i1_7 ), .ZN(
        \SB1_2_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_9/Component_Function_0/N4  ( .A1(\SB1_2_9/i0[7] ), .A2(
        \SB1_2_9/i0_3 ), .A3(\SB1_2_9/i0_0 ), .ZN(
        \SB1_2_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2229 ( .A1(\SB1_2_8/i1_7 ), .A2(\SB1_2_8/i0[8] ), .A3(
        \SB1_2_8/i0_4 ), .ZN(\SB1_2_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_20/Component_Function_4/N4  ( .A1(\SB1_2_20/i1[9] ), .A2(
        \SB1_2_20/i1_5 ), .A3(\SB1_2_20/i0_4 ), .ZN(
        \SB1_2_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1015 ( .A1(\SB1_2_5/i0_0 ), .A2(\SB1_2_5/i1_7 ), .A3(
        \SB1_2_5/i3[0] ), .ZN(n840) );
  NAND3_X1 U1702 ( .A1(\SB1_2_15/i1[9] ), .A2(\RI1[2][101] ), .A3(
        \SB1_2_15/i0[6] ), .ZN(\SB1_2_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1652 ( .A1(\SB1_2_22/i1_5 ), .A2(\SB1_2_22/i0_4 ), .A3(
        \SB1_2_22/i1[9] ), .ZN(n2604) );
  NAND3_X1 \SB1_2_4/Component_Function_4/N4  ( .A1(\SB1_2_4/i1[9] ), .A2(
        \SB1_2_4/i1_5 ), .A3(\SB1_2_4/i0_4 ), .ZN(
        \SB1_2_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_6/Component_Function_3/N2  ( .A1(\SB1_2_6/i0_0 ), .A2(
        \SB1_2_6/i0_3 ), .A3(\SB1_2_6/i0_4 ), .ZN(
        \SB1_2_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_20/Component_Function_0/N3  ( .A1(\SB1_2_20/i0[10] ), .A2(
        \SB1_2_20/i0_4 ), .A3(\SB1_2_20/i0_3 ), .ZN(
        \SB1_2_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_6/Component_Function_4/N3  ( .A1(\SB1_2_6/i0[9] ), .A2(
        \SB1_2_6/i0[10] ), .A3(\SB1_2_6/i0_3 ), .ZN(
        \SB1_2_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_1/Component_Function_4/N4  ( .A1(\SB1_2_1/i1[9] ), .A2(
        \SB1_2_1/i1_5 ), .A3(\SB1_2_1/i0_4 ), .ZN(
        \SB1_2_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_27/Component_Function_3/N1  ( .A1(\SB1_2_27/i1[9] ), .A2(
        \SB1_2_27/i0_3 ), .A3(\SB1_2_27/i0[6] ), .ZN(
        \SB1_2_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_29/Component_Function_1/N3  ( .A1(\SB1_2_29/i1_5 ), .A2(
        \SB1_2_29/i0[6] ), .A3(\SB1_2_29/i0[9] ), .ZN(
        \SB1_2_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_25/Component_Function_3/N2  ( .A1(\SB1_2_25/i0_0 ), .A2(
        \SB1_2_25/i0_3 ), .A3(\SB1_2_25/i0_4 ), .ZN(
        \SB1_2_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_26/Component_Function_4/N4  ( .A1(\SB1_2_26/i1[9] ), .A2(
        \SB1_2_26/i1_5 ), .A3(\SB1_2_26/i0_4 ), .ZN(
        \SB1_2_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2223 ( .A1(\SB1_2_30/i1[9] ), .A2(\SB1_2_30/i1_5 ), .A3(
        \SB1_2_30/i0_4 ), .ZN(\SB1_2_30/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_25/Component_Function_1/N1  ( .A1(\SB1_2_25/i0_3 ), .A2(
        \SB1_2_25/i1[9] ), .ZN(\SB1_2_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1009 ( .A1(\SB1_2_14/i0[10] ), .A2(\SB1_2_14/i1[9] ), .A3(
        \SB1_2_14/i1_7 ), .ZN(n3005) );
  NAND3_X1 \SB1_2_21/Component_Function_0/N4  ( .A1(\SB1_2_21/i0[7] ), .A2(
        \SB1_2_21/i0_3 ), .A3(\SB1_2_21/i0_0 ), .ZN(
        \SB1_2_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_29/Component_Function_0/N2  ( .A1(\SB1_2_29/i0[8] ), .A2(
        \SB1_2_29/i0[7] ), .A3(\SB1_2_29/i0[6] ), .ZN(
        \SB1_2_29/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_0/Component_Function_1/N2  ( .A1(\RI1[2][191] ), .A2(
        \SB1_2_0/i1_7 ), .A3(\SB1_2_0/i0[8] ), .ZN(
        \SB1_2_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_12/Component_Function_4/N2  ( .A1(\SB1_2_12/i3[0] ), .A2(
        \RI1[2][116] ), .A3(\SB1_2_12/i1_7 ), .ZN(
        \SB1_2_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_0/Component_Function_0/N4  ( .A1(\SB1_2_0/i0[7] ), .A2(
        \RI1[2][191] ), .A3(\SB1_2_0/i0_0 ), .ZN(
        \SB1_2_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1668 ( .A1(\SB1_2_30/i0_4 ), .A2(\SB1_2_30/i1_7 ), .A3(
        \SB1_2_30/i0[8] ), .ZN(\SB1_2_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_20/Component_Function_1/N3  ( .A1(\SB1_2_20/i1_5 ), .A2(
        \SB1_2_20/i0[6] ), .A3(\SB1_2_20/i0[9] ), .ZN(
        \SB1_2_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U5767 ( .A1(\SB1_2_24/i0[10] ), .A2(\SB1_2_24/i1[9] ), .A3(
        \SB1_2_24/i1_5 ), .ZN(n1637) );
  NAND3_X1 \SB1_2_3/Component_Function_4/N1  ( .A1(\SB1_2_3/i0[9] ), .A2(
        \SB1_2_3/i0_0 ), .A3(\SB1_2_3/i0[8] ), .ZN(
        \SB1_2_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U989 ( .A1(\SB1_2_10/i0[9] ), .A2(\SB1_2_10/i0[8] ), .A3(
        \SB1_2_10/i0_3 ), .ZN(n958) );
  NAND3_X1 U5682 ( .A1(\SB1_2_31/i0[8] ), .A2(\SB1_2_31/i0_3 ), .A3(
        \SB1_2_31/i1_7 ), .ZN(\SB1_2_31/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_19/Component_Function_2/N2  ( .A1(\SB1_2_19/i0_3 ), .A2(
        \SB1_2_19/i0[10] ), .A3(\SB1_2_19/i0[6] ), .ZN(
        \SB1_2_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1000 ( .A1(\SB1_2_6/i0[8] ), .A2(\SB1_2_6/i0_4 ), .A3(
        \SB1_2_6/i1_7 ), .ZN(n944) );
  NAND2_X1 \SB1_2_31/Component_Function_1/N1  ( .A1(\SB1_2_31/i0_3 ), .A2(
        \SB1_2_31/i1[9] ), .ZN(\SB1_2_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_2/N2  ( .A1(\SB1_2_9/i0_3 ), .A2(
        \SB1_2_9/i0[10] ), .A3(\SB1_2_9/i0[6] ), .ZN(
        \SB1_2_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_21/Component_Function_0/N3  ( .A1(\SB1_2_21/i0[10] ), .A2(
        \SB1_2_21/i0_4 ), .A3(\SB1_2_21/i0_3 ), .ZN(
        \SB1_2_21/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 U7026 ( .A1(\SB1_2_29/i1_5 ), .A2(n2210), .ZN(
        \SB1_2_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_4/Component_Function_2/N1  ( .A1(\SB1_2_4/i1_5 ), .A2(
        \SB1_2_4/i0[10] ), .A3(\SB1_2_4/i1[9] ), .ZN(
        \SB1_2_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U6911 ( .A1(\SB1_2_20/i0_4 ), .A2(\SB1_2_20/i0_3 ), .A3(
        \SB1_2_20/i1[9] ), .ZN(\SB1_2_20/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1018 ( .A1(\SB1_2_6/i0[9] ), .A2(\SB1_2_6/i0_4 ), .A3(
        \SB1_2_6/i0[6] ), .ZN(\SB1_2_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_11/Component_Function_1/N3  ( .A1(\SB1_2_11/i1_5 ), .A2(
        \SB1_2_11/i0[6] ), .A3(\MC_ARK_ARC_1_1/buf_output[120] ), .ZN(
        \SB1_2_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_9/Component_Function_3/N2  ( .A1(\SB1_2_9/i0_0 ), .A2(
        \SB1_2_9/i0_3 ), .A3(\SB1_2_9/i0_4 ), .ZN(
        \SB1_2_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_25/Component_Function_4/N3  ( .A1(\SB1_2_25/i0[9] ), .A2(
        \SB1_2_25/i0[10] ), .A3(\SB1_2_25/i0_3 ), .ZN(
        \SB1_2_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_21/Component_Function_0/N2  ( .A1(\SB1_2_21/i0[8] ), .A2(
        \SB1_2_21/i0[7] ), .A3(\SB1_2_21/i0[6] ), .ZN(
        \SB1_2_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U4757 ( .A1(n6291), .A2(\SB1_2_28/i1[9] ), .A3(\SB1_2_28/i0_4 ), 
        .ZN(n1420) );
  NAND3_X1 U1017 ( .A1(n3839), .A2(\SB1_2_29/i1[9] ), .A3(\SB1_2_29/i0[10] ), 
        .ZN(\SB1_2_29/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U2021 ( .I(\SB2_2_23/i0_4 ), .Z(n600) );
  NAND2_X1 \SB2_2_3/Component_Function_5/N1  ( .A1(\SB2_2_3/i0_0 ), .A2(
        \SB2_2_3/i3[0] ), .ZN(\SB2_2_3/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_29/Component_Function_5/N1  ( .A1(\SB2_2_29/i0_0 ), .A2(
        \SB2_2_29/i3[0] ), .ZN(\SB2_2_29/Component_Function_5/NAND4_in[0] ) );
  INV_X1 \SB2_2_17/INV_1  ( .I(\SB1_2_21/buf_output[1] ), .ZN(\SB2_2_17/i1_7 )
         );
  INV_X1 \SB2_2_11/INV_1  ( .I(\RI3[2][121] ), .ZN(\SB2_2_11/i1_7 ) );
  NAND3_X1 U6800 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0[8] ), .A3(
        \SB2_2_29/i0[9] ), .ZN(n2105) );
  NAND3_X1 \SB2_2_27/Component_Function_4/N2  ( .A1(\SB2_2_27/i3[0] ), .A2(
        \SB2_2_27/i0_0 ), .A3(\SB2_2_27/i1_7 ), .ZN(
        \SB2_2_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_2/Component_Function_0/N2  ( .A1(\SB2_2_2/i0[8] ), .A2(
        \SB2_2_2/i0[7] ), .A3(\SB2_2_2/i0[6] ), .ZN(
        \SB2_2_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U932 ( .A1(\SB2_2_2/i0_3 ), .A2(\SB2_2_2/i0[8] ), .A3(
        \SB2_2_2/i1_7 ), .ZN(\SB2_2_2/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U6125 ( .A1(\SB2_2_15/i0_0 ), .A2(\SB2_2_15/i0_3 ), .A3(
        \SB2_2_15/i0[7] ), .ZN(\SB2_2_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_11/Component_Function_0/N4  ( .A1(\SB2_2_11/i0[7] ), .A2(
        \SB2_2_11/i0_3 ), .A3(\SB2_2_11/i0_0 ), .ZN(
        \SB2_2_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_23/Component_Function_3/N4  ( .A1(\SB2_2_23/i1_5 ), .A2(
        \SB2_2_23/i0[8] ), .A3(\SB2_2_23/i3[0] ), .ZN(
        \SB2_2_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U7913 ( .A1(\SB2_2_18/i1_7 ), .A2(\SB2_2_18/i0_4 ), .A3(
        \SB2_2_18/i0[8] ), .ZN(\SB2_2_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_3/Component_Function_1/N3  ( .A1(n3994), .A2(\SB2_2_3/i0[6] ), .A3(\SB2_2_3/i0[9] ), .ZN(\SB2_2_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_1/Component_Function_1/N3  ( .A1(\SB2_2_1/i1_5 ), .A2(
        \SB2_2_1/i0[6] ), .A3(\SB2_2_1/i0[9] ), .ZN(
        \SB2_2_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_11/Component_Function_4/N3  ( .A1(\SB2_2_11/i0[9] ), .A2(
        \SB2_2_11/i0[10] ), .A3(\SB2_2_11/i0_3 ), .ZN(
        \SB2_2_11/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_3/Component_Function_1/N1  ( .A1(\SB2_2_3/i0_3 ), .A2(
        \SB2_2_3/i1[9] ), .ZN(\SB2_2_3/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_27/Component_Function_0/N1  ( .A1(\SB2_2_27/i0[10] ), .A2(
        \SB2_2_27/i0[9] ), .ZN(\SB2_2_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_9/Component_Function_0/N2  ( .A1(\SB2_2_9/i0[8] ), .A2(
        \SB2_2_9/i0[7] ), .A3(\SB2_2_9/i0[6] ), .ZN(
        \SB2_2_9/Component_Function_0/NAND4_in[1] ) );
  INV_X1 \SB2_2_20/INV_1  ( .I(\SB1_2_24/buf_output[1] ), .ZN(\SB2_2_20/i1_7 )
         );
  NAND3_X1 \SB2_2_9/Component_Function_0/N3  ( .A1(\SB2_2_9/i0[10] ), .A2(
        \SB2_2_9/i0_4 ), .A3(\SB2_2_9/i0_3 ), .ZN(
        \SB2_2_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_9/Component_Function_4/N3  ( .A1(\SB2_2_9/i0[9] ), .A2(
        \SB2_2_9/i0[10] ), .A3(\SB2_2_9/i0_3 ), .ZN(
        \SB2_2_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U7456 ( .A1(\SB2_2_27/i0[9] ), .A2(\SB2_2_27/i0_3 ), .A3(
        \SB2_2_27/i0[8] ), .ZN(n2404) );
  NAND3_X1 \SB2_2_30/Component_Function_3/N4  ( .A1(\SB2_2_30/i1_5 ), .A2(
        \SB2_2_30/i0[8] ), .A3(\SB2_2_30/i3[0] ), .ZN(
        \SB2_2_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_5/Component_Function_0/N2  ( .A1(\SB2_2_5/i0[8] ), .A2(
        \SB2_2_5/i0[7] ), .A3(\SB2_2_5/i0[6] ), .ZN(
        \SB2_2_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_21/Component_Function_1/N4  ( .A1(\SB2_2_21/i1_7 ), .A2(
        \SB2_2_21/i0[8] ), .A3(\SB1_2_22/buf_output[4] ), .ZN(
        \SB2_2_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3429 ( .A1(\SB2_2_23/i0[7] ), .A2(\SB2_2_23/i0_0 ), .A3(
        \SB2_2_23/i0_3 ), .ZN(\SB2_2_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2263 ( .A1(\SB2_2_27/i1_5 ), .A2(\SB2_2_27/i0[6] ), .A3(
        \SB2_2_27/i0[9] ), .ZN(\SB2_2_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2275 ( .A1(\SB2_2_22/i0[6] ), .A2(\SB2_2_22/i1_5 ), .A3(
        \SB2_2_22/i0[9] ), .ZN(n1959) );
  NAND3_X1 \SB2_2_3/Component_Function_3/N2  ( .A1(\SB2_2_3/i0_0 ), .A2(
        \SB1_2_3/buf_output[5] ), .A3(\SB1_2_4/buf_output[4] ), .ZN(
        \SB2_2_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_16/Component_Function_2/N4  ( .A1(\SB2_2_16/i1_5 ), .A2(
        \SB2_2_16/i0_0 ), .A3(\SB2_2_16/i0_4 ), .ZN(
        \SB2_2_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_9/Component_Function_3/N1  ( .A1(\SB2_2_9/i1[9] ), .A2(
        \SB2_2_9/i0_3 ), .A3(\SB2_2_9/i0[6] ), .ZN(
        \SB2_2_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_1/N4  ( .A1(\SB2_2_16/i1_7 ), .A2(
        \SB2_2_16/i0[8] ), .A3(\SB2_2_16/i0_4 ), .ZN(
        \SB2_2_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U5251 ( .A1(\SB2_2_27/i0[9] ), .A2(\SB2_2_27/i0_4 ), .A3(
        \SB2_2_27/i0[6] ), .ZN(n2175) );
  NAND2_X1 \SB2_2_5/Component_Function_0/N1  ( .A1(\SB2_2_5/i0[10] ), .A2(
        \SB2_2_5/i0[9] ), .ZN(\SB2_2_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U919 ( .A1(\SB2_2_17/i0_3 ), .A2(\RI3[2][88] ), .A3(
        \SB2_2_17/i0[10] ), .ZN(n1012) );
  NAND3_X1 \SB2_2_17/Component_Function_1/N2  ( .A1(\SB2_2_17/i0_3 ), .A2(
        \SB2_2_17/i1_7 ), .A3(\SB2_2_17/i0[8] ), .ZN(
        \SB2_2_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_20/Component_Function_1/N2  ( .A1(\SB2_2_20/i0_3 ), .A2(
        \SB2_2_20/i1_7 ), .A3(\SB2_2_20/i0[8] ), .ZN(
        \SB2_2_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U6108 ( .A1(\SB1_2_12/buf_output[4] ), .A2(\SB2_2_11/i1_7 ), .A3(
        \SB2_2_11/i0[8] ), .ZN(n2014) );
  NAND3_X1 U5609 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0[10] ), .A3(
        \SB2_2_22/i0_4 ), .ZN(n2416) );
  NAND3_X1 U6521 ( .A1(\RI3[2][88] ), .A2(\SB2_2_17/i1_7 ), .A3(
        \SB2_2_17/i0[8] ), .ZN(\SB2_2_17/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U1355 ( .I(\MC_ARK_ARC_1_2/buf_output[66] ), .ZN(\SB1_3_20/i3[0] ) );
  NAND3_X1 U909 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i0[9] ), .A3(
        \SB1_3_5/i0[10] ), .ZN(\SB1_3_5/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U1848 ( .I(\MC_ARK_ARC_1_2/buf_output[54] ), .ZN(\SB1_3_22/i3[0] ) );
  INV_X1 \SB1_3_10/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[126] ), .ZN(
        \SB1_3_10/i3[0] ) );
  INV_X1 \SB1_3_8/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[138] ), .ZN(
        \SB1_3_8/i3[0] ) );
  INV_X1 \SB1_3_15/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[96] ), .ZN(
        \SB1_3_15/i3[0] ) );
  INV_X1 \SB1_3_15/INV_5  ( .I(\RI1[3][101] ), .ZN(\SB1_3_15/i1_5 ) );
  BUF_X2 \SB1_3_19/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[72] ), .Z(
        \SB1_3_19/i0[9] ) );
  BUF_X2 U1775 ( .I(\MC_ARK_ARC_1_2/buf_output[13] ), .Z(\SB1_3_29/i0[6] ) );
  NAND3_X1 U2742 ( .A1(\SB1_3_13/i0[10] ), .A2(\SB1_3_13/i0[9] ), .A3(
        \SB1_3_13/i0_3 ), .ZN(\SB1_3_13/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_4/N2  ( .A1(\SB1_3_13/i3[0] ), .A2(
        \SB1_3_13/i0_0 ), .A3(\SB1_3_13/i1_7 ), .ZN(
        \SB1_3_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_2/N1  ( .A1(\SB1_3_2/i1_5 ), .A2(
        \SB1_3_2/i0[10] ), .A3(\SB1_3_2/i1[9] ), .ZN(
        \SB1_3_2/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U7836 ( .A1(\SB1_3_5/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_3_5/Component_Function_4/NAND4_in[2] ), .ZN(n2599) );
  NAND3_X1 \SB1_3_23/Component_Function_4/N4  ( .A1(\SB1_3_23/i1[9] ), .A2(
        \SB1_3_23/i1_5 ), .A3(\SB1_3_23/i0_4 ), .ZN(
        \SB1_3_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_24/Component_Function_1/N3  ( .A1(\SB1_3_24/i1_5 ), .A2(
        \SB1_3_24/i0[6] ), .A3(\SB1_3_24/i0[9] ), .ZN(
        \SB1_3_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_24/Component_Function_1/N2  ( .A1(\SB1_3_24/i0_3 ), .A2(
        \SB1_3_24/i1_7 ), .A3(\SB1_3_24/i0[8] ), .ZN(
        \SB1_3_24/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_13/Component_Function_4/N4  ( .A1(\SB1_3_13/i1[9] ), .A2(
        \SB1_3_13/i1_5 ), .A3(\SB1_3_13/i0_4 ), .ZN(
        \SB1_3_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U7893 ( .A1(\SB1_3_23/i0_0 ), .A2(\SB1_3_23/i3[0] ), .A3(
        \SB1_3_23/i1_7 ), .ZN(\SB1_3_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U7146 ( .A1(\SB1_3_23/i0[9] ), .A2(\SB1_3_23/i0_0 ), .A3(
        \SB1_3_23/i0[8] ), .ZN(n2262) );
  NAND3_X1 \SB1_3_24/Component_Function_1/N4  ( .A1(\SB1_3_24/i1_7 ), .A2(
        \SB1_3_24/i0[8] ), .A3(\SB1_3_24/i0_4 ), .ZN(
        \SB1_3_24/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_3_13/Component_Function_0/N1  ( .A1(\SB1_3_13/i0[10] ), .A2(
        \SB1_3_13/i0[9] ), .ZN(\SB1_3_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_4/N3  ( .A1(\SB1_3_18/i0[9] ), .A2(
        \SB1_3_18/i0[10] ), .A3(\SB1_3_18/i0_3 ), .ZN(
        \SB1_3_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U5908 ( .A1(\SB1_3_16/i0[10] ), .A2(\SB1_3_16/i0_3 ), .A3(
        \SB1_3_16/i0[6] ), .ZN(\SB1_3_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3074 ( .A1(\SB1_3_4/i0_0 ), .A2(\SB1_3_4/i1_7 ), .A3(
        \SB1_3_4/i3[0] ), .ZN(\SB1_3_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_9/Component_Function_3/N3  ( .A1(\SB1_3_9/i1[9] ), .A2(
        \SB1_3_9/i1_7 ), .A3(\SB1_3_9/i0[10] ), .ZN(
        \SB1_3_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_23/Component_Function_1/N3  ( .A1(\SB1_3_23/i1_5 ), .A2(
        \SB1_3_23/i0[6] ), .A3(\SB1_3_23/i0[9] ), .ZN(
        \SB1_3_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_31/Component_Function_0/N2  ( .A1(n5441), .A2(
        \SB1_3_31/i0[7] ), .A3(\SB1_3_31/i0[6] ), .ZN(
        \SB1_3_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_24/Component_Function_5/N1  ( .A1(\SB1_3_24/i0_0 ), .A2(
        \SB1_3_24/i3[0] ), .ZN(\SB1_3_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_4/N4  ( .A1(\SB1_3_16/i1[9] ), .A2(
        \SB1_3_16/i1_5 ), .A3(\SB1_3_16/i0_4 ), .ZN(
        \SB1_3_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U5226 ( .A1(\SB1_3_1/i0_0 ), .A2(\SB1_3_1/i1_5 ), .A3(
        \SB1_3_1/i0_4 ), .ZN(n2724) );
  NAND2_X1 \SB1_3_2/Component_Function_0/N1  ( .A1(\SB1_3_2/i0[10] ), .A2(
        \SB1_3_2/i0[9] ), .ZN(\SB1_3_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3909 ( .A1(\SB1_3_20/i1_5 ), .A2(\SB1_3_20/i0[6] ), .A3(
        \SB1_3_20/i0[9] ), .ZN(\SB1_3_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U863 ( .A1(\SB1_3_31/i1_5 ), .A2(\SB1_3_31/i1[9] ), .A3(
        \SB1_3_31/i0_4 ), .ZN(n2984) );
  NAND2_X1 U7130 ( .A1(n2262), .A2(\SB1_3_23/Component_Function_4/NAND4_in[1] ), .ZN(n2255) );
  NAND3_X1 \SB1_3_22/Component_Function_1/N3  ( .A1(\SB1_3_22/i1_5 ), .A2(
        \SB1_3_22/i0[6] ), .A3(\SB1_3_22/i0[9] ), .ZN(
        \SB1_3_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_27/Component_Function_5/N2  ( .A1(\SB1_3_27/i0_0 ), .A2(
        \SB1_3_27/i0[6] ), .A3(\SB1_3_27/i0[10] ), .ZN(
        \SB1_3_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U860 ( .A1(\SB1_3_18/i0[10] ), .A2(\SB1_3_18/i1[9] ), .A3(
        \SB1_3_18/i1_7 ), .ZN(n1725) );
  NAND3_X1 \SB1_3_29/Component_Function_0/N2  ( .A1(\SB1_3_29/i0[8] ), .A2(
        \SB1_3_29/i0[7] ), .A3(\SB1_3_29/i0[6] ), .ZN(
        \SB1_3_29/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_1/N2  ( .A1(\SB1_3_2/i0_3 ), .A2(
        \SB1_3_2/i1_7 ), .A3(\SB1_3_2/i0[8] ), .ZN(
        \SB1_3_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_2/Component_Function_1/N1  ( .A1(\SB1_3_2/i0_3 ), .A2(
        \SB1_3_2/i1[9] ), .ZN(\SB1_3_2/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_19/Component_Function_1/N1  ( .A1(\SB1_3_19/i0_3 ), .A2(
        \SB1_3_19/i1[9] ), .ZN(\SB1_3_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2764 ( .A1(\SB1_3_6/i0[9] ), .A2(\SB1_3_6/i0[6] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[154] ), .ZN(n684) );
  INV_X1 \SB2_3_20/INV_1  ( .I(\SB1_3_24/buf_output[1] ), .ZN(\SB2_3_20/i1_7 )
         );
  BUF_X2 U835 ( .I(\SB1_3_3/buf_output[0] ), .Z(\SB2_3_30/i0[9] ) );
  INV_X1 \SB2_3_1/INV_0  ( .I(\SB1_3_6/buf_output[0] ), .ZN(\SB2_3_1/i3[0] )
         );
  INV_X1 \SB2_3_2/INV_0  ( .I(\SB1_3_7/buf_output[0] ), .ZN(\SB2_3_2/i3[0] )
         );
  NAND2_X1 \SB2_3_7/Component_Function_5/N1  ( .A1(\SB2_3_7/i0_0 ), .A2(
        \SB2_3_7/i3[0] ), .ZN(\SB2_3_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_4/N2  ( .A1(\SB2_3_21/i3[0] ), .A2(
        \SB2_3_21/i0_0 ), .A3(\SB2_3_21/i1_7 ), .ZN(
        \SB2_3_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_24/Component_Function_1/N2  ( .A1(\SB2_3_24/i0_3 ), .A2(
        \SB2_3_24/i1_7 ), .A3(\SB2_3_24/i0[8] ), .ZN(
        \SB2_3_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_24/Component_Function_5/N1  ( .A1(\SB2_3_24/i0_0 ), .A2(
        \SB2_3_24/i3[0] ), .ZN(\SB2_3_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_31/Component_Function_2/N1  ( .A1(\SB2_3_31/i1_5 ), .A2(
        \SB2_3_31/i0[10] ), .A3(\SB2_3_31/i1[9] ), .ZN(
        \SB2_3_31/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_1/Component_Function_5/N1  ( .A1(\SB2_3_1/i0_0 ), .A2(
        \SB2_3_1/i3[0] ), .ZN(\SB2_3_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U6483 ( .A1(\SB1_3_18/buf_output[5] ), .A2(\SB2_3_18/i1[9] ), .A3(
        \SB2_3_18/i0_4 ), .ZN(\SB2_3_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U6938 ( .A1(\SB1_3_31/buf_output[4] ), .A2(\SB2_3_30/i0_3 ), .A3(
        \SB2_3_30/i1[9] ), .ZN(n2164) );
  NAND3_X1 \SB2_3_30/Component_Function_3/N1  ( .A1(\SB2_3_30/i1[9] ), .A2(
        \SB2_3_30/i0_3 ), .A3(\SB2_3_30/i0[6] ), .ZN(
        \SB2_3_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U6044 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0[8] ), .A3(
        \SB2_3_17/i1_7 ), .ZN(\SB2_3_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_0/Component_Function_3/N4  ( .A1(\SB2_3_0/i1_5 ), .A2(
        \SB2_3_0/i0[8] ), .A3(\SB2_3_0/i3[0] ), .ZN(
        \SB2_3_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_3/N3  ( .A1(\SB2_3_12/i1[9] ), .A2(
        \SB2_3_12/i1_7 ), .A3(\SB2_3_12/i0[10] ), .ZN(
        \SB2_3_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_20/Component_Function_1/N2  ( .A1(\SB2_3_20/i0_3 ), .A2(
        \SB2_3_20/i1_7 ), .A3(\SB2_3_20/i0[8] ), .ZN(
        \SB2_3_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_27/Component_Function_1/N4  ( .A1(\SB2_3_27/i1_7 ), .A2(
        \SB2_3_27/i0[8] ), .A3(\SB2_3_27/i0_4 ), .ZN(
        \SB2_3_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_5/Component_Function_2/N3  ( .A1(\SB2_3_5/i0_3 ), .A2(
        \SB2_3_5/i0[8] ), .A3(\SB2_3_5/i0[9] ), .ZN(
        \SB2_3_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_31/Component_Function_4/N4  ( .A1(\SB2_3_31/i1[9] ), .A2(
        \SB2_3_31/i1_5 ), .A3(\SB1_3_0/buf_output[4] ), .ZN(
        \SB2_3_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_2/N1  ( .A1(\SB2_3_12/i1_5 ), .A2(
        \SB2_3_12/i0[10] ), .A3(\SB2_3_12/i1[9] ), .ZN(
        \SB2_3_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_4/N4  ( .A1(\SB2_3_18/i1[9] ), .A2(
        \SB2_3_18/i1_5 ), .A3(\SB2_3_18/i0_4 ), .ZN(
        \SB2_3_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U6121 ( .A1(\SB2_3_2/i0_0 ), .A2(\SB2_3_2/i0[9] ), .A3(
        \SB2_3_2/i0[8] ), .ZN(\SB2_3_2/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_0/Component_Function_0/N1  ( .A1(\SB2_3_0/i0[10] ), .A2(
        \SB2_3_0/i0[9] ), .ZN(\SB2_3_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U4020 ( .A1(\SB2_3_11/i0[10] ), .A2(\SB2_3_11/i0_3 ), .A3(
        \SB2_3_11/i0[9] ), .ZN(n1133) );
  NAND3_X1 \SB2_3_17/Component_Function_1/N3  ( .A1(\SB2_3_17/i1_5 ), .A2(
        \SB2_3_17/i0[6] ), .A3(\SB2_3_17/i0[9] ), .ZN(
        \SB2_3_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U8313 ( .A1(n4081), .A2(\SB2_3_26/i0[8] ), .A3(\SB2_3_26/i0[6] ), 
        .ZN(\SB2_3_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_17/Component_Function_0/N2  ( .A1(\SB2_3_17/i0[8] ), .A2(
        \SB2_3_17/i0[7] ), .A3(\SB2_3_17/i0[6] ), .ZN(
        \SB2_3_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2336 ( .A1(\SB2_3_10/i1_5 ), .A2(\SB2_3_10/i0[10] ), .A3(
        \SB2_3_10/i1[9] ), .ZN(\SB2_3_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4511 ( .A1(\SB2_3_18/i0[10] ), .A2(\SB2_3_18/i1_7 ), .A3(
        \SB2_3_18/i1[9] ), .ZN(n2231) );
  NAND3_X1 \SB2_3_26/Component_Function_1/N2  ( .A1(\SB2_3_26/i0_3 ), .A2(
        \SB2_3_26/i1_7 ), .A3(\SB2_3_26/i0[8] ), .ZN(
        \SB2_3_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_22/Component_Function_2/N2  ( .A1(\SB2_3_22/i0_3 ), .A2(
        \SB2_3_22/i0[10] ), .A3(\SB2_3_22/i0[6] ), .ZN(
        \SB2_3_22/Component_Function_2/NAND4_in[1] ) );
  INV_X1 \SB1_4_31/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[1] ), .ZN(
        \SB1_4_31/i1_7 ) );
  INV_X1 U5362 ( .I(\MC_ARK_ARC_1_3/buf_output[175] ), .ZN(\SB1_4_2/i1_7 ) );
  BUF_X2 \SB1_4_20/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[66] ), .Z(
        \SB1_4_20/i0[9] ) );
  INV_X1 \SB1_4_5/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[161] ), .ZN(
        \SB1_4_5/i1_5 ) );
  INV_X1 \SB1_4_3/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[169] ), .ZN(
        \SB1_4_3/i1_7 ) );
  BUF_X2 \SB1_4_31/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[1] ), .Z(
        \SB1_4_31/i0[6] ) );
  BUF_X2 U5454 ( .I(\MC_ARK_ARC_1_3/buf_output[98] ), .Z(\SB1_4_15/i0_0 ) );
  NAND3_X1 U786 ( .A1(\SB1_4_31/i0_4 ), .A2(\SB1_4_31/i1_5 ), .A3(
        \SB1_4_31/i1[9] ), .ZN(n2346) );
  BUF_X2 \SB1_4_26/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[30] ), .Z(
        \SB1_4_26/i0[9] ) );
  NAND2_X1 \SB1_4_3/Component_Function_1/N1  ( .A1(\SB1_4_3/i0_3 ), .A2(
        \SB1_4_3/i1[9] ), .ZN(\SB1_4_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_2/Component_Function_2/N4  ( .A1(\SB1_4_2/i1_5 ), .A2(
        \SB1_4_2/i0_0 ), .A3(\SB1_4_2/i0_4 ), .ZN(
        \SB1_4_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_25/Component_Function_3/N4  ( .A1(\SB1_4_25/i1_5 ), .A2(
        \SB1_4_25/i0[8] ), .A3(\SB1_4_25/i3[0] ), .ZN(
        \SB1_4_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_22/Component_Function_2/N2  ( .A1(\RI1[4][59] ), .A2(
        \SB1_4_22/i0[10] ), .A3(\SB1_4_22/i0[6] ), .ZN(
        \SB1_4_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_5/Component_Function_2/N4  ( .A1(\SB1_4_5/i1_5 ), .A2(
        \SB1_4_5/i0_0 ), .A3(\SB1_4_5/i0_4 ), .ZN(
        \SB1_4_5/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 \SB1_4_17/Component_Function_0/N1  ( .A1(\SB1_4_17/i0[10] ), .A2(
        \SB1_4_17/i0[9] ), .ZN(\SB1_4_17/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_1/Component_Function_1/N1  ( .A1(\SB1_4_1/i0_3 ), .A2(
        \SB1_4_1/i1[9] ), .ZN(\SB1_4_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3220 ( .A1(\SB1_4_1/i0_0 ), .A2(\SB1_4_1/i0_4 ), .A3(
        \SB1_4_1/i1_5 ), .ZN(\SB1_4_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_26/Component_Function_3/N2  ( .A1(\SB1_4_26/i0_0 ), .A2(
        \SB1_4_26/i0_3 ), .A3(\SB1_4_26/i0_4 ), .ZN(
        \SB1_4_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_5/Component_Function_0/N3  ( .A1(\SB1_4_5/i0[10] ), .A2(
        \SB1_4_5/i0_4 ), .A3(\SB1_4_5/i0_3 ), .ZN(
        \SB1_4_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1552 ( .A1(\SB1_4_2/i0_3 ), .A2(\SB1_4_2/i0[10] ), .A3(
        \SB1_4_2/i0[6] ), .ZN(\SB1_4_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_4/Component_Function_4/N4  ( .A1(\SB1_4_4/i1[9] ), .A2(
        \SB1_4_4/i1_5 ), .A3(\SB1_4_4/i0_4 ), .ZN(
        \SB1_4_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_31/Component_Function_3/N3  ( .A1(\SB1_4_31/i1[9] ), .A2(
        \SB1_4_31/i1_7 ), .A3(\SB1_4_31/i0[10] ), .ZN(
        \SB1_4_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_5/Component_Function_0/N4  ( .A1(\SB1_4_5/i0[7] ), .A2(
        \SB1_4_5/i0_3 ), .A3(\SB1_4_5/i0_0 ), .ZN(
        \SB1_4_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_21/Component_Function_1/N4  ( .A1(\SB1_4_21/i1_7 ), .A2(
        \SB1_4_21/i0[8] ), .A3(\SB1_4_21/i0_4 ), .ZN(
        \SB1_4_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U6633 ( .A1(\RI1[4][59] ), .A2(\SB1_4_22/i0[7] ), .A3(
        \SB1_4_22/i0_0 ), .ZN(n2025) );
  NAND3_X1 \SB1_4_7/Component_Function_2/N2  ( .A1(\SB1_4_7/i0_3 ), .A2(
        \SB1_4_7/i0[10] ), .A3(\SB1_4_7/i0[6] ), .ZN(
        \SB1_4_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_15/Component_Function_4/N1  ( .A1(\SB1_4_15/i0[9] ), .A2(
        \SB1_4_15/i0_0 ), .A3(\SB1_4_15/i0[8] ), .ZN(
        \SB1_4_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U745 ( .A1(\SB1_4_4/i0_0 ), .A2(\SB1_4_4/i1_5 ), .A3(\SB1_4_4/i0_4 ), .ZN(n2246) );
  NAND3_X1 U707 ( .A1(\SB1_4_0/i0_3 ), .A2(\SB1_4_0/i0[7] ), .A3(
        \SB1_4_0/i0_0 ), .ZN(n2593) );
  NAND3_X1 U5792 ( .A1(\SB1_4_15/i0[9] ), .A2(\SB1_4_15/i1_5 ), .A3(
        \SB1_4_15/i0[6] ), .ZN(\SB1_4_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_30/Component_Function_1/N2  ( .A1(\SB1_4_30/i0_3 ), .A2(
        \SB1_4_30/i1_7 ), .A3(\SB1_4_30/i0[8] ), .ZN(
        \SB1_4_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4738 ( .A1(\RI1[4][59] ), .A2(\SB1_4_22/i0[9] ), .A3(
        \SB1_4_22/i0[10] ), .ZN(n1538) );
  NAND2_X1 \SB1_4_5/Component_Function_5/N1  ( .A1(\SB1_4_5/i0_0 ), .A2(
        \SB1_4_5/i3[0] ), .ZN(\SB1_4_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_11/Component_Function_3/N2  ( .A1(\SB1_4_11/i0_0 ), .A2(
        \SB1_4_11/i0_3 ), .A3(\SB1_4_11/i0_4 ), .ZN(
        \SB1_4_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U5425 ( .A1(\SB1_4_12/i0_0 ), .A2(\RI1[4][119] ), .A3(
        \SB1_4_12/i0_4 ), .ZN(\SB1_4_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U6674 ( .A1(\SB1_4_6/i0[10] ), .A2(\RI1[4][155] ), .A3(
        \SB1_4_6/i0_4 ), .ZN(n2268) );
  NAND3_X1 \SB1_4_9/Component_Function_5/N2  ( .A1(\SB1_4_9/i0_0 ), .A2(
        \SB1_4_9/i0[6] ), .A3(\SB1_4_9/i0[10] ), .ZN(
        \SB1_4_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_20/Component_Function_5/N2  ( .A1(\SB1_4_20/i0_0 ), .A2(
        \SB1_4_20/i0[6] ), .A3(\SB1_4_20/i0[10] ), .ZN(
        \SB1_4_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_12/Component_Function_2/N1  ( .A1(\SB1_4_12/i1_5 ), .A2(
        \SB1_4_12/i0[10] ), .A3(\SB1_4_12/i1[9] ), .ZN(
        \SB1_4_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_10/Component_Function_3/N3  ( .A1(\SB1_4_10/i1[9] ), .A2(
        \SB1_4_10/i1_7 ), .A3(n1491), .ZN(
        \SB1_4_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_22/Component_Function_3/N1  ( .A1(\SB1_4_22/i1[9] ), .A2(
        \RI1[4][59] ), .A3(\SB1_4_22/i0[6] ), .ZN(
        \SB1_4_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_26/Component_Function_4/N3  ( .A1(\SB1_4_26/i0[9] ), .A2(
        \SB1_4_26/i0[10] ), .A3(\SB1_4_26/i0_3 ), .ZN(
        \SB1_4_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_16/Component_Function_0/N3  ( .A1(\SB1_4_16/i0[10] ), .A2(
        \SB1_4_16/i0_4 ), .A3(\SB1_4_16/i0_3 ), .ZN(
        \SB1_4_16/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_13/Component_Function_5/N1  ( .A1(\SB2_4_13/i0_0 ), .A2(
        \SB2_4_13/i3[0] ), .ZN(\SB2_4_13/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_2/Component_Function_5/N1  ( .A1(\SB2_4_2/i0_0 ), .A2(
        \SB2_4_2/i3[0] ), .ZN(\SB2_4_2/Component_Function_5/NAND4_in[0] ) );
  INV_X1 \SB2_4_10/INV_1  ( .I(\RI3[4][127] ), .ZN(\SB2_4_10/i1_7 ) );
  INV_X1 \SB2_4_9/INV_1  ( .I(\SB1_4_13/buf_output[1] ), .ZN(\SB2_4_9/i1_7 )
         );
  INV_X1 \SB2_4_18/INV_1  ( .I(\SB1_4_22/buf_output[1] ), .ZN(\SB2_4_18/i1_7 )
         );
  BUF_X2 \SB2_4_12/BUF_0  ( .I(\SB1_4_17/buf_output[0] ), .Z(\SB2_4_12/i0[9] )
         );
  INV_X1 \SB2_4_8/INV_4  ( .I(n3183), .ZN(\SB2_4_8/i0[7] ) );
  BUF_X2 \SB2_4_26/BUF_1  ( .I(\SB1_4_30/buf_output[1] ), .Z(\SB2_4_26/i0[6] )
         );
  NAND3_X1 \SB2_4_31/Component_Function_4/N2  ( .A1(\SB2_4_31/i3[0] ), .A2(
        \SB2_4_31/i0_0 ), .A3(\SB2_4_31/i1_7 ), .ZN(
        \SB2_4_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_13/Component_Function_4/N2  ( .A1(\SB2_4_13/i3[0] ), .A2(
        \SB2_4_13/i0_0 ), .A3(\SB2_4_13/i1_7 ), .ZN(
        \SB2_4_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1536 ( .A1(\SB2_4_28/i1[9] ), .A2(\SB2_4_28/i0_3 ), .A3(
        \SB2_4_28/i0[6] ), .ZN(\SB2_4_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_26/Component_Function_4/N4  ( .A1(\SB2_4_26/i1[9] ), .A2(
        \SB2_4_26/i1_5 ), .A3(\SB2_4_26/i0_4 ), .ZN(
        \SB2_4_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_19/Component_Function_3/N4  ( .A1(\SB2_4_19/i1_5 ), .A2(
        \SB2_4_19/i0[8] ), .A3(\SB2_4_19/i3[0] ), .ZN(
        \SB2_4_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3387 ( .A1(\SB2_4_11/i0[10] ), .A2(\SB2_4_11/i1[9] ), .A3(
        \SB2_4_11/i1_7 ), .ZN(n904) );
  NAND3_X1 \SB2_4_18/Component_Function_1/N3  ( .A1(\SB2_4_18/i1_5 ), .A2(
        \SB2_4_18/i0[6] ), .A3(\SB2_4_18/i0[9] ), .ZN(
        \SB2_4_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U5515 ( .A1(\SB2_4_11/i0[10] ), .A2(\SB2_4_11/i1_5 ), .A3(
        \SB2_4_11/i1[9] ), .ZN(\SB2_4_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U7046 ( .A1(\SB2_4_6/i0_4 ), .A2(\SB2_4_6/i1[9] ), .A3(
        \SB2_4_6/i1_5 ), .ZN(n2216) );
  NAND3_X1 \SB2_4_24/Component_Function_1/N3  ( .A1(n6268), .A2(
        \SB2_4_24/i0[6] ), .A3(\SB2_4_24/i0[9] ), .ZN(
        \SB2_4_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_16/Component_Function_4/N4  ( .A1(\SB2_4_16/i1[9] ), .A2(
        \SB2_4_16/i1_5 ), .A3(\SB2_4_16/i0_4 ), .ZN(
        \SB2_4_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U7183 ( .A1(\SB2_4_9/i0_3 ), .A2(\SB2_4_9/i0[10] ), .A3(
        \SB2_4_9/i0[9] ), .ZN(\SB2_4_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4346 ( .A1(\SB2_4_2/i0_4 ), .A2(\SB2_4_2/i1_7 ), .A3(
        \SB2_4_2/i0[8] ), .ZN(\SB2_4_2/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_4_12/Component_Function_1/N1  ( .A1(\SB2_4_12/i0_3 ), .A2(
        \SB2_4_12/i1[9] ), .ZN(\SB2_4_12/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 U693 ( .A1(\SB2_4_25/i0[6] ), .A2(n1026), .ZN(n1025) );
  NAND3_X1 \SB2_4_7/Component_Function_3/N3  ( .A1(\SB2_4_7/i1[9] ), .A2(
        \SB2_4_7/i1_7 ), .A3(\SB2_4_7/i0[10] ), .ZN(
        \SB2_4_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_7/Component_Function_3/N1  ( .A1(\SB2_4_7/i1[9] ), .A2(
        \SB2_4_7/i0_3 ), .A3(\SB2_4_7/i0[6] ), .ZN(
        \SB2_4_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_18/Component_Function_1/N2  ( .A1(\SB2_4_18/i0_3 ), .A2(
        \SB2_4_18/i1_7 ), .A3(\SB2_4_18/i0[8] ), .ZN(
        \SB2_4_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U6159 ( .A1(\SB2_4_7/i0[6] ), .A2(\SB2_4_7/i0[8] ), .A3(
        \SB2_4_7/i0[7] ), .ZN(n1808) );
  NAND3_X1 U6782 ( .A1(\SB2_4_7/i0[8] ), .A2(\SB2_4_7/i3[0] ), .A3(
        \SB2_4_7/i1_5 ), .ZN(n2228) );
  BUF_X2 \MC_ARK_ARC_1_4/BUF_18  ( .I(\SB2_4_1/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[18] ) );
  BUF_X2 \SB3_29/BUF_1  ( .I(\MC_ARK_ARC_1_4/buf_output[13] ), .Z(
        \SB3_29/i0[6] ) );
  BUF_X2 U1950 ( .I(\MC_ARK_ARC_1_4/buf_output[43] ), .Z(\SB3_24/i0[6] ) );
  INV_X1 \SB3_22/INV_3  ( .I(\MC_ARK_ARC_1_4/buf_output[57] ), .ZN(
        \SB3_22/i0[8] ) );
  NAND2_X1 \SB3_27/Component_Function_5/N1  ( .A1(\SB3_27/i0_0 ), .A2(
        \SB3_27/i3[0] ), .ZN(\SB3_27/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 \SB3_3/BUF_1  ( .I(\MC_ARK_ARC_1_4/buf_output[169] ), .Z(
        \SB3_3/i0[6] ) );
  INV_X1 \SB3_25/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[36] ), .ZN(
        \SB3_25/i3[0] ) );
  BUF_X2 \SB3_3/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[168] ), .Z(
        \SB3_3/i0[9] ) );
  INV_X1 U5377 ( .I(\MC_ARK_ARC_1_4/buf_output[97] ), .ZN(\SB3_15/i1_7 ) );
  INV_X1 U1423 ( .I(\MC_ARK_ARC_1_4/buf_output[158] ), .ZN(\SB3_5/i1[9] ) );
  NAND3_X1 \SB3_30/Component_Function_2/N3  ( .A1(\RI1[5][11] ), .A2(
        \SB3_30/i0[8] ), .A3(\SB3_30/i0[9] ), .ZN(
        \SB3_30/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 \SB3_14/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[102] ), .Z(
        \SB3_14/i0[9] ) );
  BUF_X2 \SB3_29/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[12] ), .Z(
        \SB3_29/i0[9] ) );
  INV_X1 U1318 ( .I(\MC_ARK_ARC_1_4/buf_output[151] ), .ZN(\SB3_6/i1_7 ) );
  INV_X1 \SB3_5/INV_5  ( .I(n4006), .ZN(\SB3_5/i1_5 ) );
  INV_X1 \SB3_24/INV_5  ( .I(n3971), .ZN(\SB3_24/i1_5 ) );
  INV_X1 U1678 ( .I(n4001), .ZN(\SB3_13/i0[8] ) );
  NAND3_X1 \SB3_0/Component_Function_1/N2  ( .A1(\SB3_0/i0_3 ), .A2(
        \SB3_0/i1_7 ), .A3(\SB3_0/i0[8] ), .ZN(
        \SB3_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4453 ( .A1(\SB3_7/i0_3 ), .A2(\SB3_7/i0[8] ), .A3(\SB3_7/i0[9] ), 
        .ZN(\SB3_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_7/Component_Function_5/N4  ( .A1(\SB3_7/i0[9] ), .A2(
        \SB3_7/i0[6] ), .A3(\SB3_7/i0_4 ), .ZN(
        \SB3_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_2/Component_Function_4/N1  ( .A1(\SB3_2/i0[9] ), .A2(
        \SB3_2/i0_0 ), .A3(\SB3_2/i0[8] ), .ZN(
        \SB3_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U5354 ( .A1(\SB3_27/i1_7 ), .A2(\SB3_27/i0[8] ), .A3(\SB3_27/i0_4 ), 
        .ZN(\SB3_27/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB3_25/Component_Function_0/N1  ( .A1(\SB3_25/i0[10] ), .A2(
        \SB3_25/i0[9] ), .ZN(\SB3_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U4298 ( .A1(\SB3_0/i0_0 ), .A2(\SB3_0/i0_3 ), .A3(\SB3_0/i0_4 ), 
        .ZN(\SB3_0/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U4138 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i1[9] ), .ZN(n1176) );
  NAND3_X1 \SB3_12/Component_Function_1/N3  ( .A1(\SB3_12/i1_5 ), .A2(
        \SB3_12/i0[6] ), .A3(\SB3_12/i0[9] ), .ZN(
        \SB3_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U7270 ( .A1(\SB3_11/i0_3 ), .A2(\SB3_11/i1[9] ), .A3(\SB3_11/i0[6] ), .ZN(\SB3_11/Component_Function_3/NAND4_in[0] ) );
  BUF_X2 \SB4_1/BUF_0  ( .I(\SB3_6/buf_output[0] ), .Z(\SB4_1/i0[9] ) );
  BUF_X2 \SB4_17/BUF_1  ( .I(\SB3_21/buf_output[1] ), .Z(\SB4_17/i0[6] ) );
  BUF_X2 U1455 ( .I(\SB3_7/buf_output[0] ), .Z(\SB4_2/i0[9] ) );
  NAND2_X1 \SB4_29/Component_Function_1/N1  ( .A1(\SB4_29/i0_3 ), .A2(
        \SB4_29/i1[9] ), .ZN(\SB4_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U5179 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i1_7 ), .A3(
        \SB4_29/i1[9] ), .ZN(n3067) );
  NAND3_X1 U4500 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i1_5 ), .A3(
        \SB4_16/i1[9] ), .ZN(n1321) );
  NAND3_X1 U39 ( .A1(\SB4_16/i0_4 ), .A2(\SB4_16/i1_7 ), .A3(\SB4_16/i0[8] ), 
        .ZN(\SB4_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U47 ( .A1(\SB4_1/i0[10] ), .A2(\SB4_1/i1[9] ), .A3(\SB4_1/i1_7 ), 
        .ZN(n5065) );
  NAND2_X1 U613 ( .A1(\SB3_2/i0[9] ), .A2(\SB3_2/i0[10] ), .ZN(
        \SB3_2/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U620 ( .A1(\SB3_17/i0_0 ), .A2(\SB3_17/i3[0] ), .ZN(
        \SB3_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U626 ( .A1(\SB3_5/i0_0 ), .A2(\SB3_5/i0_3 ), .A3(\SB3_5/i0_4 ), 
        .ZN(\SB3_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U628 ( .A1(\SB3_21/i0[6] ), .A2(\SB3_21/i0_4 ), .A3(\SB3_21/i0[9] ), 
        .ZN(n4393) );
  NAND2_X1 U629 ( .A1(\SB3_13/i0_0 ), .A2(\SB3_13/i3[0] ), .ZN(
        \SB3_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U632 ( .A1(\SB3_27/i0[8] ), .A2(\SB3_27/i1_5 ), .A3(\SB3_27/i3[0] ), 
        .ZN(\SB3_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U633 ( .A1(\SB3_5/i0[8] ), .A2(\SB3_5/i0[7] ), .A3(\SB3_5/i0[6] ), 
        .ZN(\SB3_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U634 ( .A1(\SB3_12/i1_5 ), .A2(\SB3_12/i0_4 ), .A3(\SB3_12/i1[9] ), 
        .ZN(n1781) );
  NAND3_X1 U651 ( .A1(\RI1[5][113] ), .A2(\SB3_13/i1[9] ), .A3(\SB3_13/i0[6] ), 
        .ZN(\SB3_13/Component_Function_3/NAND4_in[0] ) );
  BUF_X2 U656 ( .I(\MC_ARK_ARC_1_4/buf_output[158] ), .Z(\SB3_5/i0_0 ) );
  BUF_X2 U666 ( .I(\MC_ARK_ARC_1_4/buf_output[55] ), .Z(\SB3_22/i0[6] ) );
  NAND2_X1 U674 ( .A1(\SB2_4_18/i0_3 ), .A2(\SB2_4_18/i1[9] ), .ZN(n3765) );
  NAND3_X1 U687 ( .A1(\SB2_4_13/i0_3 ), .A2(\SB2_4_13/i0_0 ), .A3(
        \SB2_4_13/i0_4 ), .ZN(\SB2_4_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U691 ( .A1(\SB2_4_2/i0_3 ), .A2(\SB2_4_2/i0[8] ), .A3(
        \SB2_4_2/i1_7 ), .ZN(\SB2_4_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U705 ( .A1(\SB2_4_4/i0_0 ), .A2(n3178), .ZN(n4269) );
  NAND3_X1 U708 ( .A1(\SB2_4_12/i0_0 ), .A2(\SB1_4_13/buf_output[4] ), .A3(
        \SB2_4_12/i1_5 ), .ZN(n3922) );
  NAND3_X1 U724 ( .A1(\SB2_4_10/i1[9] ), .A2(\SB2_4_10/i0_3 ), .A3(
        \SB2_4_10/i0[6] ), .ZN(\SB2_4_10/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U733 ( .A1(\SB2_4_8/i0_0 ), .A2(\SB2_4_8/i3[0] ), .ZN(n4692) );
  NAND3_X1 U735 ( .A1(\SB2_4_1/i1_7 ), .A2(\SB2_4_1/i0[8] ), .A3(
        \SB2_4_1/i0_4 ), .ZN(n3808) );
  NAND3_X1 U749 ( .A1(\SB2_4_3/i0_0 ), .A2(\SB2_4_3/i0[7] ), .A3(
        \SB2_4_3/i0_3 ), .ZN(n4985) );
  NAND3_X1 U752 ( .A1(\SB2_4_14/i0[9] ), .A2(\SB2_4_14/i0_3 ), .A3(
        \SB2_4_14/i0[10] ), .ZN(n5364) );
  INV_X1 U760 ( .I(\SB1_4_19/buf_output[1] ), .ZN(\SB2_4_15/i1_7 ) );
  INV_X1 U771 ( .I(\SB1_4_17/buf_output[1] ), .ZN(\SB2_4_13/i1_7 ) );
  INV_X1 U776 ( .I(\SB1_4_17/buf_output[0] ), .ZN(\SB2_4_12/i3[0] ) );
  NAND3_X1 U784 ( .A1(\SB1_4_13/i0_4 ), .A2(\SB1_4_13/i0[8] ), .A3(
        \SB1_4_13/i1_7 ), .ZN(n4641) );
  NAND3_X1 U792 ( .A1(\SB1_4_14/i0_4 ), .A2(\SB1_4_14/i0_3 ), .A3(
        \SB1_4_14/i1[9] ), .ZN(\SB1_4_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U827 ( .A1(\SB1_4_20/i0[9] ), .A2(\SB1_4_20/i1_5 ), .A3(
        \SB1_4_20/i0[6] ), .ZN(\SB1_4_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U831 ( .A1(\SB1_4_13/i0[10] ), .A2(\SB1_4_13/i1[9] ), .A3(
        \SB1_4_13/i1_7 ), .ZN(n4360) );
  NAND3_X1 U839 ( .A1(\SB1_4_15/i0_4 ), .A2(\SB1_4_15/i1_7 ), .A3(
        \SB1_4_15/i0[8] ), .ZN(n5306) );
  NAND3_X1 U864 ( .A1(\SB1_4_30/i0_3 ), .A2(\SB1_4_30/i0_4 ), .A3(
        \SB1_4_30/i0_0 ), .ZN(\SB1_4_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U870 ( .A1(\SB1_4_13/i0_0 ), .A2(\SB1_4_13/i0[10] ), .A3(
        \SB1_4_13/i0[6] ), .ZN(\SB1_4_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U872 ( .A1(\SB1_4_2/i0_0 ), .A2(\SB1_4_2/i1_7 ), .A3(
        \SB1_4_2/i3[0] ), .ZN(n5046) );
  NAND3_X1 U874 ( .A1(\SB1_4_4/i0[10] ), .A2(\SB1_4_4/i0_3 ), .A3(
        \SB1_4_4/i0_4 ), .ZN(n3661) );
  NAND3_X1 U903 ( .A1(\SB1_4_3/i0[9] ), .A2(\SB1_4_3/i1_5 ), .A3(
        \SB1_4_3/i0[6] ), .ZN(n4483) );
  NAND2_X1 U906 ( .A1(\SB1_4_12/i0_0 ), .A2(\SB1_4_12/i3[0] ), .ZN(
        \SB1_4_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U912 ( .A1(\SB1_4_2/i0[10] ), .A2(\SB1_4_2/i1[9] ), .A3(
        \SB1_4_2/i1_7 ), .ZN(\SB1_4_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U915 ( .A1(\SB1_4_23/i0_0 ), .A2(\SB1_4_23/i0_3 ), .A3(
        \SB1_4_23/i0[7] ), .ZN(n3847) );
  INV_X2 U927 ( .I(\SB1_4_30/i0_4 ), .ZN(\SB1_4_30/i0[7] ) );
  NAND3_X1 U935 ( .A1(\SB1_4_21/i0_3 ), .A2(\SB1_4_21/i0[9] ), .A3(
        \SB1_4_21/i0[8] ), .ZN(n4376) );
  INV_X1 U958 ( .I(\MC_ARK_ARC_1_3/buf_output[172] ), .ZN(\SB1_4_3/i0[7] ) );
  BUF_X2 U963 ( .I(\MC_ARK_ARC_1_3/buf_output[97] ), .Z(\SB1_4_15/i0[6] ) );
  INV_X1 U968 ( .I(\MC_ARK_ARC_1_3/buf_output[78] ), .ZN(\SB1_4_18/i3[0] ) );
  NAND2_X1 U979 ( .A1(\SB2_3_11/i0_3 ), .A2(\SB2_3_11/i1[9] ), .ZN(
        \SB2_3_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U993 ( .A1(\SB2_3_18/i0[10] ), .A2(\SB2_3_18/i1_5 ), .A3(
        \SB2_3_18/i1[9] ), .ZN(\SB2_3_18/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U1012 ( .A1(\SB2_3_2/i0[9] ), .A2(\SB2_3_2/i0[10] ), .ZN(n4333) );
  NAND3_X1 U1040 ( .A1(\SB2_3_11/i0_3 ), .A2(\SB2_3_11/i1_7 ), .A3(
        \SB2_3_11/i0[8] ), .ZN(n4643) );
  NAND3_X1 U1048 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i0[10] ), .A3(
        \SB2_3_23/i0[9] ), .ZN(n2996) );
  NAND3_X1 U1094 ( .A1(\SB2_3_29/i0[9] ), .A2(\SB2_3_29/i0[10] ), .A3(
        \SB2_3_29/i0_3 ), .ZN(n4027) );
  NAND3_X1 U1107 ( .A1(n6552), .A2(\SB2_3_29/i0[9] ), .A3(\SB2_3_29/i1_5 ), 
        .ZN(n4793) );
  INV_X1 U1119 ( .I(\SB1_3_4/buf_output[1] ), .ZN(\SB2_3_0/i1_7 ) );
  NAND3_X1 U1173 ( .A1(\SB1_3_24/i0_4 ), .A2(\SB1_3_24/i0_0 ), .A3(
        \SB1_3_24/i1_5 ), .ZN(n3770) );
  NAND2_X1 U1187 ( .A1(\SB1_3_29/Component_Function_4/NAND4_in[2] ), .A2(n4912), .ZN(n4524) );
  NAND3_X1 U1197 ( .A1(\SB1_3_15/i0[9] ), .A2(\SB1_3_15/i0_4 ), .A3(
        \SB1_3_15/i0[6] ), .ZN(n1537) );
  NAND3_X1 U1209 ( .A1(\SB1_3_1/i0_3 ), .A2(\SB1_3_1/i0_4 ), .A3(
        \SB1_3_1/i1[9] ), .ZN(\SB1_3_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1215 ( .A1(\SB1_3_2/i0_4 ), .A2(\SB1_3_2/i0[8] ), .A3(
        \SB1_3_2/i1_7 ), .ZN(n4756) );
  NAND2_X1 U1258 ( .A1(n4499), .A2(n4444), .ZN(n4610) );
  NAND3_X1 U1264 ( .A1(\SB1_3_10/i0[9] ), .A2(\SB1_3_10/i0[6] ), .A3(
        \SB1_3_10/i1_5 ), .ZN(n3935) );
  NAND3_X1 U1267 ( .A1(\SB1_3_13/i0[10] ), .A2(\SB1_3_13/i1[9] ), .A3(
        \SB1_3_13/i1_7 ), .ZN(n4770) );
  NAND3_X1 U1271 ( .A1(\SB1_3_10/i0[9] ), .A2(\SB1_3_10/i0_3 ), .A3(
        \SB1_3_10/i0[8] ), .ZN(n4855) );
  NAND3_X1 U1299 ( .A1(\SB1_3_21/i0[8] ), .A2(\SB1_3_21/i1_5 ), .A3(
        \SB1_3_21/i3[0] ), .ZN(\SB1_3_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1302 ( .A1(\SB1_3_24/i0[8] ), .A2(\SB1_3_24/i1_5 ), .A3(
        \SB1_3_24/i3[0] ), .ZN(\SB1_3_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1303 ( .A1(\SB1_3_26/i0[8] ), .A2(\SB1_3_26/i3[0] ), .A3(
        \SB1_3_26/i1_5 ), .ZN(n3365) );
  NAND3_X1 U1315 ( .A1(\SB1_3_27/i0[9] ), .A2(\SB1_3_27/i0_0 ), .A3(
        \SB1_3_27/i0[8] ), .ZN(n3919) );
  NAND3_X1 U1320 ( .A1(\SB1_3_27/i0[10] ), .A2(\SB1_3_27/i0_3 ), .A3(
        \SB1_3_27/i0[9] ), .ZN(n4499) );
  INV_X1 U1322 ( .I(\MC_ARK_ARC_1_2/buf_output[77] ), .ZN(\SB1_3_19/i1_5 ) );
  NAND3_X1 U1329 ( .A1(\SB1_3_10/i0[9] ), .A2(\SB1_3_10/i0_3 ), .A3(
        \SB1_3_10/i0[10] ), .ZN(n4937) );
  NAND3_X1 U1339 ( .A1(\SB1_3_1/i0[10] ), .A2(\SB1_3_1/i1[9] ), .A3(
        \SB1_3_1/i1_7 ), .ZN(\SB1_3_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1340 ( .A1(\SB1_3_27/i0_4 ), .A2(\SB1_3_27/i1[9] ), .A3(
        \SB1_3_27/i1_5 ), .ZN(n4444) );
  NAND3_X1 U1342 ( .A1(\SB1_3_22/i0[10] ), .A2(\SB1_3_22/i1[9] ), .A3(
        \SB1_3_22/i1_7 ), .ZN(\SB1_3_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1350 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i3[0] ), .A3(
        \SB1_3_27/i1_7 ), .ZN(n5218) );
  NAND3_X1 U1351 ( .A1(\SB1_3_11/i0_0 ), .A2(\SB1_3_11/i1_7 ), .A3(
        \SB1_3_11/i3[0] ), .ZN(n5160) );
  NAND3_X1 U1389 ( .A1(\SB2_2_2/i0_3 ), .A2(\SB2_2_2/i0[10] ), .A3(
        \SB2_2_2/i0[9] ), .ZN(n3912) );
  NAND3_X1 U1407 ( .A1(\SB2_2_3/i0[10] ), .A2(\SB2_2_3/i0_3 ), .A3(
        \SB2_2_3/i0[9] ), .ZN(n5208) );
  NAND3_X1 U1411 ( .A1(\SB2_2_20/i0_4 ), .A2(\SB2_2_20/i0_0 ), .A3(
        \SB2_2_20/i1_5 ), .ZN(n4901) );
  NAND3_X1 U1415 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0[8] ), .A3(
        \SB2_2_22/i1_7 ), .ZN(\SB2_2_22/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1416 ( .A1(\SB2_2_29/i0_0 ), .A2(\SB2_2_29/i3[0] ), .A3(
        \SB2_2_29/i1_7 ), .ZN(n3819) );
  NAND3_X1 U1422 ( .A1(\SB2_2_11/i0_0 ), .A2(\SB2_2_11/i0_3 ), .A3(
        \SB2_2_11/i0_4 ), .ZN(n5166) );
  NAND3_X1 U1425 ( .A1(\SB2_2_30/i0[10] ), .A2(\SB2_2_30/i0_3 ), .A3(
        \SB2_2_30/i0_4 ), .ZN(n4509) );
  NAND3_X1 U1432 ( .A1(\SB2_2_29/i0_0 ), .A2(\SB1_2_30/buf_output[4] ), .A3(
        \SB2_2_29/i1_5 ), .ZN(n3864) );
  NAND3_X1 U1445 ( .A1(\SB2_2_9/i0_0 ), .A2(\SB2_2_9/i0_3 ), .A3(
        \SB2_2_9/i0[7] ), .ZN(n5072) );
  NAND3_X1 U1450 ( .A1(\SB2_2_11/i0_3 ), .A2(\SB2_2_11/i0[6] ), .A3(
        \SB2_2_11/i1[9] ), .ZN(n3875) );
  AOI21_X1 U1461 ( .A1(\SB2_2_9/i0_0 ), .A2(n4180), .B(\SB2_2_9/i1_5 ), .ZN(
        n4249) );
  NAND3_X1 U1478 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0[10] ), .A3(
        \SB2_2_4/i0[9] ), .ZN(\SB2_2_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1479 ( .A1(\SB2_2_31/i0_0 ), .A2(\SB2_2_31/i0_3 ), .A3(
        \SB2_2_31/i0[7] ), .ZN(n1481) );
  NAND3_X1 U1508 ( .A1(\SB1_2_28/i0_3 ), .A2(\SB1_2_28/i1[9] ), .A3(
        \SB1_2_28/i0[6] ), .ZN(\SB1_2_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1528 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i0[10] ), .A3(
        \SB1_2_18/i0[9] ), .ZN(n4111) );
  NAND3_X1 U1531 ( .A1(\SB1_2_9/i0[10] ), .A2(\SB1_2_9/i1[9] ), .A3(
        \SB1_2_9/i1_5 ), .ZN(n3548) );
  NAND3_X1 U1541 ( .A1(\SB1_2_3/i0[9] ), .A2(\SB1_2_3/i0[10] ), .A3(
        \SB1_2_3/i0_3 ), .ZN(\SB1_2_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1542 ( .A1(\RI1[2][191] ), .A2(\SB1_2_0/i0[9] ), .A3(
        \SB1_2_0/i0[10] ), .ZN(\SB1_2_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1551 ( .A1(\SB1_2_20/i0[8] ), .A2(\SB1_2_20/i1_5 ), .A3(
        \SB1_2_20/i3[0] ), .ZN(n3626) );
  NAND3_X1 U1604 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i0[10] ), .A3(
        \SB1_2_18/i0[6] ), .ZN(n4390) );
  NAND3_X1 U1605 ( .A1(\SB1_2_23/i0_3 ), .A2(\SB1_2_23/i0_4 ), .A3(
        \SB1_2_23/i1[9] ), .ZN(n4604) );
  NAND3_X1 U1606 ( .A1(n3184), .A2(\SB1_2_7/i0[9] ), .A3(\RI1[2][149] ), .ZN(
        n5101) );
  NAND3_X1 U1612 ( .A1(\SB1_2_30/i0_4 ), .A2(\SB1_2_30/i1[9] ), .A3(
        \SB1_2_30/i0_3 ), .ZN(\SB1_2_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1635 ( .A1(\SB2_1_22/i0[10] ), .A2(\SB2_1_22/i0[6] ), .A3(
        \SB2_1_22/i0_3 ), .ZN(\SB2_1_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1656 ( .A1(\SB2_1_16/i0_0 ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i0[7] ), .ZN(\SB2_1_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1659 ( .A1(\SB2_1_17/i0_3 ), .A2(\SB2_1_17/i0[10] ), .A3(
        \SB2_1_17/i0_4 ), .ZN(n5287) );
  NAND3_X1 U1661 ( .A1(\SB2_1_31/i0[10] ), .A2(\SB2_1_31/i0[9] ), .A3(
        \SB2_1_31/i0_3 ), .ZN(n4460) );
  NAND3_X1 U1689 ( .A1(\SB2_1_17/i0_4 ), .A2(\SB2_1_17/i0[6] ), .A3(
        \SB2_1_17/i0[9] ), .ZN(n5418) );
  NAND3_X1 U1698 ( .A1(\SB1_1_25/i0[10] ), .A2(\SB1_1_25/i0_3 ), .A3(
        \SB1_1_25/i0_4 ), .ZN(\SB1_1_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1710 ( .A1(\SB1_1_4/i0_3 ), .A2(\SB1_1_4/i0[8] ), .A3(
        \SB1_1_4/i1_7 ), .ZN(\SB1_1_4/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1715 ( .A1(\SB1_1_3/i0_4 ), .A2(\SB1_1_3/i0[8] ), .A3(
        \SB1_1_3/i1_7 ), .ZN(n1375) );
  NAND3_X1 U1717 ( .A1(\SB1_1_7/i0_4 ), .A2(\SB1_1_7/i0[6] ), .A3(
        \SB1_1_7/i0[9] ), .ZN(n4563) );
  NAND3_X1 U1726 ( .A1(\SB1_1_7/i1_5 ), .A2(\SB1_1_7/i0[6] ), .A3(
        \SB1_1_7/i0[9] ), .ZN(\SB1_1_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1743 ( .A1(\SB1_1_27/i0[6] ), .A2(\SB1_1_27/i0_3 ), .A3(
        \SB1_1_27/i0[10] ), .ZN(n5350) );
  NAND3_X1 U1754 ( .A1(\SB1_1_6/i0[10] ), .A2(\SB1_1_6/i1[9] ), .A3(
        \SB1_1_6/i1_5 ), .ZN(n4744) );
  NAND3_X1 U1764 ( .A1(\SB1_1_11/i0_4 ), .A2(\SB1_1_11/i1_7 ), .A3(
        \SB1_1_11/i0[8] ), .ZN(n3721) );
  NAND3_X1 U1772 ( .A1(\SB1_1_1/i0[10] ), .A2(\SB1_1_1/i1_7 ), .A3(
        \SB1_1_1/i1[9] ), .ZN(\SB1_1_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1784 ( .A1(\SB1_1_10/i0[8] ), .A2(\SB1_1_10/i1_5 ), .A3(
        \SB1_1_10/i3[0] ), .ZN(n5309) );
  NAND3_X1 U1787 ( .A1(\SB1_1_23/i0_4 ), .A2(\SB1_1_23/i0[8] ), .A3(
        \SB1_1_23/i1_7 ), .ZN(n2261) );
  NAND3_X1 U1792 ( .A1(\SB1_1_1/i0[10] ), .A2(\SB1_1_1/i0_3 ), .A3(
        \SB1_1_1/i0_4 ), .ZN(\SB1_1_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1813 ( .A1(\SB1_1_7/i0_0 ), .A2(\SB1_1_7/i0[9] ), .A3(
        \SB1_1_7/i0[8] ), .ZN(\SB1_1_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1814 ( .A1(\SB1_1_4/i0[10] ), .A2(\SB1_1_4/i1[9] ), .A3(
        \SB1_1_4/i1_7 ), .ZN(n3487) );
  NAND3_X1 U1820 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i0_0 ), .A3(
        \SB1_1_14/i0_4 ), .ZN(\SB1_1_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1834 ( .A1(\SB1_1_1/i0[10] ), .A2(\SB1_1_1/i0_0 ), .A3(
        \SB1_1_1/i0[6] ), .ZN(n4950) );
  NAND3_X1 U1845 ( .A1(\SB1_1_23/i0[6] ), .A2(\MC_ARK_ARC_1_0/buf_output[52] ), 
        .A3(\SB1_1_23/i0[9] ), .ZN(n3645) );
  NAND3_X1 U1865 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0[9] ), .A3(
        \SB1_1_22/i0[10] ), .ZN(n4763) );
  NAND3_X1 U1877 ( .A1(\SB1_1_6/i0_0 ), .A2(\SB1_1_6/i0_3 ), .A3(
        \SB1_1_6/i0[7] ), .ZN(n3927) );
  NAND3_X1 U1893 ( .A1(\SB1_1_6/i0[10] ), .A2(\SB1_1_6/i0_3 ), .A3(
        \SB1_1_6/i0_4 ), .ZN(n3928) );
  NAND3_X1 U1922 ( .A1(\SB2_0_3/i0[10] ), .A2(\SB2_0_3/i0[6] ), .A3(
        \SB2_0_3/i0_3 ), .ZN(\SB2_0_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1927 ( .A1(\SB2_0_3/i0_3 ), .A2(\SB1_0_8/buf_output[0] ), .A3(
        \SB2_0_3/i0[8] ), .ZN(\SB2_0_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1931 ( .A1(\RI3[0][1] ), .A2(\RI3[0][3] ), .A3(\SB2_0_31/i0_3 ), 
        .ZN(\SB2_0_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1935 ( .A1(\RI3[0][166] ), .A2(\SB2_0_4/i1_5 ), .A3(\SB2_0_4/i0_0 ), .ZN(n5248) );
  NAND3_X1 U1936 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0[8] ), .A3(
        \SB2_0_5/i1_7 ), .ZN(\SB2_0_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1937 ( .A1(\SB2_0_18/i0[10] ), .A2(\SB2_0_18/i1_7 ), .A3(
        \SB2_0_18/i1[9] ), .ZN(n2333) );
  NAND3_X1 U1943 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i1[9] ), .A3(
        \SB2_0_4/i1_7 ), .ZN(\SB2_0_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1964 ( .A1(\SB2_0_1/i0_3 ), .A2(\SB2_0_1/i0[9] ), .A3(
        \SB2_0_1/i0[8] ), .ZN(n3465) );
  NAND3_X1 U1965 ( .A1(\SB2_0_10/i1[9] ), .A2(\SB2_0_10/i0_4 ), .A3(
        \SB2_0_10/i1_5 ), .ZN(n5018) );
  NAND3_X1 U1971 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i0_0 ), .A3(
        \RI3[0][163] ), .ZN(\SB2_0_4/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1976 ( .A1(\SB2_0_5/i0[10] ), .A2(\SB2_0_5/i0_0 ), .A3(
        \SB1_0_9/buf_output[1] ), .ZN(
        \SB2_0_5/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1988 ( .A1(\SB2_0_24/i1_5 ), .A2(\SB2_0_24/i0_0 ), .A3(
        \RI3[0][46] ), .ZN(\SB2_0_24/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1989 ( .A1(\SB2_0_1/i0_4 ), .A2(\SB2_0_1/i1_7 ), .A3(
        \SB2_0_1/i0[8] ), .ZN(n4835) );
  NAND3_X1 U2003 ( .A1(\SB2_0_1/i0[10] ), .A2(\SB2_0_1/i0[9] ), .A3(
        \SB2_0_1/i0_3 ), .ZN(\SB2_0_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2044 ( .A1(\SB1_0_7/i0[6] ), .A2(\SB1_0_7/i0[9] ), .A3(
        \SB1_0_7/i0_4 ), .ZN(n4780) );
  NAND3_X1 U2048 ( .A1(\SB1_0_14/i0_3 ), .A2(\SB1_0_14/i0[6] ), .A3(
        \SB1_0_14/i1[9] ), .ZN(n4377) );
  NAND3_X1 U2052 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0[10] ), .A3(
        \SB1_0_21/i0[9] ), .ZN(n1233) );
  NAND3_X1 U2059 ( .A1(\SB1_0_26/i0[9] ), .A2(\SB1_0_26/i0_3 ), .A3(
        \SB1_0_26/i0[8] ), .ZN(n4954) );
  NAND3_X1 U2061 ( .A1(\SB1_0_2/i0_4 ), .A2(\SB1_0_2/i0[8] ), .A3(
        \SB1_0_2/i1_7 ), .ZN(n1519) );
  NAND3_X1 U2065 ( .A1(\SB1_0_12/i0[10] ), .A2(\SB1_0_12/i1_7 ), .A3(
        \SB1_0_12/i1[9] ), .ZN(n4748) );
  NAND3_X1 U2073 ( .A1(\SB1_0_31/i0_3 ), .A2(\SB1_0_31/i0[6] ), .A3(
        \SB1_0_31/i1[9] ), .ZN(n4881) );
  NAND3_X1 U2095 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i0_0 ), .A3(
        \SB1_0_29/i0[7] ), .ZN(\SB1_0_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2104 ( .A1(\SB1_0_14/i0_3 ), .A2(\SB1_0_14/i0[10] ), .A3(
        \SB1_0_14/i0[9] ), .ZN(n4221) );
  NAND3_X1 U2128 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0[8] ), .A3(
        \SB1_0_18/i1_7 ), .ZN(n3939) );
  NOR2_X1 U2135 ( .A1(n3434), .A2(n3435), .ZN(n3286) );
  NAND3_X1 U2140 ( .A1(\SB1_0_14/i0_4 ), .A2(\SB1_0_14/i0[10] ), .A3(
        \SB1_0_14/i0_3 ), .ZN(n1460) );
  INV_X2 U2144 ( .I(\MC_ARK_ARC_1_2/buf_output[35] ), .ZN(\SB1_3_26/i1_5 ) );
  NAND2_X1 U2146 ( .A1(\SB1_3_23/Component_Function_4/NAND4_in[3] ), .A2(n3187), .ZN(n2521) );
  INV_X2 U2159 ( .I(\MC_ARK_ARC_1_0/buf_output[59] ), .ZN(\SB1_1_22/i1_5 ) );
  INV_X4 U2163 ( .I(n3370), .ZN(\SB2_4_1/i0_4 ) );
  NAND3_X2 U2165 ( .A1(\SB2_4_0/i0[9] ), .A2(\SB2_4_0/i0[6] ), .A3(
        \SB1_4_1/buf_output[4] ), .ZN(n1262) );
  NAND3_X2 U2185 ( .A1(\SB1_3_17/i0[10] ), .A2(\SB1_3_17/i0[6] ), .A3(
        \SB1_3_17/i0_0 ), .ZN(\SB1_3_17/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U2193 ( .A1(\SB2_4_20/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_20/Component_Function_0/NAND4_in[3] ), .A3(n1195), .A4(
        \SB2_4_20/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_4_20/buf_output[0] ) );
  NAND3_X2 U2204 ( .A1(\SB1_3_26/i0[10] ), .A2(\SB1_3_26/i0_0 ), .A3(
        \SB1_3_26/i0[6] ), .ZN(n4009) );
  INV_X2 U2208 ( .I(\MC_ARK_ARC_1_1/buf_output[109] ), .ZN(\SB1_2_13/i1_7 ) );
  BUF_X4 U2209 ( .I(\MC_ARK_ARC_1_2/buf_output[119] ), .Z(\SB1_3_12/i0_3 ) );
  BUF_X4 U2264 ( .I(\MC_ARK_ARC_1_0/buf_output[83] ), .Z(\SB1_1_18/i0_3 ) );
  INV_X2 U2269 ( .I(\MC_ARK_ARC_1_2/buf_output[8] ), .ZN(\SB1_3_30/i1[9] ) );
  BUF_X4 U2303 ( .I(n411), .Z(\SB1_0_1/i0_3 ) );
  NAND3_X2 U2311 ( .A1(\SB1_1_29/i0_4 ), .A2(\SB1_1_29/i0[8] ), .A3(
        \SB1_1_29/i1_7 ), .ZN(\SB1_1_29/Component_Function_1/NAND4_in[3] ) );
  NAND2_X2 U2325 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i1[9] ), .ZN(
        \SB1_1_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U2328 ( .A1(\SB1_3_27/i0[7] ), .A2(\SB1_3_27/i0[8] ), .A3(
        \SB1_3_27/i0[6] ), .ZN(n4279) );
  INV_X2 U2330 ( .I(\MC_ARK_ARC_1_2/buf_output[119] ), .ZN(\SB1_3_12/i1_5 ) );
  BUF_X2 U2341 ( .I(\SB3_31/buf_output[2] ), .Z(\SB4_28/i0_0 ) );
  NAND3_X1 U2343 ( .A1(\SB3_22/i1[9] ), .A2(\SB3_22/i0_4 ), .A3(\SB3_22/i0_3 ), 
        .ZN(\SB3_22/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2345 ( .A1(\SB3_22/i0_0 ), .A2(\SB3_22/i0_3 ), .A3(\SB3_22/i0_4 ), 
        .ZN(\SB3_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2359 ( .A1(\SB2_4_8/i0[7] ), .A2(\SB2_4_8/i0[8] ), .A3(
        \SB2_4_8/i0[6] ), .ZN(n4684) );
  NAND3_X1 U2367 ( .A1(\SB1_4_27/i0[9] ), .A2(\SB1_4_27/i1_5 ), .A3(
        \SB1_4_27/i0[6] ), .ZN(\SB1_4_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2370 ( .A1(\SB1_4_27/i0[9] ), .A2(\SB1_4_27/i0[10] ), .A3(
        \SB1_4_27/i0_3 ), .ZN(\SB1_4_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2383 ( .A1(\SB2_4_24/i0_3 ), .A2(\SB2_4_24/i1_7 ), .A3(
        \SB2_4_24/i0[8] ), .ZN(\SB2_4_24/Component_Function_1/NAND4_in[1] ) );
  INV_X1 U2385 ( .I(\SB1_3_31/buf_output[1] ), .ZN(\SB2_3_27/i1_7 ) );
  INV_X1 U2387 ( .I(\MC_ARK_ARC_1_4/buf_output[164] ), .ZN(\SB3_4/i1[9] ) );
  BUF_X2 U2388 ( .I(\MC_ARK_ARC_1_4/buf_output[164] ), .Z(\SB3_4/i0_0 ) );
  NAND3_X1 U2389 ( .A1(\SB3_10/i0_3 ), .A2(\SB3_10/i0[9] ), .A3(
        \SB3_10/i0[10] ), .ZN(n5307) );
  BUF_X2 U2404 ( .I(n294), .Z(\SB1_0_11/i0_0 ) );
  INV_X1 U2408 ( .I(n294), .ZN(\SB1_0_11/i1[9] ) );
  NAND2_X1 U2410 ( .A1(\SB3_7/i0_0 ), .A2(\SB3_7/i3[0] ), .ZN(
        \SB3_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2412 ( .A1(\SB3_7/i1_5 ), .A2(\SB3_7/i0_0 ), .A3(\SB3_7/i0_4 ), 
        .ZN(\SB3_7/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 U2421 ( .A1(\SB3_10/i0_0 ), .A2(\SB3_10/i3[0] ), .ZN(
        \SB3_10/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U2422 ( .I(\MC_ARK_ARC_1_4/buf_output[157] ), .ZN(\SB3_5/i1_7 ) );
  BUF_X2 U2423 ( .I(\MC_ARK_ARC_1_4/buf_output[157] ), .Z(\SB3_5/i0[6] ) );
  INV_X1 U2426 ( .I(\SB3_8/buf_output[2] ), .ZN(\SB4_5/i1[9] ) );
  BUF_X2 U2432 ( .I(\SB3_8/buf_output[2] ), .Z(\SB4_5/i0_0 ) );
  BUF_X2 U2434 ( .I(\SB3_16/buf_output[3] ), .Z(\SB4_14/i0[10] ) );
  NAND3_X1 U2444 ( .A1(\SB3_26/i0_0 ), .A2(\SB3_26/i0_3 ), .A3(\SB3_26/i0[7] ), 
        .ZN(n5081) );
  NAND3_X1 U2453 ( .A1(\SB3_4/i1_5 ), .A2(\SB3_4/i0_0 ), .A3(\SB3_4/i0_4 ), 
        .ZN(\SB3_4/Component_Function_2/NAND4_in[3] ) );
  BUF_X2 U2459 ( .I(\MC_ARK_ARC_1_4/buf_output[127] ), .Z(\SB3_10/i0[6] ) );
  NAND3_X1 U2461 ( .A1(\SB3_10/i1_5 ), .A2(\SB3_10/i0[10] ), .A3(
        \SB3_10/i1[9] ), .ZN(\SB3_10/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U2466 ( .I(\MC_ARK_ARC_1_4/buf_output[129] ), .ZN(\SB3_10/i0[8] ) );
  BUF_X2 U2467 ( .I(\MC_ARK_ARC_1_4/buf_output[129] ), .Z(\SB3_10/i0[10] ) );
  CLKBUF_X4 U2468 ( .I(\SB3_5/buf_output[4] ), .Z(\SB4_4/i0_4 ) );
  NAND3_X1 U2472 ( .A1(\SB2_3_23/i1_5 ), .A2(\SB2_3_23/i0[8] ), .A3(
        \SB2_3_23/i3[0] ), .ZN(\SB2_3_23/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U2474 ( .I(\SB3_15/buf_output[1] ), .ZN(\SB4_11/i1_7 ) );
  BUF_X2 U2475 ( .I(\SB3_15/buf_output[1] ), .Z(\SB4_11/i0[6] ) );
  NAND3_X1 U2476 ( .A1(\SB3_26/i0_4 ), .A2(\SB3_26/i1[9] ), .A3(\SB3_26/i0_3 ), 
        .ZN(n886) );
  BUF_X2 U2479 ( .I(\SB3_12/buf_output[0] ), .Z(\SB4_7/i0[9] ) );
  NAND3_X1 U2493 ( .A1(\SB3_24/i0_3 ), .A2(\SB3_24/i1[9] ), .A3(\SB3_24/i0_4 ), 
        .ZN(n966) );
  NAND3_X1 U2495 ( .A1(\SB3_24/i0_3 ), .A2(\SB3_24/i0[8] ), .A3(\SB3_24/i0[9] ), .ZN(\SB3_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2496 ( .A1(\SB3_24/i0_3 ), .A2(\SB3_24/i0[9] ), .A3(
        \SB3_24/i0[10] ), .ZN(n5305) );
  NAND3_X1 U2501 ( .A1(\SB3_24/i0_0 ), .A2(\SB3_24/i0_3 ), .A3(\SB3_24/i0_4 ), 
        .ZN(\SB3_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2504 ( .A1(\SB3_24/i0_3 ), .A2(\SB3_24/i0[10] ), .A3(
        \SB3_24/i0[6] ), .ZN(\SB3_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2509 ( .A1(\SB3_24/i0[6] ), .A2(\SB3_24/i0_3 ), .A3(\SB3_24/i1[9] ), .ZN(n3804) );
  NAND3_X1 U2511 ( .A1(\SB3_7/i1[9] ), .A2(\SB3_7/i0_4 ), .A3(n6270), .ZN(
        \SB3_7/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U2519 ( .I(\MC_ARK_ARC_1_4/buf_output[128] ), .ZN(\SB3_10/i1[9] ) );
  BUF_X2 U2520 ( .I(\MC_ARK_ARC_1_4/buf_output[128] ), .Z(\SB3_10/i0_0 ) );
  INV_X1 U2530 ( .I(\SB3_27/buf_output[1] ), .ZN(\SB4_23/i1_7 ) );
  NAND3_X1 U2542 ( .A1(\SB3_3/i0[8] ), .A2(\SB3_3/i0[7] ), .A3(\SB3_3/i0[6] ), 
        .ZN(\SB3_3/Component_Function_0/NAND4_in[1] ) );
  INV_X1 U2553 ( .I(\MC_ARK_ARC_1_4/buf_output[61] ), .ZN(\SB3_21/i1_7 ) );
  BUF_X2 U2555 ( .I(\MC_ARK_ARC_1_4/buf_output[61] ), .Z(\SB3_21/i0[6] ) );
  NAND3_X1 U2560 ( .A1(\SB3_18/i1_5 ), .A2(\SB3_18/i0[8] ), .A3(\SB3_18/i3[0] ), .ZN(n5138) );
  BUF_X2 U2568 ( .I(\MC_ARK_ARC_1_4/buf_output[139] ), .Z(\SB3_8/i0[6] ) );
  NAND3_X1 U2572 ( .A1(\SB4_15/i0_3 ), .A2(n1497), .A3(\SB4_15/i0[9] ), .ZN(
        \SB4_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2575 ( .A1(\SB1_4_28/i0_3 ), .A2(\SB1_4_28/i1_7 ), .A3(
        \SB1_4_28/i0[8] ), .ZN(\SB1_4_28/Component_Function_1/NAND4_in[1] ) );
  INV_X1 U2590 ( .I(\MC_ARK_ARC_1_3/buf_output[7] ), .ZN(\SB1_4_30/i1_7 ) );
  BUF_X2 U2591 ( .I(\MC_ARK_ARC_1_3/buf_output[7] ), .Z(\SB1_4_30/i0[6] ) );
  NAND3_X1 U2593 ( .A1(\SB3_21/i0[8] ), .A2(\SB3_21/i3[0] ), .A3(n3182), .ZN(
        n4856) );
  CLKBUF_X4 U2606 ( .I(\MC_ARK_ARC_1_3/buf_output[9] ), .Z(\SB1_4_30/i0[10] )
         );
  INV_X1 U2624 ( .I(\SB3_18/buf_output[2] ), .ZN(\SB4_15/i1[9] ) );
  NAND2_X1 U2634 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i3[0] ), .ZN(
        \SB4_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2635 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i0_3 ), .A3(\SB4_11/i0_4 ), 
        .ZN(\SB4_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2636 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i0_3 ), .A3(\SB4_11/i0[7] ), 
        .ZN(n1911) );
  NAND3_X1 U2638 ( .A1(\SB4_11/i0[9] ), .A2(\SB4_11/i0_0 ), .A3(\SB4_11/i0[8] ), .ZN(\SB4_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2639 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i1_5 ), .A3(\SB4_11/i0_4 ), 
        .ZN(n3023) );
  NAND3_X1 U2650 ( .A1(\SB1_4_19/i0[9] ), .A2(\SB1_4_19/i0_3 ), .A3(
        \SB1_4_19/i0[8] ), .ZN(n3551) );
  NAND2_X1 U2653 ( .A1(\SB1_4_19/i0_3 ), .A2(\SB1_4_19/i1[9] ), .ZN(
        \SB1_4_19/Component_Function_1/NAND4_in[0] ) );
  INV_X1 U2656 ( .I(\MC_ARK_ARC_1_4/buf_output[63] ), .ZN(\SB3_21/i0[8] ) );
  BUF_X2 U2658 ( .I(\MC_ARK_ARC_1_4/buf_output[63] ), .Z(\SB3_21/i0[10] ) );
  INV_X1 U2661 ( .I(\RI1[4][141] ), .ZN(\SB1_4_8/i0[8] ) );
  BUF_X2 U2662 ( .I(\RI1[4][141] ), .Z(\SB1_4_8/i0[10] ) );
  INV_X1 U2663 ( .I(\SB3_21/buf_output[5] ), .ZN(\SB4_21/i1_5 ) );
  INV_X1 U2681 ( .I(\SB3_17/buf_output[1] ), .ZN(\SB4_13/i1_7 ) );
  BUF_X2 U2683 ( .I(\SB3_17/buf_output[1] ), .Z(\SB4_13/i0[6] ) );
  NAND3_X1 U2684 ( .A1(\SB3_11/i0_0 ), .A2(\SB3_11/i0_4 ), .A3(\SB3_11/i1_5 ), 
        .ZN(n4967) );
  NAND2_X1 U2690 ( .A1(\SB3_11/i0_0 ), .A2(\SB3_11/i3[0] ), .ZN(
        \SB3_11/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U2705 ( .I(\MC_ARK_ARC_1_4/buf_output[92] ), .ZN(\SB3_16/i1[9] ) );
  BUF_X2 U2708 ( .I(\MC_ARK_ARC_1_4/buf_output[92] ), .Z(\SB3_16/i0_0 ) );
  NAND3_X1 U2711 ( .A1(\SB3_22/i0_0 ), .A2(\SB3_22/i0[6] ), .A3(
        \SB3_22/i0[10] ), .ZN(\SB3_22/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2715 ( .A1(\SB3_22/i1_5 ), .A2(\SB3_22/i0[10] ), .A3(
        \SB3_22/i1[9] ), .ZN(\SB3_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2716 ( .A1(\SB3_22/i1[9] ), .A2(\SB3_22/i1_7 ), .A3(
        \SB3_22/i0[10] ), .ZN(\SB3_22/Component_Function_3/NAND4_in[2] ) );
  BUF_X2 U2718 ( .I(\MC_ARK_ARC_1_4/buf_output[57] ), .Z(\SB3_22/i0[10] ) );
  NAND3_X1 U2721 ( .A1(\SB3_3/i0[9] ), .A2(\SB3_3/i0[6] ), .A3(\SB3_3/i0_4 ), 
        .ZN(\SB3_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2726 ( .A1(\SB2_0_2/i1[9] ), .A2(\SB2_0_2/i0_3 ), .A3(
        \SB2_0_2/i0[6] ), .ZN(\SB2_0_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2727 ( .A1(\SB2_0_2/i0_3 ), .A2(\SB2_0_2/i1[9] ), .A3(
        \RI3[0][178] ), .ZN(\SB2_0_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2730 ( .A1(\SB2_0_2/i1[9] ), .A2(\SB2_0_2/i1_5 ), .A3(
        \RI3[0][178] ), .ZN(\SB2_0_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2731 ( .A1(\SB2_0_2/i0[10] ), .A2(\SB2_0_2/i1_5 ), .A3(
        \SB2_0_2/i1[9] ), .ZN(\SB2_0_2/Component_Function_2/NAND4_in[0] ) );
  BUF_X2 U2736 ( .I(\SB3_3/buf_output[3] ), .Z(\SB4_1/i0[10] ) );
  CLKBUF_X4 U2737 ( .I(\SB2_4_6/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[165] ) );
  NAND3_X1 U2755 ( .A1(\SB1_3_23/i0_3 ), .A2(\MC_ARK_ARC_1_2/buf_output[52] ), 
        .A3(\SB1_3_23/i1[9] ), .ZN(\SB1_3_23/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U2763 ( .I(\MC_ARK_ARC_1_4/buf_output[99] ), .ZN(\SB3_15/i0[8] ) );
  BUF_X2 U2765 ( .I(\MC_ARK_ARC_1_4/buf_output[99] ), .Z(\SB3_15/i0[10] ) );
  NAND2_X1 U2780 ( .A1(\SB3_26/i0[10] ), .A2(\SB3_26/i0[9] ), .ZN(
        \SB3_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U2782 ( .A1(\SB4_14/i1[9] ), .A2(\SB4_14/i1_7 ), .A3(
        \SB4_14/i0[10] ), .ZN(\SB4_14/Component_Function_3/NAND4_in[2] ) );
  INV_X1 U2801 ( .I(\MC_ARK_ARC_1_4/buf_output[62] ), .ZN(\SB3_21/i1[9] ) );
  BUF_X2 U2802 ( .I(\MC_ARK_ARC_1_4/buf_output[62] ), .Z(\SB3_21/i0_0 ) );
  BUF_X2 U2805 ( .I(\MC_ARK_ARC_1_4/buf_output[120] ), .Z(\SB3_11/i0[9] ) );
  INV_X1 U2806 ( .I(\MC_ARK_ARC_1_4/buf_output[120] ), .ZN(\SB3_11/i3[0] ) );
  CLKBUF_X4 U2808 ( .I(\SB1_0_14/buf_output[5] ), .Z(\SB2_0_14/i0_3 ) );
  NAND3_X1 U2810 ( .A1(\SB1_4_18/i0[10] ), .A2(\SB1_4_18/i1[9] ), .A3(
        \SB1_4_18/i1_7 ), .ZN(n2577) );
  NAND2_X1 U2821 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i0[9] ), .ZN(
        \SB4_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U2823 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i0_3 ), .A3(
        \SB4_11/i0[6] ), .ZN(n5260) );
  INV_X1 U2828 ( .I(n4249), .ZN(n954) );
  NAND3_X1 U2829 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i0[8] ), .A3(
        \SB1_1_26/i0[9] ), .ZN(\SB1_1_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2830 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i0_3 ), .A3(
        \SB1_1_26/i0[6] ), .ZN(n4614) );
  NAND3_X1 U2834 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i0_4 ), .A3(
        \SB1_1_26/i0_3 ), .ZN(\SB1_1_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2835 ( .A1(\SB1_1_26/i0_0 ), .A2(\SB1_1_26/i0_3 ), .A3(
        \SB1_1_26/i0_4 ), .ZN(\SB1_1_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2842 ( .A1(\SB1_4_28/i0_0 ), .A2(\SB1_4_28/i1_5 ), .A3(
        \SB1_4_28/i0_4 ), .ZN(n2172) );
  NAND3_X1 U2858 ( .A1(n3976), .A2(\SB3_29/i1[9] ), .A3(\SB3_29/i0_4 ), .ZN(
        \SB3_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2861 ( .A1(\SB3_29/i1_5 ), .A2(\SB3_29/i1[9] ), .A3(\SB3_29/i0_4 ), 
        .ZN(n3027) );
  NAND3_X1 U2868 ( .A1(\SB4_20/i0_0 ), .A2(\SB4_20/i0[9] ), .A3(\SB4_20/i0[8] ), .ZN(n2698) );
  NAND2_X1 U2869 ( .A1(\SB4_20/i0_0 ), .A2(\SB4_20/i3[0] ), .ZN(
        \SB4_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2875 ( .A1(\SB4_20/i0_0 ), .A2(\SB4_20/i3[0] ), .A3(\SB4_20/i1_7 ), 
        .ZN(n3607) );
  INV_X1 U2876 ( .I(n351), .ZN(\SB1_0_14/i0[8] ) );
  BUF_X2 U2877 ( .I(n351), .Z(\SB1_0_14/i0[10] ) );
  CLKBUF_X4 U2878 ( .I(\SB3_13/buf_output[3] ), .Z(\SB4_11/i0[10] ) );
  NAND2_X1 U2879 ( .A1(\MC_ARK_ARC_1_2/buf_output[128] ), .A2(\SB1_3_10/i3[0] ), .ZN(\SB1_3_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2881 ( .A1(\SB1_3_10/i0_0 ), .A2(\SB1_3_10/i0_3 ), .A3(
        \SB1_3_10/i0_4 ), .ZN(\SB1_3_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2882 ( .A1(\SB1_3_10/i0_0 ), .A2(\SB1_3_10/i0_3 ), .A3(
        \SB1_3_10/i0[7] ), .ZN(n4942) );
  NAND3_X1 U2883 ( .A1(\SB1_3_10/i0_0 ), .A2(\SB1_3_10/i0[6] ), .A3(
        \SB1_3_10/i0[10] ), .ZN(\SB1_3_10/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U2899 ( .A1(n6273), .A2(\SB4_19/i0_0 ), .A3(\SB4_19/i0_4 ), .ZN(
        \SB4_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2901 ( .A1(\SB3_15/buf_output[3] ), .A2(\SB4_13/i1[9] ), .A3(
        \SB4_13/i1_7 ), .ZN(\SB4_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2902 ( .A1(n4002), .A2(\SB3_15/buf_output[3] ), .A3(\SB4_13/i1[9] ), .ZN(\SB4_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2909 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0[10] ), .A3(
        \SB2_3_31/i0[6] ), .ZN(\SB2_3_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2917 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0_0 ), .A3(
        \SB2_3_31/i0[7] ), .ZN(n1163) );
  NAND3_X1 U2922 ( .A1(\SB2_0_28/i1[9] ), .A2(\SB2_0_28/i1_5 ), .A3(
        \SB2_0_28/i0_4 ), .ZN(\SB2_0_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2923 ( .A1(\SB2_0_28/i1_5 ), .A2(\SB2_0_28/i0[10] ), .A3(
        \SB2_0_28/i1[9] ), .ZN(\SB2_0_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2924 ( .A1(\SB2_0_28/i1[9] ), .A2(\SB2_0_28/i0_3 ), .A3(
        \SB2_0_28/i0[6] ), .ZN(\SB2_0_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2948 ( .A1(\SB1_3_17/i0[9] ), .A2(\SB1_3_17/i0[6] ), .A3(
        \SB1_3_17/i1_5 ), .ZN(n3622) );
  NAND3_X1 U2953 ( .A1(\SB2_4_25/i0[10] ), .A2(\SB2_4_25/i1_7 ), .A3(
        \SB2_4_25/i1[9] ), .ZN(\SB2_4_25/Component_Function_3/NAND4_in[2] ) );
  BUF_X2 U2956 ( .I(\SB3_23/buf_output[2] ), .Z(\SB4_20/i0_0 ) );
  AND2_X1 U2957 ( .A1(\MC_ARK_ARC_1_2/buf_output[88] ), .A2(
        \MC_ARK_ARC_1_2/buf_output[85] ), .Z(n588) );
  CLKBUF_X4 U2958 ( .I(n398), .Z(\SB1_0_14/i0_3 ) );
  INV_X1 U2959 ( .I(n398), .ZN(\SB1_0_14/i1_5 ) );
  NAND3_X1 U2965 ( .A1(\SB1_0_23/i0_0 ), .A2(\SB1_0_23/i1_5 ), .A3(
        \SB1_0_23/i0_4 ), .ZN(\SB1_0_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2970 ( .A1(\SB4_23/i1_5 ), .A2(\SB4_23/i0[10] ), .A3(
        \SB4_23/i1[9] ), .ZN(\SB4_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2971 ( .A1(\SB4_23/i0[10] ), .A2(\SB4_23/i1[9] ), .A3(
        \SB4_23/i1_7 ), .ZN(n3350) );
  INV_X1 U2978 ( .I(\SB3_28/buf_output[2] ), .ZN(\SB4_25/i1[9] ) );
  NAND3_X1 U2979 ( .A1(n3998), .A2(\SB4_21/i1_7 ), .A3(\SB4_21/i0[10] ), .ZN(
        \SB4_21/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2997 ( .A1(\SB1_4_15/i0_0 ), .A2(\SB1_4_15/i0_3 ), .A3(
        \MC_ARK_ARC_1_3/buf_output[100] ), .ZN(
        \SB1_4_15/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U3009 ( .I(\SB1_2_30/buf_output[1] ), .ZN(\SB2_2_26/i1_7 ) );
  BUF_X2 U3011 ( .I(\SB1_2_30/buf_output[1] ), .Z(\SB2_2_26/i0[6] ) );
  NAND3_X1 U3012 ( .A1(\SB1_3_24/i1[9] ), .A2(\SB1_3_24/i1_5 ), .A3(
        \SB1_3_24/i0_4 ), .ZN(\SB1_3_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3014 ( .A1(\SB1_3_24/i0[10] ), .A2(\SB1_3_24/i1[9] ), .A3(
        \SB1_3_24/i1_7 ), .ZN(\SB1_3_24/Component_Function_3/NAND4_in[2] ) );
  BUF_X2 U3023 ( .I(\MC_ARK_ARC_1_3/buf_output[109] ), .Z(\SB1_4_13/i0[6] ) );
  NAND3_X1 U3028 ( .A1(\SB2_4_9/i1[9] ), .A2(\SB2_4_9/i0_3 ), .A3(
        \SB2_4_9/i0[6] ), .ZN(\SB2_4_9/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U3040 ( .A1(\SB4_25/i0[10] ), .A2(n6266), .ZN(
        \SB4_25/Component_Function_0/NAND4_in[0] ) );
  INV_X1 U3043 ( .I(\SB1_1_13/buf_output[1] ), .ZN(\SB2_1_9/i1_7 ) );
  NAND3_X1 U3048 ( .A1(\SB1_1_11/i0_3 ), .A2(\SB1_1_11/i1_7 ), .A3(
        \SB1_1_11/i0[8] ), .ZN(\SB1_1_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U3050 ( .A1(\SB1_1_11/i0_3 ), .A2(\SB1_1_11/i1[9] ), .ZN(
        \SB1_1_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3051 ( .A1(\SB1_1_11/i0_3 ), .A2(\MC_ARK_ARC_1_0/buf_output[120] ), 
        .A3(\SB1_1_11/i0[8] ), .ZN(n4016) );
  NAND3_X1 U3052 ( .A1(\SB1_1_11/i0[10] ), .A2(\SB1_1_11/i0_3 ), .A3(
        \SB1_1_11/i0_4 ), .ZN(n3292) );
  NAND2_X1 U3059 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i0[9] ), .ZN(
        \SB4_29/Component_Function_0/NAND4_in[0] ) );
  INV_X8 U3072 ( .I(\RI1[4][119] ), .ZN(\SB1_4_12/i1_5 ) );
  NAND3_X1 U3079 ( .A1(\SB1_0_17/i0[10] ), .A2(\SB1_0_17/i1[9] ), .A3(
        \SB1_0_17/i1_5 ), .ZN(n1485) );
  NAND3_X1 U3080 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i0_4 ), .A3(
        \SB1_0_17/i1[9] ), .ZN(\SB1_0_17/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U3085 ( .I(\MC_ARK_ARC_1_4/buf_output[176] ), .Z(\SB3_2/i0_0 ) );
  NAND3_X1 U3091 ( .A1(\SB2_1_19/i0_3 ), .A2(\SB2_1_19/i1_7 ), .A3(
        \SB2_1_19/i0[8] ), .ZN(\SB2_1_19/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3093 ( .A1(\SB4_21/i0_3 ), .A2(\SB4_21/i1_7 ), .A3(\SB4_21/i0[8] ), 
        .ZN(\SB4_21/Component_Function_1/NAND4_in[1] ) );
  INV_X1 U3096 ( .I(\MC_ARK_ARC_1_2/buf_output[127] ), .ZN(\SB1_3_10/i1_7 ) );
  NAND3_X1 U3113 ( .A1(\SB1_2_14/i0_0 ), .A2(\SB1_2_14/i0[6] ), .A3(
        \SB1_2_14/i0[10] ), .ZN(\SB1_2_14/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U3120 ( .A1(\SB1_0_5/i0_0 ), .A2(\SB1_0_5/i0_4 ), .A3(
        \SB1_0_5/i1_5 ), .ZN(n3938) );
  NAND3_X1 U3121 ( .A1(\SB1_0_16/i0_0 ), .A2(\SB1_0_16/i0_3 ), .A3(
        \SB1_0_16/i0_4 ), .ZN(\SB1_0_16/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U3145 ( .I(\MC_ARK_ARC_1_2/buf_output[25] ), .ZN(\SB1_3_27/i1_7 ) );
  NAND3_X1 U3154 ( .A1(\SB1_3_20/i0[10] ), .A2(\SB1_3_20/i1[9] ), .A3(
        \SB1_3_20/i1_7 ), .ZN(\SB1_3_20/Component_Function_3/NAND4_in[2] ) );
  INV_X1 U3156 ( .I(\MC_ARK_ARC_1_1/buf_output[168] ), .ZN(\SB1_2_3/i3[0] ) );
  INV_X1 U3157 ( .I(\MC_ARK_ARC_1_0/buf_output[84] ), .ZN(\SB1_1_17/i3[0] ) );
  BUF_X4 U3158 ( .I(\MC_ARK_ARC_1_0/buf_output[84] ), .Z(\SB1_1_17/i0[9] ) );
  CLKBUF_X4 U3182 ( .I(\MC_ARK_ARC_1_3/buf_output[32] ), .Z(\SB1_4_26/i0_0 )
         );
  INV_X1 U3187 ( .I(n402), .ZN(\SB1_0_10/i1_5 ) );
  INV_X1 U3196 ( .I(\MC_ARK_ARC_1_0/buf_output[138] ), .ZN(\SB1_1_8/i3[0] ) );
  CLKBUF_X4 U3209 ( .I(\SB3_23/buf_output[3] ), .Z(\SB4_21/i0[10] ) );
  NAND3_X1 U3210 ( .A1(\SB3_15/i0_0 ), .A2(\SB3_15/i0_3 ), .A3(\SB3_15/i0_4 ), 
        .ZN(\SB3_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3211 ( .A1(\SB3_15/i0[6] ), .A2(\SB3_15/i0_3 ), .A3(\SB3_15/i1[9] ), .ZN(\SB3_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3212 ( .A1(\SB3_15/i0[6] ), .A2(\SB3_15/i0_3 ), .A3(
        \SB3_15/i0[10] ), .ZN(\SB3_15/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 U3219 ( .A1(\SB1_3_22/i0_3 ), .A2(\SB1_3_22/i1[9] ), .ZN(
        \SB1_3_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3221 ( .A1(\SB1_3_22/i0[9] ), .A2(\SB1_3_22/i0[10] ), .A3(
        \SB1_3_22/i0_3 ), .ZN(\SB1_3_22/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3226 ( .A1(\SB1_2_5/i0_0 ), .A2(\SB1_2_5/i0_3 ), .A3(
        \SB1_2_5/i0_4 ), .ZN(\SB1_2_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3230 ( .A1(\SB1_2_5/i0[10] ), .A2(\SB1_2_5/i0_4 ), .A3(
        \SB1_2_5/i0_3 ), .ZN(\SB1_2_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3237 ( .A1(\SB1_2_5/i0[10] ), .A2(\SB1_2_5/i0_3 ), .A3(
        \SB1_2_5/i0[9] ), .ZN(n929) );
  NAND3_X1 U3240 ( .A1(\SB1_1_27/i0[7] ), .A2(\SB1_1_27/i0_3 ), .A3(
        \SB1_1_27/i0_0 ), .ZN(\SB1_1_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3242 ( .A1(\SB1_1_27/i0[9] ), .A2(\SB1_1_27/i0[10] ), .A3(
        \SB1_1_27/i0_3 ), .ZN(\SB1_1_27/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U3247 ( .I(n355), .ZN(\SB1_0_12/i0[8] ) );
  NAND3_X1 U3248 ( .A1(\SB1_4_30/i1_5 ), .A2(\SB1_4_30/i0[10] ), .A3(
        \SB1_4_30/i1[9] ), .ZN(\SB1_4_30/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U3251 ( .I(\SB1_3_1/buf_output[1] ), .ZN(\SB2_3_29/i1_7 ) );
  CLKBUF_X4 U3264 ( .I(\SB2_3_20/buf_output[3] ), .Z(\RI5[3][81] ) );
  NAND4_X2 U3265 ( .A1(\SB2_4_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_4_30/Component_Function_1/NAND4_in[2] ), .A3(n5172), .A4(
        \SB2_4_30/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_4_30/buf_output[1] ) );
  OR3_X2 U3269 ( .A1(\RI3[2][95] ), .A2(\SB1_2_18/buf_output[3] ), .A3(
        \SB1_2_21/buf_output[0] ), .Z(
        \SB2_2_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3272 ( .A1(\SB1_3_30/i0[10] ), .A2(\SB1_3_30/i1[9] ), .A3(
        \SB1_3_30/i1_7 ), .ZN(n5109) );
  CLKBUF_X4 U3275 ( .I(\MC_ARK_ARC_1_0/buf_output[98] ), .Z(\SB1_1_15/i0_0 )
         );
  NAND3_X1 U3284 ( .A1(\SB1_4_16/i0_0 ), .A2(\SB1_4_16/i0[9] ), .A3(
        \SB1_4_16/i0[8] ), .ZN(\SB1_4_16/Component_Function_4/NAND4_in[0] ) );
  CLKBUF_X4 U3285 ( .I(\MC_ARK_ARC_1_2/buf_output[164] ), .Z(\SB1_3_4/i0_0 )
         );
  INV_X1 U3292 ( .I(\MC_ARK_ARC_1_0/buf_output[30] ), .ZN(\SB1_1_26/i3[0] ) );
  INV_X1 U3294 ( .I(\MC_ARK_ARC_1_2/buf_output[120] ), .ZN(\SB1_3_11/i3[0] )
         );
  BUF_X2 U3295 ( .I(\MC_ARK_ARC_1_2/buf_output[120] ), .Z(\SB1_3_11/i0[9] ) );
  NAND3_X1 U3298 ( .A1(\SB2_0_27/i0_3 ), .A2(\SB2_0_27/i0[9] ), .A3(
        \SB2_0_27/i0[8] ), .ZN(\SB2_0_27/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U3300 ( .I(\MC_ARK_ARC_1_4/buf_output[111] ), .Z(\SB3_13/i0[10] ) );
  INV_X1 U3303 ( .I(\SB1_2_11/buf_output[5] ), .ZN(\SB2_2_11/i1_5 ) );
  NAND3_X1 U3326 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0[10] ), .A3(
        \SB2_2_24/i0_4 ), .ZN(\SB2_2_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3327 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0_0 ), .A3(
        \SB2_2_24/i0_4 ), .ZN(\SB2_2_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3333 ( .A1(\SB1_1_27/i0[8] ), .A2(\SB1_1_27/i0[7] ), .A3(
        \SB1_1_27/i0[6] ), .ZN(\SB1_1_27/Component_Function_0/NAND4_in[1] ) );
  CLKBUF_X4 U3337 ( .I(\MC_ARK_ARC_1_4/buf_output[177] ), .Z(\SB3_2/i0[10] )
         );
  INV_X1 U3341 ( .I(\MC_ARK_ARC_1_2/buf_output[85] ), .ZN(\SB1_3_17/i1_7 ) );
  INV_X1 U3342 ( .I(\MC_ARK_ARC_1_2/buf_output[11] ), .ZN(\SB1_3_30/i1_5 ) );
  CLKBUF_X4 U3343 ( .I(\MC_ARK_ARC_1_1/buf_output[132] ), .Z(\SB1_2_9/i0[9] )
         );
  BUF_X2 U3344 ( .I(\SB1_3_17/buf_output[1] ), .Z(\SB2_3_13/i0[6] ) );
  INV_X1 U3347 ( .I(\SB1_3_17/buf_output[1] ), .ZN(\SB2_3_13/i1_7 ) );
  INV_X1 U3351 ( .I(\MC_ARK_ARC_1_3/buf_output[18] ), .ZN(\SB1_4_28/i3[0] ) );
  BUF_X2 U3352 ( .I(\SB3_9/buf_output[1] ), .Z(\SB4_5/i0[6] ) );
  BUF_X2 U3356 ( .I(\SB3_14/buf_output[1] ), .Z(\SB4_10/i0[6] ) );
  CLKBUF_X4 U3358 ( .I(\SB3_14/buf_output[2] ), .Z(\SB4_11/i0_0 ) );
  BUF_X2 U3364 ( .I(\SB3_31/buf_output[1] ), .Z(\SB4_27/i0[6] ) );
  BUF_X2 U3366 ( .I(\SB3_5/buf_output[1] ), .Z(\SB4_1/i0[6] ) );
  BUF_X2 U3367 ( .I(\SB3_2/buf_output[1] ), .Z(\SB4_30/i0[6] ) );
  BUF_X2 U3382 ( .I(\MC_ARK_ARC_1_4/buf_output[138] ), .Z(\SB3_8/i0[9] ) );
  CLKBUF_X4 U3383 ( .I(\MC_ARK_ARC_1_4/buf_output[76] ), .Z(\SB3_19/i0_4 ) );
  CLKBUF_X4 U3385 ( .I(\MC_ARK_ARC_1_4/buf_output[170] ), .Z(\SB3_3/i0_0 ) );
  BUF_X4 U3386 ( .I(\SB2_4_30/buf_output[0] ), .Z(\RI5[4][36] ) );
  BUF_X4 U3389 ( .I(\SB2_4_3/buf_output[1] ), .Z(\RI5[4][1] ) );
  BUF_X4 U3407 ( .I(\SB1_4_14/buf_output[5] ), .Z(\SB2_4_14/i0_3 ) );
  BUF_X2 U3414 ( .I(\MC_ARK_ARC_1_3/buf_output[144] ), .Z(\SB1_4_7/i0[9] ) );
  NAND3_X2 U3418 ( .A1(\SB1_4_0/i0[8] ), .A2(\SB1_4_0/i1_7 ), .A3(
        \SB1_4_0/i0_4 ), .ZN(\SB1_4_0/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 U3435 ( .I(\SB2_3_18/buf_output[4] ), .Z(\RI5[3][88] ) );
  BUF_X4 U3436 ( .I(n2287), .Z(\SB2_3_8/i0_3 ) );
  CLKBUF_X4 U3441 ( .I(\SB1_3_20/buf_output[3] ), .Z(\SB2_3_18/i0[10] ) );
  BUF_X4 U3448 ( .I(n3986), .Z(\SB1_3_21/i0_3 ) );
  BUF_X4 U3453 ( .I(\SB2_2_25/buf_output[4] ), .Z(\RI5[2][46] ) );
  BUF_X4 U3454 ( .I(\SB2_2_28/buf_output[3] ), .Z(\RI5[2][33] ) );
  BUF_X4 U3461 ( .I(\SB2_2_11/buf_output[4] ), .Z(\RI5[2][130] ) );
  CLKBUF_X4 U3462 ( .I(\SB2_2_5/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[181] ) );
  NAND2_X1 U3466 ( .A1(\SB2_2_31/i0[8] ), .A2(n4961), .ZN(n4960) );
  NAND3_X2 U3467 ( .A1(\SB2_2_6/i0[10] ), .A2(\SB2_2_6/i1_7 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(n2983) );
  CLKBUF_X4 U3468 ( .I(\SB1_2_14/buf_output[2] ), .Z(\SB2_2_11/i0_0 ) );
  BUF_X2 U3469 ( .I(\SB1_2_31/buf_output[0] ), .Z(\SB2_2_26/i0[9] ) );
  CLKBUF_X4 U3486 ( .I(\MC_ARK_ARC_1_1/buf_output[134] ), .Z(\SB1_2_9/i0_0 )
         );
  BUF_X4 U3495 ( .I(\SB2_1_17/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[94] ) );
  BUF_X4 U3499 ( .I(\SB2_0_24/buf_output[2] ), .Z(\RI5[0][62] ) );
  BUF_X4 U3502 ( .I(\SB2_0_4/buf_output[3] ), .Z(\RI5[0][177] ) );
  CLKBUF_X4 U3510 ( .I(\SB2_0_5/buf_output[5] ), .Z(\RI5[0][161] ) );
  CLKBUF_X4 U3511 ( .I(\SB1_0_29/buf_output[2] ), .Z(\SB2_0_26/i0_0 ) );
  NAND2_X1 U3514 ( .A1(\SB1_0_18/Component_Function_4/NAND4_in[1] ), .A2(n3870), .ZN(n2326) );
  NAND2_X1 U3519 ( .A1(\SB1_0_5/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_5/Component_Function_4/NAND4_in[0] ), .ZN(n3568) );
  BUF_X2 U3529 ( .I(n309), .Z(\SB1_0_3/i0[9] ) );
  NAND2_X1 U3531 ( .A1(\SB1_0_20/i1[9] ), .A2(n4187), .ZN(
        \SB1_0_20/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3532 ( .A1(\SB1_0_29/i0[9] ), .A2(\SB1_0_29/i0[10] ), .A3(
        \SB1_0_29/i0_3 ), .ZN(\SB1_0_29/Component_Function_4/NAND4_in[2] ) );
  CLKBUF_X4 U3534 ( .I(n310), .Z(\SB1_0_3/i0_0 ) );
  INV_X1 U3535 ( .I(n326), .ZN(\SB1_0_27/i0[7] ) );
  NAND3_X1 U3537 ( .A1(\SB1_0_10/i0_0 ), .A2(\SB1_0_10/i1_5 ), .A3(
        \SB1_0_10/i0_4 ), .ZN(n1913) );
  NAND3_X1 U3540 ( .A1(\SB1_0_26/i1[9] ), .A2(\SB1_0_26/i1_7 ), .A3(
        \SB1_0_26/i0[10] ), .ZN(\SB1_0_26/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U3541 ( .A1(\SB1_0_14/i0_0 ), .A2(\SB1_0_14/i0[6] ), .A3(
        \SB1_0_14/i0[10] ), .ZN(\SB1_0_14/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U3542 ( .A1(\SB1_0_10/i0[8] ), .A2(\SB1_0_10/i0[7] ), .A3(
        \SB1_0_10/i0[6] ), .ZN(\SB1_0_10/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3543 ( .A1(\SB1_0_5/i0_3 ), .A2(\SB1_0_5/i0_0 ), .A3(
        \SB1_0_5/i0_4 ), .ZN(\SB1_0_5/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U3544 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i1[9] ), .ZN(
        \SB1_0_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3545 ( .A1(\SB1_0_9/i0[10] ), .A2(\SB1_0_9/i1[9] ), .A3(
        \SB1_0_9/i1_7 ), .ZN(n1589) );
  NAND3_X1 U3546 ( .A1(\SB1_0_7/i0_0 ), .A2(\SB1_0_7/i0[10] ), .A3(
        \SB1_0_7/i0[6] ), .ZN(\SB1_0_7/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3550 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i0[10] ), .A3(
        \SB1_0_7/i0[6] ), .ZN(\SB1_0_7/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 U3552 ( .A1(\SB1_0_21/i0[10] ), .A2(\SB1_0_21/i0[9] ), .ZN(
        \SB1_0_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3553 ( .A1(\SB1_0_21/i1_5 ), .A2(\SB1_0_21/i0[6] ), .A3(
        \SB1_0_21/i0[9] ), .ZN(\SB1_0_21/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U3554 ( .A1(\SB1_0_4/i0[10] ), .A2(\SB1_0_4/i0[9] ), .ZN(
        \SB1_0_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3555 ( .A1(\SB1_0_14/i1_5 ), .A2(\SB1_0_14/i1[9] ), .A3(
        \SB1_0_14/i0_4 ), .ZN(\SB1_0_14/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U3556 ( .I(\SB1_0_22/buf_output[3] ), .Z(\SB2_0_20/i0[10] ) );
  NAND3_X1 U3570 ( .A1(\SB2_0_9/i0[10] ), .A2(\SB2_0_9/i1_5 ), .A3(
        \SB2_0_9/i1[9] ), .ZN(\SB2_0_9/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 U3571 ( .I(\SB1_0_6/buf_output[3] ), .Z(\SB2_0_4/i0[10] ) );
  NAND2_X1 U3581 ( .A1(\SB2_0_3/i0_3 ), .A2(\SB2_0_3/i1[9] ), .ZN(
        \SB2_0_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3583 ( .A1(\SB2_0_0/i0[10] ), .A2(\SB2_0_0/i0_3 ), .A3(
        \RI3[0][190] ), .ZN(n5220) );
  NAND3_X1 U3584 ( .A1(\SB2_0_30/i0[10] ), .A2(\SB2_0_30/i1_7 ), .A3(
        \SB2_0_30/i1[9] ), .ZN(\SB2_0_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3587 ( .A1(n2886), .A2(\SB2_0_9/i0_3 ), .A3(\SB2_0_9/i0[7] ), .ZN(
        n2628) );
  NAND3_X1 U3590 ( .A1(\SB2_0_13/i1_5 ), .A2(\SB2_0_13/i0[10] ), .A3(
        \SB2_0_13/i1[9] ), .ZN(\SB2_0_13/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U3595 ( .I(\SB1_0_21/buf_output[1] ), .ZN(\SB2_0_17/i1_7 ) );
  NAND3_X1 U3597 ( .A1(\SB2_0_0/i0_0 ), .A2(\SB2_0_0/i0_3 ), .A3(\RI3[0][190] ), .ZN(\SB2_0_0/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X1 U3606 ( .I(n68), .Z(\MC_ARK_ARC_1_0/buf_keyinput[92] ) );
  CLKBUF_X4 U3608 ( .I(\SB2_0_3/buf_output[2] ), .Z(\RI5[0][188] ) );
  NAND3_X1 U3627 ( .A1(\SB1_1_10/i1[9] ), .A2(\SB1_1_10/i1_7 ), .A3(
        \SB1_1_10/i0[10] ), .ZN(\SB1_1_10/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U3628 ( .A1(\SB1_1_5/i1_5 ), .A2(\SB1_1_5/i0_0 ), .A3(
        \SB1_1_5/i0_4 ), .ZN(\SB1_1_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3629 ( .A1(\SB1_1_26/i0[9] ), .A2(\SB1_1_26/i0[10] ), .A3(
        \SB1_1_26/i0_3 ), .ZN(\SB1_1_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3631 ( .A1(\SB1_1_12/i0[9] ), .A2(\SB1_1_12/i0[10] ), .A3(
        \SB1_1_12/i0_3 ), .ZN(\SB1_1_12/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U3639 ( .A1(\SB1_1_27/i0_3 ), .A2(\SB1_1_27/i1[9] ), .ZN(
        \SB1_1_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3641 ( .A1(\SB1_1_1/i1[9] ), .A2(\SB1_1_1/i1_5 ), .A3(
        \SB1_1_1/i0_4 ), .ZN(\SB1_1_1/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U3643 ( .A1(\SB1_1_8/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_1_8/Component_Function_1/NAND4_in[0] ), .ZN(n2755) );
  NAND3_X1 U3663 ( .A1(\SB1_1_2/i0[9] ), .A2(\SB1_1_2/i1_5 ), .A3(
        \SB1_1_2/i0[6] ), .ZN(n2856) );
  NAND3_X1 U3682 ( .A1(\SB2_1_17/i0[6] ), .A2(n3990), .A3(\SB2_1_17/i0[9] ), 
        .ZN(\SB2_1_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3691 ( .A1(\SB2_1_5/i1[9] ), .A2(\SB2_1_5/i1_5 ), .A3(
        \SB2_1_5/i0_4 ), .ZN(\SB2_1_5/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U3704 ( .I(\MC_ARK_ARC_1_1/buf_output[103] ), .ZN(\SB1_2_14/i1_7 ) );
  CLKBUF_X4 U3705 ( .I(\MC_ARK_ARC_1_1/buf_output[178] ), .Z(\SB1_2_2/i0_4 )
         );
  CLKBUF_X4 U3710 ( .I(\MC_ARK_ARC_1_1/buf_output[145] ), .Z(\SB1_2_7/i0[6] )
         );
  CLKBUF_X4 U3716 ( .I(\MC_ARK_ARC_1_1/buf_output[56] ), .Z(\SB1_2_22/i0_0 )
         );
  NAND3_X1 U3717 ( .A1(\SB1_2_17/i0[7] ), .A2(\SB1_2_17/i0_3 ), .A3(
        \SB1_2_17/i0_0 ), .ZN(\SB1_2_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3721 ( .A1(\SB1_2_20/i0[8] ), .A2(\SB1_2_20/i0[7] ), .A3(
        \SB1_2_20/i0[6] ), .ZN(\SB1_2_20/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3726 ( .A1(\SB1_2_3/i3[0] ), .A2(\SB1_2_3/i0_0 ), .A3(
        \SB1_2_3/i1_7 ), .ZN(\SB1_2_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3729 ( .A1(\SB1_2_4/i0[10] ), .A2(\SB1_2_4/i0_4 ), .A3(
        \SB1_2_4/i0_3 ), .ZN(\SB1_2_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3730 ( .A1(\SB1_2_3/i0[9] ), .A2(\SB1_2_3/i1_5 ), .A3(
        \SB1_2_3/i0[6] ), .ZN(\SB1_2_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3732 ( .A1(\SB1_2_28/i1[9] ), .A2(\SB1_2_28/i1_5 ), .A3(
        \SB1_2_28/i0_4 ), .ZN(n4584) );
  NAND3_X1 U3733 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i0_3 ), .A3(
        \SB1_2_18/i0_4 ), .ZN(\SB1_2_18/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U3749 ( .I(\SB1_2_5/buf_output[0] ), .ZN(\SB2_2_0/i3[0] ) );
  CLKBUF_X4 U3750 ( .I(\SB1_2_17/buf_output[3] ), .Z(\SB2_2_15/i0[10] ) );
  CLKBUF_X4 U3754 ( .I(\SB1_2_7/buf_output[2] ), .Z(\SB2_2_4/i0_0 ) );
  CLKBUF_X4 U3758 ( .I(\SB1_2_21/buf_output[3] ), .Z(\SB2_2_19/i0[10] ) );
  NAND3_X1 U3763 ( .A1(\SB2_2_27/i0_4 ), .A2(\SB2_2_27/i0[8] ), .A3(
        \SB2_2_27/i1_7 ), .ZN(n5031) );
  NAND3_X1 U3767 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i0[9] ), .A3(
        \SB2_2_17/i0[10] ), .ZN(n1387) );
  NAND3_X1 U3769 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0[8] ), .A3(
        \SB2_2_29/i1_7 ), .ZN(\SB2_2_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U3771 ( .A1(\SB2_2_26/i0[10] ), .A2(\SB2_2_26/i0[9] ), .ZN(
        \SB2_2_26/Component_Function_0/NAND4_in[0] ) );
  CLKBUF_X4 U3773 ( .I(\SB2_2_21/buf_output[0] ), .Z(\RI5[2][90] ) );
  INV_X1 U3774 ( .I(\MC_ARK_ARC_1_2/buf_output[137] ), .ZN(\SB1_3_9/i1_5 ) );
  CLKBUF_X4 U3787 ( .I(\MC_ARK_ARC_1_2/buf_output[117] ), .Z(\SB1_3_12/i0[10] ) );
  INV_X1 U3798 ( .I(\MC_ARK_ARC_1_2/buf_output[162] ), .ZN(\SB1_3_4/i3[0] ) );
  NAND3_X1 U3813 ( .A1(\SB1_3_15/i0[8] ), .A2(\SB1_3_15/i1_5 ), .A3(
        \SB1_3_15/i3[0] ), .ZN(n2516) );
  NAND3_X1 U3839 ( .A1(\SB1_3_17/i1_7 ), .A2(\SB1_3_17/i0_3 ), .A3(
        \SB1_3_17/i0[8] ), .ZN(n4323) );
  CLKBUF_X4 U3850 ( .I(\SB1_3_25/buf_output[0] ), .Z(\SB2_3_20/i0[9] ) );
  CLKBUF_X4 U3857 ( .I(\SB1_3_2/buf_output[3] ), .Z(\SB2_3_0/i0[10] ) );
  CLKBUF_X4 U3859 ( .I(\SB1_3_27/buf_output[0] ), .Z(\SB2_3_22/i0[9] ) );
  NAND3_X1 U3867 ( .A1(\SB1_3_1/buf_output[4] ), .A2(\SB2_3_0/i0[8] ), .A3(
        \SB2_3_0/i1_7 ), .ZN(\SB2_3_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3871 ( .A1(\SB2_3_10/i3[0] ), .A2(\SB2_3_10/i0[8] ), .A3(
        \SB2_3_10/i1_5 ), .ZN(\SB2_3_10/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 U3874 ( .A1(\SB2_3_8/i0[10] ), .A2(\SB2_3_8/i0[9] ), .ZN(
        \SB2_3_8/Component_Function_0/NAND4_in[0] ) );
  CLKBUF_X4 U3878 ( .I(\SB1_3_29/buf_output[2] ), .Z(\SB2_3_26/i0_0 ) );
  INV_X1 U3895 ( .I(\MC_ARK_ARC_1_3/buf_output[66] ), .ZN(\SB1_4_20/i3[0] ) );
  NAND3_X1 U3916 ( .A1(\SB1_4_4/i1_7 ), .A2(\SB1_4_4/i0[8] ), .A3(
        \SB1_4_4/i0_4 ), .ZN(\SB1_4_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3944 ( .A1(\SB1_4_11/i3[0] ), .A2(\SB1_4_11/i0[8] ), .A3(
        \SB1_4_11/i1_5 ), .ZN(n1734) );
  NAND2_X1 U3949 ( .A1(\SB1_4_2/i0_3 ), .A2(\SB1_4_2/i1[9] ), .ZN(
        \SB1_4_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3952 ( .A1(\RI1[4][119] ), .A2(\SB1_4_12/i1[9] ), .A3(
        \SB1_4_12/i0[6] ), .ZN(\SB1_4_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3964 ( .A1(\SB1_4_31/i1_5 ), .A2(\SB1_4_31/i0[8] ), .A3(
        \SB1_4_31/i3[0] ), .ZN(\SB1_4_31/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X4 U3966 ( .I(\SB1_4_18/buf_output[0] ), .Z(\SB2_4_13/i0[9] ) );
  NAND3_X1 U3973 ( .A1(\SB2_4_7/i1_5 ), .A2(\SB2_4_7/i0[6] ), .A3(
        \SB2_4_7/i0[9] ), .ZN(\SB2_4_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3978 ( .A1(\SB2_4_10/i1_7 ), .A2(\SB2_4_10/i0[8] ), .A3(
        \SB2_4_10/i0_4 ), .ZN(\SB2_4_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3989 ( .A1(\SB2_4_11/i1[9] ), .A2(\SB2_4_11/i1_5 ), .A3(
        \SB2_4_11/i0_4 ), .ZN(\SB2_4_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3993 ( .A1(\SB2_4_25/i0[8] ), .A2(\SB2_4_25/i0[7] ), .A3(
        \SB2_4_25/i0[6] ), .ZN(\SB2_4_25/Component_Function_0/NAND4_in[1] ) );
  INV_X1 U3996 ( .I(n22), .ZN(n494) );
  NAND3_X1 U3999 ( .A1(\SB2_4_9/i0[10] ), .A2(\SB2_4_9/i1_7 ), .A3(
        \SB2_4_9/i1[9] ), .ZN(n4292) );
  CLKBUF_X4 U4025 ( .I(\MC_ARK_ARC_1_4/buf_output[25] ), .Z(\SB3_27/i0[6] ) );
  INV_X1 U4028 ( .I(\MC_ARK_ARC_1_4/buf_output[43] ), .ZN(\SB3_24/i1_7 ) );
  INV_X1 U4034 ( .I(\MC_ARK_ARC_1_4/buf_output[174] ), .ZN(\SB3_2/i3[0] ) );
  NAND3_X1 U4039 ( .A1(\SB3_15/i0[9] ), .A2(\SB3_15/i0[6] ), .A3(\SB3_15/i1_5 ), .ZN(\SB3_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4040 ( .A1(\SB3_29/i1[9] ), .A2(\SB3_29/i1_7 ), .A3(
        \SB3_29/i0[10] ), .ZN(\SB3_29/Component_Function_3/NAND4_in[2] ) );
  NAND2_X1 U4042 ( .A1(\SB3_5/i0_0 ), .A2(\SB3_5/i3[0] ), .ZN(
        \SB3_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4045 ( .A1(\SB3_24/i0[10] ), .A2(\SB3_24/i1[9] ), .A3(
        \SB3_24/i1_7 ), .ZN(n4586) );
  CLKBUF_X4 U4052 ( .I(\MC_ARK_ARC_1_4/buf_output[40] ), .Z(\SB3_25/i0_4 ) );
  NAND3_X1 U4054 ( .A1(\SB3_23/i0_0 ), .A2(\SB3_23/i0[6] ), .A3(
        \SB3_23/i0[10] ), .ZN(\SB3_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4055 ( .A1(\SB3_5/i0_0 ), .A2(\SB3_5/i1_5 ), .A3(\SB3_5/i0_4 ), 
        .ZN(n2283) );
  NAND3_X1 U4058 ( .A1(\SB3_22/i1[9] ), .A2(\SB3_22/i0_3 ), .A3(\SB3_22/i0[6] ), .ZN(\SB3_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4062 ( .A1(\SB3_10/i1_5 ), .A2(\SB3_10/i0[8] ), .A3(\SB3_10/i3[0] ), .ZN(\SB3_10/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 U4065 ( .A1(\SB3_20/i0_3 ), .A2(\SB3_20/i1[9] ), .ZN(
        \SB3_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U4069 ( .A1(\SB3_5/i1[9] ), .A2(\SB3_5/i1_5 ), .A3(\SB3_5/i0_4 ), 
        .ZN(\SB3_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4070 ( .A1(\SB3_22/i1_5 ), .A2(\SB3_22/i0[6] ), .A3(\SB3_22/i0[9] ), .ZN(\SB3_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4073 ( .A1(\SB3_5/i0_0 ), .A2(\SB3_5/i0_3 ), .A3(\SB3_5/i0[7] ), 
        .ZN(n3632) );
  INV_X1 U4080 ( .I(\SB3_26/buf_output[0] ), .ZN(\SB4_21/i3[0] ) );
  CLKBUF_X4 U4083 ( .I(\SB3_19/buf_output[4] ), .Z(\SB4_18/i0_4 ) );
  NAND3_X1 U4099 ( .A1(\SB4_13/i0_4 ), .A2(\SB4_13/i1[9] ), .A3(n4002), .ZN(
        \SB4_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4100 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i0[6] ), .A3(\SB4_28/i1[9] ), .ZN(n5237) );
  NAND3_X1 U4107 ( .A1(\SB4_5/i3[0] ), .A2(\SB4_5/i0_0 ), .A3(\SB4_5/i1_7 ), 
        .ZN(\SB4_5/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 U4109 ( .A1(\SB3_24/buf_output[2] ), .A2(\SB4_21/i3[0] ), .ZN(
        \SB4_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4113 ( .A1(\SB4_25/i1_5 ), .A2(\SB4_25/i0[6] ), .A3(n6266), .ZN(
        \SB4_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4126 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i1[9] ), .A3(\SB4_13/i0_4 ), 
        .ZN(\SB4_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4129 ( .A1(\SB4_19/i0[10] ), .A2(\SB4_19/i0[9] ), .A3(
        \SB4_19/i0_3 ), .ZN(n2092) );
  NAND3_X1 U4130 ( .A1(\SB4_5/i0[7] ), .A2(\SB4_5/i0_3 ), .A3(\SB4_5/i0_0 ), 
        .ZN(\SB4_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4135 ( .A1(\SB4_13/i0_4 ), .A2(n1498), .A3(\SB4_13/i1_7 ), .ZN(
        n2183) );
  NAND3_X1 U4140 ( .A1(\SB4_26/i0[10] ), .A2(\SB4_26/i0[6] ), .A3(
        \SB3_29/buf_output[2] ), .ZN(n960) );
  NAND2_X1 U4141 ( .A1(\SB4_22/i0[10] ), .A2(\SB4_22/i0[9] ), .ZN(
        \SB4_22/Component_Function_0/NAND4_in[0] ) );
  CLKBUF_X1 U4143 ( .I(Key[35]), .Z(n123) );
  AND2_X1 U4144 ( .A1(\SB1_2_24/Component_Function_4/NAND4_in[2] ), .A2(n919), 
        .Z(n3169) );
  NOR2_X1 U4151 ( .A1(n5959), .A2(\RI3[0][60] ), .ZN(n3171) );
  CLKBUF_X4 U4156 ( .I(\SB1_2_12/buf_output[2] ), .Z(\SB2_2_9/i0_0 ) );
  AND2_X1 U4158 ( .A1(\SB1_0_12/Component_Function_2/NAND4_in[2] ), .A2(n835), 
        .Z(n3173) );
  XNOR2_X1 U4160 ( .A1(\SB2_1_26/buf_output[2] ), .A2(n88), .ZN(n3175) );
  AND2_X1 U4165 ( .A1(\SB1_4_20/buf_output[0] ), .A2(\SB2_4_15/i0[8] ), .Z(
        n3177) );
  XNOR2_X1 U4167 ( .A1(\SB2_3_18/buf_output[5] ), .A2(n543), .ZN(n3179) );
  AND3_X1 U4169 ( .A1(\SB2_1_4/i1[9] ), .A2(\SB2_1_4/i1_5 ), .A3(
        \SB2_1_4/i0_4 ), .Z(n3180) );
  XNOR2_X1 U4173 ( .A1(n4227), .A2(n4226), .ZN(n3182) );
  OR2_X2 U4174 ( .A1(n2718), .A2(n4792), .Z(n3183) );
  XNOR2_X1 U4178 ( .A1(n3009), .A2(n5105), .ZN(n3184) );
  XOR2_X1 U4180 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[71] ), .A2(n546), .Z(n3185) );
  XOR2_X1 U4181 ( .A1(\RI5[1][101] ), .A2(\RI5[1][137] ), .Z(n3186) );
  NAND3_X2 U4184 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i0_3 ), .A3(
        \SB4_16/i0[6] ), .ZN(n3188) );
  INV_X1 U4192 ( .I(\SB1_2_25/buf_output[1] ), .ZN(\SB2_2_21/i1_7 ) );
  NAND4_X2 U4193 ( .A1(\SB1_2_25/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_25/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_2_25/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_2_25/buf_output[1] ) );
  NAND4_X2 U4194 ( .A1(\SB1_2_8/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_8/Component_Function_2/NAND4_in[3] ), .A3(n4926), .A4(n3190), 
        .ZN(\SB1_2_8/buf_output[2] ) );
  NAND3_X2 U4196 ( .A1(\SB1_2_8/i0[10] ), .A2(\SB1_2_8/i0_3 ), .A3(
        \SB1_2_8/i0[6] ), .ZN(n3190) );
  NAND4_X2 U4197 ( .A1(\SB1_1_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_25/Component_Function_0/NAND4_in[0] ), .A4(n3191), .ZN(
        \SB1_1_25/buf_output[0] ) );
  NAND3_X1 U4201 ( .A1(\SB4_24/i0_4 ), .A2(\SB4_24/i0_0 ), .A3(\SB4_24/i0_3 ), 
        .ZN(\SB4_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U4206 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i1[9] ), .A3(
        \SB1_0_22/i0[6] ), .ZN(\SB1_0_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4219 ( .A1(\SB4_5/i0[9] ), .A2(\SB4_5/i0_3 ), .A3(\SB4_5/i0[8] ), 
        .ZN(\SB4_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U4222 ( .A1(\SB2_0_20/i1_5 ), .A2(\SB2_0_20/i3[0] ), .A3(
        \SB2_0_20/i0[8] ), .ZN(\SB2_0_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U4227 ( .A1(\SB2_3_19/i0_0 ), .A2(\SB2_3_19/i0[10] ), .A3(
        \SB2_3_19/i0[6] ), .ZN(n3193) );
  NAND3_X1 U4228 ( .A1(\SB4_3/i0[10] ), .A2(\SB4_3/i1[9] ), .A3(\SB4_3/i1_7 ), 
        .ZN(n4949) );
  NAND4_X2 U4232 ( .A1(\SB2_2_17/Component_Function_3/NAND4_in[0] ), .A2(n3508), .A3(\SB2_2_17/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_2_17/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_2_17/buf_output[3] ) );
  XOR2_X1 U4233 ( .A1(n5410), .A2(n3194), .Z(\MC_ARK_ARC_1_4/temp5[40] ) );
  XOR2_X1 U4237 ( .A1(\RI5[4][10] ), .A2(\RI5[4][178] ), .Z(n3194) );
  NAND4_X2 U4241 ( .A1(\SB1_3_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_21/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_3_21/Component_Function_3/NAND4_in[2] ), .A4(n1412), .ZN(
        \SB1_3_21/buf_output[3] ) );
  XOR2_X1 U4247 ( .A1(\RI5[4][149] ), .A2(\RI5[4][143] ), .Z(n4032) );
  NAND3_X1 U4252 ( .A1(\SB1_3_10/i3[0] ), .A2(\SB1_3_10/i1_5 ), .A3(
        \SB1_3_10/i0[8] ), .ZN(n1304) );
  NAND3_X1 U4254 ( .A1(\SB4_24/i0_4 ), .A2(\SB4_24/i1_7 ), .A3(n1494), .ZN(
        \SB4_24/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U4255 ( .A1(\SB2_2_4/Component_Function_5/NAND4_in[2] ), .A2(n5379), 
        .A3(\SB2_2_4/Component_Function_5/NAND4_in[1] ), .A4(n1520), .ZN(
        \SB2_2_4/buf_output[5] ) );
  NAND3_X1 U4258 ( .A1(\SB2_1_2/i0_3 ), .A2(\SB2_1_2/i0_0 ), .A3(
        \SB2_1_2/i0_4 ), .ZN(\SB2_1_2/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U4259 ( .A1(\SB2_2_8/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_8/Component_Function_4/NAND4_in[0] ), .A3(n3359), .A4(n3196), 
        .ZN(\SB2_2_8/buf_output[4] ) );
  NAND3_X1 U4260 ( .A1(\SB2_2_8/i0_0 ), .A2(\SB2_2_8/i3[0] ), .A3(
        \SB2_2_8/i1_7 ), .ZN(n3196) );
  NAND4_X2 U4272 ( .A1(n1523), .A2(\SB1_3_2/Component_Function_5/NAND4_in[1] ), 
        .A3(n3961), .A4(\SB1_3_2/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_2/buf_output[5] ) );
  NAND4_X2 U4277 ( .A1(\SB2_1_8/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_1_8/Component_Function_5/NAND4_in[1] ), .A3(n859), .A4(
        \SB2_1_8/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_1_8/buf_output[5] ) );
  XOR2_X1 U4281 ( .A1(\MC_ARK_ARC_1_1/temp6[185] ), .A2(n3198), .Z(
        \RI1[2][185] ) );
  XOR2_X1 U4289 ( .A1(\RI5[0][122] ), .A2(\RI5[0][146] ), .Z(
        \MC_ARK_ARC_1_0/temp2[176] ) );
  XOR2_X1 U4290 ( .A1(n3200), .A2(n3199), .Z(n4787) );
  XOR2_X1 U4292 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[146] ), .A2(n74), .Z(n3199) );
  XOR2_X1 U4293 ( .A1(\RI5[1][80] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .Z(n3200) );
  NAND3_X1 U4295 ( .A1(\SB2_4_18/i0_0 ), .A2(\SB1_4_19/buf_output[4] ), .A3(
        \SB2_4_18/i1_5 ), .ZN(n3201) );
  XOR2_X1 U4297 ( .A1(\RI5[1][166] ), .A2(\RI5[1][118] ), .Z(n3202) );
  XOR2_X1 U4300 ( .A1(n578), .A2(\RI5[1][142] ), .Z(n3203) );
  XOR2_X1 U4301 ( .A1(n3205), .A2(n3204), .Z(n4750) );
  XOR2_X1 U4307 ( .A1(\RI5[3][149] ), .A2(n514), .Z(n3204) );
  NAND4_X2 U4312 ( .A1(n3725), .A2(\SB2_3_1/Component_Function_0/NAND4_in[2] ), 
        .A3(\SB2_3_1/Component_Function_0/NAND4_in[1] ), .A4(n3206), .ZN(
        \SB2_3_1/buf_output[0] ) );
  NAND2_X1 U4313 ( .A1(\SB2_3_1/i0[9] ), .A2(\SB2_3_1/i0[10] ), .ZN(n3206) );
  NAND4_X2 U4322 ( .A1(\SB1_4_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_4_2/Component_Function_3/NAND4_in[2] ), .A4(n3207), .ZN(
        \SB1_4_2/buf_output[3] ) );
  NAND3_X2 U4323 ( .A1(\SB2_1_20/i0_3 ), .A2(\SB2_1_20/i0_4 ), .A3(
        \SB2_1_20/i1[9] ), .ZN(n1490) );
  NAND4_X2 U4325 ( .A1(\SB1_1_16/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_16/Component_Function_3/NAND4_in[2] ), .A3(n4337), .A4(n3208), 
        .ZN(\SB1_1_16/buf_output[3] ) );
  INV_X1 U4326 ( .I(\SB1_2_3/buf_output[1] ), .ZN(\SB2_2_31/i1_7 ) );
  NAND4_X2 U4331 ( .A1(\SB1_2_3/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_3/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_2_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_3/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_3/buf_output[1] ) );
  NAND2_X2 U4336 ( .A1(n2387), .A2(n2001), .ZN(\RI5[4][175] ) );
  XOR2_X1 U4355 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[173] ), .A2(\RI5[4][143] ), 
        .Z(n1789) );
  NAND4_X2 U4359 ( .A1(\SB1_2_29/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_1/NAND4_in[0] ), .A4(n3212), .ZN(
        \SB1_2_29/buf_output[1] ) );
  NAND3_X2 U4362 ( .A1(\SB2_2_21/i0[10] ), .A2(\SB2_2_21/i1_7 ), .A3(
        \SB2_2_21/i1[9] ), .ZN(n1654) );
  NAND3_X1 U4365 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i3[0] ), .A3(\SB4_22/i1_7 ), 
        .ZN(n3213) );
  INV_X2 U4367 ( .I(\SB1_1_7/buf_output[2] ), .ZN(\SB2_1_4/i1[9] ) );
  XOR2_X1 U4373 ( .A1(\MC_ARK_ARC_1_4/temp1[25] ), .A2(n3214), .Z(
        \MC_ARK_ARC_1_4/temp5[25] ) );
  XOR2_X1 U4374 ( .A1(\RI5[4][187] ), .A2(\RI5[4][163] ), .Z(n3214) );
  XOR2_X1 U4375 ( .A1(n3215), .A2(n19), .Z(Ciphertext[56]) );
  XOR2_X1 U4378 ( .A1(\RI5[3][134] ), .A2(\RI5[3][110] ), .Z(n1608) );
  NAND4_X2 U4380 ( .A1(n2783), .A2(n2116), .A3(n1025), .A4(n3216), .ZN(
        \SB2_4_25/buf_output[5] ) );
  XOR2_X1 U4387 ( .A1(n3218), .A2(\MC_ARK_ARC_1_4/temp4[51] ), .Z(
        \MC_ARK_ARC_1_4/temp6[51] ) );
  XOR2_X1 U4389 ( .A1(\RI5[4][153] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[117] ), 
        .Z(n3218) );
  NAND3_X1 U4390 ( .A1(\SB4_18/i1_7 ), .A2(\SB4_18/i3[0] ), .A3(\SB4_18/i0_0 ), 
        .ZN(\SB4_18/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U4411 ( .A1(\MC_ARK_ARC_1_4/temp5[55] ), .A2(n3221), .Z(
        \MC_ARK_ARC_1_4/buf_output[55] ) );
  XOR2_X1 U4412 ( .A1(\MC_ARK_ARC_1_4/temp3[55] ), .A2(
        \MC_ARK_ARC_1_4/temp4[55] ), .Z(n3221) );
  NAND4_X2 U4413 ( .A1(\SB1_2_25/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_25/Component_Function_2/NAND4_in[0] ), .A3(n3758), .A4(n606), 
        .ZN(\SB1_2_25/buf_output[2] ) );
  INV_X8 U4422 ( .I(n3222), .ZN(\RI1[3][107] ) );
  INV_X2 U4424 ( .I(\MC_ARK_ARC_1_2/buf_output[107] ), .ZN(n3222) );
  XOR2_X1 U4425 ( .A1(\RI5[0][92] ), .A2(\RI5[0][98] ), .Z(
        \MC_ARK_ARC_1_0/temp1[98] ) );
  XOR2_X1 U4430 ( .A1(\RI5[1][126] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[162] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[60] ) );
  NAND4_X2 U4437 ( .A1(\SB2_4_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_0/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_4_0/Component_Function_2/NAND4_in[1] ), .A4(n3223), .ZN(
        \SB2_4_0/buf_output[2] ) );
  NAND3_X2 U4438 ( .A1(\SB2_4_0/i0_4 ), .A2(n3978), .A3(\SB2_4_0/i0_0 ), .ZN(
        n3223) );
  XOR2_X1 U4446 ( .A1(n3225), .A2(\MC_ARK_ARC_1_2/temp1[120] ), .Z(
        \MC_ARK_ARC_1_2/temp5[120] ) );
  XOR2_X1 U4447 ( .A1(\RI5[2][90] ), .A2(\RI5[2][66] ), .Z(n3225) );
  XOR2_X1 U4454 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[87] ), .A2(\RI5[4][123] ), 
        .Z(n3226) );
  NAND3_X1 U4457 ( .A1(\SB2_3_28/i0_0 ), .A2(\SB2_3_28/i3[0] ), .A3(
        \SB2_3_28/i1_7 ), .ZN(n3227) );
  XOR2_X1 U4458 ( .A1(\RI5[3][60] ), .A2(\RI5[3][54] ), .Z(
        \MC_ARK_ARC_1_3/temp1[60] ) );
  NAND4_X2 U4462 ( .A1(\SB1_4_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_21/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_4_21/Component_Function_3/NAND4_in[1] ), .A4(n3229), .ZN(
        \SB1_4_21/buf_output[3] ) );
  NAND3_X1 U4463 ( .A1(\SB1_4_21/i0[8] ), .A2(\SB1_4_21/i3[0] ), .A3(
        \SB1_4_21/i1_5 ), .ZN(n3229) );
  XOR2_X1 U4469 ( .A1(n3231), .A2(\MC_ARK_ARC_1_2/temp1[144] ), .Z(
        \MC_ARK_ARC_1_2/temp5[144] ) );
  XOR2_X1 U4470 ( .A1(\RI5[2][90] ), .A2(\RI5[2][114] ), .Z(n3231) );
  NAND4_X2 U4486 ( .A1(\SB2_2_31/Component_Function_0/NAND4_in[1] ), .A2(n1770), .A3(n1481), .A4(n3234), .ZN(\SB2_2_31/buf_output[0] ) );
  XOR2_X1 U4534 ( .A1(\RI5[2][85] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[121] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[19] ) );
  NAND4_X2 U4562 ( .A1(\SB2_3_12/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_3_12/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_12/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_3_12/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_3_12/buf_output[3] ) );
  NAND3_X2 U4570 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0_4 ), .A3(
        \SB2_1_10/i1[9] ), .ZN(n3287) );
  NAND4_X2 U4573 ( .A1(\SB2_0_19/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_19/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_0_19/Component_Function_1/NAND4_in[0] ), .A4(n3248), .ZN(
        \SB2_0_19/buf_output[1] ) );
  NAND3_X2 U4574 ( .A1(\SB2_0_19/i0[8] ), .A2(\RI3[0][76] ), .A3(
        \SB2_0_19/i1_7 ), .ZN(n3248) );
  XOR2_X1 U4575 ( .A1(n3249), .A2(\MC_ARK_ARC_1_0/temp4[57] ), .Z(n3103) );
  XOR2_X1 U4576 ( .A1(\SB2_0_13/buf_output[3] ), .A2(\SB2_0_7/buf_output[3] ), 
        .Z(n3249) );
  XOR2_X1 U4584 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[182] ), .A2(\RI5[1][158] ), 
        .Z(n3252) );
  XOR2_X1 U4586 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[110] ), .A2(\RI5[1][104] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[110] ) );
  XOR2_X1 U4588 ( .A1(\RI5[4][179] ), .A2(\RI5[4][185] ), .Z(n4447) );
  NAND4_X2 U4590 ( .A1(\SB2_0_21/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_21/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_21/Component_Function_3/NAND4_in[3] ), .A4(n3253), .ZN(
        \SB2_0_21/buf_output[3] ) );
  NAND4_X2 U4592 ( .A1(\SB1_4_28/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_4_28/Component_Function_3/NAND4_in[0] ), .A3(n3255), .A4(n3254), 
        .ZN(\SB1_4_28/buf_output[3] ) );
  NAND3_X2 U4594 ( .A1(\SB1_2_23/i0_0 ), .A2(\SB1_2_23/i0[10] ), .A3(
        \SB1_2_23/i0[6] ), .ZN(n3256) );
  NAND3_X1 U4603 ( .A1(\SB2_0_19/i0[6] ), .A2(\RI3[0][77] ), .A3(
        \SB2_0_19/i1[9] ), .ZN(\SB2_0_19/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U4616 ( .A1(n3141), .A2(n3257), .Z(\MC_ARK_ARC_1_3/buf_output[74] )
         );
  XOR2_X1 U4617 ( .A1(n4972), .A2(\MC_ARK_ARC_1_3/temp4[74] ), .Z(n3257) );
  XOR2_X1 U4632 ( .A1(n3263), .A2(n3262), .Z(\MC_ARK_ARC_1_2/buf_output[107] )
         );
  XOR2_X1 U4633 ( .A1(n3310), .A2(\MC_ARK_ARC_1_2/temp4[107] ), .Z(n3262) );
  XOR2_X1 U4634 ( .A1(\MC_ARK_ARC_1_2/temp2[107] ), .A2(
        \MC_ARK_ARC_1_2/temp3[107] ), .Z(n3263) );
  XOR2_X1 U4641 ( .A1(n3266), .A2(n3265), .Z(\MC_ARK_ARC_1_2/temp5[35] ) );
  XOR2_X1 U4646 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[35] ), .A2(\RI5[2][173] ), 
        .Z(n3266) );
  NAND3_X2 U4647 ( .A1(\SB2_1_25/i0[6] ), .A2(\SB2_1_25/i0_0 ), .A3(
        \SB1_1_27/buf_output[3] ), .ZN(n3436) );
  OR3_X1 U4652 ( .A1(\RI1[4][155] ), .A2(n3967), .A3(
        \MC_ARK_ARC_1_3/buf_output[150] ), .Z(n3957) );
  XOR2_X1 U4659 ( .A1(\MC_ARK_ARC_1_0/temp1[129] ), .A2(n3270), .Z(
        \MC_ARK_ARC_1_0/temp5[129] ) );
  XOR2_X1 U4660 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[75] ), .A2(\RI5[0][99] ), 
        .Z(n3270) );
  XOR2_X1 U4662 ( .A1(n3272), .A2(n3271), .Z(\MC_ARK_ARC_1_1/buf_output[95] )
         );
  XOR2_X1 U4664 ( .A1(n3588), .A2(\MC_ARK_ARC_1_1/temp4[95] ), .Z(n3272) );
  XOR2_X1 U4673 ( .A1(\MC_ARK_ARC_1_1/temp3[4] ), .A2(
        \MC_ARK_ARC_1_1/temp4[4] ), .Z(\MC_ARK_ARC_1_1/temp6[4] ) );
  NAND4_X2 U4677 ( .A1(\SB2_0_16/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_16/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_0_16/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_0_16/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_16/buf_output[0] ) );
  NAND3_X1 U4679 ( .A1(\SB1_0_15/i0_3 ), .A2(n285), .A3(\SB1_0_15/i0[8] ), 
        .ZN(\SB1_0_15/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U4687 ( .A1(\SB2_1_8/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_8/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_8/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_1_8/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB2_1_8/buf_output[2] ) );
  NAND3_X1 U4688 ( .A1(\SB1_2_14/i0[10] ), .A2(\SB1_2_14/i1_5 ), .A3(
        \SB1_2_14/i1[9] ), .ZN(\SB1_2_14/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U4689 ( .A1(\SB2_1_9/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_9/Component_Function_1/NAND4_in[2] ), .A3(n2378), .A4(
        \SB2_1_9/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_9/buf_output[1] ) );
  INV_X2 U4692 ( .I(\SB1_1_17/buf_output[2] ), .ZN(\SB2_1_14/i1[9] ) );
  NAND3_X1 U4694 ( .A1(\SB1_0_29/i0[10] ), .A2(\SB1_0_29/i1_5 ), .A3(
        \SB1_0_29/i1[9] ), .ZN(\SB1_0_29/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U4699 ( .A1(\SB2_2_18/Component_Function_0/NAND4_in[3] ), .A2(n2708), .A3(\SB2_2_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_18/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_18/buf_output[0] ) );
  NAND3_X2 U4713 ( .A1(\SB2_0_16/i0_3 ), .A2(n6976), .A3(\SB2_0_16/i0[9] ), 
        .ZN(n2600) );
  XOR2_X1 U4727 ( .A1(n3279), .A2(\MC_ARK_ARC_1_2/temp1[0] ), .Z(n877) );
  XOR2_X1 U4728 ( .A1(\RI5[2][138] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .Z(n3279) );
  XOR2_X1 U4729 ( .A1(n3280), .A2(n4385), .Z(n5385) );
  XOR2_X1 U4731 ( .A1(\RI5[1][131] ), .A2(\RI5[1][137] ), .Z(n3280) );
  XOR2_X1 U4735 ( .A1(n1546), .A2(\MC_ARK_ARC_1_2/temp6[146] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[146] ) );
  INV_X2 U4753 ( .I(\SB1_2_4/buf_output[3] ), .ZN(\SB2_2_2/i0[8] ) );
  XOR2_X1 U4756 ( .A1(\MC_ARK_ARC_1_2/temp4[146] ), .A2(
        \MC_ARK_ARC_1_2/temp3[146] ), .Z(\MC_ARK_ARC_1_2/temp6[146] ) );
  INV_X2 U4764 ( .I(\SB1_0_16/buf_output[3] ), .ZN(\SB2_0_14/i0[8] ) );
  NOR2_X2 U4775 ( .A1(n5388), .A2(n3286), .ZN(n3061) );
  NAND2_X2 U4780 ( .A1(\SB2_3_4/i0_0 ), .A2(\SB2_3_4/i3[0] ), .ZN(n3288) );
  XOR2_X1 U4782 ( .A1(n3150), .A2(n3289), .Z(\MC_ARK_ARC_1_1/temp5[131] ) );
  XOR2_X1 U4784 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[125] ), .A2(\RI5[1][131] ), 
        .Z(n3289) );
  XOR2_X1 U4785 ( .A1(n3290), .A2(\MC_ARK_ARC_1_1/temp4[171] ), .Z(n1348) );
  XOR2_X1 U4787 ( .A1(\RI5[1][81] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[45] ), 
        .Z(n3290) );
  NAND4_X2 U4791 ( .A1(\SB1_1_11/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_1_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_11/Component_Function_0/NAND4_in[0] ), .A4(n3292), .ZN(
        \SB1_1_11/buf_output[0] ) );
  NAND4_X2 U4792 ( .A1(\SB1_0_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_19/Component_Function_4/NAND4_in[1] ), .A3(n1054), .A4(n3293), 
        .ZN(\SB1_0_19/buf_output[4] ) );
  XOR2_X1 U4795 ( .A1(\MC_ARK_ARC_1_0/temp3[17] ), .A2(
        \MC_ARK_ARC_1_0/temp1[17] ), .Z(n3295) );
  XOR2_X1 U4801 ( .A1(\MC_ARK_ARC_1_1/temp2[143] ), .A2(n3298), .Z(
        \MC_ARK_ARC_1_1/temp5[143] ) );
  XOR2_X1 U4802 ( .A1(\RI5[1][143] ), .A2(\RI5[1][137] ), .Z(n3298) );
  BUF_X4 U4803 ( .I(\SB1_4_26/buf_output[5] ), .Z(\SB2_4_26/i0_3 ) );
  XOR2_X1 U4810 ( .A1(n3299), .A2(n2265), .Z(\MC_ARK_ARC_1_1/buf_output[49] )
         );
  XOR2_X1 U4811 ( .A1(\MC_ARK_ARC_1_1/temp1[49] ), .A2(
        \MC_ARK_ARC_1_1/temp2[49] ), .Z(n3299) );
  XOR2_X1 U4813 ( .A1(\RI5[3][95] ), .A2(\RI5[3][131] ), .Z(
        \MC_ARK_ARC_1_3/temp3[29] ) );
  XOR2_X1 U4816 ( .A1(\RI5[1][77] ), .A2(\RI5[1][29] ), .Z(n4561) );
  XOR2_X1 U4832 ( .A1(\MC_ARK_ARC_1_0/temp1[110] ), .A2(
        \MC_ARK_ARC_1_0/temp4[110] ), .Z(n3302) );
  NOR2_X1 U4840 ( .A1(n4734), .A2(\SB1_2_4/buf_output[0] ), .ZN(n4961) );
  NAND4_X2 U4844 ( .A1(\SB1_2_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_9/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_2_9/Component_Function_4/NAND4_in[1] ), .A4(n3305), .ZN(
        \SB1_2_9/buf_output[4] ) );
  XOR2_X1 U4847 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[24] ), .A2(\RI5[3][48] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[78] ) );
  XOR2_X1 U4848 ( .A1(\RI5[1][59] ), .A2(\RI5[1][53] ), .Z(n3424) );
  XOR2_X1 U4850 ( .A1(\RI5[2][129] ), .A2(\RI5[2][165] ), .Z(
        \MC_ARK_ARC_1_2/temp3[63] ) );
  XOR2_X1 U4851 ( .A1(\RI5[1][47] ), .A2(\RI5[1][11] ), .Z(
        \MC_ARK_ARC_1_1/temp3[137] ) );
  NAND3_X2 U4854 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0_0 ), .A3(
        \SB2_2_25/i0_4 ), .ZN(n4976) );
  NOR2_X2 U4860 ( .A1(n4524), .A2(n3311), .ZN(n3308) );
  NAND3_X2 U4861 ( .A1(\SB2_1_26/i3[0] ), .A2(\SB2_1_26/i1_5 ), .A3(
        \SB2_1_26/i0[8] ), .ZN(\SB2_1_26/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U4864 ( .A1(\RI5[2][101] ), .A2(\RI5[2][107] ), .Z(n3310) );
  NAND4_X2 U4867 ( .A1(n2912), .A2(\SB4_29/Component_Function_4/NAND4_in[0] ), 
        .A3(n3724), .A4(n3312), .ZN(n3750) );
  XOR2_X1 U4875 ( .A1(\MC_ARK_ARC_1_0/temp5[85] ), .A2(
        \MC_ARK_ARC_1_0/temp6[85] ), .Z(\MC_ARK_ARC_1_0/buf_output[85] ) );
  NAND4_X2 U4887 ( .A1(\SB2_4_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_3/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_4_3/Component_Function_2/NAND4_in[3] ), .A4(n3316), .ZN(
        \SB2_4_3/buf_output[2] ) );
  NAND3_X2 U4892 ( .A1(\SB2_4_3/i0[10] ), .A2(\SB2_4_3/i0_3 ), .A3(
        \SB2_4_3/i0[6] ), .ZN(n3316) );
  NAND3_X2 U4901 ( .A1(\SB2_2_14/i0[6] ), .A2(\SB2_2_14/i0_4 ), .A3(
        \SB2_2_14/i0[9] ), .ZN(n3317) );
  NAND4_X2 U4902 ( .A1(\SB4_15/Component_Function_1/NAND4_in[2] ), .A2(n2069), 
        .A3(\SB4_15/Component_Function_1/NAND4_in[1] ), .A4(n3318), .ZN(n3404)
         );
  NAND2_X1 U4903 ( .A1(\SB4_15/i0_3 ), .A2(\SB4_15/i1[9] ), .ZN(n3318) );
  NAND4_X2 U4905 ( .A1(\SB1_3_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_21/Component_Function_2/NAND4_in[2] ), .A4(n3448), .ZN(
        \SB1_3_21/buf_output[2] ) );
  NAND4_X2 U4919 ( .A1(\SB1_0_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_21/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_21/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_0_21/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][65] ) );
  XOR2_X1 U4927 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[156] ), .A2(\RI5[3][180] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[18] ) );
  XOR2_X1 U4931 ( .A1(\SB2_3_22/buf_output[0] ), .A2(\RI5[3][120] ), .Z(
        \MC_ARK_ARC_1_3/temp3[18] ) );
  BUF_X4 U4948 ( .I(\RI1[1][23] ), .Z(\SB1_1_28/i0_3 ) );
  XOR2_X1 U4949 ( .A1(\MC_ARK_ARC_1_3/temp4[3] ), .A2(
        \MC_ARK_ARC_1_3/temp3[3] ), .Z(\MC_ARK_ARC_1_3/temp6[3] ) );
  XOR2_X1 U4952 ( .A1(n3326), .A2(n3325), .Z(\MC_ARK_ARC_1_1/buf_output[56] )
         );
  XOR2_X1 U4958 ( .A1(n3456), .A2(n1773), .Z(n3325) );
  INV_X2 U4970 ( .I(\RI1[1][23] ), .ZN(\SB1_1_28/i1_5 ) );
  NAND3_X2 U4976 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0[10] ), .A3(
        \SB2_1_9/i0[9] ), .ZN(\SB2_1_9/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U4979 ( .A1(\MC_ARK_ARC_1_1/temp1[14] ), .A2(n3327), .Z(n3708) );
  XOR2_X1 U4980 ( .A1(\RI5[1][116] ), .A2(\RI5[1][80] ), .Z(n3327) );
  NAND3_X2 U4997 ( .A1(\SB2_1_28/i0_4 ), .A2(\SB2_1_28/i1_5 ), .A3(
        \SB2_1_28/i0_0 ), .ZN(n3329) );
  XOR2_X1 U4998 ( .A1(\MC_ARK_ARC_1_1/temp5[2] ), .A2(n3330), .Z(
        \MC_ARK_ARC_1_1/buf_output[2] ) );
  XOR2_X1 U5002 ( .A1(\MC_ARK_ARC_1_1/temp3[2] ), .A2(
        \MC_ARK_ARC_1_1/temp4[2] ), .Z(n3330) );
  XOR2_X1 U5004 ( .A1(n3331), .A2(n1548), .Z(\MC_ARK_ARC_1_0/buf_output[68] )
         );
  XOR2_X1 U5006 ( .A1(\MC_ARK_ARC_1_0/temp3[68] ), .A2(n802), .Z(n3331) );
  NAND3_X2 U5036 ( .A1(\SB1_2_26/i0_3 ), .A2(\SB1_2_26/i0_4 ), .A3(
        \SB1_2_26/i1[9] ), .ZN(\SB1_2_26/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U5054 ( .A1(n3335), .A2(n3334), .Z(\MC_ARK_ARC_1_3/temp5[29] ) );
  XOR2_X1 U5059 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[29] ), .A2(\RI5[3][191] ), 
        .Z(n3334) );
  XOR2_X1 U5063 ( .A1(\RI5[3][167] ), .A2(\RI5[3][23] ), .Z(n3335) );
  XOR2_X1 U5071 ( .A1(\RI5[1][113] ), .A2(\RI5[1][137] ), .Z(n3337) );
  XOR2_X1 U5072 ( .A1(n3338), .A2(n216), .Z(Ciphertext[11]) );
  NAND4_X2 U5073 ( .A1(\SB4_30/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_30/Component_Function_5/NAND4_in[2] ), .A3(n2594), .A4(
        \SB4_30/Component_Function_5/NAND4_in[0] ), .ZN(n3338) );
  INV_X2 U5083 ( .I(\SB1_1_17/buf_output[3] ), .ZN(\SB2_1_15/i0[8] ) );
  XOR2_X1 U5091 ( .A1(\RI5[4][116] ), .A2(\RI5[4][152] ), .Z(
        \MC_ARK_ARC_1_4/temp3[50] ) );
  NAND3_X1 U5101 ( .A1(\SB2_4_11/i0_3 ), .A2(\SB2_4_11/i1[9] ), .A3(
        \SB2_4_11/i0[6] ), .ZN(\SB2_4_11/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U5115 ( .A1(n3344), .A2(n3343), .Z(\MC_ARK_ARC_1_1/buf_output[23] )
         );
  BUF_X4 U5130 ( .I(\MC_ARK_ARC_1_2/buf_output[20] ), .Z(\SB1_3_28/i0_0 ) );
  XOR2_X1 U5141 ( .A1(\MC_ARK_ARC_1_3/temp2[120] ), .A2(n3349), .Z(
        \MC_ARK_ARC_1_3/temp5[120] ) );
  XOR2_X1 U5148 ( .A1(\RI5[3][120] ), .A2(\RI5[3][114] ), .Z(n3349) );
  XOR2_X1 U5180 ( .A1(n3355), .A2(n3354), .Z(\MC_ARK_ARC_1_0/buf_output[109] )
         );
  XOR2_X1 U5183 ( .A1(\MC_ARK_ARC_1_0/temp2[109] ), .A2(
        \MC_ARK_ARC_1_0/temp4[109] ), .Z(n3355) );
  NAND3_X2 U5187 ( .A1(\SB2_0_6/i0_3 ), .A2(\SB2_0_6/i0[8] ), .A3(
        \SB2_0_6/i0[9] ), .ZN(\SB2_0_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U5192 ( .A1(\SB2_2_24/i0[10] ), .A2(\SB2_2_24/i1_5 ), .A3(
        \SB2_2_24/i1[9] ), .ZN(\SB2_2_24/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U5195 ( .A1(\RI5[0][153] ), .A2(\RI5[0][129] ), .Z(
        \MC_ARK_ARC_1_0/temp2[183] ) );
  NAND3_X1 U5211 ( .A1(\SB1_0_10/i0_3 ), .A2(\SB1_0_10/i0_4 ), .A3(
        \SB1_0_10/i1[9] ), .ZN(n3357) );
  NAND3_X2 U5218 ( .A1(\SB2_2_12/i0[10] ), .A2(\SB2_2_12/i1_5 ), .A3(
        \SB2_2_12/i1[9] ), .ZN(\SB2_2_12/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U5220 ( .A1(\SB1_0_13/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_13/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_0_13/Component_Function_4/NAND4_in[0] ), .A4(n3358), .ZN(
        \SB1_0_13/buf_output[4] ) );
  BUF_X4 U5229 ( .I(\SB2_1_2/buf_output[2] ), .Z(\RI5[1][2] ) );
  NAND3_X1 U5236 ( .A1(\SB2_2_8/i0[10] ), .A2(\SB2_2_8/i0[9] ), .A3(
        \SB2_2_8/i0_3 ), .ZN(n3359) );
  NAND3_X1 U5240 ( .A1(\SB1_2_6/i0_0 ), .A2(\SB1_2_6/i0_3 ), .A3(
        \SB1_2_6/i0[7] ), .ZN(n4214) );
  XOR2_X1 U5260 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[75] ), .A2(\RI5[0][39] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[165] ) );
  BUF_X4 U5262 ( .I(\SB2_4_10/buf_output[5] ), .Z(\RI5[4][131] ) );
  NAND4_X2 U5271 ( .A1(\SB1_1_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_26/Component_Function_3/NAND4_in[1] ), .A3(n2392), .A4(
        \SB1_1_26/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_26/buf_output[3] ) );
  XOR2_X1 U5273 ( .A1(\RI5[2][191] ), .A2(\RI5[2][185] ), .Z(
        \MC_ARK_ARC_1_2/temp1[191] ) );
  NAND3_X2 U5276 ( .A1(\SB2_1_24/i0[10] ), .A2(\SB2_1_24/i0[6] ), .A3(
        \SB2_1_24/i0_0 ), .ZN(\SB2_1_24/Component_Function_5/NAND4_in[1] ) );
  NOR2_X2 U5279 ( .A1(n3363), .A2(n3362), .ZN(n4003) );
  NAND4_X2 U5281 ( .A1(\SB2_2_1/Component_Function_3/NAND4_in[0] ), .A2(n4526), 
        .A3(n2721), .A4(n4669), .ZN(\SB2_2_1/buf_output[3] ) );
  INV_X1 U5285 ( .I(\SB1_0_22/buf_output[1] ), .ZN(\SB2_0_18/i1_7 ) );
  NAND4_X2 U5286 ( .A1(\SB1_0_22/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_22/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_0_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_22/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_22/buf_output[1] ) );
  XOR2_X1 U5287 ( .A1(n3364), .A2(n65), .Z(Ciphertext[131]) );
  XOR2_X1 U5308 ( .A1(\RI5[3][146] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[140] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[146] ) );
  XOR2_X1 U5313 ( .A1(n3367), .A2(n3070), .Z(\MC_ARK_ARC_1_4/temp5[3] ) );
  XOR2_X1 U5314 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[3] ), .A2(\RI5[4][189] ), 
        .Z(n3367) );
  NAND3_X1 U5331 ( .A1(\SB2_4_2/i0_3 ), .A2(\SB2_4_2/i0_0 ), .A3(
        \SB2_4_2/i0[7] ), .ZN(\SB2_4_2/Component_Function_0/NAND4_in[3] ) );
  BUF_X2 U5334 ( .I(\SB3_20/buf_output[2] ), .Z(\SB4_17/i0_0 ) );
  XOR2_X1 U5347 ( .A1(n3368), .A2(\MC_ARK_ARC_1_4/temp6[66] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[66] ) );
  NOR2_X2 U5353 ( .A1(n3621), .A2(n3512), .ZN(n3370) );
  NAND3_X2 U5383 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0[10] ), .A3(
        \SB2_3_10/i0[6] ), .ZN(n3373) );
  NAND3_X1 U5404 ( .A1(\SB4_31/i0_3 ), .A2(\SB4_31/i0[10] ), .A3(
        \SB4_31/i0[6] ), .ZN(n3375) );
  NAND3_X2 U5410 ( .A1(\SB2_4_2/i0_3 ), .A2(\SB2_4_2/i0_0 ), .A3(
        \SB2_4_2/i0_4 ), .ZN(\SB2_4_2/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U5420 ( .A1(n2404), .A2(n4223), .A3(
        \SB2_2_27/Component_Function_2/NAND4_in[3] ), .A4(n3377), .ZN(
        \SB2_2_27/buf_output[2] ) );
  NAND4_X2 U5421 ( .A1(\SB2_1_26/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_1_26/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_26/Component_Function_1/NAND4_in[1] ), .A4(n3378), .ZN(
        \SB2_1_26/buf_output[1] ) );
  XOR2_X1 U5435 ( .A1(\MC_ARK_ARC_1_1/temp5[5] ), .A2(n3380), .Z(\RI1[2][5] )
         );
  XOR2_X1 U5438 ( .A1(\MC_ARK_ARC_1_1/temp3[5] ), .A2(
        \MC_ARK_ARC_1_1/temp4[5] ), .Z(n3380) );
  XOR2_X1 U5446 ( .A1(n4778), .A2(n3381), .Z(n1631) );
  NAND3_X2 U5472 ( .A1(\SB2_1_27/i1[9] ), .A2(\SB2_1_27/i0[6] ), .A3(
        \SB2_1_27/i0_3 ), .ZN(\SB2_1_27/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U5475 ( .A1(\SB1_1_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_3/NAND4_in[2] ), .A4(n4450), .ZN(
        \SB1_1_19/buf_output[3] ) );
  XOR2_X1 U5476 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[56] ), .A2(\RI5[2][20] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[146] ) );
  NAND3_X2 U5477 ( .A1(\SB3_25/i1[9] ), .A2(\SB3_25/i1_7 ), .A3(
        \SB3_25/i0[10] ), .ZN(\SB3_25/Component_Function_3/NAND4_in[2] ) );
  AND2_X1 U5481 ( .A1(\SB3_25/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_25/Component_Function_3/NAND4_in[0] ), .Z(n3386) );
  NAND3_X2 U5482 ( .A1(\SB1_1_13/i0_3 ), .A2(\SB1_1_13/i0[10] ), .A3(
        \SB1_1_13/i0[9] ), .ZN(n3528) );
  XOR2_X1 U5483 ( .A1(n3388), .A2(n3387), .Z(\MC_ARK_ARC_1_2/buf_output[152] )
         );
  XOR2_X1 U5484 ( .A1(n2957), .A2(\MC_ARK_ARC_1_2/temp4[152] ), .Z(n3387) );
  XOR2_X1 U5489 ( .A1(\RI5[1][149] ), .A2(n141), .Z(n3389) );
  XOR2_X1 U5490 ( .A1(\RI5[1][119] ), .A2(\RI5[1][185] ), .Z(n3390) );
  XOR2_X1 U5491 ( .A1(\RI5[0][10] ), .A2(\RI5[0][4] ), .Z(
        \MC_ARK_ARC_1_0/temp1[10] ) );
  XOR2_X1 U5498 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[183] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[15] ), .Z(n3391) );
  NAND4_X2 U5502 ( .A1(\SB1_3_8/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_3_8/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_3_8/Component_Function_0/NAND4_in[1] ), .A4(n3392), .ZN(
        \SB1_3_8/buf_output[0] ) );
  XOR2_X1 U5507 ( .A1(n5408), .A2(n3393), .Z(n1536) );
  XOR2_X1 U5508 ( .A1(\RI5[3][107] ), .A2(\RI5[3][77] ), .Z(n3393) );
  XOR2_X1 U5511 ( .A1(\MC_ARK_ARC_1_0/temp1[75] ), .A2(n3395), .Z(n4981) );
  XOR2_X1 U5512 ( .A1(\SB2_0_26/buf_output[3] ), .A2(\RI5[0][21] ), .Z(n3395)
         );
  INV_X2 U5517 ( .I(\SB1_2_13/buf_output[2] ), .ZN(\SB2_2_10/i1[9] ) );
  NAND3_X1 U5531 ( .A1(\SB4_5/i0_0 ), .A2(\SB4_5/i0_4 ), .A3(\SB4_5/i1_5 ), 
        .ZN(n3398) );
  XOR2_X1 U5541 ( .A1(n3403), .A2(n3402), .Z(\MC_ARK_ARC_1_2/temp6[176] ) );
  XOR2_X1 U5542 ( .A1(\RI5[2][20] ), .A2(n165), .Z(n3402) );
  XOR2_X1 U5543 ( .A1(\RI5[2][50] ), .A2(\RI5[2][86] ), .Z(n3403) );
  XOR2_X1 U5544 ( .A1(n3404), .A2(n101), .Z(Ciphertext[97]) );
  NAND4_X2 U5545 ( .A1(\SB1_1_29/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_29/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_29/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_1_29/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_29/buf_output[1] ) );
  INV_X1 U5549 ( .I(\SB1_3_29/buf_output[1] ), .ZN(\SB2_3_25/i1_7 ) );
  NAND4_X2 U5550 ( .A1(\SB1_3_29/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_3_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_29/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_29/buf_output[1] ) );
  NAND3_X2 U5553 ( .A1(\SB2_1_3/i0_4 ), .A2(\SB2_1_3/i0_0 ), .A3(
        \SB2_1_3/i1_5 ), .ZN(\SB2_1_3/Component_Function_2/NAND4_in[3] ) );
  INV_X2 U5554 ( .I(\SB1_4_25/buf_output[2] ), .ZN(\SB2_4_22/i1[9] ) );
  XOR2_X1 U5566 ( .A1(\RI5[1][191] ), .A2(\RI5[1][137] ), .Z(n3408) );
  NAND4_X2 U5575 ( .A1(\SB2_0_28/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_0_28/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_28/Component_Function_5/NAND4_in[0] ), .A4(n3411), .ZN(
        \SB2_0_28/buf_output[5] ) );
  XOR2_X1 U5576 ( .A1(n3413), .A2(n3412), .Z(n1284) );
  XOR2_X1 U5577 ( .A1(\RI5[2][159] ), .A2(n520), .Z(n3412) );
  BUF_X4 U5590 ( .I(\SB2_4_28/buf_output[3] ), .Z(\RI5[4][33] ) );
  XOR2_X1 U5598 ( .A1(n3417), .A2(n3416), .Z(n3937) );
  XOR2_X1 U5605 ( .A1(\RI5[0][29] ), .A2(n555), .Z(n3416) );
  INV_X1 U5618 ( .I(\SB3_25/buf_output[0] ), .ZN(\SB4_20/i3[0] ) );
  NAND4_X2 U5622 ( .A1(\SB3_25/Component_Function_0/NAND4_in[1] ), .A2(n2929), 
        .A3(\SB3_25/Component_Function_0/NAND4_in[0] ), .A4(
        \SB3_25/Component_Function_0/NAND4_in[2] ), .ZN(\SB3_25/buf_output[0] ) );
  NAND4_X2 U5624 ( .A1(\SB2_3_27/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_27/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_27/Component_Function_4/NAND4_in[3] ), .A4(n3421), .ZN(
        \SB2_3_27/buf_output[4] ) );
  NAND3_X2 U5626 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i0[10] ), .A3(
        \SB2_3_27/i0[9] ), .ZN(n3421) );
  NAND3_X2 U5632 ( .A1(\SB2_0_18/i0[10] ), .A2(\SB2_0_18/i0_3 ), .A3(
        \SB2_0_18/i0[6] ), .ZN(n982) );
  NAND3_X2 U5636 ( .A1(\SB1_1_24/i0[9] ), .A2(\SB1_1_24/i0_4 ), .A3(
        \SB1_1_24/i0[6] ), .ZN(n3422) );
  NAND4_X2 U5638 ( .A1(\SB2_4_31/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_31/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_4_31/Component_Function_0/NAND4_in[2] ), .A4(n3423), .ZN(
        \SB2_4_31/buf_output[0] ) );
  INV_X8 U5647 ( .I(n3425), .ZN(\RI1[3][167] ) );
  INV_X2 U5650 ( .I(\MC_ARK_ARC_1_2/buf_output[167] ), .ZN(n3425) );
  NAND4_X2 U5653 ( .A1(\SB1_4_13/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_4_13/Component_Function_1/NAND4_in[2] ), .A3(n4641), .A4(
        \SB1_4_13/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_4_13/buf_output[1] ) );
  XOR2_X1 U5663 ( .A1(\RI5[3][126] ), .A2(\RI5[3][150] ), .Z(n3428) );
  XOR2_X1 U5665 ( .A1(n3948), .A2(n3834), .Z(n3430) );
  XOR2_X1 U5666 ( .A1(n3432), .A2(n3431), .Z(\MC_ARK_ARC_1_0/temp5[179] ) );
  XOR2_X1 U5669 ( .A1(\RI5[0][125] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[173] ), 
        .Z(n3431) );
  XOR2_X1 U5674 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[149] ), .A2(\RI5[0][179] ), 
        .Z(n3432) );
  XOR2_X1 U5675 ( .A1(\MC_ARK_ARC_1_2/temp5[64] ), .A2(n3433), .Z(
        \MC_ARK_ARC_1_2/buf_output[64] ) );
  XOR2_X1 U5676 ( .A1(\MC_ARK_ARC_1_2/temp4[64] ), .A2(
        \MC_ARK_ARC_1_2/temp3[64] ), .Z(n3433) );
  NAND3_X2 U5684 ( .A1(\SB2_1_28/i0_4 ), .A2(\SB2_1_28/i0_3 ), .A3(
        \SB2_1_28/i0_0 ), .ZN(\SB2_1_28/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U5696 ( .A1(\SB1_0_4/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_4/NAND4_in[0] ), .A4(n3437), .ZN(
        \SB1_0_4/buf_output[4] ) );
  NAND3_X1 U5697 ( .A1(\SB1_0_4/i0_4 ), .A2(\SB1_0_4/i1[9] ), .A3(
        \SB1_0_4/i1_5 ), .ZN(n3437) );
  XOR2_X1 U5707 ( .A1(\MC_ARK_ARC_1_4/temp6[118] ), .A2(n3439), .Z(
        \MC_ARK_ARC_1_4/buf_output[118] ) );
  NAND4_X2 U5709 ( .A1(\SB2_3_19/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_19/Component_Function_1/NAND4_in[0] ), .A3(n4837), .A4(n2239), 
        .ZN(\SB2_3_19/buf_output[1] ) );
  XOR2_X1 U5715 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[32] ), .A2(\RI5[3][56] ), 
        .Z(n3440) );
  BUF_X4 U5717 ( .I(\MC_ARK_ARC_1_3/buf_output[185] ), .Z(\SB1_4_1/i0_3 ) );
  XOR2_X1 U5720 ( .A1(\MC_ARK_ARC_1_3/temp4[61] ), .A2(
        \MC_ARK_ARC_1_3/temp3[61] ), .Z(\MC_ARK_ARC_1_3/temp6[61] ) );
  NAND3_X1 U5730 ( .A1(\SB1_3_23/i0[10] ), .A2(\SB1_3_23/i0_3 ), .A3(
        \SB1_3_23/i0_4 ), .ZN(\SB1_3_23/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 U5733 ( .I(\SB2_3_28/buf_output[0] ), .Z(\RI5[3][48] ) );
  XOR2_X1 U5741 ( .A1(\RI5[0][5] ), .A2(\RI5[0][29] ), .Z(n3445) );
  XOR2_X1 U5742 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[35] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[173] ), .Z(n3446) );
  XOR2_X1 U5743 ( .A1(\RI5[1][64] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[58] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[64] ) );
  NAND3_X1 U5745 ( .A1(\SB4_10/i0_3 ), .A2(\SB4_10/i0[8] ), .A3(\SB4_10/i1_7 ), 
        .ZN(n3447) );
  NAND3_X2 U5746 ( .A1(\SB1_3_21/i0_4 ), .A2(\SB1_3_21/i0_0 ), .A3(
        \SB1_3_21/i1_5 ), .ZN(n3448) );
  NAND4_X2 U5750 ( .A1(\SB1_4_18/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_4_18/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_4_18/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_4_18/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_4_18/buf_output[0] ) );
  XOR2_X1 U5753 ( .A1(n3449), .A2(\MC_ARK_ARC_1_2/temp1[108] ), .Z(
        \MC_ARK_ARC_1_2/temp5[108] ) );
  XOR2_X1 U5754 ( .A1(\RI5[2][54] ), .A2(\RI5[2][78] ), .Z(n3449) );
  XOR2_X1 U5756 ( .A1(n3450), .A2(\MC_ARK_ARC_1_3/temp2[33] ), .Z(
        \MC_ARK_ARC_1_3/temp5[33] ) );
  XOR2_X1 U5757 ( .A1(\RI5[3][33] ), .A2(\RI5[3][27] ), .Z(n3450) );
  CLKBUF_X4 U5766 ( .I(\SB3_0/buf_output[2] ), .Z(\SB4_29/i0_0 ) );
  NAND4_X2 U5781 ( .A1(\SB1_0_22/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_22/Component_Function_0/NAND4_in[0] ), .A4(n3454), .ZN(
        \SB1_0_22/buf_output[0] ) );
  NAND3_X1 U5788 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i0_0 ), .A3(
        \SB1_0_22/i0[7] ), .ZN(n3454) );
  XOR2_X1 U5794 ( .A1(\RI5[1][26] ), .A2(\RI5[1][56] ), .Z(n3456) );
  XOR2_X1 U5797 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[50] ), .A2(\RI5[1][2] ), 
        .Z(n3457) );
  NAND3_X1 U5804 ( .A1(\RI3[0][148] ), .A2(\SB2_0_7/i1_5 ), .A3(
        \SB1_0_10/buf_output[2] ), .ZN(n3460) );
  XOR2_X1 U5820 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[37] ), .A2(\RI5[3][31] ), 
        .Z(n3464) );
  XOR2_X1 U5824 ( .A1(\RI5[2][51] ), .A2(\RI5[2][57] ), .Z(n2411) );
  XOR2_X1 U5825 ( .A1(\RI5[0][117] ), .A2(\RI5[0][81] ), .Z(
        \MC_ARK_ARC_1_0/temp3[15] ) );
  NAND3_X1 U5828 ( .A1(\SB2_0_1/i0_4 ), .A2(\SB2_0_1/i0_0 ), .A3(
        \SB2_0_1/i1_5 ), .ZN(n3466) );
  AND2_X1 U5830 ( .A1(n4568), .A2(n3467), .Z(n4579) );
  NAND3_X1 U5832 ( .A1(\SB1_0_10/i0_3 ), .A2(\SB1_0_10/i0[6] ), .A3(
        \SB1_0_10/i1[9] ), .ZN(n3467) );
  XOR2_X1 U5833 ( .A1(n4194), .A2(n3468), .Z(\MC_ARK_ARC_1_4/buf_output[182] )
         );
  XOR2_X1 U5834 ( .A1(\MC_ARK_ARC_1_4/temp3[182] ), .A2(
        \MC_ARK_ARC_1_4/temp4[182] ), .Z(n3468) );
  BUF_X4 U5835 ( .I(\SB2_4_25/buf_output[2] ), .Z(\RI5[4][56] ) );
  XOR2_X1 U5848 ( .A1(n3471), .A2(n163), .Z(Ciphertext[35]) );
  NAND4_X2 U5849 ( .A1(\SB4_26/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_26/Component_Function_5/NAND4_in[2] ), .A3(n960), .A4(
        \SB4_26/Component_Function_5/NAND4_in[0] ), .ZN(n3471) );
  INV_X2 U5867 ( .I(\SB1_4_21/buf_output[2] ), .ZN(\SB2_4_18/i1[9] ) );
  NAND3_X2 U5873 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i1[9] ), .A3(\SB3_1/i0[6] ), 
        .ZN(\SB3_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U5878 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i1[9] ), .A3(
        \SB4_10/i1_5 ), .ZN(n3477) );
  XOR2_X1 U5880 ( .A1(n3478), .A2(n2161), .Z(\MC_ARK_ARC_1_4/temp6[185] ) );
  NAND4_X2 U5883 ( .A1(\SB2_1_0/Component_Function_2/NAND4_in[2] ), .A2(n4270), 
        .A3(\SB2_1_0/Component_Function_2/NAND4_in[3] ), .A4(n3479), .ZN(
        \SB2_1_0/buf_output[2] ) );
  NAND3_X2 U5888 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i1_5 ), .A3(
        \SB2_1_0/i1[9] ), .ZN(n3479) );
  XOR2_X1 U5894 ( .A1(\RI5[0][160] ), .A2(\RI5[0][166] ), .Z(
        \MC_ARK_ARC_1_0/temp1[166] ) );
  NAND3_X1 U5903 ( .A1(\SB3_12/i0_0 ), .A2(\SB3_12/i0_4 ), .A3(\RI1[5][119] ), 
        .ZN(n3480) );
  XOR2_X1 U5905 ( .A1(\MC_ARK_ARC_1_1/temp5[84] ), .A2(n3481), .Z(
        \MC_ARK_ARC_1_1/buf_output[84] ) );
  XOR2_X1 U5907 ( .A1(\MC_ARK_ARC_1_1/temp4[84] ), .A2(
        \MC_ARK_ARC_1_1/temp3[84] ), .Z(n3481) );
  NAND3_X1 U5911 ( .A1(\SB2_1_27/i0_3 ), .A2(\SB2_1_27/i0[10] ), .A3(
        \SB2_1_27/i0_4 ), .ZN(\SB2_1_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U5920 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i0_0 ), .A3(
        \SB2_1_4/i0[7] ), .ZN(n4898) );
  XOR2_X1 U5933 ( .A1(\MC_ARK_ARC_1_1/temp2[159] ), .A2(n610), .Z(n3484) );
  XOR2_X1 U5937 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[184] ), .A2(\RI5[3][22] ), 
        .Z(n4030) );
  INV_X1 U5942 ( .I(\SB1_2_13/buf_output[0] ), .ZN(\SB2_2_8/i3[0] ) );
  NAND4_X2 U5946 ( .A1(\SB1_2_13/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_13/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_13/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_13/buf_output[0] ) );
  XOR2_X1 U5949 ( .A1(\MC_ARK_ARC_1_4/temp1[41] ), .A2(n3609), .Z(n3485) );
  XOR2_X1 U5950 ( .A1(\RI5[1][35] ), .A2(\RI5[1][41] ), .Z(n3486) );
  XOR2_X1 U5956 ( .A1(n3076), .A2(\MC_ARK_ARC_1_2/temp6[63] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[63] ) );
  NAND3_X1 U5961 ( .A1(\SB4_0/i1_5 ), .A2(\SB4_0/i3[0] ), .A3(\SB4_0/i0[8] ), 
        .ZN(\SB4_0/Component_Function_3/NAND4_in[3] ) );
  INV_X2 U5972 ( .I(\RI3[0][9] ), .ZN(\SB2_0_30/i0[8] ) );
  NAND4_X2 U5973 ( .A1(n1512), .A2(\SB1_0_0/Component_Function_3/NAND4_in[0] ), 
        .A3(n1169), .A4(\SB1_0_0/Component_Function_3/NAND4_in[3] ), .ZN(
        \RI3[0][9] ) );
  NAND3_X1 U5974 ( .A1(\SB2_1_7/i0[10] ), .A2(\SB2_1_7/i0_4 ), .A3(
        \SB2_1_7/i0_3 ), .ZN(\SB2_1_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U5980 ( .A1(\SB2_2_7/i0[10] ), .A2(\SB2_2_7/i1_5 ), .A3(
        \SB2_2_7/i1[9] ), .ZN(\SB2_2_7/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U5983 ( .A1(n4142), .A2(n3489), .Z(n3506) );
  XOR2_X1 U5984 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[152] ), .A2(\RI5[1][158] ), 
        .Z(n3489) );
  NAND4_X2 U5988 ( .A1(\SB2_1_0/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_0/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_0/Component_Function_1/NAND4_in[2] ), .A4(n3490), .ZN(
        \SB2_1_0/buf_output[1] ) );
  NAND3_X2 U5991 ( .A1(n590), .A2(\SB2_1_0/i1_7 ), .A3(\SB2_1_0/i0[8] ), .ZN(
        n3490) );
  XOR2_X1 U5997 ( .A1(\RI5[1][70] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[94] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[124] ) );
  XOR2_X1 U6015 ( .A1(n3495), .A2(n3494), .Z(\MC_ARK_ARC_1_3/buf_output[134] )
         );
  XOR2_X1 U6018 ( .A1(\MC_ARK_ARC_1_3/temp1[134] ), .A2(
        \MC_ARK_ARC_1_3/temp4[134] ), .Z(n3494) );
  XOR2_X1 U6020 ( .A1(n3497), .A2(n3496), .Z(\MC_ARK_ARC_1_4/temp5[14] ) );
  XOR2_X1 U6028 ( .A1(\RI5[4][14] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[176] ), 
        .Z(n3496) );
  XOR2_X1 U6029 ( .A1(\RI5[4][152] ), .A2(\RI5[4][8] ), .Z(n3497) );
  XOR2_X1 U6045 ( .A1(\RI5[1][5] ), .A2(\RI5[1][29] ), .Z(n3499) );
  NAND3_X1 U6048 ( .A1(\SB2_3_7/i0[10] ), .A2(\SB2_3_7/i0_3 ), .A3(
        \SB2_3_7/i0[9] ), .ZN(n3500) );
  BUF_X4 U6049 ( .I(\MC_ARK_ARC_1_3/buf_output[154] ), .Z(\SB1_4_6/i0_4 ) );
  XOR2_X1 U6055 ( .A1(n1014), .A2(\MC_ARK_ARC_1_3/temp4[135] ), .Z(n3501) );
  NAND3_X1 U6059 ( .A1(\SB2_1_28/i0[6] ), .A2(\SB2_1_28/i1_5 ), .A3(
        \SB2_1_28/i0[9] ), .ZN(\SB2_1_28/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U6063 ( .A1(\SB2_2_4/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_4/Component_Function_1/NAND4_in[2] ), .A4(n3503), .ZN(
        \SB2_2_4/buf_output[1] ) );
  NAND2_X1 U6065 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i1[9] ), .ZN(n3503) );
  NAND4_X2 U6089 ( .A1(n3522), .A2(\SB1_4_25/Component_Function_0/NAND4_in[2] ), .A3(n1902), .A4(\SB1_4_25/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_4_25/buf_output[0] ) );
  NAND4_X2 U6101 ( .A1(\SB1_4_10/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_4_10/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_4_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_4_10/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_4_10/buf_output[1] ) );
  NAND3_X1 U6109 ( .A1(\SB2_0_27/i0[6] ), .A2(\RI3[0][28] ), .A3(
        \SB2_0_27/i0[9] ), .ZN(n1454) );
  NAND4_X2 U6118 ( .A1(\SB2_0_27/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_27/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_0_27/Component_Function_0/NAND4_in[2] ), .A4(n3507), .ZN(
        \SB2_0_27/buf_output[0] ) );
  NAND3_X1 U6119 ( .A1(\SB1_0_0/i0[10] ), .A2(\SB1_0_0/i1_5 ), .A3(
        \SB1_0_0/i1[9] ), .ZN(\SB1_0_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U6122 ( .A1(\SB2_2_17/i3[0] ), .A2(\SB2_2_17/i1_5 ), .A3(
        \SB2_2_17/i0[8] ), .ZN(n3508) );
  XOR2_X1 U6126 ( .A1(\MC_ARK_ARC_1_1/temp4[90] ), .A2(
        \MC_ARK_ARC_1_1/temp3[90] ), .Z(n3509) );
  XOR2_X1 U6127 ( .A1(\MC_ARK_ARC_1_2/temp4[50] ), .A2(n3511), .Z(n4699) );
  XOR2_X1 U6129 ( .A1(\RI5[2][188] ), .A2(\RI5[2][20] ), .Z(n3511) );
  XOR2_X1 U6134 ( .A1(\MC_ARK_ARC_1_4/temp2[120] ), .A2(
        \MC_ARK_ARC_1_4/temp1[120] ), .Z(\MC_ARK_ARC_1_4/temp5[120] ) );
  NAND4_X2 U6135 ( .A1(\SB2_4_24/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_4_24/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_4_24/Component_Function_4/NAND4_in[0] ), .A4(n3513), .ZN(
        \SB2_4_24/buf_output[4] ) );
  NAND4_X2 U6139 ( .A1(\SB1_2_6/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_6/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_6/Component_Function_2/NAND4_in[2] ), .A4(n3515), .ZN(
        \SB1_2_6/buf_output[2] ) );
  NAND3_X2 U6142 ( .A1(\SB1_2_6/i0_0 ), .A2(\SB1_2_6/i0_4 ), .A3(
        \SB1_2_6/i1_5 ), .ZN(n3515) );
  XOR2_X1 U6148 ( .A1(\RI5[0][60] ), .A2(\RI5[0][96] ), .Z(
        \MC_ARK_ARC_1_0/temp3[186] ) );
  NAND4_X2 U6151 ( .A1(\SB2_0_11/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_11/Component_Function_4/NAND4_in[0] ), .A3(n4193), .A4(n3518), 
        .ZN(\SB2_0_11/buf_output[4] ) );
  NAND3_X1 U6157 ( .A1(\SB2_0_11/i0_0 ), .A2(\SB2_0_11/i3[0] ), .A3(
        \SB2_0_11/i1_7 ), .ZN(n3518) );
  NAND2_X2 U6177 ( .A1(\SB2_0_21/i0_0 ), .A2(n3171), .ZN(
        \SB2_0_21/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U6178 ( .A1(\SB1_1_30/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_1_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_1/NAND4_in[0] ), .A4(n1718), .ZN(
        \SB1_1_30/buf_output[1] ) );
  NAND3_X1 U6192 ( .A1(\SB4_15/i0_3 ), .A2(\SB4_15/i0[6] ), .A3(\SB4_15/i1[9] ), .ZN(n2663) );
  NAND4_X2 U6194 ( .A1(\SB2_1_24/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_24/Component_Function_1/NAND4_in[2] ), .A3(n1936), .A4(
        \SB2_1_24/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_24/buf_output[1] ) );
  BUF_X4 U6198 ( .I(\SB2_3_31/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[15] ) );
  NAND4_X2 U6203 ( .A1(\SB1_1_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_25/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_1_25/Component_Function_2/NAND4_in[1] ), .A4(n766), .ZN(
        \SB1_1_25/buf_output[2] ) );
  XOR2_X1 U6213 ( .A1(\RI5[3][41] ), .A2(\RI5[3][35] ), .Z(n2193) );
  NAND3_X1 U6215 ( .A1(\SB1_3_0/i0[10] ), .A2(\SB1_3_0/i1_7 ), .A3(
        \SB1_3_0/i1[9] ), .ZN(\SB1_3_0/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U6218 ( .A1(\RI5[3][179] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[143] ), 
        .Z(n2741) );
  XOR2_X1 U6221 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[44] ), .A2(n3167), .Z(
        n1268) );
  NAND3_X2 U6223 ( .A1(\SB1_0_9/i0_3 ), .A2(\SB1_0_9/i0_4 ), .A3(
        \SB1_0_9/i1[9] ), .ZN(\SB1_0_9/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U6230 ( .A1(\SB2_1_29/i0_3 ), .A2(\SB2_1_29/i0_4 ), .A3(
        \SB2_1_29/i1[9] ), .ZN(\SB2_1_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U6231 ( .A1(\SB2_0_1/i0[10] ), .A2(\SB2_0_1/i0_3 ), .A3(
        \SB2_0_1/i0[6] ), .ZN(\SB2_0_1/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U6232 ( .A1(n685), .A2(n3956), .Z(\MC_ARK_ARC_1_3/buf_output[32] )
         );
  NAND4_X2 U6247 ( .A1(n3734), .A2(\SB1_1_27/Component_Function_4/NAND4_in[2] ), .A3(\SB1_1_27/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_1_27/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB1_1_27/buf_output[4] ) );
  NAND3_X2 U6248 ( .A1(\SB2_3_25/i0[10] ), .A2(\SB2_3_25/i0_0 ), .A3(
        \SB2_3_25/i0[6] ), .ZN(\SB2_3_25/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U6259 ( .A1(\MC_ARK_ARC_1_2/temp2[92] ), .A2(n3519), .Z(n5395) );
  XOR2_X1 U6263 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[92] ), .A2(\RI5[2][86] ), 
        .Z(n3519) );
  XOR2_X1 U6266 ( .A1(\MC_ARK_ARC_1_0/temp5[140] ), .A2(n3521), .Z(
        \MC_ARK_ARC_1_0/buf_output[140] ) );
  NAND4_X2 U6269 ( .A1(\SB2_4_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_4_3/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_4_3/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_4_3/buf_output[4] ) );
  INV_X2 U6271 ( .I(\SB1_1_16/buf_output[1] ), .ZN(\SB2_1_12/i1_7 ) );
  NAND3_X2 U6278 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i1[9] ), .A3(
        \SB1_3_2/i1_7 ), .ZN(n3523) );
  NAND4_X2 U6279 ( .A1(\SB1_3_28/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_3_28/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_28/Component_Function_3/NAND4_in[1] ), .A4(n3524), .ZN(
        \SB1_3_28/buf_output[3] ) );
  NAND3_X2 U6283 ( .A1(\SB1_3_28/i0[8] ), .A2(\SB1_3_28/i3[0] ), .A3(
        \SB1_3_28/i1_5 ), .ZN(n3524) );
  NAND4_X2 U6286 ( .A1(\SB2_2_7/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_7/Component_Function_0/NAND4_in[2] ), .A3(n976), .A4(
        \SB2_2_7/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_7/buf_output[0] ) );
  NAND3_X2 U6288 ( .A1(\SB1_0_21/i0_0 ), .A2(\SB1_0_21/i1_5 ), .A3(
        \SB1_0_21/i0_4 ), .ZN(n5122) );
  XOR2_X1 U6290 ( .A1(n3147), .A2(n3525), .Z(n1047) );
  XOR2_X1 U6294 ( .A1(\RI5[0][165] ), .A2(\RI5[0][171] ), .Z(n3525) );
  XOR2_X1 U6295 ( .A1(n3526), .A2(\MC_ARK_ARC_1_4/temp1[150] ), .Z(
        \MC_ARK_ARC_1_4/temp5[150] ) );
  NAND4_X2 U6301 ( .A1(\SB2_4_16/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_16/Component_Function_0/NAND4_in[0] ), .A4(n3527), .ZN(
        \SB2_4_16/buf_output[0] ) );
  NAND4_X2 U6305 ( .A1(\SB1_1_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_4/NAND4_in[3] ), .A4(n3528), .ZN(
        \SB1_1_13/buf_output[4] ) );
  XOR2_X1 U6317 ( .A1(n3530), .A2(\MC_ARK_ARC_1_1/temp6[145] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[145] ) );
  XOR2_X1 U6320 ( .A1(\MC_ARK_ARC_1_1/temp1[145] ), .A2(
        \MC_ARK_ARC_1_1/temp2[145] ), .Z(n3530) );
  XOR2_X1 U6322 ( .A1(\MC_ARK_ARC_1_1/temp5[58] ), .A2(
        \MC_ARK_ARC_1_1/temp6[58] ), .Z(\MC_ARK_ARC_1_1/buf_output[58] ) );
  XOR2_X1 U6327 ( .A1(n1819), .A2(\MC_ARK_ARC_1_3/temp1[77] ), .Z(n3532) );
  NAND4_X2 U6333 ( .A1(n3535), .A2(n3534), .A3(
        \SB2_0_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_22/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_22/buf_output[0] ) );
  XOR2_X1 U6339 ( .A1(\RI5[1][186] ), .A2(\RI5[1][138] ), .Z(n2211) );
  XOR2_X1 U6341 ( .A1(\MC_ARK_ARC_1_2/temp1[184] ), .A2(n3537), .Z(
        \MC_ARK_ARC_1_2/temp5[184] ) );
  XOR2_X1 U6342 ( .A1(\RI5[2][130] ), .A2(\RI5[2][154] ), .Z(n3537) );
  NAND3_X2 U6344 ( .A1(\SB1_4_12/i0[9] ), .A2(\RI1[4][119] ), .A3(
        \SB1_4_12/i0[10] ), .ZN(n1928) );
  XOR2_X1 U6355 ( .A1(n3540), .A2(n3539), .Z(n4439) );
  XOR2_X1 U6356 ( .A1(\RI5[0][20] ), .A2(n499), .Z(n3539) );
  XOR2_X1 U6362 ( .A1(\RI5[0][86] ), .A2(\RI5[0][50] ), .Z(n3540) );
  NAND3_X1 U6363 ( .A1(\SB1_1_21/i0_3 ), .A2(\MC_ARK_ARC_1_0/buf_output[64] ), 
        .A3(\SB1_1_21/i1[9] ), .ZN(n3065) );
  XOR2_X1 U6366 ( .A1(n3542), .A2(n818), .Z(n4123) );
  XOR2_X1 U6367 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[65] ), .Z(n3542) );
  XOR2_X1 U6370 ( .A1(\RI5[1][41] ), .A2(n33), .Z(n3543) );
  XOR2_X1 U6371 ( .A1(\RI5[1][77] ), .A2(\RI5[1][11] ), .Z(n3544) );
  XOR2_X1 U6376 ( .A1(\MC_ARK_ARC_1_3/temp1[116] ), .A2(
        \MC_ARK_ARC_1_3/temp2[116] ), .Z(\MC_ARK_ARC_1_3/temp5[116] ) );
  XOR2_X1 U6386 ( .A1(\RI5[3][137] ), .A2(\RI5[3][173] ), .Z(n3546) );
  NAND4_X2 U6414 ( .A1(\SB1_2_3/Component_Function_2/NAND4_in[0] ), .A2(n1234), 
        .A3(\SB1_2_3/Component_Function_2/NAND4_in[1] ), .A4(n3552), .ZN(
        \SB1_2_3/buf_output[2] ) );
  NAND3_X1 U6415 ( .A1(\SB1_2_3/i0_0 ), .A2(\MC_ARK_ARC_1_1/buf_output[172] ), 
        .A3(\SB1_2_3/i1_5 ), .ZN(n3552) );
  NAND4_X2 U6417 ( .A1(\SB1_4_12/Component_Function_5/NAND4_in[1] ), .A2(n3907), .A3(\SB1_4_12/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_4_12/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_4_12/buf_output[5] ) );
  NAND3_X2 U6419 ( .A1(\SB2_1_14/i0_0 ), .A2(\SB2_1_14/i0_4 ), .A3(
        \SB2_1_14/i1_5 ), .ZN(n1082) );
  NAND3_X1 U6420 ( .A1(\SB1_0_10/i0_3 ), .A2(n295), .A3(\SB1_0_10/i0[8] ), 
        .ZN(\SB1_0_10/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U6425 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[23] ), .A2(\RI5[4][191] ), 
        .Z(n1259) );
  NAND3_X2 U6432 ( .A1(\SB1_3_0/i0_4 ), .A2(\SB1_3_0/i0[9] ), .A3(
        \SB1_3_0/i0[6] ), .ZN(n5278) );
  NAND3_X1 U6435 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i0_4 ), .A3(\SB4_28/i0[10] ), .ZN(\SB4_28/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U6445 ( .A1(\SB2_1_27/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_1_27/Component_Function_3/NAND4_in[0] ), .A3(n1680), .A4(
        \SB2_1_27/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_27/buf_output[3] ) );
  BUF_X4 U6451 ( .I(\SB1_4_20/buf_output[5] ), .Z(\SB2_4_20/i0_3 ) );
  NAND4_X2 U6454 ( .A1(\SB2_3_0/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_0/Component_Function_0/NAND4_in[2] ), .A3(n4064), .A4(
        \SB2_3_0/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_0/buf_output[0] ) );
  INV_X2 U6465 ( .I(\SB1_2_22/buf_output[3] ), .ZN(\SB2_2_20/i0[8] ) );
  XOR2_X1 U6469 ( .A1(\RI5[0][90] ), .A2(\RI5[0][114] ), .Z(
        \MC_ARK_ARC_1_0/temp2[144] ) );
  XOR2_X1 U6476 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[129] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[165] ), .Z(\MC_ARK_ARC_1_4/temp3[63] )
         );
  NAND4_X2 U6477 ( .A1(\SB2_2_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_18/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_18/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_18/buf_output[5] ) );
  XOR2_X1 U6479 ( .A1(\MC_ARK_ARC_1_1/temp4[136] ), .A2(
        \MC_ARK_ARC_1_1/temp3[136] ), .Z(\MC_ARK_ARC_1_1/temp6[136] ) );
  XOR2_X1 U6480 ( .A1(\MC_ARK_ARC_1_2/temp5[131] ), .A2(
        \MC_ARK_ARC_1_2/temp6[131] ), .Z(\MC_ARK_ARC_1_2/buf_output[131] ) );
  XOR2_X1 U6487 ( .A1(\RI5[3][35] ), .A2(\RI5[3][191] ), .Z(
        \MC_ARK_ARC_1_3/temp3[125] ) );
  XOR2_X1 U6488 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[39] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[15] ), .Z(n1223) );
  XOR2_X1 U6491 ( .A1(\RI5[2][182] ), .A2(\RI5[2][26] ), .Z(
        \MC_ARK_ARC_1_2/temp3[116] ) );
  XOR2_X1 U6494 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[158] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[182] ), .Z(\MC_ARK_ARC_1_3/temp2[20] )
         );
  NAND4_X2 U6500 ( .A1(\SB1_1_7/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_7/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_7/Component_Function_4/NAND4_in[3] ), .A4(n3553), .ZN(
        \SB1_1_7/buf_output[4] ) );
  XOR2_X1 U6511 ( .A1(\MC_ARK_ARC_1_2/temp3[47] ), .A2(
        \MC_ARK_ARC_1_2/temp4[47] ), .Z(n1355) );
  NAND3_X1 U6516 ( .A1(\SB2_4_12/i0_3 ), .A2(\SB2_4_12/i0[6] ), .A3(
        \SB2_4_12/i1[9] ), .ZN(\SB2_4_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U6519 ( .A1(\SB1_1_7/i0[9] ), .A2(\SB1_1_7/i0_3 ), .A3(
        \SB1_1_7/i0[8] ), .ZN(\SB1_1_7/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U6523 ( .A1(\SB1_4_3/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_4_3/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_4_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_3/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_4_3/buf_output[0] ) );
  NAND3_X1 U6528 ( .A1(\SB2_4_30/i0[9] ), .A2(\SB2_4_30/i0[10] ), .A3(
        \SB2_4_30/i0_3 ), .ZN(\SB2_4_30/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U6534 ( .A1(n3082), .A2(\SB2_2_25/Component_Function_3/NAND4_in[0] ), .A3(n4976), .A4(\SB2_2_25/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_25/buf_output[3] ) );
  XOR2_X1 U6553 ( .A1(n3735), .A2(n3556), .Z(\MC_ARK_ARC_1_0/temp5[167] ) );
  XOR2_X1 U6567 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[113] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[137] ), .Z(n3556) );
  NAND4_X2 U6570 ( .A1(\SB1_2_29/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_29/Component_Function_3/NAND4_in[2] ), .A3(n2132), .A4(n3557), 
        .ZN(\SB1_2_29/buf_output[3] ) );
  NAND3_X2 U6571 ( .A1(\SB1_2_29/i0[6] ), .A2(\SB1_2_29/i1[9] ), .A3(
        \RI1[2][17] ), .ZN(n3557) );
  NAND3_X2 U6574 ( .A1(\SB1_1_27/i0[10] ), .A2(\SB1_1_27/i1[9] ), .A3(
        \SB1_1_27/i1_5 ), .ZN(\SB1_1_27/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U6602 ( .A1(n3561), .A2(\MC_ARK_ARC_1_2/temp1[84] ), .Z(
        \MC_ARK_ARC_1_2/temp5[84] ) );
  XOR2_X1 U6603 ( .A1(\RI5[2][30] ), .A2(\RI5[2][54] ), .Z(n3561) );
  NAND4_X2 U6609 ( .A1(\SB1_4_22/Component_Function_3/NAND4_in[0] ), .A2(n4301), .A3(\SB1_4_22/Component_Function_3/NAND4_in[2] ), .A4(n3563), .ZN(
        \SB1_4_22/buf_output[3] ) );
  XOR2_X1 U6613 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[39] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[63] ), .Z(\MC_ARK_ARC_1_4/temp2[93] ) );
  NOR2_X2 U6641 ( .A1(n4099), .A2(n3568), .ZN(\SB2_0_4/i0[7] ) );
  XOR2_X1 U6662 ( .A1(\MC_ARK_ARC_1_0/temp4[3] ), .A2(
        \MC_ARK_ARC_1_0/temp3[3] ), .Z(\MC_ARK_ARC_1_0/temp6[3] ) );
  XOR2_X1 U6667 ( .A1(\MC_ARK_ARC_1_2/temp4[180] ), .A2(n3570), .Z(
        \MC_ARK_ARC_1_2/temp6[180] ) );
  XOR2_X1 U6668 ( .A1(\SB2_2_27/buf_output[0] ), .A2(\SB2_2_21/buf_output[0] ), 
        .Z(n3570) );
  XOR2_X1 U6675 ( .A1(\RI5[4][139] ), .A2(\RI5[4][163] ), .Z(n3573) );
  INV_X1 U6676 ( .I(\SB3_31/buf_output[5] ), .ZN(\SB4_31/i1_5 ) );
  NAND4_X2 U6677 ( .A1(n4751), .A2(\SB3_31/Component_Function_5/NAND4_in[2] ), 
        .A3(n3800), .A4(\SB3_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_31/buf_output[5] ) );
  XOR2_X1 U6679 ( .A1(n1935), .A2(n3574), .Z(\MC_ARK_ARC_1_1/buf_output[29] )
         );
  XOR2_X1 U6685 ( .A1(\MC_ARK_ARC_1_2/temp5[149] ), .A2(n3576), .Z(
        \MC_ARK_ARC_1_2/buf_output[149] ) );
  XOR2_X1 U6687 ( .A1(\MC_ARK_ARC_1_2/temp3[149] ), .A2(
        \MC_ARK_ARC_1_2/temp4[149] ), .Z(n3576) );
  NAND2_X2 U6700 ( .A1(n2890), .A2(n3173), .ZN(\SB2_0_9/i0_0 ) );
  NAND3_X2 U6701 ( .A1(\SB1_0_0/i0_4 ), .A2(\SB1_0_0/i0[10] ), .A3(
        \SB1_0_0/i0_3 ), .ZN(n3579) );
  NAND3_X2 U6713 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i0_4 ), .A3(
        \SB1_3_27/i1_5 ), .ZN(n3580) );
  XOR2_X1 U6716 ( .A1(n3581), .A2(\MC_ARK_ARC_1_2/temp2[20] ), .Z(
        \MC_ARK_ARC_1_2/temp5[20] ) );
  XOR2_X1 U6720 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[14] ), .A2(\RI5[2][20] ), 
        .Z(n3581) );
  NAND3_X2 U6721 ( .A1(\SB2_1_29/i0[10] ), .A2(\SB2_1_29/i1[9] ), .A3(
        \SB2_1_29/i1_7 ), .ZN(\SB2_1_29/Component_Function_3/NAND4_in[2] ) );
  INV_X4 U6722 ( .I(\SB2_1_0/i0[7] ), .ZN(n590) );
  NOR2_X2 U6724 ( .A1(n648), .A2(n646), .ZN(\SB2_1_0/i0[7] ) );
  NAND3_X1 U6726 ( .A1(\SB2_0_7/i0_0 ), .A2(\SB2_0_7/i0[9] ), .A3(
        \SB2_0_7/i0[8] ), .ZN(\SB2_0_7/Component_Function_4/NAND4_in[0] ) );
  BUF_X4 U6739 ( .I(\SB1_3_13/buf_output[5] ), .Z(\SB2_3_13/i0_3 ) );
  NAND4_X2 U6753 ( .A1(\SB2_0_10/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_0_10/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_10/Component_Function_5/NAND4_in[0] ), .A4(n3583), .ZN(
        \SB2_0_10/buf_output[5] ) );
  NAND4_X2 U6761 ( .A1(\SB1_1_11/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_1_11/Component_Function_1/NAND4_in[1] ), .A3(n3721), .A4(
        \SB1_1_11/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_11/buf_output[1] ) );
  XOR2_X1 U6786 ( .A1(\RI5[0][110] ), .A2(\RI5[0][134] ), .Z(
        \MC_ARK_ARC_1_0/temp2[164] ) );
  NAND3_X2 U6788 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0[10] ), .A3(
        \SB2_2_16/i0[6] ), .ZN(n3584) );
  NAND3_X2 U6792 ( .A1(\SB1_0_19/i0[10] ), .A2(\SB1_0_19/i0_3 ), .A3(
        \SB1_0_19/i0[6] ), .ZN(n3585) );
  NAND4_X2 U6793 ( .A1(\SB1_3_4/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_3_4/Component_Function_3/NAND4_in[0] ), .A3(n2968), .A4(n3586), 
        .ZN(\SB1_3_4/buf_output[3] ) );
  NAND3_X2 U6794 ( .A1(\SB1_3_4/i0_0 ), .A2(\SB1_3_4/i0_4 ), .A3(\RI1[3][167] ), .ZN(n3586) );
  XOR2_X1 U6801 ( .A1(\RI5[1][95] ), .A2(\RI5[1][89] ), .Z(n3588) );
  XOR2_X1 U6802 ( .A1(\RI5[0][106] ), .A2(\RI5[0][142] ), .Z(
        \MC_ARK_ARC_1_0/temp3[40] ) );
  INV_X2 U6820 ( .I(\RI3[0][86] ), .ZN(\SB2_0_17/i1[9] ) );
  XOR2_X1 U6840 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[39] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[3] ), .Z(\MC_ARK_ARC_1_4/temp3[129] ) );
  NAND4_X2 U6842 ( .A1(\SB2_3_26/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_26/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_26/Component_Function_0/NAND4_in[0] ), .A4(n3596), .ZN(
        \SB2_3_26/buf_output[0] ) );
  XOR2_X1 U6846 ( .A1(\RI5[3][135] ), .A2(\RI5[3][171] ), .Z(
        \MC_ARK_ARC_1_3/temp3[69] ) );
  NAND4_X2 U6848 ( .A1(\SB2_1_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_23/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_23/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_1_23/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_23/buf_output[1] ) );
  INV_X2 U6850 ( .I(\SB1_4_30/buf_output[2] ), .ZN(\SB2_4_27/i1[9] ) );
  XOR2_X1 U6861 ( .A1(\MC_ARK_ARC_1_0/temp3[66] ), .A2(
        \MC_ARK_ARC_1_0/temp4[66] ), .Z(n3597) );
  BUF_X4 U6863 ( .I(\SB2_4_27/buf_output[5] ), .Z(\RI5[4][29] ) );
  NAND4_X2 U6866 ( .A1(\SB3_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_5/Component_Function_3/NAND4_in[2] ), .A3(
        \SB3_5/Component_Function_3/NAND4_in[1] ), .A4(n3598), .ZN(
        \RI3[5][171] ) );
  XOR2_X1 U6879 ( .A1(\MC_ARK_ARC_1_3/temp1[75] ), .A2(n2629), .Z(
        \MC_ARK_ARC_1_3/temp5[75] ) );
  NAND3_X1 U6888 ( .A1(\SB3_21/i0[6] ), .A2(\SB3_21/i0[8] ), .A3(
        \SB3_21/i0[7] ), .ZN(\SB3_21/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U6891 ( .A1(\MC_ARK_ARC_1_4/temp6[156] ), .A2(
        \MC_ARK_ARC_1_4/temp5[156] ), .Z(\MC_ARK_ARC_1_4/buf_output[156] ) );
  XOR2_X1 U6917 ( .A1(\MC_ARK_ARC_1_0/temp4[165] ), .A2(n3605), .Z(n4625) );
  XOR2_X1 U6918 ( .A1(\RI5[0][159] ), .A2(\RI5[0][165] ), .Z(n3605) );
  NAND3_X2 U6925 ( .A1(\SB2_4_23/i0_3 ), .A2(\SB2_4_23/i1[9] ), .A3(
        \SB2_4_23/i0_4 ), .ZN(n4784) );
  INV_X1 U6929 ( .I(\SB3_15/buf_output[5] ), .ZN(\SB4_15/i1_5 ) );
  XOR2_X1 U6930 ( .A1(\MC_ARK_ARC_1_4/temp1[33] ), .A2(n3608), .Z(n2779) );
  XOR2_X1 U6933 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[171] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[3] ), .Z(n3608) );
  XOR2_X1 U6936 ( .A1(\RI5[4][179] ), .A2(\RI5[4][11] ), .Z(n3609) );
  NAND4_X2 U6942 ( .A1(\SB1_2_5/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_5/Component_Function_5/NAND4_in[1] ), .A3(n2857), .A4(n3611), 
        .ZN(\SB1_2_5/buf_output[5] ) );
  NAND2_X2 U6945 ( .A1(\SB1_2_5/i0_0 ), .A2(\SB1_2_5/i3[0] ), .ZN(n3611) );
  BUF_X4 U6953 ( .I(n260), .Z(\SB1_0_28/i0_0 ) );
  XOR2_X1 U6970 ( .A1(\MC_ARK_ARC_1_2/temp5[85] ), .A2(n790), .Z(
        \MC_ARK_ARC_1_2/buf_output[85] ) );
  XOR2_X1 U6973 ( .A1(n5412), .A2(\MC_ARK_ARC_1_1/temp5[161] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[161] ) );
  NAND3_X1 U6985 ( .A1(\SB4_29/i0[6] ), .A2(\SB4_29/i0[8] ), .A3(
        \SB4_29/i0[7] ), .ZN(\SB4_29/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U6996 ( .A1(n2274), .A2(\SB2_3_7/Component_Function_0/NAND4_in[3] ), 
        .A3(\SB2_3_7/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_3_7/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_3_7/buf_output[0] ) );
  NAND4_X2 U7001 ( .A1(\SB1_1_29/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_29/Component_Function_5/NAND4_in[2] ), .A3(n4596), .A4(
        \SB1_1_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_29/buf_output[5] ) );
  NAND4_X2 U7007 ( .A1(\SB3_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_3/NAND4_in[1] ), .A3(n5064), .A4(n3137), 
        .ZN(\SB3_31/buf_output[3] ) );
  NAND4_X2 U7008 ( .A1(\SB1_1_23/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_23/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_1_23/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_23/buf_output[0] ) );
  XOR2_X1 U7014 ( .A1(\RI5[0][116] ), .A2(\RI5[0][80] ), .Z(
        \MC_ARK_ARC_1_0/temp3[14] ) );
  NAND4_X2 U7019 ( .A1(\SB3_21/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_21/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_21/Component_Function_4/NAND4_in[1] ), .A4(n3613), .ZN(
        \SB3_21/buf_output[4] ) );
  NAND3_X1 U7020 ( .A1(\SB3_21/i0_4 ), .A2(\SB3_21/i1[9] ), .A3(n3182), .ZN(
        n3613) );
  NAND4_X2 U7022 ( .A1(\SB2_2_0/Component_Function_1/NAND4_in[2] ), .A2(n1630), 
        .A3(\SB2_2_0/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_2_0/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_0/buf_output[1] ) );
  NAND3_X1 U7023 ( .A1(\SB2_4_2/i0_3 ), .A2(\SB2_4_2/i0[10] ), .A3(
        \SB2_4_2/i0_4 ), .ZN(\SB2_4_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U7053 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0[10] ), .A3(
        \SB2_2_25/i0[6] ), .ZN(\SB2_2_25/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U7065 ( .I(\SB1_1_21/buf_output[3] ), .ZN(\SB2_1_19/i0[8] ) );
  NAND4_X2 U7069 ( .A1(\SB1_1_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_21/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_1_21/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_1_21/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_21/buf_output[3] ) );
  XOR2_X1 U7082 ( .A1(n3617), .A2(\MC_ARK_ARC_1_2/temp1[49] ), .Z(
        \MC_ARK_ARC_1_2/temp5[49] ) );
  XOR2_X1 U7085 ( .A1(\RI5[2][187] ), .A2(\RI5[2][19] ), .Z(n3617) );
  NAND4_X2 U7108 ( .A1(\SB1_3_23/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_23/Component_Function_5/NAND4_in[1] ), .A3(n4433), .A4(
        \SB1_3_23/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_23/buf_output[5] ) );
  NAND4_X2 U7112 ( .A1(\SB2_1_27/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_27/Component_Function_5/NAND4_in[0] ), .A3(
        \SB2_1_27/Component_Function_5/NAND4_in[1] ), .A4(n3620), .ZN(
        \SB2_1_27/buf_output[5] ) );
  NAND3_X2 U7113 ( .A1(\SB2_1_27/i0[9] ), .A2(\SB2_1_27/i0[6] ), .A3(
        \SB2_1_27/i0_4 ), .ZN(n3620) );
  NAND4_X2 U7120 ( .A1(\SB2_0_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_11/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_0_11/Component_Function_3/NAND4_in[1] ), .A4(n3623), .ZN(
        \SB2_0_11/buf_output[3] ) );
  NAND4_X2 U7139 ( .A1(\SB1_2_3/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_3/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_3/Component_Function_0/NAND4_in[0] ), .A4(n3625), .ZN(
        \SB1_2_3/buf_output[0] ) );
  NAND3_X1 U7141 ( .A1(\SB1_4_30/i0_0 ), .A2(\SB1_4_30/i1_7 ), .A3(
        \SB1_4_30/i3[0] ), .ZN(\SB1_4_30/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 U7142 ( .I(\SB1_3_23/buf_output[5] ), .Z(\SB2_3_23/i0_3 ) );
  BUF_X4 U7159 ( .I(\SB2_0_5/buf_output[1] ), .Z(\RI5[0][181] ) );
  NAND3_X1 U7162 ( .A1(\SB1_1_29/i0_3 ), .A2(\SB1_1_29/i0[8] ), .A3(
        \SB1_1_29/i1_7 ), .ZN(\SB1_1_29/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U7166 ( .I(\SB2_4_1/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[3] ) );
  NAND4_X2 U7167 ( .A1(\SB1_0_22/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_22/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_22/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_0_22/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_0_22/buf_output[2] ) );
  XOR2_X1 U7171 ( .A1(\MC_ARK_ARC_1_1/temp2[97] ), .A2(
        \MC_ARK_ARC_1_1/temp1[97] ), .Z(\MC_ARK_ARC_1_1/temp5[97] ) );
  INV_X2 U7172 ( .I(\SB1_0_7/buf_output[3] ), .ZN(\SB2_0_5/i0[8] ) );
  NAND4_X2 U7173 ( .A1(\SB1_0_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_7/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_7/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_0_7/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB1_0_7/buf_output[3] ) );
  XOR2_X1 U7177 ( .A1(\MC_ARK_ARC_1_0/temp2[39] ), .A2(n3629), .Z(
        \MC_ARK_ARC_1_0/temp5[39] ) );
  XOR2_X1 U7178 ( .A1(\RI5[0][33] ), .A2(\RI5[0][39] ), .Z(n3629) );
  XOR2_X1 U7187 ( .A1(n3630), .A2(n11), .Z(Ciphertext[19]) );
  XOR2_X1 U7192 ( .A1(\SB2_1_28/buf_output[1] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[7] ), .Z(\MC_ARK_ARC_1_1/temp3[133] ) );
  NAND4_X2 U7202 ( .A1(\SB3_5/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_5/Component_Function_0/NAND4_in[0] ), .A4(n3632), .ZN(
        \SB3_5/buf_output[0] ) );
  XOR2_X1 U7204 ( .A1(n3862), .A2(n3633), .Z(\RI1[1][11] ) );
  XOR2_X1 U7207 ( .A1(n4015), .A2(\MC_ARK_ARC_1_0/temp4[11] ), .Z(n3633) );
  XOR2_X1 U7210 ( .A1(\MC_ARK_ARC_1_3/temp5[53] ), .A2(n3634), .Z(\RI1[4][53] ) );
  XOR2_X1 U7211 ( .A1(\MC_ARK_ARC_1_3/temp3[53] ), .A2(
        \MC_ARK_ARC_1_3/temp4[53] ), .Z(n3634) );
  XOR2_X1 U7214 ( .A1(n4060), .A2(n3635), .Z(\MC_ARK_ARC_1_3/buf_output[154] )
         );
  XOR2_X1 U7215 ( .A1(n2088), .A2(\MC_ARK_ARC_1_3/temp2[154] ), .Z(n3635) );
  XOR2_X1 U7227 ( .A1(\MC_ARK_ARC_1_0/temp6[67] ), .A2(n3636), .Z(
        \MC_ARK_ARC_1_0/buf_output[67] ) );
  XOR2_X1 U7228 ( .A1(\MC_ARK_ARC_1_0/temp2[67] ), .A2(
        \MC_ARK_ARC_1_0/temp1[67] ), .Z(n3636) );
  NAND3_X2 U7245 ( .A1(\SB1_3_15/i0[10] ), .A2(\SB1_3_15/i0_0 ), .A3(
        \SB1_3_15/i0[6] ), .ZN(n3637) );
  NAND3_X2 U7246 ( .A1(\SB1_2_24/i0_4 ), .A2(\SB1_2_24/i0_3 ), .A3(
        \SB1_2_24/i1[9] ), .ZN(n4819) );
  XOR2_X1 U7249 ( .A1(\RI5[2][67] ), .A2(\RI5[2][103] ), .Z(
        \MC_ARK_ARC_1_2/temp3[1] ) );
  XOR2_X1 U7252 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[140] ), .Z(n5090) );
  XOR2_X1 U7266 ( .A1(\RI5[2][88] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[22] ) );
  NAND4_X2 U7267 ( .A1(\SB2_2_3/Component_Function_2/NAND4_in[2] ), .A2(n4135), 
        .A3(\SB2_2_3/Component_Function_2/NAND4_in[1] ), .A4(n687), .ZN(
        \SB2_2_3/buf_output[2] ) );
  NAND3_X1 U7269 ( .A1(\SB2_1_8/i0_0 ), .A2(\SB2_1_8/i0[9] ), .A3(
        \SB2_1_8/i0[8] ), .ZN(\SB2_1_8/Component_Function_4/NAND4_in[0] ) );
  INV_X1 U7284 ( .I(\SB1_2_8/buf_output[0] ), .ZN(\SB2_2_3/i3[0] ) );
  XOR2_X1 U7289 ( .A1(n3640), .A2(n3639), .Z(\MC_ARK_ARC_1_3/buf_output[182] )
         );
  XOR2_X1 U7294 ( .A1(\SB2_2_25/buf_output[3] ), .A2(\RI5[2][15] ), .Z(
        \MC_ARK_ARC_1_2/temp3[141] ) );
  NAND3_X1 U7296 ( .A1(\SB1_1_26/i0[8] ), .A2(\SB1_1_26/i1_7 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[34] ), .ZN(n3642) );
  XOR2_X1 U7299 ( .A1(\MC_ARK_ARC_1_0/temp1[55] ), .A2(n3643), .Z(
        \MC_ARK_ARC_1_0/temp5[55] ) );
  XOR2_X1 U7300 ( .A1(\RI5[0][1] ), .A2(\RI5[0][25] ), .Z(n3643) );
  INV_X2 U7304 ( .I(\MC_ARK_ARC_1_0/buf_output[55] ), .ZN(\SB1_1_22/i1_7 ) );
  NAND4_X2 U7306 ( .A1(\SB1_1_23/Component_Function_5/NAND4_in[2] ), .A2(n3798), .A3(n3680), .A4(n3645), .ZN(\SB1_1_23/buf_output[5] ) );
  INV_X2 U7307 ( .I(\SB1_1_11/buf_output[2] ), .ZN(\SB2_1_8/i1[9] ) );
  NAND4_X2 U7312 ( .A1(\SB2_1_12/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_12/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_12/Component_Function_0/NAND4_in[0] ), .A4(n3646), .ZN(
        \SB2_1_12/buf_output[0] ) );
  NAND4_X2 U7316 ( .A1(\SB2_0_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_2/Component_Function_2/NAND4_in[2] ), .A4(n3647), .ZN(
        \SB2_0_2/buf_output[2] ) );
  NAND3_X1 U7322 ( .A1(\SB4_5/i0_3 ), .A2(\SB4_5/i1[9] ), .A3(\SB4_5/i0[6] ), 
        .ZN(n3649) );
  INV_X2 U7329 ( .I(\SB1_4_25/buf_output[3] ), .ZN(\SB2_4_23/i0[8] ) );
  XOR2_X1 U7332 ( .A1(\RI5[0][158] ), .A2(\RI5[0][2] ), .Z(n1305) );
  XOR2_X1 U7353 ( .A1(\RI5[4][68] ), .A2(\RI5[4][92] ), .Z(n3651) );
  NAND3_X1 U7358 ( .A1(\SB4_9/i0[6] ), .A2(\SB4_9/i0[9] ), .A3(n6272), .ZN(
        \SB4_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U7362 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0_4 ), .A3(
        \SB2_2_4/i1[9] ), .ZN(\SB2_2_4/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7367 ( .A1(\MC_ARK_ARC_1_2/temp6[180] ), .A2(n3654), .Z(
        \MC_ARK_ARC_1_2/buf_output[180] ) );
  XOR2_X1 U7368 ( .A1(\MC_ARK_ARC_1_2/temp2[180] ), .A2(
        \MC_ARK_ARC_1_2/temp1[180] ), .Z(n3654) );
  NAND3_X2 U7374 ( .A1(\SB1_3_19/i0_3 ), .A2(\SB1_3_19/i0[9] ), .A3(
        \SB1_3_19/i0[8] ), .ZN(n5106) );
  NAND3_X2 U7387 ( .A1(\SB2_2_28/i0[6] ), .A2(\SB2_2_28/i0_4 ), .A3(
        \SB2_2_28/i0[9] ), .ZN(n5043) );
  BUF_X4 U7402 ( .I(\SB1_3_1/buf_output[5] ), .Z(\SB2_3_1/i0_3 ) );
  NAND4_X2 U7403 ( .A1(\SB1_4_4/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_4_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_4/Component_Function_0/NAND4_in[0] ), .A4(n3661), .ZN(
        \SB1_4_4/buf_output[0] ) );
  NAND3_X2 U7410 ( .A1(\SB2_3_20/i0[10] ), .A2(n5440), .A3(\SB2_3_20/i1[9] ), 
        .ZN(\SB2_3_20/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U7414 ( .A1(\RI5[0][159] ), .A2(\RI5[0][3] ), .Z(
        \MC_ARK_ARC_1_0/temp3[93] ) );
  NAND3_X2 U7433 ( .A1(\SB2_3_14/i0_3 ), .A2(\SB2_3_14/i0[10] ), .A3(
        \SB2_3_14/i0[6] ), .ZN(n1716) );
  XOR2_X1 U7434 ( .A1(n3666), .A2(n2168), .Z(\MC_ARK_ARC_1_2/buf_output[60] )
         );
  XOR2_X1 U7435 ( .A1(n893), .A2(\MC_ARK_ARC_1_2/temp2[60] ), .Z(n3666) );
  NAND3_X2 U7439 ( .A1(\SB1_2_27/i0[9] ), .A2(\SB1_2_27/i0_3 ), .A3(
        \SB1_2_27/i0[10] ), .ZN(n3668) );
  NAND3_X1 U7445 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0[8] ), .A3(
        \SB2_1_24/i1_7 ), .ZN(\SB2_1_24/Component_Function_1/NAND4_in[1] ) );
  INV_X2 U7446 ( .I(\SB1_3_1/buf_output[5] ), .ZN(\SB2_3_1/i1_5 ) );
  XOR2_X1 U7462 ( .A1(n3676), .A2(\MC_ARK_ARC_1_2/temp4[26] ), .Z(n3844) );
  XOR2_X1 U7465 ( .A1(\RI5[2][20] ), .A2(\RI5[2][26] ), .Z(n3676) );
  INV_X2 U7475 ( .I(\SB1_3_23/buf_output[3] ), .ZN(\SB2_3_21/i0[8] ) );
  NAND3_X2 U7488 ( .A1(\SB2_4_19/i0_4 ), .A2(\SB2_4_19/i0[6] ), .A3(
        \SB2_4_19/i0[9] ), .ZN(n3678) );
  NAND3_X2 U7493 ( .A1(\RI3[3][70] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \SB2_3_20/i1[9] ), .ZN(\SB2_3_20/Component_Function_5/NAND4_in[2] ) );
  NAND2_X2 U7494 ( .A1(\SB1_1_23/i0_0 ), .A2(\SB1_1_23/i3[0] ), .ZN(n3680) );
  NAND3_X2 U7502 ( .A1(\SB2_4_18/i0_4 ), .A2(\SB2_4_18/i0[6] ), .A3(
        \SB2_4_18/i0[9] ), .ZN(n3681) );
  NAND3_X2 U7518 ( .A1(\SB1_1_17/i0[9] ), .A2(\SB1_1_17/i0[8] ), .A3(
        \SB1_1_17/i0_0 ), .ZN(\SB1_1_17/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U7525 ( .A1(\MC_ARK_ARC_1_0/temp2[190] ), .A2(
        \MC_ARK_ARC_1_0/temp1[190] ), .Z(\MC_ARK_ARC_1_0/temp5[190] ) );
  NAND3_X2 U7539 ( .A1(\SB2_1_28/i0[6] ), .A2(\SB2_1_28/i0[9] ), .A3(n5855), 
        .ZN(n3684) );
  XOR2_X1 U7540 ( .A1(\RI5[4][65] ), .A2(\RI5[4][29] ), .Z(
        \MC_ARK_ARC_1_4/temp3[155] ) );
  NAND3_X2 U7550 ( .A1(\SB2_0_6/i0_3 ), .A2(\SB2_0_6/i0_4 ), .A3(
        \SB2_0_6/i1[9] ), .ZN(\SB2_0_6/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U7560 ( .A1(\SB1_0_26/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_26/Component_Function_1/NAND4_in[0] ), .A4(n3685), .ZN(
        \SB1_0_26/buf_output[1] ) );
  NAND3_X1 U7561 ( .A1(\SB1_0_26/i0[6] ), .A2(\SB1_0_26/i1_5 ), .A3(
        \SB1_0_26/i0[9] ), .ZN(n3685) );
  NAND3_X2 U7581 ( .A1(\SB1_4_12/i0[9] ), .A2(\SB1_4_12/i0[8] ), .A3(
        \SB1_4_12/i0_0 ), .ZN(n3730) );
  NAND3_X2 U7590 ( .A1(\SB1_3_29/i1_5 ), .A2(\SB1_3_29/i0[8] ), .A3(
        \SB1_3_29/i3[0] ), .ZN(n3756) );
  XOR2_X1 U7591 ( .A1(\RI5[1][42] ), .A2(\RI5[1][66] ), .Z(
        \MC_ARK_ARC_1_1/temp2[96] ) );
  NAND3_X2 U7592 ( .A1(\SB2_3_16/i0[6] ), .A2(\SB2_3_16/i0_4 ), .A3(
        \SB2_3_16/i0[9] ), .ZN(n4137) );
  NAND3_X2 U7595 ( .A1(\SB1_0_4/i0_0 ), .A2(\SB1_0_4/i0_4 ), .A3(
        \SB1_0_4/i1_5 ), .ZN(n3690) );
  XOR2_X1 U7600 ( .A1(\MC_ARK_ARC_1_0/temp5[74] ), .A2(n3691), .Z(
        \MC_ARK_ARC_1_0/buf_output[74] ) );
  XOR2_X1 U7604 ( .A1(\RI5[2][42] ), .A2(\RI5[2][66] ), .Z(
        \MC_ARK_ARC_1_2/temp2[96] ) );
  BUF_X4 U7605 ( .I(\MC_ARK_ARC_1_1/buf_output[95] ), .Z(\SB1_2_16/i0_3 ) );
  NAND3_X2 U7608 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i1[9] ), .A3(
        \SB2_2_16/i0[6] ), .ZN(\SB2_2_16/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U7609 ( .A1(\RI5[4][44] ), .A2(\RI5[4][80] ), .Z(
        \MC_ARK_ARC_1_4/temp3[170] ) );
  XOR2_X1 U7613 ( .A1(\MC_ARK_ARC_1_2/temp4[163] ), .A2(
        \MC_ARK_ARC_1_2/temp3[163] ), .Z(n3737) );
  INV_X2 U7616 ( .I(\SB1_2_31/buf_output[3] ), .ZN(\SB2_2_29/i0[8] ) );
  NAND4_X2 U7617 ( .A1(\SB1_0_31/Component_Function_5/NAND4_in[2] ), .A2(n1614), .A3(\SB1_0_31/Component_Function_5/NAND4_in[0] ), .A4(n1450), .ZN(
        \RI3[0][5] ) );
  NAND4_X2 U7654 ( .A1(\SB1_4_25/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_4_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_25/Component_Function_1/NAND4_in[3] ), .A4(n3698), .ZN(
        \SB1_4_25/buf_output[1] ) );
  NAND4_X2 U7662 ( .A1(\SB1_3_23/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_23/Component_Function_0/NAND4_in[0] ), .A4(n3699), .ZN(
        \SB1_3_23/buf_output[0] ) );
  NAND4_X2 U7664 ( .A1(n3700), .A2(\SB2_3_29/Component_Function_5/NAND4_in[2] ), .A3(\SB2_3_29/Component_Function_5/NAND4_in[0] ), .A4(n2407), .ZN(
        \SB2_3_29/buf_output[5] ) );
  NAND4_X2 U7668 ( .A1(\SB3_18/Component_Function_2/NAND4_in[3] ), .A2(
        \SB3_18/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_18/Component_Function_2/NAND4_in[2] ), .A4(n4626), .ZN(
        \SB3_18/buf_output[2] ) );
  XOR2_X1 U7671 ( .A1(\RI5[4][32] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[176] ), 
        .Z(n3701) );
  XOR2_X1 U7684 ( .A1(\RI5[3][86] ), .A2(n517), .Z(n3703) );
  XOR2_X1 U7687 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[20] ), .A2(\RI5[3][50] ), 
        .Z(n3704) );
  NAND3_X2 U7693 ( .A1(\SB1_1_21/i0[10] ), .A2(\SB1_1_21/i1_5 ), .A3(
        \SB1_1_21/i1[9] ), .ZN(\SB1_1_21/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U7694 ( .A1(\RI5[3][92] ), .A2(\RI5[3][56] ), .Z(
        \MC_ARK_ARC_1_3/temp3[182] ) );
  BUF_X4 U7699 ( .I(\SB1_2_29/buf_output[5] ), .Z(\SB2_2_29/i0_3 ) );
  XOR2_X1 U7701 ( .A1(n3708), .A2(n3707), .Z(n4719) );
  XOR2_X1 U7703 ( .A1(n5033), .A2(n3175), .Z(n3707) );
  NAND4_X2 U7707 ( .A1(\SB3_27/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_27/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_27/Component_Function_3/NAND4_in[3] ), .A4(n3710), .ZN(
        \SB3_27/buf_output[3] ) );
  NAND3_X2 U7708 ( .A1(\SB3_27/i0_4 ), .A2(\SB3_27/i0_3 ), .A3(\SB3_27/i0_0 ), 
        .ZN(n3710) );
  INV_X2 U7710 ( .I(\SB1_2_29/buf_output[5] ), .ZN(\SB2_2_29/i1_5 ) );
  NAND4_X2 U7720 ( .A1(\SB1_3_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_22/Component_Function_3/NAND4_in[2] ), .A3(n2310), .A4(n3711), 
        .ZN(\SB1_3_22/buf_output[3] ) );
  NAND3_X2 U7722 ( .A1(\SB1_3_22/i0[8] ), .A2(\SB1_3_22/i3[0] ), .A3(
        \SB1_3_22/i1_5 ), .ZN(n3711) );
  NAND3_X1 U7724 ( .A1(\SB1_1_31/i0[8] ), .A2(\SB1_1_31/i1_7 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[4] ), .ZN(n3712) );
  INV_X2 U7729 ( .I(\SB1_0_22/buf_output[3] ), .ZN(\SB2_0_20/i0[8] ) );
  NAND4_X2 U7730 ( .A1(\SB1_0_22/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_22/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_22/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_0_22/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_0_22/buf_output[3] ) );
  NAND4_X2 U7748 ( .A1(\SB2_3_9/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_9/Component_Function_0/NAND4_in[0] ), .A4(n3714), .ZN(
        \SB2_3_9/buf_output[0] ) );
  NAND3_X1 U7751 ( .A1(\SB4_25/i0[10] ), .A2(\SB4_25/i1[9] ), .A3(
        \SB4_25/i1_5 ), .ZN(n3716) );
  NAND4_X2 U7769 ( .A1(\SB1_3_30/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_30/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_3_30/Component_Function_5/NAND4_in[0] ), .A4(n3718), .ZN(
        \SB1_3_30/buf_output[5] ) );
  NAND3_X2 U7770 ( .A1(\SB1_3_30/i0[6] ), .A2(\SB1_3_30/i0_4 ), .A3(
        \SB1_3_30/i0[9] ), .ZN(n3718) );
  NAND3_X2 U7787 ( .A1(\SB2_1_9/i0[10] ), .A2(\SB2_1_9/i1[9] ), .A3(
        \SB2_1_9/i1_7 ), .ZN(\SB2_1_9/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U7789 ( .A1(\SB2_2_12/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_12/Component_Function_2/NAND4_in[0] ), .A4(n1266), .ZN(
        \SB2_2_12/buf_output[2] ) );
  XOR2_X1 U7791 ( .A1(\RI5[2][17] ), .A2(\RI5[2][173] ), .Z(
        \MC_ARK_ARC_1_2/temp3[107] ) );
  NAND3_X1 U7792 ( .A1(\SB2_4_9/i0_3 ), .A2(\SB2_4_9/i0[8] ), .A3(
        \SB2_4_9/i1_7 ), .ZN(\SB2_4_9/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U7793 ( .I(\MC_ARK_ARC_1_3/buf_output[179] ), .Z(\SB1_4_2/i0_3 ) );
  NAND4_X2 U7798 ( .A1(\SB1_4_8/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_4_8/Component_Function_5/NAND4_in[3] ), .A3(n2927), .A4(n1615), 
        .ZN(\SB1_4_8/buf_output[5] ) );
  NAND4_X2 U7809 ( .A1(\SB4_5/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_5/Component_Function_0/NAND4_in[3] ), .A4(
        \SB4_5/Component_Function_0/NAND4_in[0] ), .ZN(n3960) );
  NAND4_X2 U7817 ( .A1(\SB2_1_17/Component_Function_5/NAND4_in[2] ), .A2(n5418), .A3(n5178), .A4(\SB2_1_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_17/buf_output[5] ) );
  XOR2_X1 U7831 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[83] ), .A2(\RI5[1][89] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[89] ) );
  NAND4_X2 U7833 ( .A1(\SB1_0_21/Component_Function_4/NAND4_in[1] ), .A2(n1233), .A3(\SB1_0_21/Component_Function_4/NAND4_in[3] ), .A4(n3722), .ZN(
        \SB1_0_21/buf_output[4] ) );
  NAND3_X2 U7837 ( .A1(\SB1_0_21/i0_0 ), .A2(\SB1_0_21/i0[9] ), .A3(
        \SB1_0_21/i0[8] ), .ZN(n3722) );
  NAND3_X1 U7839 ( .A1(\SB1_4_20/i0[9] ), .A2(\SB1_4_20/i0_3 ), .A3(
        \SB1_4_20/i0[8] ), .ZN(\SB1_4_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U7842 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i0_3 ), .A3(
        \SB1_3_17/i1[9] ), .ZN(n1593) );
  NAND3_X1 U7847 ( .A1(\SB2_3_1/i0_0 ), .A2(\SB2_3_1/i0_3 ), .A3(
        \SB2_3_1/i0[7] ), .ZN(n3725) );
  NAND3_X2 U7850 ( .A1(\SB2_2_20/i3[0] ), .A2(\SB2_2_20/i1_5 ), .A3(
        \SB2_2_20/i0[8] ), .ZN(n4104) );
  NAND3_X1 U7854 ( .A1(\SB2_4_29/i0_0 ), .A2(\SB2_4_29/i3[0] ), .A3(
        \SB2_4_29/i1_7 ), .ZN(n3726) );
  XOR2_X1 U7869 ( .A1(\RI5[3][165] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[159] ), 
        .Z(n3728) );
  NAND4_X2 U7872 ( .A1(\SB1_3_9/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_3_9/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_3_9/Component_Function_4/NAND4_in[1] ), .A4(n3729), .ZN(
        \SB1_3_9/buf_output[4] ) );
  NAND3_X1 U7873 ( .A1(\SB1_3_9/i0[10] ), .A2(\SB1_3_9/i0_3 ), .A3(n3979), 
        .ZN(n3729) );
  NAND4_X2 U7883 ( .A1(\SB1_4_4/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_4_4/Component_Function_3/NAND4_in[0] ), .A3(n4962), .A4(n3733), 
        .ZN(\SB1_4_4/buf_output[3] ) );
  NAND3_X1 U7884 ( .A1(\SB1_1_27/i0_4 ), .A2(\SB1_1_27/i1[9] ), .A3(
        \SB1_1_27/i1_5 ), .ZN(n3734) );
  XOR2_X1 U7888 ( .A1(\RI5[0][161] ), .A2(\RI5[0][167] ), .Z(n3735) );
  XOR2_X1 U7889 ( .A1(n3079), .A2(\MC_ARK_ARC_1_4/temp4[20] ), .Z(n3736) );
  NAND4_X2 U7897 ( .A1(\SB2_2_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_2/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_2_2/Component_Function_1/NAND4_in[2] ), .A4(n3738), .ZN(
        \SB2_2_2/buf_output[1] ) );
  NAND4_X2 U7901 ( .A1(\SB3_3/Component_Function_3/NAND4_in[1] ), .A2(n4645), 
        .A3(\SB3_3/Component_Function_3/NAND4_in[0] ), .A4(
        \SB3_3/Component_Function_3/NAND4_in[3] ), .ZN(\SB3_3/buf_output[3] )
         );
  XOR2_X1 U7905 ( .A1(n869), .A2(n3740), .Z(\MC_ARK_ARC_1_0/buf_output[138] )
         );
  XOR2_X1 U7907 ( .A1(\MC_ARK_ARC_1_0/temp4[138] ), .A2(
        \MC_ARK_ARC_1_0/temp3[138] ), .Z(n3740) );
  XOR2_X1 U7910 ( .A1(\MC_ARK_ARC_1_0/temp4[43] ), .A2(n3742), .Z(
        \MC_ARK_ARC_1_0/temp6[43] ) );
  XOR2_X1 U7912 ( .A1(\RI5[0][145] ), .A2(\RI5[0][109] ), .Z(n3742) );
  NAND3_X2 U7925 ( .A1(\SB2_3_0/i0_4 ), .A2(\SB2_3_0/i0_3 ), .A3(
        \SB2_3_0/i1[9] ), .ZN(n3743) );
  NAND3_X2 U7926 ( .A1(\SB2_0_18/i0[8] ), .A2(\SB2_0_18/i1_5 ), .A3(
        \SB2_0_18/i3[0] ), .ZN(\SB2_0_18/Component_Function_3/NAND4_in[3] ) );
  INV_X2 U7927 ( .I(\SB1_4_12/buf_output[3] ), .ZN(\SB2_4_10/i0[8] ) );
  NAND4_X2 U7931 ( .A1(\SB2_1_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_4/NAND4_in[3] ), .A3(n3745), .A4(n3744), 
        .ZN(\SB2_1_12/buf_output[4] ) );
  NAND3_X1 U7932 ( .A1(\SB2_1_12/i0_0 ), .A2(\SB2_1_12/i3[0] ), .A3(
        \SB2_1_12/i1_7 ), .ZN(n3745) );
  NAND3_X1 U7933 ( .A1(\SB4_19/i0[10] ), .A2(\SB4_19/i1[9] ), .A3(
        \SB4_19/i1_7 ), .ZN(n3746) );
  XOR2_X1 U7934 ( .A1(\SB2_2_14/buf_output[0] ), .A2(\RI5[2][156] ), .Z(
        \MC_ARK_ARC_1_2/temp2[186] ) );
  BUF_X4 U7940 ( .I(n4006), .Z(\SB3_5/i0_3 ) );
  NAND3_X2 U7946 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0[9] ), .A3(
        \SB3_30/i0[10] ), .ZN(n3749) );
  XOR2_X1 U7947 ( .A1(n3750), .A2(n61), .Z(Ciphertext[16]) );
  XOR2_X1 U7952 ( .A1(\MC_ARK_ARC_1_4/temp5[61] ), .A2(n3752), .Z(
        \MC_ARK_ARC_1_4/buf_output[61] ) );
  XOR2_X1 U7955 ( .A1(\MC_ARK_ARC_1_4/temp3[61] ), .A2(
        \MC_ARK_ARC_1_4/temp4[61] ), .Z(n3752) );
  NAND4_X2 U7956 ( .A1(\SB2_3_2/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_3_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_2/Component_Function_3/NAND4_in[0] ), .A4(n3753), .ZN(
        \SB2_3_2/buf_output[3] ) );
  NAND3_X2 U7963 ( .A1(\SB2_3_2/i3[0] ), .A2(\SB2_3_2/i1_5 ), .A3(
        \SB2_3_2/i0[8] ), .ZN(n3753) );
  NAND3_X1 U7966 ( .A1(\SB2_4_20/i0[7] ), .A2(\SB2_4_20/i0[8] ), .A3(
        \SB2_4_20/i0[6] ), .ZN(\SB2_4_20/Component_Function_0/NAND4_in[1] ) );
  BUF_X2 U7984 ( .I(\RI1[3][17] ), .Z(n3757) );
  INV_X2 U7989 ( .I(\SB1_4_4/buf_output[3] ), .ZN(\SB2_4_2/i0[8] ) );
  BUF_X4 U8025 ( .I(\SB2_4_17/buf_output[3] ), .Z(\RI5[4][99] ) );
  XOR2_X1 U8027 ( .A1(\RI5[0][59] ), .A2(\RI5[0][65] ), .Z(n3762) );
  NAND3_X2 U8044 ( .A1(\SB2_2_7/i0_4 ), .A2(\SB2_2_7/i0_3 ), .A3(
        \SB2_2_7/i1[9] ), .ZN(n3766) );
  NAND3_X1 U8050 ( .A1(\SB1_0_24/i0_3 ), .A2(n332), .A3(\SB1_0_24/i1[9] ), 
        .ZN(\SB1_0_24/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U8054 ( .A1(\SB2_0_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_21/Component_Function_4/NAND4_in[3] ), .A4(n4781), .ZN(
        \SB2_0_21/buf_output[4] ) );
  XOR2_X1 U8056 ( .A1(\MC_ARK_ARC_1_3/temp6[76] ), .A2(
        \MC_ARK_ARC_1_3/temp5[76] ), .Z(\MC_ARK_ARC_1_3/buf_output[76] ) );
  NAND3_X1 U8059 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i1[9] ), .A3(
        \SB1_1_19/i0[6] ), .ZN(\SB1_1_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U8062 ( .A1(\SB1_2_31/i0_4 ), .A2(\SB1_2_31/i0_3 ), .A3(
        \SB1_2_31/i1[9] ), .ZN(n3091) );
  NAND3_X1 U8065 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i0[8] ), .A3(
        \SB1_1_14/i1_7 ), .ZN(\SB1_1_14/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U8069 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[15] ), .A2(\RI5[1][9] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[15] ) );
  XOR2_X1 U8070 ( .A1(\MC_ARK_ARC_1_1/temp5[4] ), .A2(
        \MC_ARK_ARC_1_1/temp6[4] ), .Z(\MC_ARK_ARC_1_1/buf_output[4] ) );
  XOR2_X1 U8072 ( .A1(\MC_ARK_ARC_1_1/temp5[13] ), .A2(
        \MC_ARK_ARC_1_1/temp6[13] ), .Z(\MC_ARK_ARC_1_1/buf_output[13] ) );
  XOR2_X1 U8073 ( .A1(\RI5[2][78] ), .A2(\RI5[2][102] ), .Z(
        \MC_ARK_ARC_1_2/temp2[132] ) );
  XOR2_X1 U8074 ( .A1(n4800), .A2(n4017), .Z(n4005) );
  INV_X1 U8079 ( .I(\SB1_4_2/buf_output[1] ), .ZN(\SB2_4_30/i1_7 ) );
  NAND4_X2 U8080 ( .A1(\SB1_4_2/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_4_2/Component_Function_1/NAND4_in[1] ), .A3(n5040), .A4(
        \SB1_4_2/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_4_2/buf_output[1] ) );
  NAND3_X1 U8087 ( .A1(\SB4_30/i0[6] ), .A2(\SB4_30/i0_3 ), .A3(n3973), .ZN(
        n3769) );
  NAND3_X1 U8103 ( .A1(\SB2_1_30/i0[10] ), .A2(\SB2_1_30/i0_3 ), .A3(
        \SB2_1_30/i0_4 ), .ZN(\SB2_1_30/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U8104 ( .A1(\SB1_0_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_27/Component_Function_2/NAND4_in[3] ), .A4(n3773), .ZN(
        \RI3[0][44] ) );
  XOR2_X1 U8113 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[122] ), .A2(n537), .Z(
        n3774) );
  XOR2_X1 U8114 ( .A1(\RI5[2][86] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .Z(n3775) );
  XOR2_X1 U8116 ( .A1(\MC_ARK_ARC_1_3/temp2[167] ), .A2(
        \MC_ARK_ARC_1_3/temp4[167] ), .Z(n3776) );
  XOR2_X1 U8118 ( .A1(\MC_ARK_ARC_1_3/temp1[167] ), .A2(n1433), .Z(n3777) );
  NAND3_X1 U8126 ( .A1(\SB4_14/i0[10] ), .A2(n1495), .A3(\SB4_14/i1[9] ), .ZN(
        \SB4_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U8138 ( .A1(\SB4_4/i0[10] ), .A2(\SB4_4/i0_3 ), .A3(\SB4_4/i0[6] ), 
        .ZN(n3780) );
  NAND4_X2 U8139 ( .A1(\SB1_0_16/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_16/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_16/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_0_16/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_0_16/buf_output[3] ) );
  XOR2_X1 U8144 ( .A1(\MC_ARK_ARC_1_3/temp6[65] ), .A2(n3781), .Z(\RI1[4][65] ) );
  XOR2_X1 U8147 ( .A1(\MC_ARK_ARC_1_3/temp1[65] ), .A2(
        \MC_ARK_ARC_1_3/temp2[65] ), .Z(n3781) );
  INV_X1 U8149 ( .I(\SB3_6/buf_output[1] ), .ZN(\SB4_2/i1_7 ) );
  NAND4_X2 U8153 ( .A1(\SB3_6/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_6/Component_Function_1/NAND4_in[3] ), .A3(
        \SB3_6/Component_Function_1/NAND4_in[1] ), .A4(
        \SB3_6/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_6/buf_output[1] )
         );
  NAND3_X1 U8168 ( .A1(\SB4_4/i0[10] ), .A2(\SB4_4/i1[9] ), .A3(\SB4_4/i1_7 ), 
        .ZN(n3783) );
  XOR2_X1 U8171 ( .A1(\MC_ARK_ARC_1_1/temp2[154] ), .A2(n3785), .Z(n4555) );
  XOR2_X1 U8173 ( .A1(\RI5[1][148] ), .A2(\RI5[1][154] ), .Z(n3785) );
  NAND3_X2 U8180 ( .A1(\SB2_4_6/i0_3 ), .A2(\SB2_4_6/i0_0 ), .A3(
        \SB2_4_6/i0_4 ), .ZN(n1938) );
  NAND4_X2 U8189 ( .A1(\SB4_8/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_8/Component_Function_1/NAND4_in[0] ), .ZN(n5257) );
  NAND3_X2 U8190 ( .A1(\SB3_18/i0[6] ), .A2(\SB3_18/i0[10] ), .A3(
        \SB3_18/i0_3 ), .ZN(n4626) );
  NAND3_X2 U8193 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i0_4 ), .A3(
        \SB2_0_25/i1[9] ), .ZN(n3787) );
  NAND3_X1 U8217 ( .A1(\SB4_5/i0_4 ), .A2(\SB4_5/i0[9] ), .A3(\SB4_5/i0[6] ), 
        .ZN(n3788) );
  NAND4_X2 U8220 ( .A1(n3109), .A2(\SB1_1_30/Component_Function_2/NAND4_in[0] ), .A3(\SB1_1_30/Component_Function_2/NAND4_in[2] ), .A4(n3789), .ZN(
        \SB1_1_30/buf_output[2] ) );
  NAND3_X2 U8224 ( .A1(\SB1_1_30/i0[6] ), .A2(\SB1_1_30/i0_3 ), .A3(
        \SB1_1_30/i0[10] ), .ZN(n3789) );
  XOR2_X1 U8226 ( .A1(n3790), .A2(n174), .Z(Ciphertext[23]) );
  NAND4_X2 U8233 ( .A1(n3851), .A2(\SB4_28/Component_Function_5/NAND4_in[1] ), 
        .A3(n2453), .A4(\SB4_28/Component_Function_5/NAND4_in[0] ), .ZN(n3790)
         );
  NAND3_X1 U8235 ( .A1(\SB1_4_13/i0[9] ), .A2(\SB1_4_13/i1_5 ), .A3(
        \SB1_4_13/i0[6] ), .ZN(\SB1_4_13/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U8241 ( .A1(\SB1_3_24/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_24/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_5/NAND4_in[0] ), .A4(n3792), .ZN(
        \SB1_3_24/buf_output[5] ) );
  NAND3_X1 U8249 ( .A1(\SB1_2_12/i0[9] ), .A2(\RI1[2][116] ), .A3(
        \SB1_2_12/i0[8] ), .ZN(\SB1_2_12/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U8257 ( .A1(\SB2_3_24/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_24/Component_Function_0/NAND4_in[0] ), .A4(n3794), .ZN(
        \SB2_3_24/buf_output[0] ) );
  XOR2_X1 U8269 ( .A1(n3795), .A2(n2767), .Z(\MC_ARK_ARC_1_0/buf_output[132] )
         );
  XOR2_X1 U8271 ( .A1(\MC_ARK_ARC_1_0/temp4[132] ), .A2(n2485), .Z(n3795) );
  XOR2_X1 U8289 ( .A1(\MC_ARK_ARC_1_0/temp2[183] ), .A2(n3797), .Z(n2788) );
  XOR2_X1 U8293 ( .A1(\RI5[0][183] ), .A2(\RI5[0][177] ), .Z(n3797) );
  NAND3_X2 U8302 ( .A1(\SB1_1_23/i0[10] ), .A2(\SB1_1_23/i0_0 ), .A3(
        \SB1_1_23/i0[6] ), .ZN(n3798) );
  NAND4_X2 U8308 ( .A1(\SB3_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_27/Component_Function_1/NAND4_in[3] ), .A3(
        \SB3_27/Component_Function_1/NAND4_in[0] ), .A4(n3799), .ZN(
        \SB3_27/buf_output[1] ) );
  AND2_X1 U8310 ( .A1(n3848), .A2(\SB1_0_10/Component_Function_3/NAND4_in[2] ), 
        .Z(n3802) );
  XOR2_X1 U8312 ( .A1(\RI5[4][109] ), .A2(\RI5[4][145] ), .Z(
        \MC_ARK_ARC_1_4/temp3[43] ) );
  NAND4_X2 U8318 ( .A1(\SB3_24/Component_Function_3/NAND4_in[1] ), .A2(n1398), 
        .A3(n4586), .A4(n3804), .ZN(\SB3_24/buf_output[3] ) );
  XOR2_X1 U8325 ( .A1(n2256), .A2(n3806), .Z(\MC_ARK_ARC_1_4/buf_output[24] )
         );
  XOR2_X1 U8327 ( .A1(\MC_ARK_ARC_1_4/temp1[24] ), .A2(
        \MC_ARK_ARC_1_4/temp2[24] ), .Z(n3806) );
  XOR2_X1 U8334 ( .A1(n4461), .A2(n933), .Z(\MC_ARK_ARC_1_3/buf_output[18] )
         );
  NAND3_X1 U8342 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i0[9] ), .A3(n1494), .ZN(
        n3807) );
  NAND4_X2 U8343 ( .A1(\SB2_4_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_4_1/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_4_1/Component_Function_1/NAND4_in[2] ), .A4(n3808), .ZN(
        \SB2_4_1/buf_output[1] ) );
  NAND4_X2 U8355 ( .A1(\SB2_0_31/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_31/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_31/Component_Function_4/NAND4_in[1] ), .A4(n3811), .ZN(
        \SB2_0_31/buf_output[4] ) );
  NAND3_X1 U8359 ( .A1(\SB2_0_31/i1[9] ), .A2(\RI3[0][4] ), .A3(
        \SB2_0_31/i1_5 ), .ZN(n3811) );
  NAND3_X2 U8362 ( .A1(\SB2_2_10/i0[6] ), .A2(\SB2_2_10/i0[7] ), .A3(
        \SB2_2_10/i0[8] ), .ZN(\SB2_2_10/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U8365 ( .A1(n3814), .A2(n3813), .Z(\MC_ARK_ARC_1_2/temp6[120] ) );
  XOR2_X1 U8366 ( .A1(\SB2_2_31/buf_output[0] ), .A2(n435), .Z(n3813) );
  XOR2_X1 U8367 ( .A1(\RI5[2][186] ), .A2(\RI5[2][156] ), .Z(n3814) );
  XOR2_X1 U8370 ( .A1(n3815), .A2(\MC_ARK_ARC_1_2/temp1[43] ), .Z(
        \MC_ARK_ARC_1_2/temp5[43] ) );
  XOR2_X1 U8371 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[181] ), .A2(\RI5[2][13] ), 
        .Z(n3815) );
  NAND3_X2 U8375 ( .A1(\SB2_1_15/i0[8] ), .A2(\SB2_1_15/i0[7] ), .A3(
        \SB2_1_15/i0[6] ), .ZN(\SB2_1_15/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U8376 ( .A1(\SB2_3_17/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_17/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_17/Component_Function_0/NAND4_in[0] ), .A4(n3817), .ZN(
        \SB2_3_17/buf_output[0] ) );
  NAND4_X2 U8380 ( .A1(\SB2_2_29/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_29/Component_Function_4/NAND4_in[0] ), .A3(n2429), .A4(n3819), 
        .ZN(\SB2_2_29/buf_output[4] ) );
  NAND3_X1 U8382 ( .A1(\SB4_21/i0[6] ), .A2(\SB4_21/i0[7] ), .A3(
        \SB4_21/i0[8] ), .ZN(n3820) );
  NAND3_X1 U8384 ( .A1(\SB4_20/i1_7 ), .A2(\SB4_20/i0[10] ), .A3(
        \SB4_20/i1[9] ), .ZN(\SB4_20/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U8391 ( .A1(\RI5[0][15] ), .A2(\RI5[0][51] ), .Z(n3822) );
  BUF_X4 U8395 ( .I(\SB2_4_13/buf_output[1] ), .Z(\RI5[4][133] ) );
  XOR2_X1 U8399 ( .A1(\MC_ARK_ARC_1_4/temp2[188] ), .A2(n3824), .Z(n2985) );
  XOR2_X1 U8400 ( .A1(\RI5[4][182] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[188] ), 
        .Z(n3824) );
  NAND4_X2 U8424 ( .A1(\SB2_4_4/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_4/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_4_4/Component_Function_0/NAND4_in[0] ), .A4(n3828), .ZN(
        \SB2_4_4/buf_output[0] ) );
  XOR2_X1 U8426 ( .A1(n3829), .A2(\MC_ARK_ARC_1_3/temp1[60] ), .Z(
        \MC_ARK_ARC_1_3/temp5[60] ) );
  XOR2_X1 U8428 ( .A1(\RI5[3][6] ), .A2(\RI5[3][30] ), .Z(n3829) );
  XOR2_X1 U8435 ( .A1(n796), .A2(n3830), .Z(\MC_ARK_ARC_1_4/buf_output[6] ) );
  XOR2_X1 U8440 ( .A1(n3831), .A2(n186), .Z(Ciphertext[96]) );
  NAND4_X2 U8442 ( .A1(\SB4_15/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_15/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_15/Component_Function_0/NAND4_in[3] ), .ZN(n3831) );
  NAND3_X1 U8449 ( .A1(\SB3_20/i0[10] ), .A2(\SB3_20/i1[9] ), .A3(
        \SB3_20/i1_7 ), .ZN(\SB3_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U8451 ( .A1(\SB2_2_5/i0_0 ), .A2(\SB2_2_5/i3[0] ), .A3(
        \SB2_2_5/i1_7 ), .ZN(\SB2_2_5/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U8456 ( .A1(\SB1_1_14/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_14/Component_Function_1/NAND4_in[2] ), .A3(n2081), .A4(n3833), 
        .ZN(\SB1_1_14/buf_output[1] ) );
  XOR2_X1 U8458 ( .A1(\RI5[0][4] ), .A2(\RI5[0][136] ), .Z(n3834) );
  NAND3_X1 U8462 ( .A1(\SB4_15/i0_0 ), .A2(\SB4_15/i0_4 ), .A3(\SB4_15/i1_5 ), 
        .ZN(n3880) );
  XOR2_X1 U8469 ( .A1(n3836), .A2(n4849), .Z(\MC_ARK_ARC_1_0/temp5[30] ) );
  XOR2_X1 U8471 ( .A1(\RI5[0][168] ), .A2(\RI5[0][0] ), .Z(n3836) );
  NAND3_X1 U8476 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i0[8] ), .A3(
        \SB1_1_16/i1_7 ), .ZN(\SB1_1_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U8479 ( .A1(\SB1_0_2/i0_4 ), .A2(\SB1_0_2/i0_0 ), .A3(
        \SB1_0_2/i1_5 ), .ZN(n1839) );
  BUF_X4 U8480 ( .I(\SB2_3_1/buf_output[5] ), .Z(\RI5[3][185] ) );
  NAND4_X2 U8482 ( .A1(\SB2_3_19/Component_Function_3/NAND4_in[0] ), .A2(n871), 
        .A3(n5148), .A4(\SB2_3_19/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_19/buf_output[3] ) );
  XOR2_X1 U8495 ( .A1(\MC_ARK_ARC_1_2/temp1[54] ), .A2(
        \MC_ARK_ARC_1_2/temp2[54] ), .Z(\MC_ARK_ARC_1_2/temp5[54] ) );
  NAND2_X2 U8496 ( .A1(\SB1_2_29/i1_5 ), .A2(n3838), .ZN(n2132) );
  NOR2_X1 U8497 ( .A1(\MC_ARK_ARC_1_1/buf_output[12] ), .A2(
        \MC_ARK_ARC_1_1/buf_output[15] ), .ZN(n3838) );
  NAND4_X2 U8511 ( .A1(\SB2_0_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_1/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_1/Component_Function_3/NAND4_in[2] ), .A4(n3842), .ZN(
        \SB2_0_1/buf_output[3] ) );
  XOR2_X1 U8525 ( .A1(n3843), .A2(\MC_ARK_ARC_1_0/temp4[175] ), .Z(
        \MC_ARK_ARC_1_0/temp6[175] ) );
  XOR2_X1 U8526 ( .A1(\RI5[0][49] ), .A2(\RI5[0][85] ), .Z(n3843) );
  XOR2_X1 U8529 ( .A1(n3844), .A2(n1702), .Z(\MC_ARK_ARC_1_2/buf_output[26] )
         );
  BUF_X4 U8530 ( .I(\SB2_4_31/buf_output[5] ), .Z(\RI5[4][5] ) );
  NAND4_X2 U8539 ( .A1(\SB2_0_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_27/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_0_27/Component_Function_1/NAND4_in[0] ), .A4(n4964), .ZN(
        \SB2_0_27/buf_output[1] ) );
  NAND4_X2 U8546 ( .A1(\SB2_2_7/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_7/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_7/Component_Function_4/NAND4_in[2] ), .A4(n3846), .ZN(
        \SB2_2_7/buf_output[4] ) );
  NAND3_X2 U8549 ( .A1(\SB2_2_7/i0_0 ), .A2(\SB2_2_7/i3[0] ), .A3(
        \SB2_2_7/i1_7 ), .ZN(n3846) );
  NAND4_X2 U8554 ( .A1(\SB1_4_23/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_23/Component_Function_0/NAND4_in[0] ), .A4(n3847), .ZN(
        \SB1_4_23/buf_output[0] ) );
  XOR2_X1 U8562 ( .A1(\RI5[3][190] ), .A2(\RI5[3][4] ), .Z(
        \MC_ARK_ARC_1_3/temp1[4] ) );
  XOR2_X1 U8565 ( .A1(\MC_ARK_ARC_1_0/temp3[54] ), .A2(
        \MC_ARK_ARC_1_0/temp4[54] ), .Z(\MC_ARK_ARC_1_0/temp6[54] ) );
  NAND3_X1 U8569 ( .A1(\SB1_0_10/i0_0 ), .A2(\SB1_0_10/i0_4 ), .A3(
        \SB1_0_10/i0_3 ), .ZN(n3848) );
  NAND3_X1 U8578 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i0_4 ), .A3(\SB4_28/i1[9] ), 
        .ZN(n3851) );
  NAND3_X2 U8581 ( .A1(\SB1_2_19/i0[10] ), .A2(\SB1_2_19/i1[9] ), .A3(
        \SB1_2_19/i1_7 ), .ZN(n3852) );
  XOR2_X1 U8584 ( .A1(\RI5[0][181] ), .A2(\RI5[0][13] ), .Z(
        \MC_ARK_ARC_1_0/temp2[43] ) );
  XOR2_X1 U8590 ( .A1(\MC_ARK_ARC_1_3/temp6[166] ), .A2(n3854), .Z(
        \MC_ARK_ARC_1_3/buf_output[166] ) );
  XOR2_X1 U8596 ( .A1(\MC_ARK_ARC_1_3/temp2[166] ), .A2(
        \MC_ARK_ARC_1_3/temp1[166] ), .Z(n3854) );
  XOR2_X1 U8598 ( .A1(\MC_ARK_ARC_1_2/temp3[93] ), .A2(
        \MC_ARK_ARC_1_2/temp4[93] ), .Z(n3855) );
  NAND4_X2 U8608 ( .A1(\SB1_0_10/Component_Function_4/NAND4_in[2] ), .A2(n5221), .A3(\SB1_0_10/Component_Function_4/NAND4_in[0] ), .A4(n3857), .ZN(
        \RI3[0][136] ) );
  NAND3_X1 U8611 ( .A1(\SB1_0_10/i0_4 ), .A2(\SB1_0_10/i1[9] ), .A3(
        \SB1_0_10/i1_5 ), .ZN(n3857) );
  NAND4_X2 U8612 ( .A1(\SB2_1_3/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_3/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_3/Component_Function_4/NAND4_in[3] ), .A4(n3858), .ZN(
        \SB2_1_3/buf_output[4] ) );
  XOR2_X1 U8618 ( .A1(n2948), .A2(n3860), .Z(\MC_ARK_ARC_1_2/temp5[68] ) );
  XOR2_X1 U8620 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), .A2(\RI5[2][62] ), 
        .Z(n3860) );
  NAND3_X2 U8622 ( .A1(\SB2_2_21/i1[9] ), .A2(\SB1_2_22/buf_output[4] ), .A3(
        \SB2_2_21/i0_3 ), .ZN(\SB2_2_21/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U8627 ( .I(\SB1_2_27/buf_output[2] ), .ZN(\SB2_2_24/i1[9] ) );
  NAND4_X2 U8637 ( .A1(\SB1_4_23/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_4_23/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_4_23/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_4_23/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_4_23/buf_output[4] ) );
  NAND3_X2 U8650 ( .A1(\SB2_1_20/i0[6] ), .A2(\SB2_1_20/i0[9] ), .A3(
        \SB2_1_20/i0_4 ), .ZN(n980) );
  XOR2_X1 U8676 ( .A1(\MC_ARK_ARC_1_3/temp5[60] ), .A2(n3868), .Z(
        \MC_ARK_ARC_1_3/buf_output[60] ) );
  XOR2_X1 U8677 ( .A1(\MC_ARK_ARC_1_3/temp3[60] ), .A2(
        \MC_ARK_ARC_1_3/temp4[60] ), .Z(n3868) );
  BUF_X4 U8686 ( .I(\SB1_3_15/buf_output[5] ), .Z(\SB2_3_15/i0_3 ) );
  NAND3_X2 U8699 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i0[8] ), .A3(\SB3_1/i0[9] ), 
        .ZN(\SB3_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U8702 ( .A1(n6290), .A2(\SB1_0_18/i0[9] ), .A3(\SB1_0_18/i0[8] ), 
        .ZN(n3870) );
  XOR2_X1 U8703 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[97] ), .A2(\RI5[0][91] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[97] ) );
  XOR2_X1 U8718 ( .A1(n3872), .A2(\MC_ARK_ARC_1_2/temp1[189] ), .Z(
        \MC_ARK_ARC_1_2/temp5[189] ) );
  INV_X2 U8730 ( .I(\SB1_3_0/buf_output[3] ), .ZN(\SB2_3_30/i0[8] ) );
  XOR2_X1 U8745 ( .A1(\RI5[4][42] ), .A2(\RI5[4][48] ), .Z(n3874) );
  NAND4_X2 U8750 ( .A1(\SB2_2_11/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_2_11/Component_Function_3/NAND4_in[2] ), .A3(n5166), .A4(n3875), 
        .ZN(\SB2_2_11/buf_output[3] ) );
  INV_X2 U8753 ( .I(\SB1_1_6/buf_output[2] ), .ZN(\SB2_1_3/i1[9] ) );
  NAND3_X1 U8759 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i0[10] ), .A3(
        \SB1_0_16/i0[9] ), .ZN(n3877) );
  XOR2_X1 U8760 ( .A1(\MC_ARK_ARC_1_1/temp5[73] ), .A2(n3878), .Z(
        \MC_ARK_ARC_1_1/buf_output[73] ) );
  NAND4_X2 U8762 ( .A1(\SB1_3_5/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_3_5/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_5/Component_Function_3/NAND4_in[1] ), .A4(n3879), .ZN(
        \SB1_3_5/buf_output[3] ) );
  NAND3_X2 U8768 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[6] ), .A3(
        \SB1_3_31/i1[9] ), .ZN(\SB1_3_31/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U8771 ( .A1(\SB1_0_24/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_0_24/Component_Function_0/NAND4_in[3] ), .A3(n4138), .A4(
        \SB1_0_24/Component_Function_0/NAND4_in[2] ), .ZN(\RI3[0][72] ) );
  NAND3_X1 U8774 ( .A1(\SB4_4/i0_0 ), .A2(\SB4_4/i0[9] ), .A3(\SB4_4/i0[8] ), 
        .ZN(n3882) );
  BUF_X4 U8775 ( .I(\MC_ARK_ARC_1_0/buf_output[167] ), .Z(\SB1_1_4/i0_3 ) );
  NAND3_X2 U8787 ( .A1(\SB2_1_12/i0_0 ), .A2(\SB2_1_12/i0[10] ), .A3(
        \SB2_1_12/i0[6] ), .ZN(n3883) );
  XOR2_X1 U8791 ( .A1(n3886), .A2(n3885), .Z(\MC_ARK_ARC_1_1/buf_output[57] )
         );
  XOR2_X1 U8792 ( .A1(\MC_ARK_ARC_1_1/temp2[57] ), .A2(
        \MC_ARK_ARC_1_1/temp4[57] ), .Z(n3885) );
  BUF_X4 U8793 ( .I(\SB2_1_23/buf_output[2] ), .Z(\RI5[1][68] ) );
  INV_X2 U8794 ( .I(\SB1_3_4/buf_output[2] ), .ZN(\SB2_3_1/i1[9] ) );
  NAND3_X2 U8812 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i0[10] ), .A3(
        \SB1_0_11/i0[6] ), .ZN(n3891) );
  INV_X1 U8813 ( .I(\SB1_1_6/buf_output[1] ), .ZN(\SB2_1_2/i1_7 ) );
  NAND4_X2 U8816 ( .A1(\SB1_1_6/Component_Function_1/NAND4_in[1] ), .A2(n1918), 
        .A3(\SB1_1_6/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_1_6/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_1_6/buf_output[1] ) );
  XOR2_X1 U8818 ( .A1(n3892), .A2(\MC_ARK_ARC_1_1/temp2[9] ), .Z(
        \MC_ARK_ARC_1_1/temp5[9] ) );
  XOR2_X1 U8820 ( .A1(\RI5[1][9] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[3] ), 
        .Z(n3892) );
  NAND3_X1 U8849 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i0_0 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[94] ), .ZN(
        \SB1_1_16/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U8855 ( .A1(\SB1_1_25/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_1_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_25/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_1_25/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_25/buf_output[4] ) );
  XOR2_X1 U8859 ( .A1(n4357), .A2(\MC_ARK_ARC_1_1/temp6[32] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[32] ) );
  NAND3_X2 U8863 ( .A1(\SB2_4_16/i0_3 ), .A2(\SB2_4_16/i0_4 ), .A3(
        \SB2_4_16/i1[9] ), .ZN(n3102) );
  NAND3_X1 U8865 ( .A1(\SB2_2_23/i0[6] ), .A2(\SB2_2_23/i0[7] ), .A3(
        \SB2_2_23/i0[8] ), .ZN(\SB2_2_23/Component_Function_0/NAND4_in[1] ) );
  BUF_X4 U8872 ( .I(\SB1_0_5/buf_output[5] ), .Z(\SB2_0_5/i0_3 ) );
  XOR2_X1 U8873 ( .A1(\MC_ARK_ARC_1_1/temp3[161] ), .A2(
        \MC_ARK_ARC_1_1/temp4[161] ), .Z(n5412) );
  NAND4_X2 U8892 ( .A1(n602), .A2(\SB2_3_27/Component_Function_5/NAND4_in[1] ), 
        .A3(n4718), .A4(\SB2_3_27/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_27/buf_output[5] ) );
  XOR2_X1 U8893 ( .A1(\RI5[1][134] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[164] ) );
  XOR2_X1 U8894 ( .A1(\RI5[2][187] ), .A2(\RI5[2][1] ), .Z(
        \MC_ARK_ARC_1_2/temp1[1] ) );
  XOR2_X1 U8905 ( .A1(n4030), .A2(n3898), .Z(n4628) );
  XOR2_X1 U8908 ( .A1(\RI5[3][160] ), .A2(\RI5[3][16] ), .Z(n3898) );
  NAND4_X2 U8940 ( .A1(\SB1_3_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_23/Component_Function_1/NAND4_in[2] ), .A3(n759), .A4(
        \SB1_3_23/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_23/buf_output[1] ) );
  NAND3_X2 U8943 ( .A1(\SB1_0_19/i0_3 ), .A2(\SB1_0_19/i0_4 ), .A3(
        \SB1_0_19/i1[9] ), .ZN(n3900) );
  XOR2_X1 U8945 ( .A1(\MC_ARK_ARC_1_3/temp3[89] ), .A2(
        \MC_ARK_ARC_1_3/temp4[89] ), .Z(\MC_ARK_ARC_1_3/temp6[89] ) );
  XOR2_X1 U8956 ( .A1(\MC_ARK_ARC_1_2/temp4[136] ), .A2(
        \MC_ARK_ARC_1_2/temp2[136] ), .Z(n3902) );
  NAND3_X1 U8971 ( .A1(\SB2_4_3/i0_0 ), .A2(\SB2_4_3/i3[0] ), .A3(
        \SB2_4_3/i1_7 ), .ZN(\SB2_4_3/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U8979 ( .A1(\MC_ARK_ARC_1_2/temp3[151] ), .A2(
        \MC_ARK_ARC_1_2/temp4[151] ), .Z(\MC_ARK_ARC_1_2/temp6[151] ) );
  XOR2_X1 U8987 ( .A1(\MC_ARK_ARC_1_2/temp3[12] ), .A2(
        \MC_ARK_ARC_1_2/temp4[12] ), .Z(n5123) );
  XOR2_X1 U8999 ( .A1(\RI5[4][106] ), .A2(\RI5[4][142] ), .Z(n3904) );
  NAND4_X2 U9001 ( .A1(\SB2_4_8/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_4_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_8/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_4_8/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_4_8/buf_output[1] ) );
  XOR2_X1 U9032 ( .A1(\MC_ARK_ARC_1_3/temp2[149] ), .A2(n3905), .Z(
        \MC_ARK_ARC_1_3/temp5[149] ) );
  XOR2_X1 U9035 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[143] ), .A2(\RI5[3][149] ), 
        .Z(n3905) );
  XOR2_X1 U9039 ( .A1(\MC_ARK_ARC_1_1/temp5[93] ), .A2(n3115), .Z(
        \MC_ARK_ARC_1_1/buf_output[93] ) );
  NAND3_X2 U9062 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i1_7 ), .A3(
        \SB2_1_15/i0[8] ), .ZN(\SB2_1_15/Component_Function_1/NAND4_in[1] ) );
  INV_X2 U9065 ( .I(\SB1_3_15/buf_output[5] ), .ZN(\SB2_3_15/i1_5 ) );
  NAND3_X2 U9068 ( .A1(\SB1_4_12/i0[9] ), .A2(\SB1_4_12/i0_4 ), .A3(
        \SB1_4_12/i0[6] ), .ZN(n3907) );
  NAND3_X1 U9070 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0[8] ), .A3(
        \SB1_3_23/i1_7 ), .ZN(\SB1_3_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U9073 ( .A1(\SB4_20/i0_4 ), .A2(\SB4_20/i0[10] ), .A3(\SB4_20/i0_3 ), .ZN(n3909) );
  XOR2_X1 U9085 ( .A1(\MC_ARK_ARC_1_2/temp5[2] ), .A2(n2819), .Z(
        \MC_ARK_ARC_1_2/buf_output[2] ) );
  NAND3_X2 U9089 ( .A1(\SB1_0_19/i0_3 ), .A2(\SB1_0_19/i1[9] ), .A3(
        \SB1_0_19/i0[6] ), .ZN(n4671) );
  NAND4_X2 U9092 ( .A1(\SB2_2_2/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_2/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_2/Component_Function_4/NAND4_in[3] ), .A4(n3912), .ZN(
        \SB2_2_2/buf_output[4] ) );
  NAND4_X2 U9095 ( .A1(\SB2_3_15/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_15/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_3_15/Component_Function_1/NAND4_in[1] ), .A4(n3914), .ZN(
        \SB2_3_15/buf_output[1] ) );
  NAND3_X1 U9096 ( .A1(\SB1_0_7/i1_7 ), .A2(\SB1_0_7/i0[10] ), .A3(
        \SB1_0_7/i1[9] ), .ZN(\SB1_0_7/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U9100 ( .A1(\SB2_4_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_12/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_4_12/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_4_12/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_4_12/buf_output[4] ) );
  XOR2_X1 U9107 ( .A1(\RI5[2][134] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[98] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[32] ) );
  INV_X1 U9121 ( .I(\RI3[0][5] ), .ZN(\SB2_0_31/i1_5 ) );
  NAND3_X2 U9126 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i0[9] ), .A3(
        \SB2_1_15/i0[8] ), .ZN(n865) );
  BUF_X4 U9129 ( .I(\SB1_1_13/buf_output[5] ), .Z(\SB2_1_13/i0_3 ) );
  NAND3_X1 U9132 ( .A1(\SB1_0_22/i0_3 ), .A2(\SB1_0_22/i0[9] ), .A3(
        \SB1_0_22/i0[10] ), .ZN(\SB1_0_22/Component_Function_4/NAND4_in[2] )
         );
  NAND2_X1 U9142 ( .A1(n5218), .A2(n3919), .ZN(n4130) );
  NAND3_X1 U9147 ( .A1(\SB1_4_15/i0[10] ), .A2(\SB1_4_15/i1_5 ), .A3(
        \SB1_4_15/i1[9] ), .ZN(n3920) );
  XOR2_X1 U9151 ( .A1(\RI5[1][149] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[125] ), 
        .Z(n3921) );
  XOR2_X1 U9158 ( .A1(\RI5[2][184] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[28] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[118] ) );
  NAND4_X2 U9161 ( .A1(\SB2_2_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_30/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_2_30/Component_Function_3/NAND4_in[1] ), .A4(n3923), .ZN(
        \SB2_2_30/buf_output[3] ) );
  INV_X2 U9176 ( .I(\SB1_1_13/buf_output[5] ), .ZN(\SB2_1_13/i1_5 ) );
  NAND3_X2 U9178 ( .A1(\SB2_1_15/i1_5 ), .A2(\SB2_1_15/i0[8] ), .A3(
        \SB2_1_15/i3[0] ), .ZN(\SB2_1_15/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U9183 ( .A1(\SB1_1_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_6/Component_Function_0/NAND4_in[1] ), .A3(n3928), .A4(n3927), 
        .ZN(\SB1_1_6/buf_output[0] ) );
  XOR2_X1 U9191 ( .A1(n1268), .A2(n2425), .Z(n4496) );
  NAND4_X2 U9194 ( .A1(\SB2_4_5/Component_Function_5/NAND4_in[2] ), .A2(n3002), 
        .A3(\SB2_4_5/Component_Function_5/NAND4_in[0] ), .A4(n3930), .ZN(
        \SB2_4_5/buf_output[5] ) );
  NAND3_X2 U9197 ( .A1(\SB2_4_5/i0[10] ), .A2(\SB2_4_5/i0_0 ), .A3(
        \SB2_4_5/i0[6] ), .ZN(n3930) );
  NAND3_X1 U9204 ( .A1(\SB1_0_7/i0_0 ), .A2(\SB1_0_7/i1_7 ), .A3(
        \SB1_0_7/i3[0] ), .ZN(\SB1_0_7/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U9226 ( .A1(\SB1_2_4/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_4/Component_Function_0/NAND4_in[0] ), .A4(n3931), .ZN(
        \SB1_2_4/buf_output[0] ) );
  XOR2_X1 U9227 ( .A1(\RI5[4][83] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[77] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[83] ) );
  XOR2_X1 U9228 ( .A1(\RI5[2][108] ), .A2(\RI5[2][144] ), .Z(
        \MC_ARK_ARC_1_2/temp3[42] ) );
  NAND3_X1 U9230 ( .A1(\SB4_10/i0[9] ), .A2(\SB4_10/i0_3 ), .A3(\SB4_10/i0[8] ), .ZN(n3932) );
  INV_X2 U9234 ( .I(\SB1_3_7/buf_output[5] ), .ZN(\SB2_3_7/i1_5 ) );
  NAND4_X2 U9246 ( .A1(n2476), .A2(\SB2_2_12/Component_Function_0/NAND4_in[1] ), .A3(\SB2_2_12/Component_Function_0/NAND4_in[0] ), .A4(n3933), .ZN(
        \SB2_2_12/buf_output[0] ) );
  XOR2_X1 U9259 ( .A1(n1631), .A2(n4309), .Z(\MC_ARK_ARC_1_2/buf_output[164] )
         );
  BUF_X4 U9260 ( .I(\SB2_4_28/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[23] ) );
  NAND4_X2 U9267 ( .A1(\SB1_3_10/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_3_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_1/NAND4_in[0] ), .A4(n3935), .ZN(
        \SB1_3_10/buf_output[1] ) );
  XOR2_X1 U9273 ( .A1(\RI5[1][65] ), .A2(\RI5[1][89] ), .Z(
        \MC_ARK_ARC_1_1/temp2[119] ) );
  NAND4_X2 U9274 ( .A1(\SB1_3_26/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_3_26/Component_Function_5/NAND4_in[2] ), .A3(n4009), .A4(
        \SB1_3_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_26/buf_output[5] ) );
  NAND4_X2 U9276 ( .A1(\SB1_3_4/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_4/Component_Function_1/NAND4_in[3] ), .A3(n4429), .A4(
        \SB1_3_4/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_4/buf_output[1] ) );
  NAND3_X1 U9281 ( .A1(\SB1_0_28/i0_0 ), .A2(n5433), .A3(\SB1_0_28/i1_5 ), 
        .ZN(\SB1_0_28/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U9285 ( .A1(\SB2_0_8/i0[10] ), .A2(\SB2_0_8/i0_0 ), .A3(
        \SB2_0_8/i0[6] ), .ZN(\SB2_0_8/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U9287 ( .A1(\SB4_0/i0_0 ), .A2(\SB4_0/i0[10] ), .A3(\SB4_0/i0[6] ), 
        .ZN(n3936) );
  NAND3_X2 U9291 ( .A1(\SB2_2_0/i0[8] ), .A2(\SB2_2_0/i1_5 ), .A3(
        \SB2_2_0/i3[0] ), .ZN(\SB2_2_0/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U9297 ( .A1(\SB2_0_3/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_3/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_0_3/Component_Function_2/NAND4_in[2] ), .A4(n5211), .ZN(
        \SB2_0_3/buf_output[2] ) );
  BUF_X4 U9298 ( .I(\MC_ARK_ARC_1_1/buf_output[161] ), .Z(\SB1_2_5/i0_3 ) );
  XOR2_X1 U9300 ( .A1(n3937), .A2(n3942), .Z(\MC_ARK_ARC_1_0/buf_output[29] )
         );
  NAND3_X1 U9307 ( .A1(\SB4_0/i0_0 ), .A2(\SB4_0/i1_7 ), .A3(\SB4_0/i3[0] ), 
        .ZN(n2707) );
  XOR2_X1 U9309 ( .A1(\RI5[4][116] ), .A2(\RI5[4][140] ), .Z(
        \MC_ARK_ARC_1_4/temp2[170] ) );
  NAND3_X2 U9310 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i1[9] ), .A3(
        \SB2_3_20/i1_7 ), .ZN(n3940) );
  INV_X2 U9313 ( .I(\MC_ARK_ARC_1_1/buf_output[161] ), .ZN(\SB1_2_5/i1_5 ) );
  NAND4_X2 U9315 ( .A1(\SB2_2_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_19/Component_Function_3/NAND4_in[3] ), .A4(n3943), .ZN(
        \SB2_2_19/buf_output[3] ) );
  XOR2_X1 U9320 ( .A1(\RI5[1][61] ), .A2(\RI5[1][85] ), .Z(n3946) );
  XOR2_X1 U9327 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[149] ), .A2(\RI5[0][125] ), 
        .Z(n4452) );
  XOR2_X1 U9328 ( .A1(n3951), .A2(n3950), .Z(\MC_ARK_ARC_1_2/temp5[170] ) );
  XOR2_X1 U9329 ( .A1(\RI5[2][170] ), .A2(\RI5[2][140] ), .Z(n3950) );
  NAND4_X2 U9333 ( .A1(\SB2_1_13/Component_Function_0/NAND4_in[3] ), .A2(n3954), .A3(\SB2_1_13/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_1_13/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_1_13/buf_output[0] ) );
  NAND3_X2 U9334 ( .A1(\SB2_1_13/i0[7] ), .A2(\SB2_1_13/i0[8] ), .A3(
        \SB2_1_13/i0[6] ), .ZN(n3954) );
  BUF_X4 U9337 ( .I(\SB2_2_19/buf_output[3] ), .Z(\RI5[2][87] ) );
  XOR2_X1 U9345 ( .A1(n3960), .A2(n74), .Z(Ciphertext[156]) );
  BUF_X4 U9346 ( .I(\SB2_3_30/buf_output[2] ), .Z(\RI5[3][26] ) );
  XOR2_X1 U9349 ( .A1(\RI5[4][111] ), .A2(\RI5[4][147] ), .Z(
        \MC_ARK_ARC_1_4/temp3[45] ) );
  XOR2_X1 U9352 ( .A1(\RI5[2][47] ), .A2(\RI5[2][11] ), .Z(
        \MC_ARK_ARC_1_2/temp3[137] ) );
  NAND3_X2 U9357 ( .A1(\SB2_0_30/i0_3 ), .A2(\SB2_0_30/i0[10] ), .A3(
        \SB2_0_30/i0[9] ), .ZN(n4929) );
  BUF_X4 U9359 ( .I(\SB1_1_30/buf_output[5] ), .Z(\SB2_1_30/i0_3 ) );
  BUF_X4 U9364 ( .I(n409), .Z(\SB1_0_3/i0_3 ) );
  BUF_X2 U9365 ( .I(\SB3_1/buf_output[3] ), .Z(\SB4_31/i0[10] ) );
  NAND3_X2 U9368 ( .A1(\SB2_1_15/i0_4 ), .A2(\SB2_1_15/i1_7 ), .A3(
        \SB2_1_15/i0[8] ), .ZN(n4093) );
  BUF_X4 U9370 ( .I(n407), .Z(\SB1_0_5/i0_3 ) );
  NAND3_X1 U9377 ( .A1(\SB3_8/i0[9] ), .A2(\SB3_8/i0[10] ), .A3(\SB3_8/i0_3 ), 
        .ZN(\SB3_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U9378 ( .A1(\SB3_8/i0_0 ), .A2(\SB3_8/i0[6] ), .A3(\SB3_8/i0[10] ), 
        .ZN(\SB3_8/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U9379 ( .A1(\SB3_8/i0_3 ), .A2(\SB3_8/i0[10] ), .A3(\SB3_8/i0[6] ), 
        .ZN(\SB3_8/Component_Function_2/NAND4_in[1] ) );
  INV_X1 U9382 ( .I(\MC_ARK_ARC_1_4/buf_output[141] ), .ZN(\SB3_8/i0[8] ) );
  BUF_X2 U9383 ( .I(\MC_ARK_ARC_1_4/buf_output[141] ), .Z(\SB3_8/i0[10] ) );
  CLKBUF_X4 U9385 ( .I(\SB3_23/buf_output[4] ), .Z(\SB4_22/i0_4 ) );
  CLKBUF_X4 U9386 ( .I(\MC_ARK_ARC_1_4/buf_output[146] ), .Z(\SB3_7/i0_0 ) );
  NAND3_X1 U9387 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i1_5 ), .A3(\SB4_8/i0_4 ), 
        .ZN(n4332) );
  BUF_X2 U9391 ( .I(\MC_ARK_ARC_1_3/buf_output[90] ), .Z(\SB1_4_16/i0[9] ) );
  INV_X1 U9392 ( .I(\MC_ARK_ARC_1_3/buf_output[90] ), .ZN(\SB1_4_16/i3[0] ) );
  AND4_X2 U9397 ( .A1(\SB3_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_3/NAND4_in[3] ), .Z(n3965) );
  NAND3_X1 U9401 ( .A1(\SB3_22/i0_3 ), .A2(\SB3_22/i0[8] ), .A3(
        \MC_ARK_ARC_1_4/buf_output[54] ), .ZN(
        \SB3_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U9402 ( .A1(\SB3_22/i1_7 ), .A2(\SB3_22/i0[8] ), .A3(\SB3_22/i0_4 ), 
        .ZN(\SB3_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U9403 ( .A1(\SB3_22/i0[8] ), .A2(\SB3_22/i1_5 ), .A3(\SB3_22/i3[0] ), .ZN(n694) );
  NAND3_X1 U9408 ( .A1(\SB3_10/i0_3 ), .A2(\SB3_10/i0[8] ), .A3(\SB3_10/i0[9] ), .ZN(\SB3_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U9409 ( .A1(\SB3_10/i0[7] ), .A2(\SB3_10/i0_3 ), .A3(\SB3_10/i0_0 ), 
        .ZN(\SB3_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U9413 ( .A1(\SB3_20/i0_3 ), .A2(\SB3_20/i0[9] ), .A3(\SB3_20/i0[8] ), .ZN(n5100) );
  NAND3_X1 U9417 ( .A1(\SB4_16/i0_4 ), .A2(\SB4_16/i0_3 ), .A3(\SB4_16/i1[9] ), 
        .ZN(\SB4_16/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U9424 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i1[9] ), .ZN(
        \SB3_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U9425 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i0_3 ), .A3(\SB4_22/i0[7] ), 
        .ZN(n1746) );
  CLKBUF_X4 U9430 ( .I(\SB3_4/buf_output[5] ), .Z(\SB4_4/i0_3 ) );
  BUF_X4 U9431 ( .I(n3980), .Z(\SB3_31/i0_3 ) );
  INV_X1 U9437 ( .I(\MC_ARK_ARC_1_4/buf_output[169] ), .ZN(\SB3_3/i1_7 ) );
  CLKBUF_X4 U9440 ( .I(\SB3_22/buf_output[1] ), .Z(\SB4_18/i0[6] ) );
  BUF_X4 U9443 ( .I(n3968), .Z(\SB1_4_6/i0[10] ) );
  BUF_X4 U9444 ( .I(\SB2_4_28/buf_output[2] ), .Z(\RI5[4][38] ) );
  NAND3_X1 U9445 ( .A1(\SB2_4_27/i3[0] ), .A2(\SB2_4_27/i1_5 ), .A3(
        \SB2_4_27/i0[8] ), .ZN(n1429) );
  NAND3_X1 U9446 ( .A1(\SB2_4_27/i0[8] ), .A2(\SB2_4_27/i0[7] ), .A3(
        \SB2_4_27/i0[6] ), .ZN(\SB2_4_27/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U9449 ( .A1(\SB3_5/i1[9] ), .A2(\SB3_5/i0_4 ), .A3(\SB3_5/i0_3 ), 
        .ZN(\SB3_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U9450 ( .A1(\SB3_5/i0[9] ), .A2(\SB3_5/i0[10] ), .A3(\SB3_5/i0_3 ), 
        .ZN(\SB3_5/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U9452 ( .I(\MC_ARK_ARC_1_3/buf_output[85] ), .ZN(\SB1_4_17/i1_7 ) );
  CLKBUF_X4 U9453 ( .I(\MC_ARK_ARC_1_3/buf_output[85] ), .Z(\SB1_4_17/i0[6] )
         );
  CLKBUF_X4 U9456 ( .I(\MC_ARK_ARC_1_2/buf_output[86] ), .Z(\SB1_3_17/i0_0 )
         );
  INV_X1 U9457 ( .I(\MC_ARK_ARC_1_3/buf_output[185] ), .ZN(\SB1_4_1/i1_5 ) );
  NAND3_X1 U9461 ( .A1(n5442), .A2(\SB4_1/i0[6] ), .A3(\SB4_1/i0[9] ), .ZN(
        \SB4_1/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 U9462 ( .I(\SB2_3_19/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[102] ) );
  NAND3_X1 U9465 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i0[7] ), .A3(\SB4_23/i0_3 ), 
        .ZN(\SB4_23/Component_Function_0/NAND4_in[3] ) );
  INV_X1 U9469 ( .I(\SB3_0/buf_output[0] ), .ZN(\SB4_27/i3[0] ) );
  NAND3_X1 U9470 ( .A1(\SB3_21/i0[10] ), .A2(\SB3_21/i1[9] ), .A3(
        \SB3_21/i1_7 ), .ZN(n4989) );
  INV_X1 U9475 ( .I(n3974), .ZN(n3966) );
  NAND3_X1 U9476 ( .A1(\SB4_13/i0[6] ), .A2(\SB4_13/i0_3 ), .A3(\SB4_13/i1[9] ), .ZN(n1916) );
  NAND3_X1 U9478 ( .A1(\SB4_13/i0[6] ), .A2(n4002), .A3(\SB4_13/i0[9] ), .ZN(
        \SB4_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U9479 ( .A1(\SB4_4/i0_0 ), .A2(\SB4_4/i0[6] ), .A3(\SB4_4/i0[10] ), 
        .ZN(\SB4_4/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U9480 ( .A1(\MC_ARK_ARC_1_3/temp6[153] ), .A2(
        \MC_ARK_ARC_1_3/temp5[153] ), .Z(n3967) );
  NAND3_X1 U9482 ( .A1(\SB4_1/i0_4 ), .A2(\SB4_1/i1_7 ), .A3(\SB4_1/i0[8] ), 
        .ZN(n4735) );
  NAND3_X1 U9486 ( .A1(\SB3_10/i0[10] ), .A2(\SB3_10/i1[9] ), .A3(
        \SB3_10/i1_7 ), .ZN(\SB3_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U9491 ( .A1(\SB4_4/i0_3 ), .A2(\SB4_4/i1[9] ), .A3(\SB4_4/i0[6] ), 
        .ZN(n5209) );
  CLKBUF_X4 U9494 ( .I(\MC_ARK_ARC_1_3/buf_output[118] ), .Z(\SB1_4_12/i0_4 )
         );
  NAND3_X1 U9495 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i0_4 ), .A3(\SB3_19/i1[9] ), 
        .ZN(n2337) );
  XOR2_X1 U9497 ( .A1(\MC_ARK_ARC_1_4/temp6[125] ), .A2(
        \MC_ARK_ARC_1_4/temp5[125] ), .Z(n3970) );
  NAND3_X1 U9498 ( .A1(\RI1[4][119] ), .A2(\SB1_4_12/i0[7] ), .A3(
        \SB1_4_12/i0_0 ), .ZN(\SB1_4_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U9499 ( .A1(\SB1_4_12/i0[10] ), .A2(\SB1_4_12/i0[6] ), .A3(
        \SB1_4_12/i0_0 ), .ZN(\SB1_4_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U9500 ( .A1(\SB2_4_27/i0_0 ), .A2(\SB2_4_27/i1_5 ), .A3(
        \SB1_4_28/buf_output[4] ), .ZN(
        \SB2_4_27/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 U9501 ( .A1(\SB2_4_27/i0_0 ), .A2(\SB2_4_27/i3[0] ), .ZN(
        \SB2_4_27/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U9502 ( .I(\SB1_4_30/buf_output[2] ), .Z(\SB2_4_27/i0_0 ) );
  NAND3_X1 U9504 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0[10] ), .A3(
        \SB3_30/i0[6] ), .ZN(\SB3_30/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U9505 ( .I(\SB2_4_12/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[129] ) );
  BUF_X2 U9506 ( .I(\MC_ARK_ARC_1_3/buf_output[62] ), .Z(\SB1_4_21/i0_0 ) );
  INV_X1 U9507 ( .I(\MC_ARK_ARC_1_3/buf_output[62] ), .ZN(\SB1_4_21/i1[9] ) );
  BUF_X2 U9508 ( .I(\MC_ARK_ARC_1_4/buf_output[30] ), .Z(\SB3_26/i0[9] ) );
  CLKBUF_X4 U9509 ( .I(\SB1_4_22/buf_output[2] ), .Z(\SB2_4_19/i0_0 ) );
  INV_X1 U9510 ( .I(\MC_ARK_ARC_1_4/buf_output[55] ), .ZN(\SB3_22/i1_7 ) );
  INV_X1 U9514 ( .I(\SB3_3/buf_output[5] ), .ZN(\SB4_3/i1_5 ) );
  NAND3_X1 U9516 ( .A1(\SB4_3/i0[6] ), .A2(\SB4_3/i0_0 ), .A3(\SB4_3/i0[10] ), 
        .ZN(n2522) );
  NAND3_X1 U9517 ( .A1(\SB4_3/i0_0 ), .A2(\SB4_3/i0_4 ), .A3(\SB4_3/i1_5 ), 
        .ZN(n1828) );
  NAND3_X1 U9518 ( .A1(\RI1[4][59] ), .A2(\SB1_4_22/i0[8] ), .A3(
        \SB1_4_22/i1_7 ), .ZN(\SB1_4_22/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X4 U9519 ( .I(\MC_ARK_ARC_1_1/buf_output[136] ), .Z(\SB1_2_9/i0_4 )
         );
  NAND3_X1 U9520 ( .A1(\SB3_18/i0_0 ), .A2(\SB3_18/i1_5 ), .A3(\SB3_18/i0_4 ), 
        .ZN(\SB3_18/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U9521 ( .A1(\SB1_4_8/i0[10] ), .A2(\SB1_4_8/i1[9] ), .A3(
        \SB1_4_8/i1_7 ), .ZN(\SB1_4_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U9528 ( .A1(\SB3_27/i1[9] ), .A2(\SB3_27/i1_7 ), .A3(
        \SB3_27/i0[10] ), .ZN(\SB3_27/Component_Function_3/NAND4_in[2] ) );
  INV_X1 U9529 ( .I(\SB3_5/buf_output[1] ), .ZN(\SB4_1/i1_7 ) );
  XOR2_X1 U9530 ( .A1(\MC_ARK_ARC_1_4/temp5[47] ), .A2(
        \MC_ARK_ARC_1_4/temp6[47] ), .Z(n3971) );
  CLKBUF_X4 U9536 ( .I(\SB2_2_18/buf_output[0] ), .Z(\RI5[2][108] ) );
  BUF_X4 U9537 ( .I(n3992), .Z(\SB1_4_30/i0_3 ) );
  NAND2_X1 U9539 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i3[0] ), .ZN(
        \SB4_14/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U9540 ( .I(\MC_ARK_ARC_1_3/buf_output[168] ), .ZN(\SB1_4_3/i3[0] ) );
  BUF_X2 U9541 ( .I(\MC_ARK_ARC_1_3/buf_output[168] ), .Z(\SB1_4_3/i0[9] ) );
  NAND3_X1 U9546 ( .A1(\SB4_27/i0_0 ), .A2(\SB4_27/i3[0] ), .A3(\SB4_27/i1_7 ), 
        .ZN(\SB4_27/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 U9547 ( .A1(\SB4_27/i0_0 ), .A2(\SB4_27/i3[0] ), .ZN(
        \SB4_27/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U9550 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i1[9] ), .ZN(
        \SB3_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U9551 ( .A1(\SB3_31/i1_5 ), .A2(\SB3_31/i0_4 ), .A3(\SB3_31/i1[9] ), 
        .ZN(\SB3_31/Component_Function_4/NAND4_in[3] ) );
  AND4_X2 U9553 ( .A1(\SB3_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_1/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_1/Component_Function_2/NAND4_in[1] ), .A4(n4293), .Z(n3973) );
  CLKBUF_X4 U9554 ( .I(\MC_ARK_ARC_1_3/buf_output[8] ), .Z(\SB1_4_30/i0_0 ) );
  CLKBUF_X4 U9555 ( .I(\MC_ARK_ARC_1_4/buf_output[56] ), .Z(\SB3_22/i0_0 ) );
  NAND3_X1 U9556 ( .A1(\SB4_3/i0[10] ), .A2(\SB4_3/i1_5 ), .A3(\SB4_3/i1[9] ), 
        .ZN(n4953) );
  NAND3_X2 U9558 ( .A1(\SB2_4_20/i0_3 ), .A2(\SB2_4_20/i0[10] ), .A3(
        \SB2_4_20/i0[6] ), .ZN(\SB2_4_20/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 U9559 ( .A1(n2717), .A2(n4685), .ZN(n4792) );
  NAND2_X1 U9561 ( .A1(\SB4_4/i0_0 ), .A2(\SB4_4/i3[0] ), .ZN(
        \SB4_4/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U9562 ( .A1(\SB3_15/buf_output[3] ), .A2(\SB4_13/i0[9] ), .ZN(
        \SB4_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U9563 ( .A1(\SB4_13/i0_3 ), .A2(\SB3_15/buf_output[3] ), .A3(
        \SB4_13/i0_4 ), .ZN(n729) );
  NAND3_X1 U9565 ( .A1(\SB2_4_9/i0_0 ), .A2(\SB2_4_9/i0[6] ), .A3(
        \SB2_4_9/i0[10] ), .ZN(\SB2_4_9/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X4 U9567 ( .I(\SB1_4_12/buf_output[2] ), .Z(\SB2_4_9/i0_0 ) );
  NAND3_X1 U9569 ( .A1(\RI1[2][149] ), .A2(\SB1_2_7/i1_7 ), .A3(n3184), .ZN(
        \SB1_2_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U9573 ( .A1(\SB3_0/i0[10] ), .A2(\SB3_0/i0[9] ), .ZN(
        \SB3_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U9574 ( .A1(\SB3_0/i0[10] ), .A2(\SB3_0/i0_4 ), .A3(\SB3_0/i0_3 ), 
        .ZN(\SB3_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U9577 ( .A1(\SB3_21/i0_0 ), .A2(\SB3_21/i0[6] ), .A3(
        \SB3_21/i0[10] ), .ZN(\SB3_21/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U9578 ( .A1(n3182), .A2(\SB3_21/i0[10] ), .A3(\SB3_21/i1[9] ), .ZN(
        \SB3_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U9579 ( .A1(\SB3_21/i0[9] ), .A2(\SB3_21/i0[10] ), .A3(
        \SB3_21/i0_3 ), .ZN(\SB3_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U9580 ( .A1(\SB4_17/i0[7] ), .A2(\SB4_17/i0_3 ), .A3(\SB4_17/i0_0 ), 
        .ZN(\SB4_17/Component_Function_0/NAND4_in[3] ) );
  INV_X1 U9585 ( .I(\SB1_4_15/buf_output[1] ), .ZN(\SB2_4_11/i1_7 ) );
  NAND3_X1 U9588 ( .A1(\SB2_4_6/i0[9] ), .A2(\SB2_4_6/i0[10] ), .A3(
        \SB2_4_6/i0_3 ), .ZN(\SB2_4_6/Component_Function_4/NAND4_in[2] ) );
  CLKBUF_X4 U9590 ( .I(\MC_ARK_ARC_1_4/buf_output[7] ), .Z(\SB3_30/i0[6] ) );
  INV_X1 U9591 ( .I(\MC_ARK_ARC_1_4/buf_output[7] ), .ZN(\SB3_30/i1_7 ) );
  CLKBUF_X4 U9595 ( .I(\SB2_4_9/buf_output[1] ), .Z(\RI5[4][157] ) );
  NAND3_X1 U9599 ( .A1(\SB3_30/i0[10] ), .A2(\SB3_30/i0_0 ), .A3(
        \SB3_30/i0[6] ), .ZN(\SB3_30/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X12 U9603 ( .I(\MC_ARK_ARC_1_4/buf_output[17] ), .Z(\RI1[5][17] ) );
  NAND3_X1 U9607 ( .A1(\SB3_26/i1[9] ), .A2(\SB3_26/i0_3 ), .A3(\SB3_26/i0[6] ), .ZN(\SB3_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U9608 ( .A1(\SB3_26/i0_3 ), .A2(\SB3_26/i0_0 ), .A3(\SB3_26/i0_4 ), 
        .ZN(\SB3_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U9609 ( .A1(\SB2_3_29/i0[10] ), .A2(\SB2_3_29/i1[9] ), .A3(
        \SB2_3_29/i1_7 ), .ZN(n2972) );
  BUF_X4 U9611 ( .I(\SB2_2_20/buf_output[2] ), .Z(\RI5[2][86] ) );
  NAND2_X1 U9616 ( .A1(\SB2_1_1/i0_0 ), .A2(\SB2_1_1/i3[0] ), .ZN(
        \SB2_1_1/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U9619 ( .I(\RI3[0][188] ), .Z(\SB2_0_0/i0_0 ) );
  NAND3_X1 U9622 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i1[9] ), .A3(
        \SB2_2_11/i1_5 ), .ZN(n5170) );
  NAND3_X1 U9623 ( .A1(\SB2_2_11/i1[9] ), .A2(\SB2_2_11/i1_7 ), .A3(
        \SB2_2_11/i0[10] ), .ZN(\SB2_2_11/Component_Function_3/NAND4_in[2] )
         );
  CLKBUF_X4 U9628 ( .I(\MC_ARK_ARC_1_4/buf_output[104] ), .Z(\SB3_14/i0_0 ) );
  NAND3_X1 U9630 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i3[0] ), .A3(\SB4_1/i1_7 ), 
        .ZN(n2562) );
  NAND3_X1 U9631 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i0[6] ), .A3(\SB4_1/i0[10] ), 
        .ZN(\SB4_1/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U9636 ( .I(\SB2_3_29/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[32] ) );
  CLKBUF_X4 U9637 ( .I(\SB3_18/buf_output[5] ), .Z(\SB4_18/i0_3 ) );
  BUF_X2 U9638 ( .I(\SB3_10/buf_output[2] ), .Z(\SB4_7/i0_0 ) );
  INV_X1 U9639 ( .I(\SB3_10/buf_output[2] ), .ZN(\SB4_7/i1[9] ) );
  CLKBUF_X4 U9640 ( .I(n386), .Z(\SB1_0_26/i0_3 ) );
  XOR2_X1 U9642 ( .A1(\MC_ARK_ARC_1_4/temp6[5] ), .A2(
        \MC_ARK_ARC_1_4/temp5[5] ), .Z(n3981) );
  NAND3_X1 U9645 ( .A1(\SB1_0_1/i0_0 ), .A2(\SB1_0_1/i1_5 ), .A3(
        \SB1_0_1/i0_4 ), .ZN(n2181) );
  CLKBUF_X4 U9648 ( .I(\SB3_6/buf_output[3] ), .Z(\SB4_4/i0[10] ) );
  NAND3_X1 U9649 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB2_3_19/i0[8] ), .A3(
        \SB2_3_19/i1_7 ), .ZN(\SB2_3_19/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U9652 ( .A1(\SB1_3_26/i0_0 ), .A2(\MC_ARK_ARC_1_2/buf_output[34] ), 
        .A3(\SB1_3_26/i1_5 ), .ZN(\SB1_3_26/Component_Function_2/NAND4_in[3] )
         );
  XOR2_X1 U9653 ( .A1(\MC_ARK_ARC_1_2/temp5[2] ), .A2(n2819), .Z(n3982) );
  AND4_X1 U9654 ( .A1(\SB1_4_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_4_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_3/Component_Function_0/NAND4_in[3] ), .Z(n3983) );
  NAND3_X1 U9656 ( .A1(\SB1_4_3/i0[7] ), .A2(\SB1_4_3/i0_3 ), .A3(
        \SB1_4_3/i0_0 ), .ZN(\SB1_4_3/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U9657 ( .A1(\SB4_18/i0_3 ), .A2(n1496), .ZN(
        \SB4_18/Component_Function_1/NAND4_in[0] ) );
  CLKBUF_X4 U9658 ( .I(\MC_ARK_ARC_1_4/buf_output[64] ), .Z(\SB3_21/i0_4 ) );
  XOR2_X1 U9659 ( .A1(Key[65]), .A2(Plaintext[65]), .Z(n3985) );
  NAND3_X1 U9662 ( .A1(\SB1_2_3/i1[9] ), .A2(\SB1_2_3/i0_3 ), .A3(
        \SB1_2_3/i0[6] ), .ZN(\SB1_2_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U9663 ( .A1(\SB1_1_5/i1_7 ), .A2(\SB1_1_5/i0[8] ), .A3(
        \SB1_1_5/i0_4 ), .ZN(\SB1_1_5/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 U9664 ( .I(\SB3_26/buf_output[4] ), .Z(\SB4_25/i0_4 ) );
  NAND3_X1 U9665 ( .A1(\SB2_0_7/i1[9] ), .A2(\SB2_0_7/i1_5 ), .A3(
        \RI3[0][148] ), .ZN(\SB2_0_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U9669 ( .A1(\SB1_1_28/i1_5 ), .A2(\SB1_1_28/i0[6] ), .A3(
        \SB1_1_28/i0[9] ), .ZN(\SB1_1_28/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U9671 ( .A1(\SB1_4_14/i0_3 ), .A2(\SB1_4_14/i1[9] ), .ZN(n1106) );
  NAND3_X1 U9672 ( .A1(\SB1_4_14/i0[10] ), .A2(\SB1_4_14/i0_4 ), .A3(
        \SB1_4_14/i0_3 ), .ZN(\SB1_4_14/Component_Function_0/NAND4_in[2] ) );
  INV_X1 U9682 ( .I(\MC_ARK_ARC_1_0/buf_output[168] ), .ZN(\SB1_1_3/i3[0] ) );
  XOR2_X1 U9683 ( .A1(n2936), .A2(\MC_ARK_ARC_1_2/temp6[65] ), .Z(n3986) );
  XOR2_X1 U9684 ( .A1(n2936), .A2(\MC_ARK_ARC_1_2/temp6[65] ), .Z(n3987) );
  BUF_X4 U9685 ( .I(\SB2_1_31/buf_output[2] ), .Z(\RI5[1][20] ) );
  CLKBUF_X4 U9686 ( .I(\SB2_3_26/buf_output[0] ), .Z(\RI5[3][60] ) );
  NAND3_X1 U9689 ( .A1(\SB4_30/i0[6] ), .A2(\SB4_30/i0_4 ), .A3(
        \SB3_3/buf_output[0] ), .ZN(n2594) );
  NAND3_X1 U9690 ( .A1(n5427), .A2(\SB4_30/i0[9] ), .A3(\SB4_30/i0[8] ), .ZN(
        n1424) );
  NAND3_X1 U9692 ( .A1(\SB4_22/i0[9] ), .A2(\SB4_22/i0[10] ), .A3(
        \SB4_22/i0_3 ), .ZN(\SB4_22/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U9693 ( .A1(\SB4_22/i0_4 ), .A2(\SB4_22/i0_3 ), .A3(\SB4_22/i1[9] ), 
        .ZN(\SB4_22/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U9695 ( .I(\SB1_4_6/buf_output[1] ), .Z(\SB2_4_2/i0[6] ) );
  CLKBUF_X4 U9698 ( .I(\SB1_3_19/buf_output[3] ), .Z(\SB2_3_17/i0[10] ) );
  NAND3_X1 U9699 ( .A1(\SB2_2_19/i1[9] ), .A2(\SB2_2_19/i0_3 ), .A3(
        \SB2_2_19/i0[6] ), .ZN(\SB2_2_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U9701 ( .A1(\SB2_2_19/i1[9] ), .A2(\SB2_2_19/i1_5 ), .A3(
        \SB1_2_20/buf_output[4] ), .ZN(
        \SB2_2_19/Component_Function_4/NAND4_in[3] ) );
  AND4_X2 U9704 ( .A1(n2584), .A2(\SB1_4_3/Component_Function_5/NAND4_in[1] ), 
        .A3(n1142), .A4(\SB1_4_3/Component_Function_5/NAND4_in[0] ), .Z(n3988)
         );
  INV_X1 U9706 ( .I(\SB1_1_1/buf_output[0] ), .ZN(\SB2_1_28/i3[0] ) );
  INV_X1 U9708 ( .I(\MC_ARK_ARC_1_3/buf_output[91] ), .ZN(\SB1_4_16/i1_7 ) );
  CLKBUF_X4 U9709 ( .I(\MC_ARK_ARC_1_4/buf_output[87] ), .Z(\SB3_17/i0[10] )
         );
  NAND3_X1 U9710 ( .A1(\SB1_0_14/i0_4 ), .A2(\SB1_0_14/i1[9] ), .A3(
        \SB1_0_14/i0_3 ), .ZN(\SB1_0_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U9711 ( .A1(\SB1_0_14/i0_3 ), .A2(\SB1_0_14/i0[10] ), .A3(n238), 
        .ZN(\SB1_0_14/Component_Function_2/NAND4_in[1] ) );
  AND4_X2 U9714 ( .A1(\SB1_1_17/Component_Function_5/NAND4_in[3] ), .A2(n1187), 
        .A3(\SB1_1_17/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_1_17/Component_Function_5/NAND4_in[0] ), .Z(n3990) );
  INV_X1 U9717 ( .I(n383), .ZN(\SB1_0_29/i1_5 ) );
  CLKBUF_X4 U9718 ( .I(\SB1_1_4/buf_output[1] ), .Z(\SB2_1_0/i0[6] ) );
  NAND3_X1 U9719 ( .A1(\SB4_1/i0_4 ), .A2(\SB4_1/i0_3 ), .A3(\SB4_1/i1[9] ), 
        .ZN(n4682) );
  XOR2_X1 U9720 ( .A1(n2950), .A2(\MC_ARK_ARC_1_3/temp6[11] ), .Z(n3992) );
  XOR2_X1 U9721 ( .A1(\MC_ARK_ARC_1_3/temp6[11] ), .A2(n2950), .Z(n3993) );
  AND4_X2 U9724 ( .A1(n2595), .A2(\SB1_2_3/Component_Function_5/NAND4_in[2] ), 
        .A3(n5394), .A4(\SB1_2_3/Component_Function_5/NAND4_in[0] ), .Z(n3994)
         );
  NAND3_X1 U9727 ( .A1(\SB2_2_6/i0_4 ), .A2(\SB2_2_6/i1_5 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(n641) );
  NAND3_X1 U9728 ( .A1(\SB1_2_9/i0_4 ), .A2(\SB1_2_9/i1_5 ), .A3(
        \SB1_2_9/i0_0 ), .ZN(\SB1_2_9/Component_Function_2/NAND4_in[3] ) );
  AND4_X2 U9729 ( .A1(\SB1_1_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_27/Component_Function_3/NAND4_in[3] ), .A4(n4067), .Z(n3995) );
  NAND3_X1 U9731 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i1_7 ), .A3(
        \SB2_0_11/i0[8] ), .ZN(\SB2_0_11/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U9735 ( .I(\RI3[0][173] ), .Z(\SB2_0_3/i0_3 ) );
  NAND3_X1 U9739 ( .A1(\SB2_0_4/i0[9] ), .A2(\SB2_0_4/i0[8] ), .A3(
        \SB2_0_4/i0_0 ), .ZN(n4612) );
  CLKBUF_X4 U9740 ( .I(\MC_ARK_ARC_1_0/buf_output[182] ), .Z(\SB1_1_1/i0_0 )
         );
  NAND3_X1 U9741 ( .A1(\SB4_0/i0_3 ), .A2(\SB4_0/i0[9] ), .A3(\SB4_0/i0[10] ), 
        .ZN(\SB4_0/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U9742 ( .I(\SB1_3_23/buf_output[1] ), .ZN(\SB2_3_19/i1_7 ) );
  CLKBUF_X4 U9743 ( .I(\MC_ARK_ARC_1_4/buf_output[50] ), .Z(\SB3_23/i0_0 ) );
  INV_X1 U9745 ( .I(\MC_ARK_ARC_1_2/buf_output[13] ), .ZN(\SB1_3_29/i1_7 ) );
  NAND4_X2 U9748 ( .A1(\SB2_1_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_23/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_23/Component_Function_2/NAND4_in[2] ), .A4(n1838), .ZN(
        \SB2_1_23/buf_output[2] ) );
  BUF_X2 U9749 ( .I(\MC_ARK_ARC_1_1/buf_output[51] ), .Z(\SB1_2_23/i0[10] ) );
  INV_X1 U9750 ( .I(\MC_ARK_ARC_1_1/buf_output[51] ), .ZN(\SB1_2_23/i0[8] ) );
  BUF_X2 U9753 ( .I(\MC_ARK_ARC_1_2/buf_output[98] ), .Z(\SB1_3_15/i0_0 ) );
  INV_X1 U9754 ( .I(\MC_ARK_ARC_1_2/buf_output[98] ), .ZN(\SB1_3_15/i1[9] ) );
  CLKBUF_X4 U9755 ( .I(\SB3_1/buf_output[0] ), .Z(\SB4_28/i0[9] ) );
  NAND3_X1 U9759 ( .A1(\SB3_13/i0[10] ), .A2(\SB3_13/i1[9] ), .A3(
        \SB3_13/i1_7 ), .ZN(n2579) );
  CLKBUF_X4 U9760 ( .I(\SB1_4_29/buf_output[0] ), .Z(\SB2_4_24/i0[9] ) );
  NAND2_X1 U9761 ( .A1(\SB2_4_24/i0_0 ), .A2(\SB2_4_24/i3[0] ), .ZN(
        \SB2_4_24/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U9762 ( .I(\MC_ARK_ARC_1_2/buf_output[30] ), .ZN(\SB1_3_26/i3[0] ) );
  NAND4_X2 U9764 ( .A1(\SB3_1/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_1/Component_Function_5/NAND4_in[2] ), .A3(n2627), .A4(
        \SB3_1/Component_Function_5/NAND4_in[0] ), .ZN(n3999) );
  NAND3_X2 U9766 ( .A1(\SB3_1/i0[6] ), .A2(\SB3_1/i0_4 ), .A3(\SB3_1/i0[9] ), 
        .ZN(n2627) );
  AND4_X2 U9767 ( .A1(\SB1_4_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_4_30/Component_Function_3/NAND4_in[3] ), .A4(n4125), .Z(n4000) );
  NAND3_X1 U9768 ( .A1(\SB1_1_30/i1[9] ), .A2(\SB1_1_30/i0_3 ), .A3(
        \SB1_1_30/i0[6] ), .ZN(\SB1_1_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U9769 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i1[9] ), .A3(
        \SB1_1_30/i0_4 ), .ZN(\SB1_1_30/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U9771 ( .I(\RI3[0][176] ), .Z(\SB2_0_2/i0_0 ) );
  NAND3_X1 U9774 ( .A1(\SB3_0/i1[9] ), .A2(\SB3_0/i1_5 ), .A3(\SB3_0/i0_4 ), 
        .ZN(\SB3_0/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U9775 ( .I(\SB1_3_14/buf_output[2] ), .Z(\SB2_3_11/i0_0 ) );
  CLKBUF_X4 U9781 ( .I(n6276), .Z(\SB1_3_1/i0[10] ) );
  XOR2_X1 U9784 ( .A1(\MC_ARK_ARC_1_4/temp5[111] ), .A2(
        \MC_ARK_ARC_1_4/temp6[111] ), .Z(n4001) );
  INV_X1 U9786 ( .I(\MC_ARK_ARC_1_2/buf_output[131] ), .ZN(\SB1_3_10/i1_5 ) );
  CLKBUF_X4 U9788 ( .I(n3999), .Z(\SB4_1/i0_3 ) );
  OR3_X2 U9789 ( .A1(\RI1[5][113] ), .A2(\MC_ARK_ARC_1_4/buf_output[111] ), 
        .A3(\MC_ARK_ARC_1_4/buf_output[108] ), .Z(n736) );
  INV_X1 U9794 ( .I(\MC_ARK_ARC_1_0/buf_output[48] ), .ZN(\SB1_1_23/i3[0] ) );
  XOR2_X1 U9796 ( .A1(n4124), .A2(n4123), .Z(n4004) );
  INV_X1 U9803 ( .I(n407), .ZN(\SB1_0_5/i1_5 ) );
  INV_X1 U9807 ( .I(\MC_ARK_ARC_1_3/buf_output[97] ), .ZN(\SB1_4_15/i1_7 ) );
  XOR2_X1 U9808 ( .A1(n2441), .A2(\MC_ARK_ARC_1_4/temp6[161] ), .Z(n4006) );
  INV_X1 U9810 ( .I(\SB1_1_11/buf_output[1] ), .ZN(\SB2_1_7/i1_7 ) );
  NAND3_X2 U9814 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0[8] ), .A3(
        \SB1_1_22/i1_7 ), .ZN(\SB1_1_22/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U9816 ( .A1(n4010), .A2(\MC_ARK_ARC_1_1/temp5[184] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[184] ) );
  XOR2_X1 U9817 ( .A1(\MC_ARK_ARC_1_1/temp4[184] ), .A2(
        \MC_ARK_ARC_1_1/temp3[184] ), .Z(n4010) );
  NAND4_X2 U9818 ( .A1(\SB2_2_3/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_3/Component_Function_5/NAND4_in[0] ), .A3(
        \SB2_2_3/Component_Function_5/NAND4_in[1] ), .A4(n5326), .ZN(
        \SB2_2_3/buf_output[5] ) );
  NAND4_X2 U9822 ( .A1(n3097), .A2(\SB2_4_4/Component_Function_5/NAND4_in[1] ), 
        .A3(n1682), .A4(\SB2_4_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_4_4/buf_output[5] ) );
  XOR2_X1 U9823 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[83] ), .A2(\RI5[1][113] ), 
        .Z(n4458) );
  NAND3_X2 U9824 ( .A1(\SB1_2_3/i0[6] ), .A2(\SB1_2_3/i0[10] ), .A3(
        \SB1_2_3/i0_0 ), .ZN(n5394) );
  XOR2_X1 U9826 ( .A1(\RI5[2][47] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[23] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[77] ) );
  NAND3_X2 U9828 ( .A1(\SB1_2_12/i1[9] ), .A2(\SB1_2_12/i0[6] ), .A3(
        \RI1[2][119] ), .ZN(n4012) );
  NAND2_X1 U9831 ( .A1(\SB2_2_17/i0[9] ), .A2(\SB2_2_17/i0[10] ), .ZN(
        \SB2_2_17/Component_Function_0/NAND4_in[0] ) );
  INV_X2 U9832 ( .I(\SB1_4_8/buf_output[5] ), .ZN(\SB2_4_8/i1_5 ) );
  XOR2_X1 U9837 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[149] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[173] ), .Z(n4015) );
  XOR2_X1 U9838 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[7] ), .A2(\RI5[2][13] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[13] ) );
  XOR2_X1 U9841 ( .A1(n4018), .A2(\MC_ARK_ARC_1_2/temp6[46] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[46] ) );
  XOR2_X1 U9842 ( .A1(\MC_ARK_ARC_1_2/temp2[46] ), .A2(
        \MC_ARK_ARC_1_2/temp1[46] ), .Z(n4018) );
  INV_X1 U9843 ( .I(\SB1_4_12/buf_output[1] ), .ZN(\SB2_4_8/i1_7 ) );
  NAND4_X2 U9844 ( .A1(n4824), .A2(\SB1_4_12/Component_Function_1/NAND4_in[3] ), .A3(\SB1_4_12/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_4_12/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_4_12/buf_output[1] ) );
  NAND3_X1 U9845 ( .A1(\SB1_2_28/i0_3 ), .A2(\SB1_2_28/i0[8] ), .A3(
        \SB1_2_28/i1_7 ), .ZN(\SB1_2_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U9848 ( .A1(\SB1_3_20/i0[6] ), .A2(\SB1_3_20/i0_0 ), .A3(
        \SB1_3_20/i0[10] ), .ZN(n4020) );
  XOR2_X1 U9853 ( .A1(n4022), .A2(n187), .Z(Ciphertext[113]) );
  NAND4_X2 U9854 ( .A1(\SB4_13/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_13/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_13/Component_Function_5/NAND4_in[0] ), .A4(n792), .ZN(n4022) );
  XOR2_X1 U9857 ( .A1(\SB2_0_3/buf_output[2] ), .A2(\RI5[0][182] ), .Z(
        \MC_ARK_ARC_1_0/temp1[188] ) );
  NAND3_X2 U9859 ( .A1(\SB2_1_3/i0[6] ), .A2(\SB2_1_3/i0[10] ), .A3(
        \SB2_1_3/i0_0 ), .ZN(n4023) );
  XOR2_X1 U9864 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[183] ), .A2(\RI5[2][177] ), 
        .Z(n4026) );
  INV_X2 U9865 ( .I(\SB1_3_6/buf_output[2] ), .ZN(\SB2_3_3/i1[9] ) );
  NAND4_X2 U9866 ( .A1(n1772), .A2(\SB1_3_6/Component_Function_2/NAND4_in[1] ), 
        .A3(n4449), .A4(n3068), .ZN(\SB1_3_6/buf_output[2] ) );
  NAND3_X2 U9868 ( .A1(\SB2_2_8/i0_0 ), .A2(\SB2_2_8/i1_5 ), .A3(
        \SB2_2_8/i0_4 ), .ZN(n4028) );
  XOR2_X1 U9872 ( .A1(\RI5[4][95] ), .A2(\RI5[4][119] ), .Z(n4031) );
  NAND4_X2 U9873 ( .A1(n1940), .A2(\SB1_4_10/Component_Function_0/NAND4_in[1] ), .A3(\SB1_4_10/Component_Function_0/NAND4_in[0] ), .A4(n4033), .ZN(
        \SB1_4_10/buf_output[0] ) );
  NAND4_X2 U9877 ( .A1(\SB2_0_3/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_3/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_3/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_3/Component_Function_5/NAND4_in[0] ), .ZN(\RI5[0][173] ) );
  XOR2_X1 U9878 ( .A1(n1947), .A2(\MC_ARK_ARC_1_3/temp6[119] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[119] ) );
  XOR2_X1 U9884 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[53] ), .A2(\RI5[4][89] ), 
        .Z(n4037) );
  XOR2_X1 U9885 ( .A1(\RI5[0][178] ), .A2(\RI5[0][22] ), .Z(
        \MC_ARK_ARC_1_0/temp3[112] ) );
  NAND3_X2 U9886 ( .A1(\SB2_2_8/i0_0 ), .A2(\SB2_2_8/i0_3 ), .A3(
        \SB2_2_8/i0_4 ), .ZN(n4038) );
  XOR2_X1 U9893 ( .A1(n4044), .A2(n4043), .Z(\MC_ARK_ARC_1_1/buf_output[165] )
         );
  NAND3_X1 U9895 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB1_1_27/buf_output[0] ), .A3(
        n6283), .ZN(\SB2_1_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U9896 ( .A1(\RI3[0][190] ), .A2(\SB2_0_0/i1_7 ), .A3(n4003), .ZN(
        \SB2_0_0/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U9899 ( .A1(n1890), .A2(n4046), .Z(n1544) );
  XOR2_X1 U9900 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[53] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[5] ), .Z(n4046) );
  XOR2_X1 U9901 ( .A1(\RI5[2][167] ), .A2(\RI5[2][101] ), .Z(n5085) );
  XOR2_X1 U9903 ( .A1(n1018), .A2(n4047), .Z(n2083) );
  XOR2_X1 U9906 ( .A1(\RI5[2][189] ), .A2(\RI5[2][21] ), .Z(n4048) );
  NAND3_X2 U9907 ( .A1(\SB2_3_1/i0[9] ), .A2(\SB2_3_1/i0[6] ), .A3(
        \SB2_3_1/i0_4 ), .ZN(n2115) );
  NAND3_X2 U9909 ( .A1(\SB1_0_15/i0[6] ), .A2(\SB1_0_15/i0[10] ), .A3(
        \SB1_0_15/i0_3 ), .ZN(n4049) );
  NAND3_X1 U9912 ( .A1(\SB1_2_29/i0[8] ), .A2(\RI1[2][17] ), .A3(
        \SB1_2_29/i1_7 ), .ZN(\SB1_2_29/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U9913 ( .A1(\SB1_4_6/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_4_6/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_4_6/Component_Function_5/NAND4_in[0] ), .A4(n2997), .ZN(
        \SB1_4_6/buf_output[5] ) );
  NAND4_X2 U9914 ( .A1(\SB3_8/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_8/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_8/buf_output[1] )
         );
  NAND4_X2 U9916 ( .A1(\SB1_2_3/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_2_3/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_3/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_2_3/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_2_3/buf_output[4] ) );
  XOR2_X1 U9917 ( .A1(\RI5[3][113] ), .A2(\RI5[3][77] ), .Z(
        \MC_ARK_ARC_1_3/temp3[11] ) );
  XOR2_X1 U9920 ( .A1(\MC_ARK_ARC_1_4/temp2[170] ), .A2(n4052), .Z(
        \MC_ARK_ARC_1_4/temp5[170] ) );
  XOR2_X1 U9921 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[170] ), .A2(\RI5[4][164] ), 
        .Z(n4052) );
  NAND4_X2 U9922 ( .A1(\SB2_4_6/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_6/Component_Function_0/NAND4_in[1] ), .A3(n1823), .A4(
        \SB2_4_6/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_4_6/buf_output[0] ) );
  NAND4_X2 U9923 ( .A1(\SB1_4_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_4_11/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_4_11/Component_Function_2/NAND4_in[1] ), .A4(n4053), .ZN(
        \SB1_4_11/buf_output[2] ) );
  XOR2_X1 U9927 ( .A1(n4056), .A2(\MC_ARK_ARC_1_1/temp2[148] ), .Z(n1390) );
  XOR2_X1 U9930 ( .A1(\MC_ARK_ARC_1_4/temp5[124] ), .A2(
        \MC_ARK_ARC_1_4/temp6[124] ), .Z(\MC_ARK_ARC_1_4/buf_output[124] ) );
  NAND3_X1 U9933 ( .A1(\SB2_4_27/i0[9] ), .A2(\SB2_4_27/i0[6] ), .A3(
        \SB2_4_27/i1_5 ), .ZN(\SB2_4_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U9936 ( .A1(\SB3_18/i0[6] ), .A2(\SB3_18/i0[8] ), .A3(
        \SB3_18/i0[7] ), .ZN(\SB3_18/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U9937 ( .A1(\MC_ARK_ARC_1_3/temp4[154] ), .A2(
        \MC_ARK_ARC_1_3/temp3[154] ), .Z(n4060) );
  NAND4_X2 U9938 ( .A1(n2231), .A2(\SB2_3_18/Component_Function_3/NAND4_in[0] ), .A3(\SB2_3_18/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_3_18/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_18/buf_output[3] ) );
  NAND3_X1 U9939 ( .A1(\SB4_4/i0_3 ), .A2(\SB4_4/i0[8] ), .A3(\SB4_4/i1_7 ), 
        .ZN(\SB4_4/Component_Function_1/NAND4_in[1] ) );
  INV_X2 U9942 ( .I(\SB1_3_10/buf_output[2] ), .ZN(\SB2_3_7/i1[9] ) );
  NAND4_X2 U9943 ( .A1(\SB1_3_10/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_3_10/Component_Function_2/NAND4_in[0] ), .A3(n4855), .A4(
        \SB1_3_10/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB1_3_10/buf_output[2] ) );
  NAND4_X2 U9945 ( .A1(n5340), .A2(n5339), .A3(
        \SB2_2_25/Component_Function_0/NAND4_in[0] ), .A4(n4063), .ZN(
        \SB2_2_25/buf_output[0] ) );
  INV_X2 U9948 ( .I(\SB1_4_16/buf_output[3] ), .ZN(\SB2_4_14/i0[8] ) );
  NAND4_X2 U9950 ( .A1(n4298), .A2(\SB2_2_19/Component_Function_5/NAND4_in[0] ), .A3(\SB2_2_19/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_19/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_2_19/buf_output[5] ) );
  NAND4_X2 U9952 ( .A1(\SB2_1_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_7/Component_Function_2/NAND4_in[2] ), .A3(n4065), .A4(
        \SB2_1_7/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_1_7/buf_output[2] ) );
  NAND4_X2 U9954 ( .A1(\SB1_1_9/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_9/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_9/Component_Function_4/NAND4_in[2] ), .A4(n4066), .ZN(
        \SB1_1_9/buf_output[4] ) );
  NAND3_X1 U9955 ( .A1(\SB1_1_9/i0_4 ), .A2(\SB1_1_9/i1[9] ), .A3(
        \SB1_1_9/i1_5 ), .ZN(n4066) );
  INV_X2 U9956 ( .I(\SB1_3_19/buf_output[3] ), .ZN(\SB2_3_17/i0[8] ) );
  NAND4_X2 U9959 ( .A1(\SB1_1_16/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_16/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_16/Component_Function_4/NAND4_in[3] ), .A4(n4068), .ZN(
        \SB1_1_16/buf_output[4] ) );
  NAND4_X2 U9960 ( .A1(\SB2_2_0/Component_Function_5/NAND4_in[2] ), .A2(n601), 
        .A3(n5406), .A4(n4069), .ZN(\SB2_2_0/buf_output[5] ) );
  NAND3_X1 U9961 ( .A1(n5444), .A2(\SB1_2_5/buf_output[0] ), .A3(
        \SB1_2_4/buf_output[1] ), .ZN(n4069) );
  XOR2_X1 U9962 ( .A1(\MC_ARK_ARC_1_1/temp6[86] ), .A2(n4070), .Z(
        \MC_ARK_ARC_1_1/buf_output[86] ) );
  XOR2_X1 U9964 ( .A1(\MC_ARK_ARC_1_1/temp3[183] ), .A2(
        \MC_ARK_ARC_1_1/temp4[183] ), .Z(\MC_ARK_ARC_1_1/temp6[183] ) );
  NAND3_X1 U9966 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0_0 ), .A3(
        \SB2_0_5/i0_4 ), .ZN(\SB2_0_5/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U9967 ( .A1(\MC_ARK_ARC_1_0/temp3[162] ), .A2(
        \MC_ARK_ARC_1_0/temp4[162] ), .Z(\MC_ARK_ARC_1_0/temp6[162] ) );
  XOR2_X1 U9968 ( .A1(\SB2_3_10/buf_output[4] ), .A2(\RI5[3][160] ), .Z(
        \MC_ARK_ARC_1_3/temp2[190] ) );
  XOR2_X1 U9970 ( .A1(\MC_ARK_ARC_1_2/temp5[45] ), .A2(n4073), .Z(
        \MC_ARK_ARC_1_2/buf_output[45] ) );
  XOR2_X1 U9971 ( .A1(\MC_ARK_ARC_1_2/temp3[45] ), .A2(
        \MC_ARK_ARC_1_2/temp4[45] ), .Z(n4073) );
  NAND4_X2 U9972 ( .A1(\SB2_1_20/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_20/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_20/Component_Function_1/NAND4_in[2] ), .A4(n4074), .ZN(
        \SB2_1_20/buf_output[1] ) );
  XOR2_X1 U9974 ( .A1(\RI5[1][113] ), .A2(\RI5[1][107] ), .Z(n4075) );
  NAND4_X2 U9977 ( .A1(\SB1_4_15/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_4_15/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_4_15/Component_Function_4/NAND4_in[1] ), .A4(n4350), .ZN(
        \SB1_4_15/buf_output[4] ) );
  NOR2_X2 U9984 ( .A1(n4610), .A2(n4130), .ZN(n4081) );
  XOR2_X1 U9985 ( .A1(n4082), .A2(\MC_ARK_ARC_1_0/temp6[126] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[126] ) );
  XOR2_X1 U9986 ( .A1(\MC_ARK_ARC_1_0/temp1[126] ), .A2(
        \MC_ARK_ARC_1_0/temp2[126] ), .Z(n4082) );
  XOR2_X1 U9987 ( .A1(\RI5[2][59] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[35] ), 
        .Z(n1739) );
  INV_X8 U9988 ( .I(n4083), .ZN(\RI1[2][17] ) );
  INV_X2 U9989 ( .I(\MC_ARK_ARC_1_1/buf_output[17] ), .ZN(n4083) );
  NAND4_X2 U9992 ( .A1(\SB2_0_13/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_0_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_0/NAND4_in[0] ), .A4(n4084), .ZN(
        \SB2_0_13/buf_output[0] ) );
  NAND3_X2 U9993 ( .A1(\SB2_0_13/i0_0 ), .A2(\SB2_0_13/i0_3 ), .A3(
        \SB2_0_13/i0[7] ), .ZN(n4084) );
  NAND4_X2 U9994 ( .A1(\SB1_4_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_20/Component_Function_3/NAND4_in[1] ), .A3(n1793), .A4(
        \SB1_4_20/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_4_20/buf_output[3] ) );
  NOR2_X2 U9998 ( .A1(n4089), .A2(n4087), .ZN(n630) );
  NAND2_X2 U9999 ( .A1(\SB1_0_9/Component_Function_0/NAND4_in[1] ), .A2(n4088), 
        .ZN(n4087) );
  NAND4_X2 U10002 ( .A1(\SB2_0_3/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_3/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_3/Component_Function_4/NAND4_in[1] ), .A4(n4090), .ZN(
        \SB2_0_3/buf_output[4] ) );
  NAND4_X2 U10006 ( .A1(\SB2_1_15/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_15/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_15/Component_Function_1/NAND4_in[2] ), .A4(n4093), .ZN(
        \SB2_1_15/buf_output[1] ) );
  NAND3_X2 U10007 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0[9] ), .A3(
        \SB1_1_22/i0[8] ), .ZN(\SB1_1_22/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U10008 ( .I(\SB1_4_31/buf_output[2] ), .ZN(\SB2_4_28/i1[9] ) );
  NAND4_X2 U10009 ( .A1(\SB1_4_31/Component_Function_2/NAND4_in[1] ), .A2(
        n5155), .A3(\SB1_4_31/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_4_31/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_4_31/buf_output[2] ) );
  NAND3_X2 U10020 ( .A1(\SB1_3_28/i0_3 ), .A2(\SB1_3_28/i0_4 ), .A3(
        \SB1_3_28/i1[9] ), .ZN(\SB1_3_28/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U10022 ( .A1(\SB3_15/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_15/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_15/Component_Function_4/NAND4_in[3] ), .A4(n4098), .ZN(
        \SB3_15/buf_output[4] ) );
  NAND3_X1 U10023 ( .A1(\SB3_15/i0_0 ), .A2(\SB3_15/i3[0] ), .A3(\SB3_15/i1_7 ), .ZN(n4098) );
  INV_X4 U10024 ( .I(\SB2_0_4/i0[7] ), .ZN(\RI3[0][166] ) );
  NAND2_X1 U10026 ( .A1(n4101), .A2(\SB1_0_5/Component_Function_4/NAND4_in[1] ), .ZN(n4099) );
  NAND3_X1 U10028 ( .A1(\SB1_0_5/i0_3 ), .A2(\SB1_0_5/i0[9] ), .A3(
        \SB1_0_5/i0[10] ), .ZN(n4101) );
  NOR2_X2 U10029 ( .A1(n2802), .A2(n4102), .ZN(n3000) );
  NAND3_X2 U10030 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i1[9] ), .A3(
        \SB1_1_22/i0[6] ), .ZN(\SB1_1_22/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U10031 ( .A1(\SB2_2_16/Component_Function_1/NAND4_in[3] ), .A2(
        n5374), .A3(\SB2_2_16/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_2_16/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_2_16/buf_output[1] ) );
  NAND3_X1 U10033 ( .A1(\SB2_0_14/i0[10] ), .A2(\SB2_0_14/i1_5 ), .A3(
        \SB2_0_14/i1[9] ), .ZN(\SB2_0_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U10034 ( .A1(n2381), .A2(\SB2_0_5/i0_3 ), .A3(\SB2_0_5/i0_0 ), .ZN(
        n4724) );
  XOR2_X1 U10035 ( .A1(\MC_ARK_ARC_1_4/temp5[98] ), .A2(
        \MC_ARK_ARC_1_4/temp6[98] ), .Z(\MC_ARK_ARC_1_4/buf_output[98] ) );
  NAND3_X2 U10036 ( .A1(\SB2_1_21/i0_4 ), .A2(\SB2_1_21/i0[9] ), .A3(
        \SB2_1_21/i0[6] ), .ZN(\SB2_1_21/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U10037 ( .A1(\MC_ARK_ARC_1_2/temp1[121] ), .A2(n2136), .Z(n5161) );
  XOR2_X1 U10038 ( .A1(\MC_ARK_ARC_1_0/temp1[186] ), .A2(
        \MC_ARK_ARC_1_0/temp2[186] ), .Z(n1653) );
  NAND3_X2 U10041 ( .A1(\SB2_1_19/i0_0 ), .A2(\SB2_1_19/i1_5 ), .A3(
        \SB2_1_19/i0_4 ), .ZN(n2733) );
  XOR2_X1 U10043 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[80] ), .A2(\RI5[3][56] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[110] ) );
  NAND4_X2 U10044 ( .A1(\SB2_2_20/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_2_20/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_20/Component_Function_3/NAND4_in[1] ), .A4(n4104), .ZN(
        \SB2_2_20/buf_output[3] ) );
  XOR2_X1 U10045 ( .A1(n1764), .A2(n4105), .Z(\MC_ARK_ARC_1_4/buf_output[62] )
         );
  XOR2_X1 U10046 ( .A1(\MC_ARK_ARC_1_4/temp4[62] ), .A2(n4316), .Z(n4105) );
  XOR2_X1 U10048 ( .A1(\MC_ARK_ARC_1_3/temp4[185] ), .A2(n4107), .Z(n4343) );
  XOR2_X1 U10049 ( .A1(\RI5[3][59] ), .A2(\RI5[3][95] ), .Z(n4107) );
  NAND3_X1 U10052 ( .A1(\SB2_1_22/i0_4 ), .A2(\SB2_1_22/i1[9] ), .A3(
        \SB2_1_22/i1_5 ), .ZN(\SB2_1_22/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U10053 ( .A1(\MC_ARK_ARC_1_3/temp5[100] ), .A2(n4109), .Z(
        \MC_ARK_ARC_1_3/buf_output[100] ) );
  XOR2_X1 U10054 ( .A1(\MC_ARK_ARC_1_3/temp4[100] ), .A2(n599), .Z(n4109) );
  XOR2_X1 U10058 ( .A1(\MC_ARK_ARC_1_4/temp3[191] ), .A2(
        \MC_ARK_ARC_1_4/temp4[191] ), .Z(n4113) );
  INV_X2 U10059 ( .I(\RI3[4][188] ), .ZN(\SB2_4_0/i1[9] ) );
  NAND4_X2 U10061 ( .A1(\SB1_1_16/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_16/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_1_16/Component_Function_1/NAND4_in[2] ), .A4(n4114), .ZN(
        \SB1_1_16/buf_output[1] ) );
  XOR2_X1 U10062 ( .A1(\MC_ARK_ARC_1_3/temp6[171] ), .A2(n4115), .Z(
        \MC_ARK_ARC_1_3/buf_output[171] ) );
  XOR2_X1 U10063 ( .A1(n4739), .A2(\MC_ARK_ARC_1_3/temp2[171] ), .Z(n4115) );
  NAND3_X2 U10064 ( .A1(\SB1_3_31/i0[10] ), .A2(\SB1_3_31/i1[9] ), .A3(
        \SB1_3_31/i1_5 ), .ZN(n4329) );
  NAND4_X2 U10067 ( .A1(n2121), .A2(
        \SB1_4_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_4_15/Component_Function_3/NAND4_in[2] ), .A4(n5086), .ZN(
        \SB1_4_15/buf_output[3] ) );
  NAND4_X2 U10069 ( .A1(\SB2_3_2/Component_Function_5/NAND4_in[3] ), .A2(n4768), .A3(n4143), .A4(\SB2_3_2/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_2/buf_output[5] ) );
  XOR2_X1 U10074 ( .A1(n4118), .A2(n4117), .Z(n3093) );
  XOR2_X1 U10075 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[99] ), .A2(n165), .Z(
        n4117) );
  XOR2_X1 U10079 ( .A1(\MC_ARK_ARC_1_2/temp3[23] ), .A2(
        \MC_ARK_ARC_1_2/temp2[23] ), .Z(n4120) );
  XOR2_X1 U10082 ( .A1(\MC_ARK_ARC_1_0/temp5[96] ), .A2(n4122), .Z(
        \MC_ARK_ARC_1_0/buf_output[96] ) );
  XOR2_X1 U10083 ( .A1(\MC_ARK_ARC_1_0/temp3[96] ), .A2(
        \MC_ARK_ARC_1_0/temp4[96] ), .Z(n4122) );
  XOR2_X1 U10084 ( .A1(n4124), .A2(n4123), .Z(\MC_ARK_ARC_1_2/buf_output[155] ) );
  XOR2_X1 U10087 ( .A1(n4126), .A2(\MC_ARK_ARC_1_0/temp4[152] ), .Z(n2343) );
  XOR2_X1 U10088 ( .A1(\RI5[0][26] ), .A2(\RI5[0][62] ), .Z(n4126) );
  INV_X2 U10094 ( .I(\SB1_4_6/buf_output[3] ), .ZN(\SB2_4_4/i0[8] ) );
  NAND3_X1 U10096 ( .A1(\SB1_4_18/i0_3 ), .A2(\SB1_4_18/i0_0 ), .A3(
        \SB1_4_18/i0_4 ), .ZN(\SB1_4_18/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U10098 ( .A1(\RI5[4][32] ), .A2(\RI5[4][8] ), .Z(n1339) );
  NAND3_X2 U10101 ( .A1(\SB1_2_30/i0[10] ), .A2(\SB1_2_30/i1[9] ), .A3(
        \SB1_2_30/i1_5 ), .ZN(n4129) );
  INV_X1 U10103 ( .I(\RI3[0][29] ), .ZN(\SB2_0_27/i1_5 ) );
  NAND4_X2 U10104 ( .A1(\SB1_0_27/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_0_27/Component_Function_5/NAND4_in[2] ), .A3(n4839), .A4(
        \SB1_0_27/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][29] ) );
  INV_X1 U10109 ( .I(\RI3[0][47] ), .ZN(\SB2_0_24/i1_5 ) );
  NAND4_X2 U10110 ( .A1(\SB1_0_24/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_24/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_0_24/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_24/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][47] ) );
  NAND4_X2 U10111 ( .A1(\SB2_0_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_12/Component_Function_4/NAND4_in[2] ), .A4(n4133), .ZN(
        \SB2_0_12/buf_output[4] ) );
  NAND3_X2 U10112 ( .A1(\SB2_0_12/i1_5 ), .A2(\SB2_0_12/i1[9] ), .A3(
        \RI3[0][118] ), .ZN(n4133) );
  NAND3_X2 U10114 ( .A1(\SB2_2_3/i0[10] ), .A2(n3994), .A3(\SB2_2_3/i1[9] ), 
        .ZN(n4135) );
  XOR2_X1 U10115 ( .A1(n4136), .A2(\MC_ARK_ARC_1_1/temp4[26] ), .Z(n4474) );
  XOR2_X1 U10116 ( .A1(\RI5[1][128] ), .A2(\RI5[1][92] ), .Z(n4136) );
  NAND2_X2 U10118 ( .A1(\SB1_0_24/i0[9] ), .A2(\SB1_0_24/i0[10] ), .ZN(n4138)
         );
  XOR2_X1 U10119 ( .A1(\MC_ARK_ARC_1_3/temp2[71] ), .A2(n4139), .Z(
        \MC_ARK_ARC_1_3/temp5[71] ) );
  XOR2_X1 U10120 ( .A1(\RI5[3][65] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .Z(n4139) );
  XOR2_X1 U10121 ( .A1(\RI5[1][139] ), .A2(\RI5[1][175] ), .Z(n4140) );
  NAND4_X2 U10122 ( .A1(\SB2_4_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_19/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_4_19/Component_Function_4/NAND4_in[1] ), .A4(n4141), .ZN(
        \SB2_4_19/buf_output[4] ) );
  XOR2_X1 U10124 ( .A1(\RI5[1][128] ), .A2(\RI5[1][104] ), .Z(n4142) );
  NAND3_X2 U10125 ( .A1(\SB2_3_2/i0[6] ), .A2(\SB2_3_2/i0[10] ), .A3(
        \SB2_3_2/i0_0 ), .ZN(n4143) );
  NAND4_X2 U10126 ( .A1(\SB1_0_24/Component_Function_2/NAND4_in[1] ), .A2(
        n5381), .A3(n5023), .A4(n4144), .ZN(\SB1_0_24/buf_output[2] ) );
  NAND3_X2 U10127 ( .A1(\SB1_0_24/i0[9] ), .A2(\SB1_0_24/i0[8] ), .A3(
        \SB1_0_24/i0_3 ), .ZN(n4144) );
  NAND3_X2 U10129 ( .A1(\SB1_0_19/i0_0 ), .A2(\SB1_0_19/i1_5 ), .A3(
        \SB1_0_19/i0_4 ), .ZN(n4146) );
  NAND3_X2 U10130 ( .A1(\SB1_4_25/i0_3 ), .A2(\SB1_4_25/i1[9] ), .A3(
        \SB1_4_25/i0[6] ), .ZN(n4147) );
  NAND4_X1 U10135 ( .A1(\SB2_0_27/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_27/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_27/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_0_27/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB2_0_27/buf_output[3] ) );
  XOR2_X1 U10138 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[23] ), .A2(\RI5[4][59] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[149] ) );
  NAND4_X2 U10140 ( .A1(\SB1_2_18/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_18/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_2_18/Component_Function_5/NAND4_in[0] ), .A4(n4149), .ZN(
        \SB1_2_18/buf_output[5] ) );
  NAND3_X2 U10141 ( .A1(\SB2_0_17/i0[6] ), .A2(\SB2_0_17/i0[10] ), .A3(
        \SB2_0_17/i0_0 ), .ZN(\SB2_0_17/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U10142 ( .A1(n1284), .A2(n5319), .Z(\MC_ARK_ARC_1_2/buf_output[57] )
         );
  NAND4_X2 U10143 ( .A1(\SB1_3_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_2/Component_Function_1/NAND4_in[2] ), .A3(n4756), .A4(
        \SB1_3_2/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_2/buf_output[1] ) );
  XOR2_X1 U10145 ( .A1(\MC_ARK_ARC_1_2/temp5[68] ), .A2(n1089), .Z(
        \MC_ARK_ARC_1_2/buf_output[68] ) );
  XOR2_X1 U10146 ( .A1(\RI5[1][95] ), .A2(\RI5[1][59] ), .Z(
        \MC_ARK_ARC_1_1/temp3[185] ) );
  XOR2_X1 U10147 ( .A1(\RI5[1][23] ), .A2(\RI5[1][29] ), .Z(n745) );
  XOR2_X1 U10149 ( .A1(\RI5[1][95] ), .A2(\RI5[1][131] ), .Z(n1856) );
  XOR2_X1 U10152 ( .A1(n4150), .A2(\MC_ARK_ARC_1_1/temp6[98] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[98] ) );
  NAND4_X2 U10154 ( .A1(\SB2_3_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_17/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_3_17/Component_Function_2/NAND4_in[1] ), .A4(n4151), .ZN(
        \SB2_3_17/buf_output[2] ) );
  XOR2_X1 U10156 ( .A1(\RI5[3][104] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[140] ), .Z(n4189) );
  NAND3_X1 U10157 ( .A1(\SB1_2_22/i0[8] ), .A2(\SB1_2_22/i1_7 ), .A3(
        \RI1[2][59] ), .ZN(\SB1_2_22/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U10158 ( .A1(\SB1_1_0/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_0/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_0/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_1_0/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_0/buf_output[1] ) );
  NAND4_X2 U10159 ( .A1(\SB2_3_6/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_3_6/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_6/Component_Function_3/NAND4_in[1] ), .A4(n4152), .ZN(
        \SB2_3_6/buf_output[3] ) );
  NAND3_X2 U10160 ( .A1(\SB2_3_6/i0[10] ), .A2(\SB2_3_6/i1[9] ), .A3(
        \SB2_3_6/i1_7 ), .ZN(n4152) );
  NAND3_X2 U10162 ( .A1(\SB2_4_29/i0[8] ), .A2(\SB2_4_29/i3[0] ), .A3(
        \SB2_4_29/i1_5 ), .ZN(n4153) );
  XOR2_X1 U10163 ( .A1(n4154), .A2(\MC_ARK_ARC_1_3/temp1[3] ), .Z(n2253) );
  XOR2_X1 U10164 ( .A1(\RI5[3][165] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[141] ), .Z(n4154) );
  XOR2_X1 U10165 ( .A1(\SB2_3_20/buf_output[3] ), .A2(n174), .Z(n4155) );
  NAND3_X2 U10170 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0_0 ), .A3(
        \SB2_1_9/i0_4 ), .ZN(\SB2_1_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U10171 ( .A1(\SB1_2_24/i0_3 ), .A2(\SB1_2_24/i0[8] ), .A3(
        \SB1_2_24/i1_7 ), .ZN(\SB1_2_24/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U10172 ( .A1(\MC_ARK_ARC_1_1/temp1[153] ), .A2(
        \MC_ARK_ARC_1_1/temp2[153] ), .Z(n4556) );
  XOR2_X1 U10177 ( .A1(\RI5[2][87] ), .A2(\RI5[2][51] ), .Z(
        \MC_ARK_ARC_1_2/temp3[177] ) );
  XOR2_X1 U10179 ( .A1(\MC_ARK_ARC_1_0/temp4[92] ), .A2(n1305), .Z(n4160) );
  XOR2_X1 U10180 ( .A1(\MC_ARK_ARC_1_3/temp2[112] ), .A2(n4161), .Z(
        \MC_ARK_ARC_1_3/temp5[112] ) );
  XOR2_X1 U10181 ( .A1(\RI5[3][106] ), .A2(\RI5[3][112] ), .Z(n4161) );
  XOR2_X1 U10182 ( .A1(\MC_ARK_ARC_1_2/temp3[137] ), .A2(n4162), .Z(n2360) );
  XOR2_X1 U10183 ( .A1(\RI5[2][83] ), .A2(\RI5[2][107] ), .Z(n4162) );
  XOR2_X1 U10189 ( .A1(\MC_ARK_ARC_1_1/temp6[157] ), .A2(n4165), .Z(
        \MC_ARK_ARC_1_1/buf_output[157] ) );
  NAND3_X2 U10194 ( .A1(\SB2_0_31/i0[10] ), .A2(\SB2_0_31/i1[9] ), .A3(
        \SB2_0_31/i1_5 ), .ZN(\SB2_0_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U10201 ( .A1(\SB2_0_24/i0_3 ), .A2(\SB2_0_24/i1[9] ), .A3(
        \RI3[0][46] ), .ZN(n4169) );
  XOR2_X1 U10202 ( .A1(n4171), .A2(n4170), .Z(\MC_ARK_ARC_1_0/buf_output[94] )
         );
  XOR2_X1 U10203 ( .A1(\MC_ARK_ARC_1_0/temp2[94] ), .A2(
        \MC_ARK_ARC_1_0/temp4[94] ), .Z(n4170) );
  XOR2_X1 U10204 ( .A1(\MC_ARK_ARC_1_0/temp3[94] ), .A2(
        \MC_ARK_ARC_1_0/temp1[94] ), .Z(n4171) );
  XOR2_X1 U10205 ( .A1(\MC_ARK_ARC_1_3/temp5[39] ), .A2(n4172), .Z(
        \MC_ARK_ARC_1_3/buf_output[39] ) );
  XOR2_X1 U10206 ( .A1(\MC_ARK_ARC_1_3/temp3[39] ), .A2(
        \MC_ARK_ARC_1_3/temp4[39] ), .Z(n4172) );
  NAND3_X2 U10207 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0[9] ), .A3(
        \SB2_3_17/i0[8] ), .ZN(\SB2_3_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U10210 ( .A1(\SB2_2_18/i0[6] ), .A2(\SB2_2_18/i0_3 ), .A3(
        \SB2_2_18/i0[10] ), .ZN(n4174) );
  XOR2_X1 U10214 ( .A1(\MC_ARK_ARC_1_2/temp5[5] ), .A2(
        \MC_ARK_ARC_1_2/temp6[5] ), .Z(\RI1[3][5] ) );
  XOR2_X1 U10220 ( .A1(\RI5[3][149] ), .A2(\RI5[3][173] ), .Z(n4177) );
  NAND4_X2 U10221 ( .A1(\SB1_2_22/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_22/Component_Function_0/NAND4_in[2] ), .A3(n1636), .A4(n4176), 
        .ZN(\SB1_2_22/buf_output[0] ) );
  XOR2_X1 U10222 ( .A1(n4177), .A2(n4178), .Z(n2950) );
  XOR2_X1 U10223 ( .A1(\RI5[3][11] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[5] ), 
        .Z(n4178) );
  XOR2_X1 U10225 ( .A1(n5074), .A2(n4430), .Z(\MC_ARK_ARC_1_1/temp5[171] ) );
  XOR2_X1 U10227 ( .A1(n4183), .A2(n4182), .Z(\MC_ARK_ARC_1_0/temp5[153] ) );
  XOR2_X1 U10231 ( .A1(n4185), .A2(n4184), .Z(\MC_ARK_ARC_1_0/temp6[26] ) );
  XOR2_X1 U10232 ( .A1(\SB2_0_19/buf_output[2] ), .A2(n11), .Z(n4184) );
  XOR2_X1 U10233 ( .A1(\RI5[0][128] ), .A2(\RI5[0][62] ), .Z(n4185) );
  NAND3_X1 U10234 ( .A1(\SB1_2_29/i0_0 ), .A2(\SB1_2_29/i1_7 ), .A3(
        \SB1_2_29/i3[0] ), .ZN(\SB1_2_29/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U10235 ( .A1(\SB3_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_3/NAND4_in[1] ), .A3(n4989), .A4(n4856), 
        .ZN(\SB3_21/buf_output[3] ) );
  NAND4_X2 U10236 ( .A1(\SB2_2_28/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_28/Component_Function_5/NAND4_in[1] ), .A3(n5043), .A4(
        \SB2_2_28/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_28/buf_output[5] ) );
  XOR2_X1 U10237 ( .A1(\RI5[4][178] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[22] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[112] ) );
  NAND3_X2 U10241 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i0[10] ), .A3(
        \SB2_0_11/i0[6] ), .ZN(n5052) );
  NAND4_X2 U10242 ( .A1(\SB1_4_15/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_4_15/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_4_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_15/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_4_15/buf_output[0] ) );
  NAND3_X2 U10243 ( .A1(\SB2_1_30/i0[6] ), .A2(\SB2_1_30/i1[9] ), .A3(
        \SB2_1_30/i0_3 ), .ZN(\SB2_1_30/Component_Function_3/NAND4_in[0] ) );
  AND2_X1 U10245 ( .A1(n340), .A2(n392), .Z(n4187) );
  NAND4_X2 U10246 ( .A1(n1166), .A2(
        \SB1_0_14/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_2/NAND4_in[0] ), .A4(n4917), .ZN(
        \RI3[0][122] ) );
  XOR2_X1 U10248 ( .A1(n4188), .A2(\MC_ARK_ARC_1_3/temp2[141] ), .Z(n4865) );
  XOR2_X1 U10249 ( .A1(\RI5[3][135] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[141] ), .Z(n4188) );
  NAND3_X2 U10251 ( .A1(\SB2_3_7/i0[6] ), .A2(\SB2_3_7/i0_4 ), .A3(
        \SB2_3_7/i0[9] ), .ZN(n4287) );
  XOR2_X1 U10254 ( .A1(\MC_ARK_ARC_1_4/temp6[146] ), .A2(n4191), .Z(
        \MC_ARK_ARC_1_4/buf_output[146] ) );
  NAND3_X2 U10261 ( .A1(\SB2_2_10/i0[10] ), .A2(n589), .A3(\SB2_2_10/i1[9] ), 
        .ZN(n4192) );
  NAND3_X2 U10263 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i0[10] ), .A3(
        \SB2_0_11/i0[9] ), .ZN(n4193) );
  XOR2_X1 U10264 ( .A1(\RI5[0][14] ), .A2(\RI5[0][20] ), .Z(n2601) );
  NAND3_X1 U10265 ( .A1(\SB1_0_16/i0_0 ), .A2(\SB1_0_16/i0_3 ), .A3(
        \SB1_0_16/i0[7] ), .ZN(\SB1_0_16/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U10266 ( .A1(\MC_ARK_ARC_1_4/temp2[182] ), .A2(
        \MC_ARK_ARC_1_4/temp1[182] ), .Z(n4194) );
  XOR2_X1 U10267 ( .A1(\RI5[0][185] ), .A2(\RI5[0][161] ), .Z(n3078) );
  XOR2_X1 U10271 ( .A1(\RI5[4][65] ), .A2(\RI5[4][131] ), .Z(n4197) );
  NAND4_X2 U10272 ( .A1(\SB2_0_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_4/Component_Function_3/NAND4_in[2] ), .A3(n1669), .A4(n4198), 
        .ZN(\SB2_0_4/buf_output[3] ) );
  NAND4_X2 U10273 ( .A1(\SB2_0_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_31/Component_Function_3/NAND4_in[2] ), .A3(n5066), .A4(
        \SB2_0_31/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_31/buf_output[3] ) );
  NAND3_X2 U10275 ( .A1(\SB1_1_23/i0[8] ), .A2(\SB1_1_23/i3[0] ), .A3(
        \SB1_1_23/i1_5 ), .ZN(n4199) );
  XOR2_X1 U10277 ( .A1(n5185), .A2(n4201), .Z(\MC_ARK_ARC_1_2/buf_output[186] ) );
  XOR2_X1 U10278 ( .A1(\MC_ARK_ARC_1_2/temp2[186] ), .A2(n4330), .Z(n4201) );
  XOR2_X1 U10280 ( .A1(\MC_ARK_ARC_1_0/temp4[153] ), .A2(
        \MC_ARK_ARC_1_0/temp3[153] ), .Z(n4202) );
  NAND4_X2 U10281 ( .A1(\SB2_2_6/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_6/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_2_6/Component_Function_0/NAND4_in[3] ), .A4(n4203), .ZN(
        \SB2_2_6/buf_output[0] ) );
  INV_X1 U10283 ( .I(\SB1_0_2/buf_output[0] ), .ZN(\SB2_0_29/i3[0] ) );
  NAND4_X2 U10284 ( .A1(\SB1_0_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_2/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_2/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_0_2/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_0_2/buf_output[0] ) );
  NAND3_X1 U10285 ( .A1(\SB1_1_1/i0[6] ), .A2(\SB1_1_1/i0[9] ), .A3(
        \SB1_1_1/i0_4 ), .ZN(\SB1_1_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U10286 ( .A1(\SB2_0_26/i0[8] ), .A2(\SB2_0_26/i3[0] ), .A3(
        \SB2_0_26/i1_5 ), .ZN(\SB2_0_26/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U10292 ( .A1(\RI5[0][150] ), .A2(\RI5[0][174] ), .Z(n4207) );
  XOR2_X1 U10293 ( .A1(\MC_ARK_ARC_1_3/temp2[76] ), .A2(
        \MC_ARK_ARC_1_3/temp1[76] ), .Z(\MC_ARK_ARC_1_3/temp5[76] ) );
  NAND3_X2 U10300 ( .A1(\SB1_4_29/i0[10] ), .A2(\SB1_4_29/i0_0 ), .A3(
        \SB1_4_29/i0[6] ), .ZN(n4213) );
  NAND3_X2 U10301 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i1[9] ), .A3(
        \SB1_1_14/i0_4 ), .ZN(\SB1_1_14/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U10302 ( .A1(\SB1_2_6/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_0/NAND4_in[0] ), .A4(n4214), .ZN(
        \SB1_2_6/buf_output[0] ) );
  NAND3_X1 U10304 ( .A1(\SB4_4/i0[10] ), .A2(\SB4_4/i0[9] ), .A3(\SB4_4/i0_3 ), 
        .ZN(\SB4_4/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U10310 ( .A1(\SB3_3/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_3/Component_Function_5/NAND4_in[3] ), .A3(n2498), .A4(
        \SB3_3/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_3/buf_output[5] )
         );
  NAND4_X2 U10311 ( .A1(\SB2_2_3/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_3/Component_Function_4/NAND4_in[3] ), .A3(n5208), .A4(
        \SB2_2_3/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB2_2_3/buf_output[4] ) );
  XOR2_X1 U10313 ( .A1(\RI5[3][26] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[182] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[116] ) );
  NAND3_X2 U10314 ( .A1(\SB2_2_1/i0[10] ), .A2(\SB2_2_1/i0_0 ), .A3(
        \SB2_2_1/i0[6] ), .ZN(\SB2_2_1/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U10315 ( .A1(\RI5[2][178] ), .A2(\RI5[2][184] ), .Z(
        \MC_ARK_ARC_1_2/temp1[184] ) );
  NAND4_X2 U10316 ( .A1(\SB1_4_22/Component_Function_4/NAND4_in[3] ), .A2(
        n1538), .A3(\SB1_4_22/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_4_22/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB1_4_22/buf_output[4] ) );
  NAND3_X1 U10317 ( .A1(\SB2_3_30/i0_3 ), .A2(\SB2_3_30/i0_0 ), .A3(
        \SB2_3_30/i0[7] ), .ZN(n1613) );
  NAND3_X1 U10322 ( .A1(\SB1_2_0/i0_0 ), .A2(\SB1_2_0/i3[0] ), .A3(
        \SB1_2_0/i1_7 ), .ZN(\SB1_2_0/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U10324 ( .A1(\MC_ARK_ARC_1_1/temp4[188] ), .A2(n5097), .Z(n4219) );
  NAND4_X2 U10327 ( .A1(\SB1_0_14/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_4/NAND4_in[0] ), .A4(n4221), .ZN(
        \SB1_0_14/buf_output[4] ) );
  NAND3_X1 U10328 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i0_4 ), .A3(\SB4_2/i0_0 ), 
        .ZN(n4222) );
  XOR2_X1 U10331 ( .A1(\RI5[3][63] ), .A2(\RI5[3][87] ), .Z(n4225) );
  NAND4_X2 U10335 ( .A1(\SB3_27/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_27/Component_Function_4/NAND4_in[0] ), .A3(n5419), .A4(n4229), 
        .ZN(\SB3_27/buf_output[4] ) );
  XOR2_X1 U10337 ( .A1(\MC_ARK_ARC_1_0/temp2[124] ), .A2(n4232), .Z(
        \MC_ARK_ARC_1_0/temp5[124] ) );
  XOR2_X1 U10338 ( .A1(\RI5[0][118] ), .A2(\RI5[0][124] ), .Z(n4232) );
  NAND4_X2 U10339 ( .A1(\SB2_0_13/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_0_13/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_13/Component_Function_4/NAND4_in[3] ), .A4(n4233), .ZN(
        \SB2_0_13/buf_output[4] ) );
  NAND3_X1 U10340 ( .A1(\SB2_0_13/i0_3 ), .A2(\SB2_0_13/i0[10] ), .A3(
        \SB2_0_13/i0[9] ), .ZN(n4233) );
  XOR2_X1 U10344 ( .A1(n4236), .A2(n4589), .Z(\MC_ARK_ARC_1_4/temp5[47] ) );
  XOR2_X1 U10345 ( .A1(\RI5[4][41] ), .A2(\RI5[4][185] ), .Z(n4236) );
  XOR2_X1 U10346 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[50] ), .A2(\RI5[1][14] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[140] ) );
  NAND3_X1 U10349 ( .A1(\SB4_14/i0[10] ), .A2(\SB4_14/i0[6] ), .A3(
        \SB4_14/i0_3 ), .ZN(n4238) );
  XOR2_X1 U10350 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[18] ), .A2(\RI5[4][174] ), 
        .Z(n1803) );
  NAND3_X1 U10352 ( .A1(\SB4_21/i0[8] ), .A2(\SB4_21/i3[0] ), .A3(
        \SB4_21/i1_5 ), .ZN(n4239) );
  NAND4_X2 U10353 ( .A1(\SB2_4_13/Component_Function_4/NAND4_in[0] ), .A2(
        n1850), .A3(\SB2_4_13/Component_Function_4/NAND4_in[1] ), .A4(n4240), 
        .ZN(\SB2_4_13/buf_output[4] ) );
  XOR2_X1 U10356 ( .A1(n1111), .A2(\MC_ARK_ARC_1_4/temp1[82] ), .Z(
        \MC_ARK_ARC_1_4/temp5[82] ) );
  NAND3_X1 U10357 ( .A1(\SB3_18/i0_4 ), .A2(\SB3_18/i1_7 ), .A3(\SB3_18/i0[8] ), .ZN(\SB3_18/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U10359 ( .A1(\RI5[1][35] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[71] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[161] ) );
  XOR2_X1 U10365 ( .A1(\MC_ARK_ARC_1_1/temp2[174] ), .A2(
        \MC_ARK_ARC_1_1/temp1[174] ), .Z(\MC_ARK_ARC_1_1/temp5[174] ) );
  NAND3_X2 U10370 ( .A1(\SB2_2_8/i0[10] ), .A2(\SB2_2_8/i1[9] ), .A3(
        \SB2_2_8/i1_7 ), .ZN(n4448) );
  XOR2_X1 U10373 ( .A1(\RI5[3][27] ), .A2(\RI5[3][51] ), .Z(n4248) );
  XOR2_X1 U10375 ( .A1(\MC_ARK_ARC_1_2/temp5[75] ), .A2(n4250), .Z(
        \MC_ARK_ARC_1_2/buf_output[75] ) );
  XOR2_X1 U10377 ( .A1(\RI5[2][184] ), .A2(\RI5[2][190] ), .Z(
        \MC_ARK_ARC_1_2/temp1[190] ) );
  XOR2_X1 U10379 ( .A1(n4252), .A2(\MC_ARK_ARC_1_3/temp5[110] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[110] ) );
  XOR2_X1 U10380 ( .A1(\MC_ARK_ARC_1_3/temp3[110] ), .A2(
        \MC_ARK_ARC_1_3/temp4[110] ), .Z(n4252) );
  NAND4_X2 U10389 ( .A1(\SB2_4_12/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_4_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_12/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_4_12/buf_output[1] ) );
  NAND4_X2 U10393 ( .A1(\SB2_2_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_2_19/Component_Function_2/NAND4_in[1] ), .A4(n4258), .ZN(
        \SB2_2_19/buf_output[2] ) );
  NAND3_X2 U10394 ( .A1(\SB2_2_19/i0_3 ), .A2(\SB2_2_19/i0[9] ), .A3(
        \SB2_2_19/i0[8] ), .ZN(n4258) );
  NAND3_X1 U10396 ( .A1(\SB4_27/i0[9] ), .A2(\SB4_27/i0_3 ), .A3(
        \SB4_27/i0[8] ), .ZN(n4486) );
  XOR2_X1 U10397 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[179] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[23] ), .Z(n4259) );
  NAND4_X2 U10399 ( .A1(\SB2_0_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_0_21/Component_Function_0/NAND4_in[1] ), .A3(n4261), .A4(
        \SB2_0_21/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_21/buf_output[0] ) );
  NAND3_X2 U10400 ( .A1(\RI3[0][62] ), .A2(\SB2_0_21/i0_3 ), .A3(
        \SB2_0_21/i0[7] ), .ZN(n4261) );
  XOR2_X1 U10402 ( .A1(\RI5[0][16] ), .A2(\RI5[0][184] ), .Z(n2618) );
  XOR2_X1 U10403 ( .A1(\RI5[4][124] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[160] ), .Z(\MC_ARK_ARC_1_4/temp3[58] ) );
  XOR2_X1 U10404 ( .A1(\MC_ARK_ARC_1_4/temp5[44] ), .A2(n4263), .Z(
        \MC_ARK_ARC_1_4/buf_output[44] ) );
  NAND3_X2 U10406 ( .A1(\SB1_2_6/i0_4 ), .A2(\SB1_2_6/i0_3 ), .A3(
        \SB1_2_6/i1[9] ), .ZN(n4264) );
  NAND3_X1 U10407 ( .A1(\SB1_3_14/i1_5 ), .A2(\SB1_3_14/i1[9] ), .A3(
        \SB1_3_14/i0[10] ), .ZN(\SB1_3_14/Component_Function_2/NAND4_in[0] )
         );
  NAND3_X1 U10408 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i0[9] ), .A3(
        \SB4_12/i0[6] ), .ZN(\SB4_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U10409 ( .A1(\SB2_2_0/i0_3 ), .A2(n5444), .A3(\SB2_2_0/i0[10] ), 
        .ZN(n2566) );
  NAND3_X1 U10413 ( .A1(\SB4_27/i0_4 ), .A2(\SB4_27/i1_7 ), .A3(\SB4_27/i0[8] ), .ZN(\SB4_27/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U10414 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[173] ), .A2(\RI5[4][17] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[107] ) );
  XOR2_X1 U10416 ( .A1(\RI5[1][183] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[177] ), .Z(\MC_ARK_ARC_1_1/temp1[183] ) );
  XOR2_X1 U10420 ( .A1(\RI5[4][17] ), .A2(\RI5[4][41] ), .Z(n4914) );
  XOR2_X1 U10421 ( .A1(\RI5[0][74] ), .A2(\RI5[0][104] ), .Z(n4403) );
  NAND4_X2 U10423 ( .A1(\SB2_3_31/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_31/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_31/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_31/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB2_3_31/buf_output[4] ) );
  XOR2_X1 U10424 ( .A1(\MC_ARK_ARC_1_0/temp1[10] ), .A2(
        \MC_ARK_ARC_1_0/temp3[10] ), .Z(n1579) );
  NAND3_X2 U10428 ( .A1(\SB2_2_2/i0[10] ), .A2(\SB2_2_2/i1_7 ), .A3(n6267), 
        .ZN(\SB2_2_2/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U10431 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[75] ), .A2(\RI5[4][99] ), 
        .Z(n4266) );
  XOR2_X1 U10432 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[129] ), .A2(\RI5[4][123] ), .Z(n4267) );
  NAND2_X1 U10433 ( .A1(\SB1_4_12/i1[9] ), .A2(\RI1[4][119] ), .ZN(
        \SB1_4_12/Component_Function_1/NAND4_in[0] ) );
  XOR2_X1 U10434 ( .A1(\RI5[3][44] ), .A2(\RI5[3][8] ), .Z(n4268) );
  NAND4_X2 U10435 ( .A1(\SB2_4_4/Component_Function_3/NAND4_in[0] ), .A2(n1638), .A3(\SB2_4_4/Component_Function_3/NAND4_in[2] ), .A4(n4269), .ZN(
        \SB2_4_4/buf_output[3] ) );
  XOR2_X1 U10436 ( .A1(\RI5[4][7] ), .A2(\RI5[4][31] ), .Z(
        \MC_ARK_ARC_1_4/temp2[61] ) );
  NAND3_X1 U10437 ( .A1(\SB1_1_13/buf_output[4] ), .A2(\SB2_1_12/i0[9] ), .A3(
        \SB1_1_16/buf_output[1] ), .ZN(n4405) );
  NAND3_X2 U10438 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i0_4 ), .A3(
        \SB2_2_3/i1[9] ), .ZN(\SB2_2_3/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U10440 ( .A1(\MC_ARK_ARC_1_1/temp1[183] ), .A2(n4272), .Z(n4730) );
  XOR2_X1 U10447 ( .A1(\RI5[3][63] ), .A2(\RI5[3][27] ), .Z(n4274) );
  NAND4_X2 U10448 ( .A1(\SB2_3_29/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_3_29/Component_Function_2/NAND4_in[2] ), .A3(n1876), .A4(
        \SB2_3_29/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB2_3_29/buf_output[2] ) );
  NAND4_X2 U10451 ( .A1(\SB2_0_31/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_31/Component_Function_0/NAND4_in[2] ), .A3(n1251), .A4(
        \SB2_0_31/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_31/buf_output[0] ) );
  NAND4_X2 U10452 ( .A1(n2070), .A2(n5396), .A3(n4276), .A4(n4275), .ZN(
        \SB2_1_20/buf_output[3] ) );
  NAND3_X2 U10453 ( .A1(\SB2_1_20/i0_0 ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0_4 ), .ZN(n4275) );
  NAND3_X1 U10455 ( .A1(\SB2_0_24/i3[0] ), .A2(\SB2_0_24/i0[8] ), .A3(
        \SB2_0_24/i1_5 ), .ZN(\SB2_0_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U10458 ( .A1(\SB1_1_0/i0[6] ), .A2(\SB1_1_0/i1_5 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[186] ), .ZN(
        \SB1_1_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U10460 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i0[10] ), .A3(
        \SB1_0_29/i0_4 ), .ZN(\SB1_0_29/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U10462 ( .A1(\SB1_3_27/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_3_27/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_3_27/Component_Function_0/NAND4_in[0] ), .A4(n4279), .ZN(
        \SB1_3_27/buf_output[0] ) );
  NAND4_X2 U10463 ( .A1(\SB2_2_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_5/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_5/Component_Function_4/NAND4_in[1] ), .A4(n4280), .ZN(
        \SB2_2_5/buf_output[4] ) );
  NAND3_X2 U10465 ( .A1(n4281), .A2(\SB1_2_0/Component_Function_0/NAND4_in[2] ), .A3(\SB1_2_0/Component_Function_0/NAND4_in[3] ), .ZN(\SB1_2_0/buf_output[0] ) );
  AND2_X1 U10466 ( .A1(\SB1_2_0/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_0/Component_Function_0/NAND4_in[0] ), .Z(n4281) );
  NAND3_X1 U10468 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i1_7 ), .A3(\SB3_14/i3[0] ), .ZN(n4875) );
  XOR2_X1 U10470 ( .A1(n4283), .A2(n4282), .Z(\MC_ARK_ARC_1_1/temp5[60] ) );
  XOR2_X1 U10471 ( .A1(\RI5[1][6] ), .A2(\RI5[1][54] ), .Z(n4282) );
  XOR2_X1 U10472 ( .A1(\RI5[1][30] ), .A2(\RI5[1][60] ), .Z(n4283) );
  NAND4_X2 U10474 ( .A1(n865), .A2(\SB2_1_15/Component_Function_2/NAND4_in[0] ), .A3(\SB2_1_15/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_1_15/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_1_15/buf_output[2] ) );
  NAND3_X2 U10476 ( .A1(\SB1_3_11/i0[10] ), .A2(\SB1_3_11/i0_0 ), .A3(
        \SB1_3_11/i0[6] ), .ZN(\SB1_3_11/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U10479 ( .A1(\SB1_1_21/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_21/Component_Function_1/NAND4_in[2] ), .A3(n614), .A4(
        \SB1_1_21/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_21/buf_output[1] ) );
  NAND4_X2 U10480 ( .A1(n5357), .A2(n2743), .A3(n4327), .A4(
        \SB2_0_7/Component_Function_5/NAND4_in[0] ), .ZN(\RI5[0][149] ) );
  NAND4_X2 U10481 ( .A1(\SB1_0_29/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_29/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_0_29/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_0_29/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_0_29/buf_output[1] ) );
  NAND4_X2 U10482 ( .A1(n621), .A2(\SB2_2_3/Component_Function_0/NAND4_in[1] ), 
        .A3(n5245), .A4(\SB2_2_3/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_3/buf_output[0] ) );
  NAND4_X2 U10484 ( .A1(\SB1_0_14/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_14/Component_Function_3/NAND4_in[2] ), .A3(n4377), .A4(
        \SB1_0_14/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][117] ) );
  NAND4_X2 U10486 ( .A1(\SB2_4_17/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_4_17/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_4_17/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_4_17/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_4_17/buf_output[2] ) );
  NAND4_X2 U10490 ( .A1(\SB2_3_10/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_10/Component_Function_1/NAND4_in[2] ), .A3(n1625), .A4(
        \SB2_3_10/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_10/buf_output[1] ) );
  XOR2_X1 U10491 ( .A1(n4285), .A2(n1479), .Z(\MC_ARK_ARC_1_2/buf_output[96] )
         );
  XOR2_X1 U10492 ( .A1(\MC_ARK_ARC_1_2/temp1[96] ), .A2(
        \MC_ARK_ARC_1_2/temp2[96] ), .Z(n4285) );
  NAND4_X2 U10493 ( .A1(\SB2_3_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_7/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_5/NAND4_in[0] ), .A4(n4287), .ZN(
        \SB2_3_7/buf_output[5] ) );
  NAND3_X1 U10494 ( .A1(\SB4_29/i0[8] ), .A2(\SB4_29/i3[0] ), .A3(
        \SB4_29/i1_5 ), .ZN(n4288) );
  XOR2_X1 U10498 ( .A1(\MC_ARK_ARC_1_0/temp1[99] ), .A2(
        \MC_ARK_ARC_1_0/temp4[99] ), .Z(n4291) );
  XOR2_X1 U10502 ( .A1(\MC_ARK_ARC_1_0/temp2[164] ), .A2(n4295), .Z(n4772) );
  XOR2_X1 U10503 ( .A1(\RI5[0][158] ), .A2(\RI5[0][164] ), .Z(n4295) );
  NAND4_X2 U10506 ( .A1(\SB1_1_20/Component_Function_2/NAND4_in[1] ), .A2(
        n2450), .A3(\SB1_1_20/Component_Function_2/NAND4_in[2] ), .A4(n4297), 
        .ZN(\SB1_1_20/buf_output[2] ) );
  NAND3_X2 U10507 ( .A1(\SB1_1_20/i0[10] ), .A2(\SB1_1_20/i1[9] ), .A3(
        \SB1_1_20/i1_5 ), .ZN(n4297) );
  XOR2_X1 U10508 ( .A1(\RI5[1][20] ), .A2(\RI5[1][14] ), .Z(n4299) );
  XOR2_X1 U10509 ( .A1(\RI5[3][78] ), .A2(\RI5[3][114] ), .Z(
        \MC_ARK_ARC_1_3/temp3[12] ) );
  XOR2_X1 U10512 ( .A1(\MC_ARK_ARC_1_1/temp1[127] ), .A2(
        \MC_ARK_ARC_1_1/temp2[127] ), .Z(n3154) );
  XOR2_X1 U10514 ( .A1(n4303), .A2(\MC_ARK_ARC_1_3/temp2[70] ), .Z(
        \MC_ARK_ARC_1_3/temp5[70] ) );
  XOR2_X1 U10515 ( .A1(\RI5[3][64] ), .A2(\RI5[3][70] ), .Z(n4303) );
  NAND3_X2 U10516 ( .A1(n600), .A2(\SB2_2_23/i0[9] ), .A3(\SB2_2_23/i0[6] ), 
        .ZN(\SB2_2_23/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U10519 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[62] ), .A2(\RI5[3][98] ), 
        .Z(n4304) );
  NAND4_X2 U10524 ( .A1(\SB2_1_20/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_20/Component_Function_0/NAND4_in[0] ), .A3(n4307), .A4(n1564), 
        .ZN(\SB2_1_20/buf_output[0] ) );
  XOR2_X1 U10527 ( .A1(n4846), .A2(\MC_ARK_ARC_1_2/temp4[164] ), .Z(n4309) );
  INV_X1 U10528 ( .I(\SB1_4_3/buf_output[1] ), .ZN(\SB2_4_31/i1_7 ) );
  INV_X2 U10530 ( .I(\SB1_4_7/buf_output[2] ), .ZN(\SB2_4_4/i1[9] ) );
  XOR2_X1 U10532 ( .A1(n2188), .A2(\MC_ARK_ARC_1_4/temp4[75] ), .Z(n4310) );
  NAND3_X1 U10535 ( .A1(\SB2_3_21/i0[10] ), .A2(\SB2_3_21/i1_5 ), .A3(
        \SB2_3_21/i1[9] ), .ZN(\SB2_3_21/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U10538 ( .A1(n4326), .A2(n4314), .Z(\MC_ARK_ARC_1_3/buf_output[17] )
         );
  XOR2_X1 U10539 ( .A1(\MC_ARK_ARC_1_3/temp4[17] ), .A2(
        \MC_ARK_ARC_1_3/temp2[17] ), .Z(n4314) );
  NAND2_X1 U10541 ( .A1(\SB4_19/i0[10] ), .A2(\SB4_19/i0[9] ), .ZN(n4315) );
  NAND3_X1 U10542 ( .A1(\SB1_2_3/i0[7] ), .A2(\SB1_2_3/i0_0 ), .A3(
        \SB1_2_3/i0_3 ), .ZN(\SB1_2_3/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U10545 ( .A1(\RI5[2][191] ), .A2(\RI5[2][167] ), .Z(
        \MC_ARK_ARC_1_2/temp2[29] ) );
  NAND4_X2 U10546 ( .A1(\SB2_4_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_4_1/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_4_1/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_4_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_4_1/buf_output[5] ) );
  XOR2_X1 U10548 ( .A1(\RI5[3][86] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[20] ), 
        .Z(n4650) );
  XOR2_X1 U10549 ( .A1(\RI5[4][128] ), .A2(\RI5[4][164] ), .Z(n4316) );
  NAND4_X2 U10551 ( .A1(\SB2_2_18/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_2_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_18/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_2_18/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_18/buf_output[1] ) );
  NAND4_X2 U10552 ( .A1(\SB2_0_14/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_0_14/Component_Function_5/NAND4_in[0] ), .A3(
        \SB2_0_14/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_0_14/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_0_14/buf_output[5] ) );
  XOR2_X1 U10553 ( .A1(\MC_ARK_ARC_1_3/temp4[99] ), .A2(n4317), .Z(n2747) );
  XOR2_X1 U10554 ( .A1(\RI5[3][9] ), .A2(\RI5[3][165] ), .Z(n4317) );
  NAND3_X2 U10555 ( .A1(\SB2_0_17/i0[6] ), .A2(\SB2_0_17/i1[9] ), .A3(
        \SB2_0_17/i0_3 ), .ZN(\SB2_0_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U10561 ( .A1(\SB1_0_21/i0[10] ), .A2(\SB1_0_21/i1[9] ), .A3(
        \SB1_0_21/i1_5 ), .ZN(n4406) );
  XOR2_X1 U10567 ( .A1(\MC_ARK_ARC_1_0/temp1[161] ), .A2(n4322), .Z(
        \MC_ARK_ARC_1_0/temp5[161] ) );
  XOR2_X1 U10568 ( .A1(\SB2_0_14/buf_output[5] ), .A2(\RI5[0][131] ), .Z(n4322) );
  XOR2_X1 U10569 ( .A1(\MC_ARK_ARC_1_2/temp4[15] ), .A2(n4324), .Z(n4505) );
  XOR2_X1 U10570 ( .A1(\RI5[2][117] ), .A2(\RI5[2][81] ), .Z(n4324) );
  NAND3_X2 U10572 ( .A1(\SB2_0_14/i1_7 ), .A2(\SB2_0_14/i0[10] ), .A3(
        \SB2_0_14/i1[9] ), .ZN(n4325) );
  NAND3_X2 U10573 ( .A1(\SB2_0_7/i0_0 ), .A2(\SB2_0_7/i0[6] ), .A3(
        \SB2_0_7/i0[10] ), .ZN(n4327) );
  NAND4_X2 U10574 ( .A1(\SB1_4_5/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_4_5/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_4_5/Component_Function_4/NAND4_in[3] ), .A4(n4328), .ZN(
        \SB1_4_5/buf_output[4] ) );
  XOR2_X1 U10575 ( .A1(\RI5[2][180] ), .A2(\RI5[2][186] ), .Z(n4330) );
  XOR2_X1 U10576 ( .A1(n4331), .A2(\MC_ARK_ARC_1_3/temp5[159] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[159] ) );
  XOR2_X1 U10577 ( .A1(\MC_ARK_ARC_1_3/temp3[159] ), .A2(
        \MC_ARK_ARC_1_3/temp4[159] ), .Z(n4331) );
  NAND4_X2 U10580 ( .A1(\SB2_3_2/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_2/Component_Function_0/NAND4_in[2] ), .A3(n4741), .A4(n4333), 
        .ZN(\SB2_3_2/buf_output[0] ) );
  NAND4_X2 U10583 ( .A1(\SB1_3_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_7/Component_Function_0/NAND4_in[0] ), .A4(n4336), .ZN(
        \SB1_3_7/buf_output[0] ) );
  NAND3_X1 U10584 ( .A1(\SB1_1_16/i0[8] ), .A2(\SB1_1_16/i3[0] ), .A3(
        \SB1_1_16/i1_5 ), .ZN(n4337) );
  NAND3_X1 U10585 ( .A1(\SB4_15/i0_3 ), .A2(\SB3_17/buf_output[3] ), .A3(
        \SB4_15/i0[6] ), .ZN(\SB4_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U10587 ( .A1(\SB2_1_7/i0[6] ), .A2(\SB2_1_7/i0[10] ), .A3(
        \SB2_1_7/i0_0 ), .ZN(\SB2_1_7/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U10588 ( .A1(\SB2_2_22/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_22/Component_Function_4/NAND4_in[0] ), .A3(n4708), .A4(
        \SB2_2_22/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_2_22/buf_output[4] ) );
  NAND3_X2 U10589 ( .A1(\SB1_1_29/i0_3 ), .A2(\SB1_1_29/i0_4 ), .A3(
        \SB1_1_29/i1[9] ), .ZN(\SB1_1_29/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U10591 ( .A1(\SB1_1_17/Component_Function_5/NAND4_in[3] ), .A2(
        n1187), .A3(\SB1_1_17/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_1_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_17/buf_output[5] ) );
  NAND2_X1 U10592 ( .A1(\SB1_3_4/i1[9] ), .A2(\RI1[3][167] ), .ZN(
        \SB1_3_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10594 ( .A1(\SB1_4_15/i0[6] ), .A2(\SB1_4_15/i0[10] ), .A3(
        \SB1_4_15/i0_3 ), .ZN(\SB1_4_15/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U10595 ( .A1(n4339), .A2(n4506), .Z(\MC_ARK_ARC_1_3/temp5[97] ) );
  XOR2_X1 U10596 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[43] ), .A2(\RI5[3][67] ), 
        .Z(n4339) );
  XOR2_X1 U10597 ( .A1(\MC_ARK_ARC_1_4/temp1[164] ), .A2(n4340), .Z(
        \MC_ARK_ARC_1_4/temp5[164] ) );
  XOR2_X1 U10598 ( .A1(\RI5[4][134] ), .A2(\RI5[4][110] ), .Z(n4340) );
  XOR2_X1 U10601 ( .A1(\SB2_2_0/buf_output[5] ), .A2(\SB2_2_24/buf_output[5] ), 
        .Z(n4342) );
  XOR2_X1 U10603 ( .A1(n4343), .A2(n5082), .Z(\MC_ARK_ARC_1_3/buf_output[185] ) );
  XOR2_X1 U10604 ( .A1(\RI5[1][92] ), .A2(\RI5[1][98] ), .Z(n4344) );
  XOR2_X1 U10605 ( .A1(\MC_ARK_ARC_1_1/temp5[80] ), .A2(n4345), .Z(
        \MC_ARK_ARC_1_1/buf_output[80] ) );
  XOR2_X1 U10608 ( .A1(n2553), .A2(n4346), .Z(\MC_ARK_ARC_1_1/buf_output[191] ) );
  XOR2_X1 U10609 ( .A1(\RI5[1][43] ), .A2(\RI5[1][67] ), .Z(
        \MC_ARK_ARC_1_1/temp2[97] ) );
  NAND3_X2 U10610 ( .A1(\SB1_3_22/i0[10] ), .A2(\SB1_3_22/i1[9] ), .A3(
        \SB1_3_22/i1_5 ), .ZN(n4347) );
  NAND4_X2 U10611 ( .A1(\SB2_2_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_30/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_30/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_30/buf_output[1] ) );
  XOR2_X1 U10614 ( .A1(\MC_ARK_ARC_1_2/temp6[106] ), .A2(n4348), .Z(
        \MC_ARK_ARC_1_2/buf_output[106] ) );
  XOR2_X1 U10615 ( .A1(\MC_ARK_ARC_1_2/temp1[106] ), .A2(
        \MC_ARK_ARC_1_2/temp2[106] ), .Z(n4348) );
  INV_X1 U10616 ( .I(\SB3_5/buf_output[2] ), .ZN(\SB4_2/i1[9] ) );
  NAND4_X2 U10617 ( .A1(\SB3_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_5/Component_Function_2/NAND4_in[2] ), .A3(n2283), .A4(
        \SB3_5/Component_Function_2/NAND4_in[1] ), .ZN(\SB3_5/buf_output[2] )
         );
  XOR2_X1 U10620 ( .A1(\RI5[0][157] ), .A2(\RI5[0][121] ), .Z(
        \MC_ARK_ARC_1_0/temp3[55] ) );
  NAND3_X1 U10624 ( .A1(\SB4_3/i0_3 ), .A2(\SB4_3/i0_0 ), .A3(\SB4_3/i0[7] ), 
        .ZN(\SB4_3/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U10625 ( .A1(\SB2_4_9/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_9/Component_Function_0/NAND4_in[0] ), .A4(n4355), .ZN(
        \SB2_4_9/buf_output[0] ) );
  XOR2_X1 U10627 ( .A1(\MC_ARK_ARC_1_4/temp5[170] ), .A2(n3159), .Z(
        \MC_ARK_ARC_1_4/buf_output[170] ) );
  NAND3_X1 U10630 ( .A1(\SB4_1/i3[0] ), .A2(\SB4_1/i0[8] ), .A3(n5442), .ZN(
        \SB4_1/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U10635 ( .A1(n1005), .A2(\MC_ARK_ARC_1_0/temp4[116] ), .Z(n1814) );
  XOR2_X1 U10636 ( .A1(n5300), .A2(n5301), .Z(\RI1[5][35] ) );
  XOR2_X1 U10637 ( .A1(n4359), .A2(\MC_ARK_ARC_1_3/temp6[15] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[15] ) );
  NAND3_X1 U10639 ( .A1(\SB1_4_15/i0_3 ), .A2(\SB1_4_15/i0[8] ), .A3(
        \SB1_4_15/i1_7 ), .ZN(\SB1_4_15/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U10640 ( .A1(\MC_ARK_ARC_1_0/temp2[182] ), .A2(
        \MC_ARK_ARC_1_0/temp1[182] ), .Z(\MC_ARK_ARC_1_0/temp5[182] ) );
  XOR2_X1 U10643 ( .A1(\RI5[0][59] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[113] ), 
        .Z(n4362) );
  XOR2_X1 U10645 ( .A1(\RI5[2][116] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[110] ), .Z(\MC_ARK_ARC_1_2/temp1[116] ) );
  XOR2_X1 U10648 ( .A1(n4365), .A2(\MC_ARK_ARC_1_4/temp4[89] ), .Z(n3001) );
  XOR2_X1 U10649 ( .A1(\RI5[4][191] ), .A2(\RI5[4][155] ), .Z(n4365) );
  NAND3_X1 U10650 ( .A1(\SB2_2_31/i0_4 ), .A2(\SB2_2_31/i1_7 ), .A3(
        \SB2_2_31/i0[8] ), .ZN(n4366) );
  INV_X2 U10653 ( .I(\SB1_1_16/buf_output[3] ), .ZN(\SB2_1_14/i0[8] ) );
  INV_X1 U10654 ( .I(\SB1_1_16/buf_output[0] ), .ZN(\SB2_1_11/i3[0] ) );
  NAND4_X2 U10655 ( .A1(\SB1_1_16/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_16/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_1_16/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_1_16/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_16/buf_output[0] ) );
  NAND3_X1 U10656 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i0_3 ), .A3(
        \SB2_3_19/i0[9] ), .ZN(\SB2_3_19/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U10660 ( .A1(\MC_ARK_ARC_1_0/temp5[122] ), .A2(n4456), .Z(
        \MC_ARK_ARC_1_0/buf_output[122] ) );
  NAND3_X1 U10661 ( .A1(\SB3_15/i0[6] ), .A2(\SB3_15/i0[7] ), .A3(
        \SB3_15/i0[8] ), .ZN(\SB3_15/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U10662 ( .A1(n4370), .A2(\MC_ARK_ARC_1_4/temp1[17] ), .Z(n2191) );
  XOR2_X1 U10663 ( .A1(\RI5[4][179] ), .A2(\RI5[4][155] ), .Z(n4370) );
  XOR2_X1 U10665 ( .A1(\RI5[3][150] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[144] ), .Z(n4371) );
  NAND4_X2 U10666 ( .A1(\SB2_3_11/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_11/Component_Function_0/NAND4_in[0] ), .A4(n4372), .ZN(
        \SB2_3_11/buf_output[0] ) );
  NAND4_X2 U10667 ( .A1(\SB2_4_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_4_18/Component_Function_3/NAND4_in[3] ), .A4(n4373), .ZN(
        \SB2_4_18/buf_output[3] ) );
  XOR2_X1 U10669 ( .A1(\MC_ARK_ARC_1_3/temp1[89] ), .A2(n4375), .Z(n2284) );
  XOR2_X1 U10670 ( .A1(\RI5[3][35] ), .A2(\RI5[3][59] ), .Z(n4375) );
  NAND3_X1 U10671 ( .A1(\SB4_8/i0[10] ), .A2(\SB4_8/i1_5 ), .A3(n3996), .ZN(
        n4378) );
  NAND3_X1 U10674 ( .A1(\SB3_21/i0_0 ), .A2(\SB3_21/i3[0] ), .A3(\SB3_21/i1_7 ), .ZN(\SB3_21/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U10678 ( .A1(n877), .A2(n4380), .Z(\MC_ARK_ARC_1_2/buf_output[0] )
         );
  XOR2_X1 U10679 ( .A1(\MC_ARK_ARC_1_2/temp4[0] ), .A2(
        \MC_ARK_ARC_1_2/temp3[0] ), .Z(n4380) );
  XOR2_X1 U10680 ( .A1(n993), .A2(n4381), .Z(\MC_ARK_ARC_1_0/temp5[140] ) );
  XOR2_X1 U10681 ( .A1(\RI5[0][134] ), .A2(\RI5[0][140] ), .Z(n4381) );
  NAND4_X2 U10682 ( .A1(\SB2_0_11/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_0_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_11/Component_Function_0/NAND4_in[0] ), .A4(n4382), .ZN(
        \SB2_0_11/buf_output[0] ) );
  XOR2_X1 U10685 ( .A1(n4383), .A2(\MC_ARK_ARC_1_2/temp5[124] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[124] ) );
  XOR2_X1 U10686 ( .A1(\MC_ARK_ARC_1_2/temp4[124] ), .A2(
        \MC_ARK_ARC_1_2/temp3[124] ), .Z(n4383) );
  XOR2_X1 U10692 ( .A1(\RI5[0][135] ), .A2(\RI5[0][99] ), .Z(
        \MC_ARK_ARC_1_0/temp3[33] ) );
  NAND3_X2 U10693 ( .A1(\SB2_1_27/i1[9] ), .A2(\SB2_1_27/i0_4 ), .A3(
        \SB2_1_27/i0_3 ), .ZN(\SB2_1_27/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U10699 ( .A1(\RI5[3][174] ), .A2(\RI5[3][180] ), .Z(
        \MC_ARK_ARC_1_3/temp1[180] ) );
  XOR2_X1 U10702 ( .A1(\RI5[2][44] ), .A2(\RI5[2][20] ), .Z(
        \MC_ARK_ARC_1_2/temp2[74] ) );
  XOR2_X1 U10703 ( .A1(n4388), .A2(n14), .Z(Ciphertext[81]) );
  NAND4_X2 U10704 ( .A1(\SB4_18/Component_Function_3/NAND4_in[2] ), .A2(
        \SB4_18/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_18/Component_Function_3/NAND4_in[1] ), .A4(n1689), .ZN(n4388) );
  NAND3_X1 U10708 ( .A1(\SB1_1_0/i0[10] ), .A2(\SB1_1_0/i1[9] ), .A3(
        \SB1_1_0/i1_7 ), .ZN(n4391) );
  XOR2_X1 U10709 ( .A1(\MC_ARK_ARC_1_4/temp3[153] ), .A2(
        \MC_ARK_ARC_1_4/temp4[153] ), .Z(\MC_ARK_ARC_1_4/temp6[153] ) );
  NAND3_X2 U10711 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0[8] ), .A3(
        \SB2_2_22/i0[9] ), .ZN(n2017) );
  NAND3_X2 U10712 ( .A1(\SB1_1_17/i0[9] ), .A2(\SB1_1_17/i0_3 ), .A3(
        \SB1_1_17/i0[10] ), .ZN(n4394) );
  NAND4_X2 U10713 ( .A1(n1634), .A2(
        \SB1_1_23/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_23/Component_Function_2/NAND4_in[3] ), .A4(n4395), .ZN(
        \SB1_1_23/buf_output[2] ) );
  NAND3_X2 U10714 ( .A1(\SB1_1_23/i0[10] ), .A2(\SB1_1_23/i0_3 ), .A3(
        \SB1_1_23/i0[6] ), .ZN(n4395) );
  NAND2_X1 U10715 ( .A1(\SB1_2_22/i1[9] ), .A2(\RI1[2][59] ), .ZN(
        \SB1_2_22/Component_Function_1/NAND4_in[0] ) );
  XOR2_X1 U10716 ( .A1(\MC_ARK_ARC_1_2/temp2[24] ), .A2(
        \MC_ARK_ARC_1_2/temp1[24] ), .Z(n1877) );
  OR2_X1 U10722 ( .A1(\SB1_3_13/buf_output[0] ), .A2(\SB1_3_10/buf_output[3] ), 
        .Z(n4398) );
  XOR2_X1 U10725 ( .A1(\MC_ARK_ARC_1_1/temp5[60] ), .A2(n4399), .Z(
        \MC_ARK_ARC_1_1/buf_output[60] ) );
  XOR2_X1 U10726 ( .A1(\MC_ARK_ARC_1_1/temp4[60] ), .A2(
        \MC_ARK_ARC_1_1/temp3[60] ), .Z(n4399) );
  XOR2_X1 U10729 ( .A1(\MC_ARK_ARC_1_0/temp5[73] ), .A2(n4401), .Z(
        \MC_ARK_ARC_1_0/buf_output[73] ) );
  XOR2_X1 U10730 ( .A1(\MC_ARK_ARC_1_0/temp4[73] ), .A2(
        \MC_ARK_ARC_1_0/temp3[73] ), .Z(n4401) );
  XOR2_X1 U10731 ( .A1(n4403), .A2(n4402), .Z(\MC_ARK_ARC_1_0/temp5[104] ) );
  XOR2_X1 U10733 ( .A1(n2952), .A2(n4404), .Z(\MC_ARK_ARC_1_0/buf_output[44] )
         );
  NAND3_X2 U10736 ( .A1(\SB2_2_15/i0[6] ), .A2(\SB2_2_15/i0[9] ), .A3(
        \SB2_2_15/i0_4 ), .ZN(\SB2_2_15/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U10738 ( .A1(n4409), .A2(n4408), .Z(\MC_ARK_ARC_1_4/temp6[39] ) );
  XOR2_X1 U10739 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[75] ), .A2(n434), .Z(
        n4408) );
  XOR2_X1 U10740 ( .A1(\RI5[4][105] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[141] ), .Z(n4409) );
  NAND3_X1 U10741 ( .A1(\SB1_0_14/i0_3 ), .A2(\SB1_0_14/i0_0 ), .A3(
        \SB1_0_14/i0_4 ), .ZN(\SB1_0_14/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U10743 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[147] ), .A2(\RI5[2][111] ), .Z(\MC_ARK_ARC_1_2/temp3[45] ) );
  NAND3_X2 U10744 ( .A1(\SB2_1_12/i0[10] ), .A2(\SB2_1_12/i0_3 ), .A3(
        \SB2_1_12/i0[6] ), .ZN(\SB2_1_12/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U10745 ( .A1(\SB1_0_5/Component_Function_1/NAND4_in[1] ), .A2(n4577), .A3(\SB1_0_5/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_0_5/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_0_5/buf_output[1] ) );
  NAND3_X2 U10751 ( .A1(\SB1_3_4/i0[9] ), .A2(\SB1_3_4/i0[8] ), .A3(
        \RI1[3][167] ), .ZN(n4414) );
  NAND3_X2 U10755 ( .A1(\SB2_2_6/i0_0 ), .A2(\SB2_2_6/i0[10] ), .A3(
        \SB2_2_6/i0[6] ), .ZN(n4417) );
  XOR2_X1 U10756 ( .A1(\SB2_4_25/buf_output[1] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[97] ), .Z(\MC_ARK_ARC_1_4/temp3[187] )
         );
  INV_X2 U10759 ( .I(\SB1_3_2/buf_output[3] ), .ZN(\SB2_3_0/i0[8] ) );
  XOR2_X1 U10760 ( .A1(n2109), .A2(n4419), .Z(\MC_ARK_ARC_1_3/buf_output[155] ) );
  NAND3_X2 U10762 ( .A1(\SB2_3_28/i0_3 ), .A2(\SB1_3_29/buf_output[4] ), .A3(
        \SB2_3_28/i1[9] ), .ZN(n4421) );
  NAND4_X2 U10763 ( .A1(\SB2_4_26/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_4_26/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_4_26/Component_Function_1/NAND4_in[0] ), .A4(n4422), .ZN(
        \SB2_4_26/buf_output[1] ) );
  NAND3_X1 U10764 ( .A1(\SB2_4_26/i0_4 ), .A2(\SB2_4_26/i1_7 ), .A3(
        \SB2_4_26/i0[8] ), .ZN(n4422) );
  XOR2_X1 U10766 ( .A1(\RI5[4][82] ), .A2(\RI5[4][88] ), .Z(n4424) );
  NAND4_X2 U10767 ( .A1(n1743), .A2(\SB3_17/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB3_17/Component_Function_5/NAND4_in[0] ), .A4(n4425), .ZN(
        \SB3_17/buf_output[5] ) );
  NAND3_X2 U10768 ( .A1(\SB3_17/i0_4 ), .A2(\SB3_17/i0[9] ), .A3(
        \SB3_17/i0[6] ), .ZN(n4425) );
  NAND3_X1 U10774 ( .A1(\SB3_21/i0[6] ), .A2(n3182), .A3(\SB3_21/i0[9] ), .ZN(
        \SB3_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U10779 ( .A1(\SB1_3_4/i0[8] ), .A2(\SB1_3_4/i1_7 ), .A3(
        \RI1[3][167] ), .ZN(n4429) );
  XOR2_X1 U10780 ( .A1(\RI5[1][171] ), .A2(\RI5[1][165] ), .Z(n4430) );
  INV_X2 U10781 ( .I(\SB1_1_5/buf_output[5] ), .ZN(\SB2_1_5/i1_5 ) );
  NAND3_X2 U10783 ( .A1(\SB1_4_2/i0[9] ), .A2(\SB1_4_2/i0[6] ), .A3(
        \SB1_4_2/i0_4 ), .ZN(n4431) );
  INV_X1 U10785 ( .I(\SB1_3_29/buf_output[0] ), .ZN(\SB2_3_24/i3[0] ) );
  NAND4_X2 U10786 ( .A1(n2643), .A2(
        \SB1_3_29/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_3_29/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_3_29/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_29/buf_output[0] ) );
  NAND4_X2 U10788 ( .A1(\SB3_5/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_5/Component_Function_1/NAND4_in[3] ), .A3(
        \SB3_5/Component_Function_1/NAND4_in[0] ), .A4(
        \SB3_5/Component_Function_1/NAND4_in[1] ), .ZN(\SB3_5/buf_output[1] )
         );
  XOR2_X1 U10791 ( .A1(\RI5[1][75] ), .A2(\RI5[1][51] ), .Z(
        \MC_ARK_ARC_1_1/temp2[105] ) );
  XOR2_X1 U10792 ( .A1(n4432), .A2(\MC_ARK_ARC_1_4/temp5[158] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[158] ) );
  XOR2_X1 U10793 ( .A1(\MC_ARK_ARC_1_4/temp3[158] ), .A2(
        \MC_ARK_ARC_1_4/temp4[158] ), .Z(n4432) );
  XOR2_X1 U10795 ( .A1(n5313), .A2(\MC_ARK_ARC_1_0/temp6[60] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[60] ) );
  NAND4_X2 U10798 ( .A1(\SB2_2_31/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_31/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_31/Component_Function_4/NAND4_in[2] ), .A4(n4434), .ZN(
        \SB2_2_31/buf_output[4] ) );
  NAND4_X1 U10799 ( .A1(\SB2_0_3/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_0_3/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_3/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_0_3/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_3/buf_output[0] ) );
  XOR2_X1 U10800 ( .A1(\RI5[3][145] ), .A2(\RI5[3][121] ), .Z(
        \MC_ARK_ARC_1_3/temp2[175] ) );
  XOR2_X1 U10802 ( .A1(\RI5[0][110] ), .A2(\RI5[0][146] ), .Z(
        \MC_ARK_ARC_1_0/temp3[44] ) );
  XOR2_X1 U10809 ( .A1(\RI5[3][65] ), .A2(n426), .Z(n4437) );
  XOR2_X1 U10810 ( .A1(\RI5[3][101] ), .A2(\RI5[3][35] ), .Z(n4438) );
  XOR2_X1 U10812 ( .A1(n2795), .A2(n4440), .Z(\MC_ARK_ARC_1_4/temp5[97] ) );
  XOR2_X1 U10813 ( .A1(\RI5[4][91] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[97] ), 
        .Z(n4440) );
  NAND3_X2 U10815 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i0[8] ), .A3(
        \SB2_1_5/i0[9] ), .ZN(n4441) );
  NAND3_X2 U10817 ( .A1(\SB2_2_31/i1_5 ), .A2(\SB2_2_31/i0_0 ), .A3(
        \SB2_2_31/i0_4 ), .ZN(n4443) );
  NAND3_X2 U10819 ( .A1(\SB1_0_5/i0_3 ), .A2(\SB1_0_5/i0_4 ), .A3(
        \SB1_0_5/i1[9] ), .ZN(\SB1_0_5/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U10820 ( .A1(\RI5[2][33] ), .A2(\RI5[2][69] ), .Z(
        \MC_ARK_ARC_1_2/temp3[159] ) );
  XOR2_X1 U10821 ( .A1(\MC_ARK_ARC_1_2/temp6[159] ), .A2(
        \MC_ARK_ARC_1_2/temp5[159] ), .Z(\MC_ARK_ARC_1_2/buf_output[159] ) );
  NAND3_X2 U10823 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0[10] ), .A3(
        \SB2_2_22/i0[9] ), .ZN(n4708) );
  INV_X4 U10824 ( .I(n4677), .ZN(n592) );
  NAND3_X1 U10825 ( .A1(\SB2_4_26/i0_3 ), .A2(\SB2_4_26/i0[10] ), .A3(
        \SB2_4_26/i0_4 ), .ZN(\SB2_4_26/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U10829 ( .A1(n635), .A2(\MC_ARK_ARC_1_4/temp5[97] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[97] ) );
  NAND4_X2 U10830 ( .A1(\SB1_3_10/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_10/Component_Function_5/NAND4_in[3] ), .A3(n2309), .A4(
        \SB1_3_10/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_10/buf_output[5] ) );
  XOR2_X1 U10832 ( .A1(\RI5[0][188] ), .A2(\RI5[0][2] ), .Z(n4446) );
  INV_X1 U10833 ( .I(\SB3_4/buf_output[1] ), .ZN(\SB4_0/i1_7 ) );
  NAND4_X2 U10834 ( .A1(\SB3_4/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_4/Component_Function_1/NAND4_in[3] ), .A4(
        \SB3_4/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_4/buf_output[1] )
         );
  NAND4_X2 U10835 ( .A1(\SB2_2_15/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_15/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_15/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_2_15/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_15/buf_output[0] ) );
  NAND3_X2 U10839 ( .A1(\SB2_1_8/i0_3 ), .A2(\SB2_1_8/i1[9] ), .A3(
        \SB2_1_8/i0_4 ), .ZN(n859) );
  INV_X2 U10840 ( .I(\SB1_2_11/buf_output[3] ), .ZN(\SB2_2_9/i0[8] ) );
  NAND3_X1 U10842 ( .A1(\SB2_0_26/i1[9] ), .A2(\RI3[0][33] ), .A3(
        \SB2_0_26/i1_5 ), .ZN(\SB2_0_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U10843 ( .A1(\SB2_0_0/i0[9] ), .A2(\SB2_0_0/i0_3 ), .A3(n4003), 
        .ZN(\SB2_0_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U10845 ( .A1(\SB1_0_5/i0[6] ), .A2(\SB1_0_5/i0[8] ), .A3(
        \SB1_0_5/i0[7] ), .ZN(\SB1_0_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U10846 ( .A1(\SB1_1_19/i0[8] ), .A2(\SB1_1_19/i1_5 ), .A3(
        \SB1_1_19/i3[0] ), .ZN(n4450) );
  NAND4_X2 U10849 ( .A1(n2409), .A2(\SB3_1/Component_Function_0/NAND4_in[1] ), 
        .A3(n2408), .A4(\SB3_1/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB3_1/buf_output[0] ) );
  NAND4_X2 U10850 ( .A1(\SB2_1_23/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_23/Component_Function_0/NAND4_in[0] ), .A4(n4454), .ZN(
        \SB2_1_23/buf_output[0] ) );
  XOR2_X1 U10851 ( .A1(n4455), .A2(n4715), .Z(\MC_ARK_ARC_1_1/buf_output[168] ) );
  XOR2_X1 U10852 ( .A1(\MC_ARK_ARC_1_1/temp4[168] ), .A2(
        \MC_ARK_ARC_1_1/temp3[168] ), .Z(n4455) );
  XOR2_X1 U10854 ( .A1(\MC_ARK_ARC_1_0/temp3[122] ), .A2(
        \MC_ARK_ARC_1_0/temp4[122] ), .Z(n4456) );
  XOR2_X1 U10855 ( .A1(n4555), .A2(\MC_ARK_ARC_1_1/temp6[154] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[154] ) );
  XOR2_X1 U10857 ( .A1(\RI5[1][149] ), .A2(n210), .Z(n4457) );
  NAND4_X2 U10858 ( .A1(\SB1_4_0/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_4_0/Component_Function_5/NAND4_in[2] ), .A3(n830), .A4(n4459), 
        .ZN(\SB1_4_0/buf_output[5] ) );
  NAND2_X1 U10859 ( .A1(\SB1_4_0/i3[0] ), .A2(\SB1_4_0/i0_0 ), .ZN(n4459) );
  NAND4_X2 U10860 ( .A1(\SB1_4_18/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_4_18/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_4_18/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_4_18/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_4_18/buf_output[1] ) );
  NAND4_X2 U10864 ( .A1(\SB2_1_21/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_21/Component_Function_0/NAND4_in[2] ), .A3(n1465), .A4(
        \SB2_1_21/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_21/buf_output[0] ) );
  NAND4_X2 U10866 ( .A1(\SB2_1_31/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_31/Component_Function_4/NAND4_in[0] ), .A4(n4460), .ZN(
        \SB2_1_31/buf_output[4] ) );
  NAND3_X2 U10867 ( .A1(\SB2_4_24/i0_3 ), .A2(\SB2_4_24/i0_4 ), .A3(n5443), 
        .ZN(\SB2_4_24/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U10868 ( .A1(\SB2_0_19/i0[6] ), .A2(\SB2_0_19/i0[9] ), .A3(
        \RI3[0][76] ), .ZN(\SB2_0_19/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U10869 ( .A1(\MC_ARK_ARC_1_0/temp5[181] ), .A2(n733), .Z(
        \MC_ARK_ARC_1_0/buf_output[181] ) );
  NAND4_X2 U10874 ( .A1(\SB1_0_1/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_1/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_1/Component_Function_4/NAND4_in[2] ), .A4(n4463), .ZN(
        \SB1_0_1/buf_output[4] ) );
  NAND3_X1 U10875 ( .A1(\SB1_0_1/i0_4 ), .A2(\SB1_0_1/i1_5 ), .A3(
        \SB1_0_1/i1[9] ), .ZN(n4463) );
  NAND3_X1 U10876 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0_0 ), .A3(
        \SB2_2_29/i0[7] ), .ZN(\SB2_2_29/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U10877 ( .A1(\SB2_3_6/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_6/Component_Function_0/NAND4_in[0] ), .A4(n4464), .ZN(
        \SB2_3_6/buf_output[0] ) );
  NAND3_X1 U10883 ( .A1(\SB1_2_9/i0[6] ), .A2(\SB1_2_9/i0[9] ), .A3(
        \MC_ARK_ARC_1_1/buf_output[136] ), .ZN(n4466) );
  XOR2_X1 U10884 ( .A1(\MC_ARK_ARC_1_1/temp2[166] ), .A2(n4467), .Z(
        \MC_ARK_ARC_1_1/temp5[166] ) );
  XOR2_X1 U10885 ( .A1(\RI5[1][166] ), .A2(\RI5[1][160] ), .Z(n4467) );
  NAND4_X2 U10886 ( .A1(\SB2_2_8/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_8/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_8/Component_Function_0/NAND4_in[0] ), .A4(n4469), .ZN(
        \SB2_2_8/buf_output[0] ) );
  XOR2_X1 U10890 ( .A1(n4471), .A2(\MC_ARK_ARC_1_2/temp2[131] ), .Z(
        \MC_ARK_ARC_1_2/temp5[131] ) );
  XOR2_X1 U10891 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[131] ), .A2(\RI5[2][125] ), .Z(n4471) );
  XOR2_X1 U10896 ( .A1(\MC_ARK_ARC_1_1/temp6[46] ), .A2(
        \MC_ARK_ARC_1_1/temp5[46] ), .Z(\MC_ARK_ARC_1_1/buf_output[46] ) );
  XOR2_X1 U10899 ( .A1(n4478), .A2(\MC_ARK_ARC_1_3/temp6[79] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[79] ) );
  XOR2_X1 U10900 ( .A1(n2917), .A2(n2916), .Z(n4478) );
  INV_X2 U10901 ( .I(\SB1_2_8/buf_output[2] ), .ZN(\SB2_2_5/i1[9] ) );
  NAND4_X2 U10902 ( .A1(\SB2_0_22/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_22/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_22/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_22/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB2_0_22/buf_output[2] ) );
  NAND2_X2 U10903 ( .A1(n3033), .A2(\SB1_0_0/Component_Function_0/NAND4_in[3] ), .ZN(\SB2_0_27/i0[9] ) );
  NAND3_X1 U10913 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i0[9] ), .A3(
        \SB1_0_29/i0[8] ), .ZN(\SB1_0_29/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U10916 ( .A1(n4488), .A2(\MC_ARK_ARC_1_2/temp4[25] ), .Z(
        \MC_ARK_ARC_1_2/temp6[25] ) );
  XOR2_X1 U10917 ( .A1(\RI5[2][127] ), .A2(\RI5[2][91] ), .Z(n4488) );
  NAND4_X2 U10919 ( .A1(\SB3_0/Component_Function_0/NAND4_in[1] ), .A2(
        \SB3_0/Component_Function_0/NAND4_in[3] ), .A3(
        \SB3_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_0/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_0/buf_output[0] )
         );
  XOR2_X1 U10921 ( .A1(\MC_ARK_ARC_1_4/temp2[187] ), .A2(
        \MC_ARK_ARC_1_4/temp1[187] ), .Z(\MC_ARK_ARC_1_4/temp5[187] ) );
  XOR2_X1 U10924 ( .A1(n4490), .A2(n4787), .Z(\MC_ARK_ARC_1_1/buf_output[44] )
         );
  XOR2_X1 U10926 ( .A1(n4986), .A2(\MC_ARK_ARC_1_3/temp4[59] ), .Z(n4602) );
  NAND3_X1 U10929 ( .A1(\SB4_18/i0[10] ), .A2(n1496), .A3(\SB4_18/i1_7 ), .ZN(
        \SB4_18/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U10930 ( .A1(n4563), .A2(\SB1_1_7/Component_Function_5/NAND4_in[1] ), .A3(\SB1_1_7/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_1_7/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_7/buf_output[5] ) );
  NAND3_X1 U10935 ( .A1(\SB2_2_15/i0[9] ), .A2(\RI3[2][97] ), .A3(
        \SB2_2_15/i1_5 ), .ZN(n4492) );
  NAND3_X1 U10937 ( .A1(\SB2_0_10/i0_4 ), .A2(\SB2_0_10/i1_5 ), .A3(n1501), 
        .ZN(\SB2_0_10/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U10938 ( .A1(\SB1_4_14/Component_Function_3/NAND4_in[0] ), .A2(
        n2839), .A3(n4688), .A4(n4493), .ZN(\SB1_4_14/buf_output[3] ) );
  XOR2_X1 U10939 ( .A1(n4494), .A2(\MC_ARK_ARC_1_4/temp6[174] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[174] ) );
  XOR2_X1 U10940 ( .A1(\MC_ARK_ARC_1_4/temp1[174] ), .A2(
        \MC_ARK_ARC_1_4/temp2[174] ), .Z(n4494) );
  XOR2_X1 U10941 ( .A1(n604), .A2(n603), .Z(\MC_ARK_ARC_1_3/buf_output[102] )
         );
  XOR2_X1 U10942 ( .A1(n4496), .A2(n4495), .Z(\MC_ARK_ARC_1_1/buf_output[134] ) );
  INV_X2 U10944 ( .I(\SB1_1_1/buf_output[5] ), .ZN(\SB2_1_1/i1_5 ) );
  NAND3_X2 U10946 ( .A1(\SB2_0_6/i0_3 ), .A2(\SB2_0_6/i0_0 ), .A3(
        \SB2_0_6/i0[7] ), .ZN(n4497) );
  NAND4_X2 U10948 ( .A1(\SB3_15/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_15/Component_Function_1/NAND4_in[0] ), .A4(n4500), .ZN(
        \SB3_15/buf_output[1] ) );
  NAND3_X1 U10949 ( .A1(\SB3_15/i0_4 ), .A2(\SB3_15/i1_7 ), .A3(\SB3_15/i0[8] ), .ZN(n4500) );
  XOR2_X1 U10951 ( .A1(n4501), .A2(\MC_ARK_ARC_1_2/temp5[43] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[43] ) );
  XOR2_X1 U10952 ( .A1(\MC_ARK_ARC_1_2/temp3[43] ), .A2(
        \MC_ARK_ARC_1_2/temp4[43] ), .Z(n4501) );
  XOR2_X1 U10955 ( .A1(\RI5[2][152] ), .A2(\RI5[2][188] ), .Z(
        \MC_ARK_ARC_1_2/temp3[86] ) );
  NAND4_X2 U10956 ( .A1(\SB2_3_26/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_2/NAND4_in[2] ), .A4(n4504), .ZN(
        \SB2_3_26/buf_output[2] ) );
  NAND3_X2 U10957 ( .A1(\SB2_3_26/i0_0 ), .A2(\SB2_3_26/i0_4 ), .A3(
        \SB2_3_26/i1_5 ), .ZN(n4504) );
  XOR2_X1 U10958 ( .A1(n4505), .A2(\MC_ARK_ARC_1_2/temp5[15] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[15] ) );
  XOR2_X1 U10961 ( .A1(\RI5[3][97] ), .A2(\RI5[3][91] ), .Z(n4506) );
  NAND3_X2 U10962 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i1[9] ), .A3(
        \SB2_2_3/i0[6] ), .ZN(\SB2_2_3/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U10963 ( .A1(\MC_ARK_ARC_1_0/temp3[52] ), .A2(
        \MC_ARK_ARC_1_0/temp4[52] ), .Z(\MC_ARK_ARC_1_0/temp6[52] ) );
  XOR2_X1 U10967 ( .A1(n4508), .A2(n4507), .Z(n4562) );
  XOR2_X1 U10968 ( .A1(\RI5[2][176] ), .A2(n70), .Z(n4507) );
  XOR2_X1 U10969 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[110] ), .A2(\RI5[2][140] ), .Z(n4508) );
  NAND3_X1 U10971 ( .A1(\SB1_1_4/i0_0 ), .A2(\SB1_1_4/i0[8] ), .A3(
        \SB1_1_4/i0[9] ), .ZN(n2660) );
  NAND4_X2 U10975 ( .A1(\SB1_3_13/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_13/Component_Function_3/NAND4_in[0] ), .A3(n4770), .A4(n715), 
        .ZN(\SB1_3_13/buf_output[3] ) );
  NAND3_X2 U10976 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0[9] ), .A3(
        \SB2_3_0/i0[8] ), .ZN(\SB2_3_0/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U10977 ( .A1(\SB2_2_13/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_13/Component_Function_0/NAND4_in[2] ), .A3(n4693), .A4(
        \SB2_2_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_13/buf_output[0] ) );
  NAND4_X2 U10979 ( .A1(\SB3_2/Component_Function_5/NAND4_in[1] ), .A2(n2390), 
        .A3(n2018), .A4(\SB3_2/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_2/buf_output[5] ) );
  XOR2_X1 U10982 ( .A1(\MC_ARK_ARC_1_0/temp2[147] ), .A2(n4510), .Z(n1487) );
  XOR2_X1 U10983 ( .A1(\RI5[0][147] ), .A2(\RI5[0][141] ), .Z(n4510) );
  NAND3_X1 U10986 ( .A1(\SB2_0_27/i0[10] ), .A2(\SB2_0_27/i0[9] ), .A3(
        \SB2_0_27/i0_3 ), .ZN(\SB2_0_27/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U10987 ( .A1(\RI5[2][39] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[3] ), 
        .Z(n5302) );
  XOR2_X1 U10988 ( .A1(\RI5[4][50] ), .A2(\RI5[4][74] ), .Z(
        \MC_ARK_ARC_1_4/temp2[104] ) );
  XOR2_X1 U10990 ( .A1(\MC_ARK_ARC_1_2/temp5[144] ), .A2(
        \MC_ARK_ARC_1_2/temp6[144] ), .Z(\MC_ARK_ARC_1_2/buf_output[144] ) );
  XOR2_X1 U10991 ( .A1(\MC_ARK_ARC_1_2/temp5[181] ), .A2(n5174), .Z(
        \MC_ARK_ARC_1_2/buf_output[181] ) );
  XOR2_X1 U10993 ( .A1(\RI5[1][90] ), .A2(\RI5[1][66] ), .Z(n4513) );
  NAND3_X1 U10997 ( .A1(\SB2_1_0/i0_3 ), .A2(\SB1_1_4/buf_output[1] ), .A3(
        \SB2_1_0/i1[9] ), .ZN(n4516) );
  NAND3_X1 U10998 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i0_0 ), .A3(
        \SB2_3_23/i0_4 ), .ZN(n4517) );
  XOR2_X1 U11000 ( .A1(n4519), .A2(n4518), .Z(\MC_ARK_ARC_1_4/temp6[124] ) );
  XOR2_X1 U11001 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[160] ), .A2(n98), .Z(
        n4518) );
  NAND3_X1 U11004 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i0_0 ), .A3(
        \SB1_0_29/i0_4 ), .ZN(\SB1_0_29/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U11006 ( .A1(\MC_ARK_ARC_1_3/temp3[123] ), .A2(
        \MC_ARK_ARC_1_3/temp4[123] ), .Z(\MC_ARK_ARC_1_3/temp6[123] ) );
  NAND3_X1 U11010 ( .A1(n6274), .A2(\SB1_3_1/buf_output[1] ), .A3(
        \SB2_3_29/i0[8] ), .ZN(\SB2_3_29/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U11011 ( .A1(\SB2_4_28/i0_0 ), .A2(\SB2_4_28/i0[10] ), .A3(
        \SB2_4_28/i0[6] ), .ZN(n4532) );
  NAND3_X2 U11015 ( .A1(\SB2_2_1/i0[10] ), .A2(\SB2_2_1/i1_7 ), .A3(
        \SB2_2_1/i1[9] ), .ZN(n4526) );
  XOR2_X1 U11016 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[39] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[75] ), .Z(\MC_ARK_ARC_1_4/temp3[165] )
         );
  NAND3_X2 U11017 ( .A1(\SB2_2_2/i0[10] ), .A2(\SB2_2_2/i0_0 ), .A3(
        \SB2_2_2/i0[6] ), .ZN(n4527) );
  XOR2_X1 U11018 ( .A1(n4529), .A2(n4528), .Z(\MC_ARK_ARC_1_2/temp6[33] ) );
  XOR2_X1 U11019 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), .A2(n74), .Z(n4528) );
  XOR2_X1 U11020 ( .A1(\RI5[2][69] ), .A2(\RI5[2][135] ), .Z(n4529) );
  NAND3_X1 U11021 ( .A1(\SB2_3_26/i1_5 ), .A2(\SB2_3_26/i0_4 ), .A3(
        \SB2_3_26/i1[9] ), .ZN(\SB2_3_26/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U11022 ( .A1(\SB2_4_28/Component_Function_5/NAND4_in[0] ), .A2(
        n4532), .A3(n4531), .A4(n4530), .ZN(\SB2_4_28/buf_output[5] ) );
  XOR2_X1 U11024 ( .A1(n3167), .A2(\RI5[1][14] ), .Z(
        \MC_ARK_ARC_1_1/temp1[14] ) );
  AND3_X1 U11025 ( .A1(n295), .A2(n360), .A3(n242), .Z(n4804) );
  NAND4_X2 U11026 ( .A1(\SB2_1_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_0/Component_Function_5/NAND4_in[1] ), .A3(n914), .A4(
        \SB2_1_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_0/buf_output[5] ) );
  NAND3_X1 U11030 ( .A1(\SB1_4_29/i1_5 ), .A2(\SB1_4_29/i1[9] ), .A3(
        \SB1_4_29/i0_4 ), .ZN(n4533) );
  NAND3_X2 U11031 ( .A1(\SB2_0_19/i0[8] ), .A2(\RI3[0][77] ), .A3(
        \SB2_0_19/i1_7 ), .ZN(\SB2_0_19/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U11033 ( .A1(\MC_ARK_ARC_1_2/temp3[145] ), .A2(
        \MC_ARK_ARC_1_2/temp4[145] ), .Z(n4534) );
  NAND4_X2 U11034 ( .A1(\SB1_0_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_23/Component_Function_1/NAND4_in[0] ), .A3(n1904), .A4(n1905), 
        .ZN(\SB1_0_23/buf_output[1] ) );
  NAND4_X2 U11037 ( .A1(\SB2_0_26/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_26/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_0_26/Component_Function_1/NAND4_in[2] ), .A4(n4535), .ZN(
        \SB2_0_26/buf_output[1] ) );
  NAND3_X2 U11041 ( .A1(\SB2_0_19/i0[6] ), .A2(\RI3[0][75] ), .A3(\RI3[0][77] ), .ZN(\SB2_0_19/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U11042 ( .A1(\SB2_1_5/Component_Function_0/NAND4_in[1] ), .A2(n5286), .A3(n5285), .A4(\SB2_1_5/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_5/buf_output[0] ) );
  NAND3_X2 U11044 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i1[9] ), .A3(
        \SB1_0_23/i0_4 ), .ZN(\SB1_0_23/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U11045 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i0[8] ), .A3(
        \SB1_1_0/i1_7 ), .ZN(\SB1_1_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U11048 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i0[8] ), .A3(
        \SB1_3_10/i1_7 ), .ZN(\SB1_3_10/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U11050 ( .A1(\SB1_3_27/i0_3 ), .A2(\SB1_3_27/i1[9] ), .A3(
        \SB1_3_27/i0_4 ), .ZN(n4538) );
  XOR2_X1 U11051 ( .A1(n4539), .A2(\MC_ARK_ARC_1_4/temp5[138] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[138] ) );
  XOR2_X1 U11052 ( .A1(\MC_ARK_ARC_1_4/temp3[138] ), .A2(
        \MC_ARK_ARC_1_4/temp4[138] ), .Z(n4539) );
  XOR2_X1 U11053 ( .A1(n4540), .A2(\MC_ARK_ARC_1_4/temp6[78] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[78] ) );
  XOR2_X1 U11054 ( .A1(\MC_ARK_ARC_1_4/temp2[78] ), .A2(
        \MC_ARK_ARC_1_4/temp1[78] ), .Z(n4540) );
  NAND3_X1 U11058 ( .A1(\SB1_0_24/i0_4 ), .A2(\SB1_0_24/i1_5 ), .A3(
        \SB1_0_24/i1[9] ), .ZN(n2396) );
  NAND4_X2 U11060 ( .A1(n5324), .A2(n5281), .A3(
        \SB2_0_20/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_20/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_20/buf_output[5] ) );
  NAND4_X1 U11061 ( .A1(\SB2_0_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_3/NAND4_in[1] ), .A3(n4541), .A4(
        \SB2_0_28/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_28/buf_output[3] ) );
  XOR2_X1 U11063 ( .A1(\RI5[1][17] ), .A2(\RI5[1][23] ), .Z(n4542) );
  NAND4_X2 U11067 ( .A1(\SB1_2_24/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_24/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_24/Component_Function_0/NAND4_in[1] ), .A4(n4544), .ZN(
        \SB1_2_24/buf_output[0] ) );
  INV_X2 U11069 ( .I(\SB1_2_24/buf_output[2] ), .ZN(\SB2_2_21/i1[9] ) );
  XOR2_X1 U11070 ( .A1(\RI5[0][85] ), .A2(n7134), .Z(
        \MC_ARK_ARC_1_0/temp3[19] ) );
  XOR2_X1 U11072 ( .A1(\RI5[2][123] ), .A2(\RI5[2][117] ), .Z(
        \MC_ARK_ARC_1_2/temp1[123] ) );
  XOR2_X1 U11073 ( .A1(n2914), .A2(n4545), .Z(\MC_ARK_ARC_1_0/buf_output[4] )
         );
  NAND3_X2 U11075 ( .A1(\SB2_2_26/i0[10] ), .A2(\SB2_2_26/i1[9] ), .A3(
        \SB2_2_26/i1_5 ), .ZN(\SB2_2_26/Component_Function_2/NAND4_in[0] ) );
  NOR2_X2 U11076 ( .A1(n2605), .A2(n4546), .ZN(n3104) );
  NAND3_X2 U11081 ( .A1(\SB2_2_11/i0_0 ), .A2(\SB2_2_11/i0_4 ), .A3(
        \SB2_2_11/i1_5 ), .ZN(n4549) );
  XOR2_X1 U11082 ( .A1(n4550), .A2(\MC_ARK_ARC_1_2/temp5[49] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[49] ) );
  XOR2_X1 U11083 ( .A1(\MC_ARK_ARC_1_2/temp4[49] ), .A2(
        \MC_ARK_ARC_1_2/temp3[49] ), .Z(n4550) );
  INV_X2 U11084 ( .I(n4551), .ZN(\SB1_4_10/i0[8] ) );
  XOR2_X1 U11085 ( .A1(n3025), .A2(\MC_ARK_ARC_1_3/temp6[129] ), .Z(n4551) );
  INV_X2 U11086 ( .I(\SB1_0_29/buf_output[2] ), .ZN(\SB2_0_26/i1[9] ) );
  NAND3_X1 U11088 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i1[9] ), .A3(
        \SB1_0_21/i0_4 ), .ZN(\SB1_0_21/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U11089 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0_0 ), .A3(
        \SB2_2_20/i0_4 ), .ZN(\SB2_2_20/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U11091 ( .I(\RI3[0][122] ), .ZN(\SB2_0_11/i1[9] ) );
  XOR2_X1 U11092 ( .A1(\MC_ARK_ARC_1_0/temp5[104] ), .A2(n4552), .Z(
        \MC_ARK_ARC_1_0/buf_output[104] ) );
  XOR2_X1 U11093 ( .A1(\MC_ARK_ARC_1_0/temp3[104] ), .A2(
        \MC_ARK_ARC_1_0/temp4[104] ), .Z(n4552) );
  NAND3_X1 U11094 ( .A1(\SB3_4/i0[10] ), .A2(\SB3_4/i1[9] ), .A3(\SB3_4/i1_5 ), 
        .ZN(\SB3_4/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U11095 ( .A1(n1351), .A2(n4553), .Z(\MC_ARK_ARC_1_0/buf_output[141] ) );
  XOR2_X1 U11096 ( .A1(\MC_ARK_ARC_1_0/temp1[141] ), .A2(
        \MC_ARK_ARC_1_0/temp4[141] ), .Z(n4553) );
  XOR2_X1 U11098 ( .A1(n4556), .A2(\MC_ARK_ARC_1_1/temp6[153] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[153] ) );
  NAND3_X2 U11100 ( .A1(\SB1_0_25/i0[10] ), .A2(\SB1_0_25/i1_7 ), .A3(
        \SB1_0_25/i1[9] ), .ZN(n4557) );
  XOR2_X1 U11101 ( .A1(n4559), .A2(n4558), .Z(n2780) );
  XOR2_X1 U11102 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[93] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[45] ), .Z(n4558) );
  XOR2_X1 U11103 ( .A1(\RI5[4][69] ), .A2(\RI5[4][99] ), .Z(n4559) );
  XOR2_X1 U11104 ( .A1(n4561), .A2(n4560), .Z(\MC_ARK_ARC_1_1/temp5[83] ) );
  XOR2_X1 U11105 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[83] ), .A2(\RI5[1][53] ), 
        .Z(n4560) );
  XOR2_X1 U11106 ( .A1(n4562), .A2(\MC_ARK_ARC_1_2/temp5[74] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[74] ) );
  NAND3_X1 U11112 ( .A1(\SB1_1_1/i0[10] ), .A2(\SB1_1_1/i1[9] ), .A3(
        \SB1_1_1/i1_5 ), .ZN(\SB1_1_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U11116 ( .A1(\SB1_0_10/i3[0] ), .A2(\SB1_0_10/i1_5 ), .A3(
        \SB1_0_10/i0[8] ), .ZN(n4568) );
  XOR2_X1 U11118 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[125] ), .A2(\RI5[1][161] ), .Z(n4569) );
  XOR2_X1 U11119 ( .A1(n1394), .A2(n4570), .Z(\MC_ARK_ARC_1_4/buf_output[183] ) );
  XOR2_X1 U11120 ( .A1(\MC_ARK_ARC_1_4/temp4[183] ), .A2(n4857), .Z(n4570) );
  INV_X2 U11121 ( .I(\SB1_1_6/buf_output[3] ), .ZN(\SB2_1_4/i0[8] ) );
  NAND3_X1 U11126 ( .A1(\SB1_4_20/i0_3 ), .A2(\SB1_4_20/i0[6] ), .A3(
        \SB1_4_20/i1[9] ), .ZN(\SB1_4_20/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U11131 ( .A1(\RI5[1][55] ), .A2(\RI5[1][19] ), .Z(
        \MC_ARK_ARC_1_1/temp3[145] ) );
  NAND3_X1 U11132 ( .A1(\SB3_19/i0[10] ), .A2(\SB3_19/i1[9] ), .A3(
        \SB3_19/i1_7 ), .ZN(\SB3_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U11133 ( .A1(\SB1_0_5/i0[6] ), .A2(\SB1_0_5/i0[10] ), .A3(
        \SB1_0_5/i0_3 ), .ZN(n4574) );
  XOR2_X1 U11136 ( .A1(\RI5[4][17] ), .A2(\RI5[4][47] ), .Z(n4589) );
  XOR2_X1 U11137 ( .A1(\RI5[4][149] ), .A2(\RI5[4][113] ), .Z(
        \MC_ARK_ARC_1_4/temp3[47] ) );
  NAND4_X2 U11139 ( .A1(\SB2_0_20/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_20/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_0_20/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_0_20/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_20/buf_output[0] ) );
  NAND3_X2 U11141 ( .A1(\SB1_0_1/i0_4 ), .A2(\SB1_0_1/i0_3 ), .A3(
        \SB1_0_1/i1[9] ), .ZN(n4575) );
  NAND4_X2 U11142 ( .A1(\SB4_26/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_26/Component_Function_0/NAND4_in[1] ), .A3(n702), .A4(n4576), 
        .ZN(n4611) );
  NAND2_X1 U11143 ( .A1(\SB4_26/i0[10] ), .A2(\SB4_26/i0[9] ), .ZN(n4576) );
  NAND4_X2 U11144 ( .A1(\SB1_0_5/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_5/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_5/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_5/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_0_5/buf_output[5] ) );
  INV_X1 U11146 ( .I(\SB1_1_27/buf_output[1] ), .ZN(\SB2_1_23/i1_7 ) );
  XOR2_X1 U11149 ( .A1(\RI5[4][48] ), .A2(\RI5[4][72] ), .Z(n4581) );
  XOR2_X1 U11150 ( .A1(\RI5[4][48] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[54] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[54] ) );
  NAND4_X2 U11154 ( .A1(\SB1_2_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_2_28/Component_Function_4/NAND4_in[1] ), .A4(n4584), .ZN(
        \SB1_2_28/buf_output[4] ) );
  NAND2_X1 U11157 ( .A1(\SB1_3_7/i3[0] ), .A2(\MC_ARK_ARC_1_2/buf_output[146] ), .ZN(n4585) );
  XOR2_X1 U11159 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[39] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[45] ), .Z(\MC_ARK_ARC_1_4/temp1[45] ) );
  NAND3_X2 U11160 ( .A1(\SB1_1_8/i0_3 ), .A2(\SB1_1_8/i0_4 ), .A3(
        \SB1_1_8/i1[9] ), .ZN(n4588) );
  NAND3_X1 U11161 ( .A1(\SB1_2_28/i0[10] ), .A2(\SB1_2_28/i1[9] ), .A3(
        \SB1_2_28/i1_5 ), .ZN(\SB1_2_28/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U11162 ( .A1(\MC_ARK_ARC_1_0/temp3[46] ), .A2(
        \MC_ARK_ARC_1_0/temp4[46] ), .Z(\MC_ARK_ARC_1_0/temp6[46] ) );
  NAND3_X2 U11167 ( .A1(\SB1_3_12/i0[9] ), .A2(\SB1_3_12/i0_4 ), .A3(
        \SB1_3_12/i0[6] ), .ZN(n4591) );
  NAND4_X2 U11168 ( .A1(\SB2_1_15/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_15/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_1_15/Component_Function_3/NAND4_in[3] ), .A4(n4592), .ZN(
        \SB2_1_15/buf_output[3] ) );
  NAND3_X2 U11169 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i1[9] ), .A3(
        \SB2_1_15/i0[6] ), .ZN(n4592) );
  NAND4_X2 U11173 ( .A1(\SB1_3_18/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_18/Component_Function_3/NAND4_in[0] ), .A3(n1725), .A4(n4595), 
        .ZN(\SB1_3_18/buf_output[3] ) );
  NAND4_X2 U11175 ( .A1(\SB2_0_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_23/Component_Function_4/NAND4_in[3] ), .A4(n4598), .ZN(
        \SB2_0_23/buf_output[4] ) );
  NAND3_X2 U11176 ( .A1(\SB2_0_23/i0_3 ), .A2(\SB2_0_23/i0[10] ), .A3(
        \SB2_0_23/i0[9] ), .ZN(n4598) );
  XOR2_X1 U11179 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[15] ), .A2(\RI5[1][51] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[141] ) );
  XOR2_X1 U11180 ( .A1(n1544), .A2(n4602), .Z(\MC_ARK_ARC_1_3/buf_output[59] )
         );
  NAND3_X1 U11181 ( .A1(\SB1_2_8/i0_3 ), .A2(\SB1_2_8/i0[8] ), .A3(
        \SB1_2_8/i1_7 ), .ZN(\SB1_2_8/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U11182 ( .A1(\SB1_3_25/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_3_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_25/Component_Function_3/NAND4_in[0] ), .A4(n4603), .ZN(
        \SB1_3_25/buf_output[3] ) );
  NAND3_X2 U11183 ( .A1(\SB1_3_25/i3[0] ), .A2(\SB1_3_25/i0[8] ), .A3(
        \SB1_3_25/i1_5 ), .ZN(n4603) );
  XOR2_X1 U11188 ( .A1(\MC_ARK_ARC_1_0/temp4[22] ), .A2(
        \MC_ARK_ARC_1_0/temp3[22] ), .Z(n4606) );
  XOR2_X1 U11190 ( .A1(n4607), .A2(n4608), .Z(\MC_ARK_ARC_1_0/buf_output[89] )
         );
  XOR2_X1 U11191 ( .A1(\MC_ARK_ARC_1_0/temp1[89] ), .A2(n4667), .Z(n4607) );
  NAND4_X2 U11198 ( .A1(\SB2_0_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_30/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_0_30/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_0_30/buf_output[3] ) );
  NAND3_X1 U11200 ( .A1(\SB4_18/i0_3 ), .A2(\SB4_18/i0[7] ), .A3(\SB4_18/i0_0 ), .ZN(\SB4_18/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U11201 ( .A1(\SB3_21/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_21/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_21/Component_Function_2/NAND4_in[0] ), .A4(
        \SB3_21/Component_Function_2/NAND4_in[3] ), .ZN(\SB4_18/i0_0 ) );
  XOR2_X1 U11202 ( .A1(n4611), .A2(n38), .Z(Ciphertext[30]) );
  XOR2_X1 U11206 ( .A1(\RI5[4][116] ), .A2(\RI5[4][92] ), .Z(n4613) );
  NAND4_X2 U11208 ( .A1(\SB2_4_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_19/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_4_19/Component_Function_2/NAND4_in[1] ), .A4(n4616), .ZN(
        \SB2_4_19/buf_output[2] ) );
  NAND3_X1 U11210 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i0_4 ), .A3(
        \SB1_3_10/i0[10] ), .ZN(\SB1_3_10/Component_Function_0/NAND4_in[2] )
         );
  NAND3_X1 U11211 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i0[10] ), .A3(\SB3_5/i0_4 ), 
        .ZN(\SB3_5/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U11213 ( .A1(\RI5[0][80] ), .A2(\RI5[0][104] ), .Z(n4617) );
  XOR2_X1 U11214 ( .A1(n4618), .A2(n43), .Z(Ciphertext[138]) );
  NAND4_X2 U11215 ( .A1(\SB4_8/Component_Function_0/NAND4_in[1] ), .A2(n1643), 
        .A3(n5110), .A4(n903), .ZN(n4618) );
  NAND4_X2 U11217 ( .A1(\SB2_0_0/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_0/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_0/Component_Function_3/NAND4_in[0] ), .A4(n4620), .ZN(
        \SB2_0_0/buf_output[3] ) );
  XOR2_X1 U11223 ( .A1(\MC_ARK_ARC_1_1/temp4[12] ), .A2(n4623), .Z(
        \MC_ARK_ARC_1_1/temp6[12] ) );
  XOR2_X1 U11224 ( .A1(\RI5[1][78] ), .A2(\RI5[1][114] ), .Z(n4623) );
  NAND4_X2 U11228 ( .A1(\SB1_4_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_4_1/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_4_1/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_4_1/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_4_1/buf_output[1] ) );
  NAND3_X1 U11229 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i1_7 ), .A3(
        \SB2_2_27/i0[8] ), .ZN(\SB2_2_27/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U11230 ( .A1(n315), .A2(\SB1_0_0/i0[6] ), .A3(n380), .ZN(n2810) );
  XOR2_X1 U11232 ( .A1(\MC_ARK_ARC_1_4/temp4[82] ), .A2(n4627), .Z(
        \MC_ARK_ARC_1_4/temp6[82] ) );
  XOR2_X1 U11233 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[184] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[148] ), .Z(n4627) );
  NAND3_X1 U11235 ( .A1(\SB1_4_3/i0[8] ), .A2(\SB1_4_3/i0_4 ), .A3(
        \SB1_4_3/i1_7 ), .ZN(\SB1_4_3/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U11236 ( .A1(\MC_ARK_ARC_1_4/temp2[55] ), .A2(
        \MC_ARK_ARC_1_4/temp1[55] ), .Z(\MC_ARK_ARC_1_4/temp5[55] ) );
  NAND4_X2 U11237 ( .A1(\SB3_18/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_18/Component_Function_5/NAND4_in[2] ), .A3(
        \SB3_18/Component_Function_5/NAND4_in[3] ), .A4(
        \SB3_18/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_18/buf_output[5] ) );
  NAND4_X2 U11238 ( .A1(\SB1_0_29/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_29/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_29/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_29/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_29/buf_output[0] ) );
  XOR2_X1 U11239 ( .A1(\RI5[4][48] ), .A2(\RI5[4][84] ), .Z(
        \MC_ARK_ARC_1_4/temp3[174] ) );
  XOR2_X1 U11240 ( .A1(n4628), .A2(\MC_ARK_ARC_1_3/temp6[22] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[22] ) );
  NAND3_X2 U11242 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i0_0 ), .A3(
        \SB2_3_16/i0_4 ), .ZN(n665) );
  XOR2_X1 U11243 ( .A1(n4630), .A2(n4629), .Z(\MC_ARK_ARC_1_1/temp5[80] ) );
  XOR2_X1 U11244 ( .A1(\RI5[1][26] ), .A2(\RI5[1][80] ), .Z(n4629) );
  NAND3_X2 U11247 ( .A1(\SB2_1_22/i3[0] ), .A2(n6283), .A3(\SB2_1_22/i1_5 ), 
        .ZN(n4631) );
  XOR2_X1 U11249 ( .A1(\RI5[2][104] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[110] ), .Z(n4632) );
  NAND3_X2 U11252 ( .A1(\SB2_1_7/i0_3 ), .A2(\SB2_1_7/i0_4 ), .A3(
        \SB2_1_7/i1[9] ), .ZN(\SB2_1_7/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U11253 ( .A1(n4636), .A2(\MC_ARK_ARC_1_2/temp2[74] ), .Z(
        \MC_ARK_ARC_1_2/temp5[74] ) );
  XOR2_X1 U11254 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[74] ), .Z(n4636) );
  XOR2_X1 U11255 ( .A1(\RI5[2][138] ), .A2(\RI5[2][144] ), .Z(
        \MC_ARK_ARC_1_2/temp1[144] ) );
  XOR2_X1 U11256 ( .A1(\MC_ARK_ARC_1_0/temp5[88] ), .A2(n4637), .Z(
        \MC_ARK_ARC_1_0/buf_output[88] ) );
  XOR2_X1 U11257 ( .A1(\MC_ARK_ARC_1_0/temp3[88] ), .A2(
        \MC_ARK_ARC_1_0/temp4[88] ), .Z(n4637) );
  XOR2_X1 U11258 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[60] ), .A2(\RI5[2][36] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[90] ) );
  NAND3_X1 U11261 ( .A1(\SB1_1_3/i1[9] ), .A2(\MC_ARK_ARC_1_0/buf_output[172] ), .A3(\SB1_1_3/i1_5 ), .ZN(n4640) );
  NAND4_X2 U11263 ( .A1(\SB1_3_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_11/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_11/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_3_11/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_3_11/buf_output[5] ) );
  NAND3_X2 U11264 ( .A1(\SB2_4_30/i0[10] ), .A2(\SB2_4_30/i1_7 ), .A3(
        \SB2_4_30/i1[9] ), .ZN(n2924) );
  NAND3_X2 U11269 ( .A1(\SB2_2_20/i0[6] ), .A2(\SB2_2_20/i0_3 ), .A3(
        \SB2_2_20/i0[10] ), .ZN(n1609) );
  NAND3_X1 U11271 ( .A1(\SB1_4_2/i0[6] ), .A2(\SB1_4_2/i0_3 ), .A3(
        \SB1_4_2/i1[9] ), .ZN(\SB1_4_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U11274 ( .A1(\SB2_1_16/i0_4 ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i0[10] ), .ZN(n4647) );
  XOR2_X1 U11276 ( .A1(n4650), .A2(n4649), .Z(n4657) );
  XOR2_X1 U11277 ( .A1(\RI5[3][122] ), .A2(\RI5[3][14] ), .Z(n4649) );
  NAND3_X2 U11278 ( .A1(\SB2_2_8/i0_3 ), .A2(\SB2_2_8/i0[9] ), .A3(
        \SB2_2_8/i0[8] ), .ZN(n4651) );
  XOR2_X1 U11279 ( .A1(\RI5[2][2] ), .A2(\RI5[2][140] ), .Z(n4652) );
  XOR2_X1 U11282 ( .A1(\MC_ARK_ARC_1_1/temp3[127] ), .A2(
        \MC_ARK_ARC_1_1/temp4[127] ), .Z(n4654) );
  XOR2_X1 U11283 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[44] ), .A2(\RI5[1][20] ), 
        .Z(n2221) );
  NAND4_X2 U11289 ( .A1(n2862), .A2(
        \SB2_0_31/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_0_31/Component_Function_5/NAND4_in[0] ), .A4(n2901), .ZN(
        \SB2_0_31/buf_output[5] ) );
  XOR2_X1 U11290 ( .A1(n4658), .A2(n4659), .Z(\MC_ARK_ARC_1_3/buf_output[36] )
         );
  XOR2_X1 U11291 ( .A1(\MC_ARK_ARC_1_3/temp2[36] ), .A2(
        \MC_ARK_ARC_1_3/temp4[36] ), .Z(n4658) );
  NAND4_X2 U11296 ( .A1(\SB2_0_17/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_0_17/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_0_17/Component_Function_1/NAND4_in[1] ), .A4(n4661), .ZN(
        \SB2_0_17/buf_output[1] ) );
  NAND4_X2 U11300 ( .A1(\SB2_3_10/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_10/Component_Function_0/NAND4_in[0] ), .A4(n4664), .ZN(
        \SB2_3_10/buf_output[0] ) );
  XOR2_X1 U11302 ( .A1(\MC_ARK_ARC_1_1/temp6[110] ), .A2(n4665), .Z(
        \MC_ARK_ARC_1_1/buf_output[110] ) );
  NAND3_X1 U11306 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0[10] ), .A3(
        \SB1_0_18/i0[9] ), .ZN(\SB1_0_18/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U11307 ( .A1(n1163), .A2(
        \SB2_3_31/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_31/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_3_31/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB2_3_31/buf_output[0] ) );
  NAND3_X2 U11308 ( .A1(\SB2_1_16/i0_4 ), .A2(\SB2_1_16/i1_5 ), .A3(
        \SB2_1_16/i0_0 ), .ZN(n5393) );
  XOR2_X1 U11309 ( .A1(\RI5[0][155] ), .A2(n527), .Z(n4667) );
  NAND3_X2 U11312 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0_0 ), .A3(
        \SB1_2_2/buf_output[4] ), .ZN(n4669) );
  INV_X2 U11313 ( .I(\SB1_3_22/buf_output[3] ), .ZN(\SB2_3_20/i0[8] ) );
  XOR2_X1 U11314 ( .A1(\MC_ARK_ARC_1_0/temp3[61] ), .A2(
        \MC_ARK_ARC_1_0/temp4[61] ), .Z(\MC_ARK_ARC_1_0/temp6[61] ) );
  NAND4_X2 U11315 ( .A1(\SB2_4_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_9/Component_Function_1/NAND4_in[3] ), .A4(n4670), .ZN(
        \SB2_4_9/buf_output[1] ) );
  NAND4_X2 U11316 ( .A1(\SB1_0_9/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_3/NAND4_in[0] ), .A4(n1589), .ZN(
        \RI3[0][147] ) );
  NAND4_X2 U11318 ( .A1(\SB1_0_19/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_0_19/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_0_19/Component_Function_3/NAND4_in[1] ), .A4(n4671), .ZN(
        \RI3[0][87] ) );
  NAND4_X2 U11320 ( .A1(\SB2_0_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_10/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_0_10/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_10/buf_output[3] ) );
  NAND4_X2 U11323 ( .A1(n2740), .A2(
        \SB2_0_18/Component_Function_2/NAND4_in[0] ), .A3(n4850), .A4(n982), 
        .ZN(\SB2_0_18/buf_output[2] ) );
  XOR2_X1 U11324 ( .A1(n2555), .A2(\MC_ARK_ARC_1_2/temp3[38] ), .Z(n2120) );
  NAND4_X2 U11325 ( .A1(\SB2_0_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_16/Component_Function_5/NAND4_in[1] ), .A3(n1283), .A4(
        \SB2_0_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_16/buf_output[5] ) );
  NAND4_X2 U11326 ( .A1(\SB2_4_20/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_4_20/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_4_20/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_4_20/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_4_20/buf_output[1] ) );
  NAND4_X2 U11328 ( .A1(\SB1_1_0/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_0/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_1_0/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_1_0/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_0/buf_output[0] ) );
  NAND3_X1 U11331 ( .A1(\SB2_0_17/i0_3 ), .A2(\SB2_0_17/i0[9] ), .A3(
        \SB2_0_17/i0[8] ), .ZN(\SB2_0_17/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U11333 ( .A1(\SB2_1_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_27/Component_Function_1/NAND4_in[3] ), .A4(n4673), .ZN(
        \SB2_1_27/buf_output[1] ) );
  XOR2_X1 U11334 ( .A1(n4674), .A2(\MC_ARK_ARC_1_3/temp5[21] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[21] ) );
  XOR2_X1 U11335 ( .A1(\MC_ARK_ARC_1_3/temp4[21] ), .A2(
        \MC_ARK_ARC_1_3/temp3[21] ), .Z(n4674) );
  XOR2_X1 U11337 ( .A1(n4675), .A2(n1536), .Z(\MC_ARK_ARC_1_3/buf_output[107] ) );
  XOR2_X1 U11338 ( .A1(n4827), .A2(\MC_ARK_ARC_1_3/temp4[107] ), .Z(n4675) );
  NAND3_X2 U11339 ( .A1(\SB2_4_22/i0_0 ), .A2(\SB2_4_22/i1_5 ), .A3(
        \SB2_4_22/i0_4 ), .ZN(n4676) );
  NOR2_X2 U11340 ( .A1(n1592), .A2(n1590), .ZN(n4677) );
  NAND3_X2 U11341 ( .A1(\SB2_4_16/i0_3 ), .A2(\SB2_4_16/i0[10] ), .A3(
        \SB2_4_16/i0[6] ), .ZN(n5012) );
  XOR2_X1 U11342 ( .A1(\RI5[0][190] ), .A2(\RI5[0][166] ), .Z(
        \MC_ARK_ARC_1_0/temp2[28] ) );
  XOR2_X1 U11344 ( .A1(n4678), .A2(n452), .Z(Ciphertext[73]) );
  NOR2_X1 U11345 ( .A1(n4680), .A2(n4679), .ZN(n4678) );
  NAND2_X1 U11347 ( .A1(\SB4_19/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_19/Component_Function_1/NAND4_in[3] ), .ZN(n4680) );
  NAND4_X2 U11348 ( .A1(\SB1_0_31/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_31/Component_Function_3/NAND4_in[3] ), .A3(n4881), .A4(n4681), 
        .ZN(\RI3[0][15] ) );
  NAND3_X2 U11349 ( .A1(\SB1_0_31/i0[10] ), .A2(\SB1_0_31/i1_7 ), .A3(
        \SB1_0_31/i1[9] ), .ZN(n4681) );
  NAND3_X2 U11351 ( .A1(\SB2_3_6/i0_3 ), .A2(\SB2_3_6/i0_0 ), .A3(
        \SB2_3_6/i0_4 ), .ZN(\SB2_3_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11352 ( .A1(\SB1_3_18/i0_3 ), .A2(\SB1_3_18/i0[8] ), .A3(
        \SB1_3_18/i1_7 ), .ZN(\SB1_3_18/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U11353 ( .A1(\SB2_4_8/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_4_8/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_4_8/Component_Function_0/NAND4_in[0] ), .A4(n4684), .ZN(
        \SB2_4_8/buf_output[0] ) );
  NAND3_X1 U11354 ( .A1(\SB1_4_9/i0_0 ), .A2(\SB1_4_9/i1_7 ), .A3(
        \SB1_4_9/i3[0] ), .ZN(n4685) );
  XOR2_X1 U11356 ( .A1(\MC_ARK_ARC_1_3/temp3[63] ), .A2(
        \MC_ARK_ARC_1_3/temp4[63] ), .Z(n4686) );
  NAND4_X2 U11360 ( .A1(\SB1_0_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_24/Component_Function_3/NAND4_in[2] ), .A4(n4689), .ZN(
        \SB1_0_24/buf_output[3] ) );
  NAND3_X2 U11361 ( .A1(\SB1_0_24/i0[8] ), .A2(\SB1_0_24/i1_5 ), .A3(
        \SB1_0_24/i3[0] ), .ZN(n4689) );
  NAND4_X2 U11362 ( .A1(\SB2_1_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_20/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_1_20/Component_Function_4/NAND4_in[1] ), .A4(n4690), .ZN(
        \SB2_1_20/buf_output[4] ) );
  XOR2_X1 U11367 ( .A1(\MC_ARK_ARC_1_0/temp5[158] ), .A2(n4694), .Z(
        \MC_ARK_ARC_1_0/buf_output[158] ) );
  XOR2_X1 U11368 ( .A1(\MC_ARK_ARC_1_0/temp3[158] ), .A2(
        \MC_ARK_ARC_1_0/temp4[158] ), .Z(n4694) );
  NAND4_X2 U11369 ( .A1(n916), .A2(\SB2_3_3/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_3_3/Component_Function_5/NAND4_in[0] ), .A4(n4695), .ZN(
        \SB2_3_3/buf_output[5] ) );
  NAND3_X2 U11370 ( .A1(\SB2_3_3/i0_4 ), .A2(\SB2_3_3/i0[6] ), .A3(
        \SB2_3_3/i0[9] ), .ZN(n4695) );
  XOR2_X1 U11371 ( .A1(n4696), .A2(\MC_ARK_ARC_1_4/temp6[54] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[54] ) );
  XOR2_X1 U11372 ( .A1(\MC_ARK_ARC_1_4/temp2[54] ), .A2(
        \MC_ARK_ARC_1_4/temp1[54] ), .Z(n4696) );
  NAND3_X2 U11373 ( .A1(\SB1_1_15/i0[10] ), .A2(\SB1_1_15/i1[9] ), .A3(
        \SB1_1_15/i1_5 ), .ZN(\SB1_1_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U11374 ( .A1(\SB2_4_23/i0[8] ), .A2(\SB2_4_23/i1_5 ), .A3(
        \SB2_4_23/i3[0] ), .ZN(\SB2_4_23/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U11377 ( .A1(\RI5[4][68] ), .A2(\RI5[4][104] ), .Z(n4698) );
  XOR2_X1 U11378 ( .A1(n4700), .A2(n4699), .Z(\MC_ARK_ARC_1_2/buf_output[50] )
         );
  NAND3_X1 U11384 ( .A1(\SB3_20/i0_3 ), .A2(\SB3_20/i0[8] ), .A3(\SB3_20/i1_7 ), .ZN(\SB3_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U11386 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i1_5 ), .A3(
        \SB4_29/i1[9] ), .ZN(\SB4_29/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U11388 ( .A1(\SB3_22/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_22/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_22/Component_Function_2/NAND4_in[2] ), .A4(n4702), .ZN(
        \SB3_22/buf_output[2] ) );
  NAND3_X1 U11390 ( .A1(\SB4_20/i0[6] ), .A2(\SB4_20/i0[9] ), .A3(
        \SB4_20/i1_5 ), .ZN(\SB4_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U11394 ( .A1(\SB4_19/i0[8] ), .A2(\SB4_19/i3[0] ), .A3(n6273), .ZN(
        \SB4_19/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U11395 ( .A1(\RI5[1][147] ), .A2(\RI5[1][111] ), .Z(
        \MC_ARK_ARC_1_1/temp3[45] ) );
  NAND4_X2 U11396 ( .A1(\SB1_1_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_11/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_1_11/Component_Function_3/NAND4_in[1] ), .A4(n4704), .ZN(
        \SB1_1_11/buf_output[3] ) );
  NAND3_X1 U11397 ( .A1(\SB1_1_11/i0[8] ), .A2(\SB1_1_11/i3[0] ), .A3(
        \SB1_1_11/i1_5 ), .ZN(n4704) );
  XOR2_X1 U11398 ( .A1(\MC_ARK_ARC_1_0/temp1[53] ), .A2(
        \MC_ARK_ARC_1_0/temp2[53] ), .Z(\MC_ARK_ARC_1_0/temp5[53] ) );
  XOR2_X1 U11399 ( .A1(n4705), .A2(\MC_ARK_ARC_1_2/temp2[187] ), .Z(
        \MC_ARK_ARC_1_2/temp5[187] ) );
  XOR2_X1 U11402 ( .A1(n1671), .A2(\MC_ARK_ARC_1_1/temp1[109] ), .Z(n1197) );
  XOR2_X1 U11404 ( .A1(\MC_ARK_ARC_1_4/temp2[64] ), .A2(
        \MC_ARK_ARC_1_4/temp1[64] ), .Z(\MC_ARK_ARC_1_4/temp5[64] ) );
  NAND3_X2 U11405 ( .A1(\SB1_2_19/i0[10] ), .A2(\SB1_2_19/i0_0 ), .A3(
        \SB1_2_19/i0[6] ), .ZN(\SB1_2_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U11408 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i1_7 ), .A3(
        \SB2_1_1/i1[9] ), .ZN(n1861) );
  NAND3_X2 U11410 ( .A1(\SB2_3_20/i0[8] ), .A2(\SB2_3_20/i3[0] ), .A3(n5440), 
        .ZN(\SB2_3_20/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U11413 ( .A1(\MC_ARK_ARC_1_0/temp4[28] ), .A2(n4711), .Z(n2005) );
  XOR2_X1 U11414 ( .A1(\RI5[0][94] ), .A2(\RI5[0][130] ), .Z(n4711) );
  XOR2_X1 U11415 ( .A1(\RI5[1][49] ), .A2(\RI5[1][13] ), .Z(
        \MC_ARK_ARC_1_1/temp3[139] ) );
  NAND2_X2 U11416 ( .A1(n2613), .A2(n2612), .ZN(\RI5[1][13] ) );
  XOR2_X1 U11418 ( .A1(\RI5[1][54] ), .A2(\RI5[1][18] ), .Z(n4712) );
  NAND3_X1 U11420 ( .A1(\SB3_16/i0[10] ), .A2(\SB3_16/i1_7 ), .A3(
        \SB3_16/i1[9] ), .ZN(n4713) );
  XOR2_X1 U11421 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[177] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[21] ), .Z(\MC_ARK_ARC_1_3/temp3[111] )
         );
  XOR2_X1 U11422 ( .A1(n4714), .A2(\MC_ARK_ARC_1_2/temp2[177] ), .Z(
        \MC_ARK_ARC_1_2/temp5[177] ) );
  XOR2_X1 U11423 ( .A1(\RI5[2][177] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[171] ), .Z(n4714) );
  XOR2_X1 U11424 ( .A1(\MC_ARK_ARC_1_1/temp2[168] ), .A2(
        \MC_ARK_ARC_1_1/temp1[168] ), .Z(n4715) );
  XOR2_X1 U11427 ( .A1(\RI5[4][105] ), .A2(\RI5[4][81] ), .Z(n4717) );
  NAND3_X2 U11428 ( .A1(\SB2_3_27/i0[6] ), .A2(\SB2_3_27/i0_4 ), .A3(
        \SB2_3_27/i0[9] ), .ZN(n4718) );
  INV_X2 U11429 ( .I(n4719), .ZN(\MC_ARK_ARC_1_1/buf_output[14] ) );
  NAND3_X2 U11432 ( .A1(\SB2_0_3/i0_0 ), .A2(\SB2_0_3/i1_5 ), .A3(
        \RI3[0][172] ), .ZN(n5211) );
  NAND4_X2 U11435 ( .A1(\SB1_2_5/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_5/Component_Function_3/NAND4_in[3] ), .A3(n2041), .A4(n4722), 
        .ZN(\SB1_2_5/buf_output[3] ) );
  NAND4_X2 U11438 ( .A1(\SB2_0_5/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_5/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_0_5/Component_Function_0/NAND4_in[0] ), .A4(n4724), .ZN(
        \SB2_0_5/buf_output[0] ) );
  NAND3_X1 U11440 ( .A1(\SB1_4_0/i0_0 ), .A2(\MC_ARK_ARC_1_3/buf_output[190] ), 
        .A3(\RI1[4][191] ), .ZN(n4746) );
  NAND3_X1 U11441 ( .A1(\SB1_4_17/i0[10] ), .A2(\SB1_4_17/i0_3 ), .A3(
        \SB1_4_17/i0_4 ), .ZN(\SB1_4_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11444 ( .A1(\SB1_3_26/i0[9] ), .A2(\SB1_3_26/i1_5 ), .A3(
        \SB1_3_26/i0[6] ), .ZN(n4729) );
  NAND4_X2 U11447 ( .A1(\SB2_0_11/Component_Function_5/NAND4_in[2] ), .A2(
        n1854), .A3(n5049), .A4(\SB2_0_11/Component_Function_5/NAND4_in[0] ), 
        .ZN(\SB2_0_11/buf_output[5] ) );
  XOR2_X1 U11448 ( .A1(\MC_ARK_ARC_1_0/temp2[48] ), .A2(
        \MC_ARK_ARC_1_0/temp1[48] ), .Z(\MC_ARK_ARC_1_0/temp5[48] ) );
  XOR2_X1 U11454 ( .A1(\MC_ARK_ARC_1_4/temp5[128] ), .A2(
        \MC_ARK_ARC_1_4/temp6[128] ), .Z(\MC_ARK_ARC_1_4/buf_output[128] ) );
  NAND3_X1 U11456 ( .A1(\SB4_15/i0_0 ), .A2(\SB4_15/i1_7 ), .A3(\SB4_15/i3[0] ), .ZN(n2824) );
  XOR2_X1 U11460 ( .A1(n4737), .A2(\MC_ARK_ARC_1_1/temp5[77] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[77] ) );
  XOR2_X1 U11461 ( .A1(\MC_ARK_ARC_1_1/temp3[77] ), .A2(
        \MC_ARK_ARC_1_1/temp4[77] ), .Z(n4737) );
  NAND4_X2 U11462 ( .A1(\SB2_2_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_19/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_2_19/Component_Function_0/NAND4_in[1] ), .A4(n4738), .ZN(
        \SB2_2_19/buf_output[0] ) );
  XOR2_X1 U11464 ( .A1(\RI5[3][171] ), .A2(\RI5[3][165] ), .Z(n4739) );
  XOR2_X1 U11466 ( .A1(\RI5[2][191] ), .A2(\RI5[2][5] ), .Z(n2335) );
  NAND4_X2 U11467 ( .A1(\SB2_3_26/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_26/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_26/Component_Function_4/NAND4_in[3] ), .A4(n4740), .ZN(
        \SB2_3_26/buf_output[4] ) );
  XOR2_X1 U11471 ( .A1(\MC_ARK_ARC_1_1/temp3[91] ), .A2(
        \MC_ARK_ARC_1_1/temp4[91] ), .Z(n4743) );
  NAND4_X2 U11473 ( .A1(n2389), .A2(
        \SB2_2_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_16/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_16/buf_output[5] ) );
  NAND3_X1 U11474 ( .A1(\SB4_1/i0[6] ), .A2(\SB4_1/i0[8] ), .A3(\SB4_1/i0[7] ), 
        .ZN(\SB4_1/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U11475 ( .A1(\MC_ARK_ARC_1_1/temp5[122] ), .A2(n4745), .Z(
        \MC_ARK_ARC_1_1/buf_output[122] ) );
  XOR2_X1 U11478 ( .A1(\MC_ARK_ARC_1_1/temp1[43] ), .A2(
        \MC_ARK_ARC_1_1/temp2[43] ), .Z(n4747) );
  XOR2_X1 U11481 ( .A1(\MC_ARK_ARC_1_3/temp5[83] ), .A2(n4750), .Z(
        \MC_ARK_ARC_1_3/buf_output[83] ) );
  XOR2_X1 U11482 ( .A1(\RI5[4][103] ), .A2(\RI5[4][67] ), .Z(
        \MC_ARK_ARC_1_4/temp3[1] ) );
  NAND4_X2 U11486 ( .A1(\SB1_1_13/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_1_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_13/buf_output[0] ) );
  NAND4_X2 U11487 ( .A1(\SB2_0_12/Component_Function_2/NAND4_in[2] ), .A2(
        n5163), .A3(n4755), .A4(n4754), .ZN(\SB2_0_12/buf_output[2] ) );
  NAND3_X2 U11488 ( .A1(\SB2_0_12/i1_5 ), .A2(\SB2_0_12/i0_0 ), .A3(
        \RI3[0][118] ), .ZN(n4754) );
  NAND3_X2 U11489 ( .A1(\SB2_0_12/i1_5 ), .A2(\SB2_0_12/i0[10] ), .A3(
        \SB2_0_12/i1[9] ), .ZN(n4755) );
  XOR2_X1 U11491 ( .A1(\RI5[3][11] ), .A2(\RI5[3][173] ), .Z(n2760) );
  NAND4_X2 U11494 ( .A1(\SB1_4_22/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_4_22/Component_Function_0/NAND4_in[2] ), .A3(n2025), .A4(
        \SB1_4_22/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_4_22/buf_output[0] ) );
  NAND4_X2 U11495 ( .A1(\SB3_20/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_20/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_20/Component_Function_4/NAND4_in[3] ), .A4(n4759), .ZN(
        \SB3_20/buf_output[4] ) );
  NAND4_X2 U11496 ( .A1(\SB1_1_28/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_28/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_1_28/Component_Function_2/NAND4_in[3] ), .A4(n4761), .ZN(
        \SB1_1_28/buf_output[2] ) );
  NAND3_X2 U11497 ( .A1(\SB1_1_28/i0[10] ), .A2(\SB1_1_28/i1[9] ), .A3(
        \SB1_1_28/i1_5 ), .ZN(n4761) );
  NAND4_X2 U11499 ( .A1(\SB1_1_7/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_7/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_7/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_1_7/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_7/buf_output[1] ) );
  NAND4_X2 U11501 ( .A1(\SB1_4_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_24/Component_Function_0/NAND4_in[0] ), .A4(n4764), .ZN(
        \SB1_4_24/buf_output[0] ) );
  XOR2_X1 U11502 ( .A1(n4765), .A2(n30), .Z(Ciphertext[6]) );
  XOR2_X1 U11504 ( .A1(n4767), .A2(n4766), .Z(\MC_ARK_ARC_1_3/temp6[166] ) );
  XOR2_X1 U11505 ( .A1(\RI5[3][76] ), .A2(n38), .Z(n4766) );
  NAND3_X2 U11507 ( .A1(\SB2_3_2/i0_3 ), .A2(\SB2_3_2/i0_4 ), .A3(
        \SB2_3_2/i1[9] ), .ZN(n4768) );
  NAND4_X2 U11508 ( .A1(\SB2_3_11/Component_Function_2/NAND4_in[2] ), .A2(
        n1698), .A3(n5013), .A4(n4769), .ZN(\SB2_3_11/buf_output[2] ) );
  NAND3_X2 U11509 ( .A1(\SB2_3_11/i0[10] ), .A2(\SB2_3_11/i1_5 ), .A3(
        \SB2_3_11/i1[9] ), .ZN(n4769) );
  XOR2_X1 U11510 ( .A1(n5242), .A2(\MC_ARK_ARC_1_0/temp4[95] ), .Z(
        \MC_ARK_ARC_1_0/temp6[95] ) );
  XOR2_X1 U11512 ( .A1(n4771), .A2(\MC_ARK_ARC_1_3/temp6[126] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[126] ) );
  XOR2_X1 U11513 ( .A1(\MC_ARK_ARC_1_3/temp1[126] ), .A2(
        \MC_ARK_ARC_1_3/temp2[126] ), .Z(n4771) );
  XOR2_X1 U11514 ( .A1(\MC_ARK_ARC_1_2/temp2[165] ), .A2(
        \MC_ARK_ARC_1_2/temp1[165] ), .Z(\MC_ARK_ARC_1_2/temp5[165] ) );
  XOR2_X1 U11515 ( .A1(n4772), .A2(n2049), .Z(\MC_ARK_ARC_1_0/buf_output[164] ) );
  XOR2_X1 U11516 ( .A1(\MC_ARK_ARC_1_3/temp3[118] ), .A2(n4774), .Z(n1189) );
  XOR2_X1 U11517 ( .A1(\RI5[3][64] ), .A2(\RI5[3][88] ), .Z(n4774) );
  XOR2_X1 U11518 ( .A1(n4775), .A2(\MC_ARK_ARC_1_2/temp5[54] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[54] ) );
  XOR2_X1 U11519 ( .A1(\MC_ARK_ARC_1_2/temp4[54] ), .A2(n2031), .Z(n4775) );
  NAND3_X2 U11521 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0[9] ), .A3(
        \SB2_0_21/i0[8] ), .ZN(\SB2_0_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11524 ( .A1(\SB2_1_2/i0_4 ), .A2(\SB2_1_2/i1_7 ), .A3(
        \SB2_1_2/i0[8] ), .ZN(n1694) );
  NAND4_X2 U11526 ( .A1(\SB1_0_7/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_7/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_7/Component_Function_5/NAND4_in[0] ), .A4(n4780), .ZN(
        \RI3[0][149] ) );
  NAND3_X2 U11527 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB1_2_2/buf_output[4] ), .A3(
        \SB2_2_1/i1[9] ), .ZN(\SB2_2_1/Component_Function_5/NAND4_in[2] ) );
  NOR2_X1 U11528 ( .A1(\MC_ARK_ARC_1_3/buf_output[36] ), .A2(
        \MC_ARK_ARC_1_3/buf_output[37] ), .ZN(n5117) );
  NAND4_X2 U11529 ( .A1(\SB4_0/Component_Function_0/NAND4_in[2] ), .A2(n2966), 
        .A3(\SB4_0/Component_Function_0/NAND4_in[1] ), .A4(n4801), .ZN(n2781)
         );
  XOR2_X1 U11533 ( .A1(n2191), .A2(n5200), .Z(\MC_ARK_ARC_1_4/buf_output[17] )
         );
  NAND3_X2 U11534 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i0_0 ), .A3(
        \SB2_2_15/i0_4 ), .ZN(\SB2_2_15/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U11535 ( .A1(\SB2_3_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_27/Component_Function_2/NAND4_in[1] ), .A3(n706), .A4(
        \SB2_3_27/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_3_27/buf_output[2] ) );
  XOR2_X1 U11536 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[77] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[71] ), .Z(\MC_ARK_ARC_1_0/temp1[77] ) );
  NAND3_X2 U11537 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0[10] ), .A3(
        \SB2_0_21/i0[9] ), .ZN(n4781) );
  NAND3_X1 U11538 ( .A1(\SB3_27/i0_3 ), .A2(\SB3_27/i1_7 ), .A3(\SB3_27/i0[8] ), .ZN(\SB3_27/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U11539 ( .A1(\MC_ARK_ARC_1_0/temp5[77] ), .A2(
        \MC_ARK_ARC_1_0/temp6[77] ), .Z(\MC_ARK_ARC_1_0/buf_output[77] ) );
  NAND3_X1 U11540 ( .A1(\SB2_3_20/i0[6] ), .A2(\SB2_3_20/i0[9] ), .A3(n5440), 
        .ZN(\SB2_3_20/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U11541 ( .A1(n4878), .A2(
        \SB2_4_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_25/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_4_25/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_4_25/buf_output[1] ) );
  NAND3_X1 U11544 ( .A1(\SB2_4_11/i0_4 ), .A2(\SB2_4_11/i1_7 ), .A3(
        \SB2_4_11/i0[8] ), .ZN(n4782) );
  NAND4_X2 U11548 ( .A1(\SB1_4_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_12/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_4_12/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_4_12/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_4_12/buf_output[0] ) );
  NAND4_X2 U11549 ( .A1(\SB2_3_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_20/Component_Function_4/NAND4_in[1] ), .A3(n2424), .A4(n4785), 
        .ZN(\SB2_3_20/buf_output[4] ) );
  NAND3_X2 U11550 ( .A1(\RI3[3][70] ), .A2(n5440), .A3(\SB2_3_20/i1[9] ), .ZN(
        n4785) );
  NAND3_X1 U11552 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i0[10] ), .A3(
        \SB1_0_23/i0_4 ), .ZN(\SB1_0_23/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U11556 ( .A1(\RI5[4][96] ), .A2(\RI5[4][90] ), .Z(
        \MC_ARK_ARC_1_4/temp1[96] ) );
  NAND3_X1 U11557 ( .A1(n6552), .A2(\SB2_3_29/i0_3 ), .A3(\SB2_3_29/i0[10] ), 
        .ZN(\SB2_3_29/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U11560 ( .A1(n4790), .A2(n120), .Z(Ciphertext[33]) );
  XOR2_X1 U11564 ( .A1(\MC_ARK_ARC_1_4/temp4[7] ), .A2(
        \MC_ARK_ARC_1_4/temp3[7] ), .Z(n1599) );
  NAND3_X1 U11569 ( .A1(\SB3_15/i3[0] ), .A2(\SB3_15/i0[8] ), .A3(
        \SB3_15/i1_5 ), .ZN(\SB3_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U11570 ( .A1(\SB2_4_13/i0_4 ), .A2(\SB2_4_13/i1_5 ), .A3(
        \SB2_4_13/i1[9] ), .ZN(n1850) );
  NAND4_X2 U11571 ( .A1(\SB1_0_23/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_23/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_23/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][63] ) );
  NAND4_X2 U11572 ( .A1(\SB2_3_10/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_10/Component_Function_4/NAND4_in[0] ), .A3(n4795), .A4(n4794), 
        .ZN(\SB2_3_10/buf_output[4] ) );
  NAND3_X1 U11574 ( .A1(\SB2_3_10/i0_0 ), .A2(\SB2_3_10/i1_7 ), .A3(
        \SB2_3_10/i3[0] ), .ZN(n4795) );
  NAND3_X1 U11575 ( .A1(\SB1_4_24/i0_0 ), .A2(\SB1_4_24/i0[9] ), .A3(
        \SB1_4_24/i0[8] ), .ZN(n4796) );
  XOR2_X1 U11576 ( .A1(n4798), .A2(n4797), .Z(\MC_ARK_ARC_1_4/buf_output[56] )
         );
  XOR2_X1 U11577 ( .A1(n2324), .A2(\MC_ARK_ARC_1_4/temp4[56] ), .Z(n4797) );
  XOR2_X1 U11579 ( .A1(\RI5[3][67] ), .A2(\RI5[3][73] ), .Z(n4799) );
  XOR2_X1 U11581 ( .A1(n750), .A2(n5153), .Z(n4800) );
  XOR2_X1 U11585 ( .A1(\MC_ARK_ARC_1_4/temp1[0] ), .A2(n4805), .Z(
        \MC_ARK_ARC_1_4/temp5[0] ) );
  XOR2_X1 U11586 ( .A1(\RI5[4][138] ), .A2(\RI5[4][162] ), .Z(n4805) );
  NAND3_X1 U11587 ( .A1(\SB4_22/i0[10] ), .A2(\SB4_22/i1_5 ), .A3(
        \SB4_22/i1[9] ), .ZN(n4806) );
  XOR2_X1 U11590 ( .A1(n4809), .A2(n197), .Z(Ciphertext[79]) );
  NAND4_X2 U11591 ( .A1(\SB4_18/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_18/Component_Function_1/NAND4_in[3] ), .A4(
        \SB4_18/Component_Function_1/NAND4_in[0] ), .ZN(n4809) );
  XOR2_X1 U11594 ( .A1(\MC_ARK_ARC_1_4/temp5[21] ), .A2(n4812), .Z(
        \MC_ARK_ARC_1_4/buf_output[21] ) );
  NAND3_X2 U11597 ( .A1(\RI3[0][52] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i1[9] ), .ZN(n4814) );
  NAND3_X2 U11600 ( .A1(\SB1_1_26/i0_4 ), .A2(\SB1_1_26/i0_0 ), .A3(
        \SB1_1_26/i1_5 ), .ZN(n4816) );
  NAND4_X2 U11601 ( .A1(\SB2_0_19/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_19/Component_Function_4/NAND4_in[0] ), .A3(n2254), .A4(n4817), 
        .ZN(\SB2_0_19/buf_output[4] ) );
  NAND3_X1 U11603 ( .A1(\SB4_0/i0[6] ), .A2(\SB3_5/buf_output[0] ), .A3(
        \SB4_0/i1_5 ), .ZN(n4818) );
  XOR2_X1 U11604 ( .A1(\RI5[1][147] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[141] ), .Z(n4820) );
  XOR2_X1 U11605 ( .A1(\MC_ARK_ARC_1_0/temp1[24] ), .A2(
        \MC_ARK_ARC_1_0/temp2[24] ), .Z(n1576) );
  XOR2_X1 U11606 ( .A1(n4822), .A2(n4821), .Z(\MC_ARK_ARC_1_0/buf_output[188] ) );
  XOR2_X1 U11607 ( .A1(\MC_ARK_ARC_1_0/temp1[188] ), .A2(
        \MC_ARK_ARC_1_0/temp4[188] ), .Z(n4821) );
  XOR2_X1 U11608 ( .A1(n4823), .A2(\MC_ARK_ARC_1_1/temp1[8] ), .Z(
        \MC_ARK_ARC_1_1/temp5[8] ) );
  XOR2_X1 U11609 ( .A1(\RI5[1][170] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[146] ), .Z(n4823) );
  XOR2_X1 U11611 ( .A1(n4825), .A2(\MC_ARK_ARC_1_0/temp2[43] ), .Z(
        \MC_ARK_ARC_1_0/temp5[43] ) );
  XOR2_X1 U11612 ( .A1(\RI5[0][37] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[43] ), 
        .Z(n4825) );
  NAND3_X2 U11615 ( .A1(\SB2_3_6/i0_4 ), .A2(\SB2_3_6/i1_5 ), .A3(
        \SB2_3_6/i0_0 ), .ZN(n4922) );
  XOR2_X1 U11616 ( .A1(\RI5[3][17] ), .A2(\RI5[3][173] ), .Z(n4827) );
  NAND4_X2 U11617 ( .A1(\SB1_4_31/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_31/Component_Function_0/NAND4_in[0] ), .A4(n4828), .ZN(
        \SB1_4_31/buf_output[0] ) );
  NAND4_X2 U11619 ( .A1(\SB2_3_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_20/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_3_20/Component_Function_2/NAND4_in[1] ), .A4(n4829), .ZN(
        \SB2_3_20/buf_output[2] ) );
  NAND3_X2 U11620 ( .A1(\SB2_3_20/i0_0 ), .A2(\RI3[3][70] ), .A3(n5440), .ZN(
        n4829) );
  NAND3_X1 U11622 ( .A1(\SB1_3_20/i0_4 ), .A2(\SB1_3_20/i1[9] ), .A3(
        \SB1_3_20/i1_5 ), .ZN(\SB1_3_20/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U11629 ( .A1(\RI5[3][74] ), .A2(\RI5[3][50] ), .Z(
        \MC_ARK_ARC_1_3/temp2[104] ) );
  NAND3_X1 U11633 ( .A1(\SB2_0_27/i3[0] ), .A2(\SB2_0_27/i0[8] ), .A3(
        \SB2_0_27/i1_5 ), .ZN(\SB2_0_27/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U11637 ( .A1(\RI5[0][39] ), .A2(\RI5[0][45] ), .Z(
        \MC_ARK_ARC_1_0/temp1[45] ) );
  NAND3_X2 U11638 ( .A1(\SB2_3_19/i0[6] ), .A2(\SB2_3_19/i1_5 ), .A3(
        \SB2_3_19/i0[9] ), .ZN(n4837) );
  XOR2_X1 U11640 ( .A1(\RI5[0][87] ), .A2(\RI5[0][51] ), .Z(
        \MC_ARK_ARC_1_0/temp3[177] ) );
  NAND3_X2 U11641 ( .A1(\SB1_0_27/i0[10] ), .A2(\SB1_0_27/i0[6] ), .A3(
        \SB1_0_27/i0_0 ), .ZN(n4839) );
  NAND4_X2 U11646 ( .A1(\SB1_3_4/Component_Function_5/NAND4_in[1] ), .A2(n1361), .A3(n643), .A4(\SB1_3_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_4/buf_output[5] ) );
  NAND3_X2 U11650 ( .A1(\SB2_2_22/i0_0 ), .A2(\SB2_2_22/i1_5 ), .A3(
        \SB2_2_22/i0_4 ), .ZN(\SB2_2_22/Component_Function_2/NAND4_in[3] ) );
  BUF_X2 U11654 ( .I(\SB2_0_9/i3[0] ), .Z(n4847) );
  NAND4_X2 U11656 ( .A1(\SB2_4_19/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_4_19/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_4_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_19/Component_Function_1/NAND4_in[1] ), .ZN(
        \SB2_4_19/buf_output[1] ) );
  XOR2_X1 U11659 ( .A1(\RI5[0][24] ), .A2(\RI5[0][30] ), .Z(n4849) );
  NAND3_X1 U11661 ( .A1(\SB2_0_18/i0_0 ), .A2(\SB2_0_18/i1_5 ), .A3(
        \RI3[0][82] ), .ZN(n4850) );
  NAND3_X1 U11662 ( .A1(\SB1_3_7/i0[10] ), .A2(\SB1_3_7/i1_5 ), .A3(
        \SB1_3_7/i1[9] ), .ZN(\SB1_3_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U11663 ( .A1(\SB1_2_7/i0[10] ), .A2(\SB1_2_7/i0[6] ), .A3(
        \SB1_2_7/i0_0 ), .ZN(\SB1_2_7/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U11667 ( .A1(\SB1_1_18/i0_3 ), .A2(\SB1_1_18/i0_4 ), .A3(
        \SB1_1_18/i1[9] ), .ZN(n4852) );
  XOR2_X1 U11668 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[64] ), .A2(\RI5[4][70] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[70] ) );
  XOR2_X1 U11669 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[64] ), .A2(\RI5[4][100] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[190] ) );
  INV_X2 U11670 ( .I(\SB1_1_18/buf_output[2] ), .ZN(\SB2_1_15/i1[9] ) );
  NAND3_X2 U11672 ( .A1(\SB1_3_28/i0[10] ), .A2(\SB1_3_28/i0[6] ), .A3(
        \SB1_3_28/i0_0 ), .ZN(\SB1_3_28/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U11673 ( .A1(\RI5[3][64] ), .A2(\RI5[3][100] ), .Z(
        \MC_ARK_ARC_1_3/temp3[190] ) );
  NAND3_X2 U11675 ( .A1(\SB2_2_20/i0[6] ), .A2(\SB2_2_20/i0[10] ), .A3(
        \SB2_2_20/i0_0 ), .ZN(\SB2_2_20/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U11676 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[44] ), .A2(\RI5[1][68] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[98] ) );
  NAND2_X2 U11677 ( .A1(\SB2_3_16/i0_0 ), .A2(\SB2_3_16/i3[0] ), .ZN(n4853) );
  INV_X2 U11679 ( .I(\SB3_3/buf_output[2] ), .ZN(\SB4_0/i1[9] ) );
  XOR2_X1 U11682 ( .A1(\MC_ARK_ARC_1_4/temp3[112] ), .A2(
        \MC_ARK_ARC_1_4/temp4[112] ), .Z(\MC_ARK_ARC_1_4/temp6[112] ) );
  NAND3_X1 U11683 ( .A1(\SB2_3_4/i0_4 ), .A2(\SB2_3_4/i1_7 ), .A3(
        \SB2_3_4/i0[8] ), .ZN(\SB2_3_4/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U11684 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[93] ), .A2(\RI5[4][57] ), 
        .Z(n4857) );
  NAND4_X2 U11687 ( .A1(\SB2_3_22/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_22/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_3_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_22/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_22/buf_output[1] ) );
  XOR2_X1 U11688 ( .A1(\RI5[0][26] ), .A2(\RI5[0][2] ), .Z(
        \MC_ARK_ARC_1_0/temp2[56] ) );
  NAND3_X1 U11689 ( .A1(\SB1_1_31/i0[10] ), .A2(\SB1_1_31/i0_3 ), .A3(
        \SB1_1_31/i0[6] ), .ZN(\SB1_1_31/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U11690 ( .A1(\MC_ARK_ARC_1_1/temp5[146] ), .A2(n4859), .Z(
        \MC_ARK_ARC_1_1/buf_output[146] ) );
  XOR2_X1 U11691 ( .A1(\MC_ARK_ARC_1_1/temp3[146] ), .A2(
        \MC_ARK_ARC_1_1/temp4[146] ), .Z(n4859) );
  NAND3_X1 U11694 ( .A1(\SB1_3_3/i0[10] ), .A2(\SB1_3_3/i0_0 ), .A3(
        \SB1_3_3/i0[6] ), .ZN(\SB1_3_3/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U11696 ( .A1(\SB4_6/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_6/Component_Function_4/NAND4_in[0] ), .A3(
        \SB4_6/Component_Function_4/NAND4_in[3] ), .A4(n4861), .ZN(n5279) );
  NAND3_X1 U11699 ( .A1(\SB1_3_16/i0[10] ), .A2(\SB1_3_16/i0_3 ), .A3(
        \MC_ARK_ARC_1_2/buf_output[90] ), .ZN(
        \SB1_3_16/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U11700 ( .A1(\MC_ARK_ARC_1_2/temp5[90] ), .A2(
        \MC_ARK_ARC_1_2/temp6[90] ), .Z(\MC_ARK_ARC_1_2/buf_output[90] ) );
  XOR2_X1 U11705 ( .A1(\RI5[4][34] ), .A2(\RI5[4][58] ), .Z(
        \MC_ARK_ARC_1_4/temp2[88] ) );
  XOR2_X1 U11706 ( .A1(n4868), .A2(\MC_ARK_ARC_1_4/temp5[160] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[160] ) );
  XOR2_X1 U11707 ( .A1(\MC_ARK_ARC_1_4/temp3[160] ), .A2(
        \MC_ARK_ARC_1_4/temp4[160] ), .Z(n4868) );
  XOR2_X1 U11709 ( .A1(n4869), .A2(\MC_ARK_ARC_1_4/temp4[38] ), .Z(
        \MC_ARK_ARC_1_4/temp6[38] ) );
  XOR2_X1 U11714 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[115] ), .A2(\RI5[2][109] ), .Z(n4872) );
  NAND4_X2 U11719 ( .A1(\SB3_14/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_14/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_14/Component_Function_4/NAND4_in[3] ), .A4(n4875), .ZN(
        \SB3_14/buf_output[4] ) );
  NAND3_X2 U11720 ( .A1(\RI3[0][112] ), .A2(\SB2_0_13/i0[9] ), .A3(
        \SB2_0_13/i0[6] ), .ZN(n2180) );
  XOR2_X1 U11721 ( .A1(\RI5[1][2] ), .A2(\RI5[1][158] ), .Z(
        \MC_ARK_ARC_1_1/temp3[92] ) );
  NAND3_X2 U11722 ( .A1(\SB2_2_31/i0_3 ), .A2(\SB2_2_31/i0_4 ), .A3(
        \SB2_2_31/i1[9] ), .ZN(n3131) );
  NAND4_X2 U11723 ( .A1(\SB3_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_13/Component_Function_5/NAND4_in[0] ), .A4(n4876), .ZN(
        \SB3_13/buf_output[5] ) );
  NAND3_X2 U11724 ( .A1(\SB3_13/i0[9] ), .A2(\SB3_13/i0[6] ), .A3(
        \SB3_13/i0_4 ), .ZN(n4876) );
  NAND3_X1 U11727 ( .A1(\SB4_0/i0_3 ), .A2(\SB4_0/i0_4 ), .A3(\SB4_0/i0[10] ), 
        .ZN(\SB4_0/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U11728 ( .A1(n4879), .A2(n73), .Z(Ciphertext[21]) );
  XOR2_X1 U11731 ( .A1(\MC_ARK_ARC_1_3/temp3[28] ), .A2(
        \MC_ARK_ARC_1_3/temp4[28] ), .Z(\MC_ARK_ARC_1_3/temp6[28] ) );
  NAND4_X2 U11733 ( .A1(\SB2_1_4/Component_Function_5/NAND4_in[2] ), .A2(n809), 
        .A3(\SB2_1_4/Component_Function_5/NAND4_in[3] ), .A4(n2104), .ZN(
        \SB2_1_4/buf_output[5] ) );
  INV_X2 U11734 ( .I(\SB1_3_14/buf_output[2] ), .ZN(\SB2_3_11/i1[9] ) );
  XOR2_X1 U11735 ( .A1(n1078), .A2(\MC_ARK_ARC_1_3/temp4[177] ), .Z(n1391) );
  NAND3_X2 U11737 ( .A1(\SB2_2_1/i0[10] ), .A2(\SB2_2_1/i0[6] ), .A3(
        \SB2_2_1/i0_3 ), .ZN(\SB2_2_1/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U11739 ( .A1(\MC_ARK_ARC_1_3/temp1[181] ), .A2(n5062), .Z(
        \MC_ARK_ARC_1_3/temp5[181] ) );
  XOR2_X1 U11740 ( .A1(\MC_ARK_ARC_1_0/temp6[52] ), .A2(n4882), .Z(
        \MC_ARK_ARC_1_0/buf_output[52] ) );
  NAND2_X2 U11742 ( .A1(\SB1_4_12/i1_5 ), .A2(n4883), .ZN(
        \SB1_4_12/Component_Function_3/NAND4_in[3] ) );
  NOR2_X1 U11743 ( .A1(\MC_ARK_ARC_1_3/buf_output[114] ), .A2(n3975), .ZN(
        n4883) );
  NAND3_X1 U11747 ( .A1(\SB1_3_11/i0[9] ), .A2(\SB1_3_11/i0[6] ), .A3(
        \SB1_3_11/i1_5 ), .ZN(n4885) );
  NAND3_X2 U11748 ( .A1(\SB2_1_26/i0[10] ), .A2(\SB2_1_26/i0_0 ), .A3(
        \SB2_1_26/i0[6] ), .ZN(\SB2_1_26/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U11749 ( .A1(\SB4_22/i0_4 ), .A2(\SB4_22/i0_0 ), .A3(\SB4_22/i1_5 ), 
        .ZN(n4886) );
  XOR2_X1 U11752 ( .A1(\RI5[0][190] ), .A2(\RI5[0][184] ), .Z(
        \MC_ARK_ARC_1_0/temp1[190] ) );
  XOR2_X1 U11754 ( .A1(n2037), .A2(n5169), .Z(\MC_ARK_ARC_1_4/temp5[32] ) );
  NAND3_X2 U11755 ( .A1(\SB4_16/i0_4 ), .A2(\SB4_16/i0[9] ), .A3(
        \SB4_16/i0[6] ), .ZN(\SB4_16/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U11758 ( .A1(\MC_ARK_ARC_1_4/temp3[32] ), .A2(
        \MC_ARK_ARC_1_4/temp4[32] ), .Z(\MC_ARK_ARC_1_4/temp6[32] ) );
  NAND3_X1 U11760 ( .A1(\SB2_0_14/i0_0 ), .A2(\SB2_0_14/i0_4 ), .A3(
        \SB2_0_14/i1_5 ), .ZN(n4889) );
  NAND3_X1 U11763 ( .A1(\SB1_4_15/i0[8] ), .A2(\SB1_4_15/i1_5 ), .A3(
        \SB1_4_15/i3[0] ), .ZN(n2121) );
  XOR2_X1 U11764 ( .A1(n4891), .A2(\MC_ARK_ARC_1_2/temp4[28] ), .Z(
        \MC_ARK_ARC_1_2/temp6[28] ) );
  XOR2_X1 U11765 ( .A1(\RI5[2][94] ), .A2(\RI5[2][130] ), .Z(n4891) );
  XOR2_X1 U11767 ( .A1(n4893), .A2(\MC_ARK_ARC_1_0/temp4[63] ), .Z(
        \MC_ARK_ARC_1_0/temp6[63] ) );
  NAND3_X1 U11774 ( .A1(\SB2_0_31/i0_0 ), .A2(\SB2_0_31/i0[10] ), .A3(
        \SB2_0_31/i0[6] ), .ZN(n2862) );
  XOR2_X1 U11775 ( .A1(n1931), .A2(n3113), .Z(\MC_ARK_ARC_1_3/buf_output[170] ) );
  XOR2_X1 U11776 ( .A1(\MC_ARK_ARC_1_1/temp5[129] ), .A2(
        \MC_ARK_ARC_1_1/temp6[129] ), .Z(\MC_ARK_ARC_1_1/buf_output[129] ) );
  INV_X1 U11779 ( .I(\SB3_9/buf_output[5] ), .ZN(\SB4_9/i1_5 ) );
  NAND4_X2 U11780 ( .A1(\SB3_9/Component_Function_5/NAND4_in[1] ), .A2(n1327), 
        .A3(n3038), .A4(\SB3_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_9/buf_output[5] ) );
  NAND4_X2 U11786 ( .A1(\SB2_1_4/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_4/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_4/Component_Function_0/NAND4_in[0] ), .A4(n4898), .ZN(
        \SB2_1_4/buf_output[0] ) );
  NAND3_X1 U11787 ( .A1(\SB2_4_29/i0_3 ), .A2(\SB2_4_29/i0[10] ), .A3(
        \SB2_4_29/i0_4 ), .ZN(\SB2_4_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11790 ( .A1(\SB2_0_13/i0_3 ), .A2(\SB2_0_13/i1[9] ), .A3(
        \SB2_0_13/i0[6] ), .ZN(\SB2_0_13/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U11792 ( .A1(\SB1_1_6/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_1_6/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_6/Component_Function_4/NAND4_in[1] ), .A4(n4899), .ZN(
        \SB1_1_6/buf_output[4] ) );
  NAND3_X1 U11794 ( .A1(n5450), .A2(\SB2_0_31/i0[8] ), .A3(\SB2_0_31/i1_5 ), 
        .ZN(n5066) );
  NAND4_X2 U11796 ( .A1(n2185), .A2(n5336), .A3(n1400), .A4(n4902), .ZN(
        \SB2_1_18/buf_output[5] ) );
  NAND3_X2 U11797 ( .A1(\SB2_1_18/i0[6] ), .A2(\SB2_1_18/i0_4 ), .A3(
        \SB2_1_18/i0[9] ), .ZN(n4902) );
  XOR2_X1 U11798 ( .A1(n2933), .A2(n4903), .Z(\MC_ARK_ARC_1_4/buf_output[87] )
         );
  XOR2_X1 U11799 ( .A1(n1384), .A2(n5162), .Z(n4903) );
  NAND3_X1 U11801 ( .A1(\SB2_3_20/i0_0 ), .A2(\SB2_3_20/i3[0] ), .A3(
        \SB2_3_20/i1_7 ), .ZN(\SB2_3_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U11802 ( .A1(\SB2_1_5/i0_4 ), .A2(\SB2_1_5/i0[9] ), .A3(
        \SB2_1_5/i0[6] ), .ZN(n758) );
  NAND3_X1 U11805 ( .A1(\SB1_2_21/i0_4 ), .A2(\SB1_2_21/i1[9] ), .A3(
        \SB1_2_21/i1_5 ), .ZN(\SB1_2_21/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U11806 ( .A1(n4906), .A2(\MC_ARK_ARC_1_3/temp5[51] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[51] ) );
  XOR2_X1 U11807 ( .A1(\MC_ARK_ARC_1_3/temp3[51] ), .A2(
        \MC_ARK_ARC_1_3/temp4[51] ), .Z(n4906) );
  NAND4_X2 U11808 ( .A1(\SB2_1_5/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_5/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_1_5/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_1_5/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_1_5/buf_output[4] ) );
  XOR2_X1 U11811 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[21] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[177] ), .Z(\MC_ARK_ARC_1_1/temp3[111] )
         );
  INV_X2 U11815 ( .I(\SB1_1_22/buf_output[2] ), .ZN(\SB2_1_19/i1[9] ) );
  XOR2_X1 U11816 ( .A1(n4914), .A2(\MC_ARK_ARC_1_4/temp1[71] ), .Z(
        \MC_ARK_ARC_1_4/temp5[71] ) );
  XOR2_X1 U11818 ( .A1(\MC_ARK_ARC_1_2/temp3[7] ), .A2(
        \MC_ARK_ARC_1_2/temp4[7] ), .Z(n4915) );
  XOR2_X1 U11819 ( .A1(\RI5[1][31] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[121] ) );
  NAND3_X1 U11820 ( .A1(\SB4_11/i0_3 ), .A2(\SB4_11/i0_4 ), .A3(\SB4_11/i1[9] ), .ZN(\SB4_11/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U11821 ( .A1(n1879), .A2(n4916), .Z(\MC_ARK_ARC_1_3/buf_output[125] ) );
  XOR2_X1 U11822 ( .A1(\MC_ARK_ARC_1_3/temp1[125] ), .A2(
        \MC_ARK_ARC_1_3/temp2[125] ), .Z(n4916) );
  NAND3_X1 U11823 ( .A1(\SB1_2_8/i0[8] ), .A2(\SB1_2_8/i0_3 ), .A3(
        \SB1_2_8/i0[9] ), .ZN(\SB1_2_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11825 ( .A1(\SB4_1/i0[10] ), .A2(\SB4_1/i0_3 ), .A3(\SB4_1/i0[9] ), 
        .ZN(n4919) );
  XOR2_X1 U11826 ( .A1(\MC_ARK_ARC_1_3/temp2[87] ), .A2(
        \MC_ARK_ARC_1_3/temp1[87] ), .Z(n4921) );
  NAND3_X2 U11828 ( .A1(\SB1_2_3/i0_3 ), .A2(\SB1_2_3/i0_4 ), .A3(
        \SB1_2_3/i1[9] ), .ZN(\SB1_2_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U11833 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0_4 ), .A3(
        \SB2_3_17/i1[9] ), .ZN(n2973) );
  NAND3_X1 U11834 ( .A1(\SB1_3_20/i0_0 ), .A2(\SB1_3_20/i1_5 ), .A3(
        \MC_ARK_ARC_1_2/buf_output[70] ), .ZN(
        \SB1_3_20/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U11835 ( .A1(\MC_ARK_ARC_1_3/temp3[120] ), .A2(
        \MC_ARK_ARC_1_3/temp4[120] ), .Z(\MC_ARK_ARC_1_3/temp6[120] ) );
  NAND4_X2 U11839 ( .A1(\SB1_4_3/Component_Function_3/NAND4_in[1] ), .A2(n4933), .A3(n1101), .A4(n1117), .ZN(\SB1_4_3/buf_output[3] ) );
  NAND3_X2 U11841 ( .A1(\SB2_1_10/i0[6] ), .A2(\SB2_1_10/i0_3 ), .A3(
        \SB2_1_10/i0[10] ), .ZN(\SB2_1_10/Component_Function_2/NAND4_in[1] )
         );
  NAND4_X2 U11843 ( .A1(\SB2_2_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_24/Component_Function_0/NAND4_in[1] ), .A3(n1584), .A4(
        \SB2_2_24/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_24/buf_output[0] ) );
  NAND4_X2 U11847 ( .A1(\SB2_0_30/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_30/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_30/Component_Function_4/NAND4_in[1] ), .A4(n4929), .ZN(
        \SB2_0_30/buf_output[4] ) );
  INV_X2 U11848 ( .I(\RI3[0][155] ), .ZN(\SB2_0_6/i1_5 ) );
  INV_X1 U11850 ( .I(\SB1_1_1/buf_output[1] ), .ZN(\SB2_1_29/i1_7 ) );
  NAND4_X2 U11851 ( .A1(\SB1_1_1/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_1_1/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_1/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_1_1/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_1/buf_output[1] ) );
  XOR2_X1 U11853 ( .A1(\MC_ARK_ARC_1_2/temp5[31] ), .A2(
        \MC_ARK_ARC_1_2/temp6[31] ), .Z(\MC_ARK_ARC_1_2/buf_output[31] ) );
  XOR2_X1 U11855 ( .A1(n5323), .A2(\MC_ARK_ARC_1_3/temp4[124] ), .Z(n4930) );
  NAND3_X1 U11856 ( .A1(\SB4_17/i0_4 ), .A2(\SB4_17/i1[9] ), .A3(n3984), .ZN(
        n4931) );
  XOR2_X1 U11857 ( .A1(\RI5[1][31] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[37] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[37] ) );
  NAND3_X2 U11860 ( .A1(\SB1_4_3/i0_3 ), .A2(\SB1_4_3/i0[6] ), .A3(
        \SB1_4_3/i1[9] ), .ZN(n4933) );
  XOR2_X1 U11863 ( .A1(\MC_ARK_ARC_1_2/temp1[1] ), .A2(
        \MC_ARK_ARC_1_2/temp2[1] ), .Z(n1719) );
  NOR2_X2 U11866 ( .A1(n4938), .A2(n4936), .ZN(n1953) );
  NAND2_X1 U11867 ( .A1(\SB1_3_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_4/NAND4_in[3] ), .ZN(n4938) );
  NAND4_X2 U11871 ( .A1(\SB1_3_10/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_3_10/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_3_10/Component_Function_0/NAND4_in[0] ), .A4(n4942), .ZN(
        \SB1_3_10/buf_output[0] ) );
  XOR2_X1 U11874 ( .A1(\MC_ARK_ARC_1_1/temp1[11] ), .A2(
        \MC_ARK_ARC_1_1/temp2[11] ), .Z(n4943) );
  NAND3_X1 U11875 ( .A1(\SB1_2_30/i0_3 ), .A2(\SB1_2_30/i0[9] ), .A3(
        \SB1_2_30/i0[8] ), .ZN(n4944) );
  XOR2_X1 U11878 ( .A1(n4946), .A2(\MC_ARK_ARC_1_3/temp6[94] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[94] ) );
  NAND4_X2 U11880 ( .A1(\SB3_9/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_1/NAND4_in[0] ), .A4(n4947), .ZN(
        \SB3_9/buf_output[1] ) );
  NAND3_X1 U11881 ( .A1(\SB3_9/i0_4 ), .A2(\SB3_9/i1_7 ), .A3(\SB3_9/i0[8] ), 
        .ZN(n4947) );
  XOR2_X1 U11882 ( .A1(n4948), .A2(\MC_ARK_ARC_1_1/temp5[6] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[6] ) );
  XOR2_X1 U11883 ( .A1(\MC_ARK_ARC_1_1/temp4[6] ), .A2(
        \MC_ARK_ARC_1_1/temp3[6] ), .Z(n4948) );
  NAND4_X2 U11887 ( .A1(\SB1_0_26/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_26/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_0_26/Component_Function_2/NAND4_in[1] ), .A4(n4954), .ZN(
        \RI3[0][50] ) );
  NAND3_X1 U11888 ( .A1(\SB1_1_17/i0[10] ), .A2(\SB1_1_17/i1[9] ), .A3(
        \SB1_1_17/i1_7 ), .ZN(\SB1_1_17/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U11889 ( .A1(n4955), .A2(\MC_ARK_ARC_1_0/temp4[97] ), .Z(
        \MC_ARK_ARC_1_0/temp6[97] ) );
  XOR2_X1 U11890 ( .A1(\RI5[0][7] ), .A2(\RI5[0][163] ), .Z(n4955) );
  NAND4_X2 U11891 ( .A1(\SB1_1_9/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_1_9/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_1_9/Component_Function_0/NAND4_in[1] ), .A4(n4956), .ZN(
        \SB1_1_9/buf_output[0] ) );
  NAND3_X1 U11894 ( .A1(\SB1_4_4/i0[10] ), .A2(\SB1_4_4/i1[9] ), .A3(
        \SB1_4_4/i1_7 ), .ZN(n4962) );
  XOR2_X1 U11896 ( .A1(\MC_ARK_ARC_1_0/temp2[79] ), .A2(
        \MC_ARK_ARC_1_0/temp1[79] ), .Z(n4963) );
  NAND3_X1 U11897 ( .A1(\RI3[0][28] ), .A2(\SB2_0_27/i0[8] ), .A3(
        \SB2_0_27/i1_7 ), .ZN(n4964) );
  XOR2_X1 U11899 ( .A1(\RI5[3][139] ), .A2(\RI5[3][175] ), .Z(
        \MC_ARK_ARC_1_3/temp3[73] ) );
  NAND3_X1 U11901 ( .A1(\SB1_3_16/i0_4 ), .A2(\SB1_3_16/i0_0 ), .A3(
        \SB1_3_16/i0_3 ), .ZN(\SB1_3_16/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U11903 ( .A1(n4970), .A2(n4969), .Z(n1853) );
  XOR2_X1 U11904 ( .A1(\RI5[1][143] ), .A2(n464), .Z(n4969) );
  XOR2_X1 U11905 ( .A1(\RI5[1][77] ), .A2(\RI5[1][107] ), .Z(n4970) );
  XOR2_X1 U11908 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[140] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[176] ), .Z(n4972) );
  XOR2_X1 U11909 ( .A1(n4975), .A2(n4974), .Z(\MC_ARK_ARC_1_3/temp5[131] ) );
  XOR2_X1 U11910 ( .A1(\RI5[3][101] ), .A2(\RI5[3][125] ), .Z(n4974) );
  XOR2_X1 U11911 ( .A1(\RI5[3][131] ), .A2(\RI5[3][77] ), .Z(n4975) );
  XOR2_X1 U11914 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[165] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[9] ), .Z(n4978) );
  XOR2_X1 U11918 ( .A1(n2479), .A2(n4981), .Z(\MC_ARK_ARC_1_0/buf_output[75] )
         );
  XOR2_X1 U11919 ( .A1(n4982), .A2(\MC_ARK_ARC_1_0/temp6[78] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[78] ) );
  XOR2_X1 U11920 ( .A1(\MC_ARK_ARC_1_0/temp2[78] ), .A2(
        \MC_ARK_ARC_1_0/temp1[78] ), .Z(n4982) );
  NAND3_X2 U11922 ( .A1(\SB1_4_31/i0_3 ), .A2(\SB1_4_31/i1[9] ), .A3(
        \SB1_4_31/i0_4 ), .ZN(\SB1_4_31/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U11923 ( .A1(\SB1_1_21/i0_4 ), .A2(\SB1_1_21/i1_5 ), .A3(
        \SB1_1_21/i1[9] ), .ZN(n4984) );
  NAND3_X1 U11924 ( .A1(\SB1_0_5/i0_4 ), .A2(\SB1_0_5/i1[9] ), .A3(
        \SB1_0_5/i1_5 ), .ZN(\SB1_0_5/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U11926 ( .A1(\SB2_4_3/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_3/Component_Function_0/NAND4_in[0] ), .A4(n4985), .ZN(
        \SB2_4_3/buf_output[0] ) );
  XOR2_X1 U11929 ( .A1(\MC_ARK_ARC_1_0/temp4[117] ), .A2(n4987), .Z(n5268) );
  XOR2_X1 U11930 ( .A1(\RI5[0][183] ), .A2(\RI5[0][27] ), .Z(n4987) );
  XOR2_X1 U11931 ( .A1(\RI5[1][183] ), .A2(\RI5[1][27] ), .Z(
        \MC_ARK_ARC_1_1/temp3[117] ) );
  NAND3_X1 U11932 ( .A1(n2381), .A2(\SB2_0_5/i0[8] ), .A3(\SB2_0_5/i0[6] ), 
        .ZN(\SB2_0_5/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U11933 ( .A1(\MC_ARK_ARC_1_2/temp3[1] ), .A2(
        \MC_ARK_ARC_1_2/temp4[1] ), .Z(n4988) );
  NAND3_X2 U11934 ( .A1(n571), .A2(\SB2_3_16/i3[0] ), .A3(\SB2_3_16/i0[8] ), 
        .ZN(\SB2_3_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U11935 ( .A1(\SB4_26/i0_3 ), .A2(\SB4_26/i0[6] ), .A3(n573), .ZN(
        n4990) );
  NAND4_X2 U11937 ( .A1(\SB3_3/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_3/Component_Function_4/NAND4_in[0] ), .A4(n4992), .ZN(
        \SB3_3/buf_output[4] ) );
  NAND3_X1 U11938 ( .A1(\SB3_3/i0_4 ), .A2(\SB3_3/i1[9] ), .A3(\SB3_3/i1_5 ), 
        .ZN(n4992) );
  INV_X2 U11942 ( .I(\SB1_1_25/buf_output[2] ), .ZN(\SB2_1_22/i1[9] ) );
  NAND3_X2 U11945 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i0_4 ), .A3(
        \SB2_1_5/i1[9] ), .ZN(\SB2_1_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U11946 ( .A1(\SB4_25/i0_4 ), .A2(\SB4_25/i0_3 ), .A3(\SB4_25/i0_0 ), 
        .ZN(\SB4_25/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U11948 ( .A1(\MC_ARK_ARC_1_1/temp4[186] ), .A2(
        \MC_ARK_ARC_1_1/temp3[186] ), .Z(\MC_ARK_ARC_1_1/temp6[186] ) );
  NAND3_X1 U11949 ( .A1(\SB4_14/i0[6] ), .A2(\SB4_14/i0[8] ), .A3(
        \SB4_14/i0[7] ), .ZN(n4997) );
  XOR2_X1 U11951 ( .A1(\RI5[2][51] ), .A2(\RI5[2][75] ), .Z(n4998) );
  XOR2_X1 U11953 ( .A1(n5000), .A2(\MC_ARK_ARC_1_3/temp6[130] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[130] ) );
  XOR2_X1 U11954 ( .A1(\MC_ARK_ARC_1_3/temp2[130] ), .A2(
        \MC_ARK_ARC_1_3/temp1[130] ), .Z(n5000) );
  XOR2_X1 U11955 ( .A1(\RI5[0][190] ), .A2(\RI5[0][154] ), .Z(
        \MC_ARK_ARC_1_0/temp3[88] ) );
  NAND3_X2 U11957 ( .A1(\SB1_3_14/i0[6] ), .A2(\SB1_3_14/i1[9] ), .A3(
        \RI1[3][107] ), .ZN(n5005) );
  NOR2_X1 U11958 ( .A1(\SB2_4_15/i0[8] ), .A2(\SB2_4_15/i1_7 ), .ZN(n2152) );
  XOR2_X1 U11961 ( .A1(n5003), .A2(n57), .Z(Ciphertext[7]) );
  NAND4_X2 U11962 ( .A1(\SB4_30/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_30/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_30/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_30/Component_Function_1/NAND4_in[0] ), .ZN(n5003) );
  NAND3_X1 U11963 ( .A1(n3308), .A2(\SB2_3_28/i0_3 ), .A3(\SB2_3_28/i0_0 ), 
        .ZN(\SB2_3_28/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U11964 ( .A1(\SB1_3_14/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_3_14/Component_Function_3/NAND4_in[1] ), .A3(n913), .A4(n5005), 
        .ZN(\SB1_3_14/buf_output[3] ) );
  NAND3_X2 U11966 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0_0 ), .A3(n594), 
        .ZN(n5007) );
  NAND4_X2 U11968 ( .A1(n5047), .A2(\SB2_1_1/Component_Function_4/NAND4_in[2] ), .A3(\SB2_1_1/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_1_1/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB2_1_1/buf_output[4] ) );
  NAND3_X1 U11970 ( .A1(\SB1_1_1/i0_0 ), .A2(\SB1_1_1/i3[0] ), .A3(
        \SB1_1_1/i1_7 ), .ZN(\SB1_1_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U11972 ( .A1(\SB1_0_13/i0[6] ), .A2(\SB1_0_13/i1_5 ), .A3(
        \SB1_0_13/i0[9] ), .ZN(\SB1_0_13/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U11974 ( .A1(\SB2_3_14/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_14/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_14/Component_Function_0/NAND4_in[0] ), .A4(n5009), .ZN(
        \SB2_3_14/buf_output[0] ) );
  XOR2_X1 U11975 ( .A1(n5010), .A2(n100), .Z(Ciphertext[163]) );
  NAND3_X1 U11978 ( .A1(\SB2_3_5/i1[9] ), .A2(\SB2_3_5/i0_4 ), .A3(
        \SB2_3_5/i1_5 ), .ZN(n5011) );
  NAND4_X2 U11979 ( .A1(\SB2_4_16/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_4_16/Component_Function_2/NAND4_in[0] ), .A3(n1027), .A4(n5012), 
        .ZN(\SB2_4_16/buf_output[2] ) );
  NAND4_X2 U11980 ( .A1(\SB1_4_19/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_4_19/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_4_19/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_4_19/Component_Function_1/NAND4_in[1] ), .ZN(
        \SB1_4_19/buf_output[1] ) );
  NAND3_X1 U11982 ( .A1(\SB4_9/i0[6] ), .A2(\SB4_9/i1_5 ), .A3(\SB4_9/i0[9] ), 
        .ZN(\SB4_9/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U11985 ( .A1(\MC_ARK_ARC_1_4/temp1[141] ), .A2(
        \MC_ARK_ARC_1_4/temp2[141] ), .Z(\MC_ARK_ARC_1_4/temp5[141] ) );
  NAND4_X2 U11986 ( .A1(\SB1_4_13/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_4_13/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_4_13/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_4_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_4_13/buf_output[0] ) );
  XOR2_X1 U11987 ( .A1(\MC_ARK_ARC_1_4/temp1[183] ), .A2(n5016), .Z(n1394) );
  XOR2_X1 U11988 ( .A1(\RI5[4][153] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[129] ), .Z(n5016) );
  XOR2_X1 U11989 ( .A1(n5017), .A2(\MC_ARK_ARC_1_3/temp6[138] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[138] ) );
  NAND4_X2 U11991 ( .A1(\SB2_0_10/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_0_10/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_10/Component_Function_4/NAND4_in[2] ), .A4(n5018), .ZN(
        \SB2_0_10/buf_output[4] ) );
  XOR2_X1 U11994 ( .A1(\MC_ARK_ARC_1_3/temp2[172] ), .A2(n5019), .Z(
        \MC_ARK_ARC_1_3/temp5[172] ) );
  XOR2_X1 U11995 ( .A1(\RI5[3][172] ), .A2(\RI5[3][166] ), .Z(n5019) );
  XOR2_X1 U11996 ( .A1(\MC_ARK_ARC_1_3/temp1[187] ), .A2(n5020), .Z(
        \MC_ARK_ARC_1_3/temp5[187] ) );
  XOR2_X1 U11997 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[133] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[157] ), .Z(n5020) );
  NAND3_X1 U11998 ( .A1(\SB2_3_13/i0[6] ), .A2(\SB2_3_13/i1_5 ), .A3(
        \SB2_3_13/i0[9] ), .ZN(\SB2_3_13/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U11999 ( .A1(\MC_ARK_ARC_1_2/temp1[86] ), .A2(n5021), .Z(
        \MC_ARK_ARC_1_2/temp5[86] ) );
  XOR2_X1 U12000 ( .A1(\RI5[2][32] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .Z(n5021) );
  NOR2_X2 U12001 ( .A1(n2347), .A2(n5022), .ZN(n2554) );
  NAND2_X2 U12002 ( .A1(n2960), .A2(n2346), .ZN(n5022) );
  XOR2_X1 U12007 ( .A1(n5027), .A2(\MC_ARK_ARC_1_4/temp6[42] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[42] ) );
  XOR2_X1 U12008 ( .A1(\MC_ARK_ARC_1_4/temp1[42] ), .A2(
        \MC_ARK_ARC_1_4/temp2[42] ), .Z(n5027) );
  XOR2_X1 U12009 ( .A1(n5028), .A2(n92), .Z(Ciphertext[137]) );
  NAND4_X2 U12010 ( .A1(\SB4_9/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_9/Component_Function_5/NAND4_in[3] ), .A3(n5249), .A4(
        \SB4_9/Component_Function_5/NAND4_in[0] ), .ZN(n5028) );
  NAND4_X2 U12011 ( .A1(n5223), .A2(\SB2_2_7/Component_Function_3/NAND4_in[0] ), .A3(\SB2_2_7/Component_Function_3/NAND4_in[3] ), .A4(n5029), .ZN(
        \SB2_2_7/buf_output[3] ) );
  NAND3_X2 U12012 ( .A1(\SB2_2_7/i0_0 ), .A2(\SB2_2_7/i0_3 ), .A3(
        \SB2_2_7/i0_4 ), .ZN(n5029) );
  NAND4_X2 U12015 ( .A1(\SB2_2_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_27/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_27/Component_Function_1/NAND4_in[0] ), .A4(n5031), .ZN(
        \SB2_2_27/buf_output[1] ) );
  XOR2_X1 U12017 ( .A1(\RI5[1][176] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[152] ), .Z(n5033) );
  NAND3_X1 U12019 ( .A1(\SB4_14/i0_3 ), .A2(\SB4_14/i0[9] ), .A3(
        \SB4_14/i0[10] ), .ZN(\SB4_14/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U12020 ( .A1(\MC_ARK_ARC_1_3/temp5[0] ), .A2(n5038), .Z(
        \MC_ARK_ARC_1_3/buf_output[0] ) );
  XOR2_X1 U12021 ( .A1(\MC_ARK_ARC_1_3/temp3[0] ), .A2(
        \MC_ARK_ARC_1_3/temp4[0] ), .Z(n5038) );
  XOR2_X1 U12022 ( .A1(n5039), .A2(\MC_ARK_ARC_1_4/temp6[11] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[11] ) );
  NAND3_X1 U12023 ( .A1(\SB1_4_2/i0[8] ), .A2(\SB1_4_2/i1_7 ), .A3(
        \SB1_4_2/i0_4 ), .ZN(n5040) );
  NAND4_X2 U12028 ( .A1(\SB2_2_3/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_3/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_3/Component_Function_3/NAND4_in[3] ), .A4(n5042), .ZN(
        \SB2_2_3/buf_output[3] ) );
  NAND3_X2 U12029 ( .A1(\SB2_2_3/i0[10] ), .A2(\SB2_2_3/i1[9] ), .A3(
        \SB2_2_3/i1_7 ), .ZN(n5042) );
  XOR2_X1 U12030 ( .A1(\MC_ARK_ARC_1_0/temp5[97] ), .A2(
        \MC_ARK_ARC_1_0/temp6[97] ), .Z(\MC_ARK_ARC_1_0/buf_output[97] ) );
  NAND3_X2 U12032 ( .A1(\SB2_0_11/i0[10] ), .A2(\SB2_0_11/i0_0 ), .A3(
        \SB2_0_11/i0[6] ), .ZN(n5049) );
  NAND3_X1 U12033 ( .A1(\SB2_1_1/i0_4 ), .A2(\SB2_1_1/i1[9] ), .A3(
        \SB2_1_1/i1_5 ), .ZN(n5047) );
  INV_X2 U12034 ( .I(\SB1_4_14/buf_output[3] ), .ZN(\SB2_4_12/i0[8] ) );
  NAND3_X1 U12035 ( .A1(\SB3_3/i1_7 ), .A2(\SB3_3/i3[0] ), .A3(\SB3_3/i0_0 ), 
        .ZN(\SB3_3/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U12036 ( .A1(\MC_ARK_ARC_1_1/temp5[190] ), .A2(n3133), .Z(
        \MC_ARK_ARC_1_1/buf_output[190] ) );
  NAND3_X2 U12039 ( .A1(n851), .A2(\SB2_3_10/i0[9] ), .A3(\SB2_3_10/i0[6] ), 
        .ZN(n2792) );
  XOR2_X1 U12042 ( .A1(\RI5[1][127] ), .A2(\RI5[1][133] ), .Z(
        \MC_ARK_ARC_1_1/temp1[133] ) );
  NAND4_X2 U12043 ( .A1(\SB2_4_0/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_4_0/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_4_0/Component_Function_4/NAND4_in[1] ), .A4(n5051), .ZN(
        \SB2_4_0/buf_output[4] ) );
  NAND4_X2 U12044 ( .A1(\SB2_0_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_11/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_11/Component_Function_2/NAND4_in[3] ), .A4(n5052), .ZN(
        \SB2_0_11/buf_output[2] ) );
  NAND3_X2 U12045 ( .A1(\SB1_3_25/i0_3 ), .A2(\SB1_3_25/i1[9] ), .A3(
        \SB1_3_25/i0[6] ), .ZN(\SB1_3_25/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12051 ( .A1(\RI5[0][152] ), .A2(\RI5[0][122] ), .Z(n5055) );
  XOR2_X1 U12052 ( .A1(\RI5[0][98] ), .A2(\RI5[0][146] ), .Z(n5056) );
  NAND3_X2 U12053 ( .A1(\SB1_0_13/i0[10] ), .A2(\SB1_0_13/i1[9] ), .A3(
        \SB1_0_13/i1_5 ), .ZN(\SB1_0_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U12056 ( .A1(\SB2_3_7/i0[6] ), .A2(\SB2_3_7/i0[9] ), .A3(
        \SB2_3_7/i1_5 ), .ZN(n5088) );
  NAND4_X2 U12058 ( .A1(\SB1_0_11/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_11/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_11/Component_Function_3/NAND4_in[3] ), .A4(n5059), .ZN(
        \SB1_0_11/buf_output[3] ) );
  XOR2_X1 U12060 ( .A1(\RI5[1][33] ), .A2(\RI5[1][27] ), .Z(n5060) );
  XOR2_X1 U12061 ( .A1(\RI5[0][128] ), .A2(\RI5[0][152] ), .Z(
        \MC_ARK_ARC_1_0/temp2[182] ) );
  NAND3_X1 U12062 ( .A1(n851), .A2(\SB2_3_10/i0_3 ), .A3(\SB2_3_10/i0[10] ), 
        .ZN(\SB2_3_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U12063 ( .A1(\SB3_13/i0_3 ), .A2(\SB3_13/i0[7] ), .A3(\SB3_13/i0_0 ), .ZN(n1806) );
  XOR2_X1 U12065 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[151] ), .A2(\RI5[3][127] ), .Z(n5062) );
  INV_X1 U12066 ( .I(\SB3_2/buf_output[5] ), .ZN(\SB4_2/i1_5 ) );
  INV_X2 U12069 ( .I(\SB1_4_3/buf_output[3] ), .ZN(\SB2_4_1/i0[8] ) );
  XOR2_X1 U12071 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[164] ), .A2(\RI5[3][8] ), 
        .Z(n5067) );
  XOR2_X1 U12073 ( .A1(n5069), .A2(\MC_ARK_ARC_1_2/temp2[129] ), .Z(
        \MC_ARK_ARC_1_2/temp5[129] ) );
  XOR2_X1 U12074 ( .A1(\RI5[2][123] ), .A2(\RI5[2][129] ), .Z(n5069) );
  NAND4_X2 U12076 ( .A1(\SB2_2_9/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_9/Component_Function_0/NAND4_in[0] ), .A4(n5072), .ZN(
        \SB2_2_9/buf_output[0] ) );
  XOR2_X1 U12077 ( .A1(\MC_ARK_ARC_1_3/temp2[47] ), .A2(n2462), .Z(n3060) );
  NAND3_X1 U12079 ( .A1(\SB4_0/i0[10] ), .A2(\SB4_0/i1_5 ), .A3(\SB4_0/i1[9] ), 
        .ZN(\SB4_0/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U12080 ( .A1(\MC_ARK_ARC_1_3/temp6[103] ), .A2(n5073), .Z(
        \MC_ARK_ARC_1_3/buf_output[103] ) );
  XOR2_X1 U12083 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[117] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[141] ), .Z(n5074) );
  XOR2_X1 U12084 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[151] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[157] ), .Z(\MC_ARK_ARC_1_3/temp1[157] )
         );
  XOR2_X1 U12086 ( .A1(n5076), .A2(n804), .Z(\MC_ARK_ARC_1_3/temp5[23] ) );
  XOR2_X1 U12087 ( .A1(\RI5[3][23] ), .A2(\RI5[3][161] ), .Z(n5076) );
  NAND3_X2 U12088 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i1[9] ), .A3(
        \SB1_1_14/i0[6] ), .ZN(\SB1_1_14/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12090 ( .A1(\MC_ARK_ARC_1_3/temp2[91] ), .A2(
        \MC_ARK_ARC_1_3/temp3[91] ), .Z(n5077) );
  NAND3_X2 U12091 ( .A1(\SB1_4_6/i0[10] ), .A2(\RI1[4][155] ), .A3(
        \SB1_4_6/i0[6] ), .ZN(n5079) );
  NAND4_X2 U12092 ( .A1(\SB1_4_15/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_4_15/Component_Function_5/NAND4_in[0] ), .A3(n5299), .A4(n5080), 
        .ZN(\SB1_4_15/buf_output[5] ) );
  NAND3_X2 U12093 ( .A1(\SB1_4_15/i0_4 ), .A2(\SB1_4_15/i0[6] ), .A3(
        \SB1_4_15/i0[9] ), .ZN(n5080) );
  NAND3_X1 U12094 ( .A1(\SB2_0_9/i0_4 ), .A2(\SB2_0_9/i1[9] ), .A3(
        \SB2_0_9/i1_5 ), .ZN(\SB2_0_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U12095 ( .A1(\SB2_2_14/i0_0 ), .A2(\SB2_2_14/i0_4 ), .A3(
        \SB2_2_14/i1_5 ), .ZN(n5151) );
  NAND4_X2 U12096 ( .A1(n5335), .A2(\SB3_26/Component_Function_0/NAND4_in[1] ), 
        .A3(\SB3_26/Component_Function_0/NAND4_in[0] ), .A4(n5081), .ZN(
        \SB3_26/buf_output[0] ) );
  NAND3_X1 U12098 ( .A1(\SB1_2_15/i0_0 ), .A2(\SB1_2_15/i0[9] ), .A3(
        \SB1_2_15/i0[8] ), .ZN(\SB1_2_15/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U12099 ( .A1(n5085), .A2(n5084), .Z(\MC_ARK_ARC_1_2/temp6[65] ) );
  XOR2_X1 U12100 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[131] ), .A2(n476), .Z(
        n5084) );
  XOR2_X1 U12104 ( .A1(n1999), .A2(n5108), .Z(n5087) );
  XOR2_X1 U12106 ( .A1(\RI5[2][6] ), .A2(\RI5[2][42] ), .Z(
        \MC_ARK_ARC_1_2/temp3[132] ) );
  XOR2_X1 U12108 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[162] ), .A2(\RI5[2][156] ), .Z(n5089) );
  NAND3_X1 U12110 ( .A1(\SB2_2_4/i0_4 ), .A2(\SB2_2_4/i0[8] ), .A3(
        \SB2_2_4/i1_7 ), .ZN(\SB2_2_4/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U12111 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[109] ), .A2(\RI5[3][73] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[7] ) );
  XOR2_X1 U12112 ( .A1(\RI5[2][157] ), .A2(n468), .Z(
        \MC_ARK_ARC_1_2/temp4[121] ) );
  NAND3_X1 U12118 ( .A1(\SB1_3_12/i0[10] ), .A2(\SB1_3_12/i0_3 ), .A3(
        \SB1_3_12/i0[9] ), .ZN(n5092) );
  XOR2_X1 U12119 ( .A1(n5093), .A2(\MC_ARK_ARC_1_0/temp6[32] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[32] ) );
  XOR2_X1 U12120 ( .A1(\MC_ARK_ARC_1_0/temp1[32] ), .A2(
        \MC_ARK_ARC_1_0/temp2[32] ), .Z(n5093) );
  XOR2_X1 U12121 ( .A1(n5096), .A2(n5095), .Z(\MC_ARK_ARC_1_0/temp6[155] ) );
  XOR2_X1 U12122 ( .A1(\RI5[0][29] ), .A2(n134), .Z(n5095) );
  NAND3_X2 U12126 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i1_7 ), .A3(
        \SB2_2_0/i0[8] ), .ZN(n1630) );
  XOR2_X1 U12127 ( .A1(\RI5[1][98] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .Z(n5097) );
  NAND3_X2 U12128 ( .A1(\SB2_1_24/i0_0 ), .A2(\SB2_1_24/i0_4 ), .A3(
        \SB2_1_24/i1_5 ), .ZN(n1844) );
  XOR2_X1 U12129 ( .A1(\MC_ARK_ARC_1_2/temp1[178] ), .A2(n5098), .Z(n5113) );
  XOR2_X1 U12130 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[52] ), .A2(\RI5[2][88] ), 
        .Z(n5098) );
  NAND3_X2 U12132 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0[10] ), .A3(
        \SB2_2_24/i0[9] ), .ZN(n5365) );
  NAND4_X2 U12136 ( .A1(\SB3_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_19/Component_Function_0/NAND4_in[0] ), .A4(n5103), .ZN(
        \SB3_19/buf_output[0] ) );
  NAND3_X2 U12141 ( .A1(\SB1_0_11/i0[10] ), .A2(\SB1_0_11/i0_0 ), .A3(
        \SB1_0_11/i0[6] ), .ZN(n5186) );
  XOR2_X1 U12143 ( .A1(\RI5[3][107] ), .A2(\RI5[3][137] ), .Z(n5108) );
  XOR2_X1 U12144 ( .A1(n5395), .A2(\MC_ARK_ARC_1_2/temp6[92] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[92] ) );
  NAND3_X1 U12146 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i0_3 ), .A3(\SB4_8/i0[7] ), 
        .ZN(n5110) );
  XOR2_X1 U12147 ( .A1(\RI5[2][76] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[112] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[10] ) );
  NAND3_X2 U12148 ( .A1(\SB2_4_20/i0_3 ), .A2(\SB2_4_20/i0_4 ), .A3(
        \SB2_4_20/i1[9] ), .ZN(n3135) );
  XOR2_X1 U12152 ( .A1(\MC_ARK_ARC_1_3/temp3[70] ), .A2(
        \MC_ARK_ARC_1_3/temp4[70] ), .Z(\MC_ARK_ARC_1_3/temp6[70] ) );
  XOR2_X1 U12153 ( .A1(n5113), .A2(n5112), .Z(\MC_ARK_ARC_1_2/buf_output[178] ) );
  XOR2_X1 U12154 ( .A1(\MC_ARK_ARC_1_2/temp2[178] ), .A2(
        \MC_ARK_ARC_1_2/temp4[178] ), .Z(n5112) );
  NAND3_X1 U12155 ( .A1(\SB1_3_2/i0_4 ), .A2(\SB1_3_2/i1[9] ), .A3(
        \SB1_3_2/i1_5 ), .ZN(\SB1_3_2/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U12156 ( .A1(n5115), .A2(\MC_ARK_ARC_1_3/temp1[35] ), .Z(
        \MC_ARK_ARC_1_3/temp5[35] ) );
  XOR2_X1 U12157 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[5] ), .A2(\RI5[3][173] ), 
        .Z(n5115) );
  NAND3_X2 U12160 ( .A1(\SB1_3_7/i0_0 ), .A2(\SB1_3_7/i1_5 ), .A3(
        \SB1_3_7/i0_4 ), .ZN(n1247) );
  NAND3_X2 U12161 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i1[9] ), .A3(
        \SB3_23/i0[6] ), .ZN(n5118) );
  NAND3_X2 U12163 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0_4 ), .A3(
        \SB2_2_28/i0_0 ), .ZN(n5120) );
  XOR2_X1 U12165 ( .A1(\RI5[0][185] ), .A2(\RI5[0][17] ), .Z(
        \MC_ARK_ARC_1_0/temp2[47] ) );
  XOR2_X1 U12166 ( .A1(n5123), .A2(\MC_ARK_ARC_1_2/temp5[12] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[12] ) );
  NAND4_X2 U12167 ( .A1(\SB2_3_26/Component_Function_5/NAND4_in[2] ), .A2(
        n2006), .A3(\SB2_3_26/Component_Function_5/NAND4_in[3] ), .A4(n5124), 
        .ZN(\SB2_3_26/buf_output[5] ) );
  NAND2_X2 U12168 ( .A1(\SB2_3_26/i0_0 ), .A2(\SB2_3_26/i3[0] ), .ZN(n5124) );
  NAND4_X2 U12171 ( .A1(n1970), .A2(
        \SB2_2_28/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_2_28/Component_Function_0/NAND4_in[1] ), .A4(n5126), .ZN(
        \SB2_2_28/buf_output[0] ) );
  NAND3_X2 U12172 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0[10] ), .A3(
        \SB2_2_28/i0_4 ), .ZN(n5126) );
  NAND4_X2 U12174 ( .A1(\SB1_2_18/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_18/Component_Function_0/NAND4_in[2] ), .A3(n5129), .A4(
        \SB1_2_18/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_18/buf_output[0] ) );
  XOR2_X1 U12177 ( .A1(\RI5[3][113] ), .A2(\RI5[3][149] ), .Z(
        \MC_ARK_ARC_1_3/temp3[47] ) );
  XOR2_X1 U12179 ( .A1(n5131), .A2(n157), .Z(Ciphertext[80]) );
  INV_X2 U12180 ( .I(\SB1_0_7/buf_output[2] ), .ZN(\SB2_0_4/i1[9] ) );
  NAND4_X2 U12181 ( .A1(\SB1_0_7/Component_Function_2/NAND4_in[0] ), .A2(n5338), .A3(\SB1_0_7/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_7/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB1_0_7/buf_output[2] ) );
  XOR2_X1 U12183 ( .A1(\MC_ARK_ARC_1_4/temp3[64] ), .A2(
        \MC_ARK_ARC_1_4/temp4[64] ), .Z(\MC_ARK_ARC_1_4/temp6[64] ) );
  NAND3_X1 U12184 ( .A1(\SB4_4/i0_3 ), .A2(\SB4_4/i0[9] ), .A3(\SB4_4/i0[8] ), 
        .ZN(\SB4_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U12186 ( .A1(\SB1_1_8/i0[10] ), .A2(\SB1_1_8/i1[9] ), .A3(
        \SB1_1_8/i1_7 ), .ZN(n5133) );
  XOR2_X1 U12187 ( .A1(\MC_ARK_ARC_1_0/temp6[21] ), .A2(n5134), .Z(
        \MC_ARK_ARC_1_0/buf_output[21] ) );
  INV_X2 U12189 ( .I(\SB1_3_0/buf_output[5] ), .ZN(\SB2_3_0/i1_5 ) );
  NAND3_X2 U12192 ( .A1(\SB2_1_10/i0[6] ), .A2(\SB2_1_10/i0_0 ), .A3(
        \SB2_1_10/i0[10] ), .ZN(\SB2_1_10/Component_Function_5/NAND4_in[1] )
         );
  XOR2_X1 U12195 ( .A1(n578), .A2(\RI5[1][16] ), .Z(
        \MC_ARK_ARC_1_1/temp3[106] ) );
  NAND3_X2 U12196 ( .A1(\SB1_1_14/i0[10] ), .A2(\SB1_1_14/i1[9] ), .A3(
        \SB1_1_14/i1_5 ), .ZN(\SB1_1_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U12197 ( .A1(\SB2_4_14/i0[10] ), .A2(\SB2_4_14/i0_3 ), .A3(
        \SB2_4_14/i0_4 ), .ZN(\SB2_4_14/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U12198 ( .A1(\RI5[2][11] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .Z(n5261) );
  XOR2_X1 U12199 ( .A1(\RI5[2][129] ), .A2(\RI5[2][135] ), .Z(
        \MC_ARK_ARC_1_2/temp1[135] ) );
  NAND4_X2 U12200 ( .A1(\SB2_4_29/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_4_29/Component_Function_2/NAND4_in[0] ), .A3(n1337), .A4(
        \SB2_4_29/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_4_29/buf_output[2] ) );
  XOR2_X1 U12202 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[117] ), .A2(\RI5[1][111] ), .Z(\MC_ARK_ARC_1_1/temp1[117] ) );
  XOR2_X1 U12205 ( .A1(\RI5[2][135] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[171] ), .Z(\MC_ARK_ARC_1_2/temp3[69] ) );
  XOR2_X1 U12208 ( .A1(\MC_ARK_ARC_1_4/temp5[83] ), .A2(
        \MC_ARK_ARC_1_4/temp6[83] ), .Z(\MC_ARK_ARC_1_4/buf_output[83] ) );
  NAND4_X2 U12213 ( .A1(\SB1_2_16/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_16/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_16/Component_Function_4/NAND4_in[3] ), .A4(n5142), .ZN(
        \SB1_2_16/buf_output[4] ) );
  XOR2_X1 U12215 ( .A1(n5143), .A2(\MC_ARK_ARC_1_2/temp2[10] ), .Z(
        \MC_ARK_ARC_1_2/temp5[10] ) );
  XOR2_X1 U12216 ( .A1(\RI5[2][4] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[10] ), 
        .Z(n5143) );
  XOR2_X1 U12217 ( .A1(\RI5[2][77] ), .A2(\RI5[2][113] ), .Z(
        \MC_ARK_ARC_1_2/temp3[11] ) );
  NAND4_X2 U12218 ( .A1(\SB2_1_6/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_0/NAND4_in[0] ), .A4(n5144), .ZN(
        \SB2_1_6/buf_output[0] ) );
  NAND4_X2 U12220 ( .A1(\SB2_3_18/Component_Function_2/NAND4_in[0] ), .A2(
        n2515), .A3(n1972), .A4(n5145), .ZN(\SB2_3_18/buf_output[2] ) );
  NAND3_X2 U12221 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0[10] ), .A3(
        \SB2_3_18/i0[6] ), .ZN(n5145) );
  NAND2_X2 U12222 ( .A1(\SB2_2_22/i0_0 ), .A2(\SB2_2_22/i3[0] ), .ZN(n5147) );
  NAND3_X1 U12224 ( .A1(\SB1_4_24/i0_4 ), .A2(\SB1_4_24/i1[9] ), .A3(
        \SB1_4_24/i1_5 ), .ZN(n5149) );
  XOR2_X1 U12227 ( .A1(\RI5[0][14] ), .A2(\RI5[0][170] ), .Z(
        \MC_ARK_ARC_1_0/temp3[104] ) );
  INV_X2 U12229 ( .I(\SB1_1_29/buf_output[5] ), .ZN(\SB2_1_29/i1_5 ) );
  XOR2_X1 U12230 ( .A1(\RI5[2][113] ), .A2(\RI5[2][107] ), .Z(n5153) );
  NAND3_X1 U12232 ( .A1(\SB1_4_31/i0_0 ), .A2(\SB1_4_31/i1_5 ), .A3(
        \SB1_4_31/i0_4 ), .ZN(n5155) );
  XOR2_X1 U12242 ( .A1(\RI5[4][81] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[87] ), 
        .Z(n5162) );
  XOR2_X1 U12243 ( .A1(n5165), .A2(n5164), .Z(\MC_ARK_ARC_1_1/buf_output[116] ) );
  XOR2_X1 U12244 ( .A1(n2951), .A2(n1062), .Z(n5164) );
  XOR2_X1 U12246 ( .A1(\RI5[4][26] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[2] ), 
        .Z(n5169) );
  XOR2_X1 U12248 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[120] ), .A2(\RI5[2][126] ), .Z(\MC_ARK_ARC_1_2/temp1[126] ) );
  NAND4_X2 U12249 ( .A1(\SB2_2_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_11/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_11/Component_Function_4/NAND4_in[1] ), .A4(n5170), .ZN(
        \SB2_2_11/buf_output[4] ) );
  XOR2_X1 U12251 ( .A1(\MC_ARK_ARC_1_2/temp3[35] ), .A2(
        \MC_ARK_ARC_1_2/temp4[35] ), .Z(n5171) );
  NAND3_X1 U12252 ( .A1(\SB1_4_31/buf_output[4] ), .A2(\SB2_4_30/i0[8] ), .A3(
        \SB2_4_30/i1_7 ), .ZN(n5172) );
  NAND3_X1 U12255 ( .A1(\SB4_4/i0_4 ), .A2(\SB4_4/i0[9] ), .A3(\SB4_4/i0[6] ), 
        .ZN(n5173) );
  NAND4_X2 U12256 ( .A1(\SB1_3_1/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_1/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_3_1/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_1/buf_output[1] ) );
  NAND4_X2 U12259 ( .A1(\SB1_4_17/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_4_17/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_4_17/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_4_17/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_4_17/buf_output[0] ) );
  NAND4_X2 U12263 ( .A1(\SB1_3_30/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_30/Component_Function_1/NAND4_in[0] ), .A4(n5176), .ZN(
        \SB1_3_30/buf_output[1] ) );
  NAND3_X1 U12264 ( .A1(\SB1_3_30/i0_4 ), .A2(\SB1_3_30/i1_7 ), .A3(
        \SB1_3_30/i0[8] ), .ZN(n5176) );
  NAND3_X2 U12265 ( .A1(\SB2_1_11/i0_3 ), .A2(\SB2_1_11/i0_4 ), .A3(
        \SB2_1_11/i1[9] ), .ZN(\SB2_1_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U12267 ( .A1(\SB2_1_17/i0_0 ), .A2(\SB2_1_17/i0[10] ), .A3(
        \SB2_1_17/i0[6] ), .ZN(n5178) );
  NAND3_X1 U12268 ( .A1(\SB2_4_9/i0_3 ), .A2(\SB1_4_14/buf_output[0] ), .A3(
        \SB2_4_9/i0[8] ), .ZN(\SB2_4_9/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U12271 ( .A1(n5181), .A2(n2361), .Z(\MC_ARK_ARC_1_1/buf_output[75] )
         );
  XOR2_X1 U12272 ( .A1(\MC_ARK_ARC_1_1/temp4[75] ), .A2(
        \MC_ARK_ARC_1_1/temp3[75] ), .Z(n5181) );
  XOR2_X1 U12274 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[143] ), .A2(\RI5[2][107] ), .Z(n5183) );
  XOR2_X1 U12277 ( .A1(\MC_ARK_ARC_1_2/temp3[186] ), .A2(
        \MC_ARK_ARC_1_2/temp4[186] ), .Z(n5185) );
  NAND4_X2 U12278 ( .A1(\SB1_0_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_11/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_0_11/Component_Function_5/NAND4_in[0] ), .A4(n5186), .ZN(
        \RI3[0][125] ) );
  XOR2_X1 U12280 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[147] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[171] ), .Z(\MC_ARK_ARC_1_2/temp2[9] ) );
  NAND4_X2 U12282 ( .A1(\SB2_1_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_28/Component_Function_0/NAND4_in[0] ), .A4(n5190), .ZN(
        \SB2_1_28/buf_output[0] ) );
  XOR2_X1 U12284 ( .A1(\RI5[4][44] ), .A2(\RI5[4][50] ), .Z(
        \MC_ARK_ARC_1_4/temp1[50] ) );
  XOR2_X1 U12285 ( .A1(\MC_ARK_ARC_1_2/temp4[11] ), .A2(
        \MC_ARK_ARC_1_2/temp3[11] ), .Z(\MC_ARK_ARC_1_2/temp6[11] ) );
  XOR2_X1 U12286 ( .A1(\MC_ARK_ARC_1_0/temp2[168] ), .A2(
        \MC_ARK_ARC_1_0/temp1[168] ), .Z(\MC_ARK_ARC_1_0/temp5[168] ) );
  NAND4_X2 U12289 ( .A1(\SB2_1_5/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_5/Component_Function_1/NAND4_in[3] ), .A3(n1769), .A4(
        \SB2_1_5/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_5/buf_output[1] ) );
  XOR2_X1 U12290 ( .A1(\RI5[0][118] ), .A2(\RI5[0][142] ), .Z(
        \MC_ARK_ARC_1_0/temp2[172] ) );
  NAND3_X2 U12291 ( .A1(\SB2_3_16/i0[9] ), .A2(\SB2_3_16/i0_3 ), .A3(
        \SB2_3_16/i0[8] ), .ZN(\SB2_3_16/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U12292 ( .A1(\SB1_0_20/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_20/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_20/Component_Function_1/NAND4_in[0] ), .A4(n5193), .ZN(
        \RI3[0][91] ) );
  NAND3_X1 U12293 ( .A1(\SB1_0_20/i0_4 ), .A2(\SB1_0_20/i1_7 ), .A3(
        \SB1_0_20/i0[8] ), .ZN(n5193) );
  XOR2_X1 U12297 ( .A1(\RI5[0][10] ), .A2(\RI5[0][16] ), .Z(
        \MC_ARK_ARC_1_0/temp1[16] ) );
  XOR2_X1 U12298 ( .A1(n5197), .A2(n5198), .Z(\MC_ARK_ARC_1_1/buf_output[17] )
         );
  XOR2_X1 U12299 ( .A1(\MC_ARK_ARC_1_1/temp2[17] ), .A2(
        \MC_ARK_ARC_1_1/temp4[17] ), .Z(n5197) );
  XOR2_X1 U12300 ( .A1(\MC_ARK_ARC_1_1/temp1[17] ), .A2(n2827), .Z(n5198) );
  NAND3_X1 U12302 ( .A1(\SB1_1_17/i0_0 ), .A2(\SB1_1_17/i3[0] ), .A3(
        \SB1_1_17/i1_7 ), .ZN(\SB1_1_17/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U12303 ( .A1(\MC_ARK_ARC_1_4/temp4[17] ), .A2(n2847), .Z(n5200) );
  XOR2_X1 U12307 ( .A1(\MC_ARK_ARC_1_0/temp2[151] ), .A2(
        \MC_ARK_ARC_1_0/temp1[151] ), .Z(\MC_ARK_ARC_1_0/temp5[151] ) );
  XOR2_X1 U12310 ( .A1(n5201), .A2(n107), .Z(Ciphertext[157]) );
  NAND3_X1 U12313 ( .A1(\SB4_27/i0[6] ), .A2(\SB4_27/i0_3 ), .A3(
        \SB4_27/i1[9] ), .ZN(n5204) );
  XOR2_X1 U12315 ( .A1(n5205), .A2(n6), .Z(Ciphertext[55]) );
  NAND4_X2 U12316 ( .A1(\SB4_22/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_22/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_22/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_22/Component_Function_1/NAND4_in[0] ), .ZN(n5205) );
  NAND3_X1 U12317 ( .A1(\SB3_27/i0_4 ), .A2(\SB3_27/i0[9] ), .A3(
        \SB3_27/i0[6] ), .ZN(\SB3_27/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U12319 ( .A1(\MC_ARK_ARC_1_4/temp3[58] ), .A2(
        \MC_ARK_ARC_1_4/temp4[58] ), .Z(n5206) );
  XOR2_X1 U12323 ( .A1(\RI5[4][137] ), .A2(\RI5[4][101] ), .Z(n5212) );
  NAND3_X2 U12326 ( .A1(\SB1_0_8/i0[10] ), .A2(\SB1_0_8/i1[9] ), .A3(
        \SB1_0_8/i1_5 ), .ZN(n5214) );
  NAND4_X2 U12330 ( .A1(\SB2_1_29/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_29/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_29/Component_Function_2/NAND4_in[1] ), .A4(n5217), .ZN(
        \SB2_1_29/buf_output[2] ) );
  XOR2_X1 U12332 ( .A1(n5219), .A2(\MC_ARK_ARC_1_1/temp4[158] ), .Z(
        \MC_ARK_ARC_1_1/temp6[158] ) );
  NAND4_X2 U12334 ( .A1(\SB2_0_0/Component_Function_0/NAND4_in[1] ), .A2(n2207), .A3(\SB2_0_0/Component_Function_0/NAND4_in[0] ), .A4(n5220), .ZN(
        \SB2_0_0/buf_output[0] ) );
  NAND3_X1 U12335 ( .A1(\SB1_0_10/i0_0 ), .A2(\SB1_0_10/i3[0] ), .A3(
        \SB1_0_10/i1_7 ), .ZN(n5221) );
  XOR2_X1 U12336 ( .A1(\MC_ARK_ARC_1_0/temp4[75] ), .A2(n5222), .Z(n2479) );
  XOR2_X1 U12337 ( .A1(\RI5[0][141] ), .A2(\RI5[0][177] ), .Z(n5222) );
  XOR2_X1 U12338 ( .A1(n1200), .A2(\MC_ARK_ARC_1_0/temp2[93] ), .Z(
        \MC_ARK_ARC_1_0/temp5[93] ) );
  NAND3_X2 U12339 ( .A1(\SB2_2_7/i0[10] ), .A2(\SB2_2_7/i1_7 ), .A3(
        \SB2_2_7/i1[9] ), .ZN(n5223) );
  NAND3_X2 U12340 ( .A1(\SB3_17/i0_3 ), .A2(\SB3_17/i0[8] ), .A3(
        \SB3_17/i0[9] ), .ZN(\SB3_17/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U12342 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[117] ), .A2(\RI5[1][153] ), .Z(n5224) );
  NAND3_X2 U12344 ( .A1(\SB1_2_9/i0_4 ), .A2(\SB1_2_9/i0_3 ), .A3(
        \SB1_2_9/i1[9] ), .ZN(\SB1_2_9/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U12348 ( .A1(\SB1_0_13/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_13/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_13/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_13/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][113] ) );
  NAND3_X1 U12350 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i0[9] ), .A3(
        \SB4_22/i0[8] ), .ZN(\SB4_22/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U12351 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[133] ), .A2(\RI5[2][157] ), .Z(\MC_ARK_ARC_1_2/temp2[187] ) );
  NAND3_X1 U12353 ( .A1(\SB1_3_11/i0_3 ), .A2(\SB1_3_11/i0[6] ), .A3(
        \SB1_3_11/i1[9] ), .ZN(n2134) );
  NAND4_X2 U12354 ( .A1(\SB1_3_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_0/Component_Function_5/NAND4_in[1] ), .A3(n5278), .A4(
        \SB1_3_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_0/buf_output[5] ) );
  INV_X2 U12357 ( .I(\SB1_2_2/buf_output[3] ), .ZN(\SB2_2_0/i0[8] ) );
  NAND4_X2 U12358 ( .A1(\SB1_2_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_2/Component_Function_3/NAND4_in[2] ), .A3(n2725), .A4(n1622), 
        .ZN(\SB1_2_2/buf_output[3] ) );
  NAND3_X1 U12359 ( .A1(\SB4_27/i0[9] ), .A2(\SB4_27/i1_5 ), .A3(
        \SB4_27/i0[6] ), .ZN(\SB4_27/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U12360 ( .A1(n5226), .A2(\MC_ARK_ARC_1_0/temp6[177] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[177] ) );
  XOR2_X1 U12361 ( .A1(\MC_ARK_ARC_1_0/temp2[177] ), .A2(
        \MC_ARK_ARC_1_0/temp1[177] ), .Z(n5226) );
  XOR2_X1 U12364 ( .A1(n1968), .A2(\MC_ARK_ARC_1_1/temp6[175] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[175] ) );
  NAND3_X2 U12367 ( .A1(\RI3[0][70] ), .A2(\SB2_0_20/i0[6] ), .A3(n5264), .ZN(
        n5281) );
  XOR2_X1 U12368 ( .A1(\RI5[0][80] ), .A2(\RI5[0][86] ), .Z(
        \MC_ARK_ARC_1_0/temp1[86] ) );
  NAND4_X2 U12369 ( .A1(n1116), .A2(\SB1_0_8/Component_Function_3/NAND4_in[1] ), .A3(\SB1_0_8/Component_Function_3/NAND4_in[3] ), .A4(n5228), .ZN(
        \RI3[0][153] ) );
  NAND3_X2 U12370 ( .A1(\SB1_0_8/i0[10] ), .A2(\SB1_0_8/i1[9] ), .A3(
        \SB1_0_8/i1_7 ), .ZN(n5228) );
  XOR2_X1 U12373 ( .A1(\MC_ARK_ARC_1_1/temp2[71] ), .A2(
        \MC_ARK_ARC_1_1/temp1[71] ), .Z(n5231) );
  NAND3_X1 U12374 ( .A1(n5429), .A2(\SB2_1_31/i1_7 ), .A3(\SB2_1_31/i0[8] ), 
        .ZN(\SB2_1_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U12376 ( .A1(\SB2_1_21/i0[10] ), .A2(\SB2_1_21/i1_5 ), .A3(
        \SB2_1_21/i1[9] ), .ZN(n5233) );
  NAND4_X2 U12380 ( .A1(n2382), .A2(\SB2_1_8/Component_Function_0/NAND4_in[3] ), .A3(\SB2_1_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_8/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_8/buf_output[0] ) );
  XOR2_X1 U12381 ( .A1(n912), .A2(\MC_ARK_ARC_1_0/temp6[137] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[137] ) );
  XOR2_X1 U12386 ( .A1(\RI5[0][161] ), .A2(\RI5[0][5] ), .Z(n5242) );
  XOR2_X1 U12387 ( .A1(n5244), .A2(n5243), .Z(\MC_ARK_ARC_1_3/temp6[23] ) );
  XOR2_X1 U12388 ( .A1(\RI5[3][125] ), .A2(n193), .Z(n5243) );
  NAND3_X2 U12389 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i0_0 ), .A3(
        \SB2_2_3/i0[7] ), .ZN(n5245) );
  INV_X2 U12393 ( .I(\SB1_4_15/buf_output[3] ), .ZN(\SB2_4_13/i0[8] ) );
  NAND3_X1 U12395 ( .A1(n6272), .A2(\SB4_9/i0_3 ), .A3(\SB4_9/i1[9] ), .ZN(
        n5249) );
  NAND3_X1 U12397 ( .A1(\SB2_4_8/i0_3 ), .A2(\SB2_4_8/i0[10] ), .A3(n3183), 
        .ZN(\SB2_4_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U12398 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i0[10] ), .A3(\SB4_2/i0_4 ), 
        .ZN(n5250) );
  XOR2_X1 U12399 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[168] ), .A2(\RI5[4][174] ), .Z(\MC_ARK_ARC_1_4/temp1[174] ) );
  XOR2_X1 U12400 ( .A1(\MC_ARK_ARC_1_0/temp2[72] ), .A2(
        \MC_ARK_ARC_1_0/temp1[72] ), .Z(\MC_ARK_ARC_1_0/temp5[72] ) );
  INV_X2 U12404 ( .I(\SB1_3_6/buf_output[3] ), .ZN(\SB2_3_4/i0[8] ) );
  XOR2_X1 U12405 ( .A1(n5257), .A2(n81), .Z(Ciphertext[139]) );
  NAND3_X1 U12406 ( .A1(\SB4_0/i0[10] ), .A2(\SB4_0/i1[9] ), .A3(\SB4_0/i1_7 ), 
        .ZN(n5258) );
  NAND4_X2 U12407 ( .A1(\SB2_4_18/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_4_18/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_4_18/Component_Function_4/NAND4_in[0] ), .A4(n5259), .ZN(
        \SB2_4_18/buf_output[4] ) );
  NAND4_X2 U12408 ( .A1(n675), .A2(\SB2_2_22/Component_Function_2/NAND4_in[0] ), .A3(n2017), .A4(\SB2_2_22/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_22/buf_output[2] ) );
  XOR2_X1 U12409 ( .A1(\RI5[0][11] ), .A2(\RI5[0][17] ), .Z(
        \MC_ARK_ARC_1_0/temp1[17] ) );
  NAND3_X1 U12410 ( .A1(\SB2_0_30/i0[6] ), .A2(\SB2_0_30/i0_0 ), .A3(
        \SB2_0_30/i0[10] ), .ZN(\SB2_0_30/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U12411 ( .A1(\SB1_3_1/i0_3 ), .A2(\SB1_3_1/i0_0 ), .A3(
        \SB1_3_1/i0[7] ), .ZN(n2971) );
  NAND3_X2 U12412 ( .A1(\SB2_2_16/i0[10] ), .A2(\SB2_2_16/i0_0 ), .A3(
        \SB2_2_16/i0[6] ), .ZN(\SB2_2_16/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U12413 ( .A1(n1739), .A2(n5261), .Z(n2936) );
  XOR2_X1 U12415 ( .A1(\RI5[0][5] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[41] ), 
        .Z(n5262) );
  XOR2_X1 U12416 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[41] ), .A2(\RI5[2][17] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[71] ) );
  INV_X2 U12419 ( .I(\SB1_2_15/buf_output[2] ), .ZN(\SB2_2_12/i1[9] ) );
  NAND4_X2 U12420 ( .A1(\SB1_2_15/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_2_15/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_15/Component_Function_2/NAND4_in[1] ), .A4(n2089), .ZN(
        \SB1_2_15/buf_output[2] ) );
  NAND3_X1 U12423 ( .A1(\SB2_3_10/i1_7 ), .A2(\SB2_3_10/i0[8] ), .A3(
        \SB2_3_10/i0_4 ), .ZN(n1625) );
  XOR2_X1 U12424 ( .A1(n5267), .A2(\MC_ARK_ARC_1_0/temp4[105] ), .Z(n1973) );
  XOR2_X1 U12425 ( .A1(\RI5[0][15] ), .A2(\RI5[0][171] ), .Z(n5267) );
  XOR2_X1 U12426 ( .A1(n2509), .A2(n5268), .Z(\MC_ARK_ARC_1_0/buf_output[117] ) );
  INV_X4 U12430 ( .I(\SB2_3_20/i0[7] ), .ZN(\RI3[3][70] ) );
  NOR2_X2 U12432 ( .A1(n5272), .A2(n5271), .ZN(\SB2_3_20/i0[7] ) );
  NAND4_X2 U12433 ( .A1(\SB1_3_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_21/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_3_21/Component_Function_0/NAND4_in[1] ), .A4(n5273), .ZN(
        \SB1_3_21/buf_output[0] ) );
  NAND3_X1 U12434 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0[7] ), .A3(
        \SB1_3_21/i0_0 ), .ZN(n5273) );
  NAND4_X2 U12439 ( .A1(\SB2_2_17/Component_Function_4/NAND4_in[0] ), .A2(
        n1387), .A3(\SB2_2_17/Component_Function_4/NAND4_in[3] ), .A4(n5276), 
        .ZN(\SB2_2_17/buf_output[4] ) );
  NAND3_X1 U12440 ( .A1(\SB2_2_17/i0_0 ), .A2(\SB2_2_17/i3[0] ), .A3(
        \SB2_2_17/i1_7 ), .ZN(n5276) );
  NAND3_X1 U12441 ( .A1(\SB1_3_11/i0_4 ), .A2(\SB1_3_11/i1_7 ), .A3(
        \SB1_3_11/i0[8] ), .ZN(\SB1_3_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U12442 ( .A1(\SB1_2_14/i0_4 ), .A2(\SB1_2_14/i1_7 ), .A3(
        \SB1_2_14/i0[8] ), .ZN(n5277) );
  XOR2_X1 U12443 ( .A1(n5279), .A2(n124), .Z(Ciphertext[154]) );
  XOR2_X1 U12449 ( .A1(\MC_ARK_ARC_1_2/temp1[56] ), .A2(
        \MC_ARK_ARC_1_2/temp4[56] ), .Z(n5282) );
  NAND4_X2 U12451 ( .A1(\SB1_1_8/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_8/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_8/Component_Function_2/NAND4_in[2] ), .A4(n5284), .ZN(
        \SB1_1_8/buf_output[2] ) );
  NAND3_X2 U12455 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i0_0 ), .A3(
        \SB2_1_5/i0[7] ), .ZN(n5285) );
  NAND4_X2 U12457 ( .A1(\SB2_1_17/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_17/Component_Function_0/NAND4_in[0] ), .A4(n5287), .ZN(
        \SB2_1_17/buf_output[0] ) );
  XOR2_X1 U12458 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[32] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[188] ), .Z(n5288) );
  NAND3_X1 U12459 ( .A1(\SB2_2_6/i0_0 ), .A2(\SB2_2_6/i0[9] ), .A3(
        \SB2_2_6/i0[8] ), .ZN(\SB2_2_6/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 U12460 ( .A1(\SB1_0_7/i1[9] ), .A2(\SB1_0_7/i0_3 ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[0] ) );
  XOR2_X1 U12462 ( .A1(\RI5[4][35] ), .A2(\RI5[4][29] ), .Z(
        \MC_ARK_ARC_1_4/temp1[35] ) );
  NAND4_X2 U12464 ( .A1(\SB1_0_31/Component_Function_0/NAND4_in[2] ), .A2(n634), .A3(\SB1_0_31/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_31/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][30] ) );
  NAND4_X2 U12466 ( .A1(\SB3_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_2/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_2/Component_Function_0/NAND4_in[1] ), .A4(n5290), .ZN(
        \SB3_2/buf_output[0] ) );
  NAND3_X2 U12467 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i0[7] ), .A3(\SB3_2/i0_0 ), 
        .ZN(n5290) );
  XOR2_X1 U12468 ( .A1(\MC_ARK_ARC_1_0/temp2[137] ), .A2(n945), .Z(n912) );
  NAND4_X2 U12469 ( .A1(\SB2_2_26/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_26/Component_Function_4/NAND4_in[0] ), .A4(n5291), .ZN(
        \SB2_2_26/buf_output[4] ) );
  XOR2_X1 U12471 ( .A1(\MC_ARK_ARC_1_3/temp1[85] ), .A2(n5293), .Z(
        \MC_ARK_ARC_1_3/temp5[85] ) );
  XOR2_X1 U12472 ( .A1(\RI5[3][31] ), .A2(\RI5[3][55] ), .Z(n5293) );
  XOR2_X1 U12473 ( .A1(n5294), .A2(\MC_ARK_ARC_1_3/temp5[162] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[162] ) );
  XOR2_X1 U12474 ( .A1(\MC_ARK_ARC_1_3/temp4[162] ), .A2(
        \MC_ARK_ARC_1_3/temp3[162] ), .Z(n5294) );
  NAND3_X1 U12475 ( .A1(\SB1_4_14/i1[9] ), .A2(\SB1_4_14/i0[10] ), .A3(
        \SB1_4_14/i1_5 ), .ZN(\SB1_4_14/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U12477 ( .A1(\RI5[3][145] ), .A2(\RI5[3][169] ), .Z(n5295) );
  NAND3_X1 U12479 ( .A1(\SB1_3_25/i0_3 ), .A2(\SB1_3_25/i0_0 ), .A3(
        \SB1_3_25/i0[7] ), .ZN(n739) );
  NAND3_X1 U12480 ( .A1(\SB3_15/i0[9] ), .A2(\SB3_15/i0[10] ), .A3(
        \SB3_15/i0_3 ), .ZN(\SB3_15/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U12481 ( .A1(\MC_ARK_ARC_1_4/temp1[35] ), .A2(
        \MC_ARK_ARC_1_4/temp4[35] ), .Z(n5300) );
  XOR2_X1 U12482 ( .A1(n5302), .A2(\MC_ARK_ARC_1_2/temp4[129] ), .Z(n1776) );
  INV_X2 U12483 ( .I(\SB1_2_7/buf_output[3] ), .ZN(\SB2_2_5/i0[8] ) );
  NAND3_X1 U12486 ( .A1(\SB4_28/i1_5 ), .A2(\SB4_28/i3[0] ), .A3(
        \SB4_28/i0[8] ), .ZN(n5303) );
  NAND3_X1 U12487 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i1_5 ), .A3(
        \SB4_28/i1[9] ), .ZN(n5304) );
  INV_X1 U12488 ( .I(\SB3_29/buf_output[5] ), .ZN(\SB4_29/i1_5 ) );
  NAND4_X2 U12489 ( .A1(\SB3_29/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_29/Component_Function_5/NAND4_in[2] ), .A3(
        \SB3_29/Component_Function_5/NAND4_in[3] ), .A4(
        \SB3_29/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_29/buf_output[5] ) );
  NAND4_X2 U12490 ( .A1(\SB3_24/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_24/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_24/Component_Function_4/NAND4_in[3] ), .A4(n5305), .ZN(
        \SB3_24/buf_output[4] ) );
  NAND4_X2 U12491 ( .A1(\SB1_4_15/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_4_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_15/Component_Function_1/NAND4_in[0] ), .A4(n5306), .ZN(
        \SB1_4_15/buf_output[1] ) );
  NAND3_X1 U12497 ( .A1(\SB1_3_0/i0[6] ), .A2(\SB1_3_0/i0_3 ), .A3(
        \SB1_3_0/i1[9] ), .ZN(\SB1_3_0/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12498 ( .A1(\RI5[0][47] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[71] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[101] ) );
  NAND4_X2 U12499 ( .A1(\SB1_4_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_4_8/Component_Function_3/NAND4_in[2] ), .A3(n3013), .A4(n5311), 
        .ZN(\SB1_4_8/buf_output[3] ) );
  NAND3_X1 U12500 ( .A1(\SB2_0_3/i0_3 ), .A2(\SB2_0_3/i0[10] ), .A3(
        \RI3[0][172] ), .ZN(\SB2_0_3/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U12503 ( .A1(\MC_ARK_ARC_1_0/temp1[60] ), .A2(
        \MC_ARK_ARC_1_0/temp2[60] ), .Z(n5313) );
  XOR2_X1 U12504 ( .A1(n5314), .A2(\MC_ARK_ARC_1_0/temp4[102] ), .Z(n2776) );
  XOR2_X1 U12505 ( .A1(\RI5[0][72] ), .A2(\RI5[0][48] ), .Z(n5314) );
  XOR2_X1 U12507 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[177] ), .A2(\RI5[4][21] ), 
        .Z(n5316) );
  XOR2_X1 U12509 ( .A1(n5318), .A2(\MC_ARK_ARC_1_1/temp2[144] ), .Z(
        \MC_ARK_ARC_1_1/temp5[144] ) );
  XOR2_X1 U12510 ( .A1(\RI5[1][138] ), .A2(\RI5[1][144] ), .Z(n5318) );
  XOR2_X1 U12511 ( .A1(n2411), .A2(\MC_ARK_ARC_1_2/temp2[57] ), .Z(n5319) );
  XOR2_X1 U12512 ( .A1(n575), .A2(\MC_ARK_ARC_1_3/buf_datainput[99] ), .Z(
        n5320) );
  NAND3_X1 U12513 ( .A1(\SB3_3/i0_4 ), .A2(\SB3_3/i1_7 ), .A3(\SB3_3/i0[8] ), 
        .ZN(\SB3_3/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U12514 ( .A1(\MC_ARK_ARC_1_4/temp6[172] ), .A2(
        \MC_ARK_ARC_1_4/temp5[172] ), .Z(\MC_ARK_ARC_1_4/buf_output[172] ) );
  NAND3_X1 U12516 ( .A1(\SB1_0_7/i1[9] ), .A2(\SB1_0_7/i0[10] ), .A3(
        \SB1_0_7/i1_5 ), .ZN(\SB1_0_7/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U12518 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[60] ), .A2(\RI5[2][66] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[66] ) );
  XOR2_X1 U12522 ( .A1(\RI5[3][190] ), .A2(\RI5[3][34] ), .Z(n5323) );
  NAND3_X2 U12523 ( .A1(\SB2_0_20/i0_3 ), .A2(\RI3[0][70] ), .A3(
        \SB2_0_20/i1[9] ), .ZN(n5324) );
  NAND4_X2 U12524 ( .A1(\SB2_3_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_16/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_3_16/Component_Function_2/NAND4_in[1] ), .A4(n5325), .ZN(
        \SB2_3_16/buf_output[2] ) );
  NAND3_X2 U12525 ( .A1(\SB2_3_16/i0_0 ), .A2(\SB2_3_16/i0_4 ), .A3(n571), 
        .ZN(n5325) );
  NAND3_X1 U12526 ( .A1(\SB2_2_3/i0[6] ), .A2(\SB1_2_4/buf_output[4] ), .A3(
        \SB2_2_3/i0[9] ), .ZN(n5326) );
  XOR2_X1 U12527 ( .A1(n5328), .A2(n5327), .Z(\MC_ARK_ARC_1_2/buf_output[88] )
         );
  XOR2_X1 U12528 ( .A1(\MC_ARK_ARC_1_2/temp2[88] ), .A2(
        \MC_ARK_ARC_1_2/temp1[88] ), .Z(n5327) );
  XOR2_X1 U12529 ( .A1(\MC_ARK_ARC_1_2/temp4[88] ), .A2(
        \MC_ARK_ARC_1_2/temp3[88] ), .Z(n5328) );
  NAND4_X2 U12534 ( .A1(\SB2_2_18/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_18/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_18/Component_Function_4/NAND4_in[1] ), .A4(n5331), .ZN(
        \SB2_2_18/buf_output[4] ) );
  NAND3_X1 U12535 ( .A1(\SB2_3_1/i0_0 ), .A2(\SB2_3_1/i3[0] ), .A3(
        \SB2_3_1/i1_7 ), .ZN(\SB2_3_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U12537 ( .A1(\SB2_3_3/i0[8] ), .A2(\SB2_3_3/i3[0] ), .A3(
        \SB2_3_3/i1_5 ), .ZN(n5332) );
  NAND3_X1 U12538 ( .A1(\RI3[0][140] ), .A2(\SB2_0_8/i0_3 ), .A3(\RI3[0][142] ), .ZN(\SB2_0_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U12541 ( .A1(\SB3_5/i0[6] ), .A2(\SB3_5/i1_5 ), .A3(\SB3_5/i0[9] ), 
        .ZN(\SB3_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U12543 ( .A1(\SB3_26/i0[10] ), .A2(\SB3_26/i0_3 ), .A3(
        \SB3_26/i0_4 ), .ZN(n5335) );
  NAND3_X1 U12546 ( .A1(\SB1_0_7/i0_0 ), .A2(\SB1_0_7/i1_5 ), .A3(
        \SB1_0_7/i0_4 ), .ZN(n5338) );
  XOR2_X1 U12553 ( .A1(\MC_ARK_ARC_1_2/temp1[141] ), .A2(
        \MC_ARK_ARC_1_2/temp2[141] ), .Z(\MC_ARK_ARC_1_2/temp5[141] ) );
  NAND3_X1 U12554 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0_0 ), .A3(
        \SB2_2_25/i0[7] ), .ZN(n5339) );
  NAND3_X1 U12555 ( .A1(\SB2_2_25/i0[10] ), .A2(\SB2_2_25/i0_3 ), .A3(
        \SB2_2_25/i0_4 ), .ZN(n5340) );
  XOR2_X1 U12558 ( .A1(n5342), .A2(\MC_ARK_ARC_1_2/temp4[121] ), .Z(
        \MC_ARK_ARC_1_2/temp6[121] ) );
  XOR2_X1 U12559 ( .A1(\RI5[2][187] ), .A2(\RI5[2][31] ), .Z(n5342) );
  NAND4_X2 U12563 ( .A1(\SB2_1_11/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_0/NAND4_in[0] ), .A4(n5344), .ZN(
        \SB2_1_11/buf_output[0] ) );
  NOR2_X2 U12564 ( .A1(n1775), .A2(n5345), .ZN(n1427) );
  XOR2_X1 U12566 ( .A1(\MC_ARK_ARC_1_0/temp6[183] ), .A2(n2788), .Z(
        \MC_ARK_ARC_1_0/buf_output[183] ) );
  NAND3_X1 U12569 ( .A1(\SB3_13/i0_4 ), .A2(\SB3_13/i1_7 ), .A3(\SB3_13/i0[8] ), .ZN(n2399) );
  NAND3_X1 U12570 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i0[10] ), .A3(\SB4_8/i0[6] ), 
        .ZN(n5346) );
  NAND3_X1 U12571 ( .A1(\SB3_7/i0_3 ), .A2(\SB3_7/i0_0 ), .A3(\SB3_7/i0_4 ), 
        .ZN(\SB3_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U12573 ( .A1(\SB1_4_6/i0[6] ), .A2(\SB1_4_6/i0[8] ), .A3(
        \SB1_4_6/i0[7] ), .ZN(\SB1_4_6/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U12574 ( .A1(\SB1_1_29/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_29/Component_Function_0/NAND4_in[0] ), .A4(n5348), .ZN(
        \SB1_1_29/buf_output[0] ) );
  NAND3_X1 U12576 ( .A1(\SB1_4_30/i0[9] ), .A2(\SB1_4_30/i1_5 ), .A3(
        \SB1_4_30/i0[6] ), .ZN(\SB1_4_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U12577 ( .A1(\SB3_7/i0_3 ), .A2(\SB3_7/i0[9] ), .A3(\SB3_7/i0[10] ), 
        .ZN(\SB3_7/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U12580 ( .A1(\MC_ARK_ARC_1_0/temp4[85] ), .A2(
        \MC_ARK_ARC_1_0/temp3[85] ), .Z(\MC_ARK_ARC_1_0/temp6[85] ) );
  XOR2_X1 U12583 ( .A1(\MC_ARK_ARC_1_0/temp6[19] ), .A2(
        \MC_ARK_ARC_1_0/temp5[19] ), .Z(\MC_ARK_ARC_1_0/buf_output[19] ) );
  XOR2_X1 U12585 ( .A1(\RI5[0][178] ), .A2(\RI5[0][142] ), .Z(
        \MC_ARK_ARC_1_0/temp3[76] ) );
  XOR2_X1 U12586 ( .A1(\RI5[1][92] ), .A2(\RI5[1][56] ), .Z(
        \MC_ARK_ARC_1_1/temp3[182] ) );
  XOR2_X1 U12587 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[24] ), .A2(n567), .Z(
        n5353) );
  XOR2_X1 U12589 ( .A1(\MC_ARK_ARC_1_1/temp1[122] ), .A2(n5355), .Z(
        \MC_ARK_ARC_1_1/temp5[122] ) );
  XOR2_X1 U12590 ( .A1(\RI5[1][68] ), .A2(\RI5[1][92] ), .Z(n5355) );
  NAND3_X1 U12591 ( .A1(\SB1_4_12/i0_0 ), .A2(\SB1_4_12/i1_7 ), .A3(
        \SB1_4_12/i3[0] ), .ZN(\SB1_4_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U12593 ( .A1(\SB1_1_2/i1[9] ), .A2(\SB1_1_2/i0_4 ), .A3(
        \SB1_1_2/i1_5 ), .ZN(n2507) );
  INV_X2 U12594 ( .I(\SB1_2_29/buf_output[3] ), .ZN(\SB2_2_27/i0[8] ) );
  XOR2_X1 U12595 ( .A1(\MC_ARK_ARC_1_1/temp1[13] ), .A2(
        \MC_ARK_ARC_1_1/temp2[13] ), .Z(\MC_ARK_ARC_1_1/temp5[13] ) );
  XOR2_X1 U12596 ( .A1(\MC_ARK_ARC_1_1/temp1[15] ), .A2(
        \MC_ARK_ARC_1_1/temp2[15] ), .Z(n2761) );
  NAND4_X2 U12597 ( .A1(\SB1_3_20/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_20/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_20/Component_Function_1/NAND4_in[0] ), .A4(n5356), .ZN(
        \SB1_3_20/buf_output[1] ) );
  NAND4_X2 U12599 ( .A1(\SB3_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_4/NAND4_in[3] ), .A4(n5358), .ZN(
        \SB3_17/buf_output[4] ) );
  NAND3_X1 U12600 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i0_0 ), .A3(
        \SB2_3_24/i0_4 ), .ZN(\SB2_3_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U12603 ( .A1(\SB2_1_31/i0[7] ), .A2(\SB2_1_31/i0[8] ), .A3(
        \SB2_1_31/i0[6] ), .ZN(\SB2_1_31/Component_Function_0/NAND4_in[1] ) );
  INV_X2 U12604 ( .I(\SB1_4_0/buf_output[3] ), .ZN(\SB2_4_30/i0[8] ) );
  XOR2_X1 U12607 ( .A1(\RI5[4][186] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[18] ), 
        .Z(n5362) );
  XOR2_X1 U12608 ( .A1(\MC_ARK_ARC_1_3/temp4[106] ), .A2(n5363), .Z(
        \MC_ARK_ARC_1_3/temp6[106] ) );
  XOR2_X1 U12609 ( .A1(\RI5[3][172] ), .A2(\RI5[3][16] ), .Z(n5363) );
  NAND4_X2 U12610 ( .A1(\SB2_2_24/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_24/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_24/Component_Function_4/NAND4_in[1] ), .A4(n5365), .ZN(
        \SB2_2_24/buf_output[4] ) );
  NAND3_X1 U12611 ( .A1(\SB1_1_23/i0[6] ), .A2(\SB1_1_23/i1[9] ), .A3(
        \SB1_1_23/i0_3 ), .ZN(\SB1_1_23/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12612 ( .A1(n1161), .A2(\MC_ARK_ARC_1_0/temp6[49] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[49] ) );
  NAND3_X1 U12613 ( .A1(\SB3_9/buf_output[3] ), .A2(\SB4_7/i1_5 ), .A3(
        \SB4_7/i1[9] ), .ZN(n5367) );
  XOR2_X1 U12615 ( .A1(n5370), .A2(\MC_ARK_ARC_1_1/buf_keyinput[111] ), .Z(
        Ciphertext[127]) );
  XOR2_X1 U12617 ( .A1(n1066), .A2(\MC_ARK_ARC_1_3/temp5[75] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[75] ) );
  XOR2_X1 U12618 ( .A1(\MC_ARK_ARC_1_2/temp1[151] ), .A2(
        \MC_ARK_ARC_1_2/temp2[151] ), .Z(\MC_ARK_ARC_1_2/temp5[151] ) );
  XOR2_X1 U12621 ( .A1(n5372), .A2(n41), .Z(Ciphertext[125]) );
  NAND4_X2 U12622 ( .A1(\SB4_11/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_11/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_11/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_11/Component_Function_5/NAND4_in[0] ), .ZN(n5372) );
  XOR2_X1 U12624 ( .A1(\MC_ARK_ARC_1_2/temp1[145] ), .A2(
        \MC_ARK_ARC_1_2/temp2[145] ), .Z(n5375) );
  NAND3_X1 U12625 ( .A1(\SB1_0_19/i0_3 ), .A2(\SB1_0_19/i0[8] ), .A3(
        \SB1_0_19/i1_7 ), .ZN(\SB1_0_19/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U12626 ( .A1(\SB2_0_8/i0_0 ), .A2(\SB2_0_8/i1_5 ), .A3(
        \RI3[0][142] ), .ZN(\SB2_0_8/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U12631 ( .A1(\MC_ARK_ARC_1_1/temp2[61] ), .A2(
        \MC_ARK_ARC_1_1/temp1[61] ), .Z(\MC_ARK_ARC_1_1/temp5[61] ) );
  NAND3_X2 U12632 ( .A1(\SB2_2_4/i0[9] ), .A2(\SB2_2_4/i0_4 ), .A3(
        \SB2_2_4/i0[6] ), .ZN(n5379) );
  NAND3_X1 U12633 ( .A1(\SB1_1_13/i0_0 ), .A2(\SB1_1_13/i0[8] ), .A3(
        \SB1_1_13/i0[9] ), .ZN(\SB1_1_13/Component_Function_4/NAND4_in[0] ) );
  INV_X2 U12634 ( .I(\SB1_4_16/buf_output[2] ), .ZN(\SB2_4_13/i1[9] ) );
  XOR2_X1 U12635 ( .A1(\MC_ARK_ARC_1_0/temp5[111] ), .A2(
        \MC_ARK_ARC_1_0/temp6[111] ), .Z(\MC_ARK_ARC_1_0/buf_output[111] ) );
  XOR2_X1 U12636 ( .A1(\RI5[1][93] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[117] ), 
        .Z(n5380) );
  NAND3_X1 U12637 ( .A1(\SB1_0_24/i0_0 ), .A2(\SB1_0_24/i1_5 ), .A3(
        \SB1_0_24/i0_4 ), .ZN(n5381) );
  XOR2_X1 U12640 ( .A1(\MC_ARK_ARC_1_0/temp2[175] ), .A2(
        \MC_ARK_ARC_1_0/temp1[175] ), .Z(\MC_ARK_ARC_1_0/temp5[175] ) );
  NAND2_X2 U12641 ( .A1(\SB1_1_25/i0_0 ), .A2(\SB1_1_25/i3[0] ), .ZN(n5383) );
  XOR2_X1 U12646 ( .A1(n1436), .A2(n5387), .Z(\MC_ARK_ARC_1_1/buf_output[128] ) );
  XOR2_X1 U12647 ( .A1(\MC_ARK_ARC_1_1/temp3[128] ), .A2(
        \MC_ARK_ARC_1_1/temp4[128] ), .Z(n5387) );
  NAND3_X1 U12648 ( .A1(\SB4_22/i0[8] ), .A2(\SB4_22/i1_5 ), .A3(
        \SB4_22/i3[0] ), .ZN(\SB4_22/Component_Function_3/NAND4_in[3] ) );
  NAND4_X1 U12649 ( .A1(\SB2_0_14/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_14/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_0_14/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_14/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_0_14/buf_output[1] ) );
  NAND2_X2 U12650 ( .A1(\SB1_0_19/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_0_19/Component_Function_0/NAND4_in[0] ), .ZN(n5388) );
  XOR2_X1 U12651 ( .A1(\SB2_4_14/buf_output[3] ), .A2(\SB2_4_13/buf_output[3] ), .Z(\MC_ARK_ARC_1_4/temp1[123] ) );
  XOR2_X1 U12653 ( .A1(n3011), .A2(n5389), .Z(\MC_ARK_ARC_1_2/buf_output[39] )
         );
  AND2_X1 U12654 ( .A1(\SB2_2_9/Component_Function_1/NAND4_in[2] ), .A2(n5390), 
        .Z(n955) );
  NAND3_X1 U12658 ( .A1(\SB1_0_2/i0_0 ), .A2(\SB1_0_2/i0[9] ), .A3(
        \SB1_0_2/i0[8] ), .ZN(\SB1_0_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U12659 ( .A1(\SB2_1_20/i0_3 ), .A2(\SB2_1_20/i0[6] ), .A3(
        \SB2_1_20/i1[9] ), .ZN(n5396) );
  NAND3_X1 U12661 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i1[9] ), .A3(
        \SB4_17/i0[6] ), .ZN(\SB4_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U12662 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i0[10] ), .A3(
        \SB4_17/i0_4 ), .ZN(n5397) );
  XOR2_X1 U12664 ( .A1(n1753), .A2(\MC_ARK_ARC_1_1/temp6[25] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[25] ) );
  NAND3_X2 U12668 ( .A1(\SB2_4_12/i0_0 ), .A2(\SB2_4_12/i0[10] ), .A3(
        \SB2_4_12/i0[6] ), .ZN(n5402) );
  XOR2_X1 U12671 ( .A1(\RI5[2][59] ), .A2(\RI5[2][83] ), .Z(n750) );
  XOR2_X1 U12673 ( .A1(\MC_ARK_ARC_1_4/temp5[49] ), .A2(n5405), .Z(
        \MC_ARK_ARC_1_4/buf_output[49] ) );
  XOR2_X1 U12674 ( .A1(\MC_ARK_ARC_1_4/temp4[49] ), .A2(
        \MC_ARK_ARC_1_4/temp3[49] ), .Z(n5405) );
  NAND2_X2 U12675 ( .A1(\SB2_2_0/i0_0 ), .A2(\SB2_2_0/i3[0] ), .ZN(n5406) );
  XOR2_X1 U12676 ( .A1(\RI5[3][101] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .Z(n5408) );
  XOR2_X1 U12677 ( .A1(\RI5[4][40] ), .A2(\RI5[4][34] ), .Z(n5410) );
  NAND3_X2 U12678 ( .A1(\SB1_2_2/i0_4 ), .A2(\SB1_2_2/i0[9] ), .A3(
        \SB1_2_2/i0[6] ), .ZN(\SB1_2_2/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U12683 ( .A1(n578), .A2(\RI5[1][148] ), .Z(
        \MC_ARK_ARC_1_1/temp2[10] ) );
  INV_X2 U12684 ( .I(\RI3[0][183] ), .ZN(\SB2_0_1/i0[8] ) );
  NAND3_X1 U12686 ( .A1(\SB1_0_19/i0[8] ), .A2(\SB1_0_19/i1_5 ), .A3(
        \SB1_0_19/i3[0] ), .ZN(\SB1_0_19/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U12690 ( .A1(n5414), .A2(\MC_ARK_ARC_1_4/temp5[73] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[73] ) );
  XOR2_X1 U12691 ( .A1(\MC_ARK_ARC_1_4/temp4[73] ), .A2(
        \MC_ARK_ARC_1_4/temp3[73] ), .Z(n5414) );
  XOR2_X1 U12694 ( .A1(\RI5[1][158] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[164] ), .Z(\MC_ARK_ARC_1_1/temp1[164] ) );
  XOR2_X1 U12695 ( .A1(\MC_ARK_ARC_1_1/temp3[62] ), .A2(
        \MC_ARK_ARC_1_1/temp4[62] ), .Z(\MC_ARK_ARC_1_1/temp6[62] ) );
  XOR2_X1 U12702 ( .A1(\RI5[4][109] ), .A2(\RI5[4][103] ), .Z(
        \MC_ARK_ARC_1_4/temp1[109] ) );
  XOR2_X1 U12704 ( .A1(\RI5[0][73] ), .A2(\RI5[0][109] ), .Z(
        \MC_ARK_ARC_1_0/temp3[7] ) );
  NAND3_X1 U12706 ( .A1(\SB4_26/i0_4 ), .A2(\SB4_26/i1_5 ), .A3(
        \SB3_29/buf_output[2] ), .ZN(n5421) );
  CLKBUF_X12 U12708 ( .I(Key[123]), .Z(n161) );
  AND2_X1 U12709 ( .A1(\SB1_3_14/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_3_14/Component_Function_4/NAND4_in[1] ), .Z(n5423) );
  NAND3_X2 U1417 ( .A1(\SB2_2_12/i0_4 ), .A2(\SB2_2_12/i1_5 ), .A3(
        \SB2_2_12/i1[9] ), .ZN(n3688) );
  NAND2_X2 \SB2_1_30/Component_Function_1/N1  ( .A1(\SB2_1_30/i0_3 ), .A2(
        \SB2_1_30/i1[9] ), .ZN(\SB2_1_30/Component_Function_1/NAND4_in[0] ) );
  NAND2_X2 \SB2_3_25/Component_Function_5/N1  ( .A1(\SB2_3_25/i0_0 ), .A2(
        \SB2_3_25/i3[0] ), .ZN(\SB2_3_25/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U2266 ( .I(\SB1_2_6/buf_output[4] ), .Z(\SB2_2_5/i0_4 ) );
  NAND3_X2 U2884 ( .A1(\SB2_3_8/i0[10] ), .A2(\SB2_3_8/i0[6] ), .A3(
        \SB2_3_8/i0_0 ), .ZN(\SB2_3_8/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB1_3_10/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[128] ), .ZN(
        \SB1_3_10/i1[9] ) );
  BUF_X4 U3400 ( .I(\SB1_4_3/buf_output[0] ), .Z(\SB2_4_30/i0[9] ) );
  NAND3_X2 U1687 ( .A1(\SB2_1_3/i0[6] ), .A2(\SB2_1_3/i0_3 ), .A3(
        \SB2_1_3/i1[9] ), .ZN(n3472) );
  NAND3_X2 U6658 ( .A1(\SB1_1_21/i0[6] ), .A2(\SB1_1_21/i0_3 ), .A3(
        \SB1_1_21/i0[10] ), .ZN(\SB1_1_21/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X2 U1609 ( .A1(\SB1_0_0/i0[10] ), .A2(\SB1_0_0/i0_0 ), .A3(
        \SB1_0_0/i0[6] ), .ZN(\SB1_0_0/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB2_2_8/INV_5  ( .I(\SB1_2_8/buf_output[5] ), .ZN(\SB2_2_8/i1_5 ) );
  NAND3_X2 U9874 ( .A1(\RI1[4][131] ), .A2(\SB1_4_10/i0[10] ), .A3(
        \SB1_4_10/i0_4 ), .ZN(n4033) );
  INV_X2 \SB2_1_0/INV_1  ( .I(\SB1_1_4/buf_output[1] ), .ZN(\SB2_1_0/i1_7 ) );
  NAND3_X2 U3680 ( .A1(\SB2_1_3/i1[9] ), .A2(\SB2_1_3/i1_5 ), .A3(
        \SB2_1_3/i0_4 ), .ZN(\SB2_1_3/Component_Function_4/NAND4_in[3] ) );
  NAND2_X2 U1607 ( .A1(\SB1_0_0/i0[10] ), .A2(\SB1_0_0/i0[9] ), .ZN(
        \SB1_0_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 \SB2_4_5/Component_Function_2/N3  ( .A1(\SB2_4_5/i0_3 ), .A2(
        \SB2_4_5/i0[8] ), .A3(\SB2_4_5/i0[9] ), .ZN(
        \SB2_4_5/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB3_29/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[14] ), .ZN(
        \SB3_29/i1[9] ) );
  INV_X2 \SB2_1_3/INV_1  ( .I(\SB1_1_7/buf_output[1] ), .ZN(\SB2_1_3/i1_7 ) );
  NAND3_X2 U722 ( .A1(\SB2_4_14/i0_3 ), .A2(\SB2_4_14/i0_0 ), .A3(
        \SB2_4_14/i0_4 ), .ZN(\SB2_4_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U3434 ( .A1(\SB2_2_28/i0[10] ), .A2(\SB2_2_28/i1_7 ), .A3(
        \SB2_2_28/i1[9] ), .ZN(n922) );
  NAND3_X2 \SB2_0_25/Component_Function_3/N3  ( .A1(\SB2_0_25/i1[9] ), .A2(
        \SB2_0_25/i1_7 ), .A3(\SB2_0_25/i0[10] ), .ZN(
        \SB2_0_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U965 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i1[9] ), .A3(
        \SB2_2_14/i0_4 ), .ZN(n3114) );
  BUF_X4 \SB2_3_1/BUF_1  ( .I(\SB1_3_5/buf_output[1] ), .Z(\SB2_3_1/i0[6] ) );
  INV_X2 \SB2_3_15/INV_1  ( .I(\SB1_3_19/buf_output[1] ), .ZN(\SB2_3_15/i1_7 )
         );
  INV_X2 U3163 ( .I(\SB1_2_21/buf_output[5] ), .ZN(\SB2_2_21/i1_5 ) );
  INV_X2 U5341 ( .I(\SB1_0_30/buf_output[2] ), .ZN(\SB2_0_27/i1[9] ) );
  NAND3_X2 U2939 ( .A1(\SB1_1_22/i0[9] ), .A2(\SB1_1_22/i1_5 ), .A3(
        \SB1_1_22/i0[6] ), .ZN(\SB1_1_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U5877 ( .A1(\SB2_2_9/i0_3 ), .A2(\SB2_2_9/i0_4 ), .A3(
        \SB2_2_9/i1[9] ), .ZN(n2126) );
  NAND3_X2 U3060 ( .A1(\SB4_29/i0_3 ), .A2(\SB4_29/i0[8] ), .A3(\SB4_29/i0[9] ), .ZN(\SB4_29/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U3057 ( .I(\SB3_31/buf_output[3] ), .ZN(\SB4_29/i0[8] ) );
  NAND3_X2 \SB3_23/Component_Function_5/N4  ( .A1(\SB3_23/i0[9] ), .A2(
        \SB3_23/i0[6] ), .A3(\SB3_23/i0_4 ), .ZN(
        \SB3_23/Component_Function_5/NAND4_in[3] ) );
  INV_X2 U2759 ( .I(\MC_ARK_ARC_1_3/buf_output[134] ), .ZN(\SB1_4_9/i1[9] ) );
  NAND3_X2 \SB2_3_6/Component_Function_2/N2  ( .A1(\SB2_3_6/i0_3 ), .A2(
        \SB2_3_6/i0[10] ), .A3(\SB2_3_6/i0[6] ), .ZN(
        \SB2_3_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_10/Component_Function_3/N4  ( .A1(n589), .A2(
        \SB2_2_10/i0[8] ), .A3(\SB2_2_10/i3[0] ), .ZN(
        \SB2_2_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U4155 ( .A1(\SB1_3_8/i0[10] ), .A2(\SB1_3_8/i1[9] ), .A3(
        \SB1_3_8/i1_7 ), .ZN(n1184) );
  NAND3_X2 U3958 ( .A1(\SB1_4_13/i0[10] ), .A2(\SB1_4_13/i1_5 ), .A3(
        \SB1_4_13/i1[9] ), .ZN(n5247) );
  INV_X2 \SB1_1_27/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[27] ), .ZN(
        \SB1_1_27/i0[8] ) );
  INV_X2 \SB1_4_11/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[125] ), .ZN(
        \SB1_4_11/i1_5 ) );
  INV_X2 \SB2_4_9/INV_3  ( .I(\SB1_4_11/buf_output[3] ), .ZN(\SB2_4_9/i0[8] )
         );
  NAND3_X2 U4908 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0[10] ), .A3(
        \SB2_2_14/i0_4 ), .ZN(\SB2_2_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U6172 ( .A1(\SB2_3_5/i0[9] ), .A2(\SB2_3_5/i0_4 ), .A3(
        \SB2_3_5/i0[6] ), .ZN(n2955) );
  NAND3_X2 U5569 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0_0 ), .A3(
        \SB1_0_2/i0[7] ), .ZN(\SB1_0_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 \SB2_1_22/Component_Function_3/N1  ( .A1(\SB2_1_22/i1[9] ), .A2(
        \SB2_1_22/i0_3 ), .A3(\SB2_1_22/i0[6] ), .ZN(
        \SB2_1_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB1_3_7/Component_Function_3/N1  ( .A1(\SB1_3_7/i1[9] ), .A2(
        \SB1_3_7/i0_3 ), .A3(\SB1_3_7/i0[6] ), .ZN(
        \SB1_3_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U5338 ( .A1(\SB1_2_15/i0[9] ), .A2(\SB1_2_15/i0[8] ), .A3(
        \RI1[2][101] ), .ZN(n2089) );
  BUF_X4 U1498 ( .I(\SB3_17/buf_output[5] ), .Z(\SB4_17/i0_3 ) );
  INV_X2 U3177 ( .I(\SB1_1_20/buf_output[5] ), .ZN(\SB2_1_20/i1_5 ) );
  NAND3_X2 U876 ( .A1(\SB1_4_31/i0_3 ), .A2(\SB1_4_31/i0_0 ), .A3(
        \SB1_4_31/i0_4 ), .ZN(\SB1_4_31/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB4_23/BUF_4  ( .I(\SB3_24/buf_output[4] ), .Z(\SB4_23/i0_4 ) );
  INV_X2 U5448 ( .I(\MC_ARK_ARC_1_1/buf_output[13] ), .ZN(\SB1_2_29/i1_7 ) );
  NAND3_X2 \SB1_3_12/Component_Function_5/N2  ( .A1(\SB1_3_12/i0_0 ), .A2(
        \SB1_3_12/i0[6] ), .A3(\SB1_3_12/i0[10] ), .ZN(
        \SB1_3_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U1195 ( .A1(\SB2_0_31/i0[10] ), .A2(\SB2_0_31/i1[9] ), .A3(
        \SB2_0_31/i1_7 ), .ZN(\SB2_0_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U7431 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0_4 ), .A3(
        \SB2_2_16/i1[9] ), .ZN(n2389) );
  NAND2_X2 \SB3_29/Component_Function_5/N1  ( .A1(\SB3_29/i0_0 ), .A2(
        \SB3_29/i3[0] ), .ZN(\SB3_29/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U3175 ( .I(\SB1_1_20/buf_output[5] ), .Z(\SB2_1_20/i0_3 ) );
  NAND3_X2 \SB1_1_31/Component_Function_3/N2  ( .A1(\SB1_1_31/i0_0 ), .A2(
        \SB1_1_31/i0_3 ), .A3(\SB1_1_31/i0_4 ), .ZN(
        \SB1_1_31/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB1_4_10/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[130] ), .Z(
        \SB1_4_10/i0_4 ) );
  NAND3_X2 U8321 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i0[10] ), .A3(
        \SB2_3_16/i0_4 ), .ZN(n2869) );
  NAND3_X2 U1786 ( .A1(\SB1_1_31/i0_0 ), .A2(\SB1_1_31/i0_4 ), .A3(
        \SB1_1_31/i1_5 ), .ZN(n3723) );
  NAND3_X2 \SB2_0_15/Component_Function_4/N2  ( .A1(\SB2_0_15/i3[0] ), .A2(
        \SB1_0_18/buf_output[2] ), .A3(\SB2_0_15/i1_7 ), .ZN(
        \SB2_0_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U9416 ( .A1(\SB2_3_30/i1_7 ), .A2(\SB2_3_30/i0[8] ), .A3(
        \SB2_3_30/i0_4 ), .ZN(\SB2_3_30/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U2443 ( .A1(\SB4_13/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_13/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_13/Component_Function_2/NAND4_in[0] ), .A4(n3754), .ZN(n1260) );
  NAND3_X2 U6698 ( .A1(\SB1_4_4/i0_3 ), .A2(\SB1_4_4/i0_4 ), .A3(
        \SB1_4_4/i1[9] ), .ZN(n2056) );
  NAND3_X2 U696 ( .A1(\SB2_4_4/i0_3 ), .A2(\SB2_4_4/i0[10] ), .A3(
        \SB2_4_4/i0_4 ), .ZN(n3828) );
  NAND2_X2 \SB2_0_17/Component_Function_5/N1  ( .A1(\SB2_0_17/i0_0 ), .A2(
        \SB2_0_17/i3[0] ), .ZN(\SB2_0_17/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U1492 ( .I(\MC_ARK_ARC_1_4/buf_output[93] ), .ZN(\SB3_16/i0[8] ) );
  NAND3_X2 \SB2_2_4/Component_Function_2/N1  ( .A1(\SB2_2_4/i1_5 ), .A2(
        \SB2_2_4/i0[10] ), .A3(\SB2_2_4/i1[9] ), .ZN(
        \SB2_2_4/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 \SB2_3_5/Component_Function_3/N5  ( .A1(
        \SB2_3_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_5/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_3_5/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_3_5/buf_output[3] ) );
  INV_X2 U2482 ( .I(\SB3_16/buf_output[2] ), .ZN(\SB4_13/i1[9] ) );
  NAND4_X1 \SB2_0_28/Component_Function_1/N5  ( .A1(
        \SB2_0_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_28/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_28/buf_output[1] ) );
  BUF_X4 \SB2_2_24/BUF_0  ( .I(\SB1_2_29/buf_output[0] ), .Z(\SB2_2_24/i0[9] )
         );
  NAND3_X2 U1666 ( .A1(\SB2_1_22/i0[9] ), .A2(\SB2_1_22/i0[10] ), .A3(
        \SB2_1_22/i0_3 ), .ZN(n1417) );
  NAND3_X2 U4818 ( .A1(\SB2_4_20/i0_3 ), .A2(\SB2_4_20/i0[8] ), .A3(
        \SB2_4_20/i0[9] ), .ZN(\SB2_4_20/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 U734 ( .A1(\SB2_4_16/i0_0 ), .A2(\SB2_4_16/i3[0] ), .ZN(n3602) );
  NAND3_X2 U1729 ( .A1(\SB1_1_8/i0_0 ), .A2(\SB1_1_8/i0_4 ), .A3(
        \SB1_1_8/i1_5 ), .ZN(n5284) );
  BUF_X2 U2628 ( .I(\SB3_3/buf_output[0] ), .Z(\SB4_30/i0[9] ) );
  NAND3_X2 U891 ( .A1(\SB1_4_0/i0_3 ), .A2(\SB1_4_0/i0[8] ), .A3(
        \SB1_4_0/i0[9] ), .ZN(n1765) );
  NAND4_X2 \SB2_4_24/Component_Function_1/N5  ( .A1(
        \SB2_4_24/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_24/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_4_24/buf_output[1] ) );
  NAND3_X2 U6343 ( .A1(\SB1_4_25/i0_3 ), .A2(\SB1_4_25/i0[10] ), .A3(
        \SB1_4_25/i0[9] ), .ZN(\SB1_4_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U6245 ( .A1(n592), .A2(\SB2_3_12/i1_7 ), .A3(\SB2_3_12/i0[8] ), 
        .ZN(n1845) );
  NAND3_X2 U4106 ( .A1(\SB4_28/i0[6] ), .A2(\SB4_28/i1_5 ), .A3(\SB4_28/i0[9] ), .ZN(n2379) );
  INV_X2 U2932 ( .I(\SB3_28/buf_output[5] ), .ZN(\SB4_28/i1_5 ) );
  NAND2_X2 \SB2_1_31/Component_Function_5/N1  ( .A1(\SB2_1_31/i0_0 ), .A2(
        \SB2_1_31/i3[0] ), .ZN(\SB2_1_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_9/Component_Function_2/N1  ( .A1(\SB2_3_9/i1_5 ), .A2(
        \SB2_3_9/i0[10] ), .A3(\SB2_3_9/i1[9] ), .ZN(
        \SB2_3_9/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U10789 ( .A1(\SB2_2_21/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_21/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_2_21/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_2_21/buf_output[1] ) );
  NAND3_X2 \SB1_3_12/Component_Function_2/N2  ( .A1(\SB1_3_12/i0_3 ), .A2(
        \SB1_3_12/i0[10] ), .A3(\SB1_3_12/i0[6] ), .ZN(
        \SB1_3_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_3/Component_Function_2/N2  ( .A1(\SB2_1_3/i0_3 ), .A2(
        \SB2_1_3/i0[10] ), .A3(\SB2_1_3/i0[6] ), .ZN(
        \SB2_1_3/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U3244 ( .I(\SB1_1_5/buf_output[2] ), .Z(\SB2_1_2/i0_0 ) );
  NAND3_X2 \SB2_3_28/Component_Function_3/N3  ( .A1(\SB2_3_28/i1[9] ), .A2(
        \SB2_3_28/i1_7 ), .A3(\SB2_3_28/i0[10] ), .ZN(
        \SB2_3_28/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U1626 ( .I(\MC_ARK_ARC_1_1/buf_output[146] ), .Z(\SB1_2_7/i0_0 ) );
  INV_X2 U3124 ( .I(\SB1_4_18/buf_output[5] ), .ZN(\SB2_4_18/i1_5 ) );
  NAND3_X2 \SB2_2_10/Component_Function_4/N2  ( .A1(\SB2_2_10/i3[0] ), .A2(
        \SB2_2_10/i0_0 ), .A3(\SB2_2_10/i1_7 ), .ZN(
        \SB2_2_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U1112 ( .A1(\SB1_1_3/i0[6] ), .A2(\SB1_1_3/i0[10] ), .A3(
        \SB1_1_3/i0_0 ), .ZN(\SB1_1_3/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U5361 ( .I(\SB2_3_3/buf_output[2] ), .Z(n1506) );
  NAND3_X2 U1259 ( .A1(\SB1_3_6/i0[10] ), .A2(\SB1_3_6/i1[9] ), .A3(
        \SB1_3_6/i1_5 ), .ZN(n4449) );
  NAND2_X2 U5168 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i1[9] ), .ZN(n3352) );
  NAND3_X2 U1548 ( .A1(\SB1_2_27/i0[10] ), .A2(\SB1_2_27/i1[9] ), .A3(
        \SB1_2_27/i1_5 ), .ZN(n4103) );
  INV_X2 U4024 ( .I(\MC_ARK_ARC_1_4/buf_output[3] ), .ZN(\SB3_31/i0[8] ) );
  BUF_X4 \SB1_4_15/BUF_5  ( .I(\MC_ARK_ARC_1_3/buf_output[101] ), .Z(
        \SB1_4_15/i0_3 ) );
  INV_X2 \SB2_1_20/INV_1  ( .I(\SB1_1_24/buf_output[1] ), .ZN(\SB2_1_20/i1_7 )
         );
  NAND3_X2 \SB2_4_24/Component_Function_2/N2  ( .A1(\SB2_4_24/i0_3 ), .A2(
        \SB2_4_24/i0[10] ), .A3(\SB2_4_24/i0[6] ), .ZN(
        \SB2_4_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U2631 ( .A1(\SB4_6/i1_5 ), .A2(\SB4_6/i0_0 ), .A3(\SB4_6/i0_4 ), 
        .ZN(\SB4_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U858 ( .A1(\SB1_4_3/i0[8] ), .A2(\SB1_4_3/i1_5 ), .A3(
        \SB1_4_3/i3[0] ), .ZN(n1117) );
  BUF_X4 \SB2_3_10/BUF_3  ( .I(\SB1_3_12/buf_output[3] ), .Z(\SB2_3_10/i0[10] ) );
  BUF_X4 U9189 ( .I(\SB2_4_30/buf_output[1] ), .Z(\RI5[4][31] ) );
  BUF_X4 U1310 ( .I(\MC_ARK_ARC_1_2/buf_output[80] ), .Z(\SB1_3_18/i0_0 ) );
  NAND3_X2 U9434 ( .A1(\SB2_4_18/i0[10] ), .A2(\SB2_4_18/i1_7 ), .A3(
        \SB2_4_18/i1[9] ), .ZN(n4373) );
  NAND3_X2 U1256 ( .A1(\SB1_3_13/i0_0 ), .A2(\SB1_3_13/i1_5 ), .A3(
        \SB1_3_13/i0_4 ), .ZN(n4808) );
  NAND2_X2 \SB1_1_31/Component_Function_5/N1  ( .A1(\SB1_1_31/i0_0 ), .A2(
        \SB1_1_31/i3[0] ), .ZN(\SB1_1_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U1136 ( .A1(\SB2_3_31/i0_4 ), .A2(\SB2_3_31/i0[9] ), .A3(
        \SB2_3_31/i0[6] ), .ZN(n5352) );
  INV_X2 \SB1_4_26/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[35] ), .ZN(
        \SB1_4_26/i1_5 ) );
  INV_X2 U3129 ( .I(\RI3[0][87] ), .ZN(\SB2_0_17/i0[8] ) );
  BUF_X4 U3491 ( .I(\MC_ARK_ARC_1_1/buf_output[57] ), .Z(\SB1_2_22/i0[10] ) );
  NAND3_X2 U3950 ( .A1(\SB1_4_6/i0[10] ), .A2(\SB1_4_6/i1[9] ), .A3(
        \SB1_4_6/i1_7 ), .ZN(n2911) );
  BUF_X2 U2973 ( .I(\SB3_29/buf_output[3] ), .Z(\SB4_27/i0[10] ) );
  NAND3_X2 U1045 ( .A1(\SB2_1_0/i0[8] ), .A2(\SB2_1_0/i3[0] ), .A3(
        \SB2_1_0/i1_5 ), .ZN(\SB2_1_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U1137 ( .A1(\SB2_3_14/i0_3 ), .A2(\SB2_3_14/i1[9] ), .A3(
        \SB2_3_14/i0_4 ), .ZN(\SB2_3_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_9/Component_Function_2/N2  ( .A1(\SB2_3_9/i0_3 ), .A2(
        \SB2_3_9/i0[10] ), .A3(\SB2_3_9/i0[6] ), .ZN(
        \SB2_3_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U3765 ( .A1(\SB2_2_23/i0_3 ), .A2(n600), .A3(\SB2_2_23/i1[9] ), 
        .ZN(\SB2_2_23/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U1951 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i0[9] ), .A3(
        \SB2_0_28/i0[8] ), .ZN(\SB2_0_28/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB1_3_17/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[88] ), .Z(
        \SB1_3_17/i0_4 ) );
  NAND3_X2 U3969 ( .A1(\SB2_4_7/i0[9] ), .A2(\RI3[4][148] ), .A3(
        \SB2_4_7/i0[6] ), .ZN(n988) );
  NAND2_X2 \SB1_1_5/Component_Function_5/N1  ( .A1(\SB1_1_5/i0_0 ), .A2(
        \SB1_1_5/i3[0] ), .ZN(\SB1_1_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_4_10/Component_Function_1/N3  ( .A1(\SB1_4_10/i1_5 ), .A2(
        \SB1_4_10/i0[6] ), .A3(\SB1_4_10/i0[9] ), .ZN(
        \SB1_4_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB1_4_0/Component_Function_2/N1  ( .A1(\SB1_4_0/i1_5 ), .A2(
        \SB1_4_0/i0[10] ), .A3(\SB1_4_0/i1[9] ), .ZN(
        \SB1_4_0/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U5291 ( .I(\RI1[5][167] ), .Z(\SB3_4/i0_3 ) );
  BUF_X4 \SB2_2_30/BUF_0  ( .I(\SB1_2_3/buf_output[0] ), .Z(\SB2_2_30/i0[9] )
         );
  NAND3_X2 \SB1_3_20/Component_Function_0/N2  ( .A1(\SB1_3_20/i0[8] ), .A2(
        \SB1_3_20/i0[7] ), .A3(\SB1_3_20/i0[6] ), .ZN(
        \SB1_3_20/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U9621 ( .A1(\SB2_2_11/i0[10] ), .A2(\SB2_2_11/i1_5 ), .A3(
        \SB2_2_11/i1[9] ), .ZN(\SB2_2_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U1390 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0_0 ), .A3(
        \SB2_2_12/i0[7] ), .ZN(n3933) );
  NAND3_X2 U4846 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i0[6] ), .A3(
        \SB1_2_13/i1[9] ), .ZN(\SB1_2_13/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_0  ( .I(\SB2_3_4/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[0] ) );
  NAND3_X2 U1526 ( .A1(\SB1_2_12/i1[9] ), .A2(\RI1[2][119] ), .A3(
        \SB1_2_12/i0_4 ), .ZN(\SB1_2_12/Component_Function_5/NAND4_in[2] ) );
  BUF_X2 \SB1_4_10/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[126] ), .Z(
        \SB1_4_10/i0[9] ) );
  NAND4_X2 U6903 ( .A1(\SB2_3_13/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_13/buf_output[0] ) );
  NAND3_X2 \SB2_1_12/Component_Function_2/N1  ( .A1(\SB2_1_12/i1_5 ), .A2(
        \SB2_1_12/i0[10] ), .A3(\SB2_1_12/i1[9] ), .ZN(
        \SB2_1_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U2357 ( .A1(\SB2_4_8/i0_3 ), .A2(\SB2_4_8/i0[8] ), .A3(
        \SB2_4_8/i0[9] ), .ZN(\SB2_4_8/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U3786 ( .I(\MC_ARK_ARC_1_2/buf_output[112] ), .Z(\SB1_3_13/i0_4 ) );
  BUF_X4 \SB2_0_11/BUF_3  ( .I(\RI3[0][123] ), .Z(\SB2_0_11/i0[10] ) );
  CLKBUF_X4 \SB2_1_22/BUF_2  ( .I(\SB1_1_25/buf_output[2] ), .Z(
        \SB2_1_22/i0_0 ) );
  NAND3_X2 \SB2_3_15/Component_Function_2/N1  ( .A1(\SB2_3_15/i1_5 ), .A2(
        \SB2_3_15/i0[10] ), .A3(\SB2_3_15/i1[9] ), .ZN(
        \SB2_3_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U1681 ( .A1(\SB2_1_0/i0[6] ), .A2(\SB2_1_0/i0[10] ), .A3(
        \SB2_1_0/i0_3 ), .ZN(n4270) );
  NAND3_X2 U9646 ( .A1(\SB1_0_1/i0_0 ), .A2(\SB1_0_1/i0_3 ), .A3(
        \SB1_0_1/i0_4 ), .ZN(\SB1_0_1/Component_Function_3/NAND4_in[1] ) );
  NAND4_X1 U6601 ( .A1(\SB2_2_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_11/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_11/Component_Function_1/NAND4_in[1] ), .A4(n2014), .ZN(
        \SB2_2_11/buf_output[1] ) );
  NAND2_X2 \SB1_3_12/Component_Function_5/N1  ( .A1(\SB1_3_12/i0_0 ), .A2(
        \SB1_3_12/i3[0] ), .ZN(\SB1_3_12/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_4_18/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[80] ), .ZN(
        \SB1_4_18/i1[9] ) );
  INV_X2 \SB1_1_26/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[33] ), .ZN(
        \SB1_1_26/i0[8] ) );
  NAND3_X2 U3273 ( .A1(\SB1_3_30/i1[9] ), .A2(\SB1_3_30/i0_4 ), .A3(
        \SB1_3_30/i0_3 ), .ZN(\SB1_3_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U1566 ( .A1(\SB1_2_2/i0_0 ), .A2(\SB1_2_2/i1_5 ), .A3(
        \SB1_2_2/i0_4 ), .ZN(\SB1_2_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U7459 ( .A1(\SB2_3_10/i0[10] ), .A2(\SB2_3_10/i1[9] ), .A3(
        \SB2_3_10/i1_7 ), .ZN(n2405) );
  NAND3_X2 \SB2_4_7/Component_Function_4/N2  ( .A1(\SB2_4_7/i3[0] ), .A2(
        \SB2_4_7/i0_0 ), .A3(\SB2_4_7/i1_7 ), .ZN(
        \SB2_4_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U1297 ( .A1(n3757), .A2(\SB1_3_29/i0[8] ), .A3(\SB1_3_29/i0[9] ), 
        .ZN(\SB1_3_29/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB1_3_30/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[9] ), .ZN(
        \SB1_3_30/i0[8] ) );
  NAND3_X2 U2581 ( .A1(\SB1_4_28/i0_3 ), .A2(\SB1_4_28/i0_4 ), .A3(
        \SB1_4_28/i0_0 ), .ZN(n3254) );
  NAND3_X2 U4086 ( .A1(\SB2_3_27/i0[10] ), .A2(\SB2_3_27/i1[9] ), .A3(
        \SB2_3_27/i1_7 ), .ZN(n1154) );
  NAND3_X2 U2531 ( .A1(\SB1_2_25/i0_0 ), .A2(\SB1_2_25/i0_4 ), .A3(
        \SB1_2_25/i1_5 ), .ZN(n606) );
  NAND3_X2 U1216 ( .A1(\SB2_0_19/i1_5 ), .A2(\SB2_0_19/i1[9] ), .A3(
        \RI3[0][76] ), .ZN(\SB2_0_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_26/Component_Function_3/N3  ( .A1(\SB2_2_26/i1[9] ), .A2(
        \SB2_2_26/i1_7 ), .A3(\SB2_2_26/i0[10] ), .ZN(
        \SB2_2_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_4/Component_Function_3/N2  ( .A1(\SB2_1_4/i0_0 ), .A2(
        \SB2_1_4/i0_3 ), .A3(\SB2_1_4/i0_4 ), .ZN(
        \SB2_1_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U576 ( .A1(\SB3_13/i0_3 ), .A2(\SB3_13/i1[9] ), .A3(\SB3_13/i0_4 ), 
        .ZN(\SB3_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U7611 ( .A1(\SB2_4_21/i0[10] ), .A2(\SB2_4_21/i1_5 ), .A3(
        \SB2_4_21/i1[9] ), .ZN(\SB2_4_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_4_1/Component_Function_3/N2  ( .A1(\SB2_4_1/i0_0 ), .A2(
        \SB2_4_1/i0_3 ), .A3(\SB2_4_1/i0_4 ), .ZN(
        \SB2_4_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U1060 ( .A1(\SB2_3_6/i0_3 ), .A2(\SB2_3_6/i0[10] ), .A3(
        \SB2_3_6/i0_4 ), .ZN(n4464) );
  NAND3_X2 \SB2_1_15/Component_Function_4/N1  ( .A1(\SB2_1_15/i0[9] ), .A2(
        \SB2_1_15/i0_0 ), .A3(\SB2_1_15/i0[8] ), .ZN(
        \SB2_1_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U2125 ( .A1(\SB2_0_19/i1[9] ), .A2(\SB2_0_19/i1_7 ), .A3(
        \RI3[0][75] ), .ZN(\SB2_0_19/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U3384 ( .I(\MC_ARK_ARC_1_4/buf_output[113] ), .Z(\RI1[5][113] ) );
  INV_X2 U2522 ( .I(\MC_ARK_ARC_1_2/buf_output[32] ), .ZN(\SB1_3_26/i1[9] ) );
  BUF_X4 \SB1_1_8/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[141] ), .Z(
        \SB1_1_8/i0[10] ) );
  BUF_X4 U9697 ( .I(\MC_ARK_ARC_1_1/buf_output[20] ), .Z(\SB1_2_28/i0_0 ) );
  BUF_X4 \SB2_1_24/BUF_2  ( .I(\SB1_1_27/buf_output[2] ), .Z(\SB2_1_24/i0_0 )
         );
  BUF_X4 \SB2_3_26/BUF_1_0  ( .I(\SB2_3_26/buf_output[1] ), .Z(\RI5[3][55] )
         );
  NAND4_X2 U972 ( .A1(\SB2_3_26/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_26/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_3_26/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_3_26/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_26/buf_output[1] ) );
  NAND3_X2 U580 ( .A1(\SB3_26/i1[9] ), .A2(\SB3_26/i1_7 ), .A3(\SB3_26/i0[10] ), .ZN(\SB3_26/Component_Function_3/NAND4_in[2] ) );
  INV_X2 \SB1_3_5/INV_5  ( .I(\RI1[3][161] ), .ZN(\SB1_3_5/i1_5 ) );
  INV_X2 \SB1_1_21/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[61] ), .ZN(
        \SB1_1_21/i1_7 ) );
  NAND3_X2 U2778 ( .A1(\SB3_26/i0_0 ), .A2(\SB3_26/i0[6] ), .A3(
        \SB3_26/i0[10] ), .ZN(\SB3_26/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U1486 ( .I(\SB1_2_1/buf_output[0] ), .Z(\SB2_2_28/i0[9] ) );
  INV_X2 \SB2_0_19/INV_1  ( .I(\SB1_0_23/buf_output[1] ), .ZN(\SB2_0_19/i1_7 )
         );
  NAND3_X2 U7919 ( .A1(\SB2_3_6/i0_3 ), .A2(\SB2_3_6/i0[10] ), .A3(
        \SB2_3_6/i0[9] ), .ZN(n2634) );
  NAND3_X2 U1573 ( .A1(\SB1_2_1/i0[8] ), .A2(\SB1_2_1/i3[0] ), .A3(
        \SB1_2_1/i1_5 ), .ZN(n4958) );
  INV_X2 U2907 ( .I(n389), .ZN(\SB1_0_23/i1_5 ) );
  NAND3_X2 U2594 ( .A1(\SB2_4_27/i0[10] ), .A2(\SB2_4_27/i1[9] ), .A3(
        \SB2_4_27/i1_5 ), .ZN(n4055) );
  NAND3_X2 \SB1_0_23/Component_Function_2/N3  ( .A1(\SB1_0_23/i0_3 ), .A2(
        \SB1_0_23/i0[8] ), .A3(\SB1_0_23/i0[9] ), .ZN(
        \SB1_0_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U2126 ( .A1(\SB2_0_20/i1_5 ), .A2(\SB2_0_20/i0[10] ), .A3(
        \SB2_0_20/i1[9] ), .ZN(\SB2_0_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U3425 ( .A1(\SB2_1_0/i0[7] ), .A2(\SB2_1_0/i0[8] ), .A3(
        \SB2_1_0/i0[6] ), .ZN(n917) );
  NAND3_X2 U2005 ( .A1(\SB2_0_12/i0[10] ), .A2(\SB2_0_12/i0_0 ), .A3(
        \SB2_0_12/i0[6] ), .ZN(\SB2_0_12/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB1_0_8/INV_3  ( .I(n363), .ZN(\SB1_0_8/i0[8] ) );
  NAND2_X2 \SB2_4_1/Component_Function_5/N1  ( .A1(\SB2_4_1/i0_0 ), .A2(
        \SB2_4_1/i3[0] ), .ZN(\SB2_4_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_23/Component_Function_3/N3  ( .A1(\SB2_0_23/i1[9] ), .A2(
        \SB2_0_23/i1_7 ), .A3(\SB2_0_23/i0[10] ), .ZN(
        \SB2_0_23/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB2_0_28/BUF_4_0  ( .I(\SB2_0_28/buf_output[4] ), .Z(\RI5[0][28] )
         );
  BUF_X4 U3317 ( .I(n392), .Z(\SB1_0_20/i0_3 ) );
  INV_X2 \SB1_2_26/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[31] ), .ZN(
        \SB1_2_26/i1_7 ) );
  NAND4_X2 U9119 ( .A1(\SB2_3_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_22/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_22/buf_output[3] ) );
  NAND3_X2 U6837 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i1[9] ), .A3(
        \SB2_0_25/i0[6] ), .ZN(\SB2_0_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB1_3_5/Component_Function_2/N3  ( .A1(\SB1_3_5/i0_3 ), .A2(
        \SB1_3_5/i0[8] ), .A3(\SB1_3_5/i0[9] ), .ZN(
        \SB1_3_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_2/Component_Function_2/N2  ( .A1(\SB1_1_2/i0_3 ), .A2(
        \SB1_1_2/i0[10] ), .A3(\SB1_1_2/i0[6] ), .ZN(
        \SB1_1_2/Component_Function_2/NAND4_in[1] ) );
  INV_X2 \SB2_4_20/INV_5  ( .I(\SB1_4_20/buf_output[5] ), .ZN(\SB2_4_20/i1_5 )
         );
  NAND4_X2 \SB1_0_23/Component_Function_4/N5  ( .A1(
        \SB1_0_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_23/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_0_23/buf_output[4] ) );
  INV_X2 \SB2_0_22/INV_4  ( .I(\RI3[0][58] ), .ZN(\SB2_0_22/i0[7] ) );
  NAND3_X2 U1387 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i0_0 ), .A3(
        \SB2_2_27/i0_4 ), .ZN(\SB2_2_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_3_7/Component_Function_4/N3  ( .A1(\SB1_3_7/i0[9] ), .A2(
        \SB1_3_7/i0[10] ), .A3(\SB1_3_7/i0_3 ), .ZN(
        \SB1_3_7/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U4990 ( .A1(\SB2_4_4/i1_5 ), .A2(\SB2_4_4/i0[10] ), .A3(
        \SB2_4_4/i1[9] ), .ZN(\SB2_4_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U1360 ( .A1(\SB1_3_8/i0[10] ), .A2(\SB1_3_8/i0_0 ), .A3(
        \SB1_3_8/i0[6] ), .ZN(\SB1_3_8/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_14/Component_Function_3/N1  ( .A1(\SB2_2_14/i1[9] ), .A2(
        \SB2_2_14/i0_3 ), .A3(\SB2_2_14/i0[6] ), .ZN(
        \SB2_2_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U3262 ( .A1(\SB1_3_29/i0[6] ), .A2(\SB1_3_29/i0_0 ), .A3(
        \SB1_3_29/i0[10] ), .ZN(n857) );
  BUF_X4 U9746 ( .I(\SB1_3_29/buf_output[5] ), .Z(\SB2_3_29/i0_3 ) );
  NAND3_X2 \SB2_0_25/Component_Function_4/N4  ( .A1(\SB2_0_25/i1[9] ), .A2(
        \SB2_0_25/i1_5 ), .A3(\SB2_0_25/i0_4 ), .ZN(
        \SB2_0_25/Component_Function_4/NAND4_in[3] ) );
  BUF_X2 U2625 ( .I(\SB3_18/buf_output[2] ), .Z(\SB4_15/i0_0 ) );
  NAND2_X2 \SB1_3_29/Component_Function_5/N1  ( .A1(\SB1_3_29/i0_0 ), .A2(
        \SB1_3_29/i3[0] ), .ZN(\SB1_3_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_17/Component_Function_4/N4  ( .A1(\SB2_3_17/i1[9] ), .A2(
        \SB2_3_17/i1_5 ), .A3(\SB2_3_17/i0_4 ), .ZN(
        \SB2_3_17/Component_Function_4/NAND4_in[3] ) );
  INV_X2 U8111 ( .I(\SB1_4_15/buf_output[5] ), .ZN(\SB2_4_15/i1_5 ) );
  BUF_X4 \SB2_0_22/BUF_5  ( .I(\SB1_0_22/buf_output[5] ), .Z(\SB2_0_22/i0_3 )
         );
  BUF_X4 U2906 ( .I(n389), .Z(\SB1_0_23/i0_3 ) );
  BUF_X4 \SB2_1_23/BUF_4  ( .I(\SB1_1_24/buf_output[4] ), .Z(\SB2_1_23/i0_4 )
         );
  BUF_X4 \SB2_2_26/BUF_5  ( .I(\SB1_2_26/buf_output[5] ), .Z(\SB2_2_26/i0_3 )
         );
  OR3_X2 U2921 ( .A1(\RI1[3][5] ), .A2(\MC_ARK_ARC_1_2/buf_output[3] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[0] ), .Z(
        \SB1_3_31/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 U2698 ( .I(\SB2_4_3/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[183] ) );
  CLKBUF_X2 U166 ( .I(Key[165]), .Z(n109) );
  NAND4_X2 U2548 ( .A1(\SB3_14/Component_Function_5/NAND4_in[1] ), .A2(n1628), 
        .A3(\SB3_14/Component_Function_5/NAND4_in[0] ), .A4(
        \SB3_14/Component_Function_5/NAND4_in[2] ), .ZN(\SB3_14/buf_output[5] ) );
  NAND3_X2 \SB2_2_26/Component_Function_1/N3  ( .A1(\SB2_2_26/i1_5 ), .A2(
        \SB2_2_26/i0[6] ), .A3(\SB2_2_26/i0[9] ), .ZN(
        \SB2_2_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U704 ( .A1(n3370), .A2(\SB2_4_1/i0[6] ), .A3(\SB2_4_1/i0[8] ), .ZN(
        n4302) );
  NAND3_X2 U3290 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i0_4 ), .A3(
        \SB1_2_13/i1[9] ), .ZN(\SB1_2_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U6939 ( .A1(\SB2_2_13/i0[10] ), .A2(\SB2_2_13/i0_3 ), .A3(
        \SB2_2_13/i0[6] ), .ZN(\SB2_2_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U1011 ( .A1(\SB1_2_2/i0[8] ), .A2(\SB1_2_2/i3[0] ), .A3(
        \SB1_2_2/i1_5 ), .ZN(n1622) );
  NAND3_X2 \SB2_0_16/Component_Function_3/N3  ( .A1(\SB2_0_16/i1[9] ), .A2(
        \SB2_0_16/i1_7 ), .A3(\RI3[0][93] ), .ZN(
        \SB2_0_16/Component_Function_3/NAND4_in[2] ) );
  NAND2_X2 \SB2_0_3/Component_Function_0/N1  ( .A1(\SB2_0_3/i0[10] ), .A2(
        \SB2_0_3/i0[9] ), .ZN(\SB2_0_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 U2747 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0[8] ), .A3(
        \SB1_3_23/i0[9] ), .ZN(\SB1_3_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_14/Component_Function_2/N1  ( .A1(\SB2_3_14/i1_5 ), .A2(
        \SB2_3_14/i0[10] ), .A3(\SB2_3_14/i1[9] ), .ZN(
        \SB2_3_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_4_13/Component_Function_4/N1  ( .A1(\SB1_4_13/i0[9] ), .A2(
        \SB1_4_13/i0_0 ), .A3(\SB1_4_13/i0[8] ), .ZN(
        \SB1_4_13/Component_Function_4/NAND4_in[0] ) );
  INV_X4 \SB2_4_12/INV_4  ( .I(\SB2_4_12/i0_4 ), .ZN(\SB2_4_12/i0[7] ) );
  INV_X2 U2129 ( .I(n3579), .ZN(n1782) );
  NAND3_X2 \SB1_3_1/Component_Function_2/N2  ( .A1(\SB1_3_1/i0_3 ), .A2(
        \SB1_3_1/i0[10] ), .A3(\SB1_3_1/i0[6] ), .ZN(
        \SB1_3_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_7/Component_Function_1/N2  ( .A1(\SB2_2_7/i0_3 ), .A2(
        \SB2_2_7/i1_7 ), .A3(\SB2_2_7/i0[8] ), .ZN(
        \SB2_2_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U5001 ( .A1(\SB1_3_30/i0_0 ), .A2(\SB1_3_30/i0[6] ), .A3(
        \SB1_3_30/i0[10] ), .ZN(\SB1_3_30/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X2 U9626 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i0[6] ), .A3(
        \SB3_14/i0[10] ), .ZN(\SB3_14/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U3018 ( .I(\MC_ARK_ARC_1_3/buf_output[45] ), .ZN(\SB1_4_24/i0[8] ) );
  NAND3_X2 U1452 ( .A1(\SB2_2_4/i1[9] ), .A2(\SB2_2_4/i0_4 ), .A3(
        \SB2_2_4/i1_5 ), .ZN(n5413) );
  NAND3_X2 U3645 ( .A1(\SB1_1_16/i0[10] ), .A2(\SB1_1_16/i0_3 ), .A3(
        \SB1_1_16/i0[9] ), .ZN(n4068) );
  INV_X2 \SB1_1_1/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[183] ), .ZN(
        \SB1_1_1/i0[8] ) );
  INV_X2 \SB1_4_22/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[55] ), .ZN(
        \SB1_4_22/i1_7 ) );
  NAND3_X2 U6429 ( .A1(\SB2_4_5/i3[0] ), .A2(\SB2_4_5/i1_5 ), .A3(
        \SB2_4_5/i0[8] ), .ZN(n1937) );
  NAND3_X2 U9949 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0_0 ), .A3(
        \SB2_3_0/i0[7] ), .ZN(n4064) );
  NAND2_X2 \SB1_2_14/Component_Function_5/N1  ( .A1(\SB1_2_14/i0_0 ), .A2(
        \SB1_2_14/i3[0] ), .ZN(\SB1_2_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB3_30/Component_Function_4/N1  ( .A1(\SB3_30/i0[9] ), .A2(
        \SB3_30/i0_0 ), .A3(\SB3_30/i0[8] ), .ZN(
        \SB3_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U8814 ( .A1(\SB2_2_18/i0_3 ), .A2(\SB2_2_18/i1[9] ), .A3(
        \SB2_2_18/i0_4 ), .ZN(\SB2_2_18/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U756 ( .I(\SB1_4_5/buf_output[5] ), .ZN(\SB2_4_5/i1_5 ) );
  NAND2_X2 \SB2_3_1/Component_Function_1/N1  ( .A1(\SB2_3_1/i0_3 ), .A2(
        \SB2_3_1/i1[9] ), .ZN(\SB2_3_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U9677 ( .A1(\SB2_4_11/i0_3 ), .A2(\SB2_4_11/i0[8] ), .A3(
        \SB2_4_11/i0[9] ), .ZN(\SB2_4_11/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U3218 ( .I(\SB1_3_4/buf_output[5] ), .Z(\SB2_3_4/i0_3 ) );
  NAND3_X2 \SB2_0_20/Component_Function_4/N1  ( .A1(\SB2_0_20/i0[9] ), .A2(
        \SB2_0_20/i0_0 ), .A3(\SB2_0_20/i0[8] ), .ZN(
        \SB2_0_20/Component_Function_4/NAND4_in[0] ) );
  BUF_X4 U2009 ( .I(\SB2_2_21/buf_output[1] ), .Z(\RI5[2][85] ) );
  NAND3_X2 \SB2_0_19/Component_Function_0/N2  ( .A1(\SB2_0_19/i0[8] ), .A2(
        \SB2_0_19/i0[7] ), .A3(\SB2_0_19/i0[6] ), .ZN(
        \SB2_0_19/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U1538 ( .A1(\SB1_2_27/i0[9] ), .A2(\SB1_2_27/i0[8] ), .A3(
        \SB1_2_27/i0_3 ), .ZN(n4306) );
  BUF_X4 \SB2_0_16/BUF_2  ( .I(\SB1_0_19/buf_output[2] ), .Z(\SB2_0_16/i0_0 )
         );
  CLKBUF_X2 U21 ( .I(Key[74]), .Z(n202) );
  INV_X2 U5436 ( .I(\SB1_1_3/buf_output[1] ), .ZN(\SB2_1_31/i1_7 ) );
  NAND3_X2 U1660 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i0_0 ), .A3(
        \SB2_1_28/i0[7] ), .ZN(n5190) );
  NAND3_X2 \SB3_30/Component_Function_1/N2  ( .A1(\SB3_30/i0_3 ), .A2(
        \SB3_30/i1_7 ), .A3(\SB3_30/i0[8] ), .ZN(
        \SB3_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U3621 ( .A1(\SB1_1_21/i0[10] ), .A2(\SB1_1_21/i1_7 ), .A3(
        \SB1_1_21/i1[9] ), .ZN(\SB1_1_21/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U8275 ( .A1(\SB2_0_14/i0[9] ), .A2(\SB2_0_14/i0_4 ), .A3(
        \SB2_0_14/i0[6] ), .ZN(\SB2_0_14/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \SB2_2_18/BUF_1  ( .I(\SB1_2_22/buf_output[1] ), .Z(\SB2_2_18/i0[6] )
         );
  INV_X2 U9544 ( .I(\SB1_2_17/buf_output[5] ), .ZN(\SB2_2_17/i1_5 ) );
  NAND2_X2 U3707 ( .A1(\SB1_2_17/i0_0 ), .A2(\SB1_2_17/i3[0] ), .ZN(
        \SB1_2_17/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U2142 ( .I(\SB1_0_19/i0_0 ), .ZN(n3435) );
  NAND3_X2 U1198 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i0[6] ), .A3(
        \SB1_3_2/i0_0 ), .ZN(\SB1_3_2/Component_Function_5/NAND4_in[1] ) );
  INV_X4 \SB2_0_14/INV_0  ( .I(\SB2_0_14/i0[9] ), .ZN(\SB2_0_14/i3[0] ) );
  NAND3_X2 \SB1_1_18/Component_Function_1/N4  ( .A1(\SB1_1_18/i1_7 ), .A2(
        \SB1_1_18/i0[8] ), .A3(\SB1_1_18/i0_4 ), .ZN(
        \SB1_1_18/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U11759 ( .A1(\SB2_0_14/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_14/Component_Function_2/NAND4_in[0] ), .A3(n4889), .A4(
        \SB2_0_14/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_14/buf_output[2] ) );
  NAND3_X2 U2375 ( .A1(\SB1_4_27/i0[9] ), .A2(\SB1_4_27/i0_3 ), .A3(
        \SB1_4_27/i0[8] ), .ZN(\SB1_4_27/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U1737 ( .I(n304), .Z(\SB1_0_6/i0_0 ) );
  INV_X2 U1736 ( .I(n304), .ZN(\SB1_0_6/i1[9] ) );
  NAND3_X2 U3690 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i0[9] ), .A3(
        \SB2_1_28/i0[8] ), .ZN(n942) );
  NAND3_X2 U1529 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i0[9] ), .A3(
        \SB1_0_20/i0[10] ), .ZN(n2482) );
  INV_X4 U2115 ( .I(\RI3[0][76] ), .ZN(\SB2_0_19/i0[7] ) );
  NAND3_X2 U1599 ( .A1(\SB1_2_22/i1_5 ), .A2(\SB1_2_22/i0_0 ), .A3(
        \SB1_2_22/i0_4 ), .ZN(n4582) );
  INV_X2 \SB2_1_13/INV_1  ( .I(\SB1_1_17/buf_output[1] ), .ZN(\SB2_1_13/i1_7 )
         );
  INV_X2 \SB1_3_16/INV_0  ( .I(n1500), .ZN(\SB1_3_16/i3[0] ) );
  NAND3_X2 \SB2_4_21/Component_Function_3/N1  ( .A1(\SB2_4_21/i1[9] ), .A2(
        \SB2_4_21/i0_3 ), .A3(\SB2_4_21/i0[6] ), .ZN(
        \SB2_4_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_26/Component_Function_5/N3  ( .A1(\SB2_2_26/i1[9] ), .A2(
        n6686), .A3(\SB2_2_26/i0_3 ), .ZN(
        \SB2_2_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U3047 ( .A1(\SB1_1_11/i0_0 ), .A2(\SB1_1_11/i0_3 ), .A3(
        \SB1_1_11/i0_4 ), .ZN(\SB1_1_11/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U2043 ( .I(\SB1_1_3/buf_output[1] ), .Z(\SB2_1_31/i0[6] ) );
  BUF_X4 U9451 ( .I(\SB1_3_11/buf_output[3] ), .Z(\SB2_3_9/i0[10] ) );
  INV_X8 U1836 ( .I(\RI1[1][47] ), .ZN(\SB1_1_24/i1_5 ) );
  NAND3_X2 U3799 ( .A1(\RI3[0][82] ), .A2(\SB2_0_18/i0[9] ), .A3(
        \SB2_0_18/i0[6] ), .ZN(\SB2_0_18/Component_Function_5/NAND4_in[3] ) );
  INV_X2 U3306 ( .I(\RI3[0][173] ), .ZN(\SB2_0_3/i1_5 ) );
  INV_X2 \SB2_3_16/INV_1  ( .I(\SB1_3_20/buf_output[1] ), .ZN(\SB2_3_16/i1_7 )
         );
  NAND3_X2 U2926 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i1[9] ), .A3(
        \SB2_0_28/i0_4 ), .ZN(n3411) );
  AND4_X2 U240 ( .A1(\SB3_19/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_19/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_19/Component_Function_3/NAND4_in[1] ), .A4(
        \SB3_19/Component_Function_3/NAND4_in[3] ), .Z(n1493) );
  NAND3_X2 U1457 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0[8] ), .A3(
        \SB2_2_24/i0[9] ), .ZN(\SB2_2_24/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 \SB2_3_18/Component_Function_5/N1  ( .A1(\SB2_3_18/i0_0 ), .A2(
        \SB2_3_18/i3[0] ), .ZN(\SB2_3_18/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB2_4_3/INV_1  ( .I(\SB1_4_7/buf_output[1] ), .ZN(\SB2_4_3/i1_7 ) );
  NAND3_X2 \SB2_3_9/Component_Function_3/N4  ( .A1(\SB2_3_9/i1_5 ), .A2(
        \SB2_3_9/i0[8] ), .A3(\SB2_3_9/i3[0] ), .ZN(
        \SB2_3_9/Component_Function_3/NAND4_in[3] ) );
  INV_X2 U1346 ( .I(\MC_ARK_ARC_1_3/buf_output[147] ), .ZN(\SB1_4_7/i0[8] ) );
  NAND2_X2 U4004 ( .A1(\SB2_4_4/i0_0 ), .A2(\SB2_4_4/i3[0] ), .ZN(
        \SB2_4_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_4_7/Component_Function_1/N4  ( .A1(\SB1_4_7/i1_7 ), .A2(
        \SB1_4_7/i0[8] ), .A3(\SB1_4_7/i0_4 ), .ZN(
        \SB1_4_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U721 ( .A1(\SB2_4_20/i0[10] ), .A2(\SB2_4_20/i0_0 ), .A3(
        \SB2_4_20/i0[6] ), .ZN(\SB2_4_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U955 ( .A1(\SB2_2_10/i0[10] ), .A2(\SB2_2_10/i0[9] ), .A3(
        \SB2_2_10/i0_3 ), .ZN(n2286) );
  NAND3_X2 U2691 ( .A1(\SB3_15/i0[10] ), .A2(\SB3_15/i1[9] ), .A3(
        \SB3_15/i1_5 ), .ZN(\SB3_15/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U670 ( .A1(\SB2_4_21/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_4_21/Component_Function_1/NAND4_in[1] ), .A3(n4663), .A4(
        \SB2_4_21/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_4_21/buf_output[1] ) );
  NAND2_X2 \SB1_0_1/Component_Function_5/N1  ( .A1(\SB1_0_1/i0_0 ), .A2(
        \SB1_0_1/i3[0] ), .ZN(\SB1_0_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_12/Component_Function_3/N4  ( .A1(\SB2_2_12/i1_5 ), .A2(
        \SB2_2_12/i0[8] ), .A3(\SB2_2_12/i3[0] ), .ZN(
        \SB2_2_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U946 ( .A1(\SB1_4_8/i0_3 ), .A2(\SB1_4_8/i0[6] ), .A3(
        \SB1_4_8/i1[9] ), .ZN(n5311) );
  NAND3_X2 U7583 ( .A1(\SB2_2_26/i1[9] ), .A2(n6686), .A3(\SB2_2_26/i1_5 ), 
        .ZN(n5291) );
  NAND3_X2 U3928 ( .A1(\SB1_4_17/i0_3 ), .A2(\SB1_4_17/i0[10] ), .A3(
        \SB1_4_17/i0[6] ), .ZN(\SB1_4_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U11716 ( .A1(\SB2_2_26/i0[8] ), .A2(\SB2_2_26/i3[0] ), .A3(
        \SB2_2_26/i1_5 ), .ZN(n4873) );
  INV_X2 U1722 ( .I(\RI1[4][140] ), .ZN(\SB1_4_8/i1[9] ) );
  BUF_X4 \SB2_0_18/BUF_2  ( .I(\SB1_0_21/buf_output[2] ), .Z(\SB2_0_18/i0_0 )
         );
  NAND3_X2 U622 ( .A1(\SB3_0/i0_0 ), .A2(\SB3_0/i0_4 ), .A3(\SB3_0/i1_5 ), 
        .ZN(n2676) );
  NAND3_X2 \SB2_0_7/Component_Function_3/N2  ( .A1(\SB2_0_7/i0_0 ), .A2(
        \SB2_0_7/i0_3 ), .A3(\RI3[0][148] ), .ZN(
        \SB2_0_7/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 U5823 ( .I(\SB2_2_15/buf_output[2] ), .Z(\RI5[2][116] ) );
  INV_X2 \SB2_0_7/INV_1  ( .I(\SB1_0_11/buf_output[1] ), .ZN(\SB2_0_7/i1_7 )
         );
  NAND2_X2 \SB1_2_1/Component_Function_5/N1  ( .A1(\SB1_2_1/i0_0 ), .A2(
        \SB1_2_1/i3[0] ), .ZN(\SB1_2_1/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_0_11/INV_5  ( .I(n401), .ZN(\SB1_0_11/i1_5 ) );
  NAND3_X2 U596 ( .A1(\SB3_31/i0[6] ), .A2(\SB3_31/i0_0 ), .A3(\SB3_31/i0[10] ), .ZN(n3800) );
  BUF_X4 U1364 ( .I(\MC_ARK_ARC_1_2/buf_output[137] ), .Z(\SB1_3_9/i0_3 ) );
  NAND3_X2 U1281 ( .A1(\SB1_3_22/i0[9] ), .A2(\SB1_3_22/i0[8] ), .A3(
        \SB1_3_22/i0_3 ), .ZN(n4334) );
  BUF_X4 \SB2_4_24/BUF_1_0  ( .I(\SB2_4_24/buf_output[1] ), .Z(\RI5[4][67] )
         );
  BUF_X2 \SB2_4_0/BUF_1  ( .I(\SB1_4_4/buf_output[1] ), .Z(\SB2_4_0/i0[6] ) );
  BUF_X4 U1987 ( .I(\SB2_3_13/buf_output[0] ), .Z(\RI5[3][138] ) );
  INV_X2 U3198 ( .I(\SB1_4_27/buf_output[5] ), .ZN(\SB2_4_27/i1_5 ) );
  NAND2_X2 \SB2_2_13/Component_Function_0/N1  ( .A1(\SB2_2_13/i0[10] ), .A2(
        \SB2_2_13/i0[9] ), .ZN(\SB2_2_13/Component_Function_0/NAND4_in[0] ) );
  BUF_X4 U1920 ( .I(\SB1_2_31/buf_output[5] ), .Z(\SB2_2_31/i0_3 ) );
  NAND2_X2 \SB1_2_31/Component_Function_5/N1  ( .A1(\SB1_2_31/i0_0 ), .A2(
        \SB1_2_31/i3[0] ), .ZN(\SB1_2_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_27/Component_Function_3/N2  ( .A1(\SB2_0_27/i0_0 ), .A2(
        \SB2_0_27/i0_3 ), .A3(\RI3[0][28] ), .ZN(
        \SB2_0_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_4_11/Component_Function_3/N4  ( .A1(\SB2_4_11/i1_5 ), .A2(
        \SB2_4_11/i0[8] ), .A3(\SB2_4_11/i3[0] ), .ZN(
        \SB2_4_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U1396 ( .A1(\SB2_2_9/i0_0 ), .A2(\SB2_2_9/i0_3 ), .A3(
        \SB2_2_9/i0_4 ), .ZN(\SB2_2_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U7198 ( .A1(\SB1_1_22/i0[6] ), .A2(\SB1_1_22/i0[10] ), .A3(
        \SB1_1_22/i0_3 ), .ZN(n3631) );
  NAND3_X2 U849 ( .A1(\SB1_3_22/i0[8] ), .A2(\SB1_3_22/i0_4 ), .A3(
        \SB1_3_22/i1_7 ), .ZN(n2713) );
  NAND3_X2 \SB1_1_21/Component_Function_1/N3  ( .A1(\SB1_1_21/i1_5 ), .A2(
        \SB1_1_21/i0[6] ), .A3(\SB1_1_21/i0[9] ), .ZN(
        \SB1_1_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U3987 ( .A1(\SB2_4_5/i0_3 ), .A2(\SB2_4_5/i0[10] ), .A3(
        \SB2_4_5/i0[6] ), .ZN(\SB2_4_5/Component_Function_2/NAND4_in[1] ) );
  INV_X2 \SB1_0_22/INV_3  ( .I(n335), .ZN(\SB1_0_22/i0[8] ) );
  INV_X2 U2934 ( .I(\MC_ARK_ARC_1_0/buf_output[74] ), .ZN(\SB1_1_19/i1[9] ) );
  BUF_X4 \SB2_1_19/BUF_2  ( .I(\SB1_1_22/buf_output[2] ), .Z(\SB2_1_19/i0_0 )
         );
  NAND4_X1 U969 ( .A1(n4517), .A2(n2995), .A3(n4476), .A4(
        \SB2_3_23/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_23/buf_output[3] ) );
  NAND2_X2 \SB1_3_23/Component_Function_5/N1  ( .A1(\SB1_3_23/i0_0 ), .A2(
        \SB1_3_23/i3[0] ), .ZN(\SB1_3_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U718 ( .A1(\RI1[4][26] ), .A2(\SB1_4_27/i0[10] ), .A3(
        \SB1_4_27/i0[6] ), .ZN(\SB1_4_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U3092 ( .A1(\SB2_1_19/i0[10] ), .A2(\SB2_1_19/i0_3 ), .A3(
        \SB2_1_19/i0[6] ), .ZN(\SB2_1_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U5965 ( .A1(\SB2_2_6/i0_3 ), .A2(\SB2_2_6/i0_4 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(\SB2_2_6/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U1942 ( .I(\SB3_0/buf_output[5] ), .Z(\SB4_0/i0_3 ) );
  INV_X2 U53 ( .I(n158), .ZN(n220) );
  BUF_X4 \SB2_1_0/BUF_3  ( .I(\SB1_1_2/buf_output[3] ), .Z(\SB2_1_0/i0[10] )
         );
  NAND4_X2 U7274 ( .A1(\SB2_4_15/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_4_15/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_4_15/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_4_15/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_4_15/buf_output[1] ) );
  INV_X2 U9455 ( .I(\MC_ARK_ARC_1_4/buf_output[71] ), .ZN(\SB3_20/i1_5 ) );
  NAND3_X2 U1680 ( .A1(\SB2_1_19/i0[10] ), .A2(\SB2_1_19/i0_3 ), .A3(
        \SB2_1_19/i0[9] ), .ZN(n4200) );
  NAND3_X2 U4075 ( .A1(\SB3_27/i0[10] ), .A2(\SB3_27/i0_3 ), .A3(
        \SB3_27/i0[9] ), .ZN(n5419) );
  NAND3_X2 U1296 ( .A1(\SB1_3_12/i0[9] ), .A2(\SB1_3_12/i0[8] ), .A3(
        \SB1_3_12/i0_0 ), .ZN(n4599) );
  NAND3_X2 U1700 ( .A1(\SB1_2_15/i1_5 ), .A2(\SB1_2_15/i1[9] ), .A3(
        \SB1_2_15/i0_4 ), .ZN(n1821) );
  NAND3_X2 \SB2_2_14/Component_Function_1/N4  ( .A1(\SB2_2_14/i1_7 ), .A2(
        \SB2_2_14/i0[8] ), .A3(\SB2_2_14/i0_4 ), .ZN(
        \SB2_2_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 \SB2_3_9/Component_Function_3/N2  ( .A1(\SB2_3_9/i0_0 ), .A2(
        \SB2_3_9/i0_3 ), .A3(\SB1_3_10/buf_output[4] ), .ZN(
        \SB2_3_9/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB4_15/BUF_0  ( .I(\SB3_20/buf_output[0] ), .Z(\SB4_15/i0[9] ) );
  NAND2_X2 \SB1_0_23/Component_Function_5/N1  ( .A1(\SB1_0_23/i0_0 ), .A2(
        \SB1_0_23/i3[0] ), .ZN(\SB1_0_23/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U952 ( .I(\MC_ARK_ARC_1_3/buf_output[38] ), .Z(\SB1_4_25/i0_0 ) );
  NAND3_X2 \SB2_0_10/Component_Function_3/N2  ( .A1(\RI3[0][128] ), .A2(
        \SB2_0_10/i0_3 ), .A3(\SB2_0_10/i0_4 ), .ZN(
        \SB2_0_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_8/Component_Function_2/N2  ( .A1(\SB1_0_8/i0_3 ), .A2(
        \SB1_0_8/i0[10] ), .A3(\SB1_0_8/i0[6] ), .ZN(
        \SB1_0_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U9647 ( .A1(\SB1_0_1/i1_7 ), .A2(\SB1_0_1/i0[8] ), .A3(
        \SB1_0_1/i0_4 ), .ZN(\SB1_0_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U12308 ( .A1(\SB1_0_7/i0_0 ), .A2(\SB1_0_7/i0_3 ), .A3(
        \SB1_0_7/i0_4 ), .ZN(\SB1_0_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_8/Component_Function_2/N3  ( .A1(\SB1_0_8/i0_3 ), .A2(
        \SB1_0_8/i0[8] ), .A3(\SB1_0_8/i0[9] ), .ZN(
        \SB1_0_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB1_0_19/Component_Function_2/N3  ( .A1(\SB1_0_19/i0_3 ), .A2(
        \SB1_0_19/i0[8] ), .A3(\SB1_0_19/i0[9] ), .ZN(
        \SB1_0_19/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U3513 ( .A1(\SB2_1_2/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_1_2/Component_Function_1/NAND4_in[1] ), .A3(n1694), .A4(
        \SB2_1_2/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_2/buf_output[1] ) );
  NAND3_X2 \SB2_3_31/Component_Function_3/N3  ( .A1(\SB2_3_31/i1[9] ), .A2(
        \SB2_3_31/i1_7 ), .A3(\SB2_3_31/i0[10] ), .ZN(
        \SB2_3_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U7273 ( .A1(\SB1_2_4/i0_0 ), .A2(\SB1_2_4/i0_4 ), .A3(
        \SB1_2_4/i1_5 ), .ZN(\SB1_2_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U1629 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i0_0 ), .A3(
        \SB2_1_5/i0_4 ), .ZN(\SB2_1_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U1473 ( .A1(\SB2_2_6/i0[10] ), .A2(\SB2_2_6/i1_5 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(\SB2_2_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U1699 ( .A1(\RI1[2][101] ), .A2(\SB1_2_15/i1[9] ), .A3(
        \SB1_2_15/i0_4 ), .ZN(n2833) );
  BUF_X4 \SB1_1_23/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[50] ), .Z(
        \SB1_1_23/i0_0 ) );
  BUF_X4 \SB1_3_12/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[116] ), .Z(
        \SB1_3_12/i0_0 ) );
  BUF_X4 U3076 ( .I(\SB2_0_19/buf_output[2] ), .Z(\RI5[0][92] ) );
  NAND3_X2 U6865 ( .A1(\SB1_3_13/i0[10] ), .A2(\SB1_3_13/i0[6] ), .A3(
        \SB1_3_13/i0_0 ), .ZN(\SB1_3_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U709 ( .A1(\SB2_4_18/i0_3 ), .A2(\SB2_4_18/i0[10] ), .A3(
        \SB2_4_18/i0[9] ), .ZN(n5259) );
  NAND3_X2 U2748 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0_0 ), .A3(
        \SB1_3_23/i0_4 ), .ZN(\SB1_3_23/Component_Function_3/NAND4_in[1] ) );
  NAND2_X2 \SB1_1_20/Component_Function_5/N1  ( .A1(\SB1_1_20/i0_0 ), .A2(
        \SB1_1_20/i3[0] ), .ZN(\SB1_1_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U7806 ( .A1(\SB2_3_15/i0_0 ), .A2(\SB2_3_15/i0_4 ), .A3(
        \SB2_3_15/i1_5 ), .ZN(n2578) );
  BUF_X4 U3149 ( .I(\MC_ARK_ARC_1_2/buf_output[50] ), .Z(\SB1_3_23/i0_0 ) );
  NAND3_X2 \SB1_2_29/Component_Function_5/N2  ( .A1(\SB1_2_29/i0_0 ), .A2(
        \SB1_2_29/i0[6] ), .A3(\SB1_2_29/i0[10] ), .ZN(
        \SB1_2_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U2324 ( .A1(\SB2_3_9/i1_7 ), .A2(\SB2_3_9/i0[8] ), .A3(
        \SB1_3_10/buf_output[4] ), .ZN(
        \SB2_3_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U8613 ( .A1(\SB2_1_3/i0_3 ), .A2(\SB2_1_3/i0[10] ), .A3(
        \SB2_1_3/i0[9] ), .ZN(n3858) );
  NAND3_X2 \SB1_3_30/Component_Function_0/N2  ( .A1(\SB1_3_30/i0[8] ), .A2(
        \SB1_3_30/i0[7] ), .A3(\SB1_3_30/i0[6] ), .ZN(
        \SB1_3_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X2 U2462 ( .A1(\SB4_18/i0[10] ), .A2(\SB4_18/i0[9] ), .ZN(
        \SB4_18/Component_Function_0/NAND4_in[0] ) );
  BUF_X4 U3304 ( .I(\SB1_2_11/buf_output[5] ), .Z(\SB2_2_11/i0_3 ) );
  BUF_X4 U3127 ( .I(\SB1_4_18/buf_output[5] ), .Z(\SB2_4_18/i0_3 ) );
  BUF_X4 U9420 ( .I(\SB1_4_29/buf_output[4] ), .Z(\SB2_4_28/i0_4 ) );
  CLKBUF_X4 U3106 ( .I(\RI3[0][170] ), .Z(\SB2_0_3/i0_0 ) );
  BUF_X4 U3844 ( .I(\SB1_3_15/buf_output[4] ), .Z(\SB2_3_14/i0_4 ) );
  BUF_X4 U5184 ( .I(\SB1_4_19/buf_output[2] ), .Z(\SB2_4_16/i0_0 ) );
  CLKBUF_X2 U197 ( .I(Key[140]), .Z(n140) );
  NAND3_X2 U6334 ( .A1(\SB2_0_22/i0[7] ), .A2(\SB2_0_22/i0[8] ), .A3(
        \RI3[0][55] ), .ZN(n3534) );
  NAND3_X2 U2136 ( .A1(\SB1_0_24/i0[10] ), .A2(\SB1_0_24/i1[9] ), .A3(
        \SB1_0_24/i1_7 ), .ZN(\SB1_0_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB1_4_7/Component_Function_4/N3  ( .A1(\SB1_4_7/i0[9] ), .A2(
        \SB1_4_7/i0[10] ), .A3(\SB1_4_7/i0_3 ), .ZN(
        \SB1_4_7/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 \SB2_0_9/BUF_4_0  ( .I(\SB2_0_9/buf_output[4] ), .Z(\RI5[0][142] ) );
  NAND4_X2 U6806 ( .A1(\SB2_0_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_9/Component_Function_4/NAND4_in[3] ), .A4(n3590), .ZN(
        \SB2_0_9/buf_output[4] ) );
  BUF_X4 \SB1_2_4/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[162] ), .Z(
        \SB1_2_4/i0[9] ) );
  BUF_X2 U1130 ( .I(\SB1_3_1/buf_output[0] ), .Z(\SB2_3_28/i0[9] ) );
  INV_X2 U3216 ( .I(\SB1_3_4/buf_output[5] ), .ZN(\SB2_3_4/i1_5 ) );
  NAND3_X2 U10253 ( .A1(\SB3_7/i1_5 ), .A2(\SB3_7/i1[9] ), .A3(\SB3_7/i0_4 ), 
        .ZN(n4190) );
  NAND3_X2 U1670 ( .A1(\SB2_1_12/i0[10] ), .A2(\SB2_1_12/i0_3 ), .A3(
        \SB2_1_12/i0_4 ), .ZN(n3646) );
  NAND3_X2 \SB2_2_6/Component_Function_1/N3  ( .A1(\SB2_2_6/i1_5 ), .A2(
        \SB2_2_6/i0[6] ), .A3(\SB2_2_6/i0[9] ), .ZN(
        \SB2_2_6/Component_Function_1/NAND4_in[2] ) );
  INV_X4 \SB1_0_20/INV_4  ( .I(\SB1_0_20/i0_4 ), .ZN(\SB1_0_20/i0[7] ) );
  NAND3_X2 \SB2_3_7/Component_Function_3/N3  ( .A1(\SB2_3_7/i1[9] ), .A2(
        \SB2_3_7/i1_7 ), .A3(\SB2_3_7/i0[10] ), .ZN(
        \SB2_3_7/Component_Function_3/NAND4_in[2] ) );
  INV_X2 \SB1_2_25/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[39] ), .ZN(
        \SB1_2_25/i0[8] ) );
  BUF_X4 \SB3_1/BUF_4  ( .I(\MC_ARK_ARC_1_4/buf_output[184] ), .Z(\SB3_1/i0_4 ) );
  NAND3_X2 U1598 ( .A1(\SB1_2_7/i1_5 ), .A2(\SB1_2_7/i0_4 ), .A3(
        \SB1_2_7/i0_0 ), .ZN(\SB1_2_7/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 \SB1_0_2/Component_Function_1/N1  ( .A1(\SB1_0_2/i0_3 ), .A2(
        \SB1_0_2/i1[9] ), .ZN(\SB1_0_2/Component_Function_1/NAND4_in[0] ) );
  BUF_X2 \SB2_4_7/BUF_0  ( .I(\SB1_4_12/buf_output[0] ), .Z(\SB2_4_7/i0[9] )
         );
  INV_X2 U2796 ( .I(\MC_ARK_ARC_1_4/buf_output[74] ), .ZN(\SB3_19/i1[9] ) );
  BUF_X4 U3286 ( .I(\MC_ARK_ARC_1_3/buf_output[83] ), .Z(\SB1_4_18/i0_3 ) );
  NAND3_X2 \SB2_2_27/Component_Function_2/N4  ( .A1(\SB2_2_27/i1_5 ), .A2(
        \SB2_2_27/i0_0 ), .A3(\SB2_2_27/i0_4 ), .ZN(
        \SB2_2_27/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 U3809 ( .A1(\SB1_3_8/i0_0 ), .A2(\SB1_3_8/i3[0] ), .ZN(n4392) );
  NAND3_X1 \SB2_1_29/Component_Function_4/N3  ( .A1(\SB2_1_29/i0[9] ), .A2(
        \SB2_1_29/i0[10] ), .A3(\SB2_1_29/i0_3 ), .ZN(
        \SB2_1_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U1397 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i1_5 ), .A3(
        \SB2_2_27/i1[9] ), .ZN(n3377) );
  NAND3_X2 U808 ( .A1(\SB2_3_15/i0[10] ), .A2(\SB2_3_15/i1_7 ), .A3(
        \SB2_3_15/i1[9] ), .ZN(n714) );
  BUF_X4 U2795 ( .I(\MC_ARK_ARC_1_4/buf_output[74] ), .Z(\SB3_19/i0_0 ) );
  NAND3_X2 U4318 ( .A1(\SB1_1_23/i0_0 ), .A2(\SB1_1_23/i3[0] ), .A3(
        \SB1_1_23/i1_7 ), .ZN(\SB1_1_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_6/Component_Function_3/N3  ( .A1(\SB2_0_6/i1[9] ), .A2(
        \SB2_0_6/i1_7 ), .A3(\SB2_0_6/i0[10] ), .ZN(
        \SB2_0_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U3983 ( .A1(\SB1_0_8/i0_4 ), .A2(\SB1_0_8/i0_0 ), .A3(
        \SB1_0_8/i0_3 ), .ZN(\SB1_0_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U646 ( .A1(\SB3_17/i0_3 ), .A2(\SB3_17/i0[10] ), .A3(\SB3_17/i0[9] ), .ZN(n5358) );
  NAND3_X2 \SB2_1_5/Component_Function_3/N1  ( .A1(\SB2_1_5/i1[9] ), .A2(
        \SB2_1_5/i0_3 ), .A3(\SB2_1_5/i0[6] ), .ZN(
        \SB2_1_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U8197 ( .A1(\SB1_1_5/i0[6] ), .A2(\SB1_1_5/i0[10] ), .A3(
        \SB1_1_5/i0_0 ), .ZN(\SB1_1_5/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U5747 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i0_0 ), .A3(
        \SB1_3_5/i0_4 ), .ZN(\SB1_3_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_3_21/Component_Function_5/N3  ( .A1(\SB2_3_21/i1[9] ), .A2(
        \RI3[3][64] ), .A3(\SB2_3_21/i0_3 ), .ZN(
        \SB2_3_21/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_21/Component_Function_3/N1  ( .A1(\SB2_2_21/i1[9] ), .A2(
        \SB2_2_21/i0_3 ), .A3(\SB2_2_21/i0[6] ), .ZN(
        \SB2_2_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB1_3_16/Component_Function_0/N3  ( .A1(\SB1_3_16/i0[10] ), .A2(
        \SB1_3_16/i0_4 ), .A3(\SB1_3_16/i0_3 ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_183  ( .I(\SB2_3_3/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[183] ) );
  NAND3_X2 \SB2_3_16/Component_Function_4/N4  ( .A1(\SB2_3_16/i1[9] ), .A2(
        n571), .A3(\SB2_3_16/i0_4 ), .ZN(
        \SB2_3_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U3222 ( .A1(\SB1_3_22/i0_3 ), .A2(\SB1_3_22/i0_0 ), .A3(
        \SB1_3_22/i0_4 ), .ZN(n2310) );
  NAND3_X2 \SB2_2_19/Component_Function_1/N4  ( .A1(\SB2_2_19/i1_7 ), .A2(
        \SB2_2_19/i0[8] ), .A3(\SB2_2_19/i0_4 ), .ZN(
        \SB2_2_19/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 \SB1_2_31/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[3] ), .Z(
        \SB1_2_31/i0[10] ) );
  BUF_X2 U11455 ( .I(\SB1_2_31/buf_output[5] ), .Z(n4734) );
  AOI21_X2 U2615 ( .A1(\SB1_4_19/i3[0] ), .A2(\SB1_4_19/i0_0 ), .B(n3397), 
        .ZN(n3396) );
  BUF_X2 U9305 ( .I(Key[58]), .Z(n199) );
  NAND3_X2 \SB2_3_21/Component_Function_3/N1  ( .A1(\SB2_3_21/i1[9] ), .A2(
        \SB2_3_21/i0_3 ), .A3(\SB2_3_21/i0[6] ), .ZN(
        \SB2_3_21/Component_Function_3/NAND4_in[0] ) );
  CLKBUF_X4 \SB2_0_31/BUF_2  ( .I(\SB1_0_2/buf_output[2] ), .Z(\SB2_0_31/i0_0 ) );
  INV_X2 \SB2_0_21/INV_1  ( .I(n5959), .ZN(\SB2_0_21/i1_7 ) );
  BUF_X4 U5319 ( .I(\RI1[2][125] ), .Z(\SB1_2_11/i0_3 ) );
  BUF_X4 U3677 ( .I(\SB1_1_24/buf_output[0] ), .Z(\SB2_1_19/i0[9] ) );
  NAND2_X2 \SB1_4_18/Component_Function_5/N1  ( .A1(\SB1_4_18/i0_0 ), .A2(
        \SB1_4_18/i3[0] ), .ZN(\SB1_4_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U3832 ( .A1(\SB1_3_25/i1_7 ), .A2(\SB1_3_25/i0[8] ), .A3(
        \SB1_3_25/i0_4 ), .ZN(\SB1_3_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U6114 ( .A1(\SB3_17/i0[10] ), .A2(\SB3_17/i1[9] ), .A3(
        \SB3_17/i1_5 ), .ZN(n1787) );
  NAND3_X2 \SB2_4_18/Component_Function_3/N2  ( .A1(\SB2_4_18/i0_0 ), .A2(
        \SB2_4_18/i0_3 ), .A3(\SB2_4_18/i0_4 ), .ZN(
        \SB2_4_18/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 U3340 ( .I(\MC_ARK_ARC_1_2/buf_output[85] ), .Z(\SB1_3_17/i0[6] ) );
  BUF_X4 \SB2_0_0/BUF_3_0  ( .I(\SB2_0_0/buf_output[3] ), .Z(\RI5[0][9] ) );
  NAND3_X2 U943 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0[10] ), .A3(
        \SB2_2_12/i0[9] ), .ZN(\SB2_2_12/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 U3159 ( .I(\SB1_2_21/buf_output[5] ), .Z(\SB2_2_21/i0_3 ) );
  NAND3_X2 U698 ( .A1(\SB2_4_18/i0_3 ), .A2(\SB2_4_18/i0[10] ), .A3(
        \SB2_4_18/i0[6] ), .ZN(n5315) );
  NAND4_X2 U22 ( .A1(\SB4_5/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_5/Component_Function_1/NAND4_in[0] ), .ZN(n5201) );
  BUF_X4 \SB1_4_28/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[18] ), .Z(
        \SB1_4_28/i0[9] ) );
  BUF_X2 U703 ( .I(\SB1_4_28/buf_output[0] ), .Z(\SB2_4_23/i0[9] ) );
  INV_X2 U1366 ( .I(\MC_ARK_ARC_1_4/buf_output[147] ), .ZN(\SB3_7/i0[8] ) );
  NAND3_X2 U2630 ( .A1(\SB4_6/i1[9] ), .A2(\SB4_6/i1_5 ), .A3(\SB4_6/i0_4 ), 
        .ZN(\SB4_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U2378 ( .A1(n6268), .A2(\SB2_4_24/i0[8] ), .A3(\SB2_4_24/i3[0] ), 
        .ZN(\SB2_4_24/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_1_5/BUF_3  ( .I(\SB1_1_7/buf_output[3] ), .Z(\SB2_1_5/i0[10] )
         );
  NAND3_X2 \SB2_1_13/Component_Function_3/N4  ( .A1(\SB2_1_13/i1_5 ), .A2(
        \SB2_1_13/i0[8] ), .A3(\SB2_1_13/i3[0] ), .ZN(
        \SB2_1_13/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 U1171 ( .I(\MC_ARK_ARC_1_0/buf_output[96] ), .Z(\SB1_1_15/i0[9] ) );
  INV_X8 \SB1_2_12/INV_2  ( .I(\RI1[2][116] ), .ZN(\SB1_2_12/i1[9] ) );
  NAND3_X2 \SB2_1_11/Component_Function_3/N1  ( .A1(\SB2_1_11/i1[9] ), .A2(
        \SB2_1_11/i0_3 ), .A3(\SB2_1_11/i0[6] ), .ZN(
        \SB2_1_11/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_131_1  ( .I(\MC_ARK_ARC_1_3/buf_output[131] ), 
        .Z(\RI1[4][131] ) );
  NAND3_X2 U1947 ( .A1(\SB2_0_18/i0_3 ), .A2(\SB2_0_18/i0[6] ), .A3(
        \SB2_0_18/i1[9] ), .ZN(\SB2_0_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB1_4_27/Component_Function_2/N1  ( .A1(\SB1_4_27/i1_5 ), .A2(
        \SB1_4_27/i0[10] ), .A3(\SB1_4_27/i1[9] ), .ZN(
        \SB1_4_27/Component_Function_2/NAND4_in[0] ) );
  AND4_X2 U228 ( .A1(\SB3_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_24/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_24/Component_Function_2/NAND4_in[3] ), .Z(n3998) );
  NAND3_X2 U2241 ( .A1(\RI1[2][119] ), .A2(\SB1_2_12/i0[9] ), .A3(
        \SB1_2_12/i0[10] ), .ZN(n2915) );
  NAND2_X2 U814 ( .A1(\SB1_4_27/i3[0] ), .A2(\RI1[4][26] ), .ZN(n4587) );
  NAND3_X2 \SB2_1_12/Component_Function_2/N3  ( .A1(\SB2_1_12/i0_3 ), .A2(
        \SB2_1_12/i0[8] ), .A3(\SB2_1_12/i0[9] ), .ZN(
        \SB2_1_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U4394 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i0_4 ), .A3(
        \SB1_3_8/i1[9] ), .ZN(n1271) );
  NAND3_X2 \SB2_0_31/Component_Function_3/N2  ( .A1(\SB2_0_31/i0_0 ), .A2(
        \SB2_0_31/i0_3 ), .A3(\RI3[0][4] ), .ZN(
        \SB2_0_31/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U9778 ( .I(\SB1_3_13/buf_output[5] ), .ZN(\SB2_3_13/i1_5 ) );
  NAND3_X2 \SB2_0_15/Component_Function_2/N2  ( .A1(\SB2_0_15/i0_3 ), .A2(
        \SB2_0_15/i0[10] ), .A3(\SB2_0_15/i0[6] ), .ZN(
        \SB2_0_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_25/Component_Function_2/N3  ( .A1(\SB2_0_25/i0_3 ), .A2(
        \SB2_0_25/i0[8] ), .A3(\SB2_0_25/i0[9] ), .ZN(
        \SB2_0_25/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U2798 ( .I(\SB1_4_29/buf_output[3] ), .ZN(\SB2_4_27/i0[8] ) );
  INV_X2 \SB1_0_25/INV_5  ( .I(n387), .ZN(\SB1_0_25/i1_5 ) );
  NAND3_X2 U9800 ( .A1(\SB2_3_28/i0_0 ), .A2(\SB2_3_28/i1_5 ), .A3(
        \SB1_3_29/buf_output[4] ), .ZN(
        \SB2_3_28/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 \SB2_3_6/BUF_4  ( .I(\SB1_3_7/buf_output[4] ), .Z(\SB2_3_6/i0_4 ) );
  NAND3_X2 \SB2_0_22/Component_Function_1/N3  ( .A1(\SB2_0_22/i1_5 ), .A2(
        \RI3[0][55] ), .A3(\SB2_0_22/i0[9] ), .ZN(
        \SB2_0_22/Component_Function_1/NAND4_in[2] ) );
  AND4_X2 U214 ( .A1(\SB3_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_3/NAND4_in[2] ), .A4(n863), .Z(n3989) );
  NAND3_X2 U681 ( .A1(\SB2_4_22/i0[10] ), .A2(\SB2_4_22/i1_5 ), .A3(
        \SB2_4_22/i1[9] ), .ZN(\SB2_4_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U11793 ( .A1(\SB1_1_6/i0[10] ), .A2(\SB1_1_6/i0[9] ), .A3(
        \SB1_1_6/i0_3 ), .ZN(n4899) );
  BUF_X4 \SB1_3_15/BUF_5  ( .I(\RI1[3][101] ), .Z(\SB1_3_15/i0_3 ) );
  NAND3_X2 \SB2_2_28/Component_Function_0/N2  ( .A1(\SB2_2_28/i0[8] ), .A2(
        \SB2_2_28/i0[7] ), .A3(\SB2_2_28/i0[6] ), .ZN(
        \SB2_2_28/Component_Function_0/NAND4_in[1] ) );
  BUF_X4 \SB2_1_5/BUF_4  ( .I(\SB1_1_6/buf_output[4] ), .Z(\SB2_1_5/i0_4 ) );
  NAND3_X2 U942 ( .A1(\SB2_2_7/i0_0 ), .A2(\SB2_2_7/i0_3 ), .A3(
        \SB2_2_7/i0[7] ), .ZN(n976) );
  INV_X2 U1849 ( .I(\MC_ARK_ARC_1_1/buf_output[65] ), .ZN(\SB1_2_21/i1_5 ) );
  NAND3_X2 U4123 ( .A1(\SB4_6/i0[10] ), .A2(\SB4_6/i0_3 ), .A3(\SB4_6/i0_4 ), 
        .ZN(\SB4_6/Component_Function_0/NAND4_in[2] ) );
  INV_X2 U3017 ( .I(\MC_ARK_ARC_1_2/buf_output[44] ), .ZN(\SB1_3_24/i1[9] ) );
  NAND3_X2 \SB3_30/Component_Function_2/N4  ( .A1(\SB3_30/i1_5 ), .A2(
        \SB3_30/i0_0 ), .A3(\SB3_30/i0_4 ), .ZN(
        \SB3_30/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U2413 ( .A1(\SB3_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_24/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_24/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_24/buf_output[2] ) );
  NAND3_X2 U9725 ( .A1(\SB2_2_6/i1[9] ), .A2(\SB2_2_6/i0_3 ), .A3(
        \SB2_2_6/i0[6] ), .ZN(\SB2_2_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U3413 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0[8] ), .A3(
        \SB2_2_28/i1_7 ), .ZN(\SB2_2_28/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X4 \SB2_0_12/BUF_2  ( .I(\RI3[0][116] ), .Z(\SB2_0_12/i0_0 ) );
  NAND3_X2 U2414 ( .A1(\SB2_4_19/i1_5 ), .A2(\SB2_4_19/i0[6] ), .A3(
        \SB2_4_19/i0[9] ), .ZN(\SB2_4_19/Component_Function_1/NAND4_in[2] ) );
  NAND2_X2 \SB2_4_5/Component_Function_1/N1  ( .A1(\SB2_4_5/i0_3 ), .A2(
        \SB2_4_5/i1[9] ), .ZN(\SB2_4_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U12379 ( .A1(\SB1_4_5/i0_4 ), .A2(\SB1_4_5/i0[6] ), .A3(
        \SB1_4_5/i0[9] ), .ZN(n5238) );
  NAND2_X2 \SB1_1_28/Component_Function_5/N1  ( .A1(\SB1_1_28/i0_0 ), .A2(
        \SB1_1_28/i3[0] ), .ZN(\SB1_1_28/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB1_3_13/Component_Function_5/N1  ( .A1(\SB1_3_13/i0_0 ), .A2(
        \SB1_3_13/i3[0] ), .ZN(\SB1_3_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U9797 ( .A1(\SB1_0_2/i0[10] ), .A2(\SB1_0_2/i1[9] ), .A3(
        \SB1_0_2/i1_7 ), .ZN(n1920) );
  INV_X2 \SB3_22/INV_2  ( .I(\MC_ARK_ARC_1_4/buf_output[56] ), .ZN(
        \SB3_22/i1[9] ) );
  CLKBUF_X2 U226 ( .I(Key[113]), .Z(n176) );
  NAND3_X2 \SB2_4_22/Component_Function_3/N1  ( .A1(\SB2_4_22/i1[9] ), .A2(
        \SB2_4_22/i0_3 ), .A3(\SB2_4_22/i0[6] ), .ZN(
        \SB2_4_22/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U1850 ( .I(\MC_ARK_ARC_1_1/buf_output[65] ), .Z(\SB1_2_21/i0_3 ) );
  BUF_X4 U3775 ( .I(\MC_ARK_ARC_1_2/buf_output[141] ), .Z(\SB1_3_8/i0[10] ) );
  NAND3_X2 U9557 ( .A1(\SB2_2_27/i1[9] ), .A2(\SB2_2_27/i1_7 ), .A3(
        \SB2_2_27/i0[10] ), .ZN(\SB2_2_27/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X2 \SB2_2_17/Component_Function_2/N1  ( .A1(\SB2_2_17/i1_5 ), .A2(
        \SB2_2_17/i0[10] ), .A3(\SB2_2_17/i1[9] ), .ZN(
        \SB2_2_17/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB1_2_1/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[182] ), .Z(
        \SB1_2_1/i0_0 ) );
  NAND3_X2 U4251 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i1[9] ), .A3(
        \RI3[2][88] ), .ZN(\SB2_2_17/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U1768 ( .I(\SB1_3_5/buf_output[5] ), .ZN(\SB2_3_5/i1_5 ) );
  NAND3_X2 \SB2_3_18/Component_Function_3/N4  ( .A1(\SB2_3_18/i1_5 ), .A2(
        \SB2_3_18/i0[8] ), .A3(\SB2_3_18/i3[0] ), .ZN(
        \SB2_3_18/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB1_3_25/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[37] ), .Z(
        \SB1_3_25/i0[6] ) );
  NAND3_X2 \SB2_3_2/Component_Function_1/N3  ( .A1(\SB2_3_2/i1_5 ), .A2(
        \SB2_3_2/i0[6] ), .A3(\SB2_3_2/i0[9] ), .ZN(
        \SB2_3_2/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 \SB1_2_26/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[30] ), .Z(
        \SB1_2_26/i0[9] ) );
  INV_X4 \SB1_1_30/INV_4  ( .I(\SB1_1_30/i0_4 ), .ZN(\SB1_1_30/i0[7] ) );
  NAND3_X2 \SB1_3_28/Component_Function_2/N3  ( .A1(\SB1_3_28/i0_3 ), .A2(
        \SB1_3_28/i0[8] ), .A3(\SB1_3_28/i0[9] ), .ZN(
        \SB1_3_28/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB3_11/INV_5  ( .I(n3970), .ZN(\SB3_11/i1_5 ) );
  INV_X2 U5443 ( .I(n408), .ZN(\SB1_0_4/i1_5 ) );
  NAND3_X2 \SB2_2_15/Component_Function_1/N2  ( .A1(\SB2_2_15/i0_3 ), .A2(
        \SB2_2_15/i1_7 ), .A3(\SB2_2_15/i0[8] ), .ZN(
        \SB2_2_15/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \SB1_2_23/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[50] ), .Z(
        \SB1_2_23/i0_0 ) );
  NAND3_X2 \SB1_0_4/Component_Function_2/N3  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i0[8] ), .A3(\SB1_0_4/i0[9] ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB2_0_0/BUF_4_0  ( .I(\SB2_0_0/buf_output[4] ), .Z(\RI5[0][4] ) );
  INV_X2 U2219 ( .I(n6289), .ZN(\SB1_2_14/i1_5 ) );
  NAND3_X2 U1403 ( .A1(\SB2_2_28/i0[10] ), .A2(\SB2_2_28/i0_0 ), .A3(
        \SB2_2_28/i0[6] ), .ZN(\SB2_2_28/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U3675 ( .I(\SB1_1_10/buf_output[5] ), .ZN(\SB2_1_10/i1_5 ) );
  NAND3_X2 U7041 ( .A1(\SB2_3_13/i1_5 ), .A2(n6746), .A3(\SB2_3_13/i1[9] ), 
        .ZN(\SB2_3_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB2_1_23/Component_Function_3/N3  ( .A1(\SB2_1_23/i1[9] ), .A2(
        \SB2_1_23/i1_7 ), .A3(\SB2_1_23/i0[10] ), .ZN(
        \SB2_1_23/Component_Function_3/NAND4_in[2] ) );
  NAND2_X2 U2025 ( .A1(\SB1_0_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_2/Component_Function_3/NAND4_in[3] ), .ZN(n3362) );
  NAND3_X2 U3722 ( .A1(\SB1_2_17/i0[8] ), .A2(\SB1_2_17/i3[0] ), .A3(
        \SB1_2_17/i1_5 ), .ZN(\SB1_2_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB2_1_2/Component_Function_3/N3  ( .A1(\SB2_1_2/i1[9] ), .A2(
        \SB2_1_2/i1_7 ), .A3(\SB2_1_2/i0[10] ), .ZN(
        \SB2_1_2/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U3711 ( .I(\MC_ARK_ARC_1_1/buf_output[100] ), .Z(\SB1_2_15/i0_4 ) );
  INV_X2 U1448 ( .I(\SB3_8/buf_output[3] ), .ZN(\SB4_6/i0[8] ) );
  NAND3_X2 U2605 ( .A1(\SB2_4_29/i0_0 ), .A2(\SB2_4_29/i1_5 ), .A3(
        \SB2_4_29/i0_4 ), .ZN(n1337) );
  NAND3_X2 U1679 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0[9] ), .ZN(n4690) );
  INV_X2 U3104 ( .I(\MC_ARK_ARC_1_3/buf_output[135] ), .ZN(\SB1_4_9/i0[8] ) );
  INV_X2 U1328 ( .I(\MC_ARK_ARC_1_4/buf_output[140] ), .ZN(\SB3_8/i1[9] ) );
  NAND3_X2 U3942 ( .A1(\SB1_4_12/i1_5 ), .A2(\SB1_4_12/i1[9] ), .A3(
        \SB1_4_12/i0_4 ), .ZN(n757) );
  NAND3_X2 U1414 ( .A1(\SB2_2_1/i0_0 ), .A2(\SB2_2_1/i0[9] ), .A3(
        \SB2_2_1/i0[8] ), .ZN(n3672) );
  NAND3_X2 \SB2_1_28/Component_Function_0/N2  ( .A1(\SB2_1_28/i0[8] ), .A2(
        \SB2_1_28/i0[7] ), .A3(\SB2_1_28/i0[6] ), .ZN(
        \SB2_1_28/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 \SB4_6/Component_Function_1/N2  ( .A1(\SB4_6/i0_3 ), .A2(
        \SB4_6/i1_7 ), .A3(\SB4_6/i0[8] ), .ZN(
        \SB4_6/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U1214 ( .A1(\SB1_3_24/i0[6] ), .A2(\SB1_3_24/i0_4 ), .A3(
        \SB1_3_24/i0[9] ), .ZN(n3792) );
  NAND3_X2 U1757 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0[10] ), .A3(
        \SB2_2_30/i0[6] ), .ZN(\SB2_2_30/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U5785 ( .A1(\SB2_0_10/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_10/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_0_10/Component_Function_0/NAND4_in[0] ), .A4(n1651), .ZN(
        \SB2_0_10/buf_output[0] ) );
  BUF_X4 U3214 ( .I(\MC_ARK_ARC_1_3/buf_output[149] ), .Z(\SB1_4_7/i0_3 ) );
  BUF_X2 \SB2_0_10/BUF_0  ( .I(\RI3[0][126] ), .Z(\SB2_0_10/i0[9] ) );
  INV_X2 U2863 ( .I(\MC_ARK_ARC_1_4/buf_output[189] ), .ZN(\SB3_0/i0[8] ) );
  NAND3_X2 U5021 ( .A1(\SB3_19/i0_0 ), .A2(\SB3_19/i0[6] ), .A3(
        \SB3_19/i0[10] ), .ZN(\SB3_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U3010 ( .A1(\SB1_1_25/i0_0 ), .A2(\SB1_1_25/i1_5 ), .A3(
        \SB1_1_25/i0_4 ), .ZN(n766) );
  INV_X1 \SB2_0_15/INV_1  ( .I(\RI3[0][97] ), .ZN(\SB2_0_15/i1_7 ) );
  NAND2_X2 \SB4_6/Component_Function_0/N1  ( .A1(\SB4_6/i0[10] ), .A2(
        \SB4_6/i0[9] ), .ZN(\SB4_6/Component_Function_0/NAND4_in[0] ) );
  NAND4_X2 U3564 ( .A1(\SB4_26/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_26/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_26/Component_Function_1/NAND4_in[3] ), .ZN(n1120) );
  NAND3_X2 U1664 ( .A1(\SB2_1_11/i0_3 ), .A2(\SB2_1_11/i0_0 ), .A3(
        \SB2_1_11/i0[7] ), .ZN(n5344) );
  NAND3_X2 \SB1_3_14/Component_Function_5/N4  ( .A1(\SB1_3_14/i0[9] ), .A2(
        \SB1_3_14/i0[6] ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB2_1_13/Component_Function_4/N1  ( .A1(\SB2_1_13/i0[9] ), .A2(
        \SB2_1_13/i0_0 ), .A3(\SB2_1_13/i0[8] ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U1458 ( .A1(\SB2_4_0/i0_3 ), .A2(\SB2_4_0/i0[10] ), .A3(
        \SB2_4_0/i0[6] ), .ZN(\SB2_4_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U781 ( .A1(\SB1_4_23/i0_3 ), .A2(\SB1_4_23/i1[9] ), .A3(
        \SB1_4_23/i0_4 ), .ZN(\SB1_4_23/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_2_22/BUF_2  ( .I(\SB1_2_25/buf_output[2] ), .Z(\SB2_2_22/i0_0 )
         );
  INV_X2 \SB1_2_28/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[18] ), .ZN(
        \SB1_2_28/i3[0] ) );
  BUF_X4 U2380 ( .I(\MC_ARK_ARC_1_3/buf_output[16] ), .Z(\SB1_4_29/i0_4 ) );
  BUF_X4 U3701 ( .I(\SB2_1_19/buf_output[3] ), .Z(\RI5[1][87] ) );
  NAND3_X2 \SB2_0_16/Component_Function_2/N1  ( .A1(\SB2_0_16/i1_5 ), .A2(
        n6976), .A3(\SB2_0_16/i1[9] ), .ZN(
        \SB2_0_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_4_29/Component_Function_2/N1  ( .A1(\SB2_4_29/i1_5 ), .A2(
        \SB2_4_29/i0[10] ), .A3(\SB2_4_29/i1[9] ), .ZN(
        \SB2_4_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U1469 ( .A1(\SB2_4_29/i1[9] ), .A2(\SB2_4_29/i0_3 ), .A3(
        \SB2_4_29/i0[6] ), .ZN(\SB2_4_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U9680 ( .A1(\SB3_1/i1_5 ), .A2(\SB3_1/i0[8] ), .A3(\SB3_1/i3[0] ), 
        .ZN(n2062) );
  NAND3_X2 U1243 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i1[9] ), .A3(
        \SB1_0_16/i0_4 ), .ZN(\SB1_0_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_16/Component_Function_1/N3  ( .A1(\SB2_2_16/i1_5 ), .A2(
        \SB2_2_16/i0[6] ), .A3(\SB2_2_16/i0[9] ), .ZN(
        \SB2_2_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB3_12/Component_Function_2/N1  ( .A1(\SB3_12/i1_5 ), .A2(
        \SB3_12/i0[10] ), .A3(\SB3_12/i1[9] ), .ZN(
        \SB3_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_7/Component_Function_0/N3  ( .A1(\SB2_2_7/i0[10] ), .A2(
        \SB2_2_7/i0_4 ), .A3(\SB2_2_7/i0_3 ), .ZN(
        \SB2_2_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U10166 ( .A1(\SB2_0_27/i0_0 ), .A2(\SB2_0_27/i0[9] ), .A3(
        \SB2_0_27/i0[8] ), .ZN(\SB2_0_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U9396 ( .A1(\SB2_4_13/i1_5 ), .A2(\SB2_4_13/i0[10] ), .A3(
        \SB2_4_13/i1[9] ), .ZN(\SB2_4_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_4_31/Component_Function_1/N2  ( .A1(\SB1_4_31/i0_3 ), .A2(
        \SB1_4_31/i1_7 ), .A3(\SB1_4_31/i0[8] ), .ZN(
        \SB1_4_31/Component_Function_1/NAND4_in[1] ) );
  BUF_X2 \SB2_0_31/BUF_0  ( .I(\RI3[0][0] ), .Z(\SB2_0_31/i0[9] ) );
  BUF_X4 U5442 ( .I(n408), .Z(\SB1_0_4/i0_3 ) );
  INV_X2 U769 ( .I(\SB1_4_26/buf_output[5] ), .ZN(\SB2_4_26/i1_5 ) );
  NAND3_X2 U730 ( .A1(\SB2_4_14/i0_3 ), .A2(\SB2_4_14/i0[8] ), .A3(
        \SB2_4_14/i0[9] ), .ZN(\SB2_4_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U3814 ( .A1(\SB1_3_0/i0_3 ), .A2(\SB1_3_0/i0[9] ), .A3(
        \SB1_3_0/i0[8] ), .ZN(n5114) );
  NAND3_X2 U1161 ( .A1(\SB1_3_24/i0_3 ), .A2(\SB1_3_24/i0_0 ), .A3(
        \SB1_3_24/i0_4 ), .ZN(\SB1_3_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_4/Component_Function_3/N2  ( .A1(\SB1_0_4/i0_0 ), .A2(
        \SB1_0_4/i0_3 ), .A3(\SB1_0_4/i0_4 ), .ZN(
        \SB1_0_4/Component_Function_3/NAND4_in[1] ) );
  INV_X4 U3890 ( .I(\SB1_4_19/i0_4 ), .ZN(\SB1_4_19/i0[7] ) );
  BUF_X4 U3681 ( .I(\SB1_1_23/buf_output[3] ), .Z(\SB2_1_21/i0[10] ) );
  CLKBUF_X4 \SB2_0_2/BUF_3  ( .I(\RI3[0][177] ), .Z(\SB2_0_2/i0[10] ) );
  CLKBUF_X2 U92 ( .I(Key[179]), .Z(n216) );
  NAND3_X2 \SB2_1_0/Component_Function_5/N3  ( .A1(\SB2_1_0/i1[9] ), .A2(n590), 
        .A3(\SB2_1_0/i0_3 ), .ZN(\SB2_1_0/Component_Function_5/NAND4_in[2] )
         );
  NAND4_X1 U10086 ( .A1(\SB1_4_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_4_30/Component_Function_3/NAND4_in[3] ), .A4(n4125), .ZN(
        \SB1_4_30/buf_output[3] ) );
  NAND3_X2 U2745 ( .A1(\SB3_25/i0[10] ), .A2(\SB3_25/i1[9] ), .A3(
        \SB3_25/i1_5 ), .ZN(\SB3_25/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_3_25/BUF_4  ( .I(\SB1_3_26/buf_output[4] ), .Z(\SB2_3_25/i0_4 )
         );
  NAND2_X2 \SB2_2_24/Component_Function_5/N1  ( .A1(\SB2_2_24/i0_0 ), .A2(
        \SB2_2_24/i3[0] ), .ZN(\SB2_2_24/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U3046 ( .I(\MC_ARK_ARC_1_2/buf_output[33] ), .Z(\SB1_3_26/i0[10] ) );
  INV_X2 U3045 ( .I(\MC_ARK_ARC_1_2/buf_output[33] ), .ZN(\SB1_3_26/i0[8] ) );
  NAND2_X2 U9726 ( .A1(\SB2_2_6/i0_3 ), .A2(\SB2_2_6/i1[9] ), .ZN(
        \SB2_2_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U611 ( .A1(\SB3_25/i0[8] ), .A2(\SB3_25/i3[0] ), .A3(\SB3_25/i1_5 ), 
        .ZN(n2011) );
  NAND3_X2 U1306 ( .A1(\SB1_3_0/i0[6] ), .A2(\SB1_3_0/i0_3 ), .A3(
        \SB1_3_0/i0[10] ), .ZN(n5347) );
  INV_X2 U7107 ( .I(\SB1_3_23/buf_output[5] ), .ZN(\SB2_3_23/i1_5 ) );
  BUF_X2 \SB2_3_23/BUF_3_0  ( .I(\SB2_3_23/buf_output[3] ), .Z(\RI5[3][63] )
         );
  NAND3_X2 \SB1_4_22/Component_Function_2/N4  ( .A1(\SB1_4_22/i1_5 ), .A2(
        \SB1_4_22/i0_0 ), .A3(\SB1_4_22/i0_4 ), .ZN(
        \SB1_4_22/Component_Function_2/NAND4_in[3] ) );
  INV_X2 \SB3_25/INV_5  ( .I(\RI1[5][41] ), .ZN(\SB3_25/i1_5 ) );
  NAND3_X2 U6937 ( .A1(\SB1_3_6/i0[8] ), .A2(\SB1_3_6/i3[0] ), .A3(
        \SB1_3_6/i1_5 ), .ZN(n2163) );
  NAND3_X2 U10216 ( .A1(\SB2_0_16/i0_3 ), .A2(n594), .A3(n6976), .ZN(
        \SB2_0_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U1684 ( .A1(\SB2_1_3/i0_3 ), .A2(\SB2_1_3/i0[9] ), .A3(
        \SB2_1_3/i0[8] ), .ZN(\SB2_1_3/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 \SB3_23/Component_Function_5/N1  ( .A1(\SB3_23/i0_0 ), .A2(
        \SB3_23/i3[0] ), .ZN(\SB3_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U883 ( .A1(\SB1_3_22/i0[9] ), .A2(\SB1_3_22/i0[8] ), .A3(
        \SB1_3_22/i0_0 ), .ZN(\SB1_3_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U5966 ( .A1(\SB1_3_25/i0_3 ), .A2(\SB1_3_25/i0[8] ), .A3(
        \SB1_3_25/i1_7 ), .ZN(\SB1_3_25/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X4 U351 ( .I(\SB3_21/buf_output[4] ), .Z(\SB4_20/i0_4 ) );
  NAND3_X2 \SB1_0_13/Component_Function_3/N3  ( .A1(\SB1_0_13/i1[9] ), .A2(
        \SB1_0_13/i1_7 ), .A3(\SB1_0_13/i0[10] ), .ZN(
        \SB1_0_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_18/Component_Function_1/N4  ( .A1(\SB2_3_18/i1_7 ), .A2(
        \SB2_3_18/i0[8] ), .A3(\SB2_3_18/i0_4 ), .ZN(
        \SB2_3_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U11773 ( .A1(\SB1_3_20/i0[8] ), .A2(\SB1_3_20/i1_5 ), .A3(
        \SB1_3_20/i3[0] ), .ZN(\SB1_3_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_2_0/Component_Function_3/N4  ( .A1(\SB1_2_0/i1_5 ), .A2(
        \SB1_2_0/i0[8] ), .A3(\SB1_2_0/i3[0] ), .ZN(
        \SB1_2_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U1643 ( .A1(\SB2_1_0/i0_0 ), .A2(\SB2_1_0/i0_3 ), .A3(n590), .ZN(
        n4228) );
  NAND3_X2 U8711 ( .A1(\SB2_4_22/i0[9] ), .A2(\SB2_4_22/i0_3 ), .A3(
        \SB2_4_22/i0[8] ), .ZN(n3098) );
  BUF_X4 U1617 ( .I(\SB1_2_0/buf_output[2] ), .Z(\SB2_2_29/i0_0 ) );
  INV_X2 \SB1_4_24/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[47] ), .ZN(
        \SB1_4_24/i1_5 ) );
  NAND3_X2 \SB1_1_31/Component_Function_1/N3  ( .A1(\SB1_1_31/i1_5 ), .A2(
        \SB1_1_31/i0[6] ), .A3(\SB1_1_31/i0[9] ), .ZN(
        \SB1_1_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U6723 ( .A1(\SB2_1_0/i0_0 ), .A2(\SB2_1_0/i0_3 ), .A3(
        \SB2_1_0/i0[7] ), .ZN(\SB2_1_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 \SB1_3_28/Component_Function_0/N4  ( .A1(\SB1_3_28/i0[7] ), .A2(
        \SB1_3_28/i0_3 ), .A3(\SB1_3_28/i0_0 ), .ZN(
        \SB1_3_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U743 ( .A1(\SB1_4_20/i0[10] ), .A2(\SB1_4_20/i1[9] ), .A3(
        \SB1_4_20/i1_5 ), .ZN(n2034) );
  BUF_X4 \SB2_0_8/BUF_1_0  ( .I(\SB2_0_8/buf_output[1] ), .Z(\RI5[0][163] ) );
  NAND4_X2 U10927 ( .A1(\SB2_0_8/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_0_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_8/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_0_8/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_8/buf_output[1] ) );
  NAND2_X2 U1338 ( .A1(\SB1_3_14/i0_0 ), .A2(\SB1_3_14/i3[0] ), .ZN(n5180) );
  BUF_X4 \SB1_2_0/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[190] ), .Z(
        \SB1_2_0/i0_4 ) );
  INV_X2 \SB1_1_10/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[131] ), .ZN(
        \SB1_1_10/i1_5 ) );
  NAND3_X2 U1309 ( .A1(\SB1_3_29/i0_4 ), .A2(\SB1_3_29/i1[9] ), .A3(
        \SB1_3_29/i1_5 ), .ZN(n807) );
  INV_X8 \SB1_2_0/INV_5  ( .I(\RI1[2][191] ), .ZN(\SB1_2_0/i1_5 ) );
  BUF_X4 \SB1_4_6/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[150] ), .Z(
        \SB1_4_6/i0[9] ) );
  BUF_X4 U1999 ( .I(\SB1_3_5/buf_output[5] ), .Z(\SB2_3_5/i0_3 ) );
  BUF_X4 \SB2_4_3/BUF_2  ( .I(\SB1_4_6/buf_output[2] ), .Z(\SB2_4_3/i0_0 ) );
  BUF_X4 \SB2_1_10/BUF_4  ( .I(\SB1_1_11/buf_output[4] ), .Z(\SB2_1_10/i0_4 )
         );
  BUF_X4 \SB1_1_28/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[22] ), .Z(
        \SB1_1_28/i0_4 ) );
  CLKBUF_X2 U222 ( .I(Key[159]), .Z(n172) );
  INV_X2 \SB1_2_9/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[133] ), .ZN(
        \SB1_2_9/i1_7 ) );
  NAND3_X2 U2206 ( .A1(\SB2_1_15/i1[9] ), .A2(\SB2_1_15/i1_5 ), .A3(
        \SB2_1_15/i0_4 ), .ZN(\SB2_1_15/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \SB2_2_12/BUF_4  ( .I(\SB1_2_13/buf_output[4] ), .Z(\SB2_2_12/i0_4 )
         );
  NAND3_X2 \SB1_2_24/Component_Function_3/N1  ( .A1(\SB1_2_24/i1[9] ), .A2(
        \SB1_2_24/i0_3 ), .A3(\SB1_2_24/i0[6] ), .ZN(
        \SB1_2_24/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 U2646 ( .A1(\SB1_1_1/Component_Function_4/NAND4_in[0] ), .A2(n647), 
        .ZN(n646) );
  NAND3_X2 U6303 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i1[9] ), .A3(
        \SB2_3_24/i0_4 ), .ZN(n2364) );
  NAND3_X2 U2227 ( .A1(\SB1_2_20/i1_5 ), .A2(\SB1_2_20/i0_0 ), .A3(
        \SB1_2_20/i0_4 ), .ZN(\SB1_2_20/Component_Function_2/NAND4_in[3] ) );
  INV_X2 \SB1_4_9/INV_5  ( .I(n5424), .ZN(\SB1_4_9/i1_5 ) );
  NAND3_X2 \SB2_4_17/Component_Function_2/N1  ( .A1(\SB2_4_17/i1_5 ), .A2(
        \SB2_4_17/i0[10] ), .A3(\SB2_4_17/i1[9] ), .ZN(
        \SB2_4_17/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB1_4_0/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[189] ), .Z(
        \SB1_4_0/i0[10] ) );
  INV_X2 U2607 ( .I(\SB1_3_21/buf_output[5] ), .ZN(\SB2_3_21/i1_5 ) );
  BUF_X4 U9543 ( .I(\SB1_2_17/buf_output[5] ), .Z(\SB2_2_17/i0_3 ) );
  BUF_X4 \SB2_2_10/BUF_2  ( .I(\SB1_2_13/buf_output[2] ), .Z(\SB2_2_10/i0_0 )
         );
  CLKBUF_X4 \SB1_2_22/BUF_0  ( .I(n6938), .Z(\SB1_2_22/i0[9] ) );
  BUF_X4 \SB2_3_8/BUF_2  ( .I(\SB1_3_11/buf_output[2] ), .Z(\SB2_3_8/i0_0 ) );
  BUF_X4 \SB1_2_13/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[108] ), .Z(
        \SB1_2_13/i0[9] ) );
  NAND3_X1 \SB2_2_22/Component_Function_0/N2  ( .A1(\SB2_2_22/i0[8] ), .A2(
        \SB2_2_22/i0[7] ), .A3(\SB2_2_22/i0[6] ), .ZN(
        \SB2_2_22/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U10566 ( .A1(\SB2_4_30/i0_0 ), .A2(\SB1_4_31/buf_output[4] ), .A3(
        \SB2_4_30/i1_5 ), .ZN(n4321) );
  NAND3_X2 U9596 ( .A1(\SB2_3_30/i0_3 ), .A2(\SB2_3_30/i0[8] ), .A3(
        \SB2_3_30/i0[9] ), .ZN(\SB2_3_30/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB2_1_4/BUF_4  ( .I(\SB1_1_5/buf_output[4] ), .Z(\SB2_1_4/i0_4 ) );
  BUF_X4 U9600 ( .I(\SB1_0_0/buf_output[4] ), .Z(\RI3[0][4] ) );
  NAND3_X2 \SB2_3_24/Component_Function_4/N4  ( .A1(\SB2_3_24/i1[9] ), .A2(
        \SB2_3_24/i1_5 ), .A3(\SB2_3_24/i0_4 ), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[3] ) );
  NAND2_X2 \SB1_3_0/Component_Function_5/N1  ( .A1(\SB1_3_0/i0_0 ), .A2(
        \SB1_3_0/i3[0] ), .ZN(\SB1_3_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U1025 ( .A1(\SB2_3_30/i1_5 ), .A2(\SB2_3_30/i0[8] ), .A3(
        \SB2_3_30/i3[0] ), .ZN(\SB2_3_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_4_14/Component_Function_5/N4  ( .A1(\SB1_4_14/i0[9] ), .A2(
        \SB1_4_14/i0[6] ), .A3(\SB1_4_14/i0_4 ), .ZN(
        \SB1_4_14/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U1104 ( .A1(\SB1_1_9/i0[10] ), .A2(\SB1_1_9/i0[6] ), .A3(
        \SB1_1_9/i0_0 ), .ZN(n1878) );
  INV_X2 U7644 ( .I(\SB1_3_3/buf_output[3] ), .ZN(\SB2_3_1/i0[8] ) );
  NAND3_X2 \SB2_1_21/Component_Function_3/N4  ( .A1(\SB2_1_21/i1_5 ), .A2(
        \SB2_1_21/i0[8] ), .A3(\SB2_1_21/i3[0] ), .ZN(
        \SB2_1_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_1_13/Component_Function_2/N2  ( .A1(\SB1_1_13/i0_3 ), .A2(
        \SB1_1_13/i0[10] ), .A3(\SB1_1_13/i0[6] ), .ZN(
        \SB1_1_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U5022 ( .A1(\SB3_19/i0_0 ), .A2(\SB3_19/i1_5 ), .A3(\SB3_19/i0_4 ), 
        .ZN(\SB3_19/Component_Function_2/NAND4_in[3] ) );
  INV_X2 U2442 ( .I(\MC_ARK_ARC_1_4/buf_output[117] ), .ZN(\SB3_12/i0[8] ) );
  INV_X4 \SB1_1_18/INV_4  ( .I(\SB1_1_18/i0_4 ), .ZN(\SB1_1_18/i0[7] ) );
  NAND3_X2 \SB2_4_17/Component_Function_3/N4  ( .A1(\SB2_4_17/i1_5 ), .A2(
        \SB2_4_17/i0[8] ), .A3(\SB2_4_17/i3[0] ), .ZN(
        \SB2_4_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U1657 ( .A1(\SB2_1_12/i0[10] ), .A2(\SB2_1_12/i0_3 ), .A3(
        \SB2_1_12/i0[9] ), .ZN(n3744) );
  NAND3_X2 U791 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0_0 ), .A3(
        \SB2_3_18/i0_4 ), .ZN(\SB2_3_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_2_12/Component_Function_3/N2  ( .A1(\RI1[2][116] ), .A2(
        \RI1[2][119] ), .A3(\SB1_2_12/i0_4 ), .ZN(
        \SB1_2_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_4_12/Component_Function_2/N1  ( .A1(\SB2_4_12/i1_5 ), .A2(
        \SB2_4_12/i0[10] ), .A3(\SB2_4_12/i1[9] ), .ZN(
        \SB2_4_12/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_0_3/BUF_1_0  ( .I(\SB2_0_3/buf_output[1] ), .Z(\RI5[0][1] ) );
  NAND4_X2 U7832 ( .A1(\SB2_0_3/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_3/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_0_3/Component_Function_1/NAND4_in[0] ), .A4(n1663), .ZN(
        \SB2_0_3/buf_output[1] ) );
  NAND3_X2 U4866 ( .A1(\SB1_1_23/i0_0 ), .A2(\SB1_1_23/i0[8] ), .A3(
        \SB1_1_23/i0[9] ), .ZN(\SB1_1_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_6/Component_Function_2/N2  ( .A1(\SB2_2_6/i0_3 ), .A2(
        \SB2_2_6/i0[10] ), .A3(\SB2_2_6/i0[6] ), .ZN(
        \SB2_2_6/Component_Function_2/NAND4_in[1] ) );
  BUF_X2 U69 ( .I(Key[6]), .Z(n46) );
  BUF_X2 U192 ( .I(Key[67]), .Z(n135) );
  CLKBUF_X2 U201 ( .I(Key[59]), .Z(n144) );
  NAND3_X2 U2889 ( .A1(\SB2_3_8/i1_5 ), .A2(\SB2_3_8/i0[10] ), .A3(
        \SB2_3_8/i1[9] ), .ZN(\SB2_3_8/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U6421 ( .A1(\SB2_3_5/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_5/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_5/buf_output[0] ) );
  BUF_X4 U1734 ( .I(\MC_ARK_ARC_1_0/buf_output[133] ), .Z(\SB1_1_9/i0[6] ) );
  NAND3_X2 U5407 ( .A1(\SB2_4_5/i1_5 ), .A2(\SB2_4_5/i0[10] ), .A3(
        \SB2_4_5/i1[9] ), .ZN(\SB2_4_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U8094 ( .A1(\SB4_6/i0_3 ), .A2(\SB4_6/i0_4 ), .A3(\SB4_6/i1[9] ), 
        .ZN(n2742) );
  NAND2_X2 \SB1_1_8/Component_Function_0/N1  ( .A1(\SB1_1_8/i0[10] ), .A2(
        \SB1_1_8/i0[9] ), .ZN(\SB1_1_8/Component_Function_0/NAND4_in[0] ) );
  INV_X2 U2584 ( .I(\MC_ARK_ARC_1_2/buf_output[175] ), .ZN(\SB1_3_2/i1_7 ) );
  NAND3_X2 \SB2_2_15/Component_Function_1/N4  ( .A1(\SB2_2_15/i1_7 ), .A2(
        \SB2_2_15/i0[8] ), .A3(\SB2_2_15/i0_4 ), .ZN(
        \SB2_2_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U5957 ( .A1(\SB2_1_20/i0_0 ), .A2(\SB2_1_20/i0_4 ), .A3(
        \SB2_1_20/i1_5 ), .ZN(\SB2_1_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U10870 ( .A1(\SB2_4_30/i0_3 ), .A2(\SB2_4_30/i0[6] ), .A3(
        \SB2_4_30/i1[9] ), .ZN(\SB2_4_30/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 U1750 ( .A1(\SB1_1_8/i0_0 ), .A2(\SB1_1_8/i3[0] ), .ZN(
        \SB1_1_8/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_5/Component_Function_5/N1  ( .A1(\SB2_2_5/i0_0 ), .A2(
        \SB2_2_5/i3[0] ), .ZN(\SB2_2_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U4273 ( .A1(\SB2_1_7/i0[8] ), .A2(\SB2_1_7/i3[0] ), .A3(
        \SB2_1_7/i1_5 ), .ZN(n1224) );
  NAND2_X2 \SB1_3_1/Component_Function_1/N1  ( .A1(\SB1_3_1/i0_3 ), .A2(
        \SB1_3_1/i1[9] ), .ZN(\SB1_3_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U7802 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i0_0 ), .A3(\SB4_28/i0[7] ), 
        .ZN(n3122) );
  NAND3_X2 U6631 ( .A1(\SB2_4_22/i0_0 ), .A2(\SB2_4_22/i1_7 ), .A3(
        \SB2_4_22/i3[0] ), .ZN(\SB2_4_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U9674 ( .A1(\SB1_4_14/i0[7] ), .A2(\SB1_4_14/i0_3 ), .A3(
        \SB1_4_14/i0_0 ), .ZN(\SB1_4_14/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 \SB2_2_6/BUF_1_0  ( .I(\SB2_2_6/buf_output[1] ), .Z(\RI5[2][175] ) );
  NAND4_X2 U6841 ( .A1(\SB2_2_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_6/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_6/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_2_6/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_2_6/buf_output[1] ) );
  NAND3_X2 U1311 ( .A1(\SB1_3_2/i0_3 ), .A2(\SB1_3_2/i0_0 ), .A3(
        \SB1_3_2/i0_4 ), .ZN(n4511) );
  NAND3_X2 U2299 ( .A1(\SB1_3_14/i0_0 ), .A2(\SB1_3_14/i0[9] ), .A3(
        \SB1_3_14/i0[8] ), .ZN(n2486) );
  INV_X2 U2817 ( .I(\SB1_2_26/buf_output[3] ), .ZN(\SB2_2_24/i0[8] ) );
  NAND3_X2 \SB2_2_15/Component_Function_0/N2  ( .A1(\SB2_2_15/i0[8] ), .A2(
        \SB2_2_15/i0[7] ), .A3(\SB2_2_15/i0[6] ), .ZN(
        \SB2_2_15/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U1441 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0_0 ), .A3(
        \SB2_2_12/i0_4 ), .ZN(n5330) );
  NAND4_X2 \SB2_4_31/Component_Function_1/N5  ( .A1(
        \SB2_4_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_4_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_31/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_4_31/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_4_31/buf_output[1] ) );
  NAND3_X2 U3697 ( .A1(\SB2_1_7/i0[6] ), .A2(\SB2_1_7/i1[9] ), .A3(
        \SB2_1_7/i0_3 ), .ZN(n4351) );
  NAND2_X2 \SB1_2_19/Component_Function_1/N1  ( .A1(\SB1_2_19/i0_3 ), .A2(
        \SB1_2_19/i1[9] ), .ZN(\SB1_2_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U7610 ( .A1(\SB2_1_7/i0_3 ), .A2(\SB2_1_7/i0[9] ), .A3(
        \SB2_1_7/i0[10] ), .ZN(\SB2_1_7/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U2265 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0_0 ), .A3(
        \SB2_2_29/i0_4 ), .ZN(\SB2_2_29/Component_Function_3/NAND4_in[1] ) );
  NAND2_X2 \SB1_1_0/Component_Function_1/N1  ( .A1(\SB1_1_0/i0_3 ), .A2(
        \SB1_1_0/i1[9] ), .ZN(\SB1_1_0/Component_Function_1/NAND4_in[0] ) );
  BUF_X4 \SB2_1_12/BUF_3  ( .I(\SB1_1_14/buf_output[3] ), .Z(\SB2_1_12/i0[10] ) );
  BUF_X4 \SB2_2_24/BUF_1  ( .I(\SB1_2_28/buf_output[1] ), .Z(\SB2_2_24/i0[6] )
         );
  BUF_X4 \SB2_4_16/BUF_0  ( .I(\SB1_4_21/buf_output[0] ), .Z(\SB2_4_16/i0[9] )
         );
  BUF_X4 \SB2_1_7/BUF_5  ( .I(\SB1_1_7/buf_output[5] ), .Z(\SB2_1_7/i0_3 ) );
  NAND3_X2 U2890 ( .A1(\SB2_3_8/i0[10] ), .A2(\SB2_3_8/i1[9] ), .A3(
        \SB2_3_8/i1_7 ), .ZN(\SB2_3_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB1_2_27/Component_Function_3/N3  ( .A1(\SB1_2_27/i1[9] ), .A2(
        \SB1_2_27/i1_7 ), .A3(\SB1_2_27/i0[10] ), .ZN(
        \SB1_2_27/Component_Function_3/NAND4_in[2] ) );
  NAND2_X2 U780 ( .A1(\SB1_4_16/i0_0 ), .A2(\SB1_4_16/i3[0] ), .ZN(n4361) );
  NAND2_X2 U3810 ( .A1(\SB1_3_17/i0_0 ), .A2(\SB1_3_17/i3[0] ), .ZN(
        \SB1_3_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U3700 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i0[9] ), .A3(
        \SB2_1_0/i0_3 ), .ZN(\SB2_1_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U9433 ( .A1(\SB2_4_18/i1_5 ), .A2(\SB2_4_18/i0[10] ), .A3(
        \SB2_4_18/i1[9] ), .ZN(\SB2_4_18/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB1_2_27/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[27] ), .Z(
        \SB1_2_27/i0[10] ) );
  BUF_X4 U9703 ( .I(\MC_ARK_ARC_1_3/buf_output[40] ), .Z(\SB1_4_25/i0_4 ) );
  INV_X2 \SB2_2_0/INV_1  ( .I(\SB1_2_4/buf_output[1] ), .ZN(\SB2_2_0/i1_7 ) );
  NAND3_X2 \SB2_3_7/Component_Function_3/N4  ( .A1(\SB2_3_7/i1_5 ), .A2(
        \SB2_3_7/i0[8] ), .A3(\SB2_3_7/i3[0] ), .ZN(
        \SB2_3_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_2_23/Component_Function_3/N2  ( .A1(\SB1_2_23/i0_0 ), .A2(
        \SB1_2_23/i0_3 ), .A3(\SB1_2_23/i0_4 ), .ZN(
        \SB1_2_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U1185 ( .A1(\SB2_0_7/i0_3 ), .A2(\SB2_0_7/i0[10] ), .A3(
        \SB2_0_7/i0[9] ), .ZN(\SB2_0_7/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U2854 ( .A1(\SB2_4_10/i0_0 ), .A2(\SB2_4_10/i0_3 ), .A3(
        \SB2_4_10/i0_4 ), .ZN(\SB2_4_10/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB2_0_14/BUF_2_0  ( .I(\SB2_0_14/buf_output[2] ), .Z(\RI5[0][122] )
         );
  NAND3_X2 U2619 ( .A1(\SB1_4_19/i0_0 ), .A2(\SB1_4_19/i0[6] ), .A3(
        \SB1_4_19/i0[10] ), .ZN(\SB1_4_19/Component_Function_5/NAND4_in[1] )
         );
  NAND2_X2 \SB2_2_7/Component_Function_0/N1  ( .A1(\SB2_2_7/i0[10] ), .A2(
        \SB2_2_7/i0[9] ), .ZN(\SB2_2_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_27/Component_Function_1/N2  ( .A1(\SB2_3_27/i0_3 ), .A2(
        \SB2_3_27/i1_7 ), .A3(\SB2_3_27/i0[8] ), .ZN(
        \SB2_3_27/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U6238 ( .A1(\SB1_1_25/i0_3 ), .A2(\SB1_1_25/i0[9] ), .A3(
        \SB1_1_25/i0[8] ), .ZN(\SB1_1_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U2564 ( .A1(\SB3_3/i0[10] ), .A2(\SB3_3/i1[9] ), .A3(\SB3_3/i1_5 ), 
        .ZN(n4966) );
  NAND2_X2 \SB1_2_26/Component_Function_5/N1  ( .A1(\SB1_2_26/i0_0 ), .A2(
        \SB1_2_26/i3[0] ), .ZN(\SB1_2_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U6239 ( .A1(\SB1_2_11/i0[6] ), .A2(\SB1_2_11/i1[9] ), .A3(
        \SB1_2_11/i0_3 ), .ZN(\SB1_2_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_31/Component_Function_2/N4  ( .A1(\SB2_3_31/i1_5 ), .A2(
        \SB2_3_31/i0_0 ), .A3(\SB2_3_31/i0_4 ), .ZN(
        \SB2_3_31/Component_Function_2/NAND4_in[3] ) );
  INV_X2 U9744 ( .I(n247), .ZN(\SB1_0_5/i1_7 ) );
  NAND2_X2 U6819 ( .A1(\SB1_2_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_2/Component_Function_4/NAND4_in[1] ), .ZN(n2111) );
  BUF_X4 \SB1_1_29/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[16] ), .Z(
        \SB1_1_29/i0_4 ) );
  BUF_X4 U3421 ( .I(\MC_ARK_ARC_1_3/buf_output[104] ), .Z(\SB1_4_14/i0_0 ) );
  NAND3_X2 U650 ( .A1(\SB2_4_22/i1_5 ), .A2(\SB2_4_22/i0[8] ), .A3(
        \SB2_4_22/i3[0] ), .ZN(\SB2_4_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB2_0_5/Component_Function_2/N2  ( .A1(\SB2_0_5/i0_3 ), .A2(
        \SB2_0_5/i0[10] ), .A3(\SB2_0_5/i0[6] ), .ZN(
        \SB2_0_5/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U5324 ( .I(\MC_ARK_ARC_1_0/buf_output[88] ), .Z(\SB1_1_17/i0_4 ) );
  NAND3_X2 \SB2_1_19/Component_Function_4/N4  ( .A1(\SB2_1_19/i1[9] ), .A2(
        \SB2_1_19/i1_5 ), .A3(\SB2_1_19/i0_4 ), .ZN(
        \SB2_1_19/Component_Function_4/NAND4_in[3] ) );
  INV_X2 U3283 ( .I(\MC_ARK_ARC_1_0/buf_output[171] ), .ZN(\SB1_1_3/i0[8] ) );
  INV_X2 U577 ( .I(\SB3_21/buf_output[3] ), .ZN(\SB4_19/i0[8] ) );
  NAND3_X2 \SB2_4_5/Component_Function_3/N3  ( .A1(\SB2_4_5/i1[9] ), .A2(
        \SB2_4_5/i1_7 ), .A3(\SB2_4_5/i0[10] ), .ZN(
        \SB2_4_5/Component_Function_3/NAND4_in[2] ) );
  CLKBUF_X2 U625 ( .I(Key[172]), .Z(n184) );
  NAND3_X2 U3500 ( .A1(\SB2_2_2/i3[0] ), .A2(\SB2_2_2/i1_5 ), .A3(
        \SB2_2_2/i0[8] ), .ZN(n1704) );
  NAND3_X2 \SB1_1_16/Component_Function_2/N2  ( .A1(\SB1_1_16/i0_3 ), .A2(
        \SB1_1_16/i0[10] ), .A3(\SB1_1_16/i0[6] ), .ZN(
        \SB1_1_16/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_5/Component_Function_5/N1  ( .A1(\SB1_0_5/i0_0 ), .A2(
        \SB1_0_5/i3[0] ), .ZN(\SB1_0_5/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 U3668 ( .A1(\SB2_1_1/i0[9] ), .A2(\SB2_1_1/i0[8] ), .ZN(n1666) );
  NAND3_X2 U4415 ( .A1(\SB2_4_5/i0_3 ), .A2(\SB2_4_5/i1[9] ), .A3(
        \SB1_4_6/buf_output[4] ), .ZN(
        \SB2_4_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U2779 ( .A1(\SB3_26/i0[10] ), .A2(\SB3_26/i0_3 ), .A3(
        \SB3_26/i0[6] ), .ZN(\SB3_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U1705 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i0_4 ), .A3(
        \SB1_1_16/i1[9] ), .ZN(\SB1_1_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U3657 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i0[6] ), .A3(
        \SB1_1_16/i1[9] ), .ZN(n3208) );
  NAND3_X2 \SB2_2_16/Component_Function_5/N4  ( .A1(\SB2_2_16/i0[9] ), .A2(
        \SB2_2_16/i0[6] ), .A3(\SB1_2_17/buf_output[4] ), .ZN(
        \SB2_2_16/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U2329 ( .A1(\SB2_3_31/i1_7 ), .A2(\SB2_3_31/i0[8] ), .A3(
        \SB2_3_31/i0_4 ), .ZN(\SB2_3_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U3619 ( .A1(\SB1_1_0/i1[9] ), .A2(\SB1_1_0/i0_3 ), .A3(
        \SB1_1_0/i0[6] ), .ZN(\SB1_1_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U2910 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0_0 ), .A3(
        \SB2_3_31/i0_4 ), .ZN(\SB2_3_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U584 ( .A1(\SB3_25/i0[6] ), .A2(\SB3_25/i1[9] ), .A3(\SB3_25/i0_3 ), 
        .ZN(\SB3_25/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_4_29/BUF_5  ( .I(\SB1_4_29/buf_output[5] ), .Z(\SB2_4_29/i0_3 )
         );
  BUF_X4 U2807 ( .I(\SB1_3_31/buf_output[5] ), .Z(\SB2_3_31/i0_3 ) );
  CLKBUF_X4 U9435 ( .I(\MC_ARK_ARC_1_4/buf_output[28] ), .Z(\SB3_27/i0_4 ) );
  CLKBUF_X4 \SB2_4_6/BUF_4  ( .I(\SB1_4_7/buf_output[4] ), .Z(\SB2_4_6/i0_4 )
         );
  CLKBUF_X8 U3416 ( .I(\RI1[4][5] ), .Z(\SB1_4_31/i0_3 ) );
  CLKBUF_X2 U212 ( .I(Key[119]), .Z(n159) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_37  ( .I(\SB2_3_29/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[37] ) );
  NAND3_X2 \SB2_0_25/Component_Function_5/N2  ( .A1(\SB2_0_25/i0_0 ), .A2(
        \SB2_0_25/i0[6] ), .A3(\SB2_0_25/i0[10] ), .ZN(
        \SB2_0_25/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U9428 ( .A1(\SB2_3_13/i1[9] ), .A2(n6746), .A3(\SB2_3_13/i0_3 ), 
        .ZN(\SB2_3_13/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_0_25/BUF_3  ( .I(\RI3[0][39] ), .Z(\SB2_0_25/i0[10] ) );
  NAND3_X2 \SB3_25/Component_Function_3/N2  ( .A1(\SB3_25/i0_0 ), .A2(
        \SB3_25/i0_3 ), .A3(\SB3_25/i0_4 ), .ZN(
        \SB3_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U8411 ( .A1(\SB1_0_6/i0_0 ), .A2(\SB1_0_6/i1_5 ), .A3(
        \SB1_0_6/i0_4 ), .ZN(n2918) );
  NAND3_X2 U826 ( .A1(\SB2_3_8/i0[6] ), .A2(\SB2_3_8/i0_3 ), .A3(
        \SB2_3_8/i1[9] ), .ZN(\SB2_3_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_19/Component_Function_1/N3  ( .A1(\SB2_2_19/i1_5 ), .A2(
        \SB2_2_19/i0[6] ), .A3(\SB2_2_19/i0[9] ), .ZN(
        \SB2_2_19/Component_Function_1/NAND4_in[2] ) );
  INV_X2 \SB2_2_19/INV_5  ( .I(\SB1_2_19/buf_output[5] ), .ZN(\SB2_2_19/i1_5 )
         );
  NAND3_X2 U2202 ( .A1(\SB2_1_31/i0[9] ), .A2(\SB2_1_31/i0_3 ), .A3(
        \SB2_1_31/i0[8] ), .ZN(\SB2_1_31/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X2 U245 ( .I(Key[15]), .Z(n204) );
  BUF_X4 U5204 ( .I(\SB2_3_8/buf_output[1] ), .Z(\RI5[3][163] ) );
  NAND4_X2 U1008 ( .A1(\SB2_3_8/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_8/Component_Function_1/NAND4_in[1] ), .A3(n4512), .A4(
        \SB2_3_8/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_8/buf_output[1] ) );
  NAND3_X2 U3232 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i0[10] ), .A3(
        \SB1_2_5/i0[6] ), .ZN(\SB1_2_5/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U1151 ( .I(\SB1_3_5/buf_output[0] ), .Z(\SB2_3_0/i0[9] ) );
  NAND3_X2 U3899 ( .A1(\SB1_4_3/i0[9] ), .A2(\SB1_4_3/i0[10] ), .A3(
        \SB1_4_3/i0_3 ), .ZN(\SB1_4_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_14/Component_Function_1/N4  ( .A1(\SB2_1_14/i1_7 ), .A2(
        \SB2_1_14/i0[8] ), .A3(\SB2_1_14/i0_4 ), .ZN(
        \SB2_1_14/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 U5427 ( .I(\SB2_1_16/buf_output[0] ), .Z(\RI5[1][120] ) );
  NAND3_X2 U2915 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0[8] ), .A3(
        \SB2_3_31/i0[9] ), .ZN(\SB2_3_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U1818 ( .A1(\SB2_4_25/i0[10] ), .A2(\SB2_4_25/i1_5 ), .A3(
        \SB2_4_25/i1[9] ), .ZN(\SB2_4_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_0_4/Component_Function_0/N3  ( .A1(\SB1_0_4/i0[10] ), .A2(
        \SB1_0_4/i0_4 ), .A3(\SB1_0_4/i0_3 ), .ZN(
        \SB1_0_4/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 U3354 ( .I(\SB3_21/buf_output[3] ), .Z(\SB4_19/i0[10] ) );
  NAND3_X2 U675 ( .A1(\SB2_4_25/i0[9] ), .A2(\SB2_4_25/i0_3 ), .A3(
        \SB2_4_25/i0[8] ), .ZN(n935) );
  NAND3_X2 U682 ( .A1(\SB2_4_25/i1_5 ), .A2(\SB2_4_25/i3[0] ), .A3(
        \SB2_4_25/i0[8] ), .ZN(n3039) );
  BUF_X4 \SB2_4_30/BUF_3_0  ( .I(\SB2_4_30/buf_output[3] ), .Z(\RI5[4][21] )
         );
  NAND4_X2 U8020 ( .A1(\SB2_4_30/Component_Function_3/NAND4_in[3] ), .A2(n2924), .A3(n2683), .A4(\SB2_4_30/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB2_4_30/buf_output[3] ) );
  NAND3_X2 U9419 ( .A1(\SB3_13/i0[10] ), .A2(\SB3_13/i1_5 ), .A3(
        \SB3_13/i1[9] ), .ZN(\SB3_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB3_13/Component_Function_2/N2  ( .A1(\SB3_13/i0_3 ), .A2(
        \SB3_13/i0[10] ), .A3(\SB3_13/i0[6] ), .ZN(
        \SB3_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U1139 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i1[9] ), .A3(
        \SB2_3_31/i0_4 ), .ZN(n3162) );
  NAND3_X2 U12349 ( .A1(\SB2_2_26/i0[8] ), .A2(\SB2_2_26/i0_3 ), .A3(
        \SB2_2_26/i0[9] ), .ZN(\SB2_2_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_13/Component_Function_2/N1  ( .A1(\SB2_1_13/i1_5 ), .A2(
        \SB2_1_13/i0[10] ), .A3(\SB2_1_13/i1[9] ), .ZN(
        \SB2_1_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_4_16/Component_Function_2/N1  ( .A1(\SB2_4_16/i1_5 ), .A2(
        \SB2_4_16/i0[10] ), .A3(\SB2_4_16/i1[9] ), .ZN(
        \SB2_4_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_6/Component_Function_0/N2  ( .A1(\SB2_1_6/i0[8] ), .A2(
        \SB2_1_6/i0[7] ), .A3(\SB2_1_6/i0[6] ), .ZN(
        \SB2_1_6/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U7276 ( .A1(\SB1_3_14/i0_0 ), .A2(\SB1_3_14/i1_7 ), .A3(
        \SB1_3_14/i3[0] ), .ZN(\SB1_3_14/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 U3195 ( .I(\MC_ARK_ARC_1_2/buf_output[104] ), .Z(\SB1_3_14/i0_0 ) );
  CLKBUF_X4 U3291 ( .I(\SB1_0_5/buf_output[0] ), .Z(\SB2_0_0/i0[9] ) );
  BUF_X4 \SB1_2_21/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[60] ), .Z(
        \SB1_2_21/i0[9] ) );
  BUF_X4 U9523 ( .I(\MC_ARK_ARC_1_4/buf_output[183] ), .Z(\SB3_1/i0[10] ) );
  NAND3_X2 U1241 ( .A1(\SB1_0_7/i0[10] ), .A2(\SB1_0_7/i0_3 ), .A3(
        \SB1_0_7/i0[9] ), .ZN(n1333) );
  NAND3_X2 U3032 ( .A1(\SB1_2_26/i0_0 ), .A2(\SB1_2_26/i0_4 ), .A3(
        \SB1_2_26/i1_5 ), .ZN(\SB1_2_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB1_2_26/Component_Function_1/N4  ( .A1(\SB1_2_26/i1_7 ), .A2(
        \SB1_2_26/i0[8] ), .A3(\SB1_2_26/i0_4 ), .ZN(
        \SB1_2_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U2272 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0[10] ), .A3(
        \SB2_2_29/i0[9] ), .ZN(n2429) );
  NAND3_X2 U3731 ( .A1(\SB2_4_16/i0_0 ), .A2(\SB2_4_16/i0_4 ), .A3(
        \SB2_4_16/i1_5 ), .ZN(n1027) );
  NAND3_X2 \SB2_3_25/Component_Function_4/N1  ( .A1(n5432), .A2(
        \SB2_3_25/i0_0 ), .A3(\SB2_3_25/i0[8] ), .ZN(
        \SB2_3_25/Component_Function_4/NAND4_in[0] ) );
  INV_X4 \SB2_2_7/INV_5  ( .I(n6737), .ZN(\SB2_2_7/i1_5 ) );
  NAND3_X2 U7263 ( .A1(\SB2_3_1/i0[9] ), .A2(\SB2_3_1/i0_3 ), .A3(
        \SB2_3_1/i0[8] ), .ZN(\SB2_3_1/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB1_1_28/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[20] ), .Z(
        \SB1_1_28/i0_0 ) );
  BUF_X4 \SB1_0_14/BUF_4_0  ( .I(\SB1_0_14/buf_output[4] ), .Z(\RI3[0][112] )
         );
  BUF_X4 U645 ( .I(\SB2_4_31/buf_output[1] ), .Z(\RI5[4][25] ) );
  NAND4_X2 \SB2_0_1/Component_Function_4/N5  ( .A1(
        \SB2_0_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_1/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_0_1/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_0_1/buf_output[4] ) );
  NAND3_X2 U8232 ( .A1(\SB2_3_30/i0[10] ), .A2(\SB2_3_30/i0_3 ), .A3(
        \SB2_3_30/i0[6] ), .ZN(\SB2_3_30/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_0_1/BUF_4_0  ( .I(\SB2_0_1/buf_output[4] ), .Z(\RI5[0][190] ) );
  NAND3_X2 U1087 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0_4 ), .A3(
        \SB2_3_15/i1[9] ), .ZN(n4672) );
  INV_X4 \SB2_0_16/INV_4  ( .I(n594), .ZN(\SB2_0_16/i0[7] ) );
  NAND3_X2 U2435 ( .A1(\SB3_18/i0[7] ), .A2(\SB3_18/i0_3 ), .A3(\SB3_18/i0_0 ), 
        .ZN(\SB3_18/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 \SB1_0_17/BUF_2  ( .I(n282), .Z(\SB1_0_17/i0_0 ) );
  CLKBUF_X2 U234 ( .I(Key[34]), .Z(n189) );
  NAND3_X2 \SB2_3_9/Component_Function_0/N2  ( .A1(\SB2_3_9/i0[8] ), .A2(n1953), .A3(\SB2_3_9/i0[6] ), .ZN(\SB2_3_9/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_25/Component_Function_3/N4  ( .A1(\SB2_2_25/i1_5 ), .A2(
        \SB2_2_25/i0[8] ), .A3(\SB2_2_25/i3[0] ), .ZN(
        \SB2_2_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U1828 ( .A1(\SB2_2_13/i1[9] ), .A2(\SB2_2_13/i1_7 ), .A3(
        \SB2_2_13/i0[10] ), .ZN(\SB2_2_13/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X2 U1371 ( .A1(\SB1_3_12/i0[8] ), .A2(\SB1_3_12/i3[0] ), .A3(
        \SB1_3_12/i1_5 ), .ZN(\SB1_3_12/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB1_2_8/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[141] ), .Z(
        \SB1_2_8/i0[10] ) );
  BUF_X4 U5076 ( .I(\MC_ARK_ARC_1_2/buf_output[15] ), .Z(\SB1_3_29/i0[10] ) );
  NAND3_X2 U2918 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0[10] ), .A3(
        \SB2_3_31/i0[9] ), .ZN(\SB2_3_31/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 U3348 ( .I(\RI5[1][8] ), .Z(n3167) );
  CLKBUF_X4 U2954 ( .I(\SB1_4_27/buf_output[3] ), .Z(\SB2_4_25/i0[10] ) );
  NAND4_X2 U9104 ( .A1(\SB2_3_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_3/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_3/buf_output[1] ) );
  NAND3_X2 \SB2_0_2/Component_Function_3/N2  ( .A1(\SB2_0_2/i0_0 ), .A2(
        \SB2_0_2/i0_3 ), .A3(\RI3[0][178] ), .ZN(
        \SB2_0_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_4_26/Component_Function_2/N1  ( .A1(\SB1_4_26/i1_5 ), .A2(
        \SB1_4_26/i0[10] ), .A3(\SB1_4_26/i1[9] ), .ZN(
        \SB1_4_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U3855 ( .A1(\SB2_3_28/i0[8] ), .A2(\SB2_3_28/i3[0] ), .A3(
        \SB2_3_28/i1_5 ), .ZN(n5296) );
  BUF_X4 \SB1_1_18/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[82] ), .Z(
        \SB1_1_18/i0_4 ) );
  INV_X2 U3215 ( .I(\MC_ARK_ARC_1_3/buf_output[149] ), .ZN(\SB1_4_7/i1_5 ) );
  NAND3_X2 \SB2_4_5/Component_Function_4/N3  ( .A1(\SB2_4_5/i0[9] ), .A2(
        \SB2_4_5/i0[10] ), .A3(\SB2_4_5/i0_3 ), .ZN(
        \SB2_4_5/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 \SB1_1_4/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[166] ), .Z(
        \SB1_1_4/i0_4 ) );
  BUF_X4 \SB1_3_12/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[118] ), .Z(
        \SB1_3_12/i0_4 ) );
  CLKBUF_X4 \SB2_0_29/BUF_3  ( .I(\RI3[0][15] ), .Z(\SB2_0_29/i0[10] ) );
  NAND3_X2 U9979 ( .A1(\SB2_4_28/i0_4 ), .A2(\SB1_4_28/buf_output[5] ), .A3(
        \SB2_4_28/i1[9] ), .ZN(n4531) );
  BUF_X4 U9375 ( .I(\MC_ARK_ARC_1_2/buf_output[9] ), .Z(\SB1_3_30/i0[10] ) );
  BUF_X4 \SB1_3_20/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[68] ), .Z(
        \SB1_3_20/i0_0 ) );
  INV_X2 \SB1_0_16/INV_0  ( .I(n6149), .ZN(\SB1_0_16/i3[0] ) );
  NAND3_X1 U7636 ( .A1(\SB2_2_6/i0_0 ), .A2(\SB2_2_6/i1_5 ), .A3(
        \SB2_2_6/i0_4 ), .ZN(\SB2_2_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U7484 ( .A1(\SB2_0_12/i0[9] ), .A2(\SB2_0_12/i0[6] ), .A3(
        \RI3[0][118] ), .ZN(n2418) );
  NAND3_X2 U1682 ( .A1(\SB2_1_8/i0_0 ), .A2(\SB2_1_8/i1_7 ), .A3(
        \SB2_1_8/i3[0] ), .ZN(\SB2_1_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_4/Component_Function_0/N3  ( .A1(\SB2_0_4/i0[10] ), .A2(
        \RI3[0][166] ), .A3(\SB2_0_4/i0_3 ), .ZN(
        \SB2_0_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_5/Component_Function_4/N4  ( .A1(\SB2_0_5/i1[9] ), .A2(n6282), .A3(\SB2_0_5/i0_4 ), .ZN(\SB2_0_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB1_3_30/Component_Function_2/N3  ( .A1(\SB1_3_30/i0_3 ), .A2(
        \SB1_3_30/i0[8] ), .A3(\SB1_3_30/i0[9] ), .ZN(
        \SB1_3_30/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 \SB2_4_28/BUF_3  ( .I(\SB1_4_30/buf_output[3] ), .Z(\SB2_4_28/i0[10] ) );
  NAND3_X2 U9388 ( .A1(\SB2_4_6/i0_3 ), .A2(\SB2_4_6/i0[8] ), .A3(
        \SB2_4_6/i0[9] ), .ZN(\SB2_4_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U1101 ( .A1(\SB2_3_30/i1_5 ), .A2(\SB2_3_30/i0[10] ), .A3(
        \SB2_3_30/i1[9] ), .ZN(\SB2_3_30/Component_Function_2/NAND4_in[0] ) );
  INV_X2 \SB2_0_29/INV_5  ( .I(\SB1_0_29/buf_output[5] ), .ZN(\SB2_0_29/i1_5 )
         );
  NAND3_X2 U1703 ( .A1(\SB1_1_16/i0_4 ), .A2(\SB1_1_16/i0[9] ), .A3(
        \SB1_1_16/i0[6] ), .ZN(n2764) );
  NAND3_X2 U12309 ( .A1(\SB1_0_29/i0[10] ), .A2(\SB1_0_29/i0_0 ), .A3(
        \SB1_0_29/i0[6] ), .ZN(\SB1_0_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_29/Component_Function_3/N2  ( .A1(\SB2_0_29/i0_0 ), .A2(
        \SB2_0_29/i0_3 ), .A3(\SB2_0_29/i0_4 ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U2793 ( .I(n6286), .ZN(\SB3_11/i0[8] ) );
  BUF_X4 \SB1_2_14/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[106] ), .Z(
        \SB1_2_14/i0_4 ) );
  NAND3_X2 U5648 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0_0 ), .A3(
        \SB2_2_24/i0[7] ), .ZN(n1584) );
  BUF_X4 U2790 ( .I(\MC_ARK_ARC_1_4/buf_output[123] ), .Z(\SB3_11/i0[10] ) );
  NAND3_X2 \SB2_1_31/Component_Function_2/N4  ( .A1(\SB2_1_31/i1_5 ), .A2(
        \SB2_1_31/i0_0 ), .A3(n5429), .ZN(
        \SB2_1_31/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 \SB1_0_29/Component_Function_5/N1  ( .A1(\SB1_0_29/i0_0 ), .A2(
        \SB1_0_29/i3[0] ), .ZN(\SB1_0_29/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_1_28/BUF_4  ( .I(\SB1_1_29/buf_output[4] ), .Z(\SB2_1_28/i0_4 )
         );
  CLKBUF_X4 U5030 ( .I(\SB1_4_19/buf_output[4] ), .Z(\SB2_4_18/i0_4 ) );
  NAND3_X2 \SB2_4_18/Component_Function_3/N1  ( .A1(\SB2_4_18/i1[9] ), .A2(
        \SB2_4_18/i0_3 ), .A3(\SB2_4_18/i0[6] ), .ZN(
        \SB2_4_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB1_3_30/Component_Function_0/N4  ( .A1(\SB1_3_30/i0[7] ), .A2(
        \SB1_3_30/i0_3 ), .A3(\SB1_3_30/i0_0 ), .ZN(
        \SB1_3_30/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 \SB1_4_9/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[132] ), .Z(
        \SB1_4_9/i0[9] ) );
  NAND3_X2 U1378 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i0_3 ), .A3(
        \SB2_2_27/i0[6] ), .ZN(n4223) );
  NAND3_X2 U3155 ( .A1(\SB1_3_20/i1_5 ), .A2(\SB1_3_20/i0[10] ), .A3(
        \SB1_3_20/i1[9] ), .ZN(\SB1_3_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_17/Component_Function_2/N4  ( .A1(\SB2_2_17/i1_5 ), .A2(
        \SB2_2_17/i0_0 ), .A3(\RI3[2][88] ), .ZN(
        \SB2_2_17/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 \SB2_3_27/BUF_0  ( .I(\SB1_3_0/buf_output[0] ), .Z(\SB2_3_27/i0[9] )
         );
  NAND3_X2 U5026 ( .A1(\SB1_4_15/i1[9] ), .A2(\SB1_4_15/i1_7 ), .A3(
        \SB1_4_15/i0[10] ), .ZN(\SB1_4_15/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X2 U1880 ( .A1(\SB2_1_2/i1[9] ), .A2(\SB2_1_2/i0_4 ), .A3(
        \SB2_1_2/i0_3 ), .ZN(\SB2_1_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB1_0_4/Component_Function_5/N2  ( .A1(\SB1_0_4/i0_0 ), .A2(
        \SB1_0_4/i0[6] ), .A3(\SB1_0_4/i0[10] ), .ZN(
        \SB1_0_4/Component_Function_5/NAND4_in[1] ) );
  INV_X4 U1150 ( .I(n6746), .ZN(\SB2_3_13/i0[7] ) );
  NAND3_X2 U1401 ( .A1(\SB4_0/i0_4 ), .A2(\SB4_0/i0[9] ), .A3(\SB4_0/i0[6] ), 
        .ZN(\SB4_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U5329 ( .A1(\SB3_11/i1_5 ), .A2(\SB3_11/i0[10] ), .A3(
        \SB3_11/i1[9] ), .ZN(\SB3_11/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U3917 ( .I(\MC_ARK_ARC_1_3/buf_output[89] ), .ZN(\SB1_4_17/i1_5 ) );
  BUF_X4 \SB2_3_9/BUF_2  ( .I(\SB1_3_12/buf_output[2] ), .Z(\SB2_3_9/i0_0 ) );
  BUF_X2 U593 ( .I(Key[46]), .Z(n181) );
  CLKBUF_X2 U195 ( .I(Key[68]), .Z(n138) );
  CLKBUF_X2 U204 ( .I(Key[110]), .Z(n149) );
  CLKBUF_X12 \SB2_0_20/BUF_0  ( .I(\SB1_0_25/buf_output[0] ), .Z(
        \SB2_0_20/i0[9] ) );
  NAND3_X2 \SB2_0_29/Component_Function_2/N1  ( .A1(\SB2_0_29/i1_5 ), .A2(
        \SB2_0_29/i0[10] ), .A3(\SB2_0_29/i1[9] ), .ZN(
        \SB2_0_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_29/Component_Function_3/N3  ( .A1(\SB2_0_29/i1[9] ), .A2(
        \SB2_0_29/i1_7 ), .A3(\SB2_0_29/i0[10] ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U1177 ( .A1(\SB2_0_26/i0_0 ), .A2(\RI3[0][33] ), .A3(
        \SB2_0_26/i0[6] ), .ZN(\SB2_0_26/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_142  ( .I(\SB2_3_9/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[142] ) );
  NAND3_X2 U5929 ( .A1(\SB2_0_22/i0[8] ), .A2(\SB2_0_22/i0_3 ), .A3(
        \SB2_0_22/i1_7 ), .ZN(\SB2_0_22/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U1098 ( .A1(\SB2_3_6/i0_4 ), .A2(\SB2_3_6/i1_7 ), .A3(
        \SB2_3_6/i0[8] ), .ZN(\SB2_3_6/Component_Function_1/NAND4_in[3] ) );
  INV_X2 U1336 ( .I(\MC_ARK_ARC_1_2/buf_output[145] ), .ZN(\SB1_3_7/i1_7 ) );
  NAND3_X2 U7522 ( .A1(\SB2_0_6/i0_3 ), .A2(\SB2_0_6/i1[9] ), .A3(
        \SB2_0_6/i0[6] ), .ZN(\SB2_0_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_17/Component_Function_3/N1  ( .A1(\SB2_2_17/i1[9] ), .A2(
        \SB2_2_17/i0_3 ), .A3(\SB2_2_17/i0[6] ), .ZN(
        \SB2_2_17/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_0_4/BUF_5  ( .I(\RI3[0][167] ), .Z(\SB2_0_4/i0_3 ) );
  NAND3_X2 U7749 ( .A1(\SB2_3_9/i0_3 ), .A2(\SB2_3_9/i0[10] ), .A3(
        \SB1_3_10/buf_output[4] ), .ZN(n3714) );
  INV_X2 U1618 ( .I(\MC_ARK_ARC_1_4/buf_output[181] ), .ZN(\SB3_1/i1_7 ) );
  NAND3_X2 \SB2_0_29/Component_Function_4/N4  ( .A1(\SB2_0_29/i1[9] ), .A2(
        \SB2_0_29/i1_5 ), .A3(\SB2_0_29/i0_4 ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB2_4_18/Component_Function_2/N3  ( .A1(\SB2_4_18/i0_3 ), .A2(
        \SB2_4_18/i0[8] ), .A3(\SB2_4_18/i0[9] ), .ZN(
        \SB2_4_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U1760 ( .A1(\SB1_1_11/i0[10] ), .A2(\SB1_1_11/i1[9] ), .A3(
        \SB1_1_11/i1_5 ), .ZN(\SB1_1_11/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U9406 ( .I(\SB1_4_6/buf_output[5] ), .Z(\SB2_4_6/i0_3 ) );
  INV_X2 U2695 ( .I(\SB3_27/buf_output[2] ), .ZN(\SB4_24/i1[9] ) );
  NAND3_X2 U10499 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i1_5 ), .A3(\SB3_1/i0_4 ), 
        .ZN(n4293) );
  NAND2_X2 \SB1_1_14/Component_Function_5/N1  ( .A1(\SB1_1_14/i0_0 ), .A2(
        \SB1_1_14/i3[0] ), .ZN(\SB1_1_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U649 ( .A1(\SB3_25/i1[9] ), .A2(\SB3_25/i0_4 ), .A3(\SB3_25/i0_3 ), 
        .ZN(\SB3_25/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U5175 ( .I(\SB3_25/buf_output[1] ), .Z(\SB4_21/i0[6] ) );
  BUF_X4 \SB2_3_25/BUF_1  ( .I(\SB1_3_29/buf_output[1] ), .Z(\SB2_3_25/i0[6] )
         );
  NAND3_X2 \SB1_2_0/Component_Function_5/N3  ( .A1(\SB1_2_0/i1[9] ), .A2(
        \SB1_2_0/i0_4 ), .A3(\RI1[2][191] ), .ZN(
        \SB1_2_0/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB3_22/Component_Function_0/N4  ( .A1(\SB3_22/i0[7] ), .A2(
        \SB3_22/i0_3 ), .A3(\SB3_22/i0_0 ), .ZN(
        \SB3_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 \SB2_4_16/Component_Function_2/N3  ( .A1(\SB2_4_16/i0_3 ), .A2(
        \SB2_4_16/i0[8] ), .A3(\SB2_4_16/i0[9] ), .ZN(
        \SB2_4_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U887 ( .A1(\SB1_3_8/i0[9] ), .A2(\SB1_3_8/i0[6] ), .A3(
        \SB1_3_8/i0_4 ), .ZN(n2306) );
  NAND3_X2 \SB1_0_13/Component_Function_3/N2  ( .A1(\SB1_0_13/i0_0 ), .A2(
        \SB1_0_13/i0_3 ), .A3(\SB1_0_13/i0_4 ), .ZN(
        \SB1_0_13/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB1_0_23/BUF_4_0  ( .I(\SB1_0_23/buf_output[4] ), .Z(\RI3[0][58] )
         );
  NAND2_X2 \SB1_1_18/Component_Function_5/N1  ( .A1(\SB1_1_18/i0_0 ), .A2(
        \SB1_1_18/i3[0] ), .ZN(\SB1_1_18/Component_Function_5/NAND4_in[0] ) );
  INV_X4 U8507 ( .I(n2978), .ZN(\SB2_0_25/i0_4 ) );
  NAND2_X2 U1494 ( .A1(\SB2_2_9/i0[8] ), .A2(\SB2_2_9/i1_7 ), .ZN(n4180) );
  INV_X2 U1842 ( .I(\MC_ARK_ARC_1_3/buf_output[67] ), .ZN(\SB1_4_20/i1_7 ) );
  INV_X2 \SB1_1_30/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[6] ), .ZN(
        \SB1_1_30/i3[0] ) );
  CLKBUF_X2 U156 ( .I(Key[89]), .Z(n98) );
  NAND3_X2 U2326 ( .A1(\SB2_3_26/i1_5 ), .A2(\SB2_3_26/i0[10] ), .A3(
        \SB2_3_26/i1[9] ), .ZN(\SB2_3_26/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U11543 ( .A1(\SB2_4_11/Component_Function_1/NAND4_in[0] ), .A2(
        n2648), .A3(\SB2_4_11/Component_Function_1/NAND4_in[1] ), .A4(n4782), 
        .ZN(\SB2_4_11/buf_output[1] ) );
  NAND3_X2 U8617 ( .A1(\SB1_2_26/i0[10] ), .A2(\SB1_2_26/i1[9] ), .A3(
        \SB1_2_26/i1_5 ), .ZN(\SB1_2_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U3401 ( .A1(\SB1_0_18/i0[6] ), .A2(\SB1_0_18/i1_5 ), .A3(
        \SB1_0_18/i0[9] ), .ZN(n910) );
  INV_X2 \SB1_0_18/INV_5  ( .I(n394), .ZN(\SB1_0_18/i1_5 ) );
  INV_X4 U11297 ( .I(n4662), .ZN(\SB1_0_18/buf_output[2] ) );
  NAND3_X2 \SB1_1_11/Component_Function_3/N3  ( .A1(\SB1_1_11/i1[9] ), .A2(
        \SB1_1_11/i1_7 ), .A3(\SB1_1_11/i0[10] ), .ZN(
        \SB1_1_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_2/Component_Function_3/N1  ( .A1(\SB2_1_2/i1[9] ), .A2(
        \SB2_1_2/i0_3 ), .A3(\SB2_1_2/i0[6] ), .ZN(
        \SB2_1_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U11520 ( .A1(\SB1_2_11/i0[8] ), .A2(\SB1_2_11/i0[9] ), .A3(
        \SB1_2_11/i0_3 ), .ZN(n4777) );
  NAND3_X2 U2173 ( .A1(\SB1_1_23/i0[10] ), .A2(\SB1_1_23/i1[9] ), .A3(
        \SB1_1_23/i1_7 ), .ZN(n2401) );
  INV_X2 \SB1_0_18/INV_1  ( .I(n234), .ZN(\SB1_0_18/i1_7 ) );
  BUF_X4 \SB2_3_5/BUF_3_0  ( .I(\SB2_3_5/buf_output[3] ), .Z(\RI5[3][171] ) );
  NAND2_X2 \SB1_4_27/Component_Function_1/N1  ( .A1(\SB1_4_27/i0_3 ), .A2(
        \SB1_4_27/i1[9] ), .ZN(\SB1_4_27/Component_Function_1/NAND4_in[0] ) );
  NAND2_X2 U2783 ( .A1(\SB2_0_25/i0_0 ), .A2(\SB2_0_25/i3[0] ), .ZN(
        \SB2_0_25/Component_Function_5/NAND4_in[0] ) );
  INV_X4 U1228 ( .I(\SB2_0_17/i0[7] ), .ZN(\RI3[0][88] ) );
  NAND3_X2 \SB1_4_17/Component_Function_1/N3  ( .A1(\SB1_4_17/i1_5 ), .A2(
        \SB1_4_17/i0[6] ), .A3(\SB1_4_17/i0[9] ), .ZN(
        \SB1_4_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_13/Component_Function_0/N3  ( .A1(\SB2_3_13/i0[10] ), .A2(
        n6746), .A3(\SB2_3_13/i0_3 ), .ZN(
        \SB2_3_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_17/Component_Function_1/N3  ( .A1(\SB2_2_17/i1_5 ), .A2(
        \SB2_2_17/i0[6] ), .A3(\SB2_2_17/i0[9] ), .ZN(
        \SB2_2_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB1_3_5/Component_Function_2/N2  ( .A1(\SB1_3_5/i0_3 ), .A2(
        \SB1_3_5/i0[10] ), .A3(\SB1_3_5/i0[6] ), .ZN(
        \SB1_3_5/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_2_31/BUF_4  ( .I(\SB1_2_0/buf_output[4] ), .Z(\SB2_2_31/i0_4 )
         );
  BUF_X2 U3144 ( .I(\RI5[4][175] ), .Z(n3166) );
  BUF_X4 \SB1_0_4/BUF_4  ( .I(n372), .Z(\SB1_0_4/i0_4 ) );
  BUF_X4 \SB2_3_10/BUF_1  ( .I(\SB1_3_14/buf_output[1] ), .Z(\SB2_3_10/i0[6] )
         );
  NAND3_X2 U12137 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i0_0 ), .A3(\SB3_19/i0[7] ), .ZN(n5103) );
  NAND3_X2 U10889 ( .A1(\SB2_1_30/i3[0] ), .A2(\SB2_1_30/i0[8] ), .A3(
        \SB2_1_30/i1_5 ), .ZN(n4470) );
  INV_X2 U4859 ( .I(n3308), .ZN(\SB1_3_29/buf_output[4] ) );
  NAND2_X2 \SB2_1_23/Component_Function_1/N1  ( .A1(\SB2_1_23/i0_3 ), .A2(
        \SB2_1_23/i1[9] ), .ZN(\SB2_1_23/Component_Function_1/NAND4_in[0] ) );
  INV_X1 \SB2_0_26/INV_1  ( .I(\SB1_0_30/buf_output[1] ), .ZN(\SB2_0_26/i1_7 )
         );
  NAND4_X2 U1039 ( .A1(\SB2_1_3/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_3/Component_Function_1/NAND4_in[0] ), .A3(n1612), .A4(
        \SB2_1_3/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_3/buf_output[1] ) );
  NAND3_X2 U1982 ( .A1(\RI3[0][52] ), .A2(\SB2_0_23/i1_5 ), .A3(
        \SB2_0_23/i0_0 ), .ZN(\SB2_0_23/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 U3614 ( .I(\MC_ARK_ARC_1_0/buf_output[71] ), .Z(\SB1_1_20/i0_3 ) );
  NAND3_X2 \SB2_1_31/Component_Function_3/N4  ( .A1(\SB2_1_31/i1_5 ), .A2(
        \SB2_1_31/i0[8] ), .A3(\SB2_1_31/i3[0] ), .ZN(
        \SB2_1_31/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB1_1_31/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[1] ), .Z(
        \SB1_1_31/i0[6] ) );
  AND2_X1 U6585 ( .A1(\SB2_1_1/Component_Function_2/NAND4_in[3] ), .A2(n5001), 
        .Z(n2530) );
  NAND4_X2 U5827 ( .A1(\SB2_0_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_1/Component_Function_2/NAND4_in[1] ), .A3(n3466), .A4(n3465), 
        .ZN(\SB2_0_1/buf_output[2] ) );
  NAND2_X2 \SB1_2_20/Component_Function_5/N1  ( .A1(\SB1_2_20/i0_0 ), .A2(
        \SB1_2_20/i3[0] ), .ZN(\SB1_2_20/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_20/Component_Function_1/N1  ( .A1(\SB2_2_20/i0_3 ), .A2(
        \SB2_2_20/i1[9] ), .ZN(\SB2_2_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U42 ( .A1(\SB4_3/i0_0 ), .A2(\SB4_3/i3[0] ), .A3(\SB4_3/i1_7 ), 
        .ZN(n2026) );
  BUF_X4 U9676 ( .I(\SB1_4_11/buf_output[5] ), .Z(\SB2_4_11/i0_3 ) );
  BUF_X4 \SB2_1_15/BUF_1  ( .I(\SB1_1_19/buf_output[1] ), .Z(\SB2_1_15/i0[6] )
         );
  BUF_X2 U210 ( .I(Key[96]), .Z(n156) );
  CLKBUF_X8 \SB3_23/BUF_5  ( .I(\RI1[5][53] ), .Z(\SB3_23/i0_3 ) );
  NAND3_X1 U7618 ( .A1(\SB2_1_13/i0[10] ), .A2(\SB2_1_13/i1_7 ), .A3(
        \SB2_1_13/i1[9] ), .ZN(n2878) );
  BUF_X4 \SB1_3_8/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[138] ), .Z(
        \SB1_3_8/i0[9] ) );
  BUF_X2 U2196 ( .I(\SB1_1_25/buf_output[0] ), .Z(\SB2_1_20/i0[9] ) );
  INV_X2 \SB2_4_29/INV_1  ( .I(\SB1_4_1/buf_output[1] ), .ZN(\SB2_4_29/i1_7 )
         );
  NAND3_X2 U1164 ( .A1(\SB1_1_3/i0_0 ), .A2(\SB1_1_3/i3[0] ), .A3(
        \SB1_1_3/i1_7 ), .ZN(\SB1_1_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U1193 ( .A1(\SB2_0_22/i0[8] ), .A2(\SB2_0_22/i1_7 ), .A3(
        \RI3[0][58] ), .ZN(\SB2_0_22/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U11627 ( .A1(\SB2_4_29/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_4_29/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_4_29/Component_Function_1/NAND4_in[0] ), .A4(n4832), .ZN(
        \SB2_4_29/buf_output[1] ) );
  NAND3_X2 U3090 ( .A1(\SB2_1_19/i1[9] ), .A2(\SB2_1_19/i0_3 ), .A3(
        \SB2_1_19/i0[6] ), .ZN(\SB2_1_19/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U1695 ( .I(\SB1_2_1/buf_output[3] ), .Z(\SB2_2_31/i0[10] ) );
  BUF_X2 U1886 ( .I(\MC_ARK_ARC_1_0/buf_output[168] ), .Z(\SB1_1_3/i0[9] ) );
  BUF_X4 U5453 ( .I(\MC_ARK_ARC_1_1/buf_output[33] ), .Z(\SB1_2_26/i0[10] ) );
  BUF_X4 U1561 ( .I(\MC_ARK_ARC_1_0/buf_output[31] ), .Z(\SB1_1_26/i0[6] ) );
  CLKBUF_X4 U2936 ( .I(\MC_ARK_ARC_1_0/buf_output[74] ), .Z(\SB1_1_19/i0_0 )
         );
  CLKBUF_X4 U2054 ( .I(\SB2_0_18/buf_output[5] ), .Z(\RI5[0][83] ) );
  NAND3_X2 U1062 ( .A1(\SB2_1_3/i0_4 ), .A2(\SB2_1_3/i0[9] ), .A3(
        \SB2_1_3/i0[6] ), .ZN(n1061) );
  NAND3_X2 \SB1_2_27/Component_Function_4/N4  ( .A1(\SB1_2_27/i1[9] ), .A2(
        \SB1_2_27/i1_5 ), .A3(\SB1_2_27/i0_4 ), .ZN(
        \SB1_2_27/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 U3116 ( .I(\SB1_1_2/buf_output[5] ), .Z(\SB2_1_2/i0_3 ) );
  INV_X4 \SB1_2_29/INV_5  ( .I(\RI1[2][17] ), .ZN(\SB1_2_29/i1_5 ) );
  NAND3_X2 \SB1_0_13/Component_Function_4/N1  ( .A1(\SB1_0_13/i0[9] ), .A2(
        \SB1_0_13/i0_0 ), .A3(n5428), .ZN(
        \SB1_0_13/Component_Function_4/NAND4_in[0] ) );
  BUF_X4 \SB1_1_3/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[170] ), .Z(
        \SB1_1_3/i0_0 ) );
  NAND3_X2 U12515 ( .A1(\SB1_1_22/i0[10] ), .A2(\SB1_1_22/i1[9] ), .A3(
        \SB1_1_22/i1_7 ), .ZN(\SB1_1_22/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB2_0_10/BUF_2_0  ( .I(\SB2_0_10/buf_output[2] ), .Z(\RI5[0][146] )
         );
  INV_X4 U6186 ( .I(\SB2_0_28/i0[7] ), .ZN(\SB2_0_28/i0_4 ) );
  CLKBUF_X4 U9644 ( .I(n374), .Z(\SB1_0_3/i0_4 ) );
  NAND3_X2 U1088 ( .A1(\SB2_3_2/i0_3 ), .A2(\SB2_3_2/i0_0 ), .A3(
        \SB2_3_2/i0_4 ), .ZN(\SB2_3_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U848 ( .A1(\SB1_3_2/i0_3 ), .A2(\SB1_3_2/i0_4 ), .A3(
        \SB1_3_2/i1[9] ), .ZN(n1523) );
  NAND2_X2 U1236 ( .A1(\SB1_3_17/i0_3 ), .A2(\SB1_3_17/i1[9] ), .ZN(n4420) );
  INV_X2 U2673 ( .I(\MC_ARK_ARC_1_1/buf_output[110] ), .ZN(\SB1_2_13/i1[9] )
         );
  BUF_X4 U7087 ( .I(\SB2_4_15/buf_output[1] ), .Z(\RI5[4][121] ) );
  BUF_X4 \SB2_0_6/BUF_1  ( .I(\RI3[0][151] ), .Z(\SB2_0_6/i0[6] ) );
  NAND3_X2 \SB2_2_19/Component_Function_2/N2  ( .A1(\SB2_2_19/i0_3 ), .A2(
        \SB2_2_19/i0[10] ), .A3(\SB2_2_19/i0[6] ), .ZN(
        \SB2_2_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB1_1_14/Component_Function_2/N4  ( .A1(\SB1_1_14/i1_5 ), .A2(
        \SB1_1_14/i0_0 ), .A3(\SB1_1_14/i0_4 ), .ZN(
        \SB1_1_14/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 \SB1_2_7/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[147] ), .Z(
        \SB1_2_7/i0[10] ) );
  BUF_X4 U2252 ( .I(\SB1_2_20/buf_output[2] ), .Z(\SB2_2_17/i0_0 ) );
  CLKBUF_X4 U2008 ( .I(\SB2_2_9/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[147] ) );
  BUF_X2 U79 ( .I(Key[54]), .Z(n38) );
  BUF_X4 U9410 ( .I(\RI1[4][105] ), .Z(\SB1_4_14/i0[10] ) );
  CLKBUF_X4 \SB1_0_25/BUF_4  ( .I(n330), .Z(\SB1_0_25/i0_4 ) );
  NAND2_X1 \SB1_4_26/Component_Function_5/N1  ( .A1(\SB1_4_26/i0_0 ), .A2(
        \SB1_4_26/i3[0] ), .ZN(\SB1_4_26/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_2_11/BUF_1  ( .I(\RI3[2][121] ), .Z(\SB2_2_11/i0[6] ) );
  NAND2_X2 U3694 ( .A1(\SB2_1_0/i0_0 ), .A2(\SB2_1_0/i3[0] ), .ZN(
        \SB2_1_0/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U2927 ( .I(\MC_ARK_ARC_1_3/buf_output[183] ), .Z(\SB1_4_1/i0[10] ) );
  INV_X2 U2928 ( .I(\MC_ARK_ARC_1_3/buf_output[183] ), .ZN(\SB1_4_1/i0[8] ) );
  NAND3_X2 U3988 ( .A1(\SB4_11/i0_3 ), .A2(\SB4_11/i0[9] ), .A3(\SB4_11/i0[8] ), .ZN(\SB4_11/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 U3664 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i1[9] ), .ZN(
        \SB1_1_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB1_3_25/Component_Function_5/N4  ( .A1(\SB1_3_25/i0[9] ), .A2(
        \SB1_3_25/i0[6] ), .A3(\SB1_3_25/i0_4 ), .ZN(
        \SB1_3_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U612 ( .A1(\SB3_27/i0[9] ), .A2(\SB3_27/i0[6] ), .A3(\SB3_27/i1_5 ), 
        .ZN(n3799) );
  NAND3_X2 U627 ( .A1(\SB3_20/i0_3 ), .A2(\SB3_20/i0_4 ), .A3(\SB3_20/i1[9] ), 
        .ZN(n4913) );
  BUF_X2 U1349 ( .I(\SB3_24/buf_output[0] ), .Z(\SB4_19/i0[9] ) );
  NAND3_X2 U2895 ( .A1(\SB1_1_13/i0[8] ), .A2(\SB1_1_13/i3[0] ), .A3(
        \SB1_1_13/i1_5 ), .ZN(\SB1_1_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_1_5/Component_Function_2/N2  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i0[10] ), .A3(\SB1_1_5/i0[6] ), .ZN(
        \SB1_1_5/Component_Function_2/NAND4_in[1] ) );
  INV_X2 \SB1_1_30/INV_5  ( .I(\RI1[1][11] ), .ZN(\SB1_1_30/i1_5 ) );
  NAND3_X2 U2989 ( .A1(\SB4_21/i0[9] ), .A2(\SB4_21/i0_3 ), .A3(
        \SB4_21/i0[10] ), .ZN(n4352) );
  BUF_X4 U3559 ( .I(\RI3[0][47] ), .Z(\SB2_0_24/i0_3 ) );
  BUF_X4 U2236 ( .I(\MC_ARK_ARC_1_1/buf_output[31] ), .Z(\SB1_2_26/i0[6] ) );
  BUF_X4 \SB2_0_26/BUF_1_0  ( .I(\SB2_0_26/buf_output[1] ), .Z(\RI5[0][55] )
         );
  BUF_X4 \SB2_0_11/BUF_3_0  ( .I(\SB2_0_11/buf_output[3] ), .Z(\RI5[0][135] )
         );
  NAND3_X2 \SB2_3_31/Component_Function_3/N4  ( .A1(\SB2_3_31/i1_5 ), .A2(
        \SB2_3_31/i0[8] ), .A3(\SB2_3_31/i3[0] ), .ZN(
        \SB2_3_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U2244 ( .A1(\SB1_2_5/i1_5 ), .A2(\SB1_2_5/i0[10] ), .A3(
        \SB1_2_5/i1[9] ), .ZN(\SB1_2_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U2344 ( .A1(\SB3_22/i0_0 ), .A2(\SB3_22/i1_5 ), .A3(\SB3_22/i0_4 ), 
        .ZN(n4702) );
  NAND3_X2 \SB2_3_22/Component_Function_1/N3  ( .A1(\SB2_3_22/i1_5 ), .A2(
        \SB2_3_22/i0[6] ), .A3(\SB2_3_22/i0[9] ), .ZN(
        \SB2_3_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U6526 ( .A1(\SB1_2_1/i0[6] ), .A2(\SB1_2_1/i0_3 ), .A3(
        \SB1_2_1/i0[10] ), .ZN(\SB1_2_1/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U3339 ( .I(\MC_ARK_ARC_1_1/buf_output[165] ), .Z(\SB1_2_4/i0[10] ) );
  NAND3_X2 \SB4_6/Component_Function_3/N4  ( .A1(\SB4_6/i1_5 ), .A2(
        \SB4_6/i0[8] ), .A3(\SB4_6/i3[0] ), .ZN(
        \SB4_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U1611 ( .A1(\SB1_2_5/i0[10] ), .A2(\SB1_2_5/i1[9] ), .A3(
        \SB1_2_5/i1_7 ), .ZN(n2041) );
  NAND3_X2 \SB1_1_6/Component_Function_1/N3  ( .A1(\SB1_1_6/i1_5 ), .A2(
        \SB1_1_6/i0[6] ), .A3(\SB1_1_6/i0[9] ), .ZN(
        \SB1_1_6/Component_Function_1/NAND4_in[2] ) );
  NAND2_X2 \SB2_4_25/Component_Function_1/N1  ( .A1(\SB2_4_25/i0_3 ), .A2(
        \SB2_4_25/i1[9] ), .ZN(\SB2_4_25/Component_Function_1/NAND4_in[0] ) );
  BUF_X2 U194 ( .I(Key[146]), .Z(n137) );
  NAND3_X2 \SB2_4_0/Component_Function_2/N3  ( .A1(\SB2_4_0/i0_3 ), .A2(
        \SB2_4_0/i0[8] ), .A3(\SB2_4_0/i0[9] ), .ZN(
        \SB2_4_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U1949 ( .A1(\SB2_0_3/i0[10] ), .A2(\SB2_0_3/i0_3 ), .A3(
        \SB2_0_3/i0[9] ), .ZN(n4090) );
  BUF_X4 U3607 ( .I(\SB2_0_26/buf_output[3] ), .Z(\RI5[0][45] ) );
  NAND3_X2 U1061 ( .A1(\SB2_1_30/i0[6] ), .A2(\SB2_1_30/i1_5 ), .A3(
        \SB2_1_30/i0[9] ), .ZN(n1950) );
  NAND3_X2 \SB1_0_30/Component_Function_1/N3  ( .A1(\SB1_0_30/i1_5 ), .A2(
        \SB1_0_30/i0[6] ), .A3(\SB1_0_30/i0[9] ), .ZN(
        \SB1_0_30/Component_Function_1/NAND4_in[2] ) );
  NAND2_X2 U766 ( .A1(\SB1_4_23/i3[0] ), .A2(\SB1_4_23/i0_0 ), .ZN(
        \SB1_4_23/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_30/Component_Function_1/N1  ( .A1(\SB2_2_30/i0_3 ), .A2(
        \SB2_2_30/i1[9] ), .ZN(\SB2_2_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_12/Component_Function_3/N2  ( .A1(\SB1_1_12/i0_0 ), .A2(
        \SB1_1_12/i0_3 ), .A3(\SB1_1_12/i0_4 ), .ZN(
        \SB1_1_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_28/Component_Function_3/N1  ( .A1(\SB1_0_28/i1[9] ), .A2(
        \SB1_0_28/i0_3 ), .A3(\SB1_0_28/i0[6] ), .ZN(
        \SB1_0_28/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U2051 ( .I(\MC_ARK_ARC_1_0/buf_output[37] ), .Z(\SB1_1_25/i0[6] ) );
  CLKBUF_X2 U76 ( .I(Key[100]), .Z(n213) );
  NAND2_X2 U2031 ( .A1(\SB1_0_3/i0_3 ), .A2(\SB1_0_3/i1[9] ), .ZN(
        \SB1_0_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U1034 ( .A1(\SB1_2_10/i0[8] ), .A2(\SB1_2_10/i3[0] ), .A3(
        \SB1_2_10/i1_5 ), .ZN(n1956) );
  BUF_X4 \SB1_3_3/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[172] ), .Z(
        \SB1_3_3/i0_4 ) );
  NAND2_X2 \SB3_22/Component_Function_5/N1  ( .A1(\SB3_22/i0_0 ), .A2(
        \SB3_22/i3[0] ), .ZN(\SB3_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_28/Component_Function_3/N4  ( .A1(\SB2_2_28/i1_5 ), .A2(
        \SB2_2_28/i0[8] ), .A3(\SB2_2_28/i3[0] ), .ZN(
        \SB2_2_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_4_1/Component_Function_5/N3  ( .A1(\SB1_4_1/i1[9] ), .A2(
        \SB1_4_1/i0_4 ), .A3(\SB1_4_1/i0_3 ), .ZN(
        \SB1_4_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U1592 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i0_4 ), .A3(
        \SB1_2_5/i1[9] ), .ZN(\SB1_2_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U6272 ( .A1(\SB1_1_23/i0[10] ), .A2(\SB1_1_23/i1[9] ), .A3(
        \SB1_1_23/i1_5 ), .ZN(\SB1_1_23/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_26/Component_Function_5/N1  ( .A1(\SB2_2_26/i0_0 ), .A2(
        \SB2_2_26/i3[0] ), .ZN(\SB2_2_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U9946 ( .A1(\SB2_2_25/i0[6] ), .A2(\SB2_2_25/i0[8] ), .A3(
        \SB2_2_25/i0[7] ), .ZN(n4063) );
  NAND2_X2 \SB3_17/Component_Function_1/N1  ( .A1(\SB3_17/i0_3 ), .A2(
        \SB3_17/i1[9] ), .ZN(\SB3_17/Component_Function_1/NAND4_in[0] ) );
  NAND2_X2 U9418 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i3[0] ), .ZN(n5037) );
  NAND3_X2 U11299 ( .A1(\SB2_4_21/i0[6] ), .A2(\SB2_4_21/i1_5 ), .A3(
        \SB2_4_21/i0[9] ), .ZN(n4663) );
  BUF_X2 U162 ( .I(Key[70]), .Z(n106) );
  BUF_X4 \SB3_28/BUF_4  ( .I(\MC_ARK_ARC_1_4/buf_output[22] ), .Z(
        \SB3_28/i0_4 ) );
  CLKBUF_X4 \SB2_3_30/BUF_4  ( .I(\SB1_3_31/buf_output[4] ), .Z(
        \SB2_3_30/i0_4 ) );
  NAND3_X2 \SB2_3_18/Component_Function_1/N2  ( .A1(\SB2_3_18/i0_3 ), .A2(
        \SB2_3_18/i1_7 ), .A3(\SB2_3_18/i0[8] ), .ZN(
        \SB2_3_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X2 U7170 ( .A1(n929), .A2(\SB1_2_5/Component_Function_4/NAND4_in[3] ), 
        .ZN(n5015) );
  NAND3_X2 \SB2_0_31/Component_Function_1/N3  ( .A1(\SB2_0_31/i1_5 ), .A2(
        \SB2_0_31/i0[6] ), .A3(\SB2_0_31/i0[9] ), .ZN(
        \SB2_0_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U7697 ( .A1(\SB3_23/i0_0 ), .A2(\SB3_23/i1_5 ), .A3(\SB3_23/i0_4 ), 
        .ZN(\SB3_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_4_15/Component_Function_3/N1  ( .A1(\SB2_4_15/i1[9] ), .A2(
        \SB2_4_15/i0_3 ), .A3(\SB2_4_15/i0[6] ), .ZN(
        \SB2_4_15/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U9737 ( .I(\MC_ARK_ARC_1_4/buf_output[75] ), .ZN(\SB3_19/i0[8] ) );
  BUF_X4 U1621 ( .I(\MC_ARK_ARC_1_3/buf_output[96] ), .Z(\SB1_4_15/i0[9] ) );
  NAND3_X2 \SB4_6/Component_Function_2/N1  ( .A1(\SB4_6/i1_5 ), .A2(
        \SB4_6/i0[10] ), .A3(\SB4_6/i1[9] ), .ZN(
        \SB4_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_31/Component_Function_3/N1  ( .A1(\SB2_0_31/i1[9] ), .A2(
        \SB2_0_31/i0_3 ), .A3(\SB2_0_31/i0[6] ), .ZN(
        \SB2_0_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB4_6/Component_Function_3/N3  ( .A1(\SB4_6/i1[9] ), .A2(
        \SB4_6/i1_7 ), .A3(\SB4_6/i0[10] ), .ZN(
        \SB4_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U3437 ( .A1(\SB2_4_16/i0[10] ), .A2(\SB2_4_16/i1[9] ), .A3(
        \SB2_4_16/i1_7 ), .ZN(n920) );
  INV_X2 \SB2_4_16/INV_1  ( .I(\SB1_4_20/buf_output[1] ), .ZN(\SB2_4_16/i1_7 )
         );
  BUF_X4 \SB1_4_20/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[67] ), .Z(
        \SB1_4_20/i0[6] ) );
  NAND2_X2 \SB2_2_9/Component_Function_5/N1  ( .A1(\SB2_2_9/i0_0 ), .A2(
        \SB2_2_9/i3[0] ), .ZN(\SB2_2_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U2577 ( .A1(\SB1_4_28/i0_3 ), .A2(\SB1_4_28/i1[9] ), .A3(
        \SB1_4_28/i0[6] ), .ZN(\SB1_4_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U8169 ( .A1(\SB2_2_13/i0[10] ), .A2(\SB2_2_13/i0[6] ), .A3(
        \SB2_2_13/i0_0 ), .ZN(\SB2_2_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_13/Component_Function_2/N1  ( .A1(\SB2_2_13/i1_5 ), .A2(
        \SB2_2_13/i0[10] ), .A3(\SB2_2_13/i1[9] ), .ZN(
        \SB2_2_13/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U8211 ( .I(\SB2_1_22/buf_output[1] ), .Z(\RI5[1][79] ) );
  NAND3_X2 U4960 ( .A1(\SB3_20/i1[9] ), .A2(\SB3_20/i1_5 ), .A3(\SB3_20/i0_4 ), 
        .ZN(\SB3_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_30/Component_Function_1/N3  ( .A1(\SB2_2_30/i1_5 ), .A2(
        \SB2_2_30/i0[6] ), .A3(\SB2_2_30/i0[9] ), .ZN(
        \SB2_2_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U7977 ( .A1(\SB2_1_4/i0_4 ), .A2(\SB2_1_4/i0[9] ), .A3(
        \SB1_1_8/buf_output[1] ), .ZN(
        \SB2_1_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U1523 ( .A1(\SB1_2_9/i0_3 ), .A2(\SB1_2_9/i1[9] ), .A3(
        \SB1_2_9/i0[6] ), .ZN(\SB1_2_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U8524 ( .A1(\SB2_3_13/i0[7] ), .A2(\SB2_3_13/i0[6] ), .A3(
        \SB2_3_13/i0[8] ), .ZN(\SB2_3_13/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 \SB1_4_22/Component_Function_2/N1  ( .A1(\SB1_4_22/i1_5 ), .A2(
        \SB1_4_22/i0[10] ), .A3(\SB1_4_22/i1[9] ), .ZN(
        \SB1_4_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U7549 ( .A1(\SB1_0_24/i0_4 ), .A2(\SB1_0_24/i1_7 ), .A3(
        \SB1_0_24/i0[8] ), .ZN(n2447) );
  NAND3_X2 \SB2_3_13/Component_Function_0/N4  ( .A1(\SB2_3_13/i0[7] ), .A2(
        \SB2_3_13/i0_3 ), .A3(\SB2_3_13/i0_0 ), .ZN(
        \SB2_3_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 \SB1_3_17/Component_Function_1/N4  ( .A1(\SB1_3_17/i1_7 ), .A2(
        \SB1_3_17/i0[8] ), .A3(\SB1_3_17/i0_4 ), .ZN(
        \SB1_3_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 \SB2_3_13/Component_Function_3/N4  ( .A1(\SB2_3_13/i1_5 ), .A2(
        \SB2_3_13/i0[8] ), .A3(\SB2_3_13/i3[0] ), .ZN(
        \SB2_3_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U8475 ( .A1(\SB2_4_21/i0_0 ), .A2(\SB2_4_21/i0_4 ), .A3(
        \SB2_4_21/i1_5 ), .ZN(n4159) );
  NAND2_X2 \SB3_18/Component_Function_5/N1  ( .A1(\SB3_18/i0_0 ), .A2(
        \SB3_18/i3[0] ), .ZN(\SB3_18/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 U244 ( .I(Key[141]), .Z(n203) );
  NAND2_X1 U2597 ( .A1(\SB2_4_29/i0_0 ), .A2(\SB2_4_29/i3[0] ), .ZN(
        \SB2_4_29/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 U2950 ( .A1(\SB2_0_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_27/Component_Function_2/NAND4_in[1] ), .A3(n748), .A4(
        \SB2_0_27/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_27/buf_output[2] ) );
  NAND3_X2 U1066 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0[10] ), .A3(
        \SB2_3_18/i0[9] ), .ZN(\SB2_3_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_22/Component_Function_5/N2  ( .A1(\SB2_0_22/i0_0 ), .A2(
        \RI3[0][55] ), .A3(\RI3[0][57] ), .ZN(
        \SB2_0_22/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_2_13/BUF_3  ( .I(\SB1_2_15/buf_output[3] ), .Z(\SB2_2_13/i0[10] ) );
  BUF_X4 \SB2_1_5/BUF_1  ( .I(\SB1_1_9/buf_output[1] ), .Z(\SB2_1_5/i0[6] ) );
  CLKBUF_X4 U6179 ( .I(\RI3[0][189] ), .Z(\SB2_0_0/i0[10] ) );
  BUF_X4 \SB1_4_31/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[3] ), .Z(
        \SB1_4_31/i0[10] ) );
  BUF_X2 U20 ( .I(Key[45]), .Z(n198) );
  CLKBUF_X4 \SB2_3_18/BUF_1  ( .I(\SB1_3_22/buf_output[1] ), .Z(
        \SB2_3_18/i0[6] ) );
  CLKBUF_X2 U243 ( .I(Key[33]), .Z(n201) );
  CLKBUF_X2 U248 ( .I(Key[39]), .Z(n210) );
  CLKBUF_X2 U172 ( .I(Key[152]), .Z(n114) );
  NAND2_X2 \SB2_1_3/Component_Function_5/N1  ( .A1(\SB2_1_3/i0_0 ), .A2(
        \SB2_1_3/i3[0] ), .ZN(\SB2_1_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U11366 ( .A1(\SB2_2_13/i0_3 ), .A2(\SB2_2_13/i0_0 ), .A3(
        \SB2_2_13/i0[7] ), .ZN(n4693) );
  INV_X2 U4955 ( .I(\MC_ARK_ARC_1_4/buf_output[145] ), .ZN(\SB3_7/i1_7 ) );
  NAND3_X2 U7621 ( .A1(\SB2_4_25/i0_4 ), .A2(\SB2_4_25/i0[8] ), .A3(
        \SB2_4_25/i1_7 ), .ZN(n4878) );
  NAND3_X2 \SB2_4_5/Component_Function_1/N2  ( .A1(\SB2_4_5/i0_3 ), .A2(
        \SB2_4_5/i1_7 ), .A3(\SB2_4_5/i0[8] ), .ZN(
        \SB2_4_5/Component_Function_1/NAND4_in[1] ) );
  INV_X2 U12453 ( .I(\SB1_0_14/buf_output[5] ), .ZN(\SB2_0_14/i1_5 ) );
  NAND3_X2 U3568 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i0_4 ), .A3(
        \SB2_0_11/i1[9] ), .ZN(\SB2_0_11/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 \SB2_2_11/BUF_4  ( .I(\SB1_2_12/buf_output[4] ), .Z(
        \SB2_2_11/i0_4 ) );
  CLKBUF_X4 \SB2_4_19/BUF_4  ( .I(\SB1_4_20/buf_output[4] ), .Z(
        \SB2_4_19/i0_4 ) );
  CLKBUF_X4 U4036 ( .I(\MC_ARK_ARC_1_4/buf_output[72] ), .Z(\SB3_19/i0[9] ) );
  BUF_X2 U2004 ( .I(\SB1_3_3/buf_output[1] ), .Z(\SB2_3_31/i0[6] ) );
  BUF_X4 U9716 ( .I(n383), .Z(\SB1_0_29/i0_3 ) );
  NAND3_X2 \SB2_3_5/Component_Function_3/N1  ( .A1(\SB2_3_5/i1[9] ), .A2(
        \SB2_3_5/i0_3 ), .A3(\SB2_3_5/i0[6] ), .ZN(
        \SB2_3_5/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_0_27/BUF_2_0  ( .I(\SB2_0_27/buf_output[2] ), .Z(\RI5[0][44] )
         );
  NAND3_X2 \SB2_0_6/Component_Function_0/N2  ( .A1(\SB2_0_6/i0[8] ), .A2(
        \SB2_0_6/i0[7] ), .A3(\SB2_0_6/i0[6] ), .ZN(
        \SB2_0_6/Component_Function_0/NAND4_in[1] ) );
  CLKBUF_X4 U5165 ( .I(\SB1_4_16/buf_output[2] ), .Z(\SB2_4_13/i0_0 ) );
  NAND2_X2 \SB2_3_2/Component_Function_5/N1  ( .A1(\SB2_3_2/i0_0 ), .A2(
        \SB2_3_2/i3[0] ), .ZN(\SB2_3_2/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U8500 ( .I(\RI1[2][17] ), .ZN(n3839) );
  NAND4_X1 U11976 ( .A1(\SB4_4/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_4/Component_Function_1/NAND4_in[0] ), .ZN(n5010) );
  NAND3_X2 U3068 ( .A1(\SB2_4_10/i0_3 ), .A2(\SB2_4_10/i0[9] ), .A3(
        \SB2_4_10/i0[8] ), .ZN(n788) );
  NAND3_X2 U6678 ( .A1(\SB1_0_25/i0[6] ), .A2(\SB1_0_25/i0[9] ), .A3(
        \SB1_0_25/i0_4 ), .ZN(\SB1_0_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB2_0_5/Component_Function_2/N1  ( .A1(n6282), .A2(
        \SB2_0_5/i0[10] ), .A3(\SB2_0_5/i1[9] ), .ZN(
        \SB2_0_5/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_2_9/BUF_4  ( .I(\SB1_2_10/buf_output[4] ), .Z(\SB2_2_9/i0_4 ) );
  BUF_X4 U1170 ( .I(\MC_ARK_ARC_1_0/buf_output[115] ), .Z(\SB1_1_12/i0[6] ) );
  INV_X2 U3070 ( .I(\MC_ARK_ARC_1_3/buf_output[75] ), .ZN(\SB1_4_19/i0[8] ) );
  NAND3_X1 U11262 ( .A1(\RI3[0][28] ), .A2(\SB2_0_27/i1[9] ), .A3(
        \SB2_0_27/i1_5 ), .ZN(\SB2_0_27/Component_Function_4/NAND4_in[3] ) );
  INV_X2 \SB1_1_27/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[24] ), .ZN(
        \SB1_1_27/i3[0] ) );
  NAND3_X2 U10694 ( .A1(\SB2_2_28/i0_4 ), .A2(\SB2_2_28/i0[8] ), .A3(
        \SB2_2_28/i1_7 ), .ZN(n2237) );
  NAND3_X2 U8300 ( .A1(\SB1_4_16/i0[9] ), .A2(\SB1_4_16/i0_4 ), .A3(
        \SB1_4_16/i0[6] ), .ZN(n3136) );
  NAND3_X2 \SB1_4_1/Component_Function_4/N2  ( .A1(\SB1_4_1/i3[0] ), .A2(
        \SB1_4_1/i0_0 ), .A3(\SB1_4_1/i1_7 ), .ZN(
        \SB1_4_1/Component_Function_4/NAND4_in[1] ) );
  NAND2_X2 \SB1_3_15/Component_Function_5/N1  ( .A1(\SB1_3_15/i0_0 ), .A2(
        \SB1_3_15/i3[0] ), .ZN(\SB1_3_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U3824 ( .A1(\SB1_3_15/i1_5 ), .A2(\SB1_3_15/i0_0 ), .A3(
        \SB1_3_15/i0_4 ), .ZN(\SB1_3_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_28/Component_Function_4/N1  ( .A1(\SB2_2_28/i0[9] ), .A2(
        \SB2_2_28/i0_0 ), .A3(\SB2_2_28/i0[8] ), .ZN(
        \SB2_2_28/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 U2175 ( .A1(n2645), .A2(\SB1_1_20/Component_Function_4/NAND4_in[3] ), .ZN(n2458) );
  NAND2_X2 \SB2_4_17/Component_Function_1/N1  ( .A1(\SB2_4_17/i0_3 ), .A2(
        \SB2_4_17/i1[9] ), .ZN(\SB2_4_17/Component_Function_1/NAND4_in[0] ) );
  BUF_X4 \SB2_0_1/BUF_2_0  ( .I(\SB2_0_1/buf_output[2] ), .Z(\RI5[0][8] ) );
  CLKBUF_X4 \SB2_1_26/BUF_0  ( .I(\SB1_1_31/buf_output[0] ), .Z(
        \SB2_1_26/i0[9] ) );
  CLKBUF_X4 \SB3_6/BUF_5  ( .I(\RI1[5][155] ), .Z(\SB3_6/i0_3 ) );
  NAND3_X2 \SB4_11/Component_Function_5/N4  ( .A1(\SB4_11/i0[9] ), .A2(
        \SB4_11/i0[6] ), .A3(\SB4_11/i0_4 ), .ZN(
        \SB4_11/Component_Function_5/NAND4_in[3] ) );
  INV_X4 U3678 ( .I(\SB2_1_20/i0_4 ), .ZN(\SB2_1_20/i0[7] ) );
  NAND3_X2 U12700 ( .A1(\SB2_4_17/i0_3 ), .A2(\SB2_4_17/i1_7 ), .A3(
        \SB2_4_17/i0[8] ), .ZN(\SB2_4_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_12/Component_Function_3/N1  ( .A1(\SB2_0_12/i1[9] ), .A2(
        \RI3[0][119] ), .A3(\SB2_0_12/i0[6] ), .ZN(
        \SB2_0_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U10386 ( .A1(\SB1_4_30/i0[7] ), .A2(\SB1_4_30/i0_3 ), .A3(
        \SB1_4_30/i0_0 ), .ZN(n4848) );
  NAND3_X2 U8434 ( .A1(\SB2_2_26/i0[10] ), .A2(\SB2_2_26/i0_3 ), .A3(
        \SB2_2_26/i0[6] ), .ZN(\SB2_2_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U2456 ( .A1(\SB4_11/i1_7 ), .A2(\SB4_11/i0[8] ), .A3(\SB4_11/i0_4 ), 
        .ZN(\SB4_11/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 \SB2_0_1/BUF_1_0  ( .I(\SB2_0_1/buf_output[1] ), .Z(\RI5[0][13] ) );
  NAND4_X2 U11634 ( .A1(\SB2_0_1/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_0_1/Component_Function_1/NAND4_in[1] ), .A3(n4835), .A4(
        \SB2_0_1/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_0_1/buf_output[1] ) );
  NAND3_X2 \SB2_3_15/Component_Function_0/N2  ( .A1(\SB2_3_15/i0[8] ), .A2(
        \SB2_3_15/i0[7] ), .A3(\SB2_3_15/i0[6] ), .ZN(
        \SB2_3_15/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U10672 ( .A1(\SB2_0_9/i0[6] ), .A2(\SB2_0_9/i0_3 ), .A3(
        \SB2_0_9/i0[10] ), .ZN(\SB2_0_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U1864 ( .A1(\SB1_1_4/i0[8] ), .A2(\SB1_1_4/i3[0] ), .A3(
        \SB1_1_4/i1_5 ), .ZN(n1693) );
  NAND3_X2 U2669 ( .A1(\SB1_1_24/i0_0 ), .A2(\SB1_1_24/i0[7] ), .A3(
        \RI1[1][47] ), .ZN(n656) );
  NAND3_X2 \SB2_3_15/Component_Function_4/N1  ( .A1(\SB2_3_15/i0[9] ), .A2(
        \SB2_3_15/i0_0 ), .A3(\SB2_3_15/i0[8] ), .ZN(
        \SB2_3_15/Component_Function_4/NAND4_in[0] ) );
  BUF_X4 U1769 ( .I(\MC_ARK_ARC_1_0/buf_output[177] ), .Z(\SB1_1_2/i0[10] ) );
  BUF_X4 U2083 ( .I(n292), .Z(\SB1_0_12/i0_0 ) );
  NAND3_X1 \SB2_1_15/Component_Function_2/N4  ( .A1(\SB2_1_15/i1_5 ), .A2(
        \SB2_1_15/i0_0 ), .A3(\SB2_1_15/i0_4 ), .ZN(
        \SB2_1_15/Component_Function_2/NAND4_in[3] ) );
  CLKBUF_X4 U8664 ( .I(\SB2_2_26/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[60] ) );
  INV_X2 \SB2_1_28/INV_4  ( .I(n5855), .ZN(\SB2_1_28/i0[7] ) );
  NAND3_X2 U10467 ( .A1(\SB2_3_11/i0_0 ), .A2(\SB2_3_11/i0_4 ), .A3(
        \SB2_3_11/i1_5 ), .ZN(n5013) );
  NAND3_X2 U1593 ( .A1(\SB1_4_25/i1[9] ), .A2(\SB1_4_25/i0_4 ), .A3(
        \RI1[4][41] ), .ZN(n3117) );
  BUF_X4 \SB1_1_31/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[4] ), .Z(
        \SB1_1_31/i0_4 ) );
  INV_X2 \SB2_3_25/INV_0  ( .I(n5432), .ZN(\SB2_3_25/i3[0] ) );
  NAND3_X2 U7144 ( .A1(\SB1_1_23/i0_4 ), .A2(\SB1_1_23/i1[9] ), .A3(
        \SB1_1_23/i1_5 ), .ZN(\SB1_1_23/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_151  ( .I(\SB2_3_10/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[151] ) );
  NAND3_X2 U8109 ( .A1(\SB1_0_27/i0_3 ), .A2(\SB1_0_27/i0[9] ), .A3(
        \SB1_0_27/i0[8] ), .ZN(n3773) );
  NAND3_X2 \SB1_3_15/Component_Function_1/N4  ( .A1(\SB1_3_15/i1_7 ), .A2(
        \SB1_3_15/i0[8] ), .A3(\SB1_3_15/i0_4 ), .ZN(
        \SB1_3_15/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_21/Component_Function_5/N1  ( .A1(\SB1_2_21/i0_0 ), .A2(
        \SB1_2_21/i3[0] ), .ZN(\SB1_2_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U10102 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i0[6] ), .A3(
        \SB2_2_27/i1[9] ), .ZN(\SB2_2_27/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_14/Component_Function_5/N1  ( .A1(\SB2_4_14/i0_0 ), .A2(
        \SB2_4_14/i3[0] ), .ZN(\SB2_4_14/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U10974 ( .I(\MC_ARK_ARC_1_1/buf_output[116] ), .Z(\RI1[2][116] )
         );
  BUF_X2 U188 ( .I(Key[137]), .Z(n131) );
  BUF_X2 U158 ( .I(Key[169]), .Z(n101) );
  CLKBUF_X2 U207 ( .I(Key[38]), .Z(n152) );
  CLKBUF_X2 U216 ( .I(Key[11]), .Z(n163) );
  NAND4_X2 U11265 ( .A1(\SB2_3_11/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_11/Component_Function_1/NAND4_in[2] ), .A3(n4643), .A4(
        \SB2_3_11/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_11/buf_output[1] ) );
  BUF_X4 U3318 ( .I(\SB2_1_9/buf_output[4] ), .Z(\RI5[1][142] ) );
  INV_X8 U9361 ( .I(\RI1[3][107] ), .ZN(\SB1_3_14/i1_5 ) );
  BUF_X4 \SB2_2_29/BUF_1  ( .I(\SB1_2_1/buf_output[1] ), .Z(\SB2_2_29/i0[6] )
         );
  CLKBUF_X4 \MC_ARK_ARC_1_4/BUF_63  ( .I(\SB2_4_23/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[63] ) );
  BUF_X4 \SB2_4_18/BUF_0  ( .I(\SB1_4_23/buf_output[0] ), .Z(\SB2_4_18/i0[9] )
         );
  CLKBUF_X4 \SB2_0_15/BUF_3_0  ( .I(\SB2_0_15/buf_output[3] ), .Z(
        \RI5[0][111] ) );
  CLKBUF_X4 U1493 ( .I(\MC_ARK_ARC_1_4/buf_output[93] ), .Z(\SB3_16/i0[10] )
         );
  BUF_X4 \SB2_3_24/BUF_4  ( .I(\SB1_3_25/buf_output[4] ), .Z(\SB2_3_24/i0_4 )
         );
  NAND3_X2 \SB2_0_8/Component_Function_3/N1  ( .A1(\SB2_0_8/i1[9] ), .A2(
        \SB2_0_8/i0_3 ), .A3(\SB2_0_8/i0[6] ), .ZN(
        \SB2_0_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U11124 ( .A1(\SB2_0_8/i3[0] ), .A2(\SB2_0_8/i0[8] ), .A3(
        \SB2_0_8/i1_5 ), .ZN(n4571) );
  NAND3_X2 \SB1_3_15/Component_Function_3/N2  ( .A1(\SB1_3_15/i0_0 ), .A2(
        \SB1_3_15/i0_3 ), .A3(\SB1_3_15/i0_4 ), .ZN(
        \SB1_3_15/Component_Function_3/NAND4_in[1] ) );
  NAND2_X2 \SB1_2_19/Component_Function_5/N1  ( .A1(\SB1_2_19/i0_0 ), .A2(
        \SB1_2_19/i3[0] ), .ZN(\SB1_2_19/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB1_1_5/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[159] ), .Z(
        \SB1_1_5/i0[10] ) );
  BUF_X4 \SB1_1_30/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[10] ), .Z(
        \SB1_1_30/i0_4 ) );
  NAND3_X2 U1509 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i1[9] ), .A3(
        \SB1_2_18/i0[6] ), .ZN(\SB1_2_18/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_2_13/BUF_2  ( .I(\SB1_2_16/buf_output[2] ), .Z(\SB2_2_13/i0_0 )
         );
  BUF_X2 U3557 ( .I(n2611), .Z(n3510) );
  BUF_X4 \SB2_1_15/BUF_4  ( .I(\SB1_1_16/buf_output[4] ), .Z(\SB2_1_15/i0_4 )
         );
  BUF_X2 U3512 ( .I(\RI3[0][90] ), .Z(n5157) );
  INV_X1 U291 ( .I(n46), .ZN(n563) );
  CLKBUF_X4 \SB2_4_20/BUF_0  ( .I(\SB1_4_25/buf_output[0] ), .Z(
        \SB2_4_20/i0[9] ) );
  BUF_X2 U199 ( .I(Key[52]), .Z(n142) );
  CLKBUF_X4 \SB2_1_31/BUF_0_0  ( .I(\SB2_1_31/buf_output[0] ), .Z(\RI5[1][30] ) );
  NAND3_X1 \SB2_0_25/Component_Function_3/N4  ( .A1(\SB2_0_25/i1_5 ), .A2(
        \SB2_0_25/i0[8] ), .A3(\SB2_0_25/i3[0] ), .ZN(
        \SB2_0_25/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X2 U190 ( .I(Key[9]), .Z(n133) );
  NAND3_X2 U2561 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0_0 ), .A3(
        \RI3[0][58] ), .ZN(\SB2_0_22/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 U259 ( .I(\SB3_4/buf_output[1] ), .Z(\SB4_0/i0[6] ) );
  NAND3_X2 \SB2_1_16/Component_Function_2/N1  ( .A1(\SB2_1_16/i1_5 ), .A2(
        \SB2_1_16/i0[10] ), .A3(\SB2_1_16/i1[9] ), .ZN(
        \SB2_1_16/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 \SB1_4_28/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[19] ), .Z(
        \SB1_4_28/i0[6] ) );
  NAND3_X2 U9678 ( .A1(\SB2_4_11/i0_3 ), .A2(\SB2_4_11/i0[10] ), .A3(
        \SB2_4_11/i0[6] ), .ZN(\SB2_4_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U2920 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i1_7 ), .A3(
        \SB2_3_31/i0[8] ), .ZN(\SB2_3_31/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U2041 ( .I(\SB2_1_6/buf_output[2] ), .Z(\RI5[1][170] ) );
  BUF_X4 U5231 ( .I(\MC_ARK_ARC_1_1/buf_output[124] ), .Z(\SB1_2_11/i0_4 ) );
  CLKBUF_X4 \SB2_0_22/BUF_2_0  ( .I(\SB2_0_22/buf_output[2] ), .Z(\RI5[0][74] ) );
  NAND3_X2 \SB2_4_1/Component_Function_2/N3  ( .A1(\SB2_4_1/i0_3 ), .A2(
        \SB2_4_1/i0[8] ), .A3(\SB2_4_1/i0[9] ), .ZN(
        \SB2_4_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_6/Component_Function_3/N4  ( .A1(\SB2_3_6/i1_5 ), .A2(
        \SB2_3_6/i0[8] ), .A3(\SB2_3_6/i3[0] ), .ZN(
        \SB2_3_6/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_3_15/BUF_4  ( .I(\SB1_3_16/buf_output[4] ), .Z(\SB2_3_15/i0_4 )
         );
  NAND3_X2 \SB2_3_5/Component_Function_1/N3  ( .A1(\SB2_3_5/i1_5 ), .A2(
        \SB2_3_5/i0[6] ), .A3(\SB2_3_5/i0[9] ), .ZN(
        \SB2_3_5/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 U5234 ( .I(\SB3_12/buf_output[4] ), .Z(\SB4_11/i0_4 ) );
  NAND2_X1 \SB2_3_14/Component_Function_5/N1  ( .A1(\SB2_3_14/i0_0 ), .A2(
        \SB2_3_14/i3[0] ), .ZN(\SB2_3_14/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_0_7/BUF_5  ( .I(\RI3[0][149] ), .Z(\SB2_0_7/i0_3 ) );
  NAND2_X1 \SB2_1_19/Component_Function_5/N1  ( .A1(\SB2_1_19/i0_0 ), .A2(
        \SB2_1_19/i3[0] ), .ZN(\SB2_1_19/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 U16 ( .I(Key[106]), .Z(n191) );
  CLKBUF_X2 U239 ( .I(Key[184]), .Z(n195) );
  NAND3_X2 U2205 ( .A1(\SB2_1_8/i1[9] ), .A2(\SB2_1_8/i1_5 ), .A3(
        \SB2_1_8/i0_4 ), .ZN(\SB2_1_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U8301 ( .A1(\SB1_3_1/i0[10] ), .A2(\SB1_3_1/i1[9] ), .A3(
        \SB1_3_1/i1_5 ), .ZN(\SB1_3_1/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 \SB2_4_15/BUF_2  ( .I(\SB1_4_18/buf_output[2] ), .Z(
        \SB2_4_15/i0_0 ) );
  BUF_X2 U2488 ( .I(Key[142]), .Z(n217) );
  NAND3_X2 \SB1_3_22/Component_Function_0/N3  ( .A1(\SB1_3_22/i0[10] ), .A2(
        \SB1_3_22/i0_4 ), .A3(\SB1_3_22/i0_3 ), .ZN(
        \SB1_3_22/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 \SB2_3_17/BUF_0  ( .I(\SB1_3_22/buf_output[0] ), .Z(\SB2_3_17/i0[9] )
         );
  NAND2_X2 U6738 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i1[9] ), .ZN(n2081) );
  NAND2_X2 \SB2_0_8/Component_Function_5/N1  ( .A1(\SB2_0_8/i0_0 ), .A2(
        \SB2_0_8/i3[0] ), .ZN(\SB2_0_8/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 \SB2_1_14/BUF_1  ( .I(\SB1_1_18/buf_output[1] ), .Z(
        \SB2_1_14/i0[6] ) );
  CLKBUF_X4 \SB2_4_7/BUF_1  ( .I(\SB1_4_11/buf_output[1] ), .Z(\SB2_4_7/i0[6] ) );
  NAND3_X2 U8066 ( .A1(\SB2_2_1/i0[8] ), .A2(\SB2_2_1/i3[0] ), .A3(
        \SB2_2_1/i1_5 ), .ZN(n2721) );
  NAND3_X2 \SB1_3_26/Component_Function_2/N1  ( .A1(\SB1_3_26/i1_5 ), .A2(
        \SB1_3_26/i0[10] ), .A3(\SB1_3_26/i1[9] ), .ZN(
        \SB1_3_26/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 \SB2_0_18/Component_Function_1/N1  ( .A1(\SB2_0_18/i0_3 ), .A2(
        \SB2_0_18/i1[9] ), .ZN(\SB2_0_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U3908 ( .A1(\SB1_4_19/i3[0] ), .A2(\SB1_4_19/i1_5 ), .A3(
        \SB1_4_19/i0[8] ), .ZN(n1035) );
  NAND3_X2 \SB1_0_1/Component_Function_5/N2  ( .A1(\SB1_0_1/i0_0 ), .A2(
        \SB1_0_1/i0[6] ), .A3(\SB1_0_1/i0[10] ), .ZN(
        \SB1_0_1/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_0_1/BUF_0_0  ( .I(\SB2_0_1/buf_output[0] ), .Z(\RI5[0][18] ) );
  INV_X2 \SB2_0_29/INV_1  ( .I(\SB1_0_1/buf_output[1] ), .ZN(\SB2_0_29/i1_7 )
         );
  INV_X2 \SB1_0_1/INV_1  ( .I(n251), .ZN(\SB1_0_1/i1_7 ) );
  NAND3_X2 U1217 ( .A1(\SB2_0_28/i0[6] ), .A2(\SB2_0_28/i0_4 ), .A3(
        \SB2_0_28/i0[9] ), .ZN(\SB2_0_28/Component_Function_5/NAND4_in[3] ) );
  BUF_X2 U205 ( .I(Key[71]), .Z(n150) );
  BUF_X4 \SB4_16/BUF_1  ( .I(\SB3_20/buf_output[1] ), .Z(\SB4_16/i0[6] ) );
  CLKBUF_X2 U221 ( .I(Key[125]), .Z(n170) );
  NAND3_X2 \SB2_4_16/Component_Function_3/N4  ( .A1(\SB2_4_16/i1_5 ), .A2(
        \SB2_4_16/i0[8] ), .A3(\SB2_4_16/i3[0] ), .ZN(
        \SB2_4_16/Component_Function_3/NAND4_in[3] ) );
  NAND2_X2 \SB1_1_19/Component_Function_5/N1  ( .A1(\SB1_1_19/i0_0 ), .A2(
        \SB1_1_19/i3[0] ), .ZN(\SB1_1_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_9/Component_Function_1/N2  ( .A1(\SB2_3_9/i0_3 ), .A2(
        \SB2_3_9/i1_7 ), .A3(\SB2_3_9/i0[8] ), .ZN(
        \SB2_3_9/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_47_1  ( .I(\MC_ARK_ARC_1_0/buf_output[47] ), .Z(
        \RI1[1][47] ) );
  CLKBUF_X4 U1780 ( .I(\SB1_0_22/buf_output[2] ), .Z(\SB2_0_19/i0_0 ) );
  NAND2_X2 U4098 ( .A1(\SB4_0/i0[9] ), .A2(\SB4_0/i0[10] ), .ZN(n4801) );
  NAND2_X1 U977 ( .A1(\SB1_2_2/Component_Function_4/NAND4_in[3] ), .A2(n2445), 
        .ZN(n2444) );
  NAND2_X1 U2064 ( .A1(\SB1_0_27/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_27/Component_Function_4/NAND4_in[2] ), .ZN(n1470) );
  BUF_X4 U5075 ( .I(\MC_ARK_ARC_1_4/buf_output[6] ), .Z(\SB3_30/i0[9] ) );
  CLKBUF_X8 \SB2_1_27/BUF_5  ( .I(\SB1_1_27/buf_output[5] ), .Z(
        \SB2_1_27/i0_3 ) );
  BUF_X4 \SB2_4_25/BUF_4  ( .I(\SB1_4_26/buf_output[4] ), .Z(\SB2_4_25/i0_4 )
         );
  NAND2_X1 \SB1_2_24/Component_Function_5/N1  ( .A1(\SB1_2_24/i0_0 ), .A2(
        \SB1_2_24/i3[0] ), .ZN(\SB1_2_24/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_4_15/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[99] ), .ZN(
        \SB1_4_15/i0[8] ) );
  BUF_X4 U1755 ( .I(\MC_ARK_ARC_1_1/buf_output[101] ), .Z(\RI1[2][101] ) );
  BUF_X4 U3069 ( .I(\MC_ARK_ARC_1_3/buf_output[75] ), .Z(\SB1_4_19/i0[10] ) );
  BUF_X4 \SB2_3_5/BUF_0_0  ( .I(\SB2_3_5/buf_output[0] ), .Z(\RI5[3][186] ) );
  BUF_X4 U3397 ( .I(\SB1_4_25/buf_output[4] ), .Z(\SB2_4_24/i0_4 ) );
  BUF_X8 \SB2_0_21/BUF_2  ( .I(\RI3[0][62] ), .Z(\SB2_0_21/i0_0 ) );
  CLKBUF_X4 U4745 ( .I(\SB2_4_21/buf_output[1] ), .Z(\RI5[4][85] ) );
  NAND3_X2 U7929 ( .A1(n5444), .A2(\SB2_2_0/i0[8] ), .A3(\SB2_2_0/i1_7 ), .ZN(
        \SB2_2_0/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 \SB1_0_12/BUF_4  ( .I(n356), .Z(\SB1_0_12/i0_4 ) );
  CLKBUF_X4 \SB1_0_9/BUF_4  ( .I(n362), .Z(\SB1_0_9/i0_4 ) );
  CLKBUF_X4 \SB1_0_19/BUF_1  ( .I(n233), .Z(\SB1_0_19/i0[6] ) );
  INV_X1 U326 ( .I(n132), .ZN(n502) );
  CLKBUF_X4 U2082 ( .I(n243), .Z(\SB1_0_9/i0[6] ) );
  BUF_X1 \MC_ARK_ARC_1_1/BUF_148_0  ( .I(n166), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[148] ) );
  INV_X1 U2 ( .I(n4), .ZN(n490) );
  INV_X1 U58 ( .I(n57), .ZN(n426) );
  INV_X1 U322 ( .I(n65), .ZN(n485) );
  INV_X1 U38 ( .I(n16), .ZN(n509) );
  INV_X1 U35 ( .I(n60), .ZN(n483) );
  CLKBUF_X4 U1521 ( .I(n337), .Z(\SB1_0_21/i0[10] ) );
  CLKBUF_X4 \SB1_0_15/BUF_4  ( .I(n350), .Z(\SB1_0_15/i0_4 ) );
  CLKBUF_X4 \SB1_0_1/BUF_1  ( .I(n251), .Z(\SB1_0_1/i0[6] ) );
  CLKBUF_X4 \SB1_0_1/BUF_2  ( .I(n314), .Z(\SB1_0_1/i0_0 ) );
  INV_X1 U29 ( .I(n54), .ZN(n488) );
  INV_X1 U26 ( .I(n34), .ZN(n434) );
  CLKBUF_X4 \SB1_0_16/BUF_1  ( .I(n236), .Z(\SB1_0_16/i0[6] ) );
  INV_X1 U6 ( .I(n73), .ZN(n493) );
  CLKBUF_X4 \SB1_0_2/BUF_3  ( .I(n375), .Z(\SB1_0_2/i0[10] ) );
  CLKBUF_X4 U9358 ( .I(n367), .Z(\SB1_0_6/i0[10] ) );
  CLKBUF_X1 \MC_ARK_ARC_1_3/BUF_132_0  ( .I(n162), .Z(
        \MC_ARK_ARC_1_3/buf_keyinput[132] ) );
  CLKBUF_X4 \SB1_0_4/BUF_3  ( .I(n371), .Z(\SB1_0_4/i0[10] ) );
  CLKBUF_X1 U3995 ( .I(n125), .Z(\MC_ARK_ARC_1_3/buf_keyinput[183] ) );
  INV_X1 U64 ( .I(n31), .ZN(n556) );
  CLKBUF_X4 \SB1_0_19/BUF_3  ( .I(n341), .Z(\SB1_0_19/i0[10] ) );
  CLKBUF_X4 U6752 ( .I(n247), .Z(\SB1_0_5/i0[6] ) );
  CLKBUF_X4 U2096 ( .I(n234), .Z(\SB1_0_18/i0[6] ) );
  CLKBUF_X4 \SB1_0_3/BUF_3  ( .I(n373), .Z(\SB1_0_3/i0[10] ) );
  CLKBUF_X4 \SB1_0_25/BUF_2  ( .I(n266), .Z(\SB1_0_25/i0_0 ) );
  CLKBUF_X4 \SB1_0_30/BUF_4  ( .I(n320), .Z(\SB1_0_30/i0_4 ) );
  INV_X1 U45 ( .I(n2), .ZN(n418) );
  CLKBUF_X4 U2080 ( .I(n252), .Z(\SB1_0_0/i0[6] ) );
  INV_X1 U337 ( .I(n30), .ZN(n544) );
  INV_X1 U293 ( .I(n192), .ZN(n99) );
  CLKBUF_X4 \SB1_0_31/BUF_5  ( .I(n381), .Z(\SB1_0_31/i0_3 ) );
  CLKBUF_X4 \SB1_0_31/BUF_1  ( .I(n221), .Z(\SB1_0_31/i0[6] ) );
  INV_X1 U313 ( .I(n122), .ZN(n414) );
  CLKBUF_X4 \SB1_0_31/BUF_3  ( .I(n317), .Z(\SB1_0_31/i0[10] ) );
  INV_X1 U49 ( .I(n35), .ZN(n444) );
  INV_X1 U4003 ( .I(n117), .ZN(n528) );
  INV_X1 U367 ( .I(n176), .ZN(n479) );
  CLKBUF_X4 \SB1_0_20/BUF_2  ( .I(n276), .Z(\SB1_0_20/i0_0 ) );
  CLKBUF_X4 \SB1_0_24/BUF_3  ( .I(n331), .Z(\SB1_0_24/i0[10] ) );
  CLKBUF_X4 U3193 ( .I(n402), .Z(\SB1_0_10/i0_3 ) );
  INV_X1 U2351 ( .I(n170), .ZN(n467) );
  NAND2_X1 U6468 ( .A1(\SB1_0_11/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_11/Component_Function_4/NAND4_in[2] ), .ZN(n2626) );
  NAND2_X1 U7887 ( .A1(\SB1_0_11/Component_Function_4/NAND4_in[1] ), .A2(n2625), .ZN(n2624) );
  NAND2_X1 U7747 ( .A1(\SB1_0_30/Component_Function_4/NAND4_in[2] ), .A2(n2547), .ZN(n2546) );
  BUF_X4 \SB1_0_9/BUF_4_0  ( .I(\SB1_0_9/buf_output[4] ), .Z(\RI3[0][142] ) );
  CLKBUF_X4 \SB2_0_13/BUF_2  ( .I(\RI3[0][110] ), .Z(\SB2_0_13/i0_0 ) );
  CLKBUF_X4 \SB2_0_25/BUF_2  ( .I(\RI3[0][38] ), .Z(\SB2_0_25/i0_0 ) );
  CLKBUF_X4 \SB2_0_1/BUF_1  ( .I(\SB1_0_5/buf_output[1] ), .Z(\SB2_0_1/i0[6] )
         );
  CLKBUF_X4 U3567 ( .I(\SB1_0_11/buf_output[1] ), .Z(\SB2_0_7/i0[6] ) );
  CLKBUF_X4 \SB2_0_1/BUF_5  ( .I(\SB1_0_1/buf_output[5] ), .Z(\SB2_0_1/i0_3 )
         );
  CLKBUF_X4 U5445 ( .I(\RI3[0][187] ), .Z(\SB2_0_0/i0[6] ) );
  CLKBUF_X4 \SB2_0_21/BUF_3  ( .I(\RI3[0][63] ), .Z(\SB2_0_21/i0[10] ) );
  CLKBUF_X4 \SB2_0_23/BUF_2  ( .I(\RI3[0][50] ), .Z(\SB2_0_23/i0_0 ) );
  CLKBUF_X4 \SB2_0_23/BUF_3  ( .I(\SB1_0_25/buf_output[3] ), .Z(
        \SB2_0_23/i0[10] ) );
  CLKBUF_X4 \SB2_0_15/BUF_1  ( .I(\RI3[0][97] ), .Z(\SB2_0_15/i0[6] ) );
  BUF_X2 \SB1_0_29/BUF_0_0  ( .I(\SB1_0_29/buf_output[0] ), .Z(\RI3[0][42] )
         );
  CLKBUF_X4 \SB1_0_21/BUF_4_0  ( .I(\SB1_0_21/buf_output[4] ), .Z(\RI3[0][70] ) );
  CLKBUF_X4 \SB2_0_28/BUF_5  ( .I(\SB1_0_28/buf_output[5] ), .Z(
        \SB2_0_28/i0_3 ) );
  BUF_X4 \SB2_0_22/BUF_2  ( .I(\RI3[0][56] ), .Z(\SB2_0_22/i0_0 ) );
  CLKBUF_X4 \SB2_0_17/BUF_2  ( .I(\RI3[0][86] ), .Z(\SB2_0_17/i0_0 ) );
  CLKBUF_X4 \SB2_0_30/BUF_1  ( .I(\SB1_0_2/buf_output[1] ), .Z(
        \SB2_0_30/i0[6] ) );
  BUF_X2 U2113 ( .I(\RI3[0][90] ), .Z(\SB2_0_16/i0[9] ) );
  CLKBUF_X4 \SB2_0_30/BUF_4  ( .I(\RI3[0][10] ), .Z(\SB2_0_30/i0_4 ) );
  CLKBUF_X4 \SB1_0_3/BUF_4_0  ( .I(\SB1_0_3/buf_output[4] ), .Z(\RI3[0][178] )
         );
  CLKBUF_X4 \SB2_0_29/BUF_1  ( .I(\SB1_0_1/buf_output[1] ), .Z(
        \SB2_0_29/i0[6] ) );
  BUF_X2 \SB2_0_2/BUF_0  ( .I(\RI3[0][174] ), .Z(\SB2_0_2/i0[9] ) );
  CLKBUF_X4 \SB2_0_3/BUF_3  ( .I(\RI3[0][171] ), .Z(\SB2_0_3/i0[10] ) );
  CLKBUF_X4 \SB2_0_18/BUF_1  ( .I(\SB1_0_22/buf_output[1] ), .Z(
        \SB2_0_18/i0[6] ) );
  CLKBUF_X4 U5342 ( .I(\SB1_0_30/buf_output[2] ), .Z(\SB2_0_27/i0_0 ) );
  CLKBUF_X4 U2119 ( .I(\SB1_0_7/buf_output[3] ), .Z(\SB2_0_5/i0[10] ) );
  CLKBUF_X4 U5250 ( .I(\RI3[0][29] ), .Z(\SB2_0_27/i0_3 ) );
  CLKBUF_X4 U7666 ( .I(\SB2_0_9/i0_0 ), .Z(n2886) );
  CLKBUF_X4 U9776 ( .I(\SB1_0_10/buf_output[0] ), .Z(\SB2_0_5/i0[9] ) );
  INV_X2 \SB2_0_27/INV_0  ( .I(\SB2_0_27/i0[9] ), .ZN(\SB2_0_27/i3[0] ) );
  CLKBUF_X4 \SB2_0_31/BUF_2_0  ( .I(\SB2_0_31/buf_output[2] ), .Z(\RI5[0][20] ) );
  CLKBUF_X4 U3506 ( .I(\SB2_0_2/buf_output[0] ), .Z(\RI5[0][12] ) );
  CLKBUF_X4 \SB2_0_5/BUF_2_0  ( .I(\SB2_0_5/buf_output[2] ), .Z(\RI5[0][176] )
         );
  CLKBUF_X4 \SB2_0_14/BUF_1_0  ( .I(\SB2_0_14/buf_output[1] ), .Z(
        \RI5[0][127] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_0/BUF_84  ( .I(\SB2_0_22/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[84] ) );
  BUF_X4 \SB2_0_10/BUF_0_0  ( .I(\SB2_0_10/buf_output[0] ), .Z(\RI5[0][156] )
         );
  CLKBUF_X4 U3609 ( .I(\SB2_0_7/buf_output[4] ), .Z(\RI5[0][154] ) );
  CLKBUF_X4 \SB2_0_23/BUF_4_0  ( .I(\SB2_0_23/buf_output[4] ), .Z(\RI5[0][58] ) );
  CLKBUF_X4 U3257 ( .I(\SB2_0_14/buf_output[5] ), .Z(\RI5[0][107] ) );
  CLKBUF_X4 \SB2_0_16/BUF_0_0  ( .I(\SB2_0_16/buf_output[0] ), .Z(
        \RI5[0][120] ) );
  CLKBUF_X4 U1881 ( .I(\MC_ARK_ARC_1_0/buf_output[91] ), .Z(\SB1_1_16/i0[6] )
         );
  CLKBUF_X4 U2157 ( .I(\MC_ARK_ARC_1_0/buf_output[178] ), .Z(\SB1_1_2/i0_4 )
         );
  CLKBUF_X4 \SB1_1_28/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[21] ), .Z(
        \SB1_1_28/i0[10] ) );
  CLKBUF_X4 \SB1_1_4/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[164] ), .Z(
        \SB1_1_4/i0_0 ) );
  CLKBUF_X4 \SB1_1_1/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[183] ), .Z(
        \SB1_1_1/i0[10] ) );
  CLKBUF_X4 \SB1_1_25/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[38] ), .Z(
        \SB1_1_25/i0_0 ) );
  CLKBUF_X4 U9747 ( .I(\MC_ARK_ARC_1_0/buf_output[57] ), .Z(\SB1_1_22/i0[10] )
         );
  CLKBUF_X4 \SB1_1_8/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[138] ), .Z(
        \SB1_1_8/i0[9] ) );
  CLKBUF_X4 U3276 ( .I(\MC_ARK_ARC_1_0/buf_output[134] ), .Z(\SB1_1_9/i0_0 )
         );
  CLKBUF_X4 \SB1_1_26/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[33] ), .Z(
        \SB1_1_26/i0[10] ) );
  CLKBUF_X4 \SB1_1_15/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[100] ), .Z(
        \SB1_1_15/i0_4 ) );
  CLKBUF_X4 \SB1_1_6/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[152] ), .Z(
        \SB1_1_6/i0_0 ) );
  CLKBUF_X4 \SB1_1_30/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[6] ), .Z(
        \SB1_1_30/i0[9] ) );
  CLKBUF_X4 U3330 ( .I(\MC_ARK_ARC_1_0/buf_output[105] ), .Z(\SB1_1_14/i0[10] ) );
  CLKBUF_X4 \SB1_1_19/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[76] ), .Z(
        \SB1_1_19/i0_4 ) );
  CLKBUF_X4 U9756 ( .I(\MC_ARK_ARC_1_0/buf_output[147] ), .Z(\SB1_1_7/i0[10] )
         );
  CLKBUF_X4 \SB1_1_12/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[116] ), .Z(
        \SB1_1_12/i0_0 ) );
  CLKBUF_X4 U3612 ( .I(\MC_ARK_ARC_1_0/buf_output[2] ), .Z(\SB1_1_31/i0_0 ) );
  CLKBUF_X4 U9694 ( .I(\MC_ARK_ARC_1_0/buf_output[165] ), .Z(\SB1_1_4/i0[10] )
         );
  CLKBUF_X4 \SB1_1_13/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[111] ), .Z(
        \SB1_1_13/i0[10] ) );
  CLKBUF_X4 \SB1_1_16/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[94] ), .Z(
        \SB1_1_16/i0_4 ) );
  CLKBUF_X4 \SB1_1_0/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[190] ), .Z(
        \SB1_1_0/i0_4 ) );
  CLKBUF_X4 \SB1_1_13/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[109] ), .Z(
        \SB1_1_13/i0[6] ) );
  CLKBUF_X4 \SB1_1_29/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[12] ), .Z(
        \SB1_1_29/i0[9] ) );
  CLKBUF_X4 \SB1_1_18/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[80] ), .Z(
        \SB1_1_18/i0_0 ) );
  CLKBUF_X4 \SB1_1_7/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[146] ), .Z(
        \SB1_1_7/i0_0 ) );
  CLKBUF_X4 \SB1_1_10/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[127] ), .Z(
        \SB1_1_10/i0[6] ) );
  CLKBUF_X4 \SB1_1_21/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[63] ), .Z(
        \SB1_1_21/i0[10] ) );
  CLKBUF_X4 \SB1_1_2/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[174] ), .Z(
        \SB1_1_2/i0[9] ) );
  CLKBUF_X4 \SB1_1_22/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[56] ), .Z(
        \SB1_1_22/i0_0 ) );
  CLKBUF_X4 U3497 ( .I(\MC_ARK_ARC_1_0/buf_output[55] ), .Z(\SB1_1_22/i0[6] )
         );
  CLKBUF_X4 \SB1_1_21/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[64] ), .Z(
        \SB1_1_21/i0_4 ) );
  CLKBUF_X4 U2944 ( .I(\MC_ARK_ARC_1_0/buf_output[58] ), .Z(\SB1_1_22/i0_4 )
         );
  CLKBUF_X4 \SB1_1_22/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[54] ), .Z(
        \SB1_1_22/i0[9] ) );
  CLKBUF_X4 \SB1_1_7/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[148] ), .Z(
        \SB1_1_7/i0_4 ) );
  CLKBUF_X4 \SB1_1_4/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[163] ), .Z(
        \SB1_1_4/i0[6] ) );
  CLKBUF_X4 \SB1_1_24/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[45] ), .Z(
        \SB1_1_24/i0[10] ) );
  CLKBUF_X4 \SB1_1_12/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[117] ), .Z(
        \SB1_1_12/i0[10] ) );
  CLKBUF_X4 \SB1_1_26/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[34] ), .Z(
        \SB1_1_26/i0_4 ) );
  CLKBUF_X4 U3282 ( .I(\MC_ARK_ARC_1_0/buf_output[171] ), .Z(\SB1_1_3/i0[10] )
         );
  CLKBUF_X4 U1712 ( .I(\MC_ARK_ARC_1_0/buf_output[32] ), .Z(\SB1_1_26/i0_0 )
         );
  CLKBUF_X4 U1911 ( .I(\MC_ARK_ARC_1_0/buf_output[104] ), .Z(\SB1_1_14/i0_0 )
         );
  CLKBUF_X4 U3498 ( .I(\MC_ARK_ARC_1_0/buf_output[153] ), .Z(\SB1_1_6/i0[10] )
         );
  CLKBUF_X4 \SB1_1_9/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[132] ), .Z(
        \SB1_1_9/i0[9] ) );
  CLKBUF_X4 \SB1_1_5/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[156] ), .Z(
        \SB1_1_5/i0[9] ) );
  CLKBUF_X4 \SB1_1_1/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[184] ), .Z(
        \SB1_1_1/i0_4 ) );
  CLKBUF_X4 \SB1_1_11/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[123] ), .Z(
        \SB1_1_11/i0[10] ) );
  CLKBUF_X4 U3213 ( .I(\MC_ARK_ARC_1_0/buf_output[172] ), .Z(\SB1_1_3/i0_4 )
         );
  CLKBUF_X4 U9722 ( .I(\MC_ARK_ARC_1_0/buf_output[93] ), .Z(\SB1_1_16/i0[10] )
         );
  CLKBUF_X4 \SB1_1_16/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[92] ), .Z(
        \SB1_1_16/i0_0 ) );
  CLKBUF_X4 \SB1_1_14/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[106] ), .Z(
        \SB1_1_14/i0_4 ) );
  CLKBUF_X4 \SB2_1_9/BUF_0  ( .I(\SB1_1_14/buf_output[0] ), .Z(\SB2_1_9/i0[9] ) );
  CLKBUF_X4 \SB2_1_9/BUF_4  ( .I(\SB1_1_10/buf_output[4] ), .Z(\SB2_1_9/i0_4 )
         );
  CLKBUF_X4 \SB2_1_13/BUF_4  ( .I(\SB1_1_14/buf_output[4] ), .Z(
        \SB2_1_13/i0_4 ) );
  CLKBUF_X4 \SB2_1_9/BUF_2  ( .I(\SB1_1_12/buf_output[2] ), .Z(\SB2_1_9/i0_0 )
         );
  CLKBUF_X4 \SB2_1_7/BUF_2  ( .I(\SB1_1_10/buf_output[2] ), .Z(\SB2_1_7/i0_0 )
         );
  INV_X1 \SB2_1_7/INV_4  ( .I(\SB1_1_8/buf_output[4] ), .ZN(\SB2_1_7/i0[7] )
         );
  CLKBUF_X4 \SB2_1_9/BUF_3  ( .I(\SB1_1_11/buf_output[3] ), .Z(
        \SB2_1_9/i0[10] ) );
  CLKBUF_X4 U3044 ( .I(\SB1_1_13/buf_output[1] ), .Z(\SB2_1_9/i0[6] ) );
  CLKBUF_X4 U3197 ( .I(\SB1_1_18/buf_output[3] ), .Z(\SB2_1_16/i0[10] ) );
  CLKBUF_X4 \SB2_1_25/BUF_4  ( .I(\SB1_1_26/buf_output[4] ), .Z(
        \SB2_1_25/i0_4 ) );
  CLKBUF_X4 \SB2_1_4/BUF_0  ( .I(\SB1_1_9/buf_output[0] ), .Z(\SB2_1_4/i0[9] )
         );
  CLKBUF_X4 U9795 ( .I(\SB1_1_30/buf_output[3] ), .Z(\SB2_1_28/i0[10] ) );
  CLKBUF_X4 U2199 ( .I(\SB1_1_3/buf_output[3] ), .Z(\SB2_1_1/i0[10] ) );
  CLKBUF_X4 U3496 ( .I(\SB1_1_16/buf_output[1] ), .Z(\SB2_1_12/i0[6] ) );
  CLKBUF_X4 \SB2_1_13/BUF_2  ( .I(\SB1_1_16/buf_output[2] ), .Z(
        \SB2_1_13/i0_0 ) );
  CLKBUF_X4 \SB2_1_21/BUF_0  ( .I(\SB1_1_26/buf_output[0] ), .Z(
        \SB2_1_21/i0[9] ) );
  CLKBUF_X4 U4176 ( .I(\SB1_1_1/buf_output[5] ), .Z(\SB2_1_1/i0_3 ) );
  CLKBUF_X4 \SB2_1_7/BUF_3  ( .I(\SB1_1_9/buf_output[3] ), .Z(\SB2_1_7/i0[10] ) );
  CLKBUF_X4 U2195 ( .I(\SB1_1_29/buf_output[5] ), .Z(\SB2_1_29/i0_3 ) );
  CLKBUF_X4 \SB2_1_17/BUF_4  ( .I(\SB1_1_18/buf_output[4] ), .Z(
        \SB2_1_17/i0_4 ) );
  CLKBUF_X4 \SB2_1_24/BUF_0  ( .I(\SB1_1_29/buf_output[0] ), .Z(
        \SB2_1_24/i0[9] ) );
  CLKBUF_X4 \SB2_1_3/BUF_3  ( .I(\SB1_1_5/buf_output[3] ), .Z(\SB2_1_3/i0[10] ) );
  CLKBUF_X4 \SB2_1_3/BUF_4  ( .I(\SB1_1_4/buf_output[4] ), .Z(\SB2_1_3/i0_4 )
         );
  CLKBUF_X4 \SB2_1_23/BUF_2  ( .I(\SB1_1_26/buf_output[2] ), .Z(
        \SB2_1_23/i0_0 ) );
  CLKBUF_X4 \SB2_1_21/BUF_1  ( .I(\SB1_1_25/buf_output[1] ), .Z(
        \SB2_1_21/i0[6] ) );
  CLKBUF_X4 \SB2_1_12/BUF_2  ( .I(\SB1_1_15/buf_output[2] ), .Z(
        \SB2_1_12/i0_0 ) );
  CLKBUF_X4 \SB2_1_28/BUF_2  ( .I(\SB1_1_31/buf_output[2] ), .Z(
        \SB2_1_28/i0_0 ) );
  CLKBUF_X4 U1802 ( .I(\SB1_1_29/buf_output[3] ), .Z(\SB2_1_27/i0[10] ) );
  CLKBUF_X4 \SB2_1_17/BUF_1  ( .I(\SB1_1_21/buf_output[1] ), .Z(
        \SB2_1_17/i0[6] ) );
  CLKBUF_X4 \SB2_1_10/BUF_1  ( .I(\SB1_1_14/buf_output[1] ), .Z(
        \SB2_1_10/i0[6] ) );
  CLKBUF_X4 \SB2_1_21/BUF_2  ( .I(\SB1_1_24/buf_output[2] ), .Z(
        \SB2_1_21/i0_0 ) );
  CLKBUF_X4 \SB2_1_19/BUF_3  ( .I(\SB1_1_21/buf_output[3] ), .Z(
        \SB2_1_19/i0[10] ) );
  CLKBUF_X4 U1793 ( .I(\SB1_1_15/buf_output[0] ), .Z(\SB2_1_10/i0[9] ) );
  CLKBUF_X4 U5450 ( .I(\SB1_1_0/buf_output[2] ), .Z(\SB2_1_29/i0_0 ) );
  CLKBUF_X4 U3679 ( .I(\SB1_1_24/buf_output[1] ), .Z(\SB2_1_20/i0[6] ) );
  CLKBUF_X4 \SB2_1_17/BUF_3  ( .I(\SB1_1_19/buf_output[3] ), .Z(
        \SB2_1_17/i0[10] ) );
  CLKBUF_X4 \SB2_1_3/BUF_2  ( .I(\SB1_1_6/buf_output[2] ), .Z(\SB2_1_3/i0_0 )
         );
  CLKBUF_X4 \SB2_1_17/BUF_0  ( .I(\SB1_1_22/buf_output[0] ), .Z(
        \SB2_1_17/i0[9] ) );
  CLKBUF_X4 \SB2_1_11/BUF_2  ( .I(\SB1_1_14/buf_output[2] ), .Z(
        \SB2_1_11/i0_0 ) );
  CLKBUF_X4 \SB2_1_30/BUF_1  ( .I(\SB1_1_2/buf_output[1] ), .Z(
        \SB2_1_30/i0[6] ) );
  CLKBUF_X4 U2198 ( .I(\SB1_1_23/buf_output[0] ), .Z(\SB2_1_18/i0[9] ) );
  CLKBUF_X4 \SB2_1_26/BUF_1  ( .I(\SB1_1_30/buf_output[1] ), .Z(
        \SB2_1_26/i0[6] ) );
  CLKBUF_X4 \SB2_1_30/BUF_3  ( .I(\SB1_1_0/buf_output[3] ), .Z(
        \SB2_1_30/i0[10] ) );
  BUF_X4 \SB2_1_26/BUF_4  ( .I(\SB1_1_27/buf_output[4] ), .Z(\SB2_1_26/i0_4 )
         );
  CLKBUF_X4 \SB2_1_16/BUF_4  ( .I(\SB1_1_17/buf_output[4] ), .Z(
        \SB2_1_16/i0_4 ) );
  CLKBUF_X4 \SB2_1_18/BUF_2  ( .I(\SB1_1_21/buf_output[2] ), .Z(
        \SB2_1_18/i0_0 ) );
  CLKBUF_X4 \SB2_1_16/BUF_2  ( .I(\SB1_1_19/buf_output[2] ), .Z(
        \SB2_1_16/i0_0 ) );
  CLKBUF_X4 \SB2_1_22/BUF_1  ( .I(\SB1_1_26/buf_output[1] ), .Z(
        \SB2_1_22/i0[6] ) );
  CLKBUF_X4 U5326 ( .I(\SB1_1_8/buf_output[4] ), .Z(\SB2_1_7/i0_4 ) );
  CLKBUF_X4 \SB2_1_6/BUF_1  ( .I(\SB1_1_10/buf_output[1] ), .Z(\SB2_1_6/i0[6] ) );
  CLKBUF_X4 \SB2_1_18/BUF_1  ( .I(\SB1_1_22/buf_output[1] ), .Z(
        \SB2_1_18/i0[6] ) );
  CLKBUF_X4 \SB2_1_6/BUF_0  ( .I(\SB1_1_11/buf_output[0] ), .Z(\SB2_1_6/i0[9] ) );
  CLKBUF_X4 \SB2_1_6/BUF_3  ( .I(\SB1_1_8/buf_output[3] ), .Z(\SB2_1_6/i0[10] ) );
  CLKBUF_X4 \SB2_1_11/BUF_4  ( .I(\SB1_1_12/buf_output[4] ), .Z(
        \SB2_1_11/i0_4 ) );
  CLKBUF_X4 \SB2_1_11/BUF_1  ( .I(\SB1_1_15/buf_output[1] ), .Z(
        \SB2_1_11/i0[6] ) );
  CLKBUF_X4 \SB2_1_11/BUF_3  ( .I(\SB1_1_13/buf_output[3] ), .Z(
        \SB2_1_11/i0[10] ) );
  CLKBUF_X4 \SB2_1_30/BUF_4  ( .I(\SB1_1_31/buf_output[4] ), .Z(
        \SB2_1_30/i0_4 ) );
  CLKBUF_X4 U9790 ( .I(\SB1_1_1/buf_output[2] ), .Z(\SB2_1_30/i0_0 ) );
  CLKBUF_X4 U1773 ( .I(\SB1_1_2/buf_output[2] ), .Z(\SB2_1_31/i0_0 ) );
  CLKBUF_X4 \SB2_1_10/BUF_3  ( .I(\SB1_1_12/buf_output[3] ), .Z(
        \SB2_1_10/i0[10] ) );
  CLKBUF_X4 U2186 ( .I(\SB1_1_1/buf_output[3] ), .Z(\SB2_1_31/i0[10] ) );
  NAND2_X2 \SB2_1_10/Component_Function_0/N1  ( .A1(\SB2_1_10/i0[10] ), .A2(
        \SB2_1_10/i0[9] ), .ZN(\SB2_1_10/Component_Function_0/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_1  ( .I(\SB2_1_3/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[1] ) );
  CLKBUF_X4 U8709 ( .I(\SB2_1_9/buf_output[3] ), .Z(\RI5[1][147] ) );
  CLKBUF_X4 U3202 ( .I(\SB2_1_14/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[122] ) );
  CLKBUF_X4 U8898 ( .I(\SB2_1_1/buf_output[4] ), .Z(\RI5[1][190] ) );
  CLKBUF_X4 U2040 ( .I(\SB2_1_30/buf_output[1] ), .Z(\RI5[1][31] ) );
  CLKBUF_X4 U5667 ( .I(\SB2_1_10/buf_output[4] ), .Z(\RI5[1][136] ) );
  CLKBUF_X4 \SB2_1_22/BUF_3_0  ( .I(\SB2_1_22/buf_output[3] ), .Z(\RI5[1][69] ) );
  CLKBUF_X4 U1367 ( .I(\SB2_1_31/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[15] ) );
  CLKBUF_X4 \SB2_1_22/BUF_4_0  ( .I(\SB2_1_22/buf_output[4] ), .Z(\RI5[1][64] ) );
  CLKBUF_X4 U3493 ( .I(\SB2_1_29/buf_output[5] ), .Z(\RI5[1][17] ) );
  CLKBUF_X4 \SB1_2_17/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[88] ), .Z(
        \SB1_2_17/i0_4 ) );
  CLKBUF_X4 \SB1_2_24/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[43] ), .Z(
        \SB1_2_24/i0[6] ) );
  CLKBUF_X4 U2230 ( .I(\MC_ARK_ARC_1_1/buf_output[112] ), .Z(\SB1_2_13/i0_4 )
         );
  CLKBUF_X4 \SB1_2_0/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[187] ), .Z(
        \SB1_2_0/i0[6] ) );
  CLKBUF_X4 \SB1_2_14/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[104] ), .Z(
        \SB1_2_14/i0_0 ) );
  CLKBUF_X4 U1472 ( .I(\MC_ARK_ARC_1_1/buf_output[105] ), .Z(\SB1_2_14/i0[10] ) );
  CLKBUF_X4 \SB1_2_6/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[154] ), .Z(
        \SB1_2_6/i0_4 ) );
  CLKBUF_X4 \SB1_2_21/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[64] ), .Z(
        \SB1_2_21/i0_4 ) );
  CLKBUF_X4 \SB1_2_6/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[155] ), .Z(
        \SB1_2_6/i0_3 ) );
  CLKBUF_X4 \SB1_2_20/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[69] ), .Z(
        \SB1_2_20/i0[10] ) );
  BUF_X2 \SB1_2_6/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[151] ), .Z(
        \SB1_2_6/i0[6] ) );
  CLKBUF_X4 \SB1_2_28/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[18] ), .Z(
        \SB1_2_28/i0[9] ) );
  CLKBUF_X4 U5456 ( .I(\MC_ARK_ARC_1_1/buf_output[122] ), .Z(\SB1_2_11/i0_0 )
         );
  CLKBUF_X4 \SB1_2_1/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[180] ), .Z(
        \SB1_2_1/i0[9] ) );
  CLKBUF_X4 U9660 ( .I(\MC_ARK_ARC_1_1/buf_output[94] ), .Z(\SB1_2_16/i0_4 )
         );
  CLKBUF_X4 U1036 ( .I(\MC_ARK_ARC_1_1/buf_output[4] ), .Z(\SB1_2_31/i0_4 ) );
  CLKBUF_X4 \SB1_2_16/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[91] ), .Z(
        \SB1_2_16/i0[6] ) );
  CLKBUF_X4 \SB1_2_22/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[58] ), .Z(
        \SB1_2_22/i0_4 ) );
  CLKBUF_X4 \SB1_2_10/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[129] ), .Z(
        \SB1_2_10/i0[10] ) );
  CLKBUF_X4 \SB1_2_3/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[171] ), .Z(
        \SB1_2_3/i0[10] ) );
  CLKBUF_X4 \SB1_2_27/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[24] ), .Z(
        \SB1_2_27/i0[9] ) );
  CLKBUF_X4 \SB1_2_3/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[169] ), .Z(
        \SB1_2_3/i0[6] ) );
  CLKBUF_X4 \SB1_2_9/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[135] ), .Z(
        \SB1_2_9/i0[10] ) );
  CLKBUF_X4 \SB1_2_5/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[160] ), .Z(
        \SB1_2_5/i0_4 ) );
  CLKBUF_X4 U1804 ( .I(\MC_ARK_ARC_1_1/buf_output[7] ), .Z(\SB1_2_30/i0[6] )
         );
  CLKBUF_X4 U5455 ( .I(\MC_ARK_ARC_1_1/buf_output[99] ), .Z(\SB1_2_15/i0[10] )
         );
  CLKBUF_X4 \SB1_2_14/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[103] ), .Z(
        \SB1_2_14/i0[6] ) );
  INV_X1 \SB1_2_23/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[48] ), .ZN(
        \SB1_2_23/i3[0] ) );
  CLKBUF_X4 \SB1_2_8/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[139] ), .Z(
        \SB1_2_8/i0[6] ) );
  CLKBUF_X4 \SB1_2_18/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[80] ), .Z(
        \SB1_2_18/i0_0 ) );
  CLKBUF_X4 \SB1_2_18/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[82] ), .Z(
        \SB1_2_18/i0_4 ) );
  CLKBUF_X4 \SB1_2_2/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[177] ), .Z(
        \SB1_2_2/i0[10] ) );
  CLKBUF_X4 \SB1_2_15/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[98] ), .Z(
        \SB1_2_15/i0_0 ) );
  CLKBUF_X4 U5458 ( .I(\MC_ARK_ARC_1_1/buf_output[38] ), .Z(\SB1_2_25/i0_0 )
         );
  CLKBUF_X4 U9805 ( .I(\MC_ARK_ARC_1_1/buf_output[8] ), .Z(\SB1_2_30/i0_0 ) );
  CLKBUF_X4 \SB1_2_0/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[186] ), .Z(
        \SB1_2_0/i0[9] ) );
  CLKBUF_X4 \SB1_2_5/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[156] ), .Z(
        \SB1_2_5/i0[9] ) );
  BUF_X2 \SB1_2_10/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[126] ), .Z(
        \SB1_2_10/i0[9] ) );
  CLKBUF_X4 \SB1_2_20/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[70] ), .Z(
        \SB1_2_20/i0_4 ) );
  CLKBUF_X4 U2243 ( .I(\MC_ARK_ARC_1_1/buf_output[84] ), .Z(\SB1_2_17/i0[9] )
         );
  OR3_X1 U9798 ( .A1(\SB1_2_11/i0_3 ), .A2(\SB1_2_11/i0[10] ), .A3(
        \MC_ARK_ARC_1_1/buf_output[120] ), .Z(n5189) );
  NAND3_X2 \SB1_2_6/Component_Function_2/N3  ( .A1(\SB1_2_6/i0_3 ), .A2(
        \SB1_2_6/i0[8] ), .A3(\SB1_2_6/i0[9] ), .ZN(
        \SB1_2_6/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 \SB2_2_19/BUF_1  ( .I(\SB1_2_23/buf_output[1] ), .Z(\SB2_2_19/i0[6] )
         );
  CLKBUF_X4 \SB2_2_25/BUF_2  ( .I(\SB1_2_28/buf_output[2] ), .Z(
        \SB2_2_25/i0_0 ) );
  CLKBUF_X4 \SB2_2_23/BUF_1  ( .I(\SB1_2_27/buf_output[1] ), .Z(
        \SB2_2_23/i0[6] ) );
  CLKBUF_X4 U5106 ( .I(\SB1_2_28/buf_output[3] ), .Z(\SB2_2_26/i0[10] ) );
  CLKBUF_X4 \SB2_2_12/BUF_1  ( .I(\SB1_2_16/buf_output[1] ), .Z(
        \SB2_2_12/i0[6] ) );
  CLKBUF_X4 \SB2_2_14/BUF_1  ( .I(\SB1_2_18/buf_output[1] ), .Z(
        \SB2_2_14/i0[6] ) );
  CLKBUF_X4 \SB2_2_16/BUF_3  ( .I(\SB1_2_18/buf_output[3] ), .Z(
        \SB2_2_16/i0[10] ) );
  BUF_X4 \SB2_2_2/BUF_4  ( .I(\SB1_2_3/buf_output[4] ), .Z(\SB2_2_2/i0_4 ) );
  CLKBUF_X4 U5411 ( .I(\SB1_2_11/buf_output[3] ), .Z(\SB2_2_9/i0[10] ) );
  CLKBUF_X4 \SB2_2_14/BUF_3  ( .I(\SB1_2_16/buf_output[3] ), .Z(
        \SB2_2_14/i0[10] ) );
  CLKBUF_X4 \SB2_2_14/BUF_0  ( .I(\SB1_2_19/buf_output[0] ), .Z(
        \SB2_2_14/i0[9] ) );
  CLKBUF_X4 U2276 ( .I(\SB1_2_23/buf_output[4] ), .Z(\SB2_2_22/i0_4 ) );
  CLKBUF_X4 \SB2_2_28/BUF_2  ( .I(\SB1_2_31/buf_output[2] ), .Z(
        \SB2_2_28/i0_0 ) );
  CLKBUF_X4 \SB2_2_22/BUF_0  ( .I(\SB1_2_27/buf_output[0] ), .Z(
        \SB2_2_22/i0[9] ) );
  CLKBUF_X4 U3470 ( .I(\SB1_2_3/buf_output[2] ), .Z(\SB2_2_0/i0_0 ) );
  CLKBUF_X4 U5237 ( .I(\SB1_2_8/buf_output[2] ), .Z(\SB2_2_5/i0_0 ) );
  CLKBUF_X4 \SB2_2_0/BUF_1  ( .I(\SB1_2_4/buf_output[1] ), .Z(\SB2_2_0/i0[6] )
         );
  CLKBUF_X4 U2255 ( .I(\SB1_2_12/buf_output[0] ), .Z(\SB2_2_7/i0[9] ) );
  CLKBUF_X4 \SB2_2_13/BUF_4  ( .I(\SB1_2_14/buf_output[4] ), .Z(
        \SB2_2_13/i0_4 ) );
  CLKBUF_X4 \SB2_2_13/BUF_1  ( .I(\SB1_2_17/buf_output[1] ), .Z(
        \SB2_2_13/i0[6] ) );
  CLKBUF_X4 \SB2_2_13/BUF_0  ( .I(\SB1_2_18/buf_output[0] ), .Z(
        \SB2_2_13/i0[9] ) );
  CLKBUF_X4 \SB2_2_5/BUF_0  ( .I(\SB1_2_10/buf_output[0] ), .Z(\SB2_2_5/i0[9] ) );
  CLKBUF_X4 U2818 ( .I(\SB1_2_26/buf_output[3] ), .Z(\SB2_2_24/i0[10] ) );
  CLKBUF_X4 \SB2_2_16/BUF_4  ( .I(\SB1_2_17/buf_output[4] ), .Z(
        \SB2_2_16/i0_4 ) );
  CLKBUF_X4 U2250 ( .I(\SB1_2_20/buf_output[0] ), .Z(\SB2_2_15/i0[9] ) );
  CLKBUF_X4 \SB2_2_25/BUF_4  ( .I(\SB1_2_26/buf_output[4] ), .Z(
        \SB2_2_25/i0_4 ) );
  CLKBUF_X4 \SB2_2_19/BUF_4  ( .I(\SB1_2_20/buf_output[4] ), .Z(
        \SB2_2_19/i0_4 ) );
  CLKBUF_X4 \SB2_2_24/BUF_4  ( .I(\SB1_2_25/buf_output[4] ), .Z(
        \SB2_2_24/i0_4 ) );
  INV_X2 \SB2_2_27/INV_4  ( .I(\SB2_2_27/i0_4 ), .ZN(\SB2_2_27/i0[7] ) );
  CLKBUF_X4 U2251 ( .I(\SB1_2_26/buf_output[2] ), .Z(\SB2_2_23/i0_0 ) );
  CLKBUF_X4 \SB2_2_5/BUF_3  ( .I(\SB1_2_7/buf_output[3] ), .Z(\SB2_2_5/i0[10] ) );
  CLKBUF_X4 U9752 ( .I(\SB1_2_9/buf_output[1] ), .Z(\SB2_2_5/i0[6] ) );
  CLKBUF_X4 \SB2_2_23/BUF_3  ( .I(\SB1_2_25/buf_output[3] ), .Z(
        \SB2_2_23/i0[10] ) );
  CLKBUF_X4 \SB2_2_0/BUF_3  ( .I(\SB1_2_2/buf_output[3] ), .Z(\SB2_2_0/i0[10] ) );
  CLKBUF_X4 \SB2_2_17/BUF_1  ( .I(\SB1_2_21/buf_output[1] ), .Z(
        \SB2_2_17/i0[6] ) );
  CLKBUF_X4 \SB2_2_20/BUF_0  ( .I(\SB1_2_25/buf_output[0] ), .Z(
        \SB2_2_20/i0[9] ) );
  CLKBUF_X4 \SB2_2_8/BUF_4  ( .I(\SB1_2_9/buf_output[4] ), .Z(\SB2_2_8/i0_4 )
         );
  CLKBUF_X4 \SB2_2_1/BUF_3  ( .I(\SB1_2_3/buf_output[3] ), .Z(\SB2_2_1/i0[10] ) );
  CLKBUF_X4 \SB2_2_2/BUF_3  ( .I(\SB1_2_4/buf_output[3] ), .Z(\SB2_2_2/i0[10] ) );
  CLKBUF_X4 \SB2_2_3/BUF_2  ( .I(\SB1_2_6/buf_output[2] ), .Z(\SB2_2_3/i0_0 )
         );
  CLKBUF_X4 \SB2_2_2/BUF_1  ( .I(\SB1_2_6/buf_output[1] ), .Z(\SB2_2_2/i0[6] )
         );
  CLKBUF_X4 \SB2_2_6/BUF_4  ( .I(\SB1_2_7/buf_output[4] ), .Z(\SB2_2_6/i0_4 )
         );
  CLKBUF_X4 \SB2_2_31/BUF_0  ( .I(\SB1_2_4/buf_output[0] ), .Z(
        \SB2_2_31/i0[9] ) );
  CLKBUF_X4 \SB2_2_21/BUF_1  ( .I(\SB1_2_25/buf_output[1] ), .Z(
        \SB2_2_21/i0[6] ) );
  CLKBUF_X4 \SB2_2_12/BUF_3  ( .I(\SB1_2_14/buf_output[3] ), .Z(
        \SB2_2_12/i0[10] ) );
  CLKBUF_X4 \SB2_2_10/BUF_3  ( .I(\SB1_2_12/buf_output[3] ), .Z(
        \SB2_2_10/i0[10] ) );
  CLKBUF_X4 \SB2_2_27/BUF_3  ( .I(\SB1_2_29/buf_output[3] ), .Z(
        \SB2_2_27/i0[10] ) );
  CLKBUF_X4 \SB2_2_26/BUF_2  ( .I(\SB1_2_29/buf_output[2] ), .Z(
        \SB2_2_26/i0_0 ) );
  CLKBUF_X4 \SB2_2_28/BUF_1  ( .I(\SB1_2_0/buf_output[1] ), .Z(
        \SB2_2_28/i0[6] ) );
  CLKBUF_X4 \SB2_2_25/BUF_1  ( .I(\SB1_2_29/buf_output[1] ), .Z(
        \SB2_2_25/i0[6] ) );
  CLKBUF_X4 \SB2_2_8/BUF_1  ( .I(\SB1_2_12/buf_output[1] ), .Z(\SB2_2_8/i0[6] ) );
  CLKBUF_X4 U3772 ( .I(\SB2_2_13/buf_output[0] ), .Z(\RI5[2][138] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_2/BUF_183  ( .I(\SB2_2_3/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[183] ) );
  CLKBUF_X4 U4414 ( .I(\SB2_2_22/buf_output[3] ), .Z(\RI5[2][69] ) );
  CLKBUF_X4 U2019 ( .I(\SB2_2_3/buf_output[0] ), .Z(\RI5[2][6] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_2/BUF_84  ( .I(\SB2_2_22/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[84] ) );
  CLKBUF_X4 U2012 ( .I(\SB2_2_5/buf_output[2] ), .Z(\RI5[2][176] ) );
  CLKBUF_X4 U3465 ( .I(\SB2_2_22/buf_output[4] ), .Z(\RI5[2][64] ) );
  CLKBUF_X4 U3130 ( .I(\SB2_2_14/buf_output[3] ), .Z(\RI5[2][117] ) );
  CLKBUF_X4 U9021 ( .I(\SB2_2_14/buf_output[1] ), .Z(\RI5[2][127] ) );
  CLKBUF_X4 \SB2_2_31/BUF_0_0  ( .I(\SB2_2_31/buf_output[0] ), .Z(\RI5[2][30] ) );
  CLKBUF_X4 U3131 ( .I(\SB2_2_10/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[141] ) );
  CLKBUF_X4 U9598 ( .I(\SB2_2_18/buf_output[3] ), .Z(\RI5[2][93] ) );
  CLKBUF_X4 U3455 ( .I(\SB2_2_11/buf_output[5] ), .Z(\RI5[2][125] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_2/BUF_25  ( .I(\SB2_2_31/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[25] ) );
  CLKBUF_X4 U2290 ( .I(\MC_ARK_ARC_1_2/buf_output[52] ), .Z(\SB1_3_23/i0_4 )
         );
  CLKBUF_X4 U5242 ( .I(\MC_ARK_ARC_1_2/buf_output[103] ), .Z(\SB1_3_14/i0[6] )
         );
  CLKBUF_X4 U2284 ( .I(\MC_ARK_ARC_1_2/buf_output[150] ), .Z(\SB1_3_6/i0[9] )
         );
  CLKBUF_X4 \SB1_3_5/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[157] ), .Z(
        \SB1_3_5/i0[6] ) );
  CLKBUF_X4 \SB1_3_2/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[174] ), .Z(
        \SB1_3_2/i0[9] ) );
  CLKBUF_X4 \SB1_3_28/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[21] ), .Z(
        \SB1_3_28/i0[10] ) );
  CLKBUF_X4 \SB1_3_29/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[12] ), .Z(
        \SB1_3_29/i0[9] ) );
  CLKBUF_X4 \SB1_3_19/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[74] ), .Z(
        \SB1_3_19/i0_0 ) );
  CLKBUF_X4 \SB1_3_1/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[180] ), .Z(
        \SB1_3_1/i0[9] ) );
  CLKBUF_X4 U2288 ( .I(\MC_ARK_ARC_1_2/buf_output[1] ), .Z(\SB1_3_31/i0[6] )
         );
  CLKBUF_X4 \SB1_3_22/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[58] ), .Z(
        \SB1_3_22/i0_4 ) );
  CLKBUF_X4 \SB1_3_7/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[147] ), .Z(
        \SB1_3_7/i0[10] ) );
  CLKBUF_X4 \SB1_3_24/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[46] ), .Z(
        \SB1_3_24/i0_4 ) );
  CLKBUF_X4 \SB1_3_21/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[62] ), .Z(
        \SB1_3_21/i0_0 ) );
  CLKBUF_X4 \SB1_3_31/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[0] ), .Z(
        \SB1_3_31/i0[9] ) );
  CLKBUF_X4 U1759 ( .I(\MC_ARK_ARC_1_2/buf_output[60] ), .Z(\SB1_3_21/i0[9] )
         );
  CLKBUF_X4 \SB1_3_13/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[108] ), .Z(
        \SB1_3_13/i0[9] ) );
  CLKBUF_X4 U3777 ( .I(\MC_ARK_ARC_1_2/buf_output[36] ), .Z(\SB1_3_25/i0[9] )
         );
  CLKBUF_X4 U2523 ( .I(\MC_ARK_ARC_1_2/buf_output[32] ), .Z(\SB1_3_26/i0_0 )
         );
  CLKBUF_X4 \SB1_3_25/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[38] ), .Z(
        \SB1_3_25/i0_0 ) );
  CLKBUF_X4 U1515 ( .I(\MC_ARK_ARC_1_2/buf_output[177] ), .Z(\SB1_3_2/i0[10] )
         );
  CLKBUF_X4 \SB1_3_11/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[122] ), .Z(
        \SB1_3_11/i0_0 ) );
  CLKBUF_X4 \SB1_3_11/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[123] ), .Z(
        \SB1_3_11/i0[10] ) );
  CLKBUF_X4 \SB1_3_23/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[51] ), .Z(
        \SB1_3_23/i0[10] ) );
  CLKBUF_X4 \SB1_3_5/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[158] ), .Z(
        \SB1_3_5/i0_0 ) );
  CLKBUF_X4 \SB1_3_0/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[188] ), .Z(
        \SB1_3_0/i0_0 ) );
  CLKBUF_X4 \SB1_3_4/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[162] ), .Z(
        \SB1_3_4/i0[9] ) );
  CLKBUF_X4 \SB1_3_4/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[163] ), .Z(
        \SB1_3_4/i0[6] ) );
  CLKBUF_X4 \SB1_3_0/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[189] ), .Z(
        \SB1_3_0/i0[10] ) );
  CLKBUF_X4 \SB1_3_30/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[6] ), .Z(
        \SB1_3_30/i0[9] ) );
  CLKBUF_X4 \SB1_3_9/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[136] ), .Z(
        \SB1_3_9/i0_4 ) );
  CLKBUF_X4 \SB1_3_26/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[31] ), .Z(
        \SB1_3_26/i0[6] ) );
  CLKBUF_X4 U2289 ( .I(\MC_ARK_ARC_1_2/buf_output[26] ), .Z(\SB1_3_27/i0_0 )
         );
  CLKBUF_X4 U1368 ( .I(\MC_ARK_ARC_1_2/buf_output[115] ), .Z(\SB1_3_12/i0[6] )
         );
  CLKBUF_X4 \SB1_3_24/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[44] ), .Z(
        \SB1_3_24/i0_0 ) );
  CLKBUF_X4 \SB1_3_25/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[39] ), .Z(
        \SB1_3_25/i0[10] ) );
  CLKBUF_X4 \SB1_3_19/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[75] ), .Z(
        \SB1_3_19/i0[10] ) );
  CLKBUF_X4 \SB1_3_20/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[70] ), .Z(
        \SB1_3_20/i0_4 ) );
  CLKBUF_X4 U2585 ( .I(\MC_ARK_ARC_1_2/buf_output[175] ), .Z(\SB1_3_2/i0[6] )
         );
  CLKBUF_X4 U9583 ( .I(\MC_ARK_ARC_1_2/buf_output[110] ), .Z(\SB1_3_13/i0_0 )
         );
  CLKBUF_X4 \SB2_3_23/BUF_2  ( .I(\SB1_3_26/buf_output[2] ), .Z(
        \SB2_3_23/i0_0 ) );
  NAND2_X1 U10964 ( .A1(\SB1_3_22/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_3_22/Component_Function_4/NAND4_in[0] ), .ZN(n5345) );
  CLKBUF_X4 \SB2_3_3/BUF_1  ( .I(\SB1_3_7/buf_output[1] ), .Z(\SB2_3_3/i0[6] )
         );
  CLKBUF_X4 \SB2_3_1/BUF_3  ( .I(\SB1_3_3/buf_output[3] ), .Z(\SB2_3_1/i0[10] ) );
  CLKBUF_X4 \SB2_3_13/BUF_3  ( .I(\SB1_3_15/buf_output[3] ), .Z(
        \SB2_3_13/i0[10] ) );
  CLKBUF_X4 \SB2_3_6/BUF_3  ( .I(\SB1_3_8/buf_output[3] ), .Z(\SB2_3_6/i0[10] ) );
  CLKBUF_X4 \SB2_3_6/BUF_0  ( .I(\SB1_3_11/buf_output[0] ), .Z(\SB2_3_6/i0[9] ) );
  CLKBUF_X4 \SB2_3_4/BUF_3  ( .I(\SB1_3_6/buf_output[3] ), .Z(\SB2_3_4/i0[10] ) );
  CLKBUF_X4 U3845 ( .I(\SB1_3_28/buf_output[2] ), .Z(\SB2_3_25/i0_0 ) );
  CLKBUF_X4 U9782 ( .I(\SB1_3_21/buf_output[3] ), .Z(\SB2_3_19/i0[10] ) );
  CLKBUF_X4 \SB2_3_19/BUF_2  ( .I(\SB1_3_22/buf_output[2] ), .Z(
        \SB2_3_19/i0_0 ) );
  CLKBUF_X4 U2001 ( .I(\SB1_3_17/buf_output[3] ), .Z(\SB2_3_15/i0[10] ) );
  CLKBUF_X4 \SB2_3_31/BUF_4  ( .I(\SB1_3_0/buf_output[4] ), .Z(\SB2_3_31/i0_4 ) );
  CLKBUF_X4 U3914 ( .I(\SB1_3_2/buf_output[2] ), .Z(\SB2_3_31/i0_0 ) );
  CLKBUF_X4 \SB2_3_23/BUF_0  ( .I(\SB1_3_28/buf_output[0] ), .Z(
        \SB2_3_23/i0[9] ) );
  CLKBUF_X4 \SB2_3_13/BUF_2  ( .I(\SB1_3_16/buf_output[2] ), .Z(
        \SB2_3_13/i0_0 ) );
  CLKBUF_X4 \SB2_3_4/BUF_1  ( .I(\SB1_3_8/buf_output[1] ), .Z(\SB2_3_4/i0[6] )
         );
  CLKBUF_X4 U6175 ( .I(\SB1_3_23/buf_output[1] ), .Z(\SB2_3_19/i0[6] ) );
  CLKBUF_X4 \SB2_3_3/BUF_2  ( .I(\SB1_3_6/buf_output[2] ), .Z(\SB2_3_3/i0_0 )
         );
  CLKBUF_X4 \SB2_3_23/BUF_4  ( .I(\SB1_3_24/buf_output[4] ), .Z(
        \SB2_3_23/i0_4 ) );
  CLKBUF_X4 \SB2_3_14/BUF_1  ( .I(\SB1_3_18/buf_output[1] ), .Z(
        \SB2_3_14/i0[6] ) );
  CLKBUF_X4 \SB2_3_23/BUF_3  ( .I(\SB1_3_25/buf_output[3] ), .Z(
        \SB2_3_23/i0[10] ) );
  CLKBUF_X4 U2768 ( .I(\SB1_3_15/buf_output[2] ), .Z(\SB2_3_12/i0_0 ) );
  CLKBUF_X4 U3442 ( .I(\SB1_3_0/buf_output[3] ), .Z(\SB2_3_30/i0[10] ) );
  CLKBUF_X4 \SB2_3_23/BUF_1  ( .I(\SB1_3_27/buf_output[1] ), .Z(
        \SB2_3_23/i0[6] ) );
  CLKBUF_X4 \SB2_3_30/BUF_5  ( .I(\SB1_3_30/buf_output[5] ), .Z(
        \SB2_3_30/i0_3 ) );
  CLKBUF_X4 \SB2_3_16/BUF_1  ( .I(\SB1_3_20/buf_output[1] ), .Z(
        \SB2_3_16/i0[6] ) );
  CLKBUF_X4 \SB2_3_26/BUF_5  ( .I(\SB1_3_26/buf_output[5] ), .Z(
        \SB2_3_26/i0_3 ) );
  CLKBUF_X4 U1124 ( .I(\SB1_3_2/buf_output[1] ), .Z(\SB2_3_30/i0[6] ) );
  CLKBUF_X4 U2002 ( .I(\SB1_3_3/buf_output[2] ), .Z(\SB2_3_0/i0_0 ) );
  CLKBUF_X4 \SB2_3_16/BUF_3  ( .I(\SB1_3_18/buf_output[3] ), .Z(
        \SB2_3_16/i0[10] ) );
  CLKBUF_X4 U3848 ( .I(\SB1_3_29/buf_output[3] ), .Z(\SB2_3_27/i0[10] ) );
  CLKBUF_X4 \SB2_3_14/BUF_3  ( .I(\SB1_3_16/buf_output[3] ), .Z(
        \SB2_3_14/i0[10] ) );
  CLKBUF_X4 U5207 ( .I(\SB1_3_31/buf_output[0] ), .Z(\SB2_3_26/i0[9] ) );
  CLKBUF_X4 U2386 ( .I(\SB1_3_31/buf_output[1] ), .Z(\SB2_3_27/i0[6] ) );
  CLKBUF_X4 \SB2_3_8/BUF_0  ( .I(\SB1_3_13/buf_output[0] ), .Z(\SB2_3_8/i0[9] ) );
  CLKBUF_X4 U4218 ( .I(\SB1_3_28/buf_output[3] ), .Z(\SB2_3_26/i0[10] ) );
  CLKBUF_X4 U1128 ( .I(\SB1_3_15/buf_output[1] ), .Z(\SB2_3_11/i0[6] ) );
  CLKBUF_X4 U1132 ( .I(\SB1_3_17/buf_output[0] ), .Z(\SB2_3_12/i0[9] ) );
  CLKBUF_X4 \SB2_3_26/BUF_1  ( .I(\SB1_3_30/buf_output[1] ), .Z(
        \SB2_3_26/i0[6] ) );
  CLKBUF_X4 \SB2_3_24/BUF_3  ( .I(\SB1_3_26/buf_output[3] ), .Z(
        \SB2_3_24/i0[10] ) );
  CLKBUF_X4 \SB2_3_2/BUF_4  ( .I(\SB1_3_3/buf_output[4] ), .Z(\SB2_3_2/i0_4 )
         );
  CLKBUF_X4 U1129 ( .I(\SB1_3_15/buf_output[0] ), .Z(\SB2_3_10/i0[9] ) );
  CLKBUF_X4 \SB2_3_5/BUF_3  ( .I(\SB1_3_7/buf_output[3] ), .Z(\SB2_3_5/i0[10] ) );
  CLKBUF_X4 U9381 ( .I(\SB1_3_30/buf_output[3] ), .Z(\SB2_3_28/i0[10] ) );
  CLKBUF_X4 U3440 ( .I(\SB1_3_10/buf_output[1] ), .Z(\SB2_3_6/i0[6] ) );
  CLKBUF_X4 \SB2_3_24/BUF_0  ( .I(\SB1_3_29/buf_output[0] ), .Z(
        \SB2_3_24/i0[9] ) );
  CLKBUF_X4 U5038 ( .I(\SB1_3_31/buf_output[2] ), .Z(\SB2_3_28/i0_0 ) );
  CLKBUF_X4 \SB2_3_27/BUF_4  ( .I(\SB1_3_28/buf_output[4] ), .Z(
        \SB2_3_27/i0_4 ) );
  CLKBUF_X4 \SB2_3_10/BUF_2  ( .I(\SB1_3_13/buf_output[2] ), .Z(
        \SB2_3_10/i0_0 ) );
  CLKBUF_X4 \SB2_3_29/BUF_2  ( .I(\SB1_3_0/buf_output[2] ), .Z(\SB2_3_29/i0_0 ) );
  CLKBUF_X4 \SB2_3_19/BUF_0  ( .I(\SB1_3_24/buf_output[0] ), .Z(
        \SB2_3_19/i0[9] ) );
  CLKBUF_X4 U3849 ( .I(\SB1_3_4/buf_output[3] ), .Z(\SB2_3_2/i0[10] ) );
  CLKBUF_X4 \SB2_3_12/BUF_3  ( .I(\SB1_3_14/buf_output[3] ), .Z(
        \SB2_3_12/i0[10] ) );
  CLKBUF_X4 \SB2_3_1/BUF_2  ( .I(\SB1_3_4/buf_output[2] ), .Z(\SB2_3_1/i0_0 )
         );
  CLKBUF_X4 U4736 ( .I(\SB2_3_29/buf_output[3] ), .Z(\RI5[3][27] ) );
  CLKBUF_X4 \SB2_3_31/BUF_4_0  ( .I(\SB2_3_31/buf_output[4] ), .Z(\RI5[3][10] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_3/BUF_49  ( .I(\SB2_3_27/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[49] ) );
  CLKBUF_X4 U2350 ( .I(\SB2_3_10/buf_output[4] ), .Z(\RI5[3][136] ) );
  CLKBUF_X4 U8828 ( .I(\SB2_3_21/buf_output[1] ), .Z(\RI5[3][85] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_3/BUF_46  ( .I(\SB2_3_25/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[46] ) );
  CLKBUF_X4 \SB2_3_22/BUF_4_0  ( .I(\SB2_3_22/buf_output[4] ), .Z(\RI5[3][64] ) );
  CLKBUF_X4 U3199 ( .I(\SB2_3_4/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[177] ) );
  CLKBUF_X4 \SB2_3_20/BUF_4_0  ( .I(\SB2_3_20/buf_output[4] ), .Z(\RI5[3][76] ) );
  BUF_X4 U6241 ( .I(\SB2_3_11/buf_output[1] ), .Z(\RI5[3][145] ) );
  CLKBUF_X4 U6225 ( .I(\SB2_3_19/buf_output[1] ), .Z(\RI5[3][97] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_3/BUF_43  ( .I(\SB2_3_28/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[43] ) );
  CLKBUF_X4 U1990 ( .I(\SB2_3_3/buf_output[0] ), .Z(\RI5[3][6] ) );
  CLKBUF_X4 U9423 ( .I(\MC_ARK_ARC_1_3/buf_output[99] ), .Z(\SB1_4_15/i0[10] )
         );
  CLKBUF_X4 \SB1_4_12/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[117] ), .Z(
        \SB1_4_12/i0[10] ) );
  CLKBUF_X4 U2363 ( .I(\MC_ARK_ARC_1_3/buf_output[68] ), .Z(\SB1_4_20/i0_0 )
         );
  CLKBUF_X4 \SB1_4_5/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[159] ), .Z(
        \SB1_4_5/i0[10] ) );
  CLKBUF_X4 U1986 ( .I(\MC_ARK_ARC_1_3/buf_output[69] ), .Z(\SB1_4_20/i0[10] )
         );
  CLKBUF_X4 U3020 ( .I(\MC_ARK_ARC_1_3/buf_output[45] ), .Z(\SB1_4_24/i0[10] )
         );
  CLKBUF_X4 \SB1_4_0/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[186] ), .Z(
        \SB1_4_0/i0[9] ) );
  CLKBUF_X4 U4567 ( .I(\MC_ARK_ARC_1_3/buf_output[46] ), .Z(\SB1_4_24/i0_4 )
         );
  CLKBUF_X4 \SB1_4_18/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[79] ), .Z(
        \SB1_4_18/i0[6] ) );
  CLKBUF_X4 \SB1_4_27/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[28] ), .Z(
        \SB1_4_27/i0_4 ) );
  CLKBUF_X4 \SB1_4_2/BUF_2  ( .I(\MC_ARK_ARC_1_3/buf_output[176] ), .Z(
        \SB1_4_2/i0_0 ) );
  CLKBUF_X4 U3424 ( .I(\MC_ARK_ARC_1_3/buf_output[86] ), .Z(\SB1_4_17/i0_0 )
         );
  CLKBUF_X4 U9687 ( .I(\MC_ARK_ARC_1_3/buf_output[25] ), .Z(\SB1_4_27/i0[6] )
         );
  CLKBUF_X4 \SB1_4_1/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[180] ), .Z(
        \SB1_4_1/i0[9] ) );
  CLKBUF_X4 \SB1_4_31/BUF_2  ( .I(\MC_ARK_ARC_1_3/buf_output[2] ), .Z(
        \SB1_4_31/i0_0 ) );
  CLKBUF_X4 \SB1_4_31/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[4] ), .Z(
        \SB1_4_31/i0_4 ) );
  CLKBUF_X4 \SB1_4_11/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[120] ), .Z(
        \SB1_4_11/i0[9] ) );
  CLKBUF_X4 U8571 ( .I(\MC_ARK_ARC_1_3/buf_output[95] ), .Z(\SB1_4_16/i0_3 )
         );
  CLKBUF_X4 U8404 ( .I(\MC_ARK_ARC_1_3/buf_output[166] ), .Z(\SB1_4_4/i0_4 )
         );
  CLKBUF_X4 U783 ( .I(\MC_ARK_ARC_1_3/buf_output[37] ), .Z(\SB1_4_25/i0[6] )
         );
  CLKBUF_X4 U2358 ( .I(\MC_ARK_ARC_1_3/buf_output[115] ), .Z(\SB1_4_12/i0[6] )
         );
  CLKBUF_X4 \SB1_4_2/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[174] ), .Z(
        \SB1_4_2/i0[9] ) );
  CLKBUF_X4 U1345 ( .I(\MC_ARK_ARC_1_3/buf_output[147] ), .Z(\SB1_4_7/i0[10] )
         );
  CLKBUF_X4 \SB1_4_21/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[64] ), .Z(
        \SB1_4_21/i0_4 ) );
  CLKBUF_X4 U3105 ( .I(\MC_ARK_ARC_1_3/buf_output[135] ), .Z(\SB1_4_9/i0[10] )
         );
  CLKBUF_X4 U3861 ( .I(\MC_ARK_ARC_1_3/buf_output[22] ), .Z(\SB1_4_28/i0_4 )
         );
  CLKBUF_X4 U785 ( .I(\MC_ARK_ARC_1_3/buf_output[103] ), .Z(\SB1_4_14/i0[6] )
         );
  CLKBUF_X4 \SB1_4_21/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[63] ), .Z(
        \SB1_4_21/i0[10] ) );
  CLKBUF_X4 \SB1_4_8/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[142] ), .Z(
        \SB1_4_8/i0_4 ) );
  CLKBUF_X4 U2760 ( .I(\MC_ARK_ARC_1_3/buf_output[134] ), .Z(\SB1_4_9/i0_0 )
         );
  CLKBUF_X4 U5034 ( .I(\MC_ARK_ARC_1_3/buf_output[21] ), .Z(\SB1_4_28/i0[10] )
         );
  CLKBUF_X4 U1899 ( .I(\MC_ARK_ARC_1_3/buf_output[128] ), .Z(\SB1_4_10/i0_0 )
         );
  CLKBUF_X8 U9076 ( .I(\RI1[4][41] ), .Z(\SB1_4_25/i0_3 ) );
  CLKBUF_X4 \SB1_4_2/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[177] ), .Z(
        \SB1_4_2/i0[10] ) );
  CLKBUF_X4 U3409 ( .I(\MC_ARK_ARC_1_3/buf_output[36] ), .Z(\SB1_4_25/i0[9] )
         );
  CLKBUF_X4 U2819 ( .I(\MC_ARK_ARC_1_3/buf_output[82] ), .Z(\SB1_4_18/i0_4 )
         );
  CLKBUF_X4 \SB1_4_21/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[60] ), .Z(
        \SB1_4_21/i0[9] ) );
  CLKBUF_X4 \SB1_4_23/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[52] ), .Z(
        \SB1_4_23/i0_4 ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_119_1  ( .I(\MC_ARK_ARC_1_3/buf_output[119] ), 
        .Z(\RI1[4][119] ) );
  CLKBUF_X4 \SB1_4_22/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[57] ), .Z(
        \SB1_4_22/i0[10] ) );
  CLKBUF_X4 \SB1_4_14/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[102] ), .Z(
        \SB1_4_14/i0[9] ) );
  CLKBUF_X4 U5406 ( .I(\MC_ARK_ARC_1_3/buf_output[138] ), .Z(\SB1_4_8/i0[9] )
         );
  CLKBUF_X4 U3967 ( .I(\SB1_4_26/buf_output[3] ), .Z(\SB2_4_24/i0[10] ) );
  CLKBUF_X4 \SB2_4_20/BUF_3  ( .I(\SB1_4_22/buf_output[3] ), .Z(
        \SB2_4_20/i0[10] ) );
  CLKBUF_X4 \SB2_4_1/BUF_1  ( .I(\SB1_4_5/buf_output[1] ), .Z(\SB2_4_1/i0[6] )
         );
  CLKBUF_X4 \SB2_4_25/BUF_0  ( .I(\SB1_4_30/buf_output[0] ), .Z(
        \SB2_4_25/i0[9] ) );
  CLKBUF_X4 U1972 ( .I(\SB1_4_9/buf_output[3] ), .Z(\SB2_4_7/i0[10] ) );
  CLKBUF_X4 U2394 ( .I(\SB1_4_26/buf_output[1] ), .Z(\SB2_4_22/i0[6] ) );
  CLKBUF_X4 U1446 ( .I(\SB1_4_28/buf_output[5] ), .Z(\SB2_4_28/i0_3 ) );
  CLKBUF_X4 \SB2_4_21/BUF_4  ( .I(\SB1_4_22/buf_output[4] ), .Z(
        \SB2_4_21/i0_4 ) );
  CLKBUF_X4 \SB2_4_14/BUF_3  ( .I(\SB1_4_16/buf_output[3] ), .Z(
        \SB2_4_14/i0[10] ) );
  CLKBUF_X4 \SB2_4_17/BUF_1  ( .I(\SB1_4_21/buf_output[1] ), .Z(
        \SB2_4_17/i0[6] ) );
  CLKBUF_X4 U702 ( .I(\SB1_4_1/buf_output[1] ), .Z(\SB2_4_29/i0[6] ) );
  CLKBUF_X4 \SB2_4_13/BUF_1  ( .I(\SB1_4_17/buf_output[1] ), .Z(
        \SB2_4_13/i0[6] ) );
  CLKBUF_X4 U2517 ( .I(\SB1_4_28/buf_output[1] ), .Z(\SB2_4_24/i0[6] ) );
  CLKBUF_X4 \SB2_4_17/BUF_0  ( .I(\SB1_4_22/buf_output[0] ), .Z(
        \SB2_4_17/i0[9] ) );
  CLKBUF_X4 \SB2_4_22/BUF_4  ( .I(\SB1_4_23/buf_output[4] ), .Z(
        \SB2_4_22/i0_4 ) );
  CLKBUF_X4 U9723 ( .I(\SB1_4_10/buf_output[0] ), .Z(\SB2_4_5/i0[9] ) );
  CLKBUF_X4 \SB2_4_3/BUF_4  ( .I(\SB1_4_4/buf_output[4] ), .Z(\SB2_4_3/i0_4 )
         );
  CLKBUF_X4 \SB2_4_3/BUF_3  ( .I(\SB1_4_5/buf_output[3] ), .Z(\SB2_4_3/i0[10] ) );
  CLKBUF_X4 U2670 ( .I(\SB1_4_9/buf_output[5] ), .Z(\SB2_4_9/i0_3 ) );
  CLKBUF_X4 \SB2_4_18/BUF_1  ( .I(\SB1_4_22/buf_output[1] ), .Z(
        \SB2_4_18/i0[6] ) );
  CLKBUF_X4 \SB2_4_15/BUF_4  ( .I(\SB1_4_16/buf_output[4] ), .Z(
        \SB2_4_15/i0_4 ) );
  CLKBUF_X4 \SB2_4_14/BUF_4  ( .I(\SB1_4_15/buf_output[4] ), .Z(
        \SB2_4_14/i0_4 ) );
  CLKBUF_X4 U5390 ( .I(\SB1_4_11/buf_output[4] ), .Z(\SB2_4_10/i0_4 ) );
  CLKBUF_X4 \SB2_4_4/BUF_3  ( .I(\SB1_4_6/buf_output[3] ), .Z(\SB2_4_4/i0[10] ) );
  CLKBUF_X4 U1973 ( .I(\SB1_4_10/buf_output[4] ), .Z(\SB2_4_9/i0_4 ) );
  CLKBUF_X4 U2579 ( .I(\SB1_4_16/buf_output[1] ), .Z(\SB2_4_12/i0[6] ) );
  CLKBUF_X4 \SB2_4_9/BUF_1  ( .I(\SB1_4_13/buf_output[1] ), .Z(\SB2_4_9/i0[6] ) );
  CLKBUF_X4 \SB2_4_19/BUF_1  ( .I(\SB1_4_23/buf_output[1] ), .Z(
        \SB2_4_19/i0[6] ) );
  CLKBUF_X4 U9398 ( .I(\SB1_4_26/buf_output[0] ), .Z(\SB2_4_21/i0[9] ) );
  CLKBUF_X4 \SB2_4_6/BUF_0  ( .I(\SB1_4_11/buf_output[0] ), .Z(\SB2_4_6/i0[9] ) );
  CLKBUF_X4 U9164 ( .I(\SB1_4_21/buf_output[2] ), .Z(\SB2_4_18/i0_0 ) );
  CLKBUF_X4 \SB2_4_10/BUF_2  ( .I(\SB1_4_13/buf_output[2] ), .Z(
        \SB2_4_10/i0_0 ) );
  CLKBUF_X4 \SB2_4_11/BUF_3  ( .I(\SB1_4_13/buf_output[3] ), .Z(
        \SB2_4_11/i0[10] ) );
  CLKBUF_X4 \SB2_4_11/BUF_0  ( .I(\SB1_4_16/buf_output[0] ), .Z(
        \SB2_4_11/i0[9] ) );
  CLKBUF_X4 U2395 ( .I(\SB1_4_10/buf_output[1] ), .Z(\SB2_4_6/i0[6] ) );
  CLKBUF_X4 \SB2_4_16/BUF_1  ( .I(\SB1_4_20/buf_output[1] ), .Z(
        \SB2_4_16/i0[6] ) );
  CLKBUF_X4 U5185 ( .I(\SB1_4_8/buf_output[3] ), .Z(\SB2_4_6/i0[10] ) );
  CLKBUF_X4 \SB2_4_6/BUF_2  ( .I(\SB1_4_9/buf_output[2] ), .Z(\SB2_4_6/i0_0 )
         );
  CLKBUF_X4 U761 ( .I(\SB1_4_17/buf_output[2] ), .Z(\SB2_4_14/i0_0 ) );
  CLKBUF_X4 U2975 ( .I(\SB1_4_18/buf_output[1] ), .Z(\SB2_4_14/i0[6] ) );
  CLKBUF_X4 \SB2_4_16/BUF_3  ( .I(\SB1_4_18/buf_output[3] ), .Z(
        \SB2_4_16/i0[10] ) );
  CLKBUF_X4 \SB2_4_30/BUF_3  ( .I(\SB1_4_0/buf_output[3] ), .Z(
        \SB2_4_30/i0[10] ) );
  CLKBUF_X4 U5216 ( .I(\SB1_4_13/buf_output[4] ), .Z(\SB2_4_12/i0_4 ) );
  CLKBUF_X4 \SB2_4_17/BUF_2  ( .I(\SB1_4_20/buf_output[2] ), .Z(
        \SB2_4_17/i0_0 ) );
  CLKBUF_X4 \SB2_4_29/BUF_2  ( .I(\SB1_4_0/buf_output[2] ), .Z(\SB2_4_29/i0_0 ) );
  CLKBUF_X4 U5143 ( .I(\SB1_4_26/buf_output[2] ), .Z(\SB2_4_23/i0_0 ) );
  CLKBUF_X4 U5466 ( .I(\RI3[4][188] ), .Z(\SB2_4_0/i0_0 ) );
  CLKBUF_X4 U5332 ( .I(\SB1_4_24/buf_output[3] ), .Z(\SB2_4_22/i0[10] ) );
  CLKBUF_X4 U5278 ( .I(\SB1_4_31/buf_output[1] ), .Z(\SB2_4_27/i0[6] ) );
  CLKBUF_X4 \SB2_4_22/BUF_0  ( .I(\SB1_4_27/buf_output[0] ), .Z(
        \SB2_4_22/i0[9] ) );
  CLKBUF_X4 \SB2_4_2/BUF_0  ( .I(\SB1_4_7/buf_output[0] ), .Z(\SB2_4_2/i0[9] )
         );
  CLKBUF_X4 \SB2_4_20/BUF_1  ( .I(\SB1_4_24/buf_output[1] ), .Z(
        \SB2_4_20/i0[6] ) );
  CLKBUF_X4 \SB2_4_23/BUF_4  ( .I(\SB1_4_24/buf_output[4] ), .Z(
        \SB2_4_23/i0_4 ) );
  CLKBUF_X4 \SB2_4_3/BUF_1  ( .I(\SB1_4_7/buf_output[1] ), .Z(\SB2_4_3/i0[6] )
         );
  CLKBUF_X4 \SB2_4_2/BUF_4  ( .I(\SB1_4_3/buf_output[4] ), .Z(\SB2_4_2/i0_4 )
         );
  CLKBUF_X4 \SB2_4_10/BUF_1  ( .I(\RI3[4][127] ), .Z(\SB2_4_10/i0[6] ) );
  CLKBUF_X4 \SB2_4_4/BUF_2  ( .I(\SB1_4_7/buf_output[2] ), .Z(\SB2_4_4/i0_0 )
         );
  CLKBUF_X4 \SB2_4_10/BUF_3  ( .I(\SB1_4_12/buf_output[3] ), .Z(
        \SB2_4_10/i0[10] ) );
  CLKBUF_X4 \SB2_4_26/BUF_4  ( .I(\SB1_4_27/buf_output[4] ), .Z(
        \SB2_4_26/i0_4 ) );
  CLKBUF_X4 U700 ( .I(\SB1_4_27/buf_output[2] ), .Z(\SB2_4_24/i0_0 ) );
  CLKBUF_X4 U5136 ( .I(\SB2_4_22/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[64] ) );
  CLKBUF_X4 U9376 ( .I(\SB2_4_7/buf_output[3] ), .Z(\RI5[4][159] ) );
  CLKBUF_X4 U9238 ( .I(\SB2_4_23/buf_output[2] ), .Z(\RI5[4][68] ) );
  CLKBUF_X4 U2611 ( .I(\SB2_4_27/buf_output[2] ), .Z(\RI5[4][44] ) );
  CLKBUF_X4 U4681 ( .I(\RI1[5][59] ), .Z(\SB3_22/i0_3 ) );
  CLKBUF_X4 U2346 ( .I(\MC_ARK_ARC_1_4/buf_output[58] ), .Z(\SB3_22/i0_4 ) );
  CLKBUF_X4 U2424 ( .I(\MC_ARK_ARC_1_4/buf_output[2] ), .Z(\SB3_31/i0_0 ) );
  CLKBUF_X4 \SB3_26/BUF_4  ( .I(\MC_ARK_ARC_1_4/buf_output[34] ), .Z(
        \SB3_26/i0_4 ) );
  CLKBUF_X4 U1948 ( .I(\MC_ARK_ARC_1_4/buf_output[109] ), .Z(\SB3_13/i0[6] )
         );
  CLKBUF_X4 U4038 ( .I(\MC_ARK_ARC_1_4/buf_output[160] ), .Z(\SB3_5/i0_4 ) );
  CLKBUF_X4 \SB3_28/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[18] ), .Z(
        \SB3_28/i0[9] ) );
  CLKBUF_X4 \SB3_3/BUF_4  ( .I(\MC_ARK_ARC_1_4/buf_output[172] ), .Z(
        \SB3_3/i0_4 ) );
  BUF_X2 \SB3_5/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[156] ), .Z(
        \SB3_5/i0[9] ) );
  CLKBUF_X4 U9738 ( .I(\MC_ARK_ARC_1_4/buf_output[75] ), .Z(\SB3_19/i0[10] )
         );
  CLKBUF_X4 U3103 ( .I(\MC_ARK_ARC_1_4/buf_output[16] ), .Z(\SB3_29/i0_4 ) );
  CLKBUF_X4 \SB3_26/BUF_1  ( .I(\MC_ARK_ARC_1_4/buf_output[31] ), .Z(
        \SB3_26/i0[6] ) );
  CLKBUF_X4 U4944 ( .I(\MC_ARK_ARC_1_4/buf_output[100] ), .Z(\SB3_15/i0_4 ) );
  CLKBUF_X4 U1365 ( .I(\MC_ARK_ARC_1_4/buf_output[147] ), .Z(\SB3_7/i0[10] )
         );
  CLKBUF_X4 U623 ( .I(\MC_ARK_ARC_1_4/buf_output[52] ), .Z(\SB3_23/i0_4 ) );
  CLKBUF_X4 U4954 ( .I(\MC_ARK_ARC_1_4/buf_output[145] ), .Z(\SB3_7/i0[6] ) );
  CLKBUF_X4 U640 ( .I(\MC_ARK_ARC_1_4/buf_output[136] ), .Z(\SB3_9/i0_4 ) );
  CLKBUF_X4 U2392 ( .I(\MC_ARK_ARC_1_4/buf_output[131] ), .Z(\SB3_10/i0_3 ) );
  CLKBUF_X4 \SB3_26/BUF_3  ( .I(\MC_ARK_ARC_1_4/buf_output[33] ), .Z(
        \SB3_26/i0[10] ) );
  CLKBUF_X4 U1887 ( .I(n6287), .Z(\SB3_25/i0_0 ) );
  CLKBUF_X4 U1953 ( .I(\MC_ARK_ARC_1_4/buf_output[103] ), .Z(\SB3_14/i0[6] )
         );
  CLKBUF_X4 U657 ( .I(\MC_ARK_ARC_1_4/buf_output[130] ), .Z(\SB3_10/i0_4 ) );
  CLKBUF_X4 U5048 ( .I(\MC_ARK_ARC_1_4/buf_output[190] ), .Z(\SB3_0/i0_4 ) );
  CLKBUF_X4 \SB3_24/BUF_4  ( .I(\MC_ARK_ARC_1_4/buf_output[46] ), .Z(
        \SB3_24/i0_4 ) );
  INV_X2 \SB3_29/INV_5  ( .I(n3976), .ZN(\SB3_29/i1_5 ) );
  CLKBUF_X8 \SB3_17/BUF_5  ( .I(\RI1[5][89] ), .Z(\SB3_17/i0_3 ) );
  CLKBUF_X8 U3380 ( .I(\RI1[5][179] ), .Z(\SB3_2/i0_3 ) );
  BUF_X2 \SB4_17/BUF_0  ( .I(\SB3_22/buf_output[0] ), .Z(\SB4_17/i0[9] ) );
  CLKBUF_X4 U1313 ( .I(\SB3_9/buf_output[4] ), .Z(\SB4_8/i0_4 ) );
  CLKBUF_X4 U9584 ( .I(\SB3_18/buf_output[3] ), .Z(\SB4_16/i0[10] ) );
  CLKBUF_X4 U9535 ( .I(\SB3_22/buf_output[5] ), .Z(\SB4_22/i0_3 ) );
  CLKBUF_X4 \SB4_2/BUF_4  ( .I(\SB3_3/buf_output[4] ), .Z(\SB4_2/i0_4 ) );
  BUF_X2 U1930 ( .I(\SB3_8/buf_output[1] ), .Z(\SB4_4/i0[6] ) );
  CLKBUF_X4 U9474 ( .I(\SB3_22/buf_output[4] ), .Z(\SB4_21/i0_4 ) );
  CLKBUF_X4 \SB4_11/BUF_0  ( .I(\SB3_16/buf_output[0] ), .Z(\SB4_11/i0[9] ) );
  CLKBUF_X4 U261 ( .I(\SB3_28/buf_output[0] ), .Z(\SB4_23/i0[9] ) );
  CLKBUF_X4 U2451 ( .I(\SB3_3/buf_output[2] ), .Z(\SB4_0/i0_0 ) );
  CLKBUF_X4 U247 ( .I(\SB3_6/buf_output[4] ), .Z(\SB4_5/i0_4 ) );
  CLKBUF_X4 U1547 ( .I(\SB3_30/buf_output[3] ), .Z(\SB4_28/i0[10] ) );
  CLKBUF_X4 U1326 ( .I(\SB3_31/buf_output[4] ), .Z(\SB4_30/i0_4 ) );
  CLKBUF_X4 U3063 ( .I(\SB3_2/buf_output[0] ), .Z(\SB4_29/i0[9] ) );
  CLKBUF_X4 U9503 ( .I(\SB3_2/buf_output[4] ), .Z(\SB4_1/i0_4 ) );
  BUF_X4 U654 ( .I(\RI1[5][35] ), .Z(\SB3_26/i0_3 ) );
  NAND2_X2 U1268 ( .A1(\SB1_0_6/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_6/Component_Function_0/NAND4_in[1] ), .ZN(n1986) );
  NAND2_X2 U1203 ( .A1(\SB1_3_10/Component_Function_4/NAND4_in[1] ), .A2(n4937), .ZN(n4936) );
  BUF_X4 \SB2_1_1/BUF_4  ( .I(\SB1_1_2/buf_output[4] ), .Z(\SB2_1_1/i0_4 ) );
  BUF_X4 U2291 ( .I(\MC_ARK_ARC_1_2/buf_output[40] ), .Z(\SB1_3_25/i0_4 ) );
  INV_X2 U3042 ( .I(\RI1[5][35] ), .ZN(\SB3_26/i1_5 ) );
  BUF_X4 U9780 ( .I(\MC_ARK_ARC_1_1/buf_output[44] ), .Z(\SB1_2_24/i0_0 ) );
  NAND3_X2 \SB2_1_20/Component_Function_4/N2  ( .A1(\SB2_1_20/i3[0] ), .A2(
        \SB2_1_20/i0_0 ), .A3(\SB2_1_20/i1_7 ), .ZN(
        \SB2_1_20/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 \SB2_3_11/BUF_3_0  ( .I(\SB2_3_11/buf_output[3] ), .Z(\RI5[3][135] )
         );
  NAND3_X2 \SB2_2_2/Component_Function_1/N3  ( .A1(\SB2_2_2/i1_5 ), .A2(
        \SB2_2_2/i0[6] ), .A3(\SB2_2_2/i0[9] ), .ZN(
        \SB2_2_2/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 U1894 ( .I(\MC_ARK_ARC_1_0/buf_output[44] ), .Z(\SB1_1_24/i0_0 ) );
  BUF_X4 \SB1_3_0/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[190] ), .Z(
        \SB1_3_0/i0_4 ) );
  NAND3_X2 \SB1_4_13/Component_Function_2/N4  ( .A1(\SB1_4_13/i1_5 ), .A2(
        \SB1_4_13/i0_0 ), .A3(\SB1_4_13/i0_4 ), .ZN(
        \SB1_4_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U7651 ( .A1(\SB1_3_19/i0[8] ), .A2(\SB1_3_19/i0_4 ), .A3(
        \SB1_3_19/i1_7 ), .ZN(n2497) );
  NAND3_X2 \SB1_1_30/Component_Function_2/N1  ( .A1(\SB1_1_30/i1_5 ), .A2(
        \SB1_1_30/i0[10] ), .A3(\SB1_1_30/i1[9] ), .ZN(
        \SB1_1_30/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB3_13/BUF_4  ( .I(\MC_ARK_ARC_1_4/buf_output[112] ), .Z(
        \SB3_13/i0_4 ) );
  NAND3_X2 U1179 ( .A1(\SB1_3_19/i0_3 ), .A2(\SB1_3_19/i1_7 ), .A3(
        \SB1_3_19/i0[8] ), .ZN(\SB1_3_19/Component_Function_1/NAND4_in[1] ) );
  BUF_X2 U9602 ( .I(\MC_ARK_ARC_1_4/buf_output[17] ), .Z(n3976) );
  NAND3_X2 U1208 ( .A1(\SB2_0_31/i0[6] ), .A2(\SB2_0_31/i0[9] ), .A3(
        \RI3[0][4] ), .ZN(n2901) );
  NAND2_X2 \SB2_1_0/Component_Function_0/N1  ( .A1(\SB2_1_0/i0[10] ), .A2(
        \SB2_1_0/i0[9] ), .ZN(\SB2_1_0/Component_Function_0/NAND4_in[0] ) );
  BUF_X2 \SB1_0_19/BUF_0  ( .I(n277), .Z(\SB1_0_19/i0[9] ) );
  BUF_X2 \SB1_0_6/BUF_1  ( .I(n246), .Z(\SB1_0_6/i0[6] ) );
  BUF_X2 \SB1_0_0/BUF_4  ( .I(n380), .Z(\SB1_0_0/i0_4 ) );
  BUF_X2 \SB1_0_27/BUF_4  ( .I(n326), .Z(\SB1_0_27/i0_4 ) );
  BUF_X2 \SB1_0_12/BUF_3  ( .I(n355), .Z(\SB1_0_12/i0[10] ) );
  NAND3_X1 U10936 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0_4 ), .A3(
        \SB1_0_6/i1[9] ), .ZN(\SB1_0_6/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1246 ( .A1(\SB1_0_6/i0_0 ), .A2(\SB1_0_6/i0[10] ), .A3(
        \SB1_0_6/i0[6] ), .ZN(\SB1_0_6/Component_Function_5/NAND4_in[1] ) );
  BUF_X2 \SB1_0_10/BUF_4  ( .I(n360), .Z(\SB1_0_10/i0_4 ) );
  BUF_X2 \SB1_0_5/BUF_2  ( .I(n6281), .Z(\SB1_0_5/i0_0 ) );
  BUF_X2 U9792 ( .I(n357), .Z(\SB1_0_11/i0[10] ) );
  INV_X1 \SB1_0_26/INV_2  ( .I(n264), .ZN(\SB1_0_26/i1[9] ) );
  INV_X1 \SB1_0_0/INV_2  ( .I(n316), .ZN(\SB1_0_0/i1[9] ) );
  NAND3_X1 \SB1_0_13/Component_Function_4/N4  ( .A1(\SB1_0_13/i1[9] ), .A2(
        \SB1_0_13/i1_5 ), .A3(\SB1_0_13/i0_4 ), .ZN(
        \SB1_0_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1277 ( .A1(\SB1_0_6/i0_0 ), .A2(\SB1_0_6/i0[7] ), .A3(
        \SB1_0_6/i0_3 ), .ZN(\SB1_0_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3854 ( .A1(\SB1_0_8/i0[10] ), .A2(\SB1_0_8/i0_3 ), .A3(
        \SB1_0_8/i0[9] ), .ZN(n1076) );
  NAND3_X1 U10000 ( .A1(\SB1_0_9/i0_0 ), .A2(\SB1_0_9/i0_3 ), .A3(
        \SB1_0_9/i0[7] ), .ZN(n4088) );
  BUF_X2 \SB1_0_25/BUF_1  ( .I(n227), .Z(\SB1_0_25/i0[6] ) );
  NAND3_X1 U6171 ( .A1(\SB1_0_18/i0[8] ), .A2(\SB1_0_18/i1_5 ), .A3(
        \SB1_0_18/i3[0] ), .ZN(\SB1_0_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U12508 ( .A1(\SB1_0_12/i0_0 ), .A2(\SB1_0_12/i1_5 ), .A3(
        \SB1_0_12/i0_4 ), .ZN(n5317) );
  NAND3_X1 U1274 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0[10] ), .A3(
        \SB1_0_15/i0[9] ), .ZN(n2609) );
  NAND3_X1 \SB1_0_10/Component_Function_3/N3  ( .A1(\SB1_0_10/i1[9] ), .A2(
        \SB1_0_10/i1_7 ), .A3(\SB1_0_10/i0[10] ), .ZN(
        \SB1_0_10/Component_Function_3/NAND4_in[2] ) );
  BUF_X2 \SB1_0_7/BUF_1  ( .I(n245), .Z(\SB1_0_7/i0[6] ) );
  NAND3_X1 U5599 ( .A1(\SB1_0_24/i0_3 ), .A2(\SB1_0_24/i0_0 ), .A3(
        \SB1_0_24/i0_4 ), .ZN(\SB1_0_24/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 \SB1_0_7/BUF_0  ( .I(n301), .Z(\SB1_0_7/i0[9] ) );
  CLKBUF_X2 \SB1_0_23/BUF_1  ( .I(n229), .Z(\SB1_0_23/i0[6] ) );
  BUF_X2 \SB1_0_2/BUF_4  ( .I(n376), .Z(\SB1_0_2/i0_4 ) );
  BUF_X2 \SB1_0_30/BUF_1  ( .I(n222), .Z(\SB1_0_30/i0[6] ) );
  INV_X1 \SB1_0_14/INV_2  ( .I(n288), .ZN(\SB1_0_14/i1[9] ) );
  INV_X1 \SB1_0_31/INV_3  ( .I(n317), .ZN(\SB1_0_31/i0[8] ) );
  NAND3_X1 U2141 ( .A1(\SB1_0_6/i0[10] ), .A2(\SB1_0_6/i0_3 ), .A3(
        \SB1_0_6/i0[9] ), .ZN(n4727) );
  NAND3_X1 U3549 ( .A1(\SB1_0_21/i1[9] ), .A2(\SB1_0_21/i1_5 ), .A3(
        \SB1_0_21/i0_4 ), .ZN(\SB1_0_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2098 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i1[9] ), .A3(
        \SB1_0_23/i0[6] ), .ZN(\SB1_0_23/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_4/Component_Function_1/N1  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i1[9] ), .ZN(\SB1_0_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U9295 ( .A1(\SB1_0_15/i0[6] ), .A2(\SB1_0_15/i1_5 ), .A3(
        \SB1_0_15/i0[9] ), .ZN(\SB1_0_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_28/Component_Function_2/N1  ( .A1(\SB1_0_28/i1_5 ), .A2(
        \SB1_0_28/i0[10] ), .A3(\SB1_0_28/i1[9] ), .ZN(
        \SB1_0_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_0/N4  ( .A1(\SB1_0_20/i0[7] ), .A2(
        \SB1_0_20/i0_3 ), .A3(\SB1_0_20/i0_0 ), .ZN(
        \SB1_0_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_16/Component_Function_3/N3  ( .A1(\SB1_0_16/i1[9] ), .A2(
        \SB1_0_16/i1_7 ), .A3(\SB1_0_16/i0[10] ), .ZN(
        \SB1_0_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2077 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0_4 ), .A3(
        \SB1_0_6/i0_0 ), .ZN(\SB1_0_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_24/Component_Function_5/N2  ( .A1(\SB1_0_24/i0_0 ), .A2(
        \SB1_0_24/i0[6] ), .A3(\SB1_0_24/i0[10] ), .ZN(
        \SB1_0_24/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_1/Component_Function_2/N2  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i0[10] ), .A3(\SB1_0_1/i0[6] ), .ZN(
        \SB1_0_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3523 ( .A1(\SB1_0_4/i0[10] ), .A2(\SB1_0_4/i1[9] ), .A3(
        \SB1_0_4/i1_7 ), .ZN(n2622) );
  NAND3_X1 \SB1_0_4/Component_Function_1/N4  ( .A1(\SB1_0_4/i1_7 ), .A2(
        \SB1_0_4/i0[8] ), .A3(\SB1_0_4/i0_4 ), .ZN(
        \SB1_0_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_11/Component_Function_3/N1  ( .A1(\SB1_0_11/i1[9] ), .A2(
        \SB1_0_11/i0_3 ), .A3(\SB1_0_11/i0[6] ), .ZN(
        \SB1_0_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_1/N4  ( .A1(\SB1_0_21/i1_7 ), .A2(
        \SB1_0_21/i0[8] ), .A3(\SB1_0_21/i0_4 ), .ZN(
        \SB1_0_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_5/Component_Function_1/N4  ( .A1(\SB1_0_5/i1_7 ), .A2(
        \SB1_0_5/i0[8] ), .A3(\SB1_0_5/i0_4 ), .ZN(
        \SB1_0_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_23/Component_Function_2/N1  ( .A1(\SB1_0_23/i1_5 ), .A2(
        \SB1_0_23/i0[10] ), .A3(\SB1_0_23/i1[9] ), .ZN(
        \SB1_0_23/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_13/Component_Function_1/N1  ( .A1(\SB1_0_13/i0_3 ), .A2(
        \SB1_0_13/i1[9] ), .ZN(\SB1_0_13/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_0/Component_Function_5/N1  ( .A1(\SB1_0_0/i0_0 ), .A2(
        \SB1_0_0/i3[0] ), .ZN(\SB1_0_0/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_15/Component_Function_5/N1  ( .A1(\SB1_0_15/i0_0 ), .A2(
        \SB1_0_15/i3[0] ), .ZN(\SB1_0_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3278 ( .A1(\SB1_0_16/i0_3 ), .A2(n6149), .A3(\SB1_0_16/i0[8] ), 
        .ZN(n864) );
  NAND3_X1 \SB1_0_2/Component_Function_1/N2  ( .A1(\SB1_0_2/i0_3 ), .A2(
        \SB1_0_2/i1_7 ), .A3(\SB1_0_2/i0[8] ), .ZN(
        \SB1_0_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_13/Component_Function_5/N1  ( .A1(\SB1_0_13/i0_0 ), .A2(
        \SB1_0_13/i3[0] ), .ZN(\SB1_0_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_5/N4  ( .A1(\SB1_0_23/i0[9] ), .A2(
        \SB1_0_23/i0[6] ), .A3(\SB1_0_23/i0_4 ), .ZN(
        \SB1_0_23/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_28/Component_Function_5/N1  ( .A1(\SB1_0_28/i0_0 ), .A2(
        \SB1_0_28/i3[0] ), .ZN(\SB1_0_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_3/N1  ( .A1(\SB1_0_16/i1[9] ), .A2(
        \SB1_0_16/i0_3 ), .A3(\SB1_0_16/i0[6] ), .ZN(
        \SB1_0_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_3/N1  ( .A1(\SB1_0_27/i1[9] ), .A2(
        \SB1_0_27/i0_3 ), .A3(\SB1_0_27/i0[6] ), .ZN(
        \SB1_0_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_1/N4  ( .A1(\SB1_0_13/i1_7 ), .A2(
        n5428), .A3(\SB1_0_13/i0_4 ), .ZN(
        \SB1_0_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_2/N2  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i0[10] ), .A3(\SB1_0_31/i0[6] ), .ZN(
        \SB1_0_31/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_16/Component_Function_5/N1  ( .A1(\SB1_0_16/i0_0 ), .A2(
        \SB1_0_16/i3[0] ), .ZN(\SB1_0_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U11219 ( .A1(\SB1_0_29/i0_3 ), .A2(\SB1_0_29/i0[10] ), .A3(
        \SB1_0_29/i0[6] ), .ZN(n4621) );
  AOI21_X1 U11584 ( .A1(\SB1_0_10/i3[0] ), .A2(\SB1_0_10/i0_0 ), .B(n4804), 
        .ZN(n4803) );
  NAND2_X1 \SB1_0_15/Component_Function_0/N1  ( .A1(\SB1_0_15/i0[10] ), .A2(
        \SB1_0_15/i0[9] ), .ZN(\SB1_0_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_5/N4  ( .A1(\SB1_0_24/i0[9] ), .A2(
        \SB1_0_24/i0[6] ), .A3(\SB1_0_24/i0_4 ), .ZN(
        \SB1_0_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_28/Component_Function_2/N2  ( .A1(\SB1_0_28/i0_3 ), .A2(
        \SB1_0_28/i0[10] ), .A3(\SB1_0_28/i0[6] ), .ZN(
        \SB1_0_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_30/Component_Function_1/N4  ( .A1(\SB1_0_30/i1_7 ), .A2(
        \SB1_0_30/i0[8] ), .A3(\SB1_0_30/i0_4 ), .ZN(
        \SB1_0_30/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 U10001 ( .A1(\SB1_0_9/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_9/Component_Function_0/NAND4_in[0] ), .ZN(n4089) );
  NAND3_X1 \SB1_0_24/Component_Function_0/N2  ( .A1(\SB1_0_24/i0[8] ), .A2(
        \SB1_0_24/i0[7] ), .A3(\SB1_0_24/i0[6] ), .ZN(
        \SB1_0_24/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_29/Component_Function_5/N3  ( .A1(\SB1_0_29/i1[9] ), .A2(
        \SB1_0_29/i0_4 ), .A3(\SB1_0_29/i0_3 ), .ZN(
        \SB1_0_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_13/Component_Function_2/N4  ( .A1(\SB1_0_13/i1_5 ), .A2(
        \SB1_0_13/i0_0 ), .A3(\SB1_0_13/i0_4 ), .ZN(
        \SB1_0_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_5/N2  ( .A1(\SB1_0_9/i0_0 ), .A2(
        \SB1_0_9/i0[6] ), .A3(\SB1_0_9/i0[10] ), .ZN(
        \SB1_0_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_25/Component_Function_2/N1  ( .A1(\SB1_0_25/i1_5 ), .A2(
        \SB1_0_25/i0[10] ), .A3(\SB1_0_25/i1[9] ), .ZN(
        \SB1_0_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_0/N2  ( .A1(\SB1_0_15/i0[8] ), .A2(
        \SB1_0_15/i0[7] ), .A3(\SB1_0_15/i0[6] ), .ZN(
        \SB1_0_15/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U11545 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i0[10] ), .A3(
        \SB1_0_23/i0[9] ), .ZN(\SB1_0_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_15/Component_Function_1/N4  ( .A1(\SB1_0_15/i1_7 ), .A2(
        \SB1_0_15/i0[8] ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_24/Component_Function_5/N1  ( .A1(\SB1_0_24/i0_0 ), .A2(
        \SB1_0_24/i3[0] ), .ZN(\SB1_0_24/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_5/Component_Function_1/N1  ( .A1(\SB1_0_5/i0_3 ), .A2(
        \SB1_0_5/i1[9] ), .ZN(\SB1_0_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_3/N1  ( .A1(\SB1_0_1/i1[9] ), .A2(
        \SB1_0_1/i0_3 ), .A3(\SB1_0_1/i0[6] ), .ZN(
        \SB1_0_1/Component_Function_3/NAND4_in[0] ) );
  INV_X1 \SB2_0_9/INV_5  ( .I(\SB1_0_9/buf_output[5] ), .ZN(\SB2_0_9/i1_5 ) );
  INV_X2 \SB2_0_12/INV_4  ( .I(\RI3[0][118] ), .ZN(\SB2_0_12/i0[7] ) );
  BUF_X2 U12418 ( .I(\SB1_0_25/buf_output[0] ), .Z(n5264) );
  BUF_X2 \SB2_0_25/BUF_0  ( .I(\SB1_0_30/buf_output[0] ), .Z(\SB2_0_25/i0[9] )
         );
  BUF_X2 \SB2_0_10/BUF_1  ( .I(\RI3[0][127] ), .Z(\SB2_0_10/i0[6] ) );
  BUF_X2 \SB2_0_11/BUF_0  ( .I(\RI3[0][120] ), .Z(\SB2_0_11/i0[9] ) );
  INV_X4 \SB2_0_19/INV_5  ( .I(\RI3[0][77] ), .ZN(\SB2_0_19/i1_5 ) );
  CLKBUF_X2 \SB2_0_28/BUF_1  ( .I(\RI3[0][19] ), .Z(\SB2_0_28/i0[6] ) );
  INV_X2 U6466 ( .I(n2965), .ZN(\SB2_0_10/i0_4 ) );
  BUF_X2 \SB2_0_2/BUF_1  ( .I(\RI3[0][175] ), .Z(\SB2_0_2/i0[6] ) );
  BUF_X2 \SB2_0_27/BUF_3  ( .I(\RI3[0][27] ), .Z(\SB2_0_27/i0[10] ) );
  CLKBUF_X2 \SB2_0_14/BUF_2  ( .I(\SB1_0_17/buf_output[2] ), .Z(
        \SB2_0_14/i0_0 ) );
  BUF_X2 U2062 ( .I(\RI3[0][30] ), .Z(\SB2_0_26/i0[9] ) );
  BUF_X2 \SB2_0_24/BUF_1  ( .I(\SB1_0_28/buf_output[1] ), .Z(\SB2_0_24/i0[6] )
         );
  CLKBUF_X2 \SB2_0_21/BUF_1  ( .I(\SB1_0_25/buf_output[1] ), .Z(
        \SB2_0_21/i0[6] ) );
  BUF_X2 \SB2_0_17/BUF_1  ( .I(\SB1_0_21/buf_output[1] ), .Z(\SB2_0_17/i0[6] )
         );
  INV_X1 \SB2_0_8/INV_4  ( .I(\RI3[0][142] ), .ZN(\SB2_0_8/i0[7] ) );
  INV_X2 U7230 ( .I(n2822), .ZN(\SB2_0_14/i0_4 ) );
  INV_X1 \SB2_0_30/INV_5  ( .I(\SB1_0_30/buf_output[5] ), .ZN(\SB2_0_30/i1_5 )
         );
  INV_X1 \SB2_0_28/INV_5  ( .I(\SB1_0_28/buf_output[5] ), .ZN(\SB2_0_28/i1_5 )
         );
  INV_X1 \SB2_0_26/INV_5  ( .I(\RI3[0][35] ), .ZN(\SB2_0_26/i1_5 ) );
  INV_X1 U5444 ( .I(\RI3[0][187] ), .ZN(\SB2_0_0/i1_7 ) );
  INV_X1 \SB2_0_27/INV_4  ( .I(\RI3[0][28] ), .ZN(\SB2_0_27/i0[7] ) );
  BUF_X2 \SB2_0_23/BUF_0  ( .I(\SB1_0_28/buf_output[0] ), .Z(\SB2_0_23/i0[9] )
         );
  NAND3_X1 \SB2_0_4/Component_Function_5/N3  ( .A1(\SB2_0_4/i1[9] ), .A2(
        \RI3[0][166] ), .A3(\SB2_0_4/i0_3 ), .ZN(
        \SB2_0_4/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_0/Component_Function_1/N1  ( .A1(\SB2_0_0/i0_3 ), .A2(
        \SB2_0_0/i1[9] ), .ZN(\SB2_0_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2925 ( .A1(\SB2_0_28/i0[10] ), .A2(\SB2_0_28/i1_7 ), .A3(
        \SB2_0_28/i1[9] ), .ZN(n4541) );
  NAND3_X1 \SB2_0_29/Component_Function_2/N2  ( .A1(\SB2_0_29/i0_3 ), .A2(
        \SB2_0_29/i0[10] ), .A3(\SB2_0_29/i0[6] ), .ZN(
        \SB2_0_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3259 ( .A1(\SB2_0_13/i0_3 ), .A2(\RI3[0][112] ), .A3(
        \SB2_0_13/i1[9] ), .ZN(n2431) );
  NAND3_X1 U10826 ( .A1(\SB2_0_3/i0[10] ), .A2(\SB2_0_3/i1[9] ), .A3(
        \SB2_0_3/i1_7 ), .ZN(n4465) );
  NAND3_X1 \SB2_0_19/Component_Function_5/N2  ( .A1(\SB2_0_19/i0_0 ), .A2(
        \SB2_0_19/i0[6] ), .A3(\RI3[0][75] ), .ZN(
        \SB2_0_19/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_21/Component_Function_1/N1  ( .A1(\SB2_0_21/i0_3 ), .A2(
        \SB2_0_21/i1[9] ), .ZN(\SB2_0_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3575 ( .A1(\SB2_0_2/i0_3 ), .A2(\SB2_0_2/i0[10] ), .A3(
        \SB2_0_2/i0[6] ), .ZN(\SB2_0_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U6807 ( .A1(\SB2_0_9/i0_3 ), .A2(\SB2_0_9/i0[10] ), .A3(
        \SB2_0_9/i0[9] ), .ZN(n3590) );
  NAND3_X1 U1205 ( .A1(\SB2_0_18/i0[10] ), .A2(\SB2_0_18/i0_3 ), .A3(
        \RI3[0][82] ), .ZN(\SB2_0_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_6/Component_Function_2/N1  ( .A1(\SB2_0_6/i1_5 ), .A2(
        \SB2_0_6/i0[10] ), .A3(\SB2_0_6/i1[9] ), .ZN(
        \SB2_0_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_4/N1  ( .A1(\SB2_0_15/i0[9] ), .A2(
        \SB1_0_18/buf_output[2] ), .A3(\SB2_0_15/i0[8] ), .ZN(
        \SB2_0_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U10683 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i0_0 ), .A3(
        \SB2_0_11/i0[7] ), .ZN(n4382) );
  NAND3_X1 \SB2_0_6/Component_Function_1/N2  ( .A1(\SB2_0_6/i0_3 ), .A2(
        \SB2_0_6/i1_7 ), .A3(\SB2_0_6/i0[8] ), .ZN(
        \SB2_0_6/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_0/Component_Function_0/N2  ( .A1(n4003), .A2(\SB2_0_0/i0[7] ), .A3(\SB2_0_0/i0[6] ), .ZN(\SB2_0_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3596 ( .A1(\SB2_0_24/i0_0 ), .A2(\RI3[0][46] ), .A3(
        \SB2_0_24/i0_3 ), .ZN(n1794) );
  NAND3_X1 U5723 ( .A1(\SB2_0_22/i0[10] ), .A2(\SB2_0_22/i1[9] ), .A3(
        \SB2_0_22/i1_7 ), .ZN(n1617) );
  NAND2_X1 \SB2_0_13/Component_Function_5/N1  ( .A1(\SB2_0_13/i0_0 ), .A2(
        \SB2_0_13/i3[0] ), .ZN(\SB2_0_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U8040 ( .A1(n2886), .A2(n4847), .A3(\SB2_0_9/i1_7 ), .ZN(
        \SB2_0_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1180 ( .A1(\SB2_0_16/i0[8] ), .A2(n594), .A3(\SB2_0_16/i1_7 ), 
        .ZN(\SB2_0_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1941 ( .A1(\SB2_0_27/i0[7] ), .A2(\SB2_0_27/i0[8] ), .A3(
        \SB2_0_27/i0[6] ), .ZN(n3507) );
  NAND3_X1 \SB2_0_26/Component_Function_3/N3  ( .A1(\SB2_0_26/i1[9] ), .A2(
        \SB2_0_26/i1_7 ), .A3(\RI3[0][33] ), .ZN(
        \SB2_0_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_3/N1  ( .A1(\SB2_0_24/i1[9] ), .A2(
        \SB2_0_24/i0_3 ), .A3(\SB2_0_24/i0[6] ), .ZN(
        \SB2_0_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_0/N2  ( .A1(\SB2_0_26/i0[8] ), .A2(
        n3510), .A3(\SB2_0_26/i0[6] ), .ZN(
        \SB2_0_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_13/Component_Function_3/N3  ( .A1(\SB2_0_13/i1[9] ), .A2(
        \SB2_0_13/i1_7 ), .A3(\SB2_0_13/i0[10] ), .ZN(
        \SB2_0_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1957 ( .A1(\SB2_0_4/i1_7 ), .A2(\SB2_0_4/i0[8] ), .A3(
        \RI3[0][166] ), .ZN(\SB2_0_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_29/Component_Function_3/N4  ( .A1(\SB2_0_29/i1_5 ), .A2(
        \SB2_0_29/i0[8] ), .A3(\SB2_0_29/i3[0] ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_20/Component_Function_0/N2  ( .A1(\SB2_0_20/i0[8] ), .A2(
        \SB2_0_20/i0[7] ), .A3(\SB2_0_20/i0[6] ), .ZN(
        \SB2_0_20/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U12162 ( .A1(\SB2_0_9/i0[9] ), .A2(\SB2_0_9/i0_3 ), .A3(
        \SB2_0_9/i0[8] ), .ZN(n5119) );
  NAND3_X1 \SB2_0_28/Component_Function_3/N4  ( .A1(\SB2_0_28/i1_5 ), .A2(
        \SB2_0_28/i0[8] ), .A3(\SB2_0_28/i3[0] ), .ZN(
        \SB2_0_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U7317 ( .A1(\SB2_0_2/i0_0 ), .A2(\SB2_0_2/i1_5 ), .A3(\RI3[0][178] ), .ZN(n3647) );
  NAND3_X1 U8522 ( .A1(n2592), .A2(\SB2_0_1/i0[8] ), .A3(\SB2_0_1/i1_5 ), .ZN(
        n3842) );
  NAND3_X1 \SB2_0_15/Component_Function_2/N4  ( .A1(\SB2_0_15/i1_5 ), .A2(
        \SB1_0_18/buf_output[2] ), .A3(\RI3[0][100] ), .ZN(
        \SB2_0_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U10723 ( .A1(\SB2_0_17/i0[9] ), .A2(\SB2_0_17/i0[6] ), .A3(
        \SB2_0_17/i1_5 ), .ZN(n4661) );
  NAND3_X1 U7623 ( .A1(\SB2_0_12/i0[7] ), .A2(\SB2_0_12/i0[8] ), .A3(
        \SB2_0_12/i0[6] ), .ZN(n2682) );
  NAND3_X1 U1960 ( .A1(\SB2_0_22/i0[9] ), .A2(\RI3[0][55] ), .A3(\RI3[0][58] ), 
        .ZN(\SB2_0_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U6540 ( .A1(\SB2_0_30/i0_3 ), .A2(\SB2_0_30/i0[8] ), .A3(
        \SB2_0_30/i1_7 ), .ZN(\SB2_0_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_22/Component_Function_4/N2  ( .A1(\SB2_0_22/i3[0] ), .A2(
        \SB2_0_22/i0_0 ), .A3(\SB2_0_22/i1_7 ), .ZN(
        \SB2_0_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_23/Component_Function_1/N4  ( .A1(\SB2_0_23/i1_7 ), .A2(
        \SB2_0_23/i0[8] ), .A3(\RI3[0][52] ), .ZN(
        \SB2_0_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_16/Component_Function_1/N3  ( .A1(\SB2_0_16/i1_5 ), .A2(
        \SB2_0_16/i0[6] ), .A3(n5157), .ZN(
        \SB2_0_16/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_6/Component_Function_5/N1  ( .A1(\SB2_0_6/i0_0 ), .A2(
        \SB2_0_6/i3[0] ), .ZN(\SB2_0_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U6650 ( .A1(\SB2_0_20/i0_3 ), .A2(\SB2_0_20/i0[7] ), .A3(
        \SB2_0_20/i0_0 ), .ZN(\SB2_0_20/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_16/Component_Function_1/N1  ( .A1(\SB2_0_16/i0_3 ), .A2(
        \SB2_0_16/i1[9] ), .ZN(\SB2_0_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_3/N1  ( .A1(\SB2_0_5/i1[9] ), .A2(
        \SB2_0_5/i0_3 ), .A3(\SB2_0_5/i0[6] ), .ZN(
        \SB2_0_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_1/N3  ( .A1(\SB2_0_19/i1_5 ), .A2(
        \SB2_0_19/i0[6] ), .A3(\SB2_0_19/i0[9] ), .ZN(
        \SB2_0_19/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_18/Component_Function_5/N1  ( .A1(\SB2_0_18/i0_0 ), .A2(
        \SB2_0_18/i3[0] ), .ZN(\SB2_0_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_0/Component_Function_4/N1  ( .A1(\SB2_0_0/i0[9] ), .A2(
        \SB2_0_0/i0_0 ), .A3(n4003), .ZN(
        \SB2_0_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1211 ( .A1(\RI3[0][71] ), .A2(\SB2_0_20/i0[9] ), .A3(
        \SB2_0_20/i0[10] ), .ZN(\SB2_0_20/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 \SB2_0_31/Component_Function_0/N4  ( .A1(\SB2_0_31/i0[7] ), .A2(
        \SB2_0_31/i0_3 ), .A3(\SB2_0_31/i0_0 ), .ZN(
        \SB2_0_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U5851 ( .A1(n630), .A2(\SB2_0_4/i1_5 ), .A3(\SB2_0_4/i0[8] ), .ZN(
        n4198) );
  NAND3_X1 \SB2_0_2/Component_Function_3/N4  ( .A1(\SB2_0_2/i1_5 ), .A2(
        \SB2_0_2/i0[8] ), .A3(\SB2_0_2/i3[0] ), .ZN(
        \SB2_0_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_17/Component_Function_4/N3  ( .A1(\SB2_0_17/i0[9] ), .A2(
        \SB2_0_17/i0[10] ), .A3(\SB2_0_17/i0_3 ), .ZN(
        \SB2_0_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_11/Component_Function_2/N1  ( .A1(\SB2_0_11/i1_5 ), .A2(
        \SB2_0_11/i0[10] ), .A3(\SB2_0_11/i1[9] ), .ZN(
        \SB2_0_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_27/Component_Function_5/N3  ( .A1(\SB2_0_27/i1[9] ), .A2(
        \RI3[0][28] ), .A3(\SB2_0_27/i0_3 ), .ZN(
        \SB2_0_27/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1932 ( .A1(\SB2_0_12/i0[10] ), .A2(\SB2_0_12/i0[6] ), .A3(
        \RI3[0][119] ), .ZN(n5163) );
  NAND2_X1 \SB2_0_8/Component_Function_0/N1  ( .A1(\SB2_0_8/i0[10] ), .A2(
        \SB2_0_8/i0[9] ), .ZN(\SB2_0_8/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_11/Component_Function_0/N1  ( .A1(\SB2_0_11/i0[10] ), .A2(
        \SB2_0_11/i0[9] ), .ZN(\SB2_0_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_5/N3  ( .A1(\SB2_0_12/i1[9] ), .A2(
        \RI3[0][118] ), .A3(\RI3[0][119] ), .ZN(
        \SB2_0_12/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_19/Component_Function_2/N4  ( .A1(\SB2_0_19/i1_5 ), .A2(
        \SB2_0_19/i0_0 ), .A3(\RI3[0][76] ), .ZN(
        \SB2_0_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1220 ( .A1(\SB2_0_30/i0_4 ), .A2(\SB2_0_30/i0[9] ), .A3(
        \SB2_0_30/i0[6] ), .ZN(\SB2_0_30/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U9666 ( .A1(\SB2_0_7/i1[9] ), .A2(\SB2_0_7/i0_3 ), .A3(
        \SB2_0_7/i0[6] ), .ZN(\SB2_0_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_16/Component_Function_4/N2  ( .A1(\SB2_0_16/i3[0] ), .A2(
        \SB2_0_16/i0_0 ), .A3(\SB2_0_16/i1_7 ), .ZN(
        \SB2_0_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_5/Component_Function_2/N4  ( .A1(n6282), .A2(\SB2_0_5/i0_0 ), 
        .A3(\SB2_0_5/i0_4 ), .ZN(\SB2_0_5/Component_Function_2/NAND4_in[3] )
         );
  NAND2_X1 \SB2_0_3/Component_Function_5/N1  ( .A1(\SB2_0_3/i0_0 ), .A2(
        \SB2_0_3/i3[0] ), .ZN(\SB2_0_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4502 ( .A1(\SB2_0_11/i0_0 ), .A2(\SB2_0_11/i0_4 ), .A3(
        \SB2_0_11/i1_5 ), .ZN(\SB2_0_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_22/Component_Function_4/N4  ( .A1(\SB2_0_22/i1[9] ), .A2(
        \SB2_0_22/i1_5 ), .A3(\RI3[0][58] ), .ZN(
        \SB2_0_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4962 ( .A1(\SB2_0_30/i0_3 ), .A2(\SB2_0_30/i0_0 ), .A3(
        \SB2_0_30/i0_4 ), .ZN(\SB2_0_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_18/Component_Function_4/N4  ( .A1(\SB2_0_18/i1[9] ), .A2(
        \SB2_0_18/i1_5 ), .A3(\RI3[0][82] ), .ZN(
        \SB2_0_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U12447 ( .A1(\SB2_0_0/i0[10] ), .A2(\SB2_0_0/i0_0 ), .A3(
        \SB2_0_0/i0[6] ), .ZN(\SB2_0_0/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_29/Component_Function_4/N3  ( .A1(\SB2_0_29/i0[9] ), .A2(
        \SB2_0_29/i0[10] ), .A3(\SB2_0_29/i0_3 ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3569 ( .A1(\SB2_0_7/i0_0 ), .A2(\SB2_0_7/i0[7] ), .A3(
        \SB2_0_7/i0_3 ), .ZN(n1243) );
  NAND3_X1 U12663 ( .A1(\SB2_0_6/i0[8] ), .A2(\SB2_0_6/i1_7 ), .A3(
        \RI3[0][154] ), .ZN(\SB2_0_6/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 U10582 ( .A1(\SB2_0_27/i3[0] ), .A2(\SB2_0_27/i0_0 ), .ZN(n4335) );
  NAND3_X1 U2211 ( .A1(\SB2_0_16/i1_5 ), .A2(\SB2_0_16/i1[9] ), .A3(n594), 
        .ZN(\SB2_0_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_16/Component_Function_1/N2  ( .A1(\SB2_0_16/i0_3 ), .A2(
        \SB2_0_16/i1_7 ), .A3(\SB2_0_16/i0[8] ), .ZN(
        \SB2_0_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_16/Component_Function_0/N4  ( .A1(\SB2_0_16/i0[7] ), .A2(
        \SB2_0_16/i0_3 ), .A3(\SB2_0_16/i0_0 ), .ZN(
        \SB2_0_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U10947 ( .A1(\SB2_0_6/i0_4 ), .A2(\SB2_0_6/i0_3 ), .A3(
        \SB2_0_6/i0[10] ), .ZN(n4498) );
  NAND3_X1 \SB2_0_2/Component_Function_2/N3  ( .A1(\SB2_0_2/i0_3 ), .A2(
        \SB2_0_2/i0[8] ), .A3(\SB2_0_2/i0[9] ), .ZN(
        \SB2_0_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1991 ( .A1(\SB2_0_3/i0[10] ), .A2(\SB2_0_3/i0_0 ), .A3(
        \SB2_0_3/i0[6] ), .ZN(\SB2_0_3/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U7508 ( .A1(\SB2_0_6/i0_3 ), .A2(\SB2_0_6/i0[10] ), .A3(
        \SB2_0_6/i0[9] ), .ZN(\SB2_0_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U6543 ( .A1(\SB2_0_2/i0_3 ), .A2(\SB2_0_2/i0[10] ), .A3(
        \RI3[0][178] ), .ZN(\SB2_0_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1176 ( .A1(\SB2_0_0/i0_3 ), .A2(\SB2_0_0/i1[9] ), .A3(
        \RI3[0][190] ), .ZN(n1518) );
  NAND3_X1 \SB2_0_24/Component_Function_5/N4  ( .A1(\RI3[0][42] ), .A2(
        \SB2_0_24/i0[6] ), .A3(\RI3[0][46] ), .ZN(
        \SB2_0_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_16/Component_Function_4/N1  ( .A1(\SB2_0_16/i0[9] ), .A2(
        \SB2_0_16/i0_0 ), .A3(\SB2_0_16/i0[8] ), .ZN(
        \SB2_0_16/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 U3561 ( .A1(\SB2_0_7/i0_0 ), .A2(\SB2_0_7/i3[0] ), .ZN(
        \SB2_0_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U11218 ( .A1(n4003), .A2(\SB2_0_0/i1_5 ), .A3(\SB2_0_0/i3[0] ), 
        .ZN(n4620) );
  NAND3_X1 \SB2_0_29/Component_Function_1/N4  ( .A1(\SB2_0_29/i1_7 ), .A2(
        \SB2_0_29/i0[8] ), .A3(\SB2_0_29/i0_4 ), .ZN(
        \SB2_0_29/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U376 ( .I(n29), .ZN(n472) );
  INV_X1 U43 ( .I(n3), .ZN(n441) );
  BUF_X2 U2076 ( .I(Key[91]), .Z(n192) );
  BUF_X2 U196 ( .I(Key[126]), .Z(n139) );
  BUF_X2 U200 ( .I(Key[40]), .Z(n143) );
  INV_X1 U51 ( .I(n98), .ZN(n496) );
  INV_X1 U62 ( .I(n6), .ZN(n543) );
  INV_X1 U59 ( .I(n27), .ZN(n471) );
  INV_X1 U50 ( .I(n42), .ZN(n567) );
  INV_X1 U32 ( .I(n86), .ZN(n501) );
  INV_X1 U2418 ( .I(n15), .ZN(n475) );
  INV_X1 U3611 ( .I(\MC_ARK_ARC_1_0/buf_output[187] ), .ZN(\SB1_1_0/i1_7 ) );
  INV_X1 U9347 ( .I(\MC_ARK_ARC_1_0/buf_output[7] ), .ZN(\SB1_1_30/i1_7 ) );
  NAND3_X1 U6359 ( .A1(\SB1_1_3/i0_3 ), .A2(\SB1_1_3/i0_0 ), .A3(
        \SB1_1_3/i0_4 ), .ZN(\SB1_1_3/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U2148 ( .I(\SB1_1_4/i0_4 ), .ZN(\SB1_1_4/i0[7] ) );
  INV_X2 \SB1_1_0/INV_4  ( .I(\SB1_1_0/i0_4 ), .ZN(\SB1_1_0/i0[7] ) );
  NAND3_X1 U6810 ( .A1(\SB1_1_0/i0_0 ), .A2(\SB1_1_0/i0[9] ), .A3(
        \SB1_1_0/i0[8] ), .ZN(n3591) );
  INV_X1 \SB1_1_18/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[79] ), .ZN(
        \SB1_1_18/i1_7 ) );
  CLKBUF_X2 \SB1_1_0/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[187] ), .Z(
        \SB1_1_0/i0[6] ) );
  INV_X1 \SB1_1_11/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[121] ), .ZN(
        \SB1_1_11/i1_7 ) );
  INV_X1 \SB1_1_10/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[127] ), .ZN(
        \SB1_1_10/i1_7 ) );
  INV_X1 \SB1_1_6/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[152] ), .ZN(
        \SB1_1_6/i1[9] ) );
  INV_X1 \SB1_1_25/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[37] ), .ZN(
        \SB1_1_25/i1_7 ) );
  BUF_X2 \SB1_1_18/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[81] ), .Z(
        \SB1_1_18/i0[10] ) );
  INV_X1 \SB1_1_15/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[97] ), .ZN(
        \SB1_1_15/i1_7 ) );
  BUF_X2 U3613 ( .I(\MC_ARK_ARC_1_0/buf_output[42] ), .Z(\SB1_1_24/i0[9] ) );
  INV_X1 \SB1_1_4/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[163] ), .ZN(
        \SB1_1_4/i1_7 ) );
  BUF_X2 \SB1_1_27/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[25] ), .Z(
        \SB1_1_27/i0[6] ) );
  INV_X1 \SB1_1_13/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[109] ), .ZN(
        \SB1_1_13/i1_7 ) );
  AND2_X1 U3321 ( .A1(\MC_ARK_ARC_1_0/buf_output[61] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[64] ), .Z(n2355) );
  NAND3_X1 U10477 ( .A1(\SB1_1_0/i0_0 ), .A2(\SB1_1_0/i3[0] ), .A3(
        \SB1_1_0/i1_7 ), .ZN(n4996) );
  INV_X1 \SB1_1_4/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[162] ), .ZN(
        \SB1_1_4/i3[0] ) );
  INV_X1 \SB1_1_18/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[78] ), .ZN(
        \SB1_1_18/i3[0] ) );
  INV_X1 \SB1_1_29/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[12] ), .ZN(
        \SB1_1_29/i3[0] ) );
  INV_X2 U2147 ( .I(\SB1_1_10/i0_4 ), .ZN(\SB1_1_10/i0[7] ) );
  BUF_X2 \SB1_1_19/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[72] ), .Z(
        \SB1_1_19/i0[9] ) );
  BUF_X2 \SB1_1_20/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[66] ), .Z(
        \SB1_1_20/i0[9] ) );
  BUF_X2 \SB1_1_23/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[49] ), .Z(
        \SB1_1_23/i0[6] ) );
  BUF_X2 \SB1_1_28/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[19] ), .Z(
        \SB1_1_28/i0[6] ) );
  BUF_X2 \SB1_1_10/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[126] ), .Z(
        \SB1_1_10/i0[9] ) );
  CLKBUF_X2 \SB1_1_2/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[175] ), .Z(
        \SB1_1_2/i0[6] ) );
  INV_X1 \SB1_1_24/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[43] ), .ZN(
        \SB1_1_24/i1_7 ) );
  INV_X2 \SB1_1_23/INV_4  ( .I(\SB1_1_23/i0_4 ), .ZN(\SB1_1_23/i0[7] ) );
  INV_X2 \SB1_1_31/INV_4  ( .I(\SB1_1_31/i0_4 ), .ZN(\SB1_1_31/i0[7] ) );
  INV_X1 U2282 ( .I(\MC_ARK_ARC_1_0/buf_output[83] ), .ZN(\SB1_1_18/i1_5 ) );
  INV_X1 \SB1_1_19/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[77] ), .ZN(
        \SB1_1_19/i1_5 ) );
  INV_X1 \SB1_1_29/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[17] ), .ZN(
        \SB1_1_29/i1_5 ) );
  NAND3_X1 U4493 ( .A1(\SB1_1_0/i1[9] ), .A2(\SB1_1_0/i0_4 ), .A3(
        \SB1_1_0/i1_5 ), .ZN(\SB1_1_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1165 ( .A1(\SB1_1_30/i0_0 ), .A2(\SB1_1_30/i3[0] ), .A3(
        \SB1_1_30/i1_7 ), .ZN(\SB1_1_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3637 ( .A1(\SB1_1_30/i0[10] ), .A2(\SB1_1_30/i0_3 ), .A3(
        \SB1_1_30/i0[9] ), .ZN(n1922) );
  BUF_X2 \SB1_1_7/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[145] ), .Z(
        \SB1_1_7/i0[6] ) );
  BUF_X2 \SB1_1_7/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[144] ), .Z(
        \SB1_1_7/i0[9] ) );
  NAND3_X1 U1788 ( .A1(\SB1_1_2/i0[10] ), .A2(\SB1_1_2/i1[9] ), .A3(
        \SB1_1_2/i1_5 ), .ZN(\SB1_1_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_3/N2  ( .A1(\SB1_1_28/i0_0 ), .A2(
        \SB1_1_28/i0_3 ), .A3(\SB1_1_28/i0_4 ), .ZN(
        \SB1_1_28/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_11/Component_Function_0/N1  ( .A1(\SB1_1_11/i0[10] ), .A2(
        \SB1_1_11/i0[9] ), .ZN(\SB1_1_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_2/N3  ( .A1(\SB1_1_15/i0_3 ), .A2(
        \SB1_1_15/i0[8] ), .A3(\SB1_1_15/i0[9] ), .ZN(
        \SB1_1_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4354 ( .A1(\SB1_1_15/i0[10] ), .A2(\SB1_1_15/i1[9] ), .A3(
        \SB1_1_15/i1_7 ), .ZN(\SB1_1_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_5/Component_Function_2/N3  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i0[8] ), .A3(\SB1_1_5/i0[9] ), .ZN(
        \SB1_1_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_19/Component_Function_2/N3  ( .A1(\SB1_1_19/i0_3 ), .A2(
        \SB1_1_19/i0[8] ), .A3(\SB1_1_19/i0[9] ), .ZN(
        \SB1_1_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1852 ( .A1(\SB1_1_9/i0[10] ), .A2(\SB1_1_9/i0_3 ), .A3(
        \SB1_1_9/i0_4 ), .ZN(n4956) );
  NAND3_X1 U8331 ( .A1(\SB1_1_13/i0_3 ), .A2(\SB1_1_13/i0_4 ), .A3(
        \SB1_1_13/i1[9] ), .ZN(\SB1_1_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_4/Component_Function_2/N3  ( .A1(\SB1_1_4/i0_3 ), .A2(
        \SB1_1_4/i0[8] ), .A3(\SB1_1_4/i0[9] ), .ZN(
        \SB1_1_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U6510 ( .A1(\SB1_1_7/i0[9] ), .A2(\SB1_1_7/i0_3 ), .A3(
        \SB1_1_7/i0[10] ), .ZN(n3553) );
  NAND3_X1 U1105 ( .A1(\SB1_1_28/i0[10] ), .A2(\SB1_1_28/i1[9] ), .A3(
        \SB1_1_28/i1_7 ), .ZN(n1717) );
  NAND3_X1 U3167 ( .A1(\SB1_1_0/i0_0 ), .A2(\SB1_1_0/i0_4 ), .A3(
        \SB1_1_0/i1_5 ), .ZN(\SB1_1_0/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U6328 ( .A1(\SB1_1_6/i0[8] ), .A2(\SB1_1_6/i3[0] ), .A3(
        \SB1_1_6/i1_5 ), .ZN(n1883) );
  NAND3_X1 U1120 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i0_3 ), .A3(
        \SB1_1_2/i0[7] ), .ZN(n2928) );
  NAND3_X1 \SB1_1_14/Component_Function_0/N2  ( .A1(\SB1_1_14/i0[8] ), .A2(
        \SB1_1_14/i0[7] ), .A3(\SB1_1_14/i0[6] ), .ZN(
        \SB1_1_14/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1855 ( .A1(\SB1_1_31/i0[8] ), .A2(\SB1_1_31/i1_5 ), .A3(
        \SB1_1_31/i3[0] ), .ZN(\SB1_1_31/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_17/Component_Function_5/N1  ( .A1(\SB1_1_17/i0_0 ), .A2(
        \SB1_1_17/i3[0] ), .ZN(\SB1_1_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_3/N3  ( .A1(\SB1_1_25/i1[9] ), .A2(
        \SB1_1_25/i1_7 ), .A3(\SB1_1_25/i0[10] ), .ZN(
        \SB1_1_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_25/Component_Function_1/N4  ( .A1(\SB1_1_25/i1_7 ), .A2(
        \SB1_1_25/i0[8] ), .A3(\SB1_1_25/i0_4 ), .ZN(
        \SB1_1_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_10/Component_Function_1/N4  ( .A1(\SB1_1_10/i1_7 ), .A2(
        \SB1_1_10/i0[8] ), .A3(\SB1_1_10/i0_4 ), .ZN(
        \SB1_1_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1156 ( .A1(\SB1_1_1/i0_3 ), .A2(\SB1_1_1/i0_4 ), .A3(
        \SB1_1_1/i1[9] ), .ZN(\SB1_1_1/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_13/Component_Function_5/N1  ( .A1(\SB1_1_13/i0_0 ), .A2(
        \SB1_1_13/i3[0] ), .ZN(\SB1_1_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1133 ( .A1(\SB1_1_20/i0[10] ), .A2(\SB1_1_20/i1[9] ), .A3(
        \SB1_1_20/i1_7 ), .ZN(\SB1_1_20/Component_Function_3/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_22/Component_Function_5/N1  ( .A1(\SB1_1_22/i0_0 ), .A2(
        \SB1_1_22/i3[0] ), .ZN(\SB1_1_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U6219 ( .A1(\SB1_1_24/i0[10] ), .A2(\SB1_1_24/i1[9] ), .A3(
        \SB1_1_24/i1_7 ), .ZN(n1833) );
  NAND3_X1 U4245 ( .A1(\SB1_1_20/i0[8] ), .A2(\SB1_1_20/i3[0] ), .A3(
        \SB1_1_20/i1_5 ), .ZN(\SB1_1_20/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_21/Component_Function_1/N1  ( .A1(\SB1_1_21/i0_3 ), .A2(
        \SB1_1_21/i1[9] ), .ZN(\SB1_1_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_1/N3  ( .A1(\SB1_1_20/i1_5 ), .A2(
        \SB1_1_20/i0[6] ), .A3(\SB1_1_20/i0[9] ), .ZN(
        \SB1_1_20/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_15/Component_Function_5/N1  ( .A1(\SB1_1_15/i0_0 ), .A2(
        \SB1_1_15/i3[0] ), .ZN(\SB1_1_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U6401 ( .A1(\SB1_1_26/i0_4 ), .A2(\SB1_1_26/i0[9] ), .A3(
        \SB1_1_26/i0[6] ), .ZN(n4683) );
  NAND3_X1 U10134 ( .A1(\SB1_1_18/i0[6] ), .A2(\SB1_1_18/i0_3 ), .A3(
        \SB1_1_18/i1[9] ), .ZN(n1892) );
  NAND3_X1 \SB1_1_15/Component_Function_1/N3  ( .A1(\SB1_1_15/i1_5 ), .A2(
        \SB1_1_15/i0[6] ), .A3(\SB1_1_15/i0[9] ), .ZN(
        \SB1_1_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_4/Component_Function_1/N3  ( .A1(\SB1_1_4/i1_5 ), .A2(
        \SB1_1_4/i0[6] ), .A3(\SB1_1_4/i0[9] ), .ZN(
        \SB1_1_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U11485 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i1[9] ), .A3(
        \SB1_1_15/i0[6] ), .ZN(n4752) );
  NAND3_X1 U3049 ( .A1(\SB1_1_11/i0_3 ), .A2(\SB1_1_11/i1[9] ), .A3(
        \SB1_1_11/i0_4 ), .ZN(n4427) );
  NAND3_X1 \SB1_1_10/Component_Function_1/N3  ( .A1(\SB1_1_10/i1_5 ), .A2(
        \SB1_1_10/i0[6] ), .A3(\SB1_1_10/i0[9] ), .ZN(
        \SB1_1_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2177 ( .A1(\SB1_1_22/i1_7 ), .A2(\SB1_1_22/i0[8] ), .A3(
        \SB1_1_22/i0_4 ), .ZN(\SB1_1_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4445 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0[8] ), .A3(
        \SB1_1_20/i0[9] ), .ZN(\SB1_1_20/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_3/Component_Function_1/N1  ( .A1(\SB1_1_3/i0_3 ), .A2(
        \SB1_1_3/i1[9] ), .ZN(\SB1_1_3/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_31/Component_Function_1/N1  ( .A1(\SB1_1_31/i0_3 ), .A2(
        \SB1_1_31/i1[9] ), .ZN(\SB1_1_31/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_15/Component_Function_1/N1  ( .A1(\SB1_1_15/i0_3 ), .A2(
        \SB1_1_15/i1[9] ), .ZN(\SB1_1_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U7563 ( .A1(\SB1_1_15/i0_0 ), .A2(\SB1_1_15/i1_5 ), .A3(
        \SB1_1_15/i0_4 ), .ZN(n2455) );
  NAND2_X1 \SB1_1_26/Component_Function_5/N1  ( .A1(\SB1_1_26/i0_0 ), .A2(
        \SB1_1_26/i3[0] ), .ZN(\SB1_1_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_5/N4  ( .A1(\SB1_1_31/i0[9] ), .A2(
        \SB1_1_31/i0[6] ), .A3(\SB1_1_31/i0_4 ), .ZN(
        \SB1_1_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_18/Component_Function_5/N2  ( .A1(\SB1_1_18/i0_0 ), .A2(
        \SB1_1_18/i0[6] ), .A3(\SB1_1_18/i0[10] ), .ZN(
        \SB1_1_18/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U12046 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i0[10] ), .A3(
        \SB1_1_10/i0[9] ), .ZN(\SB1_1_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1837 ( .A1(\SB1_1_29/i0_4 ), .A2(\SB1_1_29/i0[9] ), .A3(
        \SB1_1_29/i0[6] ), .ZN(n4596) );
  NAND3_X1 \SB1_1_2/Component_Function_4/N3  ( .A1(\SB1_1_2/i0[9] ), .A2(
        \SB1_1_2/i0[10] ), .A3(\SB1_1_2/i0_3 ), .ZN(
        \SB1_1_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2170 ( .A1(\SB1_1_2/i0[10] ), .A2(\SB1_1_2/i0_4 ), .A3(
        \SB1_1_2/i0_3 ), .ZN(\SB1_1_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_13/Component_Function_1/N3  ( .A1(\SB1_1_13/i1_5 ), .A2(
        \SB1_1_13/i0[6] ), .A3(\SB1_1_13/i0[9] ), .ZN(
        \SB1_1_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U11151 ( .A1(\SB1_1_27/i0[6] ), .A2(\SB1_1_27/i0_0 ), .A3(
        \SB1_1_27/i0[10] ), .ZN(\SB1_1_27/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U1153 ( .A1(\SB1_1_4/i0_3 ), .A2(\SB1_1_4/i1[9] ), .A3(
        \SB1_1_4/i0_4 ), .ZN(n2588) );
  NAND3_X1 U6076 ( .A1(\SB1_1_12/i0[10] ), .A2(\SB1_1_12/i0[6] ), .A3(
        \SB1_1_12/i0_0 ), .ZN(\SB1_1_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U12048 ( .A1(\SB1_1_18/i0[9] ), .A2(\SB1_1_18/i0[6] ), .A3(
        \SB1_1_18/i0_4 ), .ZN(n5053) );
  NAND3_X1 \SB1_1_29/Component_Function_3/N2  ( .A1(\SB1_1_29/i0_0 ), .A2(
        \SB1_1_29/i0_3 ), .A3(\SB1_1_29/i0_4 ), .ZN(
        \SB1_1_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U7415 ( .A1(\SB1_1_24/i1_5 ), .A2(\SB1_1_24/i0_4 ), .A3(
        \SB1_1_24/i0_0 ), .ZN(n2380) );
  INV_X2 \SB1_1_8/INV_4  ( .I(\SB1_1_8/i0_4 ), .ZN(\SB1_1_8/i0[7] ) );
  NAND3_X1 \SB1_1_4/Component_Function_3/N1  ( .A1(\SB1_1_4/i1[9] ), .A2(
        \SB1_1_4/i0_3 ), .A3(\SB1_1_4/i0[6] ), .ZN(
        \SB1_1_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U8523 ( .A1(\SB1_1_0/i0[8] ), .A2(\SB1_1_0/i3[0] ), .A3(
        \SB1_1_0/i1_5 ), .ZN(n2496) );
  NAND3_X1 U1858 ( .A1(\SB1_1_16/i0_4 ), .A2(\SB1_1_16/i0[8] ), .A3(
        \SB1_1_16/i1_7 ), .ZN(n4114) );
  NAND3_X1 U6597 ( .A1(\SB1_1_1/i0_0 ), .A2(\SB1_1_1/i0_4 ), .A3(
        \SB1_1_1/i1_5 ), .ZN(\SB1_1_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1154 ( .A1(\SB1_1_25/i0[9] ), .A2(\SB1_1_25/i1_5 ), .A3(
        \SB1_1_25/i0[6] ), .ZN(\SB1_1_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1127 ( .A1(\SB1_1_1/i0[6] ), .A2(\SB1_1_1/i1[9] ), .A3(
        \SB1_1_1/i0_3 ), .ZN(n2861) );
  NAND3_X1 \SB1_1_7/Component_Function_3/N2  ( .A1(\SB1_1_7/i0_0 ), .A2(
        \SB1_1_7/i0_3 ), .A3(\SB1_1_7/i0_4 ), .ZN(
        \SB1_1_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U8244 ( .A1(\SB1_1_4/i0[9] ), .A2(\SB1_1_4/i0_4 ), .A3(
        \SB1_1_4/i0[6] ), .ZN(n2826) );
  NAND3_X1 U1724 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i0_0 ), .A3(
        \SB1_1_26/i0[6] ), .ZN(\SB1_1_26/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_2/Component_Function_1/N4  ( .A1(\SB1_1_2/i1_7 ), .A2(
        \SB1_1_2/i0[8] ), .A3(\SB1_1_2/i0_4 ), .ZN(
        \SB1_1_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U12266 ( .A1(\SB1_1_9/i0_3 ), .A2(\SB1_1_9/i0_4 ), .A3(
        \SB1_1_9/i1[9] ), .ZN(\SB1_1_9/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U11055 ( .A1(\SB1_1_15/i0[10] ), .A2(\SB1_1_15/i0_0 ), .A3(
        \SB1_1_15/i0[6] ), .ZN(\SB1_1_15/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_13/Component_Function_0/N4  ( .A1(\SB1_1_13/i0[7] ), .A2(
        \SB1_1_13/i0_3 ), .A3(\SB1_1_13/i0_0 ), .ZN(
        \SB1_1_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1697 ( .A1(\SB1_1_25/i0_3 ), .A2(\SB1_1_25/i0_0 ), .A3(
        \SB1_1_25/i0[7] ), .ZN(n3191) );
  NAND3_X1 \SB1_1_9/Component_Function_4/N3  ( .A1(\SB1_1_9/i0[9] ), .A2(
        \SB1_1_9/i0[10] ), .A3(\SB1_1_9/i0_3 ), .ZN(
        \SB1_1_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3054 ( .A1(\SB1_1_11/i0[9] ), .A2(\SB1_1_11/i0[10] ), .A3(
        \SB1_1_11/i0_3 ), .ZN(\SB1_1_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1747 ( .A1(\SB1_1_29/i0_4 ), .A2(\SB1_1_29/i1[9] ), .A3(
        \SB1_1_29/i1_5 ), .ZN(n3747) );
  NAND3_X1 \SB1_1_7/Component_Function_1/N4  ( .A1(\SB1_1_7/i1_7 ), .A2(
        \SB1_1_7/i0[8] ), .A3(\SB1_1_7/i0_4 ), .ZN(
        \SB1_1_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_5/Component_Function_3/N2  ( .A1(\SB1_1_5/i0_0 ), .A2(
        \SB1_1_5/i0_3 ), .A3(\SB1_1_5/i0_4 ), .ZN(
        \SB1_1_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U9770 ( .A1(\SB1_1_30/i0[10] ), .A2(\SB1_1_30/i1[9] ), .A3(
        \SB1_1_30/i1_7 ), .ZN(n5132) );
  NAND3_X1 \SB1_1_26/Component_Function_4/N4  ( .A1(\SB1_1_26/i1[9] ), .A2(
        \SB1_1_26/i1_5 ), .A3(\SB1_1_26/i0_4 ), .ZN(
        \SB1_1_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_2/N3  ( .A1(\SB1_1_27/i0_3 ), .A2(
        \SB1_1_27/i0[8] ), .A3(\SB1_1_27/i0[9] ), .ZN(
        \SB1_1_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_28/Component_Function_2/N4  ( .A1(\SB1_1_28/i1_5 ), .A2(
        \SB1_1_28/i0_0 ), .A3(\SB1_1_28/i0_4 ), .ZN(
        \SB1_1_28/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_28/Component_Function_2/N3  ( .A1(\SB1_1_28/i0_3 ), .A2(
        \SB1_1_28/i0[8] ), .A3(\SB1_1_28/i0[9] ), .ZN(
        \SB1_1_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U8184 ( .A1(\SB1_1_14/i0[8] ), .A2(\SB1_1_14/i1_7 ), .A3(
        \SB1_1_14/i0_4 ), .ZN(n3833) );
  NAND3_X1 U7530 ( .A1(\SB1_1_0/i0_4 ), .A2(\SB1_1_0/i0[8] ), .A3(
        \SB1_1_0/i1_7 ), .ZN(\SB1_1_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_25/Component_Function_0/N2  ( .A1(\SB1_1_25/i0[8] ), .A2(
        \SB1_1_25/i0[7] ), .A3(\SB1_1_25/i0[6] ), .ZN(
        \SB1_1_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U12575 ( .A1(\SB1_1_29/i0_0 ), .A2(\SB1_1_29/i0[7] ), .A3(
        \SB1_1_29/i0_3 ), .ZN(n5348) );
  NAND3_X1 \SB1_1_14/Component_Function_1/N3  ( .A1(\SB1_1_14/i1_5 ), .A2(
        \SB1_1_14/i0[6] ), .A3(\SB1_1_14/i0[9] ), .ZN(
        \SB1_1_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_18/Component_Function_1/N2  ( .A1(\SB1_1_18/i0_3 ), .A2(
        \SB1_1_18/i1_7 ), .A3(\SB1_1_18/i0[8] ), .ZN(
        \SB1_1_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1704 ( .A1(\SB1_1_19/i0[9] ), .A2(\SB1_1_19/i0_4 ), .A3(
        \SB1_1_19/i0[6] ), .ZN(n5251) );
  NAND3_X1 U7000 ( .A1(\SB1_1_15/i0[10] ), .A2(\SB1_1_15/i0_3 ), .A3(
        \SB1_1_15/i0_4 ), .ZN(n2196) );
  NAND2_X1 \SB1_1_7/Component_Function_1/N1  ( .A1(\SB1_1_7/i0_3 ), .A2(
        \SB1_1_7/i1[9] ), .ZN(\SB1_1_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_4/N1  ( .A1(\SB1_1_15/i0[9] ), .A2(
        \SB1_1_15/i0_0 ), .A3(\SB1_1_15/i0[8] ), .ZN(
        \SB1_1_15/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_24/Component_Function_1/N1  ( .A1(\RI1[1][47] ), .A2(
        \SB1_1_24/i1[9] ), .ZN(\SB1_1_24/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 U1716 ( .A1(n4984), .A2(n2801), .ZN(n4102) );
  NAND3_X1 \SB1_1_12/Component_Function_1/N3  ( .A1(\SB1_1_12/i1_5 ), .A2(
        \SB1_1_12/i0[6] ), .A3(\SB1_1_12/i0[9] ), .ZN(
        \SB1_1_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_21/Component_Function_3/N1  ( .A1(\SB1_1_21/i1[9] ), .A2(
        \SB1_1_21/i0_3 ), .A3(\SB1_1_21/i0[6] ), .ZN(
        \SB1_1_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U6406 ( .A1(\SB1_1_8/i0[10] ), .A2(\SB1_1_8/i0_0 ), .A3(
        \SB1_1_8/i0[6] ), .ZN(\SB1_1_8/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_24/Component_Function_1/N3  ( .A1(\SB1_1_24/i1_5 ), .A2(
        \SB1_1_24/i0[6] ), .A3(\SB1_1_24/i0[9] ), .ZN(
        \SB1_1_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_20/Component_Function_5/N2  ( .A1(\SB1_1_20/i0_0 ), .A2(
        \SB1_1_20/i0[6] ), .A3(\SB1_1_20/i0[10] ), .ZN(
        \SB1_1_20/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X2 \SB2_1_1/BUF_0  ( .I(\SB1_1_6/buf_output[0] ), .Z(\SB2_1_1/i0[9] )
         );
  BUF_X2 \SB2_1_1/BUF_1  ( .I(\SB1_1_5/buf_output[1] ), .Z(\SB2_1_1/i0[6] ) );
  NAND3_X1 U1781 ( .A1(\SB1_1_27/i0[10] ), .A2(\SB1_1_27/i1_7 ), .A3(
        \SB1_1_27/i1[9] ), .ZN(n4067) );
  NAND3_X1 U8198 ( .A1(\SB1_1_5/i0[10] ), .A2(\SB1_1_5/i0[9] ), .A3(
        \SB1_1_5/i0_3 ), .ZN(\SB1_1_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_27/Component_Function_3/N4  ( .A1(\SB1_1_27/i1_5 ), .A2(
        \SB1_1_27/i0[8] ), .A3(\SB1_1_27/i3[0] ), .ZN(
        \SB1_1_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_3/N1  ( .A1(\SB1_1_27/i1[9] ), .A2(
        \SB1_1_27/i0_3 ), .A3(\SB1_1_27/i0[6] ), .ZN(
        \SB1_1_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U8871 ( .A1(\SB1_1_25/i0[10] ), .A2(\SB1_1_25/i0_0 ), .A3(
        \SB1_1_25/i0[6] ), .ZN(\SB1_1_25/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_28/Component_Function_5/N2  ( .A1(\SB1_1_28/i0_0 ), .A2(
        \SB1_1_28/i0[6] ), .A3(\SB1_1_28/i0[10] ), .ZN(
        \SB1_1_28/Component_Function_5/NAND4_in[1] ) );
  BUF_X2 \SB2_1_29/BUF_1  ( .I(\SB1_1_1/buf_output[1] ), .Z(\SB2_1_29/i0[6] )
         );
  CLKBUF_X2 \SB2_1_23/BUF_0  ( .I(\SB1_1_28/buf_output[0] ), .Z(
        \SB2_1_23/i0[9] ) );
  CLKBUF_X2 \SB2_1_30/BUF_0  ( .I(\SB1_1_3/buf_output[0] ), .Z(
        \SB2_1_30/i0[9] ) );
  CLKBUF_X2 \SB2_1_5/BUF_0  ( .I(\SB1_1_10/buf_output[0] ), .Z(\SB2_1_5/i0[9] ) );
  BUF_X2 U3746 ( .I(\SB1_1_6/buf_output[1] ), .Z(\SB2_1_2/i0[6] ) );
  BUF_X2 \SB2_1_16/BUF_1  ( .I(\SB1_1_20/buf_output[1] ), .Z(\SB2_1_16/i0[6] )
         );
  INV_X1 \SB2_1_23/INV_0  ( .I(\SB1_1_28/buf_output[0] ), .ZN(\SB2_1_23/i3[0] ) );
  NAND2_X1 \SB2_1_26/Component_Function_5/N1  ( .A1(\SB2_1_26/i0_0 ), .A2(
        \SB2_1_26/i3[0] ), .ZN(\SB2_1_26/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_17/Component_Function_5/N1  ( .A1(\SB2_1_17/i0_0 ), .A2(
        \SB2_1_17/i3[0] ), .ZN(\SB2_1_17/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_13/Component_Function_5/N1  ( .A1(\SB2_1_13/i0_0 ), .A2(
        \SB2_1_13/i3[0] ), .ZN(\SB2_1_13/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U4064 ( .A1(\SB2_1_12/i0_0 ), .A2(\SB2_1_12/i3[0] ), .ZN(n1148) );
  NAND2_X1 U2187 ( .A1(\SB2_1_23/i0_0 ), .A2(\SB2_1_23/i3[0] ), .ZN(
        \SB2_1_23/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_2/Component_Function_5/N1  ( .A1(\SB2_1_2/i0_0 ), .A2(
        \SB2_1_2/i3[0] ), .ZN(\SB2_1_2/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_30/Component_Function_5/N1  ( .A1(\SB2_1_30/i0_0 ), .A2(
        \SB2_1_30/i3[0] ), .ZN(\SB2_1_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U12151 ( .A1(\SB2_1_22/i0[10] ), .A2(\SB2_1_22/i0_0 ), .A3(
        \SB2_1_22/i0[6] ), .ZN(\SB2_1_22/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3779 ( .A1(\SB2_1_17/i0_4 ), .A2(\SB2_1_17/i0_3 ), .A3(
        \SB2_1_17/i1[9] ), .ZN(\SB2_1_17/Component_Function_5/NAND4_in[2] ) );
  INV_X1 \SB2_1_16/INV_1  ( .I(\SB1_1_20/buf_output[1] ), .ZN(\SB2_1_16/i1_7 )
         );
  INV_X1 \SB2_1_28/INV_1  ( .I(\SB1_1_0/buf_output[1] ), .ZN(\SB2_1_28/i1_7 )
         );
  INV_X1 \SB2_1_6/INV_1  ( .I(\SB1_1_10/buf_output[1] ), .ZN(\SB2_1_6/i1_7 )
         );
  CLKBUF_X2 \SB2_1_25/BUF_1  ( .I(\SB1_1_29/buf_output[1] ), .Z(
        \SB2_1_25/i0[6] ) );
  BUF_X2 U9705 ( .I(\SB1_1_1/buf_output[0] ), .Z(\SB2_1_28/i0[9] ) );
  BUF_X2 \SB2_1_24/BUF_1  ( .I(\SB1_1_28/buf_output[1] ), .Z(\SB2_1_24/i0[6] )
         );
  INV_X2 U1078 ( .I(\SB2_1_19/i0[7] ), .ZN(\SB2_1_19/i0_4 ) );
  INV_X1 \SB2_1_10/INV_1  ( .I(\SB1_1_14/buf_output[1] ), .ZN(\SB2_1_10/i1_7 )
         );
  INV_X1 \SB2_1_30/INV_1  ( .I(\SB1_1_2/buf_output[1] ), .ZN(\SB2_1_30/i1_7 )
         );
  INV_X1 U2183 ( .I(\SB1_1_25/buf_output[1] ), .ZN(\SB2_1_21/i1_7 ) );
  INV_X1 \SB2_1_31/INV_3  ( .I(\SB1_1_1/buf_output[3] ), .ZN(\SB2_1_31/i0[8] )
         );
  INV_X1 \SB2_1_27/INV_1  ( .I(\SB1_1_31/buf_output[1] ), .ZN(\SB2_1_27/i1_7 )
         );
  NAND3_X1 \SB2_1_0/Component_Function_4/N1  ( .A1(\SB2_1_0/i0[9] ), .A2(
        \SB2_1_0/i0_0 ), .A3(\SB2_1_0/i0[8] ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1054 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0[10] ), .A3(
        \SB2_1_24/i0[9] ), .ZN(\SB2_1_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U12496 ( .A1(\SB2_1_11/i0_3 ), .A2(\SB2_1_11/i0[9] ), .A3(
        \SB2_1_11/i0[10] ), .ZN(\SB2_1_11/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1655 ( .A1(\SB2_1_1/i1_5 ), .A2(\SB2_1_1/i0[8] ), .A3(
        \SB2_1_1/i3[0] ), .ZN(\SB2_1_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1688 ( .A1(\SB2_1_28/i0[9] ), .A2(\SB2_1_28/i0_3 ), .A3(
        \SB2_1_28/i0[10] ), .ZN(\SB2_1_28/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 \SB2_1_8/Component_Function_2/N2  ( .A1(\SB2_1_8/i0_3 ), .A2(
        \SB2_1_8/i0[10] ), .A3(\SB2_1_8/i0[6] ), .ZN(
        \SB2_1_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U6581 ( .A1(\SB2_1_21/i0_3 ), .A2(\SB2_1_21/i0[10] ), .A3(
        \SB2_1_21/i0[9] ), .ZN(\SB2_1_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1639 ( .A1(\SB2_1_1/i0_3 ), .A2(\SB2_1_1/i0_4 ), .A3(
        \SB2_1_1/i0_0 ), .ZN(n4597) );
  NAND3_X1 U1651 ( .A1(\SB2_1_18/i1_7 ), .A2(\SB2_1_18/i0[8] ), .A3(
        \SB2_1_18/i0_4 ), .ZN(\SB2_1_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U12219 ( .A1(\SB2_1_12/i0[10] ), .A2(\SB2_1_12/i1_7 ), .A3(
        \SB2_1_12/i1[9] ), .ZN(n5298) );
  NAND3_X1 U1669 ( .A1(\SB2_1_19/i0_0 ), .A2(\SB2_1_19/i0_3 ), .A3(n5883), 
        .ZN(n5289) );
  NAND3_X1 \SB2_1_10/Component_Function_0/N2  ( .A1(\SB2_1_10/i0[8] ), .A2(
        \SB2_1_10/i0[7] ), .A3(\SB2_1_10/i0[6] ), .ZN(
        \SB2_1_10/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U7400 ( .A1(\SB2_1_13/i0_4 ), .A2(\SB2_1_13/i0_0 ), .A3(
        \SB2_1_13/i1_5 ), .ZN(n3660) );
  NAND3_X1 \SB2_1_18/Component_Function_1/N3  ( .A1(\SB2_1_18/i1_5 ), .A2(
        \SB2_1_18/i0[6] ), .A3(\SB2_1_18/i0[9] ), .ZN(
        \SB2_1_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4031 ( .A1(\SB2_1_16/i3[0] ), .A2(\SB2_1_16/i1_5 ), .A3(
        \SB2_1_16/i0[8] ), .ZN(n1210) );
  NAND3_X1 \SB2_1_30/Component_Function_1/N4  ( .A1(\SB2_1_30/i1_7 ), .A2(
        \SB2_1_30/i0[8] ), .A3(\SB2_1_30/i0_4 ), .ZN(
        \SB2_1_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U6979 ( .A1(\SB2_1_12/i0_0 ), .A2(\SB2_1_12/i0[7] ), .A3(
        \SB2_1_12/i0_3 ), .ZN(\SB2_1_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_28/Component_Function_4/N4  ( .A1(\SB2_1_28/i1[9] ), .A2(
        \SB2_1_28/i1_5 ), .A3(\SB2_1_28/i0_4 ), .ZN(
        \SB2_1_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U11655 ( .A1(\SB2_1_26/i0[10] ), .A2(\SB2_1_26/i1_7 ), .A3(
        \SB2_1_26/i1[9] ), .ZN(\SB2_1_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_9/Component_Function_3/N4  ( .A1(\SB2_1_9/i1_5 ), .A2(
        \SB2_1_9/i0[8] ), .A3(\SB2_1_9/i3[0] ), .ZN(
        \SB2_1_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U7566 ( .A1(\SB2_1_19/i0[6] ), .A2(n5883), .A3(\SB2_1_19/i0[8] ), 
        .ZN(\SB2_1_19/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_13/Component_Function_4/N4  ( .A1(\SB2_1_13/i1[9] ), .A2(
        \SB2_1_13/i1_5 ), .A3(\SB2_1_13/i0_4 ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_24/Component_Function_5/N1  ( .A1(\SB2_1_24/i0_0 ), .A2(
        \SB2_1_24/i3[0] ), .ZN(\SB2_1_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_16/Component_Function_3/N1  ( .A1(\SB2_1_16/i1[9] ), .A2(
        \SB2_1_16/i0_3 ), .A3(\SB2_1_16/i0[6] ), .ZN(
        \SB2_1_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_4/N1  ( .A1(\SB2_1_6/i0[9] ), .A2(
        \SB2_1_6/i0_0 ), .A3(\SB2_1_6/i0[8] ), .ZN(
        \SB2_1_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_2/N1  ( .A1(\SB2_1_5/i1_5 ), .A2(
        \SB2_1_5/i0[10] ), .A3(\SB2_1_5/i1[9] ), .ZN(
        \SB2_1_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_2/N1  ( .A1(n3990), .A2(
        \SB2_1_17/i0[10] ), .A3(\SB2_1_17/i1[9] ), .ZN(
        \SB2_1_17/Component_Function_2/NAND4_in[0] ) );
  INV_X1 \SB2_1_5/INV_4  ( .I(\SB1_1_6/buf_output[4] ), .ZN(\SB2_1_5/i0[7] )
         );
  NAND3_X1 \SB2_1_14/Component_Function_1/N2  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i1_7 ), .A3(\SB2_1_14/i0[8] ), .ZN(
        \SB2_1_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_2/Component_Function_2/N4  ( .A1(\SB2_1_2/i1_5 ), .A2(
        \SB2_1_2/i0_0 ), .A3(\SB2_1_2/i0_4 ), .ZN(
        \SB2_1_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_4/Component_Function_2/N1  ( .A1(\SB2_1_4/i1_5 ), .A2(
        \SB2_1_4/i0[10] ), .A3(\SB2_1_4/i1[9] ), .ZN(
        \SB2_1_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_9/Component_Function_1/N4  ( .A1(\SB2_1_9/i1_7 ), .A2(
        \SB2_1_9/i0[8] ), .A3(\SB2_1_9/i0_4 ), .ZN(
        \SB2_1_9/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_6/Component_Function_0/N1  ( .A1(\SB2_1_6/i0[10] ), .A2(
        \SB2_1_6/i0[9] ), .ZN(\SB2_1_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U7936 ( .A1(\SB2_1_16/i0[9] ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i0[8] ), .ZN(\SB2_1_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2191 ( .A1(\SB2_1_12/i1_5 ), .A2(\SB2_1_12/i0[8] ), .A3(
        \SB2_1_12/i3[0] ), .ZN(\SB2_1_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4945 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i1[9] ), .A3(
        \SB2_1_9/i0[6] ), .ZN(\SB2_1_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_2/N2  ( .A1(\SB2_1_17/i0_3 ), .A2(
        \SB2_1_17/i0[10] ), .A3(\SB2_1_17/i0[6] ), .ZN(
        \SB2_1_17/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_10/Component_Function_1/N1  ( .A1(\SB2_1_10/i0_3 ), .A2(
        \SB2_1_10/i1[9] ), .ZN(\SB2_1_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_20/Component_Function_4/N1  ( .A1(\SB2_1_20/i0[9] ), .A2(
        \SB2_1_20/i0_0 ), .A3(\SB2_1_20/i0[8] ), .ZN(
        \SB2_1_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U4706 ( .A1(\SB2_1_10/i0_0 ), .A2(\SB2_1_10/i0_3 ), .A3(
        \SB2_1_10/i0[7] ), .ZN(\SB2_1_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_20/Component_Function_4/N4  ( .A1(\SB2_1_20/i1[9] ), .A2(
        \SB2_1_20/i1_5 ), .A3(\SB2_1_20/i0_4 ), .ZN(
        \SB2_1_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1064 ( .A1(\SB2_1_23/i0_0 ), .A2(\SB2_1_23/i0_4 ), .A3(
        \SB2_1_23/i1_5 ), .ZN(n1838) );
  NAND3_X1 \SB2_1_9/Component_Function_1/N3  ( .A1(\SB2_1_9/i1_5 ), .A2(
        \SB2_1_9/i0[6] ), .A3(\SB2_1_9/i0[9] ), .ZN(
        \SB2_1_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4188 ( .A1(\SB2_1_16/i0_4 ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i0_0 ), .ZN(n1211) );
  INV_X2 U2181 ( .I(\SB2_1_8/i0_4 ), .ZN(\SB2_1_8/i0[7] ) );
  NAND3_X1 U3696 ( .A1(\SB2_1_8/i0_3 ), .A2(\SB2_1_8/i0[10] ), .A3(
        \SB2_1_8/i0[9] ), .ZN(\SB2_1_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_13/Component_Function_4/N2  ( .A1(\SB2_1_13/i3[0] ), .A2(
        \SB2_1_13/i0_0 ), .A3(\SB2_1_13/i1_7 ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_19/Component_Function_4/N2  ( .A1(\SB2_1_19/i3[0] ), .A2(
        \SB2_1_19/i0_0 ), .A3(\SB2_1_19/i1_7 ), .ZN(
        \SB2_1_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4333 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0[8] ), .A3(
        \SB2_1_10/i1_7 ), .ZN(n1359) );
  NAND3_X1 U2174 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i0[10] ), .A3(
        \SB2_1_15/i0_4 ), .ZN(\SB2_1_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U6949 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0[9] ), .A3(
        \SB2_1_24/i0[8] ), .ZN(\SB2_1_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_4/Component_Function_1/N2  ( .A1(\SB2_1_4/i0_3 ), .A2(n2656), 
        .A3(\SB2_1_4/i0[8] ), .ZN(\SB2_1_4/Component_Function_1/NAND4_in[1] )
         );
  NAND3_X1 U12178 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i0[10] ), .A3(
        \SB2_1_5/i0[9] ), .ZN(\SB2_1_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_24/Component_Function_3/N1  ( .A1(\SB2_1_24/i1[9] ), .A2(
        \SB2_1_24/i0_3 ), .A3(\SB2_1_24/i0[6] ), .ZN(
        \SB2_1_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_3/N1  ( .A1(\SB2_1_23/i1[9] ), .A2(
        \SB2_1_23/i0_3 ), .A3(\SB2_1_23/i0[6] ), .ZN(
        \SB2_1_23/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_19/Component_Function_1/N1  ( .A1(\SB2_1_19/i0_3 ), .A2(
        \SB2_1_19/i1[9] ), .ZN(\SB2_1_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_3/Component_Function_0/N4  ( .A1(\SB2_1_3/i0[7] ), .A2(
        \SB2_1_3/i0_3 ), .A3(\SB2_1_3/i0_0 ), .ZN(
        \SB2_1_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1043 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0[10] ), .A3(
        \SB2_1_9/i0_4 ), .ZN(n2270) );
  NAND3_X1 \SB2_1_29/Component_Function_3/N4  ( .A1(\SB2_1_29/i1_5 ), .A2(
        \SB2_1_29/i0[8] ), .A3(\SB2_1_29/i3[0] ), .ZN(
        \SB2_1_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_6/Component_Function_2/N2  ( .A1(\SB2_1_6/i0_3 ), .A2(
        \SB2_1_6/i0[10] ), .A3(\SB2_1_6/i0[6] ), .ZN(
        \SB2_1_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1644 ( .A1(\SB2_1_7/i0[6] ), .A2(\SB2_1_7/i0[9] ), .A3(
        \SB2_1_7/i1_5 ), .ZN(\SB2_1_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_18/Component_Function_3/N4  ( .A1(\SB2_1_18/i1_5 ), .A2(
        \SB2_1_18/i0[8] ), .A3(\SB2_1_18/i3[0] ), .ZN(
        \SB2_1_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_11/Component_Function_3/N4  ( .A1(\SB2_1_11/i1_5 ), .A2(
        \SB2_1_11/i0[8] ), .A3(\SB2_1_11/i3[0] ), .ZN(
        \SB2_1_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1753 ( .A1(\SB2_1_2/i0[8] ), .A2(\SB2_1_2/i3[0] ), .A3(
        \SB2_1_2/i1_5 ), .ZN(n2098) );
  NAND3_X1 U9484 ( .A1(\SB1_1_27/buf_output[3] ), .A2(\SB2_1_25/i1_7 ), .A3(
        \SB2_1_25/i1[9] ), .ZN(\SB2_1_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_23/Component_Function_3/N4  ( .A1(\SB2_1_23/i1_5 ), .A2(
        \SB2_1_23/i0[8] ), .A3(\SB2_1_23/i3[0] ), .ZN(
        \SB2_1_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_27/Component_Function_1/N2  ( .A1(\SB2_1_27/i0_3 ), .A2(
        \SB2_1_27/i1_7 ), .A3(\SB2_1_27/i0[8] ), .ZN(
        \SB2_1_27/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_6/Component_Function_3/N3  ( .A1(\SB2_1_6/i1[9] ), .A2(
        \SB2_1_6/i1_7 ), .A3(\SB2_1_6/i0[10] ), .ZN(
        \SB2_1_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_13/Component_Function_1/N3  ( .A1(\SB2_1_13/i1_5 ), .A2(
        \SB2_1_13/i0[6] ), .A3(\SB2_1_13/i0[9] ), .ZN(
        \SB2_1_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_17/Component_Function_3/N3  ( .A1(\SB2_1_17/i1[9] ), .A2(
        \SB2_1_17/i1_7 ), .A3(\SB2_1_17/i0[10] ), .ZN(
        \SB2_1_17/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_6/Component_Function_1/N4  ( .A1(\SB2_1_6/i1_7 ), .A2(
        \SB2_1_6/i0[8] ), .A3(\SB2_1_6/i0_4 ), .ZN(
        \SB2_1_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_8/Component_Function_1/N2  ( .A1(\SB2_1_8/i0_3 ), .A2(
        \SB2_1_8/i1_7 ), .A3(\SB2_1_8/i0[8] ), .ZN(
        \SB2_1_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_10/Component_Function_3/N4  ( .A1(\SB2_1_10/i1_5 ), .A2(
        \SB2_1_10/i0[8] ), .A3(\SB2_1_10/i3[0] ), .ZN(
        \SB2_1_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_19/Component_Function_1/N3  ( .A1(\SB2_1_19/i1_5 ), .A2(
        \SB2_1_19/i0[6] ), .A3(\SB2_1_19/i0[9] ), .ZN(
        \SB2_1_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U11772 ( .A1(\SB2_1_22/i0[9] ), .A2(\SB2_1_22/i0[6] ), .A3(
        \SB2_1_22/i1_5 ), .ZN(n4983) );
  NAND3_X1 \SB2_1_14/Component_Function_4/N2  ( .A1(\SB2_1_14/i3[0] ), .A2(
        \SB2_1_14/i0_0 ), .A3(\SB2_1_14/i1_7 ), .ZN(
        \SB2_1_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U5422 ( .A1(\SB2_1_26/i0_4 ), .A2(\SB2_1_26/i1_7 ), .A3(
        \SB2_1_26/i0[8] ), .ZN(n3378) );
  NAND3_X1 \SB2_1_14/Component_Function_0/N2  ( .A1(\SB2_1_14/i0[8] ), .A2(
        \SB2_1_14/i0[7] ), .A3(\SB2_1_14/i0[6] ), .ZN(
        \SB2_1_14/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_12/Component_Function_1/N4  ( .A1(\SB2_1_12/i1_7 ), .A2(
        \SB2_1_12/i0[8] ), .A3(\SB2_1_12/i0_4 ), .ZN(
        \SB2_1_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U6184 ( .A1(\SB2_1_4/i0[10] ), .A2(n2656), .A3(\SB2_1_4/i1[9] ), 
        .ZN(n2986) );
  NAND3_X1 U6694 ( .A1(\SB2_1_27/i0_3 ), .A2(\RI3[1][26] ), .A3(
        \SB2_1_27/i0[7] ), .ZN(n2909) );
  NAND3_X1 U8659 ( .A1(\SB2_1_21/i0[6] ), .A2(\SB2_1_21/i0[9] ), .A3(
        \SB2_1_21/i1_5 ), .ZN(\SB2_1_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1648 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB2_1_18/i0[9] ), .A3(
        \SB2_1_18/i0[8] ), .ZN(n5054) );
  NAND3_X1 \SB2_1_20/Component_Function_1/N2  ( .A1(\SB2_1_20/i0_3 ), .A2(
        \SB2_1_20/i1_7 ), .A3(\SB2_1_20/i0[8] ), .ZN(
        \SB2_1_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1074 ( .A1(\SB2_1_11/i0_0 ), .A2(\SB2_1_11/i1_5 ), .A3(
        \SB2_1_11/i0_4 ), .ZN(\SB2_1_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N4  ( .A1(\SB2_1_23/i1[9] ), .A2(
        \SB2_1_23/i1_5 ), .A3(\SB2_1_23/i0_4 ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U8284 ( .A1(\SB2_1_18/i0[10] ), .A2(\SB2_1_18/i0_3 ), .A3(
        \SB2_1_18/i0[6] ), .ZN(\SB2_1_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_28/Component_Function_0/N3  ( .A1(\SB2_1_28/i0[10] ), .A2(
        \SB2_1_28/i0_4 ), .A3(\SB2_1_28/i0_3 ), .ZN(
        \SB2_1_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1632 ( .A1(\SB2_1_8/i0_3 ), .A2(\SB2_1_8/i0[10] ), .A3(
        \SB2_1_8/i0_4 ), .ZN(\SB2_1_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3698 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0_4 ), .ZN(n1564) );
  NAND3_X1 \SB2_1_5/Component_Function_3/N4  ( .A1(\SB2_1_5/i1_5 ), .A2(
        \SB2_1_5/i0[8] ), .A3(\SB2_1_5/i3[0] ), .ZN(
        \SB2_1_5/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_21/Component_Function_0/N1  ( .A1(\SB2_1_21/i0[10] ), .A2(
        \SB2_1_21/i0[9] ), .ZN(\SB2_1_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U2749 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i0_0 ), .A3(
        \SB2_1_14/i0_4 ), .ZN(\SB2_1_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3695 ( .A1(\SB2_1_10/i1[9] ), .A2(\SB2_1_10/i1_5 ), .A3(
        \SB2_1_10/i0_4 ), .ZN(\SB2_1_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_0/Component_Function_1/N2  ( .A1(\SB2_1_0/i0_3 ), .A2(
        \SB2_1_0/i1_7 ), .A3(\SB2_1_0/i0[8] ), .ZN(
        \SB2_1_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_17/Component_Function_3/N1  ( .A1(\SB2_1_17/i1[9] ), .A2(
        \SB2_1_17/i0_3 ), .A3(\SB2_1_17/i0[6] ), .ZN(
        \SB2_1_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_3/N3  ( .A1(\SB2_1_5/i1[9] ), .A2(
        \SB2_1_5/i1_7 ), .A3(\SB2_1_5/i0[10] ), .ZN(
        \SB2_1_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_7/Component_Function_2/N1  ( .A1(\SB2_1_7/i1_5 ), .A2(
        \SB2_1_7/i0[10] ), .A3(\SB2_1_7/i1[9] ), .ZN(
        \SB2_1_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_14/Component_Function_2/N1  ( .A1(\SB2_1_14/i1_5 ), .A2(
        \SB2_1_14/i0[10] ), .A3(\SB2_1_14/i1[9] ), .ZN(
        \SB2_1_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_14/Component_Function_2/N3  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i0[8] ), .A3(\SB2_1_14/i0[9] ), .ZN(
        \SB2_1_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1063 ( .A1(\SB2_1_7/i0[9] ), .A2(\SB2_1_7/i0_3 ), .A3(
        \SB2_1_7/i0[8] ), .ZN(\SB2_1_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U8701 ( .A1(\RI3[1][26] ), .A2(\SB2_1_27/i1_5 ), .A3(
        \SB2_1_27/i0_4 ), .ZN(\SB2_1_27/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_27/Component_Function_2/N3  ( .A1(\SB2_1_27/i0_3 ), .A2(
        \SB2_1_27/i0[8] ), .A3(\SB2_1_27/i0[9] ), .ZN(
        \SB2_1_27/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_27/Component_Function_0/N1  ( .A1(\SB2_1_27/i0[10] ), .A2(
        \SB2_1_27/i0[9] ), .ZN(\SB2_1_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U9834 ( .A1(\SB2_1_21/i0_4 ), .A2(\SB2_1_21/i1_7 ), .A3(
        \SB2_1_21/i0[8] ), .ZN(\SB2_1_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4555 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0[10] ), .A3(
        \SB2_1_24/i0_4 ), .ZN(n1341) );
  NAND3_X1 U1046 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0_0 ), .A3(
        \SB2_1_9/i0[7] ), .ZN(n1714) );
  NAND3_X1 U12456 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i0[10] ), .A3(
        \SB2_1_5/i0_4 ), .ZN(n5286) );
  NAND3_X1 U9953 ( .A1(\SB2_1_7/i0[6] ), .A2(\SB2_1_7/i0_3 ), .A3(
        \SB2_1_7/i0[10] ), .ZN(n4065) );
  NAND3_X1 \SB2_1_27/Component_Function_1/N4  ( .A1(\SB2_1_27/i1_7 ), .A2(
        \SB2_1_27/i0[8] ), .A3(\SB2_1_27/i0_4 ), .ZN(
        \SB2_1_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_21/Component_Function_1/N2  ( .A1(\SB2_1_21/i0_3 ), .A2(
        \SB2_1_21/i1_7 ), .A3(\SB2_1_21/i0[8] ), .ZN(
        \SB2_1_21/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_10/Component_Function_4/N1  ( .A1(\SB2_1_10/i0[9] ), .A2(
        \SB2_1_10/i0_0 ), .A3(\SB2_1_10/i0[8] ), .ZN(
        \SB2_1_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2617 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i0[6] ), .A3(
        \SB2_1_14/i1[9] ), .ZN(\SB2_1_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1654 ( .A1(\SB2_1_27/i0[9] ), .A2(\SB2_1_27/i1_5 ), .A3(
        \SB2_1_27/i0[6] ), .ZN(n4673) );
  NAND3_X1 U1069 ( .A1(\SB2_1_21/i0[10] ), .A2(\SB2_1_21/i0_3 ), .A3(
        \SB2_1_21/i0_4 ), .ZN(\SB2_1_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_24/Component_Function_0/N4  ( .A1(\SB2_1_24/i0[7] ), .A2(
        \SB2_1_24/i0_3 ), .A3(\SB2_1_24/i0_0 ), .ZN(
        \SB2_1_24/Component_Function_0/NAND4_in[3] ) );
  INV_X1 U7 ( .I(n164), .ZN(n188) );
  INV_X1 U5 ( .I(n18), .ZN(n466) );
  NAND3_X1 U12552 ( .A1(\SB1_2_5/i0_4 ), .A2(\SB1_2_5/i1[9] ), .A3(
        \SB1_2_5/i1_5 ), .ZN(\SB1_2_5/Component_Function_4/NAND4_in[3] ) );
  INV_X4 \SB1_2_11/INV_5  ( .I(\SB1_2_11/i0_3 ), .ZN(\SB1_2_11/i1_5 ) );
  INV_X1 U1803 ( .I(\MC_ARK_ARC_1_1/buf_output[7] ), .ZN(\SB1_2_30/i1_7 ) );
  CLKBUF_X2 \SB1_2_8/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[138] ), .Z(
        \SB1_2_8/i0[9] ) );
  INV_X1 \SB1_2_27/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[24] ), .ZN(
        \SB1_2_27/i3[0] ) );
  INV_X1 \SB1_2_27/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[25] ), .ZN(
        \SB1_2_27/i1_7 ) );
  INV_X1 \SB1_2_26/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[30] ), .ZN(
        \SB1_2_26/i3[0] ) );
  INV_X1 \SB1_2_0/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[186] ), .ZN(
        \SB1_2_0/i3[0] ) );
  BUF_X2 \SB1_2_15/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[97] ), .Z(
        \SB1_2_15/i0[6] ) );
  INV_X1 \SB1_2_17/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[84] ), .ZN(
        \SB1_2_17/i3[0] ) );
  BUF_X2 \SB1_2_6/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[150] ), .Z(
        \SB1_2_6/i0[9] ) );
  INV_X1 U2213 ( .I(\MC_ARK_ARC_1_1/buf_output[73] ), .ZN(\SB1_2_19/i1_7 ) );
  BUF_X2 \SB1_2_31/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[0] ), .Z(
        \SB1_2_31/i0[9] ) );
  BUF_X2 \SB1_2_3/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[168] ), .Z(
        \SB1_2_3/i0[9] ) );
  BUF_X2 U7593 ( .I(\MC_ARK_ARC_1_1/buf_output[96] ), .Z(\SB1_2_15/i0[9] ) );
  BUF_X2 U5290 ( .I(\MC_ARK_ARC_1_1/buf_output[144] ), .Z(\SB1_2_7/i0[9] ) );
  CLKBUF_X2 U3703 ( .I(\MC_ARK_ARC_1_1/buf_output[90] ), .Z(\SB1_2_16/i0[9] )
         );
  CLKBUF_X2 \SB1_2_2/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[175] ), .Z(
        \SB1_2_2/i0[6] ) );
  BUF_X2 U2032 ( .I(\MC_ARK_ARC_1_1/buf_output[61] ), .Z(\SB1_2_21/i0[6] ) );
  BUF_X2 U1672 ( .I(\MC_ARK_ARC_1_1/buf_output[10] ), .Z(\SB1_2_30/i0_4 ) );
  BUF_X2 \SB1_2_10/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[127] ), .Z(
        \SB1_2_10/i0[6] ) );
  INV_X1 \SB1_2_1/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[180] ), .ZN(
        \SB1_2_1/i3[0] ) );
  INV_X2 \SB1_2_29/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[14] ), .ZN(
        \SB1_2_29/i1[9] ) );
  NAND3_X1 U7871 ( .A1(\SB1_2_6/i0[10] ), .A2(\SB1_2_6/i1[9] ), .A3(
        \SB1_2_6/i1_7 ), .ZN(n2616) );
  NAND3_X1 U12214 ( .A1(\SB1_2_16/i0[10] ), .A2(\SB1_2_16/i0_3 ), .A3(
        \SB1_2_16/i0[9] ), .ZN(n5142) );
  NAND3_X1 U5713 ( .A1(\SB1_2_16/i0_0 ), .A2(\SB1_2_16/i1_5 ), .A3(
        \SB1_2_16/i0_4 ), .ZN(\SB1_2_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_0/N3  ( .A1(\SB1_2_2/i0[10] ), .A2(
        \SB1_2_2/i0_4 ), .A3(\SB1_2_2/i0_3 ), .ZN(
        \SB1_2_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U5500 ( .A1(\SB1_2_13/i0[6] ), .A2(\SB1_2_13/i0[8] ), .A3(
        \SB1_2_13/i0[7] ), .ZN(\SB1_2_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 U11068 ( .A1(\SB1_2_24/i0[10] ), .A2(\SB1_2_24/i0[9] ), .ZN(n4544)
         );
  NAND3_X1 \SB1_2_28/Component_Function_4/N3  ( .A1(\SB1_2_28/i0[9] ), .A2(
        \SB1_2_28/i0[10] ), .A3(\SB1_2_28/i0_3 ), .ZN(
        \SB1_2_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_10/Component_Function_0/N3  ( .A1(\SB1_2_10/i0[10] ), .A2(
        \SB1_2_10/i0_4 ), .A3(\SB1_2_10/i0_3 ), .ZN(
        \SB1_2_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1002 ( .A1(\SB1_2_6/i3[0] ), .A2(\SB1_2_6/i1_5 ), .A3(
        \SB1_2_6/i0[8] ), .ZN(\SB1_2_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1550 ( .A1(\SB1_2_1/i0_0 ), .A2(\SB1_2_1/i1_7 ), .A3(
        \SB1_2_1/i3[0] ), .ZN(n4077) );
  NAND3_X1 \SB1_2_10/Component_Function_4/N2  ( .A1(\SB1_2_10/i3[0] ), .A2(
        \SB1_2_10/i0_0 ), .A3(\SB1_2_10/i1_7 ), .ZN(
        \SB1_2_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1613 ( .A1(\SB1_2_21/i0[8] ), .A2(\SB1_2_21/i3[0] ), .A3(
        \SB1_2_21/i1_5 ), .ZN(\SB1_2_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_10/Component_Function_0/N2  ( .A1(\SB1_2_10/i0[8] ), .A2(
        \SB1_2_10/i0[7] ), .A3(\SB1_2_10/i0[6] ), .ZN(
        \SB1_2_10/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_0/Component_Function_2/N1  ( .A1(\SB1_2_0/i1_5 ), .A2(
        \SB1_2_0/i0[10] ), .A3(\SB1_2_0/i1[9] ), .ZN(
        \SB1_2_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1614 ( .A1(\SB1_2_28/i3[0] ), .A2(\SB1_2_28/i0_0 ), .A3(
        \SB1_2_28/i1_7 ), .ZN(\SB1_2_28/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_29/Component_Function_5/N1  ( .A1(\SB1_2_29/i0_0 ), .A2(
        \SB1_2_29/i3[0] ), .ZN(\SB1_2_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U11295 ( .A1(\SB1_2_26/i0_0 ), .A2(\SB1_2_26/i3[0] ), .A3(
        \SB1_2_26/i1_7 ), .ZN(\SB1_2_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_0/Component_Function_2/N3  ( .A1(\RI1[2][191] ), .A2(
        \SB1_2_0/i0[8] ), .A3(\SB1_2_0/i0[9] ), .ZN(
        \SB1_2_0/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_7/Component_Function_5/N1  ( .A1(\SB1_2_7/i0_0 ), .A2(
        \SB1_2_7/i3[0] ), .ZN(\SB1_2_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3713 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i1_7 ), .A3(
        \SB1_2_13/i0[8] ), .ZN(\SB1_2_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_8/Component_Function_0/N4  ( .A1(\SB1_2_8/i0[7] ), .A2(
        \SB1_2_8/i0_3 ), .A3(\SB1_2_8/i0_0 ), .ZN(
        \SB1_2_8/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_13/Component_Function_5/N1  ( .A1(\SB1_2_13/i0_0 ), .A2(
        \SB1_2_13/i3[0] ), .ZN(\SB1_2_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_1/N3  ( .A1(\SB1_2_1/i1_5 ), .A2(
        \SB1_2_1/i0[6] ), .A3(\SB1_2_1/i0[9] ), .ZN(
        \SB1_2_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_18/Component_Function_2/N3  ( .A1(\SB1_2_18/i0_3 ), .A2(
        \SB1_2_18/i0[8] ), .A3(\SB1_2_18/i0[9] ), .ZN(
        \SB1_2_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_31/Component_Function_5/N4  ( .A1(\SB1_2_31/i0[9] ), .A2(
        \SB1_2_31/i0[6] ), .A3(\SB1_2_31/i0_4 ), .ZN(
        \SB1_2_31/Component_Function_5/NAND4_in[3] ) );
  INV_X1 \SB1_2_3/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[169] ), .ZN(
        \SB1_2_3/i1_7 ) );
  NAND3_X1 U3110 ( .A1(\SB1_2_14/i0[7] ), .A2(\RI1[2][107] ), .A3(
        \SB1_2_14/i0_0 ), .ZN(\SB1_2_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_17/Component_Function_1/N3  ( .A1(\SB1_2_17/i1_5 ), .A2(
        \SB1_2_17/i0[6] ), .A3(\SB1_2_17/i0[9] ), .ZN(
        \SB1_2_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4845 ( .A1(\SB1_2_9/i0[9] ), .A2(\SB1_2_9/i0_3 ), .A3(
        \SB1_2_9/i0[10] ), .ZN(n3305) );
  NAND3_X1 \SB1_2_17/Component_Function_2/N3  ( .A1(\SB1_2_17/i0_3 ), .A2(
        \SB1_2_17/i0[8] ), .A3(\SB1_2_17/i0[9] ), .ZN(
        \SB1_2_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3728 ( .A1(\SB1_2_20/i0[10] ), .A2(\SB1_2_20/i0[9] ), .A3(
        \SB1_2_20/i0_3 ), .ZN(\SB1_2_20/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U5986 ( .A1(\SB1_2_16/i0[10] ), .A2(\SB1_2_16/i0_3 ), .A3(
        \SB1_2_16/i0[6] ), .ZN(\SB1_2_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U974 ( .A1(\SB1_2_27/i0_0 ), .A2(\SB1_2_27/i0_3 ), .A3(
        \SB1_2_27/i0_4 ), .ZN(\SB1_2_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_14/Component_Function_4/N4  ( .A1(\SB1_2_14/i1[9] ), .A2(
        \SB1_2_14/i1_5 ), .A3(\SB1_2_14/i0_4 ), .ZN(
        \SB1_2_14/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U2503 ( .A1(\SB1_2_12/i1[9] ), .A2(\RI1[2][119] ), .ZN(n598) );
  NAND3_X1 U10213 ( .A1(\SB1_2_7/i1_5 ), .A2(\SB1_2_7/i0[10] ), .A3(
        \SB1_2_7/i1[9] ), .ZN(\SB1_2_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1624 ( .A1(\SB1_2_3/i0_4 ), .A2(\SB1_2_3/i0[10] ), .A3(
        \SB1_2_3/i0_3 ), .ZN(n3625) );
  NAND3_X1 U3725 ( .A1(\RI1[2][191] ), .A2(\SB1_2_0/i0_0 ), .A3(\SB1_2_0/i0_4 ), .ZN(\SB1_2_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1596 ( .A1(\SB1_2_9/i0[9] ), .A2(\SB1_2_9/i1_5 ), .A3(
        \SB1_2_9/i0[6] ), .ZN(n3832) );
  NAND2_X1 U3480 ( .A1(n2991), .A2(n840), .ZN(n4642) );
  NAND3_X1 \SB1_2_15/Component_Function_5/N4  ( .A1(\SB1_2_15/i0[9] ), .A2(
        \SB1_2_15/i0[6] ), .A3(\SB1_2_15/i0_4 ), .ZN(
        \SB1_2_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_26/Component_Function_2/N3  ( .A1(\SB1_2_26/i0_3 ), .A2(
        \SB1_2_26/i0[8] ), .A3(\SB1_2_26/i0[9] ), .ZN(
        \SB1_2_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_4/Component_Function_5/N3  ( .A1(\SB1_2_4/i1[9] ), .A2(
        \SB1_2_4/i0_4 ), .A3(\SB1_2_4/i0_3 ), .ZN(
        \SB1_2_4/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4769 ( .A1(\SB1_2_7/i0[9] ), .A2(\SB1_2_7/i0_4 ), .A3(
        \SB1_2_7/i0[6] ), .ZN(n3284) );
  NAND3_X1 U10392 ( .A1(\SB1_2_19/i0[6] ), .A2(\SB1_2_19/i0[9] ), .A3(
        \SB1_2_19/i0_4 ), .ZN(n4257) );
  NAND3_X1 U1589 ( .A1(\SB1_2_29/i0_4 ), .A2(\SB1_2_29/i1[9] ), .A3(
        \RI1[2][17] ), .ZN(n5035) );
  NAND3_X1 U8303 ( .A1(\SB1_2_5/i0[6] ), .A2(\SB1_2_5/i0_4 ), .A3(
        \SB1_2_5/i0[9] ), .ZN(n2857) );
  NAND3_X1 \SB1_2_14/Component_Function_0/N3  ( .A1(\SB1_2_14/i0[10] ), .A2(
        \SB1_2_14/i0_4 ), .A3(\RI1[2][107] ), .ZN(
        \SB1_2_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1527 ( .A1(\SB1_2_12/i1_5 ), .A2(\SB1_2_12/i0[10] ), .A3(
        \SB1_2_12/i1[9] ), .ZN(\SB1_2_12/Component_Function_2/NAND4_in[0] ) );
  AND2_X1 U5412 ( .A1(\MC_ARK_ARC_1_1/buf_output[16] ), .A2(
        \MC_ARK_ARC_1_1/buf_output[14] ), .Z(n2210) );
  NAND3_X1 \SB1_2_26/Component_Function_2/N2  ( .A1(\SB1_2_26/i0_3 ), .A2(
        \SB1_2_26/i0[10] ), .A3(\SB1_2_26/i0[6] ), .ZN(
        \SB1_2_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_16/Component_Function_2/N3  ( .A1(\SB1_2_16/i0_3 ), .A2(
        \SB1_2_16/i0[8] ), .A3(\SB1_2_16/i0[9] ), .ZN(
        \SB1_2_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1027 ( .A1(\SB1_2_2/i0_0 ), .A2(\SB1_2_2/i0[7] ), .A3(
        \SB1_2_2/i0_3 ), .ZN(n1777) );
  NAND3_X1 U11580 ( .A1(\SB1_2_28/i0_0 ), .A2(\SB1_2_28/i0[9] ), .A3(
        \SB1_2_28/i0[8] ), .ZN(\SB1_2_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U10556 ( .A1(\RI1[2][191] ), .A2(\SB1_2_0/i0[6] ), .A3(
        \SB1_2_0/i0[10] ), .ZN(\SB1_2_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_0/Component_Function_2/N4  ( .A1(\SB1_2_0/i1_5 ), .A2(
        \SB1_2_0/i0_0 ), .A3(\SB1_2_0/i0_4 ), .ZN(
        \SB1_2_0/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4561 ( .A1(\SB1_2_16/i0_3 ), .A2(\SB1_2_16/i0_4 ), .A3(
        \SB1_2_16/i1[9] ), .ZN(\SB1_2_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U6187 ( .A1(\SB1_2_8/i0[8] ), .A2(\SB1_2_8/i3[0] ), .A3(
        \SB1_2_8/i1_5 ), .ZN(\SB1_2_8/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 U3231 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i1[9] ), .ZN(
        \SB1_2_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1502 ( .A1(\SB1_2_29/i0[10] ), .A2(\RI1[2][17] ), .A3(
        \SB1_2_29/i0[6] ), .ZN(n3949) );
  NAND3_X1 U7988 ( .A1(\SB1_2_25/i0[10] ), .A2(\SB1_2_25/i0_3 ), .A3(
        \SB1_2_25/i0[6] ), .ZN(n3758) );
  NAND3_X1 U1580 ( .A1(\SB1_2_4/i0_0 ), .A2(\SB1_2_4/i0_3 ), .A3(
        \SB1_2_4/i0[7] ), .ZN(n3931) );
  NAND3_X1 U7572 ( .A1(\SB1_2_11/i1[9] ), .A2(\SB1_2_11/i0_4 ), .A3(
        \SB1_2_11/i0_3 ), .ZN(n2797) );
  NAND3_X1 U7938 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i0_0 ), .A3(
        \SB1_2_31/i0[7] ), .ZN(n2641) );
  NAND3_X1 \SB1_2_4/Component_Function_2/N2  ( .A1(\SB1_2_4/i0_3 ), .A2(
        \SB1_2_4/i0[10] ), .A3(\SB1_2_4/i0[6] ), .ZN(
        \SB1_2_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_13/Component_Function_3/N4  ( .A1(\SB1_2_13/i1_5 ), .A2(
        \SB1_2_13/i0[8] ), .A3(\SB1_2_13/i3[0] ), .ZN(
        \SB1_2_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_17/Component_Function_4/N3  ( .A1(\SB1_2_17/i0[9] ), .A2(
        \SB1_2_17/i0[10] ), .A3(\SB1_2_17/i0_3 ), .ZN(
        \SB1_2_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U8137 ( .A1(\SB1_2_17/i0_0 ), .A2(\SB1_2_17/i1_7 ), .A3(
        \SB1_2_17/i3[0] ), .ZN(\SB1_2_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U6489 ( .A1(\SB1_2_30/i0[8] ), .A2(\SB1_2_30/i1_5 ), .A3(
        \SB1_2_30/i3[0] ), .ZN(\SB1_2_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1510 ( .A1(\SB1_2_11/i0[8] ), .A2(\SB1_2_11/i1_7 ), .A3(
        \SB1_2_11/i0_4 ), .ZN(n3276) );
  NAND3_X1 U9825 ( .A1(\SB1_2_29/i0_0 ), .A2(\RI1[2][17] ), .A3(
        \SB1_2_29/i0[7] ), .ZN(n1805) );
  NAND3_X1 U7232 ( .A1(\SB1_2_11/i0_0 ), .A2(\SB1_2_11/i0[7] ), .A3(
        \SB1_2_11/i0_3 ), .ZN(n2297) );
  NAND2_X1 \SB1_2_0/Component_Function_1/N1  ( .A1(\RI1[2][191] ), .A2(
        \SB1_2_0/i1[9] ), .ZN(\SB1_2_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_2/N1  ( .A1(\SB1_2_23/i1_5 ), .A2(
        \SB1_2_23/i0[10] ), .A3(\SB1_2_23/i1[9] ), .ZN(
        \SB1_2_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U992 ( .A1(\SB1_2_2/i0[10] ), .A2(\SB1_2_2/i1[9] ), .A3(
        \SB1_2_2/i1_7 ), .ZN(\SB1_2_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U6995 ( .A1(\SB1_2_3/i0[9] ), .A2(\SB1_2_3/i0_3 ), .A3(
        \SB1_2_3/i0[8] ), .ZN(n1234) );
  NAND3_X1 U3718 ( .A1(\SB1_2_24/i0[10] ), .A2(\SB1_2_24/i1[9] ), .A3(
        \SB1_2_24/i1_7 ), .ZN(n1019) );
  NAND3_X1 U1001 ( .A1(\SB1_2_28/i0[8] ), .A2(\SB1_2_28/i0_4 ), .A3(
        \SB1_2_28/i1_7 ), .ZN(n2135) );
  NAND3_X1 \SB1_2_21/Component_Function_1/N3  ( .A1(\SB1_2_21/i1_5 ), .A2(
        \SB1_2_21/i0[6] ), .A3(\SB1_2_21/i0[9] ), .ZN(
        \SB1_2_21/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U1563 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i3[0] ), .ZN(
        \SB1_2_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_1/N3  ( .A1(\SB1_2_30/i1_5 ), .A2(
        \SB1_2_30/i0[6] ), .A3(\SB1_2_30/i0[9] ), .ZN(
        \SB1_2_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_2/Component_Function_2/N3  ( .A1(\SB1_2_2/i0_3 ), .A2(
        \SB1_2_2/i0[8] ), .A3(\SB1_2_2/i0[9] ), .ZN(
        \SB1_2_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U7804 ( .A1(\SB1_2_11/i0[10] ), .A2(\SB1_2_11/i0_0 ), .A3(
        \SB1_2_11/i0[6] ), .ZN(\SB1_2_11/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_29/Component_Function_2/N3  ( .A1(\RI1[2][17] ), .A2(
        \SB1_2_29/i0[8] ), .A3(\SB1_2_29/i0[9] ), .ZN(
        \SB1_2_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1576 ( .A1(\SB1_2_9/i0[9] ), .A2(\SB1_2_9/i0_3 ), .A3(
        \SB1_2_9/i0[8] ), .ZN(n4411) );
  NAND3_X1 \SB1_2_21/Component_Function_4/N1  ( .A1(\SB1_2_21/i0[9] ), .A2(
        \SB1_2_21/i0_0 ), .A3(\SB1_2_21/i0[8] ), .ZN(
        \SB1_2_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_4/N3  ( .A1(\SB1_2_8/i0[9] ), .A2(
        \SB1_2_8/i0[10] ), .A3(\SB1_2_8/i0_3 ), .ZN(
        \SB1_2_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_30/Component_Function_3/N1  ( .A1(\SB1_2_30/i1[9] ), .A2(
        \SB1_2_30/i0_3 ), .A3(\SB1_2_30/i0[6] ), .ZN(
        \SB1_2_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U7455 ( .A1(\SB1_2_23/i0_0 ), .A2(\SB1_2_23/i1_5 ), .A3(
        \SB1_2_23/i0_4 ), .ZN(n2403) );
  NAND3_X1 \SB1_2_13/Component_Function_2/N3  ( .A1(\SB1_2_13/i0_3 ), .A2(
        \SB1_2_13/i0[8] ), .A3(\SB1_2_13/i0[9] ), .ZN(
        \SB1_2_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4338 ( .A1(\SB1_2_1/i0[6] ), .A2(\SB1_2_1/i0[9] ), .A3(
        \SB1_2_1/i0_4 ), .ZN(n3209) );
  NAND3_X1 U1500 ( .A1(\SB1_2_22/i1_5 ), .A2(\SB1_2_22/i0[9] ), .A3(
        \SB1_2_22/i0[6] ), .ZN(n3863) );
  NAND2_X1 \SB1_2_28/Component_Function_5/N1  ( .A1(\SB1_2_28/i0_0 ), .A2(
        \SB1_2_28/i3[0] ), .ZN(\SB1_2_28/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_28/Component_Function_1/N1  ( .A1(\SB1_2_28/i0_3 ), .A2(
        \SB1_2_28/i1[9] ), .ZN(\SB1_2_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U6944 ( .A1(\RI1[2][101] ), .A2(\SB1_2_15/i0[7] ), .A3(
        \SB1_2_15/i0_0 ), .ZN(n2167) );
  NAND3_X1 \SB1_2_12/Component_Function_5/N4  ( .A1(\SB1_2_12/i0[9] ), .A2(
        \SB1_2_12/i0[6] ), .A3(\SB1_2_12/i0_4 ), .ZN(
        \SB1_2_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_13/Component_Function_4/N3  ( .A1(\SB1_2_13/i0[9] ), .A2(
        \SB1_2_13/i0[10] ), .A3(\SB1_2_13/i0_3 ), .ZN(
        \SB1_2_13/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U1540 ( .A1(\SB1_2_3/i0_3 ), .A2(\SB1_2_3/i1[9] ), .ZN(
        \SB1_2_3/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_0/Component_Function_5/N1  ( .A1(\SB1_2_0/i0_0 ), .A2(
        \SB1_2_0/i3[0] ), .ZN(\SB1_2_0/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_21/Component_Function_0/N1  ( .A1(\SB1_2_21/i0[10] ), .A2(
        \SB1_2_21/i0[9] ), .ZN(\SB1_2_21/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U1554 ( .A1(\SB1_2_22/i0[9] ), .A2(\SB1_2_22/i0[10] ), .ZN(n4176)
         );
  NAND3_X1 U2234 ( .A1(\SB1_2_0/i1_7 ), .A2(\SB1_2_0/i0[8] ), .A3(
        \SB1_2_0/i0_4 ), .ZN(\SB1_2_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U981 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i1[9] ), .A3(
        \SB1_2_21/i0_4 ), .ZN(n2981) );
  NAND3_X1 \SB1_2_19/Component_Function_3/N1  ( .A1(\SB1_2_19/i1[9] ), .A2(
        \SB1_2_19/i0_3 ), .A3(\SB1_2_19/i0[6] ), .ZN(
        \SB1_2_19/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U2027 ( .A1(\SB1_2_22/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_22/Component_Function_4/NAND4_in[0] ), .ZN(n2605) );
  NAND3_X1 \SB1_2_2/Component_Function_5/N2  ( .A1(\SB1_2_2/i0_0 ), .A2(
        \SB1_2_2/i0[6] ), .A3(\SB1_2_2/i0[10] ), .ZN(
        \SB1_2_2/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U988 ( .A1(\SB1_2_14/i0[10] ), .A2(\RI1[2][107] ), .A3(
        \SB1_2_14/i0[6] ), .ZN(n1855) );
  NAND3_X1 \SB1_2_19/Component_Function_3/N2  ( .A1(\SB1_2_19/i0_0 ), .A2(
        \SB1_2_19/i0_3 ), .A3(\SB1_2_19/i0_4 ), .ZN(
        \SB1_2_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_13/Component_Function_2/N2  ( .A1(\SB1_2_13/i0_3 ), .A2(
        \SB1_2_13/i0[10] ), .A3(\SB1_2_13/i0[6] ), .ZN(
        \SB1_2_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1013 ( .A1(\SB1_2_26/i0[6] ), .A2(\SB1_2_26/i0_4 ), .A3(
        \SB1_2_26/i0[9] ), .ZN(n1710) );
  NAND3_X1 \SB1_2_0/Component_Function_1/N3  ( .A1(\SB1_2_0/i1_5 ), .A2(
        \SB1_2_0/i0[6] ), .A3(\SB1_2_0/i0[9] ), .ZN(
        \SB1_2_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U8024 ( .A1(\SB1_2_5/i0_0 ), .A2(\SB1_2_5/i1_5 ), .A3(
        \SB1_2_5/i0_4 ), .ZN(n2685) );
  NAND3_X1 U1524 ( .A1(\SB1_2_24/i0[6] ), .A2(\SB1_2_24/i0[10] ), .A3(
        \SB1_2_24/i0_3 ), .ZN(n4951) );
  NAND3_X1 \SB1_2_26/Component_Function_3/N1  ( .A1(\SB1_2_26/i1[9] ), .A2(
        \SB1_2_26/i0_3 ), .A3(\SB1_2_26/i0[6] ), .ZN(
        \SB1_2_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_26/Component_Function_3/N2  ( .A1(\SB1_2_26/i0_0 ), .A2(
        \SB1_2_26/i0_3 ), .A3(\SB1_2_26/i0_4 ), .ZN(
        \SB1_2_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U6735 ( .A1(\SB1_2_29/i0_4 ), .A2(\RI1[2][17] ), .A3(
        \SB1_2_29/i0[10] ), .ZN(\SB1_2_29/Component_Function_0/NAND4_in[2] )
         );
  NAND2_X1 \SB1_2_4/Component_Function_0/N1  ( .A1(\SB1_2_4/i0[10] ), .A2(
        \SB1_2_4/i0[9] ), .ZN(\SB1_2_4/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_29/Component_Function_0/N1  ( .A1(\SB1_2_29/i0[10] ), .A2(
        \SB1_2_29/i0[9] ), .ZN(\SB1_2_29/Component_Function_0/NAND4_in[0] ) );
  NAND4_X1 U4190 ( .A1(\SB1_2_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_5/Component_Function_2/NAND4_in[1] ), .A3(n2685), .A4(
        \SB1_2_5/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_2_5/buf_output[2] ) );
  BUF_X2 \SB2_2_8/BUF_0  ( .I(\SB1_2_13/buf_output[0] ), .Z(\SB2_2_8/i0[9] )
         );
  BUF_X2 \SB2_2_4/BUF_0  ( .I(\SB1_2_9/buf_output[0] ), .Z(\SB2_2_4/i0[9] ) );
  BUF_X2 \SB2_2_23/BUF_0  ( .I(\SB1_2_28/buf_output[0] ), .Z(\SB2_2_23/i0[9] )
         );
  NAND3_X1 U9702 ( .A1(\SB2_2_19/i0_4 ), .A2(\SB2_2_19/i0_3 ), .A3(
        \SB2_2_19/i1[9] ), .ZN(n4298) );
  NAND3_X1 U3190 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0_4 ), .A3(
        \SB2_2_25/i1[9] ), .ZN(\SB2_2_25/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_15/Component_Function_5/N1  ( .A1(\SB2_2_15/i0_0 ), .A2(
        \SB2_2_15/i3[0] ), .ZN(\SB2_2_15/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_14/Component_Function_5/N1  ( .A1(\SB2_2_14/i0_0 ), .A2(
        \SB2_2_14/i3[0] ), .ZN(\SB2_2_14/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_23/Component_Function_5/N1  ( .A1(\SB2_2_23/i0_0 ), .A2(
        \SB2_2_23/i3[0] ), .ZN(\SB2_2_23/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U5492 ( .A1(\SB2_2_4/i0_0 ), .A2(\SB2_2_4/i3[0] ), .ZN(n1520) );
  NAND2_X1 \SB2_2_8/Component_Function_5/N1  ( .A1(\SB2_2_8/i0_0 ), .A2(
        \SB2_2_8/i3[0] ), .ZN(\SB2_2_8/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_30/Component_Function_5/N1  ( .A1(\SB2_2_30/i0_0 ), .A2(
        \SB2_2_30/i3[0] ), .ZN(\SB2_2_30/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U9802 ( .I(\SB1_2_22/buf_output[0] ), .ZN(\SB2_2_17/i3[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_5/N2  ( .A1(\SB2_2_29/i0_0 ), .A2(
        \SB2_2_29/i0[6] ), .A3(\SB2_2_29/i0[10] ), .ZN(
        \SB2_2_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U5990 ( .A1(\SB2_2_3/i0[10] ), .A2(\SB2_2_3/i0_0 ), .A3(
        \SB2_2_3/i0[6] ), .ZN(\SB2_2_3/Component_Function_5/NAND4_in[1] ) );
  BUF_X2 U2026 ( .I(\SB1_2_16/buf_output[0] ), .Z(\SB2_2_11/i0[9] ) );
  INV_X1 \SB2_2_10/INV_1  ( .I(\SB1_2_14/buf_output[1] ), .ZN(\SB2_2_10/i1_7 )
         );
  CLKBUF_X2 \SB2_2_6/BUF_1  ( .I(\SB1_2_10/buf_output[1] ), .Z(\SB2_2_6/i0[6] ) );
  CLKBUF_X2 \SB2_2_6/BUF_0  ( .I(\SB1_2_11/buf_output[0] ), .Z(\SB2_2_6/i0[9] ) );
  BUF_X2 \SB2_2_18/BUF_0  ( .I(\SB1_2_23/buf_output[0] ), .Z(\SB2_2_18/i0[9] )
         );
  BUF_X2 \SB2_2_2/BUF_2  ( .I(\SB1_2_5/buf_output[2] ), .Z(\SB2_2_2/i0_0 ) );
  CLKBUF_X2 \SB2_2_1/BUF_1  ( .I(\SB1_2_5/buf_output[1] ), .Z(\SB2_2_1/i0[6] )
         );
  INV_X1 \SB2_2_2/INV_0  ( .I(\SB1_2_7/buf_output[0] ), .ZN(\SB2_2_2/i3[0] )
         );
  INV_X1 \SB2_2_22/INV_0  ( .I(\SB1_2_27/buf_output[0] ), .ZN(\SB2_2_22/i3[0] ) );
  INV_X1 \SB2_2_13/INV_1  ( .I(\SB1_2_17/buf_output[1] ), .ZN(\SB2_2_13/i1_7 )
         );
  INV_X1 \SB2_2_7/INV_1  ( .I(\SB1_2_11/buf_output[1] ), .ZN(\SB2_2_7/i1_7 )
         );
  INV_X1 \SB2_2_31/INV_3  ( .I(\SB1_2_1/buf_output[3] ), .ZN(\SB2_2_31/i0[8] )
         );
  INV_X1 \SB2_2_12/INV_1  ( .I(\SB1_2_16/buf_output[1] ), .ZN(\SB2_2_12/i1_7 )
         );
  NAND2_X1 \SB2_2_27/Component_Function_1/N1  ( .A1(\SB2_2_27/i0_3 ), .A2(
        \SB2_2_27/i1[9] ), .ZN(\SB2_2_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U5514 ( .A1(\SB2_2_15/i0[10] ), .A2(\SB2_2_15/i0_3 ), .A3(
        \SB2_2_15/i0[9] ), .ZN(n1529) );
  NAND3_X1 \SB2_2_24/Component_Function_3/N4  ( .A1(\SB2_2_24/i1_5 ), .A2(
        \SB2_2_24/i0[8] ), .A3(\SB2_2_24/i3[0] ), .ZN(
        \SB2_2_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U7881 ( .A1(\SB2_2_10/i0_4 ), .A2(\SB2_2_10/i1[9] ), .A3(n589), 
        .ZN(n2620) );
  NAND3_X1 \SB2_2_18/Component_Function_3/N4  ( .A1(\SB2_2_18/i1_5 ), .A2(
        \SB2_2_18/i0[8] ), .A3(\SB2_2_18/i3[0] ), .ZN(
        \SB2_2_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2803 ( .A1(\SB2_2_9/i0_4 ), .A2(\SB2_2_9/i0[8] ), .A3(
        \SB2_2_9/i1_7 ), .ZN(n5390) );
  NAND2_X1 \SB2_2_31/Component_Function_5/N1  ( .A1(\SB2_2_31/i0_0 ), .A2(
        \SB2_2_31/i3[0] ), .ZN(\SB2_2_31/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_2/Component_Function_5/N1  ( .A1(\SB2_2_2/i0_0 ), .A2(
        \SB2_2_2/i3[0] ), .ZN(\SB2_2_2/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_18/Component_Function_5/N1  ( .A1(\SB2_2_18/i0_0 ), .A2(
        \SB2_2_18/i3[0] ), .ZN(\SB2_2_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_12/Component_Function_4/N2  ( .A1(\SB2_2_12/i3[0] ), .A2(
        \SB2_2_12/i0_0 ), .A3(\SB2_2_12/i1_7 ), .ZN(
        \SB2_2_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U6291 ( .A1(\SB2_2_4/i0[7] ), .A2(\SB2_2_4/i0[6] ), .A3(
        \SB2_2_4/i0[8] ), .ZN(\SB2_2_4/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_20/Component_Function_1/N3  ( .A1(\SB2_2_20/i1_5 ), .A2(
        \SB2_2_20/i0[6] ), .A3(\SB2_2_20/i0[9] ), .ZN(
        \SB2_2_20/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_16/Component_Function_5/N1  ( .A1(\SB2_2_16/i0_0 ), .A2(
        \SB2_2_16/i3[0] ), .ZN(\SB2_2_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U9700 ( .A1(\SB2_2_19/i0[10] ), .A2(\SB2_2_19/i1_5 ), .A3(
        \SB2_2_19/i1[9] ), .ZN(\SB2_2_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U9696 ( .A1(\SB2_2_21/i1[9] ), .A2(\SB2_2_21/i1_5 ), .A3(
        \SB1_2_22/buf_output[4] ), .ZN(
        \SB2_2_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_24/Component_Function_4/N4  ( .A1(\SB2_2_24/i1[9] ), .A2(
        \SB2_2_24/i1_5 ), .A3(\SB2_2_24/i0_4 ), .ZN(
        \SB2_2_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_30/Component_Function_4/N4  ( .A1(\SB2_2_30/i1[9] ), .A2(
        \SB2_2_30/i1_5 ), .A3(\SB2_2_30/i0_4 ), .ZN(
        \SB2_2_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U5796 ( .A1(\SB2_2_1/i0_0 ), .A2(\SB2_2_1/i1_5 ), .A3(
        \SB1_2_2/buf_output[4] ), .ZN(n1655) );
  NAND3_X1 U9813 ( .A1(\SB2_2_22/i0_0 ), .A2(\SB2_2_22/i0[8] ), .A3(
        \SB2_2_22/i0[9] ), .ZN(\SB2_2_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1431 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0[10] ), .A3(
        \SB2_2_4/i0_4 ), .ZN(\SB2_2_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11155 ( .A1(\SB2_2_11/i0_3 ), .A2(\SB2_2_11/i1[9] ), .A3(
        \SB2_2_11/i0_4 ), .ZN(n1766) );
  NAND3_X1 U8687 ( .A1(\SB2_2_25/i0[10] ), .A2(\SB2_2_25/i1[9] ), .A3(
        \SB2_2_25/i1_7 ), .ZN(n3082) );
  NAND3_X1 U913 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0[10] ), .A3(
        \SB2_2_16/i0_4 ), .ZN(n1067) );
  NAND3_X1 \SB2_2_23/Component_Function_4/N3  ( .A1(\SB2_2_23/i0[9] ), .A2(
        \SB2_2_23/i0[10] ), .A3(\SB2_2_23/i0_3 ), .ZN(
        \SB2_2_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U11038 ( .A1(\SB2_2_7/i0_3 ), .A2(\SB2_2_7/i0[9] ), .A3(
        \SB2_2_7/i0[8] ), .ZN(n4536) );
  INV_X1 U3115 ( .I(\SB2_2_26/i0_4 ), .ZN(\SB2_2_26/i0[7] ) );
  NAND2_X1 \SB2_2_16/Component_Function_0/N1  ( .A1(\SB2_2_16/i0[10] ), .A2(
        \SB2_2_16/i0[9] ), .ZN(\SB2_2_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_0/Component_Function_4/N1  ( .A1(\SB2_2_0/i0[9] ), .A2(
        \SB2_2_0/i0_0 ), .A3(\SB2_2_0/i0[8] ), .ZN(
        \SB2_2_0/Component_Function_4/NAND4_in[0] ) );
  BUF_X2 U8983 ( .I(\SB1_2_18/buf_output[4] ), .Z(\RI3[2][88] ) );
  INV_X1 \SB2_2_14/INV_1  ( .I(\SB1_2_18/buf_output[1] ), .ZN(\SB2_2_14/i1_7 )
         );
  NAND3_X1 \SB2_2_12/Component_Function_4/N1  ( .A1(\SB2_2_12/i0[9] ), .A2(
        \SB2_2_12/i0_0 ), .A3(\SB2_2_12/i0[8] ), .ZN(
        \SB2_2_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U3770 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i1_7 ), .A3(
        \SB2_2_24/i0[8] ), .ZN(\SB2_2_24/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3759 ( .A1(\SB2_2_30/i1[9] ), .A2(\SB2_2_30/i0_3 ), .A3(
        \SB2_2_30/i0[6] ), .ZN(\SB2_2_30/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_12/Component_Function_1/N1  ( .A1(\SB2_2_12/i0_3 ), .A2(
        \SB2_2_12/i1[9] ), .ZN(\SB2_2_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_4/N3  ( .A1(\SB2_2_19/i0[9] ), .A2(
        \SB2_2_19/i0[10] ), .A3(\SB2_2_19/i0_3 ), .ZN(
        \SB2_2_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3578 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0_0 ), .A3(
        \SB2_2_14/i0[7] ), .ZN(\SB2_2_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1427 ( .A1(\SB2_2_2/i0_4 ), .A2(\SB2_2_2/i0_3 ), .A3(
        \SB2_2_2/i0[10] ), .ZN(n4387) );
  NAND3_X1 \SB2_2_4/Component_Function_2/N3  ( .A1(\SB2_2_4/i0_3 ), .A2(
        \SB2_2_4/i0[8] ), .A3(\SB2_2_4/i0[9] ), .ZN(
        \SB2_2_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_25/Component_Function_4/N2  ( .A1(\SB2_2_25/i3[0] ), .A2(
        \SB2_2_25/i0_0 ), .A3(\SB2_2_25/i1_7 ), .ZN(
        \SB2_2_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U957 ( .A1(\SB2_2_20/i0[10] ), .A2(\SB2_2_20/i0_3 ), .A3(
        \SB2_2_20/i0_4 ), .ZN(n2165) );
  NAND2_X1 \SB2_2_16/Component_Function_1/N1  ( .A1(\SB2_2_16/i0_3 ), .A2(
        \SB2_2_16/i1[9] ), .ZN(\SB2_2_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10422 ( .A1(\SB2_2_6/i0_3 ), .A2(\SB2_2_6/i0_0 ), .A3(
        \SB2_2_6/i0_4 ), .ZN(\SB2_2_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1483 ( .A1(\SB2_2_31/i1_5 ), .A2(\SB2_2_31/i0_4 ), .A3(
        \SB2_2_31/i1[9] ), .ZN(n4434) );
  NAND3_X1 U2257 ( .A1(\SB2_2_27/i0[9] ), .A2(\SB2_2_27/i0[10] ), .A3(
        \SB2_2_27/i0_3 ), .ZN(\SB2_2_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U5826 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0[10] ), .A3(
        \SB2_2_25/i0[9] ), .ZN(\SB2_2_25/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_28/Component_Function_5/N1  ( .A1(\SB2_2_28/i0_0 ), .A2(
        \SB2_2_28/i3[0] ), .ZN(\SB2_2_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_11/Component_Function_2/N3  ( .A1(\SB2_2_11/i0_3 ), .A2(
        \SB2_2_11/i0[8] ), .A3(\SB2_2_11/i0[9] ), .ZN(
        \SB2_2_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_29/Component_Function_0/N2  ( .A1(\SB2_2_29/i0[8] ), .A2(
        \SB2_2_29/i0[7] ), .A3(\SB2_2_29/i0[6] ), .ZN(
        \SB2_2_29/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_17/Component_Function_0/N2  ( .A1(\SB2_2_17/i0[8] ), .A2(
        \SB2_2_17/i0[7] ), .A3(\SB2_2_17/i0[6] ), .ZN(
        \SB2_2_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_20/Component_Function_0/N2  ( .A1(\SB2_2_20/i0[8] ), .A2(
        \SB2_2_20/i0[7] ), .A3(\SB2_2_20/i0[6] ), .ZN(
        \SB2_2_20/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3762 ( .A1(\SB2_2_13/i0[9] ), .A2(\SB2_2_13/i0_0 ), .A3(
        \SB2_2_13/i0[8] ), .ZN(\SB2_2_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1738 ( .A1(\SB2_2_9/i1_5 ), .A2(\SB2_2_9/i0[8] ), .A3(
        \SB2_2_9/i3[0] ), .ZN(\SB2_2_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_28/Component_Function_2/N1  ( .A1(\SB2_2_28/i1_5 ), .A2(
        \SB2_2_28/i0[10] ), .A3(\SB2_2_28/i1[9] ), .ZN(
        \SB2_2_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_5/Component_Function_1/N4  ( .A1(\SB2_2_5/i1_7 ), .A2(
        \SB2_2_5/i0[8] ), .A3(\SB2_2_5/i0_4 ), .ZN(
        \SB2_2_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_1/Component_Function_1/N2  ( .A1(\SB2_2_1/i0_3 ), .A2(
        \SB2_2_1/i1_7 ), .A3(\SB2_2_1/i0[8] ), .ZN(
        \SB2_2_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_21/Component_Function_3/N4  ( .A1(\SB2_2_21/i1_5 ), .A2(
        \SB2_2_21/i0[8] ), .A3(\SB2_2_21/i3[0] ), .ZN(
        \SB2_2_21/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_21/Component_Function_5/N1  ( .A1(\SB2_2_21/i0_0 ), .A2(
        \SB2_2_21/i3[0] ), .ZN(\SB2_2_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_4/N4  ( .A1(\SB2_2_25/i1[9] ), .A2(
        \SB2_2_25/i1_5 ), .A3(\SB2_2_25/i0_4 ), .ZN(
        \SB2_2_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_3/Component_Function_0/N2  ( .A1(n3991), .A2(\SB2_2_3/i0[7] ), .A3(\SB2_2_3/i0[6] ), .ZN(\SB2_2_3/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U10258 ( .A1(\SB2_2_15/i0_0 ), .A2(\SB2_2_15/i1_5 ), .A3(
        \SB2_2_15/i0_4 ), .ZN(\SB2_2_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U10219 ( .A1(\SB2_2_7/i0_0 ), .A2(\SB2_2_7/i0[9] ), .A3(
        \SB2_2_7/i0[8] ), .ZN(\SB2_2_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2866 ( .A1(\SB2_2_22/i1_5 ), .A2(\SB2_2_22/i0[8] ), .A3(
        \SB2_2_22/i3[0] ), .ZN(\SB2_2_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_0/Component_Function_1/N3  ( .A1(\SB2_2_0/i1_5 ), .A2(
        \SB2_2_0/i0[6] ), .A3(\SB2_2_0/i0[9] ), .ZN(
        \SB2_2_0/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_20/Component_Function_5/N1  ( .A1(\SB2_2_20/i0_0 ), .A2(
        \SB2_2_20/i3[0] ), .ZN(\SB2_2_20/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U2267 ( .A1(\SB2_2_1/i0_0 ), .A2(\SB2_2_1/i3[0] ), .ZN(
        \SB2_2_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2537 ( .A1(\SB2_2_18/i0[6] ), .A2(\SB2_2_18/i1_5 ), .A3(
        \SB2_2_18/i0[9] ), .ZN(\SB2_2_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_10/Component_Function_1/N2  ( .A1(\SB2_2_10/i0_3 ), .A2(
        \SB2_2_10/i1_7 ), .A3(\SB2_2_10/i0[8] ), .ZN(
        \SB2_2_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U10367 ( .A1(\SB2_2_10/i0_0 ), .A2(\SB2_2_10/i3[0] ), .ZN(n4245) );
  NAND3_X1 U8589 ( .A1(\SB2_2_21/i0[10] ), .A2(\SB2_2_21/i1_5 ), .A3(
        \SB2_2_21/i1[9] ), .ZN(\SB2_2_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_1/N3  ( .A1(\SB2_2_25/i1_5 ), .A2(
        \SB2_2_25/i0[6] ), .A3(\SB2_2_25/i0[9] ), .ZN(
        \SB2_2_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U12652 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i1[9] ), .A3(
        \SB2_2_0/i0[6] ), .ZN(\SB2_2_0/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U4489 ( .A1(\SB2_2_31/i0[9] ), .A2(\SB2_2_31/i0[10] ), .ZN(n3234)
         );
  NAND3_X1 \SB2_2_7/Component_Function_0/N2  ( .A1(\SB2_2_7/i0[8] ), .A2(
        \SB2_2_7/i0[7] ), .A3(\SB2_2_7/i0[6] ), .ZN(
        \SB2_2_7/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2259 ( .A1(\SB2_2_9/i1[9] ), .A2(\SB2_2_9/i1_5 ), .A3(
        \SB2_2_9/i0_4 ), .ZN(\SB2_2_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3747 ( .A1(\SB2_2_2/i0_4 ), .A2(\SB2_2_2/i1_7 ), .A3(
        \SB2_2_2/i0[8] ), .ZN(n3738) );
  NAND3_X1 \SB2_2_24/Component_Function_2/N4  ( .A1(\SB2_2_24/i1_5 ), .A2(
        \SB2_2_24/i0_0 ), .A3(\SB2_2_24/i0_4 ), .ZN(
        \SB2_2_24/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U6078 ( .A1(\SB2_2_31/i0_3 ), .A2(\SB2_2_31/i0[10] ), .A3(
        \SB2_2_31/i0_4 ), .ZN(n1770) );
  NAND3_X1 \SB2_2_8/Component_Function_1/N3  ( .A1(\SB2_2_8/i1_5 ), .A2(
        \SB2_2_8/i0[6] ), .A3(\SB2_2_8/i0[9] ), .ZN(
        \SB2_2_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_13/Component_Function_1/N3  ( .A1(\SB2_2_13/i1_5 ), .A2(
        \SB2_2_13/i0[6] ), .A3(\SB2_2_13/i0[9] ), .ZN(
        \SB2_2_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_0/Component_Function_3/N3  ( .A1(\SB2_2_0/i1[9] ), .A2(
        \SB2_2_0/i1_7 ), .A3(\SB2_2_0/i0[10] ), .ZN(
        \SB2_2_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U966 ( .A1(\SB2_2_10/i0_3 ), .A2(\SB2_2_10/i1[9] ), .A3(
        \SB2_2_10/i0_4 ), .ZN(\SB2_2_10/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_14/Component_Function_3/N4  ( .A1(\SB2_2_14/i1_5 ), .A2(
        \SB2_2_14/i0[8] ), .A3(\SB2_2_14/i3[0] ), .ZN(
        \SB2_2_14/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_14/Component_Function_0/N1  ( .A1(\SB2_2_14/i0[10] ), .A2(
        \SB2_2_14/i0[9] ), .ZN(\SB2_2_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_20/Component_Function_4/N4  ( .A1(\SB2_2_20/i1[9] ), .A2(
        \SB2_2_20/i1_5 ), .A3(\SB2_2_20/i0_4 ), .ZN(
        \SB2_2_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_27/Component_Function_4/N4  ( .A1(\SB2_2_27/i1[9] ), .A2(
        \SB2_2_27/i1_5 ), .A3(\SB2_2_27/i0_4 ), .ZN(
        \SB2_2_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_1/Component_Function_4/N4  ( .A1(\SB2_2_1/i1[9] ), .A2(
        \SB2_2_1/i1_5 ), .A3(\SB1_2_2/buf_output[4] ), .ZN(
        \SB2_2_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_14/Component_Function_1/N3  ( .A1(\SB2_2_14/i1_5 ), .A2(
        \SB2_2_14/i0[6] ), .A3(\SB2_2_14/i0[9] ), .ZN(
        \SB2_2_14/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_25/Component_Function_1/N1  ( .A1(\SB2_2_25/i0_3 ), .A2(
        \SB2_2_25/i1[9] ), .ZN(\SB2_2_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10282 ( .A1(\SB2_2_6/i0_3 ), .A2(\SB2_2_6/i0[10] ), .A3(
        \SB2_2_6/i0_4 ), .ZN(n4203) );
  NAND3_X1 U11463 ( .A1(\SB2_2_19/i0_0 ), .A2(\SB2_2_19/i0_3 ), .A3(
        \SB2_2_19/i0[7] ), .ZN(n4738) );
  NAND3_X1 \SB2_2_11/Component_Function_1/N2  ( .A1(\SB2_2_11/i0_3 ), .A2(
        \SB2_2_11/i1_7 ), .A3(\SB2_2_11/i0[8] ), .ZN(
        \SB2_2_11/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_12/Component_Function_0/N2  ( .A1(\SB2_2_12/i0[8] ), .A2(
        \SB2_2_12/i0[7] ), .A3(\SB2_2_12/i0[6] ), .ZN(
        \SB2_2_12/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_12/Component_Function_1/N2  ( .A1(\SB2_2_12/i0_3 ), .A2(
        \SB2_2_12/i1_7 ), .A3(\SB2_2_12/i0[8] ), .ZN(
        \SB2_2_12/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_6/Component_Function_0/N4  ( .A1(\SB2_2_6/i0[7] ), .A2(
        \SB2_2_6/i0_3 ), .A3(\SB2_2_6/i0_0 ), .ZN(
        \SB2_2_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_16/Component_Function_2/N3  ( .A1(\SB2_2_16/i0_3 ), .A2(
        \SB2_2_16/i0[8] ), .A3(\SB2_2_16/i0[9] ), .ZN(
        \SB2_2_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_11/Component_Function_2/N2  ( .A1(\SB2_2_11/i0_3 ), .A2(
        \SB2_2_11/i0[10] ), .A3(\SB2_2_11/i0[6] ), .ZN(
        \SB2_2_11/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_13/Component_Function_1/N1  ( .A1(\SB2_2_13/i0_3 ), .A2(
        \SB2_2_13/i1[9] ), .ZN(\SB2_2_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3101 ( .A1(\SB2_2_13/i0[10] ), .A2(\SB2_2_13/i0[9] ), .A3(
        \SB2_2_13/i0_3 ), .ZN(\SB2_2_13/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_17/Component_Function_2/N2  ( .A1(\SB2_2_17/i0_3 ), .A2(
        \SB2_2_17/i0[10] ), .A3(\SB2_2_17/i0[6] ), .ZN(
        \SB2_2_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U12623 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0[8] ), .A3(
        \SB2_2_16/i1_7 ), .ZN(n5374) );
  INV_X1 \SB1_3_4/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[163] ), .ZN(
        \SB1_3_4/i1_7 ) );
  BUF_X2 \SB1_3_28/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[18] ), .Z(
        \SB1_3_28/i0[9] ) );
  BUF_X2 U2006 ( .I(\MC_ARK_ARC_1_2/buf_output[168] ), .Z(\SB1_3_3/i0[9] ) );
  INV_X1 \SB1_3_1/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[180] ), .ZN(
        \SB1_3_1/i3[0] ) );
  INV_X1 \SB1_3_15/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[97] ), .ZN(
        \SB1_3_15/i1_7 ) );
  INV_X1 \SB1_3_20/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[71] ), .ZN(
        \SB1_3_20/i1_5 ) );
  INV_X1 \SB1_3_5/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[156] ), .ZN(
        \SB1_3_5/i3[0] ) );
  INV_X1 \SB1_3_23/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[49] ), .ZN(
        \SB1_3_23/i1_7 ) );
  INV_X1 \SB1_3_5/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[157] ), .ZN(
        \SB1_3_5/i1_7 ) );
  BUF_X2 U9763 ( .I(\MC_ARK_ARC_1_2/buf_output[30] ), .Z(\SB1_3_26/i0[9] ) );
  INV_X1 \SB1_3_29/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[12] ), .ZN(
        \SB1_3_29/i3[0] ) );
  BUF_X2 U5033 ( .I(\MC_ARK_ARC_1_2/buf_output[67] ), .Z(\SB1_3_20/i0[6] ) );
  INV_X1 U2825 ( .I(\MC_ARK_ARC_1_2/buf_output[19] ), .ZN(\SB1_3_28/i1_7 ) );
  CLKBUF_X2 U2007 ( .I(\MC_ARK_ARC_1_2/buf_output[127] ), .Z(\SB1_3_10/i0[6] )
         );
  BUF_X2 U9624 ( .I(\MC_ARK_ARC_1_2/buf_output[49] ), .Z(\SB1_3_23/i0[6] ) );
  BUF_X2 U1374 ( .I(\MC_ARK_ARC_1_2/buf_output[187] ), .Z(\SB1_3_0/i0[6] ) );
  CLKBUF_X2 U5206 ( .I(\MC_ARK_ARC_1_2/buf_output[184] ), .Z(\SB1_3_1/i0_4 )
         );
  BUF_X2 U9804 ( .I(\MC_ARK_ARC_1_2/buf_output[92] ), .Z(\SB1_3_16/i0_0 ) );
  BUF_X2 U3450 ( .I(\MC_ARK_ARC_1_2/buf_output[182] ), .Z(\SB1_3_1/i0_0 ) );
  BUF_X2 U3279 ( .I(\MC_ARK_ARC_1_2/buf_output[133] ), .Z(\SB1_3_9/i0[6] ) );
  BUF_X2 \SB1_3_24/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[47] ), .Z(
        \SB1_3_24/i0_3 ) );
  INV_X1 U5241 ( .I(\MC_ARK_ARC_1_2/buf_output[103] ), .ZN(\SB1_3_14/i1_7 ) );
  NAND3_X1 U896 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i0[7] ), .A3(
        \SB1_3_5/i0_0 ), .ZN(n2273) );
  NAND3_X1 U7212 ( .A1(\SB1_3_18/i0_3 ), .A2(\SB1_3_18/i0[8] ), .A3(
        \SB1_3_18/i0[9] ), .ZN(\SB1_3_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_9/Component_Function_3/N1  ( .A1(\SB1_3_9/i1[9] ), .A2(
        \SB1_3_9/i0_3 ), .A3(\SB1_3_9/i0[6] ), .ZN(
        \SB1_3_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1372 ( .A1(\SB1_3_12/i0[8] ), .A2(\SB1_3_12/i0[7] ), .A3(
        \SB1_3_12/i0[6] ), .ZN(\SB1_3_12/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N3  ( .A1(\SB1_3_28/i0[9] ), .A2(
        \SB1_3_28/i0[10] ), .A3(\SB1_3_28/i0_3 ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[2] ) );
  INV_X2 \SB1_3_17/INV_4  ( .I(\SB1_3_17/i0_4 ), .ZN(\SB1_3_17/i0[7] ) );
  NAND3_X1 \SB1_3_16/Component_Function_4/N2  ( .A1(\SB1_3_16/i3[0] ), .A2(
        \SB1_3_16/i0_0 ), .A3(\SB1_3_16/i1_7 ), .ZN(
        \SB1_3_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_17/Component_Function_3/N4  ( .A1(\SB1_3_17/i1_5 ), .A2(
        \SB1_3_17/i0[8] ), .A3(\SB1_3_17/i3[0] ), .ZN(
        \SB1_3_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3800 ( .A1(\SB1_3_9/i1_5 ), .A2(\SB1_3_9/i0[8] ), .A3(
        \SB1_3_9/i3[0] ), .ZN(\SB1_3_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1300 ( .A1(\SB1_3_17/i1[9] ), .A2(\SB1_3_17/i1_7 ), .A3(
        \SB1_3_17/i0[10] ), .ZN(\SB1_3_17/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 \SB1_3_29/Component_Function_3/N2  ( .A1(\SB1_3_29/i0_0 ), .A2(
        \SB1_3_29/i0_3 ), .A3(\SB1_3_29/i0_4 ), .ZN(
        \SB1_3_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N4  ( .A1(\SB1_3_28/i1[9] ), .A2(
        \SB1_3_28/i1_5 ), .A3(\SB1_3_28/i0_4 ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U3806 ( .A1(\SB1_3_6/i0_0 ), .A2(\SB1_3_6/i3[0] ), .ZN(
        \SB1_3_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U11500 ( .A1(\SB1_3_31/i0[9] ), .A2(\SB1_3_31/i1_5 ), .A3(
        \SB1_3_31/i0[6] ), .ZN(n4762) );
  NAND2_X1 \SB1_3_11/Component_Function_5/N1  ( .A1(\SB1_3_11/i0_0 ), .A2(
        \SB1_3_11/i3[0] ), .ZN(\SB1_3_11/Component_Function_5/NAND4_in[0] ) );
  INV_X1 \SB1_3_30/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[7] ), .ZN(
        \SB1_3_30/i1_7 ) );
  NAND3_X1 U857 ( .A1(\SB1_3_7/i0_4 ), .A2(\SB1_3_7/i1[9] ), .A3(
        \SB1_3_7/i1_5 ), .ZN(n1825) );
  NAND3_X1 U8468 ( .A1(\SB1_3_1/i0_0 ), .A2(\SB1_3_1/i0[9] ), .A3(
        \SB1_3_1/i0[8] ), .ZN(\SB1_3_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_15/Component_Function_1/N3  ( .A1(\SB1_3_15/i1_5 ), .A2(
        \SB1_3_15/i0[6] ), .A3(\SB1_3_15/i0[9] ), .ZN(
        \SB1_3_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U859 ( .A1(\SB1_3_6/i0_3 ), .A2(\SB1_3_6/i0_4 ), .A3(
        \SB1_3_6/i1[9] ), .ZN(n2150) );
  NAND3_X1 \SB1_3_15/Component_Function_5/N3  ( .A1(n5431), .A2(
        \SB1_3_15/i0_4 ), .A3(\SB1_3_15/i0_3 ), .ZN(
        \SB1_3_15/Component_Function_5/NAND4_in[2] ) );
  INV_X1 \SB1_3_25/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[36] ), .ZN(
        \SB1_3_25/i3[0] ) );
  BUF_X2 \SB1_3_22/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[55] ), .Z(
        \SB1_3_22/i0[6] ) );
  BUF_X2 U5239 ( .I(\MC_ARK_ARC_1_2/buf_output[181] ), .Z(\SB1_3_1/i0[6] ) );
  NAND3_X1 U8014 ( .A1(\SB1_3_7/i0_3 ), .A2(\SB1_3_7/i0_4 ), .A3(
        \SB1_3_7/i1[9] ), .ZN(\SB1_3_7/Component_Function_5/NAND4_in[2] ) );
  INV_X1 \SB1_3_6/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[151] ), .ZN(
        \SB1_3_6/i1_7 ) );
  NAND3_X1 \SB1_3_9/Component_Function_2/N2  ( .A1(\SB1_3_9/i0_3 ), .A2(
        \SB1_3_9/i0[10] ), .A3(\SB1_3_9/i0[6] ), .ZN(
        \SB1_3_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_15/Component_Function_4/N1  ( .A1(\SB1_3_15/i0[9] ), .A2(
        \SB1_3_15/i0_0 ), .A3(\SB1_3_15/i0[8] ), .ZN(
        \SB1_3_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U7657 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i1[9] ), .A3(
        \SB1_3_5/i0[6] ), .ZN(\SB1_3_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U8038 ( .A1(\SB1_3_7/i0_0 ), .A2(\SB1_3_7/i0_3 ), .A3(
        \SB1_3_7/i0[7] ), .ZN(n4336) );
  NAND3_X1 U1692 ( .A1(\SB1_3_3/i0[8] ), .A2(\SB1_3_3/i0_4 ), .A3(
        \SB1_3_3/i1_7 ), .ZN(\SB1_3_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_13/Component_Function_0/N4  ( .A1(\SB1_3_13/i0[7] ), .A2(
        \SB1_3_13/i0_3 ), .A3(\SB1_3_13/i0_0 ), .ZN(
        \SB1_3_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_18/Component_Function_1/N4  ( .A1(\SB1_3_18/i1_7 ), .A2(
        \SB1_3_18/i0[8] ), .A3(\SB1_3_18/i0_4 ), .ZN(
        \SB1_3_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2750 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0_0 ), .A3(
        \SB1_3_23/i0[7] ), .ZN(n3699) );
  NAND3_X1 \SB1_3_7/Component_Function_1/N4  ( .A1(\SB1_3_7/i1_7 ), .A2(
        \SB1_3_7/i0[8] ), .A3(\SB1_3_7/i0_4 ), .ZN(
        \SB1_3_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_19/Component_Function_4/N3  ( .A1(\SB1_3_19/i0[9] ), .A2(
        \SB1_3_19/i0[10] ), .A3(\SB1_3_19/i0_3 ), .ZN(
        \SB1_3_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1166 ( .A1(\SB1_3_0/i0_3 ), .A2(\SB1_3_0/i0_4 ), .A3(
        \SB1_3_0/i0_0 ), .ZN(n3697) );
  NAND2_X1 \SB1_3_23/Component_Function_0/N1  ( .A1(\SB1_3_23/i0[10] ), .A2(
        \SB1_3_23/i0[9] ), .ZN(\SB1_3_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U4357 ( .A1(\SB1_3_27/i3[0] ), .A2(\SB1_3_27/i0[8] ), .A3(
        \SB1_3_27/i1_5 ), .ZN(n3887) );
  NAND3_X1 U897 ( .A1(\SB1_3_6/i0[10] ), .A2(\SB1_3_6/i1[9] ), .A3(
        \SB1_3_6/i1_7 ), .ZN(n3053) );
  NAND3_X1 U2312 ( .A1(\SB1_3_1/i1_7 ), .A2(\SB1_3_1/i0[8] ), .A3(
        \SB1_3_1/i0_4 ), .ZN(\SB1_3_1/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 U5504 ( .A1(\SB1_3_8/i0[9] ), .A2(\SB1_3_8/i0[10] ), .ZN(n3392) );
  NAND3_X1 \SB1_3_19/Component_Function_4/N4  ( .A1(\SB1_3_19/i1[9] ), .A2(
        \SB1_3_19/i1_5 ), .A3(\SB1_3_19/i0_4 ), .ZN(
        \SB1_3_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3636 ( .A1(\SB1_3_19/i0_0 ), .A2(\SB1_3_19/i0[7] ), .A3(
        \SB1_3_19/i0_3 ), .ZN(n996) );
  NAND3_X1 U3439 ( .A1(\SB1_3_18/i0[9] ), .A2(\SB1_3_18/i1_5 ), .A3(
        \SB1_3_18/i0[6] ), .ZN(\SB1_3_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U8605 ( .A1(\SB1_3_31/i0[9] ), .A2(n5441), .A3(\SB1_3_31/i0_0 ), 
        .ZN(\SB1_3_31/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_31/Component_Function_5/N1  ( .A1(\SB1_3_31/i0_0 ), .A2(
        \SB1_3_31/i3[0] ), .ZN(\SB1_3_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1317 ( .A1(\SB1_3_29/i0_0 ), .A2(\SB1_3_29/i3[0] ), .A3(
        \SB1_3_29/i1_7 ), .ZN(\SB1_3_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1184 ( .A1(\SB1_3_1/i1_5 ), .A2(\SB1_3_1/i0[6] ), .A3(
        \SB1_3_1/i0[9] ), .ZN(\SB1_3_1/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_25/Component_Function_5/N1  ( .A1(\SB1_3_25/i0_0 ), .A2(
        \SB1_3_25/i3[0] ), .ZN(\SB1_3_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U7070 ( .A1(\SB1_3_8/i0[9] ), .A2(\SB1_3_8/i1_5 ), .A3(
        \SB1_3_8/i0[6] ), .ZN(\SB1_3_8/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_19/Component_Function_5/N1  ( .A1(\SB1_3_19/i0_0 ), .A2(
        \SB1_3_19/i3[0] ), .ZN(\SB1_3_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U893 ( .A1(\SB1_3_6/i0_4 ), .A2(\SB1_3_6/i1[9] ), .A3(
        \SB1_3_6/i1_5 ), .ZN(\SB1_3_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3796 ( .A1(\SB1_3_29/i1_5 ), .A2(\SB1_3_29/i0[6] ), .A3(
        \SB1_3_29/i0[9] ), .ZN(\SB1_3_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1361 ( .A1(\SB1_3_16/i0[6] ), .A2(\SB1_3_16/i1[9] ), .A3(
        \SB1_3_16/i0_3 ), .ZN(n4732) );
  NAND3_X1 U1370 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i0[8] ), .A3(
        \SB1_3_12/i1_7 ), .ZN(\SB1_3_12/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1373 ( .A1(\SB1_3_12/i1_7 ), .A2(\SB1_3_12/i0[8] ), .A3(
        \SB1_3_12/i0_4 ), .ZN(\SB1_3_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U7658 ( .A1(\SB1_3_19/i0_3 ), .A2(\SB1_3_19/i0_4 ), .A3(
        \SB1_3_19/i1[9] ), .ZN(n2502) );
  NAND3_X1 U3842 ( .A1(\SB1_3_6/i0[6] ), .A2(\SB1_3_6/i1_5 ), .A3(
        \SB1_3_6/i0[9] ), .ZN(\SB1_3_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U6416 ( .A1(\SB1_3_6/i0_3 ), .A2(\SB1_3_6/i1[9] ), .A3(
        \SB1_3_6/i0[6] ), .ZN(\SB1_3_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U11207 ( .A1(\SB1_3_27/i0_3 ), .A2(\SB1_3_27/i0[9] ), .A3(
        \SB1_3_27/i0[8] ), .ZN(n4615) );
  NAND3_X1 \SB1_3_17/Component_Function_2/N2  ( .A1(\SB1_3_17/i0_3 ), .A2(
        \SB1_3_17/i0[10] ), .A3(\SB1_3_17/i0[6] ), .ZN(
        \SB1_3_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_25/Component_Function_4/N4  ( .A1(\SB1_3_25/i1[9] ), .A2(
        \SB1_3_25/i1_5 ), .A3(\SB1_3_25/i0_4 ), .ZN(
        \SB1_3_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U8174 ( .A1(\RI1[3][167] ), .A2(\SB1_3_4/i0[9] ), .A3(
        \SB1_3_4/i0[10] ), .ZN(n2786) );
  NAND3_X1 U2587 ( .A1(\SB1_3_7/i0[6] ), .A2(\SB1_3_7/i1_5 ), .A3(
        \SB1_3_7/i0[9] ), .ZN(\SB1_3_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3803 ( .A1(\SB1_3_0/i0[9] ), .A2(\SB1_3_0/i0[10] ), .A3(
        \SB1_3_0/i0_3 ), .ZN(\SB1_3_0/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_29/Component_Function_1/N1  ( .A1(\SB1_3_29/i0_3 ), .A2(
        \SB1_3_29/i1[9] ), .ZN(\SB1_3_29/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 U2756 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i1[9] ), .ZN(
        \SB1_3_23/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_16/Component_Function_1/N1  ( .A1(\SB1_3_16/i0_3 ), .A2(
        \SB1_3_16/i1[9] ), .ZN(\SB1_3_16/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_6/Component_Function_1/N1  ( .A1(\SB1_3_6/i0_3 ), .A2(
        \SB1_3_6/i1[9] ), .ZN(\SB1_3_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10395 ( .A1(\SB1_3_11/i0_4 ), .A2(\SB1_3_11/i0_0 ), .A3(
        \SB1_3_11/i1_5 ), .ZN(\SB1_3_11/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 U1312 ( .A1(\SB1_3_21/Component_Function_4/NAND4_in[1] ), .A2(n4710), .ZN(n5271) );
  NAND2_X1 \SB1_3_27/Component_Function_1/N1  ( .A1(\SB1_3_27/i0_3 ), .A2(
        \SB1_3_27/i1[9] ), .ZN(\SB1_3_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1331 ( .A1(\SB1_3_30/i0[10] ), .A2(\SB1_3_30/i0[9] ), .A3(
        \SB1_3_30/i0_3 ), .ZN(n5187) );
  NAND3_X1 U11621 ( .A1(\SB1_3_20/i0_4 ), .A2(\SB1_3_20/i0_3 ), .A3(
        \SB1_3_20/i1[9] ), .ZN(n4830) );
  NAND3_X1 U854 ( .A1(\SB1_3_29/i0_3 ), .A2(\SB1_3_29/i0[9] ), .A3(
        \SB1_3_29/i0[10] ), .ZN(\SB1_3_29/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 \SB1_3_21/Component_Function_2/N3  ( .A1(\SB1_3_21/i0_3 ), .A2(
        \SB1_3_21/i0[8] ), .A3(\SB1_3_21/i0[9] ), .ZN(
        \SB1_3_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_5/N3  ( .A1(\SB1_3_13/i1[9] ), .A2(
        \SB1_3_13/i0_4 ), .A3(\SB1_3_13/i0_3 ), .ZN(
        \SB1_3_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1223 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i0_4 ), .A3(
        \SB1_3_12/i1[9] ), .ZN(n4477) );
  NAND3_X1 U8815 ( .A1(\SB1_3_4/i0[10] ), .A2(\SB1_3_4/i0_0 ), .A3(
        \SB1_3_4/i0[6] ), .ZN(\SB1_3_4/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB1_3_27/INV_4  ( .I(\SB1_3_27/i0_4 ), .ZN(\SB1_3_27/i0[7] ) );
  NAND3_X1 U867 ( .A1(\SB1_3_27/i0[9] ), .A2(\SB1_3_27/i1_5 ), .A3(
        \SB1_3_27/i0[6] ), .ZN(n2030) );
  NAND3_X1 U1337 ( .A1(\SB1_3_17/i0[10] ), .A2(\SB1_3_17/i1[9] ), .A3(
        \SB1_3_17/i1_5 ), .ZN(n5215) );
  NAND3_X1 \SB1_3_3/Component_Function_3/N2  ( .A1(\SB1_3_3/i0_0 ), .A2(
        \SB1_3_3/i0_3 ), .A3(\SB1_3_3/i0_4 ), .ZN(
        \SB1_3_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U10688 ( .A1(\SB1_3_28/i0[6] ), .A2(\SB1_3_28/i0_3 ), .A3(
        \SB1_3_28/i1[9] ), .ZN(\SB1_3_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_13/Component_Function_2/N3  ( .A1(\SB1_3_13/i0_3 ), .A2(
        \SB1_3_13/i0[8] ), .A3(\SB1_3_13/i0[9] ), .ZN(
        \SB1_3_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2286 ( .A1(\SB1_3_5/i1_7 ), .A2(\SB1_3_5/i0[8] ), .A3(
        \SB1_3_5/i0_4 ), .ZN(\SB1_3_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1693 ( .A1(\SB1_3_3/i0[8] ), .A2(\SB1_3_3/i3[0] ), .A3(
        \SB1_3_3/i1_5 ), .ZN(\SB1_3_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_14/Component_Function_0/N4  ( .A1(\SB1_3_14/i0[7] ), .A2(
        \RI1[3][107] ), .A3(\SB1_3_14/i0_0 ), .ZN(
        \SB1_3_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U850 ( .A1(\SB1_3_21/i0_4 ), .A2(\SB1_3_21/i0[8] ), .A3(
        \SB1_3_21/i1_7 ), .ZN(n2880) );
  NAND3_X1 U3808 ( .A1(\SB1_3_7/i0[8] ), .A2(\SB1_3_7/i3[0] ), .A3(
        \SB1_3_7/i1_5 ), .ZN(n2884) );
  NAND3_X1 U10687 ( .A1(\SB1_3_18/i0[8] ), .A2(\SB1_3_18/i1_5 ), .A3(
        \SB1_3_18/i3[0] ), .ZN(n4595) );
  NAND3_X1 U6446 ( .A1(\SB1_3_8/i0[10] ), .A2(\SB1_3_8/i1[9] ), .A3(
        \SB1_3_8/i1_5 ), .ZN(\SB1_3_8/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_1/Component_Function_5/N1  ( .A1(\SB1_3_1/i0_0 ), .A2(
        \SB1_3_1/i3[0] ), .ZN(\SB1_3_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1294 ( .A1(\SB1_3_19/i0[10] ), .A2(\SB1_3_19/i1[9] ), .A3(
        \SB1_3_19/i1_7 ), .ZN(\SB1_3_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1221 ( .A1(\SB1_3_10/i0[9] ), .A2(\SB1_3_10/i0[6] ), .A3(
        \SB1_3_10/i0_4 ), .ZN(\SB1_3_10/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U866 ( .A1(\SB1_3_22/i0_0 ), .A2(\SB1_3_22/i3[0] ), .ZN(n895) );
  NAND2_X1 U11199 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i3[0] ), .ZN(
        \SB1_3_18/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U3843 ( .A1(\SB1_3_16/i3[0] ), .A2(\SB1_3_16/i0_0 ), .ZN(
        \SB1_3_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_5/N4  ( .A1(\SB1_3_26/i0[9] ), .A2(
        \SB1_3_26/i0[6] ), .A3(\SB1_3_26/i0_4 ), .ZN(
        \SB1_3_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1225 ( .A1(\SB1_3_30/i1[9] ), .A2(\SB1_3_30/i0_3 ), .A3(
        \SB1_3_30/i0[6] ), .ZN(\SB1_3_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U11813 ( .A1(\SB1_3_19/i0[10] ), .A2(\SB1_3_19/i0_3 ), .A3(
        \SB1_3_19/i0[6] ), .ZN(n4911) );
  NAND3_X1 \SB1_3_19/Component_Function_3/N2  ( .A1(\SB1_3_19/i0_0 ), .A2(
        \SB1_3_19/i0_3 ), .A3(\SB1_3_19/i0_4 ), .ZN(
        \SB1_3_19/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U2287 ( .A1(\SB1_3_20/i0_3 ), .A2(\SB1_3_20/i1[9] ), .ZN(
        \SB1_3_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U8661 ( .A1(\SB1_3_25/i0_0 ), .A2(\SB1_3_25/i1_5 ), .A3(
        \SB1_3_25/i0_4 ), .ZN(n3866) );
  NAND3_X1 U1260 ( .A1(\SB1_3_0/i1_7 ), .A2(\SB1_3_0/i0[8] ), .A3(
        \SB1_3_0/i0_4 ), .ZN(\SB1_3_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U6618 ( .A1(\SB1_3_16/i0[10] ), .A2(\SB1_3_16/i0_0 ), .A3(
        \SB1_3_16/i0[6] ), .ZN(\SB1_3_16/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_9/Component_Function_1/N4  ( .A1(\SB1_3_9/i1_7 ), .A2(
        \SB1_3_9/i0[8] ), .A3(\SB1_3_9/i0_4 ), .ZN(
        \SB1_3_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3819 ( .A1(\SB1_3_14/i1_5 ), .A2(\SB1_3_14/i0[6] ), .A3(
        \SB1_3_14/i0[9] ), .ZN(\SB1_3_14/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U1244 ( .A1(\SB1_3_29/Component_Function_4/NAND4_in[1] ), .A2(n807), 
        .ZN(n3311) );
  NAND3_X1 U5077 ( .A1(\SB1_3_29/i1_5 ), .A2(\SB1_3_29/i0[10] ), .A3(
        \SB1_3_29/i1[9] ), .ZN(\SB1_3_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2967 ( .A1(\SB1_3_29/i0_0 ), .A2(\SB1_3_29/i1_5 ), .A3(
        \SB1_3_29/i0_4 ), .ZN(n756) );
  NAND3_X1 \SB1_3_29/Component_Function_2/N2  ( .A1(\SB1_3_29/i0_3 ), .A2(
        \SB1_3_29/i0[10] ), .A3(\SB1_3_29/i0[6] ), .ZN(
        \SB1_3_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_11/Component_Function_3/N2  ( .A1(\SB1_3_11/i0_0 ), .A2(
        \SB1_3_11/i0_3 ), .A3(\SB1_3_11/i0_4 ), .ZN(
        \SB1_3_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_12/Component_Function_3/N2  ( .A1(\SB1_3_12/i0_0 ), .A2(
        \SB1_3_12/i0_3 ), .A3(\SB1_3_12/i0_4 ), .ZN(
        \SB1_3_12/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X2 U5221 ( .I(\SB1_3_12/buf_output[4] ), .Z(\SB2_3_11/i0_4 ) );
  BUF_X2 \SB2_3_21/BUF_3  ( .I(\SB1_3_23/buf_output[3] ), .Z(\SB2_3_21/i0[10] ) );
  NAND3_X1 U6847 ( .A1(\SB1_3_8/i0[9] ), .A2(\SB1_3_8/i0[8] ), .A3(
        \SB1_3_8/i0_3 ), .ZN(\SB1_3_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U12598 ( .A1(\SB1_3_20/i0_4 ), .A2(\SB1_3_20/i0[8] ), .A3(
        \SB1_3_20/i1_7 ), .ZN(n5356) );
  NAND3_X1 \SB1_3_13/Component_Function_1/N4  ( .A1(\SB1_3_13/i1_7 ), .A2(
        \SB1_3_13/i0[8] ), .A3(\SB1_3_13/i0_4 ), .ZN(
        \SB1_3_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_8/Component_Function_2/N2  ( .A1(\SB1_3_8/i0_3 ), .A2(
        \SB1_3_8/i0[10] ), .A3(\SB1_3_8/i0[6] ), .ZN(
        \SB1_3_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U10878 ( .A1(\SB1_3_28/i0_3 ), .A2(\SB1_3_28/i0_0 ), .A3(
        \SB1_3_28/i0_4 ), .ZN(\SB1_3_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11164 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB2_3_7/i1[9] ), .A3(
        \SB2_3_7/i0_4 ), .ZN(\SB2_3_7/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_6/Component_Function_5/N1  ( .A1(\SB2_3_6/i0_0 ), .A2(
        \SB2_3_6/i3[0] ), .ZN(\SB2_3_6/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U7071 ( .I(\SB2_3_4/i0[7] ), .ZN(\SB2_3_4/i0_4 ) );
  NAND2_X1 \SB2_3_11/Component_Function_5/N1  ( .A1(\SB2_3_11/i0_0 ), .A2(
        \SB2_3_11/i3[0] ), .ZN(\SB2_3_11/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_0/Component_Function_5/N1  ( .A1(\SB2_3_0/i0_0 ), .A2(
        \SB2_3_0/i3[0] ), .ZN(\SB2_3_0/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_27/Component_Function_5/N1  ( .A1(\SB2_3_27/i0_0 ), .A2(
        \SB2_3_27/i3[0] ), .ZN(\SB2_3_27/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 \SB2_3_14/BUF_0  ( .I(\SB1_3_19/buf_output[0] ), .Z(\SB2_3_14/i0[9] )
         );
  BUF_X2 \SB2_3_3/BUF_0  ( .I(\SB1_3_8/buf_output[0] ), .Z(\SB2_3_3/i0[9] ) );
  BUF_X2 \SB2_3_4/BUF_0  ( .I(\SB1_3_9/buf_output[0] ), .Z(\SB2_3_4/i0[9] ) );
  CLKBUF_X2 \SB2_3_13/BUF_0  ( .I(\SB1_3_18/buf_output[0] ), .Z(
        \SB2_3_13/i0[9] ) );
  CLKBUF_X2 \SB2_3_12/BUF_1  ( .I(\SB1_3_16/buf_output[1] ), .Z(
        \SB2_3_12/i0[6] ) );
  INV_X1 U1861 ( .I(\SB1_3_3/buf_output[5] ), .ZN(\SB2_3_3/i1_5 ) );
  INV_X1 \SB2_3_23/INV_0  ( .I(\SB1_3_28/buf_output[0] ), .ZN(\SB2_3_23/i3[0] ) );
  INV_X2 \SB2_3_3/INV_4  ( .I(\SB2_3_3/i0_4 ), .ZN(\SB2_3_3/i0[7] ) );
  NAND2_X1 U2471 ( .A1(\SB2_3_23/i0_0 ), .A2(\SB2_3_23/i3[0] ), .ZN(
        \SB2_3_23/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_30/Component_Function_5/N1  ( .A1(\SB2_3_30/i0_0 ), .A2(
        \SB2_3_30/i3[0] ), .ZN(\SB2_3_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_2/N1  ( .A1(\SB2_3_7/i1_5 ), .A2(
        \SB2_3_7/i0[10] ), .A3(\SB2_3_7/i1[9] ), .ZN(
        \SB2_3_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U10150 ( .A1(\SB2_3_29/i0_3 ), .A2(\SB2_3_29/i0_4 ), .A3(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_5/NAND4_in[2] ) );
  INV_X1 \SB2_3_14/INV_1  ( .I(\SB1_3_18/buf_output[1] ), .ZN(\SB2_3_14/i1_7 )
         );
  NAND3_X1 \SB2_3_14/Component_Function_5/N4  ( .A1(\SB2_3_14/i0[9] ), .A2(
        \SB2_3_14/i0[6] ), .A3(\SB2_3_14/i0_4 ), .ZN(
        \SB2_3_14/Component_Function_5/NAND4_in[3] ) );
  INV_X1 \SB2_3_17/INV_1  ( .I(\SB1_3_21/buf_output[1] ), .ZN(\SB2_3_17/i1_7 )
         );
  NAND2_X1 \SB2_3_29/Component_Function_5/N1  ( .A1(\SB2_3_29/i0_0 ), .A2(
        \SB2_3_29/i3[0] ), .ZN(\SB2_3_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U7712 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i1_5 ), .A3(
        \SB2_3_19/i1[9] ), .ZN(\SB2_3_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U11993 ( .A1(\SB2_3_19/i0_0 ), .A2(\SB2_3_19/i1_5 ), .A3(
        \SB1_3_20/buf_output[4] ), .ZN(n5075) );
  NAND3_X1 U7667 ( .A1(n6552), .A2(\SB2_3_29/i0_0 ), .A3(\SB2_3_29/i0[10] ), 
        .ZN(n3700) );
  NAND3_X1 U4314 ( .A1(\SB2_3_12/i0_3 ), .A2(\SB2_3_12/i1[9] ), .A3(n592), 
        .ZN(\SB2_3_12/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U9787 ( .I(\SB1_3_2/buf_output[1] ), .ZN(\SB2_3_30/i1_7 ) );
  INV_X1 \SB2_3_11/INV_1  ( .I(\SB1_3_15/buf_output[1] ), .ZN(\SB2_3_11/i1_7 )
         );
  CLKBUF_X2 \SB2_3_5/BUF_0  ( .I(\SB1_3_10/buf_output[0] ), .Z(\SB2_3_5/i0[9] ) );
  CLKBUF_X2 \SB2_3_22/BUF_1  ( .I(\SB1_3_26/buf_output[1] ), .Z(
        \SB2_3_22/i0[6] ) );
  BUF_X2 \SB2_3_16/BUF_0  ( .I(\SB1_3_21/buf_output[0] ), .Z(\SB2_3_16/i0[9] )
         );
  BUF_X2 U2313 ( .I(\SB1_3_9/buf_output[1] ), .Z(\SB2_3_5/i0[6] ) );
  INV_X2 U6053 ( .I(n1763), .ZN(\RI3[3][58] ) );
  INV_X2 U9160 ( .I(n4081), .ZN(\SB2_3_26/i0_4 ) );
  INV_X1 \SB2_3_6/INV_1  ( .I(\SB1_3_10/buf_output[1] ), .ZN(\SB2_3_6/i1_7 )
         );
  INV_X1 \SB2_3_11/INV_5  ( .I(\SB1_3_11/buf_output[5] ), .ZN(\SB2_3_11/i1_5 )
         );
  NAND3_X1 U6090 ( .A1(\SB2_3_22/i0_3 ), .A2(\SB2_3_22/i0[10] ), .A3(
        \RI3[3][58] ), .ZN(n2033) );
  NAND3_X1 U801 ( .A1(\SB2_3_29/i0[9] ), .A2(\SB2_3_29/i0_3 ), .A3(
        \SB2_3_29/i0[8] ), .ZN(\SB2_3_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U10602 ( .A1(\SB2_3_25/i0[10] ), .A2(\SB2_3_25/i1_5 ), .A3(
        \SB2_3_25/i1[9] ), .ZN(\SB2_3_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_4/N1  ( .A1(\SB2_3_12/i0[9] ), .A2(
        \SB2_3_12/i0_0 ), .A3(\SB2_3_12/i0[8] ), .ZN(
        \SB2_3_12/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_15/Component_Function_1/N1  ( .A1(\SB2_3_15/i0_3 ), .A2(
        \SB2_3_15/i1[9] ), .ZN(\SB2_3_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_3/N1  ( .A1(\SB2_3_7/i1[9] ), .A2(
        \SB2_3_7/i0_3 ), .A3(\SB2_3_7/i0[6] ), .ZN(
        \SB2_3_7/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_5/Component_Function_0/N1  ( .A1(\SB2_3_5/i0[10] ), .A2(
        \SB2_3_5/i0[9] ), .ZN(\SB2_3_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3875 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0_0 ), .A3(
        \SB2_3_18/i0[7] ), .ZN(n2061) );
  NAND3_X1 \SB2_3_18/Component_Function_0/N2  ( .A1(\SB2_3_18/i0[8] ), .A2(
        \SB2_3_18/i0[7] ), .A3(\SB2_3_18/i0[6] ), .ZN(
        \SB2_3_18/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1118 ( .A1(\SB2_3_14/i0[9] ), .A2(\SB2_3_14/i0_3 ), .A3(
        \SB2_3_14/i0[10] ), .ZN(\SB2_3_14/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 \SB2_3_8/Component_Function_4/N2  ( .A1(\SB2_3_8/i3[0] ), .A2(
        \SB2_3_8/i0_0 ), .A3(\SB2_3_8/i1_7 ), .ZN(
        \SB2_3_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U9168 ( .A1(\SB2_3_24/i3[0] ), .A2(\SB2_3_24/i1_5 ), .A3(
        \SB2_3_24/i0[8] ), .ZN(n3924) );
  NAND3_X1 U11812 ( .A1(\SB2_3_16/i0[10] ), .A2(\SB2_3_16/i0_0 ), .A3(
        \SB2_3_16/i0[6] ), .ZN(n4909) );
  NAND3_X1 \SB2_3_22/Component_Function_3/N4  ( .A1(\SB2_3_22/i1_5 ), .A2(
        \SB2_3_22/i0[8] ), .A3(\SB2_3_22/i3[0] ), .ZN(
        \SB2_3_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U793 ( .A1(\SB2_3_12/i0_3 ), .A2(n592), .A3(\SB2_3_12/i0[10] ), 
        .ZN(\SB2_3_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U5429 ( .A1(\SB2_3_21/i0[6] ), .A2(n6716), .A3(\SB2_3_21/i0[8] ), 
        .ZN(\SB2_3_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_14/Component_Function_4/N4  ( .A1(\SB2_3_14/i1[9] ), .A2(
        \SB2_3_14/i1_5 ), .A3(\SB2_3_14/i0_4 ), .ZN(
        \SB2_3_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1006 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0[9] ), .A3(
        \SB2_3_10/i0[8] ), .ZN(\SB2_3_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U6533 ( .A1(\SB2_3_21/i0[8] ), .A2(\SB2_3_21/i1_7 ), .A3(
        \RI3[3][64] ), .ZN(\SB2_3_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_16/Component_Function_0/N2  ( .A1(\SB2_3_16/i0[8] ), .A2(
        \SB2_3_16/i0[7] ), .A3(\SB2_3_16/i0[6] ), .ZN(
        \SB2_3_16/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_25/Component_Function_1/N4  ( .A1(\SB2_3_25/i1_7 ), .A2(
        \SB2_3_25/i0[8] ), .A3(\SB2_3_25/i0_4 ), .ZN(
        \SB2_3_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U6229 ( .A1(\SB2_3_19/i1_7 ), .A2(\SB1_3_20/buf_output[4] ), .A3(
        \SB2_3_19/i0[8] ), .ZN(n2239) );
  NAND3_X1 U10257 ( .A1(n6274), .A2(\SB2_3_29/i0_0 ), .A3(\SB2_3_29/i0_3 ), 
        .ZN(\SB2_3_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U11301 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0_0 ), .A3(
        \SB2_3_10/i0[7] ), .ZN(n4664) );
  NAND2_X1 \SB2_3_10/Component_Function_5/N1  ( .A1(\SB2_3_10/i0_0 ), .A2(
        \SB2_3_10/i3[0] ), .ZN(\SB2_3_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_4/N1  ( .A1(\SB2_3_21/i0[9] ), .A2(
        \SB2_3_21/i0_0 ), .A3(\SB2_3_21/i0[8] ), .ZN(
        \SB2_3_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_1/N3  ( .A1(\SB2_3_14/i1_5 ), .A2(
        \SB2_3_14/i0[6] ), .A3(\SB2_3_14/i0[9] ), .ZN(
        \SB2_3_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4048 ( .A1(\SB2_3_21/i1[9] ), .A2(\RI3[3][64] ), .A3(
        \SB2_3_21/i1_5 ), .ZN(n1144) );
  NAND3_X1 \SB2_3_13/Component_Function_3/N3  ( .A1(\SB2_3_13/i1[9] ), .A2(
        \SB2_3_13/i1_7 ), .A3(\SB2_3_13/i0[10] ), .ZN(
        \SB2_3_13/Component_Function_3/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_9/Component_Function_5/N1  ( .A1(\SB2_3_9/i0_0 ), .A2(
        \SB2_3_9/i3[0] ), .ZN(\SB2_3_9/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_13/Component_Function_5/N1  ( .A1(\SB2_3_13/i0_0 ), .A2(
        \SB2_3_13/i3[0] ), .ZN(\SB2_3_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_4/N4  ( .A1(\SB2_3_9/i1[9] ), .A2(
        \SB2_3_9/i1_5 ), .A3(\SB1_3_10/buf_output[4] ), .ZN(
        \SB2_3_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4265 ( .A1(\SB2_3_29/i3[0] ), .A2(\SB2_3_29/i0[8] ), .A3(
        \SB2_3_29/i1_5 ), .ZN(\SB2_3_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2800 ( .A1(\SB2_3_23/i0_4 ), .A2(\SB2_3_23/i0_0 ), .A3(
        \SB2_3_23/i1_5 ), .ZN(n1389) );
  NAND3_X1 \SB2_3_12/Component_Function_0/N4  ( .A1(n7586), .A2(
        \SB2_3_12/i0_3 ), .A3(\SB2_3_12/i0_0 ), .ZN(
        \SB2_3_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_9/Component_Function_1/N3  ( .A1(\SB2_3_9/i1_5 ), .A2(
        \SB2_3_9/i0[6] ), .A3(\SB2_3_9/i0[9] ), .ZN(
        \SB2_3_9/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_13/Component_Function_0/N1  ( .A1(\SB2_3_13/i0[10] ), .A2(
        \SB2_3_13/i0[9] ), .ZN(\SB2_3_13/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_12/Component_Function_1/N1  ( .A1(\SB2_3_12/i0_3 ), .A2(
        \SB2_3_12/i1[9] ), .ZN(\SB2_3_12/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_28/Component_Function_1/N1  ( .A1(\SB2_3_28/i0_3 ), .A2(
        \SB2_3_28/i1[9] ), .ZN(\SB2_3_28/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_24/Component_Function_1/N1  ( .A1(\SB2_3_24/i0_3 ), .A2(
        \SB2_3_24/i1[9] ), .ZN(\SB2_3_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3422 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i1[9] ), .A3(
        \SB2_3_10/i0[6] ), .ZN(\SB2_3_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_2/Component_Function_1/N4  ( .A1(\SB2_3_2/i1_7 ), .A2(
        \SB2_3_2/i0[8] ), .A3(\SB2_3_2/i0_4 ), .ZN(
        \SB2_3_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_3/N1  ( .A1(\SB2_3_12/i1[9] ), .A2(
        \SB2_3_12/i0_3 ), .A3(\SB2_3_12/i0[6] ), .ZN(
        \SB2_3_12/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_22/Component_Function_0/N1  ( .A1(\SB2_3_22/i0[10] ), .A2(
        \SB2_3_22/i0[9] ), .ZN(\SB2_3_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U2916 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0[10] ), .A3(
        \SB2_3_31/i0_4 ), .ZN(\SB2_3_31/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_10/Component_Function_1/N1  ( .A1(\SB2_3_10/i0_3 ), .A2(
        \SB2_3_10/i1[9] ), .ZN(\SB2_3_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3851 ( .A1(\SB2_3_6/i1_5 ), .A2(\SB2_3_6/i0[6] ), .A3(
        \SB2_3_6/i0[9] ), .ZN(\SB2_3_6/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_19/Component_Function_0/N1  ( .A1(\SB2_3_19/i0[10] ), .A2(
        \SB2_3_19/i0[9] ), .ZN(\SB2_3_19/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_29/Component_Function_0/N1  ( .A1(\SB2_3_29/i0[10] ), .A2(
        \SB2_3_29/i0[9] ), .ZN(\SB2_3_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U822 ( .A1(\SB2_3_22/i0[9] ), .A2(\SB2_3_22/i0[6] ), .A3(
        \RI3[3][58] ), .ZN(n2694) );
  NAND3_X1 \SB2_3_25/Component_Function_0/N2  ( .A1(\SB2_3_25/i0[8] ), .A2(
        \SB2_3_25/i0[7] ), .A3(\SB2_3_25/i0[6] ), .ZN(
        \SB2_3_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U8258 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i0[10] ), .A3(
        \SB2_3_24/i0_4 ), .ZN(n3794) );
  NAND3_X1 U1085 ( .A1(\SB2_3_28/i0_0 ), .A2(\SB2_3_28/i0[6] ), .A3(
        \SB2_3_28/i0[10] ), .ZN(\SB2_3_28/Component_Function_5/NAND4_in[1] )
         );
  NAND2_X1 \SB2_3_12/Component_Function_0/N1  ( .A1(\SB2_3_12/i0[10] ), .A2(
        \SB2_3_12/i0[9] ), .ZN(\SB2_3_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U4939 ( .A1(\SB2_3_14/i0_4 ), .A2(\SB2_3_14/i1_7 ), .A3(
        \SB2_3_14/i0[8] ), .ZN(\SB2_3_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_5/Component_Function_2/N1  ( .A1(\SB2_3_5/i1_5 ), .A2(
        \SB2_3_5/i0[10] ), .A3(\SB2_3_5/i1[9] ), .ZN(
        \SB2_3_5/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_9/Component_Function_1/N1  ( .A1(\SB2_3_9/i0_3 ), .A2(
        \SB2_3_9/i1[9] ), .ZN(\SB2_3_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_1/N3  ( .A1(\SB2_3_10/i1_5 ), .A2(
        \SB2_3_10/i0[6] ), .A3(\SB2_3_10/i0[9] ), .ZN(
        \SB2_3_10/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_10/Component_Function_0/N1  ( .A1(\SB2_3_10/i0[10] ), .A2(
        \SB2_3_10/i0[9] ), .ZN(\SB2_3_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_17/Component_Function_5/N1  ( .A1(\SB2_3_17/i0_0 ), .A2(
        \SB2_3_17/i3[0] ), .ZN(\SB2_3_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_3/N3  ( .A1(\SB2_3_26/i1[9] ), .A2(
        \SB2_3_26/i1_7 ), .A3(\SB2_3_26/i0[10] ), .ZN(
        \SB2_3_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_12/Component_Function_2/N2  ( .A1(\SB2_3_12/i0_3 ), .A2(
        \SB2_3_12/i0[10] ), .A3(\SB2_3_12/i0[6] ), .ZN(
        \SB2_3_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_5/Component_Function_1/N2  ( .A1(\SB2_3_5/i0_3 ), .A2(
        \SB2_3_5/i1_7 ), .A3(\SB2_3_5/i0[8] ), .ZN(
        \SB2_3_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_14/Component_Function_3/N1  ( .A1(\SB2_3_14/i1[9] ), .A2(
        \SB2_3_14/i0_3 ), .A3(\SB2_3_14/i0[6] ), .ZN(
        \SB2_3_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U805 ( .A1(\SB2_3_2/i0_0 ), .A2(\SB2_3_2/i3[0] ), .A3(
        \SB2_3_2/i1_7 ), .ZN(\SB2_3_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_2/Component_Function_4/N4  ( .A1(\SB2_3_2/i1[9] ), .A2(
        \SB2_3_2/i1_5 ), .A3(\SB2_3_2/i0_4 ), .ZN(
        \SB2_3_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_13/Component_Function_4/N2  ( .A1(\SB2_3_13/i3[0] ), .A2(
        \SB2_3_13/i0_0 ), .A3(\SB2_3_13/i1_7 ), .ZN(
        \SB2_3_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_14/Component_Function_0/N2  ( .A1(\SB2_3_14/i0[8] ), .A2(
        \SB2_3_14/i0[7] ), .A3(\SB2_3_14/i0[6] ), .ZN(
        \SB2_3_14/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3881 ( .A1(\SB2_3_24/i0[9] ), .A2(\SB2_3_24/i0[10] ), .A3(
        \SB2_3_24/i0_3 ), .ZN(\SB2_3_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1055 ( .A1(\SB2_3_11/i0[10] ), .A2(\SB2_3_11/i1_7 ), .A3(
        \SB2_3_11/i1[9] ), .ZN(n5239) );
  NAND3_X1 U12394 ( .A1(\SB2_3_5/i0[10] ), .A2(\SB2_3_5/i1_7 ), .A3(
        \SB2_3_5/i1[9] ), .ZN(\SB2_3_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_12/Component_Function_2/N4  ( .A1(\SB2_3_12/i1_5 ), .A2(
        \SB2_3_12/i0_0 ), .A3(n592), .ZN(
        \SB2_3_12/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_4/Component_Function_2/N1  ( .A1(\SB2_3_4/i1_5 ), .A2(
        \SB2_3_4/i0[10] ), .A3(\SB2_3_4/i1[9] ), .ZN(
        \SB2_3_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1068 ( .A1(\SB2_3_1/i0[9] ), .A2(\SB2_3_1/i1_5 ), .A3(
        \SB2_3_1/i0[6] ), .ZN(n3674) );
  NAND3_X1 \SB2_3_3/Component_Function_3/N1  ( .A1(\SB2_3_3/i1[9] ), .A2(
        \SB2_3_3/i0_3 ), .A3(\SB2_3_3/i0[6] ), .ZN(
        \SB2_3_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_3/N1  ( .A1(\SB2_3_0/i1[9] ), .A2(
        \SB2_3_0/i0_3 ), .A3(\SB2_3_0/i0[6] ), .ZN(
        \SB2_3_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10517 ( .A1(\SB2_3_0/i0[10] ), .A2(\SB2_3_0/i1[9] ), .A3(
        \SB2_3_0/i1_7 ), .ZN(\SB2_3_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_3/Component_Function_3/N2  ( .A1(\SB2_3_3/i0_0 ), .A2(
        \SB2_3_3/i0_3 ), .A3(\SB2_3_3/i0_4 ), .ZN(
        \SB2_3_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11573 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0[10] ), .A3(
        \SB2_3_10/i0[9] ), .ZN(n4794) );
  NAND2_X1 \SB2_3_5/Component_Function_1/N1  ( .A1(\SB2_3_5/i0_3 ), .A2(
        \SB2_3_5/i1[9] ), .ZN(\SB2_3_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1030 ( .A1(\SB2_3_2/i0_0 ), .A2(\SB2_3_2/i0_3 ), .A3(
        \SB2_3_2/i0[7] ), .ZN(n4741) );
  NAND3_X1 \SB2_3_14/Component_Function_0/N3  ( .A1(\SB2_3_14/i0[10] ), .A2(
        \SB2_3_14/i0_4 ), .A3(\SB2_3_14/i0_3 ), .ZN(
        \SB2_3_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U10838 ( .A1(\SB2_3_2/i0[10] ), .A2(\SB2_3_2/i0_3 ), .A3(
        \SB2_3_2/i0_4 ), .ZN(\SB2_3_2/Component_Function_0/NAND4_in[2] ) );
  BUF_X2 U9134 ( .I(\SB2_3_29/buf_output[0] ), .Z(\RI5[3][42] ) );
  BUF_X2 U8283 ( .I(\SB2_3_23/buf_output[4] ), .Z(\RI5[3][58] ) );
  BUF_X2 U789 ( .I(\SB2_3_5/buf_output[1] ), .Z(\RI5[3][181] ) );
  BUF_X2 U2377 ( .I(\MC_ARK_ARC_1_3/buf_output[24] ), .Z(\SB1_4_27/i0[9] ) );
  NAND3_X1 \SB1_4_6/Component_Function_4/N1  ( .A1(\SB1_4_6/i0[9] ), .A2(
        \SB1_4_6/i0_0 ), .A3(\SB1_4_6/i0[8] ), .ZN(
        \SB1_4_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U8483 ( .A1(\SB1_4_31/i0_3 ), .A2(\SB1_4_31/i0[9] ), .A3(
        \SB1_4_31/i0[10] ), .ZN(n2960) );
  NAND3_X1 \SB1_4_17/Component_Function_0/N4  ( .A1(\SB1_4_17/i0[7] ), .A2(
        \SB1_4_17/i0_3 ), .A3(\SB1_4_17/i0_0 ), .ZN(
        \SB1_4_17/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X2 \SB1_4_4/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[163] ), .Z(
        \SB1_4_4/i0[6] ) );
  INV_X1 U7037 ( .I(\MC_ARK_ARC_1_3/buf_output[179] ), .ZN(\SB1_4_2/i1_5 ) );
  NAND3_X1 \SB1_4_16/Component_Function_1/N4  ( .A1(\SB1_4_16/i1_7 ), .A2(
        \SB1_4_16/i0[8] ), .A3(\SB1_4_16/i0_4 ), .ZN(
        \SB1_4_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U844 ( .A1(\SB1_4_6/i0_0 ), .A2(\SB1_4_6/i3[0] ), .A3(
        \SB1_4_6/i1_7 ), .ZN(n4186) );
  INV_X1 U3148 ( .I(\MC_ARK_ARC_1_3/buf_output[79] ), .ZN(\SB1_4_18/i1_7 ) );
  INV_X1 U1925 ( .I(\MC_ARK_ARC_1_3/buf_output[103] ), .ZN(\SB1_4_14/i1_7 ) );
  INV_X1 U2168 ( .I(\MC_ARK_ARC_1_3/buf_output[174] ), .ZN(\SB1_4_2/i3[0] ) );
  INV_X1 \SB1_4_1/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[180] ), .ZN(
        \SB1_4_1/i3[0] ) );
  BUF_X2 U3427 ( .I(\MC_ARK_ARC_1_3/buf_output[121] ), .Z(\SB1_4_11/i0[6] ) );
  NAND2_X1 \SB1_4_16/Component_Function_1/N1  ( .A1(\SB1_4_16/i0_3 ), .A2(
        \SB1_4_16/i1[9] ), .ZN(\SB1_4_16/Component_Function_1/NAND4_in[0] ) );
  INV_X1 \SB1_4_0/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[186] ), .ZN(
        \SB1_4_0/i3[0] ) );
  INV_X1 \SB1_4_30/INV_5  ( .I(n3993), .ZN(\SB1_4_30/i1_5 ) );
  INV_X1 U3923 ( .I(\MC_ARK_ARC_1_3/buf_output[31] ), .ZN(\SB1_4_26/i1_7 ) );
  BUF_X2 U1721 ( .I(\MC_ARK_ARC_1_3/buf_output[61] ), .Z(\SB1_4_21/i0[6] ) );
  BUF_X2 U5086 ( .I(\MC_ARK_ARC_1_3/buf_output[175] ), .Z(\SB1_4_2/i0[6] ) );
  BUF_X2 \SB1_4_7/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[145] ), .Z(
        \SB1_4_7/i0[6] ) );
  BUF_X2 \SB1_4_8/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[139] ), .Z(
        \SB1_4_8/i0[6] ) );
  BUF_X2 \SB1_4_29/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[12] ), .Z(
        \SB1_4_29/i0[9] ) );
  BUF_X2 \SB1_4_5/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[156] ), .Z(
        \SB1_4_5/i0[9] ) );
  BUF_X2 \SB1_4_23/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[51] ), .Z(
        \SB1_4_23/i0[10] ) );
  INV_X2 \SB1_4_29/INV_5  ( .I(\RI1[4][17] ), .ZN(\SB1_4_29/i1_5 ) );
  CLKBUF_X2 \SB1_4_3/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[169] ), .Z(
        \SB1_4_3/i0[6] ) );
  CLKBUF_X2 \SB1_4_2/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[178] ), .Z(
        \SB1_4_2/i0_4 ) );
  BUF_X2 U5191 ( .I(\MC_ARK_ARC_1_3/buf_output[50] ), .Z(\SB1_4_23/i0_0 ) );
  BUF_X2 U962 ( .I(\MC_ARK_ARC_1_3/buf_output[170] ), .Z(\SB1_4_3/i0_0 ) );
  BUF_X2 \SB1_4_1/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[184] ), .Z(
        \SB1_4_1/i0_4 ) );
  INV_X1 \SB1_4_27/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[25] ), .ZN(
        \SB1_4_27/i1_7 ) );
  INV_X1 \SB1_4_2/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[176] ), .ZN(
        \SB1_4_2/i1[9] ) );
  INV_X1 \SB1_4_18/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[81] ), .ZN(
        \SB1_4_18/i0[8] ) );
  INV_X1 \SB1_4_21/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[63] ), .ZN(
        \SB1_4_21/i0[8] ) );
  INV_X1 \SB1_4_11/INV_3  ( .I(n1504), .ZN(\SB1_4_11/i0[8] ) );
  INV_X1 \SB1_4_17/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[86] ), .ZN(
        \SB1_4_17/i1[9] ) );
  NAND3_X1 U3900 ( .A1(\SB1_4_4/i0[8] ), .A2(\SB1_4_4/i3[0] ), .A3(
        \SB1_4_4/i1_5 ), .ZN(n3733) );
  NAND3_X1 U11359 ( .A1(\SB1_4_14/i0[10] ), .A2(\SB1_4_14/i1[9] ), .A3(
        \SB1_4_14/i1_7 ), .ZN(n4688) );
  NAND3_X1 U755 ( .A1(\SB1_4_5/i0[10] ), .A2(\SB1_4_5/i0[6] ), .A3(
        \SB1_4_5/i0_3 ), .ZN(n2078) );
  NAND3_X1 U3894 ( .A1(\SB1_4_1/i0_0 ), .A2(\SB1_4_1/i0_3 ), .A3(
        \SB1_4_1/i0_4 ), .ZN(\SB1_4_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U875 ( .A1(\SB1_4_20/i0[9] ), .A2(\SB1_4_20/i0[10] ), .A3(
        \SB1_4_20/i0_3 ), .ZN(\SB1_4_20/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2993 ( .A1(\SB1_4_15/i0_4 ), .A2(\SB1_4_15/i0_3 ), .A3(
        \SB1_4_15/i1[9] ), .ZN(n5299) );
  NAND3_X1 U911 ( .A1(\SB1_4_2/i3[0] ), .A2(\SB1_4_2/i0[8] ), .A3(
        \SB1_4_2/i1_5 ), .ZN(n3207) );
  NAND3_X1 \SB1_4_30/Component_Function_3/N4  ( .A1(\SB1_4_30/i1_5 ), .A2(
        \SB1_4_30/i0[8] ), .A3(\SB1_4_30/i3[0] ), .ZN(
        \SB1_4_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_1/Component_Function_0/N2  ( .A1(\SB1_4_1/i0[8] ), .A2(
        \SB1_4_1/i0[7] ), .A3(\SB1_4_1/i0[6] ), .ZN(
        \SB1_4_1/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U772 ( .A1(\SB1_4_20/i0[8] ), .A2(\SB1_4_20/i3[0] ), .A3(
        \SB1_4_20/i1_5 ), .ZN(\SB1_4_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_0/Component_Function_4/N2  ( .A1(\SB1_4_0/i3[0] ), .A2(
        \SB1_4_0/i0_0 ), .A3(\SB1_4_0/i1_7 ), .ZN(
        \SB1_4_0/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 \SB1_4_3/Component_Function_5/N1  ( .A1(\SB1_4_3/i0_0 ), .A2(
        \SB1_4_3/i3[0] ), .ZN(\SB1_4_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U8880 ( .A1(\SB1_4_17/i0[6] ), .A2(\SB1_4_17/i0_3 ), .A3(
        \SB1_4_17/i1[9] ), .ZN(n5373) );
  NAND3_X1 U765 ( .A1(\SB1_4_6/i0[8] ), .A2(\SB1_4_6/i1_7 ), .A3(
        \SB1_4_6/i0_4 ), .ZN(n3153) );
  NAND3_X1 U2812 ( .A1(\SB1_4_18/i0[10] ), .A2(\SB1_4_18/i1[9] ), .A3(
        \SB1_4_18/i1_5 ), .ZN(\SB1_4_18/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_0/Component_Function_1/N1  ( .A1(\SB1_4_0/i0_3 ), .A2(
        \SB1_4_0/i1[9] ), .ZN(\SB1_4_0/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_2/Component_Function_5/N1  ( .A1(\SB1_4_2/i0_0 ), .A2(
        \SB1_4_2/i3[0] ), .ZN(\SB1_4_2/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U3926 ( .I(\MC_ARK_ARC_1_3/buf_output[120] ), .ZN(\SB1_4_11/i3[0] )
         );
  NAND3_X1 \SB1_4_10/Component_Function_2/N3  ( .A1(\RI1[4][131] ), .A2(
        \SB1_4_10/i0[8] ), .A3(\SB1_4_10/i0[9] ), .ZN(
        \SB1_4_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U869 ( .A1(\SB1_4_30/i0[10] ), .A2(\SB1_4_30/i1_7 ), .A3(
        \SB1_4_30/i1[9] ), .ZN(n4125) );
  NAND3_X1 U6098 ( .A1(\SB1_4_11/i0[9] ), .A2(\SB1_4_11/i0[6] ), .A3(
        \SB1_4_11/i1_5 ), .ZN(n1778) );
  NAND3_X1 U4205 ( .A1(\SB1_4_2/i0[9] ), .A2(\SB1_4_2/i0[8] ), .A3(
        \SB1_4_2/i0_3 ), .ZN(n1115) );
  INV_X1 \SB1_4_22/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[54] ), .ZN(
        \SB1_4_22/i3[0] ) );
  NAND3_X1 U4284 ( .A1(\SB1_4_9/i0_3 ), .A2(\SB1_4_9/i1[9] ), .A3(
        \SB1_4_9/i0[6] ), .ZN(n1228) );
  NAND3_X1 \SB1_4_9/Component_Function_2/N3  ( .A1(\SB1_4_9/i0_3 ), .A2(
        \SB1_4_9/i0[8] ), .A3(\SB1_4_9/i0[9] ), .ZN(
        \SB1_4_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_1/Component_Function_2/N2  ( .A1(\SB1_4_1/i0_3 ), .A2(
        \SB1_4_1/i0[10] ), .A3(\SB1_4_1/i0[6] ), .ZN(
        \SB1_4_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U10070 ( .A1(\SB1_4_30/i0[6] ), .A2(\SB1_4_30/i0[10] ), .A3(
        \SB1_4_30/i0_0 ), .ZN(\SB1_4_30/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U10847 ( .A1(\SB1_4_29/i0[9] ), .A2(\SB1_4_29/i0[6] ), .A3(
        \SB1_4_29/i0_4 ), .ZN(n4451) );
  NAND3_X1 U2992 ( .A1(\SB1_4_17/i0[10] ), .A2(\SB1_4_17/i0_0 ), .A3(
        \SB1_4_17/i0[6] ), .ZN(\SB1_4_17/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_4/Component_Function_4/N3  ( .A1(\SB1_4_4/i0[9] ), .A2(
        \SB1_4_4/i0[10] ), .A3(\SB1_4_4/i0_3 ), .ZN(
        \SB1_4_4/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB1_4_29/Component_Function_0/N1  ( .A1(\SB1_4_29/i0[10] ), .A2(
        \SB1_4_29/i0[9] ), .ZN(\SB1_4_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_4_20/Component_Function_3/N2  ( .A1(\SB1_4_20/i0_0 ), .A2(
        \SB1_4_20/i0_3 ), .A3(\SB1_4_20/i0_4 ), .ZN(
        \SB1_4_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U879 ( .A1(\SB1_4_0/i0[6] ), .A2(\SB1_4_0/i1[9] ), .A3(
        \RI1[4][191] ), .ZN(n4462) );
  NAND2_X1 U12159 ( .A1(n5117), .A2(\SB1_4_25/i0_0 ), .ZN(
        \SB1_4_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_22/Component_Function_1/N3  ( .A1(\SB1_4_22/i1_5 ), .A2(
        \SB1_4_22/i0[6] ), .A3(\SB1_4_22/i0[9] ), .ZN(
        \SB1_4_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3941 ( .A1(\SB1_4_10/i0[8] ), .A2(\SB1_4_10/i1_7 ), .A3(
        \SB1_4_10/i0_4 ), .ZN(\SB1_4_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U757 ( .A1(\SB1_4_26/i0_0 ), .A2(\SB1_4_26/i1_5 ), .A3(
        \SB1_4_26/i0_4 ), .ZN(n1261) );
  NAND3_X1 U9635 ( .A1(\RI1[4][191] ), .A2(\SB1_4_0/i0[6] ), .A3(
        \SB1_4_0/i0[10] ), .ZN(\SB1_4_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_7/Component_Function_0/N3  ( .A1(\SB1_4_7/i0[10] ), .A2(
        \SB1_4_7/i0_4 ), .A3(\SB1_4_7/i0_3 ), .ZN(
        \SB1_4_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U7759 ( .A1(\SB1_4_2/i0[9] ), .A2(\SB1_4_2/i0[10] ), .A3(
        \SB1_4_2/i0_3 ), .ZN(n4423) );
  NAND3_X1 U717 ( .A1(\SB1_4_0/i0[9] ), .A2(\SB1_4_0/i0[6] ), .A3(
        \SB1_4_0/i1_5 ), .ZN(\SB1_4_0/Component_Function_1/NAND4_in[2] ) );
  INV_X1 \SB1_4_27/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[24] ), .ZN(
        \SB1_4_27/i3[0] ) );
  NAND3_X1 U5032 ( .A1(\SB1_4_16/i3[0] ), .A2(\SB1_4_16/i0_0 ), .A3(
        \SB1_4_16/i1_7 ), .ZN(\SB1_4_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_4_17/Component_Function_1/N2  ( .A1(\SB1_4_17/i0_3 ), .A2(
        \SB1_4_17/i1_7 ), .A3(\SB1_4_17/i0[8] ), .ZN(
        \SB1_4_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U12102 ( .A1(\SB1_4_15/i0[6] ), .A2(\SB1_4_15/i1[9] ), .A3(
        \SB1_4_15/i0_3 ), .ZN(n5086) );
  NAND3_X1 U8324 ( .A1(\SB1_4_2/i0[9] ), .A2(\SB1_4_2/i0_0 ), .A3(
        \SB1_4_2/i0[8] ), .ZN(n3805) );
  NAND3_X1 U9673 ( .A1(\SB1_4_14/i0_4 ), .A2(\SB1_4_14/i0_0 ), .A3(
        \SB1_4_14/i0_3 ), .ZN(n2839) );
  NAND3_X1 \SB1_4_23/Component_Function_4/N1  ( .A1(\SB1_4_23/i0[9] ), .A2(
        \SB1_4_23/i0_0 ), .A3(\SB1_4_23/i0[8] ), .ZN(
        \SB1_4_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U3943 ( .A1(\SB1_4_14/i0[9] ), .A2(\SB1_4_14/i0_3 ), .A3(
        \SB1_4_14/i0[8] ), .ZN(\SB1_4_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_4_28/Component_Function_3/N3  ( .A1(\SB1_4_28/i1[9] ), .A2(
        \SB1_4_28/i1_7 ), .A3(\SB1_4_28/i0[10] ), .ZN(
        \SB1_4_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3393 ( .A1(\SB1_4_26/i0[9] ), .A2(\SB1_4_26/i1_5 ), .A3(
        \SB1_4_26/i0[6] ), .ZN(\SB1_4_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U9606 ( .A1(\SB1_4_24/i1_7 ), .A2(\SB1_4_24/i0[8] ), .A3(
        \SB1_4_24/i0_4 ), .ZN(\SB1_4_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U12149 ( .A1(\SB1_4_20/i0_3 ), .A2(\SB1_4_20/i0_4 ), .A3(
        \SB1_4_20/i1[9] ), .ZN(n5111) );
  NAND3_X1 U9581 ( .A1(\SB1_4_20/i0[7] ), .A2(\SB1_4_20/i0_3 ), .A3(
        \SB1_4_20/i0_0 ), .ZN(\SB1_4_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3933 ( .A1(\SB1_4_25/i0_3 ), .A2(\SB1_4_25/i0_0 ), .A3(
        \SB1_4_25/i0[7] ), .ZN(n1902) );
  NAND3_X1 U778 ( .A1(\SB1_4_29/i0_4 ), .A2(\SB1_4_29/i1_7 ), .A3(
        \SB1_4_29/i0[8] ), .ZN(\SB1_4_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_11/Component_Function_3/N3  ( .A1(\SB1_4_11/i1[9] ), .A2(
        \SB1_4_11/i1_7 ), .A3(\SB1_4_11/i0[10] ), .ZN(
        \SB1_4_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U9849 ( .A1(\SB1_4_19/i0[6] ), .A2(\SB1_4_19/i0[9] ), .A3(
        \SB1_4_19/i1_5 ), .ZN(\SB1_4_19/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U12572 ( .A1(\SB1_4_11/i0_0 ), .A2(\SB1_4_11/i3[0] ), .ZN(
        \SB1_4_11/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_4/Component_Function_5/N1  ( .A1(\SB1_4_4/i0_0 ), .A2(
        \SB1_4_4/i3[0] ), .ZN(\SB1_4_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U6277 ( .A1(\SB1_4_25/i0[6] ), .A2(\SB1_4_25/i0[8] ), .A3(
        \SB1_4_25/i0[7] ), .ZN(n3522) );
  NAND3_X1 U2733 ( .A1(\SB1_4_18/i0[9] ), .A2(\SB1_4_18/i1_5 ), .A3(
        \SB1_4_18/i0[6] ), .ZN(\SB1_4_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U9208 ( .A1(\SB1_4_7/i1[9] ), .A2(\SB1_4_7/i0[10] ), .A3(
        \SB1_4_7/i1_5 ), .ZN(n4062) );
  NAND3_X1 U1522 ( .A1(\SB1_4_8/i0[9] ), .A2(\SB1_4_8/i0_4 ), .A3(
        \SB1_4_8/i0[6] ), .ZN(\SB1_4_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U812 ( .A1(\SB1_4_30/i0[6] ), .A2(\SB1_4_30/i0_3 ), .A3(
        \SB1_4_30/i0[10] ), .ZN(n3562) );
  NAND2_X1 \SB1_4_10/Component_Function_5/N1  ( .A1(\SB1_4_10/i0_0 ), .A2(
        \SB1_4_10/i3[0] ), .ZN(\SB1_4_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U855 ( .A1(\SB1_4_5/i0[10] ), .A2(\SB1_4_5/i0[9] ), .A3(
        \SB1_4_5/i0_3 ), .ZN(n4328) );
  NAND3_X1 \SB1_4_29/Component_Function_2/N4  ( .A1(\SB1_4_29/i1_5 ), .A2(
        \SB1_4_29/i0_0 ), .A3(\SB1_4_29/i0_4 ), .ZN(
        \SB1_4_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_4_9/Component_Function_1/N3  ( .A1(\SB1_4_9/i1_5 ), .A2(
        \SB1_4_9/i0[6] ), .A3(\SB1_4_9/i0[9] ), .ZN(
        \SB1_4_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U12579 ( .A1(\SB1_4_6/i0[6] ), .A2(\SB1_4_6/i1[9] ), .A3(
        \RI1[4][155] ), .ZN(\SB1_4_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U728 ( .A1(\SB1_4_21/i0[6] ), .A2(\SB1_4_21/i0[9] ), .A3(
        \SB1_4_21/i0_4 ), .ZN(n2463) );
  NAND3_X1 U3927 ( .A1(\SB1_4_17/i0_0 ), .A2(\SB1_4_17/i1_5 ), .A3(
        \SB1_4_17/i0_4 ), .ZN(n4548) );
  NAND3_X1 U795 ( .A1(\SB1_4_12/i0[10] ), .A2(\RI1[4][119] ), .A3(
        \SB1_4_12/i0[6] ), .ZN(\SB1_4_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U712 ( .A1(\SB1_4_31/i0[9] ), .A2(\SB1_4_31/i0[6] ), .A3(
        \SB1_4_31/i1_5 ), .ZN(n1610) );
  NAND3_X1 \SB1_4_25/Component_Function_1/N4  ( .A1(\SB1_4_25/i1_7 ), .A2(
        \SB1_4_25/i0[8] ), .A3(\SB1_4_25/i0_4 ), .ZN(
        \SB1_4_25/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_4_31/Component_Function_0/N1  ( .A1(\SB1_4_31/i0[10] ), .A2(
        \SB1_4_31/i0[9] ), .ZN(\SB1_4_31/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_4_14/Component_Function_0/N1  ( .A1(\SB1_4_14/i0[10] ), .A2(
        \SB1_4_14/i0[9] ), .ZN(\SB1_4_14/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U6957 ( .A1(n3805), .A2(n4423), .ZN(n3621) );
  NAND3_X1 U787 ( .A1(\SB1_4_28/i0_3 ), .A2(\SB1_4_28/i1[9] ), .A3(
        \SB1_4_28/i0_4 ), .ZN(\SB1_4_28/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2576 ( .A1(\SB1_4_28/i0_3 ), .A2(\SB1_4_28/i0[9] ), .A3(
        \SB1_4_28/i0[10] ), .ZN(\SB1_4_28/Component_Function_4/NAND4_in[2] )
         );
  NAND2_X1 \SB1_4_1/Component_Function_5/N1  ( .A1(\SB1_4_1/i0_0 ), .A2(
        \SB1_4_1/i3[0] ), .ZN(\SB1_4_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U713 ( .A1(\SB1_4_26/i0_4 ), .A2(\SB1_4_26/i0[9] ), .A3(
        \SB1_4_26/i0[6] ), .ZN(n2199) );
  BUF_X4 U1978 ( .I(\SB1_4_24/buf_output[5] ), .Z(\SB2_4_24/i0_3 ) );
  CLKBUF_X2 \SB2_4_31/BUF_0  ( .I(\SB1_4_4/buf_output[0] ), .Z(
        \SB2_4_31/i0[9] ) );
  BUF_X2 U5382 ( .I(\SB1_4_2/buf_output[0] ), .Z(\SB2_4_29/i0[9] ) );
  INV_X1 U6099 ( .I(\SB1_4_10/buf_output[1] ), .ZN(\SB2_4_6/i1_7 ) );
  CLKBUF_X2 \SB2_4_0/BUF_0  ( .I(\SB1_4_5/buf_output[0] ), .Z(\SB2_4_0/i0[9] )
         );
  CLKBUF_X2 \SB2_4_2/BUF_2  ( .I(\SB1_4_5/buf_output[2] ), .Z(\SB2_4_2/i0_0 )
         );
  BUF_X2 \SB2_4_28/BUF_0  ( .I(\SB1_4_1/buf_output[0] ), .Z(\SB2_4_28/i0[9] )
         );
  BUF_X2 U3201 ( .I(\SB1_4_24/buf_output[0] ), .Z(\SB2_4_19/i0[9] ) );
  BUF_X2 \SB2_4_29/BUF_4  ( .I(\SB1_4_30/buf_output[4] ), .Z(\SB2_4_29/i0_4 )
         );
  INV_X1 \SB2_4_6/INV_2  ( .I(\SB1_4_9/buf_output[2] ), .ZN(\SB2_4_6/i1[9] )
         );
  INV_X1 U4882 ( .I(\SB1_4_26/buf_output[2] ), .ZN(\SB2_4_23/i1[9] ) );
  NAND2_X1 U2900 ( .A1(\SB2_4_30/i0_0 ), .A2(n3983), .ZN(
        \SB2_4_30/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_3/Component_Function_5/N1  ( .A1(\SB2_4_3/i0_0 ), .A2(
        \SB2_4_3/i3[0] ), .ZN(\SB2_4_3/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_23/Component_Function_5/N1  ( .A1(\SB2_4_23/i0_0 ), .A2(
        \SB2_4_23/i3[0] ), .ZN(\SB2_4_23/Component_Function_5/NAND4_in[0] ) );
  INV_X1 \SB2_4_25/INV_1  ( .I(\SB1_4_29/buf_output[1] ), .ZN(\SB2_4_25/i1_7 )
         );
  INV_X1 \SB2_4_11/INV_0  ( .I(\SB1_4_16/buf_output[0] ), .ZN(\SB2_4_11/i3[0] ) );
  INV_X1 \SB2_4_26/INV_0  ( .I(\SB1_4_31/buf_output[0] ), .ZN(\SB2_4_26/i3[0] ) );
  INV_X1 \SB2_4_20/INV_1  ( .I(\SB1_4_24/buf_output[1] ), .ZN(\SB2_4_20/i1_7 )
         );
  INV_X1 \SB2_4_7/INV_1  ( .I(\SB1_4_11/buf_output[1] ), .ZN(\SB2_4_7/i1_7 )
         );
  INV_X2 U5367 ( .I(\SB2_4_31/i0_4 ), .ZN(\SB2_4_31/i0[7] ) );
  INV_X1 \SB2_4_19/INV_1  ( .I(\SB1_4_23/buf_output[1] ), .ZN(\SB2_4_19/i1_7 )
         );
  INV_X1 U1829 ( .I(\SB1_4_6/buf_output[1] ), .ZN(\SB2_4_2/i1_7 ) );
  NAND3_X1 U7944 ( .A1(\SB2_4_31/i0[10] ), .A2(\SB2_4_31/i0_0 ), .A3(
        \SB2_4_31/i0[6] ), .ZN(\SB2_4_31/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X2 U5154 ( .I(\SB1_4_13/buf_output[0] ), .Z(\SB2_4_8/i0[9] ) );
  CLKBUF_X2 U9688 ( .I(\SB1_4_28/buf_output[2] ), .Z(\SB2_4_25/i0_0 ) );
  BUF_X2 U1727 ( .I(\SB1_4_6/buf_output[0] ), .Z(\SB2_4_1/i0[9] ) );
  BUF_X2 \SB2_4_8/BUF_2  ( .I(\SB1_4_11/buf_output[2] ), .Z(\SB2_4_8/i0_0 ) );
  CLKBUF_X2 \SB2_4_5/BUF_1  ( .I(\SB1_4_9/buf_output[1] ), .Z(\SB2_4_5/i0[6] )
         );
  CLKBUF_X2 U3405 ( .I(\SB1_4_15/buf_output[1] ), .Z(\SB2_4_11/i0[6] ) );
  BUF_X2 \SB2_4_25/BUF_1  ( .I(\SB1_4_29/buf_output[1] ), .Z(\SB2_4_25/i0[6] )
         );
  INV_X1 U2974 ( .I(\SB1_4_18/buf_output[1] ), .ZN(\SB2_4_14/i1_7 ) );
  INV_X1 U7315 ( .I(\SB1_4_23/buf_output[5] ), .ZN(\SB2_4_23/i1_5 ) );
  AND4_X1 U9615 ( .A1(\SB1_4_0/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_4_0/Component_Function_5/NAND4_in[2] ), .A3(n830), .A4(n4459), 
        .Z(n3978) );
  INV_X1 \SB2_4_28/INV_5  ( .I(\SB1_4_28/buf_output[5] ), .ZN(\SB2_4_28/i1_5 )
         );
  NAND3_X1 \SB2_4_7/Component_Function_2/N1  ( .A1(\SB2_4_7/i1_5 ), .A2(
        \SB2_4_7/i0[10] ), .A3(\SB2_4_7/i1[9] ), .ZN(
        \SB2_4_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_21/Component_Function_0/N2  ( .A1(\SB2_4_21/i0[8] ), .A2(
        \SB2_4_21/i0[7] ), .A3(\SB2_4_21/i0[6] ), .ZN(
        \SB2_4_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_26/Component_Function_2/N1  ( .A1(\SB2_4_26/i1_5 ), .A2(
        \SB2_4_26/i0[10] ), .A3(\SB2_4_26/i1[9] ), .ZN(
        \SB2_4_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U6136 ( .A1(\SB2_4_24/i0[10] ), .A2(\SB2_4_24/i0_3 ), .A3(
        \SB2_4_24/i0[9] ), .ZN(n3513) );
  NAND3_X1 \SB2_4_8/Component_Function_2/N2  ( .A1(\SB2_4_8/i0_3 ), .A2(
        \SB2_4_8/i0[10] ), .A3(\SB2_4_8/i0[6] ), .ZN(
        \SB2_4_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_31/Component_Function_3/N1  ( .A1(\SB2_4_31/i1[9] ), .A2(
        \SB2_4_31/i0_3 ), .A3(\SB2_4_31/i0[6] ), .ZN(
        \SB2_4_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4368 ( .A1(\SB2_4_5/i1_7 ), .A2(\SB1_4_6/buf_output[4] ), .A3(
        \SB2_4_5/i0[8] ), .ZN(\SB2_4_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U6302 ( .A1(\SB2_4_16/i0_0 ), .A2(\SB2_4_16/i0_3 ), .A3(
        \SB2_4_16/i0[7] ), .ZN(n3527) );
  NAND3_X1 U10807 ( .A1(\SB2_4_0/i0_3 ), .A2(\SB2_4_0/i0[10] ), .A3(
        \SB2_4_0/i0[9] ), .ZN(n5051) );
  NAND3_X1 \SB2_4_2/Component_Function_3/N1  ( .A1(\SB2_4_2/i1[9] ), .A2(
        \SB2_4_2/i0_3 ), .A3(\SB2_4_2/i0[6] ), .ZN(
        \SB2_4_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U669 ( .A1(\SB2_4_4/i0_3 ), .A2(\SB2_4_4/i1[9] ), .A3(
        \SB2_4_4/i0[6] ), .ZN(\SB2_4_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_12/Component_Function_0/N3  ( .A1(\SB2_4_12/i0[10] ), .A2(
        \SB2_4_12/i0_4 ), .A3(\SB2_4_12/i0_3 ), .ZN(
        \SB2_4_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U6204 ( .A1(\SB2_4_6/i0_3 ), .A2(\SB2_4_6/i0_0 ), .A3(
        \SB2_4_6/i0[7] ), .ZN(n1823) );
  NAND3_X1 U2598 ( .A1(\SB2_4_29/i0_0 ), .A2(\SB2_4_29/i0_3 ), .A3(
        \SB2_4_29/i0[7] ), .ZN(n795) );
  NAND3_X1 \SB2_4_30/Component_Function_0/N4  ( .A1(n6265), .A2(
        \SB2_4_30/i0_3 ), .A3(\SB2_4_30/i0_0 ), .ZN(
        \SB2_4_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2853 ( .A1(n6269), .A2(\SB2_4_10/i0_0 ), .A3(\SB2_4_10/i0_4 ), 
        .ZN(\SB2_4_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_1/Component_Function_0/N3  ( .A1(\SB2_4_1/i0[10] ), .A2(
        \SB2_4_1/i0_4 ), .A3(\SB2_4_1/i0_3 ), .ZN(
        \SB2_4_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_4_14/Component_Function_4/N2  ( .A1(\SB2_4_14/i3[0] ), .A2(
        \SB2_4_14/i0_0 ), .A3(\SB2_4_14/i1_7 ), .ZN(
        \SB2_4_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_6/Component_Function_3/N4  ( .A1(\SB2_4_6/i1_5 ), .A2(
        \SB2_4_6/i0[8] ), .A3(\SB2_4_6/i3[0] ), .ZN(
        \SB2_4_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_3/Component_Function_4/N4  ( .A1(\SB2_4_3/i1[9] ), .A2(n3988), .A3(\SB2_4_3/i0_4 ), .ZN(\SB2_4_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U739 ( .A1(\SB2_4_12/i3[0] ), .A2(\SB2_4_12/i1_5 ), .A3(
        \SB2_4_12/i0[8] ), .ZN(n5127) );
  NAND3_X1 U746 ( .A1(\SB2_4_3/i0_3 ), .A2(\SB2_4_3/i0[10] ), .A3(
        \SB2_4_3/i0[9] ), .ZN(\SB2_4_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U9713 ( .A1(\SB2_4_28/i1_7 ), .A2(n4000), .A3(\SB2_4_28/i0_4 ), 
        .ZN(\SB2_4_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_21/Component_Function_3/N4  ( .A1(\SB2_4_21/i1_5 ), .A2(
        \SB2_4_21/i0[8] ), .A3(\SB2_4_21/i3[0] ), .ZN(
        \SB2_4_21/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 U6829 ( .A1(\SB2_4_25/i0_0 ), .A2(\SB2_4_25/i3[0] ), .ZN(n2116) );
  NAND3_X1 U1532 ( .A1(\SB2_4_28/i0_3 ), .A2(n4000), .A3(\SB2_4_28/i0[9] ), 
        .ZN(\SB2_4_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3974 ( .A1(\SB2_4_22/i0[7] ), .A2(\SB2_4_22/i0_3 ), .A3(
        \SB2_4_22/i0_0 ), .ZN(\SB2_4_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_29/Component_Function_1/N2  ( .A1(\SB2_4_29/i0_3 ), .A2(
        \SB2_4_29/i1_7 ), .A3(\SB2_4_29/i0[8] ), .ZN(
        \SB2_4_29/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2947 ( .A1(\SB2_4_25/i0_0 ), .A2(\SB2_4_25/i1_5 ), .A3(
        \SB2_4_25/i0_4 ), .ZN(n746) );
  NAND3_X1 U677 ( .A1(\SB2_4_23/i0_0 ), .A2(\SB2_4_23/i0[9] ), .A3(
        \SB2_4_23/i0[8] ), .ZN(n4918) );
  NAND2_X1 \SB2_4_5/Component_Function_5/N1  ( .A1(\SB2_4_5/i0_0 ), .A2(
        \SB2_4_5/i3[0] ), .ZN(\SB2_4_5/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_21/Component_Function_5/N1  ( .A1(\SB2_4_21/i0_0 ), .A2(
        \SB2_4_21/i3[0] ), .ZN(\SB2_4_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_15/Component_Function_5/N4  ( .A1(\SB2_4_15/i0[9] ), .A2(
        \SB2_4_15/i0[6] ), .A3(\SB2_4_15/i0_4 ), .ZN(
        \SB2_4_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2400 ( .A1(\SB2_4_13/i0_4 ), .A2(\SB2_4_13/i1_7 ), .A3(
        \SB2_4_13/i0[8] ), .ZN(n639) );
  NAND3_X1 \SB2_4_14/Component_Function_2/N1  ( .A1(\SB2_4_14/i1_5 ), .A2(
        \SB2_4_14/i0[10] ), .A3(\SB2_4_14/i1[9] ), .ZN(
        \SB2_4_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U10888 ( .A1(\SB2_4_9/i0[6] ), .A2(\SB2_4_9/i1_5 ), .A3(
        \SB2_4_9/i0[9] ), .ZN(n4670) );
  NAND3_X1 U653 ( .A1(\SB2_4_10/i0[8] ), .A2(\SB2_4_10/i3[0] ), .A3(n6269), 
        .ZN(n2731) );
  NAND3_X1 \SB2_4_21/Component_Function_4/N4  ( .A1(\SB2_4_21/i1[9] ), .A2(
        \SB2_4_21/i1_5 ), .A3(\SB2_4_21/i0_4 ), .ZN(
        \SB2_4_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_1/Component_Function_0/N4  ( .A1(n3370), .A2(\SB2_4_1/i0_3 ), 
        .A3(\SB2_4_1/i0_0 ), .ZN(\SB2_4_1/Component_Function_0/NAND4_in[3] )
         );
  NAND3_X1 \SB2_4_3/Component_Function_2/N3  ( .A1(\SB2_4_3/i0_3 ), .A2(
        \SB2_4_3/i0[8] ), .A3(\SB2_4_3/i0[9] ), .ZN(
        \SB2_4_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3965 ( .A1(\SB2_4_21/i0_3 ), .A2(\SB2_4_21/i0[8] ), .A3(
        \SB2_4_21/i0[9] ), .ZN(\SB2_4_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U7685 ( .A1(\SB2_4_16/i0[6] ), .A2(\SB2_4_16/i1_5 ), .A3(
        \SB2_4_16/i0[9] ), .ZN(\SB2_4_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U5935 ( .A1(\SB2_4_7/i0[10] ), .A2(\SB2_4_7/i0_3 ), .A3(
        \SB2_4_7/i0[6] ), .ZN(n1712) );
  NAND3_X1 \SB2_4_17/Component_Function_2/N2  ( .A1(\SB2_4_17/i0_3 ), .A2(
        \SB2_4_17/i0[10] ), .A3(\SB2_4_17/i0[6] ), .ZN(
        \SB2_4_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_4_23/Component_Function_3/N2  ( .A1(\SB2_4_23/i0_0 ), .A2(
        \SB2_4_23/i0_3 ), .A3(\SB2_4_23/i0_4 ), .ZN(
        \SB2_4_23/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 \SB2_4_15/Component_Function_0/N1  ( .A1(\SB2_4_15/i0[10] ), .A2(
        \SB2_4_15/i0[9] ), .ZN(\SB2_4_15/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_4_26/Component_Function_0/N1  ( .A1(\SB2_4_26/i0[10] ), .A2(
        \SB2_4_26/i0[9] ), .ZN(\SB2_4_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U11967 ( .A1(\SB2_4_20/i0[9] ), .A2(\SB2_4_20/i0_4 ), .A3(
        \SB2_4_20/i0[6] ), .ZN(n5024) );
  NAND3_X1 U2784 ( .A1(\SB2_4_11/i0[9] ), .A2(\SB2_4_11/i0[10] ), .A3(
        \SB2_4_11/i0_3 ), .ZN(\SB2_4_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3980 ( .A1(\SB2_4_14/i1_5 ), .A2(\SB2_4_14/i0_0 ), .A3(
        \SB2_4_14/i0_4 ), .ZN(\SB2_4_14/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_4/Component_Function_4/N4  ( .A1(\SB2_4_4/i1[9] ), .A2(
        \SB2_4_4/i1_5 ), .A3(\SB2_4_4/i0_4 ), .ZN(
        \SB2_4_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_21/Component_Function_3/N2  ( .A1(\SB2_4_21/i0_0 ), .A2(
        \SB2_4_21/i0_3 ), .A3(\SB2_4_21/i0_4 ), .ZN(
        \SB2_4_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4382 ( .A1(\SB2_4_25/i0[9] ), .A2(\SB2_4_25/i0[6] ), .A3(
        \SB2_4_25/i0_4 ), .ZN(n3216) );
  NAND3_X1 \SB2_4_16/Component_Function_1/N4  ( .A1(\SB2_4_16/i1_7 ), .A2(
        \SB2_4_16/i0[8] ), .A3(\SB2_4_16/i0_4 ), .ZN(
        \SB2_4_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_4_12/Component_Function_4/N4  ( .A1(\SB2_4_12/i1[9] ), .A2(
        \SB2_4_12/i1_5 ), .A3(\SB2_4_12/i0_4 ), .ZN(
        \SB2_4_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U738 ( .A1(\SB2_4_0/i0[10] ), .A2(\SB2_4_0/i1_7 ), .A3(
        \SB2_4_0/i1[9] ), .ZN(n4145) );
  NAND3_X1 \SB2_4_16/Component_Function_1/N2  ( .A1(\SB2_4_16/i0_3 ), .A2(
        \SB2_4_16/i1_7 ), .A3(\SB2_4_16/i0[8] ), .ZN(
        \SB2_4_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1815 ( .A1(\SB2_4_25/i0_3 ), .A2(\SB2_4_25/i0[6] ), .A3(
        \SB2_4_25/i1[9] ), .ZN(\SB2_4_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_3/Component_Function_1/N4  ( .A1(\SB2_4_3/i1_7 ), .A2(
        \SB2_4_3/i0[8] ), .A3(\SB2_4_3/i0_4 ), .ZN(
        \SB2_4_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U9549 ( .A1(\SB2_4_14/i0_3 ), .A2(\SB2_4_14/i1[9] ), .A3(
        \SB2_4_14/i0_4 ), .ZN(n2993) );
  NAND3_X1 U9589 ( .A1(\SB2_4_6/i0_3 ), .A2(\SB2_4_6/i0[10] ), .A3(
        \SB2_4_6/i0[6] ), .ZN(\SB2_4_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U7473 ( .A1(\SB2_4_16/i0[6] ), .A2(\SB2_4_16/i0_4 ), .A3(
        \SB2_4_16/i0[9] ), .ZN(n2410) );
  NAND3_X1 \SB2_4_19/Component_Function_2/N2  ( .A1(\SB2_4_19/i0_3 ), .A2(
        \SB2_4_19/i0[10] ), .A3(\SB2_4_19/i0[6] ), .ZN(
        \SB2_4_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U716 ( .A1(\SB2_4_10/i0[9] ), .A2(\SB2_4_10/i0_4 ), .A3(
        \SB2_4_10/i0[6] ), .ZN(n1043) );
  NAND3_X1 \SB2_4_12/Component_Function_2/N3  ( .A1(\SB2_4_12/i0_3 ), .A2(
        \SB2_4_12/i0[8] ), .A3(\SB2_4_12/i0[9] ), .ZN(
        \SB2_4_12/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 \SB2_4_26/Component_Function_1/N1  ( .A1(\SB2_4_26/i0_3 ), .A2(
        \SB2_4_26/i1[9] ), .ZN(\SB2_4_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_4_2/Component_Function_2/N2  ( .A1(\SB2_4_2/i0_3 ), .A2(
        \SB2_4_2/i0[10] ), .A3(\SB2_4_2/i0[6] ), .ZN(
        \SB2_4_2/Component_Function_2/NAND4_in[1] ) );
  NAND4_X1 U2629 ( .A1(\SB2_4_13/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_4_13/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_4_13/Component_Function_1/NAND4_in[0] ), .A4(n639), .ZN(
        \SB2_4_13/buf_output[1] ) );
  BUF_X2 U8560 ( .I(\SB2_4_19/buf_output[0] ), .Z(\RI5[4][102] ) );
  INV_X1 \SB3_28/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[18] ), .ZN(
        \SB3_28/i3[0] ) );
  BUF_X2 \SB3_27/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[24] ), .Z(
        \SB3_27/i0[9] ) );
  BUF_X2 U9421 ( .I(n3971), .Z(\SB3_24/i0_3 ) );
  INV_X1 \SB3_28/INV_5  ( .I(\MC_ARK_ARC_1_4/buf_output[23] ), .ZN(
        \SB3_28/i1_5 ) );
  NAND2_X1 \SB3_6/Component_Function_5/N1  ( .A1(\SB3_6/i0_0 ), .A2(
        \SB3_6/i3[0] ), .ZN(\SB3_6/Component_Function_5/NAND4_in[0] ) );
  INV_X1 \SB3_16/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[90] ), .ZN(
        \SB3_16/i3[0] ) );
  BUF_X2 U638 ( .I(\MC_ARK_ARC_1_4/buf_output[97] ), .Z(\SB3_15/i0[6] ) );
  INV_X1 U2391 ( .I(\MC_ARK_ARC_1_4/buf_output[131] ), .ZN(\SB3_10/i1_5 ) );
  INV_X1 \SB3_19/INV_0  ( .I(\MC_ARK_ARC_1_4/buf_output[72] ), .ZN(
        \SB3_19/i3[0] ) );
  INV_X1 U5144 ( .I(\MC_ARK_ARC_1_4/buf_output[186] ), .ZN(\SB3_0/i3[0] ) );
  INV_X1 U5200 ( .I(\RI1[5][137] ), .ZN(\SB3_9/i1_5 ) );
  BUF_X2 U8225 ( .I(\MC_ARK_ARC_1_4/buf_output[19] ), .Z(\SB3_28/i0[6] ) );
  BUF_X2 U661 ( .I(\MC_ARK_ARC_1_4/buf_output[124] ), .Z(\SB3_11/i0_4 ) );
  BUF_X2 \SB3_25/BUF_0  ( .I(\MC_ARK_ARC_1_4/buf_output[36] ), .Z(
        \SB3_25/i0[9] ) );
  CLKBUF_X2 U624 ( .I(\MC_ARK_ARC_1_4/buf_output[148] ), .Z(\SB3_7/i0_4 ) );
  INV_X1 \SB3_22/INV_5  ( .I(\RI1[5][59] ), .ZN(\SB3_22/i1_5 ) );
  CLKBUF_X2 U5008 ( .I(\MC_ARK_ARC_1_4/buf_output[175] ), .Z(\SB3_2/i0[6] ) );
  NAND3_X1 U2454 ( .A1(\SB3_4/i0_3 ), .A2(\SB3_4/i1[9] ), .A3(\SB3_4/i0_4 ), 
        .ZN(n3118) );
  NAND3_X1 U9373 ( .A1(\SB3_4/i0[9] ), .A2(\SB3_4/i0[6] ), .A3(\SB3_4/i0_4 ), 
        .ZN(\SB3_4/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U648 ( .A1(\SB3_5/i3[0] ), .A2(\SB3_5/i0[8] ), .A3(\SB3_5/i1_5 ), 
        .ZN(n3598) );
  NAND3_X1 \SB3_25/Component_Function_0/N2  ( .A1(\SB3_25/i0[8] ), .A2(
        \SB3_25/i0[7] ), .A3(\SB3_25/i0[6] ), .ZN(
        \SB3_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB3_2/Component_Function_0/N2  ( .A1(\SB3_2/i0[8] ), .A2(
        \SB3_2/i0[7] ), .A3(\SB3_2/i0[6] ), .ZN(
        \SB3_2/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_19/Component_Function_5/N1  ( .A1(\SB3_19/i0_0 ), .A2(
        \SB3_19/i3[0] ), .ZN(\SB3_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_6/Component_Function_0/N4  ( .A1(\SB3_6/i0[7] ), .A2(
        \SB3_6/i0_3 ), .A3(\SB3_6/i0_0 ), .ZN(
        \SB3_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U9103 ( .A1(\SB3_20/i0_4 ), .A2(\SB3_20/i1_7 ), .A3(\SB3_20/i0[8] ), 
        .ZN(n3916) );
  NAND3_X1 U617 ( .A1(\SB3_2/i0[10] ), .A2(\SB3_2/i1[9] ), .A3(\SB3_2/i1_7 ), 
        .ZN(n1080) );
  NAND3_X1 U2589 ( .A1(\SB3_6/i0_3 ), .A2(\SB3_6/i0[8] ), .A3(\SB3_6/i0[9] ), 
        .ZN(\SB3_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U9380 ( .A1(\SB3_8/i1[9] ), .A2(\SB3_8/i1_7 ), .A3(\SB3_8/i0[10] ), 
        .ZN(\SB3_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U599 ( .A1(\SB3_16/i0_3 ), .A2(\SB3_16/i0[10] ), .A3(\SB3_16/i0_4 ), 
        .ZN(n1721) );
  NAND3_X1 \SB3_22/Component_Function_4/N4  ( .A1(\SB3_22/i1[9] ), .A2(
        \SB3_22/i1_5 ), .A3(\SB3_22/i0_4 ), .ZN(
        \SB3_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U5210 ( .A1(\SB3_7/i1_7 ), .A2(\SB3_7/i0[8] ), .A3(\SB3_7/i0_4 ), 
        .ZN(\SB3_7/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB3_2/Component_Function_5/N1  ( .A1(\SB3_2/i0_0 ), .A2(
        \SB3_2/i3[0] ), .ZN(\SB3_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_0/N2  ( .A1(\SB3_16/i0[8] ), .A2(
        \SB3_16/i0[7] ), .A3(\SB3_16/i0[6] ), .ZN(
        \SB3_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 U4957 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i3[0] ), .ZN(
        \SB3_1/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB3_3/Component_Function_5/N1  ( .A1(\SB3_3/i0_0 ), .A2(
        \SB3_3/i3[0] ), .ZN(\SB3_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U10748 ( .A1(\SB3_14/i0[10] ), .A2(\SB3_14/i0_3 ), .A3(
        \SB3_14/i0[6] ), .ZN(n4412) );
  NAND3_X1 U5151 ( .A1(\SB3_27/i0_3 ), .A2(\SB3_27/i0[10] ), .A3(
        \SB3_27/i0[6] ), .ZN(\SB3_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U9627 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i0_3 ), .A3(\SB3_14/i0_4 ), 
        .ZN(\SB3_14/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U12016 ( .A1(\SB3_13/i0_3 ), .A2(\SB3_13/i1[9] ), .ZN(n5032) );
  NAND3_X1 \SB3_25/Component_Function_2/N3  ( .A1(\SB3_25/i0_3 ), .A2(
        \SB3_25/i0[8] ), .A3(\SB3_25/i0[9] ), .ZN(
        \SB3_25/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 \SB3_31/Component_Function_0/N1  ( .A1(\SB3_31/i0[10] ), .A2(
        \SB3_31/i0[9] ), .ZN(\SB3_31/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB3_7/Component_Function_1/N1  ( .A1(\SB3_7/i0_3 ), .A2(
        \SB3_7/i1[9] ), .ZN(\SB3_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3183 ( .A1(\SB3_31/i0[10] ), .A2(\SB3_31/i1[9] ), .A3(
        \SB3_31/i1_7 ), .ZN(n5064) );
  NAND2_X1 \SB3_30/Component_Function_5/N1  ( .A1(\SB3_30/i0_0 ), .A2(
        \SB3_30/i3[0] ), .ZN(\SB3_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U9524 ( .A1(\SB3_1/i1[9] ), .A2(\SB3_1/i1_7 ), .A3(\SB3_1/i0[10] ), 
        .ZN(\SB3_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_3/Component_Function_3/N2  ( .A1(\SB3_3/i0_0 ), .A2(
        \SB3_3/i0_3 ), .A3(\SB3_3/i0_4 ), .ZN(
        \SB3_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_1/Component_Function_2/N1  ( .A1(\SB3_1/i1_5 ), .A2(
        \SB3_1/i0[10] ), .A3(\SB3_1/i1[9] ), .ZN(
        \SB3_1/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 \SB3_11/Component_Function_0/N1  ( .A1(\SB3_11/i0[10] ), .A2(
        \SB3_11/i0[9] ), .ZN(\SB3_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U9422 ( .A1(\SB3_3/i0[10] ), .A2(\SB3_3/i1[9] ), .A3(\SB3_3/i1_7 ), 
        .ZN(n4645) );
  NAND3_X1 U3277 ( .A1(\SB3_28/i0[8] ), .A2(\SB3_28/i3[0] ), .A3(\SB3_28/i1_5 ), .ZN(n863) );
  NAND3_X1 U591 ( .A1(\SB3_28/i0[10] ), .A2(\SB3_28/i1[9] ), .A3(\SB3_28/i1_7 ), .ZN(\SB3_28/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U12492 ( .A1(\SB3_10/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_10/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_10/Component_Function_4/NAND4_in[3] ), .A4(n5307), .ZN(
        \SB3_10/buf_output[4] ) );
  NAND3_X1 U3031 ( .A1(\SB3_26/i1_5 ), .A2(\SB3_26/i0[8] ), .A3(\SB3_26/i3[0] ), .ZN(\SB3_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U9390 ( .A1(\SB3_11/i1_5 ), .A2(\SB3_11/i0[8] ), .A3(\SB3_11/i3[0] ), .ZN(\SB3_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4678 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0[7] ), .A3(\SB3_30/i0_0 ), 
        .ZN(\SB3_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U5023 ( .A1(\SB3_19/i0_0 ), .A2(\SB3_19/i0_3 ), .A3(\SB3_19/i0_4 ), 
        .ZN(\SB3_19/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 \SB4_27/BUF_4  ( .I(\SB3_28/buf_output[4] ), .Z(\SB4_27/i0_4 ) );
  NAND3_X1 \SB3_29/Component_Function_2/N4  ( .A1(\SB3_29/i1_5 ), .A2(
        \SB3_29/i0_0 ), .A3(\SB3_29/i0_4 ), .ZN(
        \SB3_29/Component_Function_2/NAND4_in[3] ) );
  BUF_X2 U9438 ( .I(\SB3_3/buf_output[1] ), .Z(\SB4_31/i0[6] ) );
  INV_X1 \SB4_20/INV_1  ( .I(\SB3_24/buf_output[1] ), .ZN(\SB4_20/i1_7 ) );
  INV_X1 U3457 ( .I(\SB3_24/buf_output[5] ), .ZN(\SB4_24/i1_5 ) );
  BUF_X2 U304 ( .I(\SB3_27/buf_output[0] ), .Z(\SB4_22/i0[9] ) );
  BUF_X2 U9532 ( .I(\SB3_11/buf_output[1] ), .Z(\SB4_7/i0[6] ) );
  CLKBUF_X2 \SB4_9/BUF_0  ( .I(\SB3_14/buf_output[0] ), .Z(\SB4_9/i0[9] ) );
  CLKBUF_X2 \SB4_2/BUF_1  ( .I(\SB3_6/buf_output[1] ), .Z(\SB4_2/i0[6] ) );
  CLKBUF_X2 U9612 ( .I(\SB3_29/buf_output[1] ), .Z(\SB4_25/i0[6] ) );
  CLKBUF_X2 U1430 ( .I(\SB3_8/buf_output[0] ), .Z(\SB4_3/i0[9] ) );
  CLKBUF_X2 U2452 ( .I(\SB3_16/buf_output[1] ), .Z(\SB4_12/i0[6] ) );
  CLKBUF_X2 U241 ( .I(\SB3_15/buf_output[4] ), .Z(\SB4_14/i0_4 ) );
  CLKBUF_X2 \SB4_7/BUF_4  ( .I(\SB3_8/buf_output[4] ), .Z(\SB4_7/i0_4 ) );
  BUF_X2 U5043 ( .I(\SB3_16/buf_output[4] ), .Z(\SB4_15/i0_4 ) );
  CLKBUF_X2 \SB4_3/BUF_4  ( .I(\SB3_4/buf_output[4] ), .Z(\SB4_3/i0_4 ) );
  CLKBUF_X2 U1383 ( .I(\SB3_0/buf_output[4] ), .Z(\SB4_31/i0_4 ) );
  BUF_X2 U9625 ( .I(\SB3_14/buf_output[5] ), .Z(\SB4_14/i0_3 ) );
  INV_X1 U4291 ( .I(\SB3_20/buf_output[5] ), .ZN(\SB4_20/i1_5 ) );
  INV_X1 U9265 ( .I(\SB3_12/buf_output[5] ), .ZN(\SB4_12/i1_5 ) );
  INV_X1 U1579 ( .I(\SB3_0/buf_output[2] ), .ZN(\SB4_29/i1[9] ) );
  INV_X1 U6560 ( .I(\SB3_26/buf_output[2] ), .ZN(\SB4_23/i1[9] ) );
  INV_X1 U2734 ( .I(\SB3_3/buf_output[3] ), .ZN(\SB4_1/i0[8] ) );
  AND4_X1 U9655 ( .A1(n1743), .A2(\SB3_17/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB3_17/Component_Function_5/NAND4_in[0] ), .A4(n4425), .Z(n3984)
         );
  AND4_X1 U5107 ( .A1(\SB3_14/Component_Function_5/NAND4_in[1] ), .A2(n1628), 
        .A3(\SB3_14/Component_Function_5/NAND4_in[0] ), .A4(
        \SB3_14/Component_Function_5/NAND4_in[2] ), .Z(n1495) );
  NAND3_X1 U5503 ( .A1(\SB4_16/i0_4 ), .A2(\SB4_16/i1[9] ), .A3(\SB4_16/i1_5 ), 
        .ZN(n2923) );
  NAND3_X1 U4856 ( .A1(\SB4_20/i0_0 ), .A2(\SB4_20/i1_5 ), .A3(\SB4_20/i0_4 ), 
        .ZN(n1457) );
  NAND3_X1 U5027 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i1_5 ), .A3(\SB4_23/i0_4 ), 
        .ZN(n2778) );
  NAND2_X1 \SB4_23/Component_Function_5/N1  ( .A1(\SB4_23/i0_0 ), .A2(
        \SB4_23/i3[0] ), .ZN(\SB4_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_23/Component_Function_2/N3  ( .A1(\SB4_23/i0_3 ), .A2(n3974), 
        .A3(\SB4_23/i0[9] ), .ZN(\SB4_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U5092 ( .A1(\SB4_28/i0[6] ), .A2(\SB4_28/i0[9] ), .A3(\SB4_28/i0_4 ), .ZN(n2453) );
  NAND3_X1 \SB4_23/Component_Function_3/N2  ( .A1(\SB4_23/i0_0 ), .A2(
        \SB4_23/i0_3 ), .A3(\SB4_23/i0_4 ), .ZN(
        \SB4_23/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U3099 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i1[9] ), .ZN(
        \SB4_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U4974 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i0_4 ), .A3(n5442), .ZN(n2558) );
  NAND4_X1 U3 ( .A1(\SB4_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_14/Component_Function_3/NAND4_in[3] ), .A4(
        \SB4_14/Component_Function_3/NAND4_in[2] ), .ZN(n6643) );
  NAND3_X1 U24 ( .A1(\SB4_20/i0_4 ), .A2(\SB4_20/i0_0 ), .A3(\SB4_20/i0_3 ), 
        .ZN(n6574) );
  NAND3_X1 U36 ( .A1(\SB4_18/i0[10] ), .A2(\SB4_18/i0_3 ), .A3(\SB4_18/i0[6] ), 
        .ZN(n5130) );
  NAND2_X1 U52 ( .A1(\SB4_0/i0_3 ), .A2(\SB4_0/i1[9] ), .ZN(
        \SB4_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U54 ( .A1(\SB4_12/i0_3 ), .A2(\SB4_12/i0[10] ), .A3(\SB4_12/i0[6] ), 
        .ZN(n4051) );
  NAND3_X1 U95 ( .A1(\SB4_23/i0_0 ), .A2(n3974), .A3(\SB4_23/i0[9] ), .ZN(
        n5252) );
  NAND2_X1 U149 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i3[0] ), .ZN(n5547) );
  NAND3_X1 U163 ( .A1(\SB4_28/i0_4 ), .A2(\SB4_28/i0_0 ), .A3(\SB4_28/i1_5 ), 
        .ZN(n6751) );
  NAND3_X1 U169 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i0[6] ), .A3(\SB4_23/i0[10] ), .ZN(\SB4_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U181 ( .A1(\SB4_6/i0_0 ), .A2(\SB4_6/i1_7 ), .A3(\SB4_6/i3[0] ), 
        .ZN(n4861) );
  NAND3_X1 U208 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i1_7 ), .A3(\SB4_23/i3[0] ), 
        .ZN(n2775) );
  NAND3_X1 U235 ( .A1(\SB4_29/i0_0 ), .A2(\SB4_29/i3[0] ), .A3(\SB4_29/i1_7 ), 
        .ZN(n3312) );
  NAND3_X1 U250 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0_3 ), .A3(\SB4_16/i0[7] ), 
        .ZN(n4957) );
  NAND3_X1 U270 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i1[9] ), .A3(\SB4_12/i1_5 ), 
        .ZN(\SB4_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U314 ( .A1(\SB4_25/i0[10] ), .A2(\SB4_25/i0_3 ), .A3(n6266), .ZN(
        n7566) );
  NAND3_X1 U333 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i0_3 ), .A3(\SB4_10/i0[7] ), 
        .ZN(n3158) );
  INV_X1 U361 ( .I(\SB3_16/buf_output[5] ), .ZN(\SB4_16/i1_5 ) );
  AND4_X1 U572 ( .A1(\SB3_30/Component_Function_0/NAND4_in[1] ), .A2(
        \SB3_30/Component_Function_0/NAND4_in[3] ), .A3(
        \SB3_30/Component_Function_0/NAND4_in[0] ), .A4(n1183), .Z(n5438) );
  CLKBUF_X2 U573 ( .I(\SB3_11/buf_output[4] ), .Z(\SB4_10/i0_4 ) );
  CLKBUF_X2 U579 ( .I(\SB3_26/buf_output[0] ), .Z(\SB4_21/i0[9] ) );
  CLKBUF_X2 U581 ( .I(\SB3_24/buf_output[1] ), .Z(\SB4_20/i0[6] ) );
  BUF_X2 U583 ( .I(\SB3_0/buf_output[1] ), .Z(\SB4_28/i0[6] ) );
  BUF_X2 U585 ( .I(\SB3_13/buf_output[1] ), .Z(\SB4_9/i0[6] ) );
  BUF_X2 U586 ( .I(\SB3_28/buf_output[1] ), .Z(\SB4_24/i0[6] ) );
  NAND3_X1 U587 ( .A1(\SB3_19/i0[6] ), .A2(\SB3_19/i1[9] ), .A3(\SB3_19/i0_3 ), 
        .ZN(\SB3_19/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U589 ( .A1(\SB3_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_13/Component_Function_5/NAND4_in[1] ), .ZN(n5815) );
  NAND2_X1 U594 ( .A1(\SB3_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_2/NAND4_in[1] ), .ZN(n5864) );
  NAND2_X1 U595 ( .A1(n4967), .A2(\SB3_11/Component_Function_2/NAND4_in[2] ), 
        .ZN(n5865) );
  NAND3_X1 U597 ( .A1(\SB3_2/i0[10] ), .A2(\SB3_2/i1_5 ), .A3(\SB3_2/i1[9] ), 
        .ZN(n7428) );
  NAND3_X1 U598 ( .A1(\SB3_3/i1[9] ), .A2(\SB3_3/i0_3 ), .A3(\SB3_3/i0[6] ), 
        .ZN(\SB3_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U600 ( .A1(\SB3_0/i0[9] ), .A2(\SB3_0/i0[10] ), .A3(\SB3_0/i0_3 ), 
        .ZN(\SB3_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U602 ( .A1(\SB3_19/i0[6] ), .A2(\SB3_19/i0_3 ), .A3(\SB3_19/i0[10] ), .ZN(\SB3_19/Component_Function_2/NAND4_in[1] ) );
  AOI21_X1 U603 ( .A1(\SB3_20/i3[0] ), .A2(\SB3_20/i0_0 ), .B(n5670), .ZN(
        n5669) );
  NAND3_X1 U604 ( .A1(\SB3_8/i0_0 ), .A2(\SB3_8/i0_3 ), .A3(\SB3_8/i0_4 ), 
        .ZN(\SB3_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U605 ( .A1(\SB3_28/i0[9] ), .A2(\SB3_28/i0[6] ), .A3(\SB3_28/i0_4 ), 
        .ZN(n5479) );
  NAND3_X1 U606 ( .A1(\SB3_22/i0[9] ), .A2(\SB3_22/i0_4 ), .A3(\SB3_22/i0[6] ), 
        .ZN(n7364) );
  NAND3_X1 U608 ( .A1(\SB3_0/i0[8] ), .A2(\SB3_0/i1_5 ), .A3(\SB3_0/i3[0] ), 
        .ZN(n1475) );
  NAND3_X1 U614 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i0[6] ), .A3(\SB3_7/i0_0 ), 
        .ZN(n1594) );
  NAND3_X1 U615 ( .A1(\SB3_13/i0[8] ), .A2(\SB3_13/i0[7] ), .A3(\SB3_13/i0[6] ), .ZN(\SB3_13/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U618 ( .A1(\SB3_0/i0[9] ), .A2(\SB3_0/i0[6] ), .A3(\SB3_0/i0_4 ), 
        .ZN(n7145) );
  NAND3_X1 U619 ( .A1(\SB3_14/i0[6] ), .A2(\SB3_14/i0_3 ), .A3(\SB3_14/i1[9] ), 
        .ZN(n4050) );
  NAND3_X1 U621 ( .A1(\SB3_16/i0_3 ), .A2(\SB3_16/i0[8] ), .A3(\SB3_16/i0[9] ), 
        .ZN(\SB3_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U630 ( .A1(\SB3_23/i0[10] ), .A2(\SB3_23/i1_5 ), .A3(\SB3_23/i1[9] ), .ZN(n5728) );
  NAND3_X1 U631 ( .A1(\SB3_27/i0_4 ), .A2(\SB3_27/i0_0 ), .A3(\SB3_27/i1_5 ), 
        .ZN(n7452) );
  NAND3_X1 U635 ( .A1(\SB3_30/i0[9] ), .A2(\SB3_30/i1_5 ), .A3(\SB3_30/i0[6] ), 
        .ZN(n6204) );
  NAND3_X1 U636 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i0[6] ), .A3(\SB3_0/i1[9] ), 
        .ZN(n7176) );
  NAND2_X1 U637 ( .A1(\SB3_26/i0_0 ), .A2(\SB3_26/i3[0] ), .ZN(n7344) );
  NAND3_X1 U639 ( .A1(\SB3_1/i0_4 ), .A2(\SB3_1/i1_7 ), .A3(\SB3_1/i0[8] ), 
        .ZN(n6589) );
  NAND2_X1 U641 ( .A1(\SB3_16/i0_0 ), .A2(\SB3_16/i3[0] ), .ZN(
        \SB3_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U642 ( .A1(\SB3_8/i0_0 ), .A2(\SB3_8/i0[7] ), .A3(\SB3_8/i0_3 ), 
        .ZN(\SB3_8/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U643 ( .A1(\SB3_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_25/Component_Function_3/NAND4_in[1] ), .ZN(n7500) );
  NAND3_X1 U647 ( .A1(\SB3_2/i1_5 ), .A2(\SB3_2/i0[8] ), .A3(\SB3_2/i3[0] ), 
        .ZN(n6915) );
  NAND3_X1 U652 ( .A1(\SB3_5/i0[10] ), .A2(\SB3_5/i1[9] ), .A3(\SB3_5/i1_7 ), 
        .ZN(\SB3_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U655 ( .A1(\SB3_11/i0[10] ), .A2(\SB3_11/i0[6] ), .A3(\SB3_11/i0_0 ), .ZN(\SB3_11/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 U659 ( .A1(\SB3_13/i0[10] ), .A2(\SB3_13/i0[9] ), .ZN(
        \SB3_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U662 ( .A1(\SB3_0/i0[10] ), .A2(\SB3_0/i1[9] ), .A3(\SB3_0/i1_7 ), 
        .ZN(n4096) );
  NAND3_X1 U664 ( .A1(\SB3_3/i1[9] ), .A2(\SB3_3/i0_4 ), .A3(\SB3_3/i0_3 ), 
        .ZN(n2498) );
  NAND3_X1 U665 ( .A1(\SB3_27/i0_0 ), .A2(\SB3_27/i0[6] ), .A3(\SB3_27/i0[10] ), .ZN(\SB3_27/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X2 U671 ( .I(\MC_ARK_ARC_1_4/buf_output[114] ), .Z(\SB3_12/i0[9] ) );
  CLKBUF_X2 U672 ( .I(\MC_ARK_ARC_1_4/buf_output[4] ), .Z(\SB3_31/i0_4 ) );
  BUF_X2 U673 ( .I(\MC_ARK_ARC_1_4/buf_output[151] ), .Z(\SB3_6/i0[6] ) );
  OAI21_X1 U676 ( .A1(n3177), .A2(n2152), .B(\SB2_4_15/i0_3 ), .ZN(n6347) );
  NAND3_X1 U680 ( .A1(\SB2_4_25/i0[10] ), .A2(\SB2_4_25/i0_3 ), .A3(
        \SB2_4_25/i0[9] ), .ZN(n7044) );
  NAND3_X1 U684 ( .A1(\SB2_4_25/i0[10] ), .A2(\SB2_4_25/i0_3 ), .A3(
        \SB2_4_25/i0_4 ), .ZN(n7446) );
  NAND3_X1 U685 ( .A1(\SB2_4_16/i0_0 ), .A2(\SB2_4_16/i0_3 ), .A3(
        \SB2_4_16/i0_4 ), .ZN(n6809) );
  NAND3_X1 U686 ( .A1(\SB2_4_22/i0[10] ), .A2(\SB2_4_22/i0[9] ), .A3(
        \SB2_4_22/i0_3 ), .ZN(n6797) );
  NAND3_X1 U688 ( .A1(\SB2_4_14/i0_3 ), .A2(\SB2_4_14/i1[9] ), .A3(
        \SB2_4_14/i0[6] ), .ZN(\SB2_4_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U689 ( .A1(\SB2_4_2/i0[9] ), .A2(\SB2_4_2/i0[10] ), .A3(
        \SB2_4_2/i0_3 ), .ZN(n5941) );
  NAND3_X1 U690 ( .A1(\SB2_4_6/i0_4 ), .A2(\SB2_4_6/i0_0 ), .A3(\SB2_4_6/i1_5 ), .ZN(\SB2_4_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U692 ( .A1(\SB2_4_3/i1[9] ), .A2(\SB2_4_3/i0_3 ), .A3(
        \SB2_4_3/i0[6] ), .ZN(\SB2_4_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U694 ( .A1(\SB2_4_26/i0_3 ), .A2(\SB2_4_26/i0[9] ), .A3(
        \SB2_4_26/i0[10] ), .ZN(\SB2_4_26/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U695 ( .A1(\SB2_4_16/i0_3 ), .A2(\SB2_4_16/i0[10] ), .A3(
        \SB2_4_16/i0[9] ), .ZN(n7388) );
  NAND3_X1 U697 ( .A1(\SB2_4_10/i0[10] ), .A2(\SB2_4_10/i0[9] ), .A3(
        \SB2_4_10/i0_3 ), .ZN(\SB2_4_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U699 ( .A1(\SB2_4_7/i0_3 ), .A2(\SB2_4_7/i0[8] ), .A3(
        \SB2_4_7/i0[9] ), .ZN(n5762) );
  NAND3_X1 U701 ( .A1(\SB2_4_28/i0_3 ), .A2(\SB2_4_28/i0[9] ), .A3(
        \SB2_4_28/i0[10] ), .ZN(\SB2_4_28/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U706 ( .A1(\SB2_4_23/i0_0 ), .A2(\SB2_4_23/i1_5 ), .A3(
        \SB2_4_23/i0_4 ), .ZN(\SB2_4_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U711 ( .A1(\SB2_4_2/i3[0] ), .A2(\SB2_4_2/i0[8] ), .A3(
        \SB2_4_2/i1_5 ), .ZN(\SB2_4_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U719 ( .A1(\SB2_4_15/i0[10] ), .A2(\SB2_4_15/i1[9] ), .A3(
        \SB2_4_15/i1_7 ), .ZN(\SB2_4_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U723 ( .A1(\SB2_4_22/i0[10] ), .A2(\SB2_4_22/i0_4 ), .A3(
        \SB2_4_22/i0_3 ), .ZN(n7019) );
  NAND3_X1 U725 ( .A1(\SB2_4_19/i0_3 ), .A2(\SB2_4_19/i1_7 ), .A3(
        \SB2_4_19/i0[8] ), .ZN(\SB2_4_19/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U726 ( .A1(\SB2_4_18/i0_3 ), .A2(\SB2_4_18/i0_4 ), .A3(
        \SB2_4_18/i0[10] ), .ZN(n6127) );
  NAND3_X1 U727 ( .A1(\SB2_4_26/i0_0 ), .A2(\SB2_4_26/i1_5 ), .A3(
        \SB2_4_26/i0_4 ), .ZN(n7151) );
  NAND3_X1 U731 ( .A1(\SB2_4_25/i0_3 ), .A2(\SB2_4_25/i0_4 ), .A3(
        \SB2_4_25/i1[9] ), .ZN(n2783) );
  NAND3_X1 U737 ( .A1(\SB2_4_28/i0_3 ), .A2(\SB2_4_28/i0_4 ), .A3(
        \SB2_4_28/i0_0 ), .ZN(\SB2_4_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U740 ( .A1(\SB2_4_31/i1_5 ), .A2(\SB2_4_31/i0[8] ), .A3(
        \SB2_4_31/i3[0] ), .ZN(\SB2_4_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U742 ( .A1(\SB2_4_29/i0_4 ), .A2(\SB2_4_29/i1_7 ), .A3(
        \SB2_4_29/i0[8] ), .ZN(n4832) );
  NAND3_X1 U744 ( .A1(\SB2_4_14/i0_3 ), .A2(\SB2_4_14/i0_0 ), .A3(
        \SB2_4_14/i0[7] ), .ZN(n7462) );
  INV_X1 U747 ( .I(\SB1_4_29/buf_output[5] ), .ZN(\SB2_4_29/i1_5 ) );
  CLKBUF_X2 U748 ( .I(\SB1_4_25/buf_output[1] ), .Z(\SB2_4_21/i0[6] ) );
  BUF_X2 U750 ( .I(\SB1_4_23/buf_output[3] ), .Z(\SB2_4_21/i0[10] ) );
  BUF_X2 U754 ( .I(\SB1_4_8/buf_output[1] ), .Z(\SB2_4_4/i0[6] ) );
  CLKBUF_X2 U758 ( .I(\SB1_4_9/buf_output[0] ), .Z(\SB2_4_4/i0[9] ) );
  NAND3_X1 U759 ( .A1(\SB2_4_19/i1[9] ), .A2(\SB2_4_19/i0_4 ), .A3(
        \SB2_4_19/i0_3 ), .ZN(\SB2_4_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U763 ( .A1(\SB2_4_29/i0[6] ), .A2(\SB2_4_29/i0[10] ), .A3(
        \SB2_4_29/i0_0 ), .ZN(n6257) );
  NAND3_X1 U767 ( .A1(\SB2_4_2/i0[6] ), .A2(\SB1_4_7/buf_output[0] ), .A3(
        \SB2_4_2/i0_4 ), .ZN(n6087) );
  CLKBUF_X2 U768 ( .I(\SB1_4_0/buf_output[1] ), .Z(\SB2_4_28/i0[6] ) );
  NAND3_X1 U770 ( .A1(\SB1_4_20/i0[6] ), .A2(\SB1_4_20/i0_4 ), .A3(
        \SB1_4_20/i0[9] ), .ZN(n6134) );
  NAND2_X1 U774 ( .A1(\SB1_4_20/i0_0 ), .A2(\SB1_4_20/i3[0] ), .ZN(n6502) );
  NAND3_X1 U775 ( .A1(\SB1_4_14/i0[6] ), .A2(\SB1_4_14/i0[8] ), .A3(
        \SB1_4_14/i0[7] ), .ZN(\SB1_4_14/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U777 ( .A1(\SB1_4_31/i0_3 ), .A2(\SB1_4_31/i0[10] ), .A3(
        \SB1_4_31/i0_4 ), .ZN(\SB1_4_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U779 ( .A1(\SB1_4_25/i0_0 ), .A2(\SB1_4_25/i1_5 ), .A3(
        \SB1_4_25/i0_4 ), .ZN(n890) );
  NAND2_X1 U782 ( .A1(\SB1_4_27/i0[6] ), .A2(n6701), .ZN(
        \SB1_4_27/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U794 ( .A1(\SB1_4_27/i0[10] ), .A2(\SB1_4_27/i0[9] ), .ZN(n6931) );
  NAND3_X1 U796 ( .A1(\SB1_4_9/i0[9] ), .A2(\SB1_4_9/i0_4 ), .A3(
        \SB1_4_9/i0[6] ), .ZN(n6788) );
  NAND3_X1 U797 ( .A1(\SB1_4_29/i0[10] ), .A2(\SB1_4_29/i1[9] ), .A3(
        \SB1_4_29/i1_7 ), .ZN(n4132) );
  NAND3_X1 U798 ( .A1(\SB1_4_23/i0_3 ), .A2(\SB1_4_23/i0[9] ), .A3(
        \SB1_4_23/i0[8] ), .ZN(n7016) );
  NAND3_X1 U800 ( .A1(\SB1_4_14/i0[9] ), .A2(\SB1_4_14/i0[6] ), .A3(
        \SB1_4_14/i1_5 ), .ZN(n6829) );
  NAND3_X1 U803 ( .A1(\SB1_4_4/i0_4 ), .A2(\SB1_4_4/i0[6] ), .A3(
        \SB1_4_4/i0[9] ), .ZN(n6872) );
  NAND3_X1 U806 ( .A1(\SB1_4_18/i0[6] ), .A2(\SB1_4_18/i0_3 ), .A3(
        \SB1_4_18/i1[9] ), .ZN(n5775) );
  NAND3_X1 U811 ( .A1(\SB1_4_24/i0[9] ), .A2(\SB1_4_24/i1_5 ), .A3(
        \SB1_4_24/i0[6] ), .ZN(\SB1_4_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U817 ( .A1(\SB1_4_20/i0[8] ), .A2(\SB1_4_20/i0_4 ), .A3(
        \SB1_4_20/i1_7 ), .ZN(n7517) );
  NAND3_X1 U819 ( .A1(\SB1_4_15/i0_4 ), .A2(\SB1_4_15/i1_5 ), .A3(
        \SB1_4_15/i1[9] ), .ZN(n4350) );
  NAND3_X1 U824 ( .A1(\SB1_4_16/i0[10] ), .A2(\SB1_4_16/i1[9] ), .A3(
        \SB1_4_16/i1_7 ), .ZN(n7081) );
  NAND3_X1 U825 ( .A1(\SB1_4_8/i0_0 ), .A2(\SB1_4_8/i1_5 ), .A3(\SB1_4_8/i0_4 ), .ZN(\SB1_4_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U828 ( .A1(\SB1_4_27/i3[0] ), .A2(\SB1_4_27/i0[8] ), .A3(
        \SB1_4_27/i1_5 ), .ZN(n6800) );
  NAND3_X1 U829 ( .A1(\SB1_4_7/i0[8] ), .A2(\SB1_4_7/i3[0] ), .A3(
        \SB1_4_7/i1_5 ), .ZN(n6129) );
  NAND3_X1 U830 ( .A1(\SB1_4_14/i0_4 ), .A2(\SB1_4_14/i0_0 ), .A3(
        \SB1_4_14/i1_5 ), .ZN(n6220) );
  NAND3_X1 U832 ( .A1(\SB1_4_27/i1_7 ), .A2(\SB1_4_27/i3[0] ), .A3(
        \RI1[4][26] ), .ZN(n7001) );
  NAND3_X1 U833 ( .A1(\SB1_4_20/i0[10] ), .A2(\SB1_4_20/i0[6] ), .A3(
        \SB1_4_20/i0_3 ), .ZN(n6485) );
  NAND3_X1 U836 ( .A1(\SB1_4_14/i0_3 ), .A2(\SB1_4_14/i0[10] ), .A3(
        \SB1_4_14/i0[9] ), .ZN(n6778) );
  NAND3_X1 U838 ( .A1(\SB1_4_21/i0[6] ), .A2(\SB1_4_21/i1_5 ), .A3(
        \SB1_4_21/i0[9] ), .ZN(n7540) );
  NAND3_X1 U841 ( .A1(\SB1_4_4/i0[8] ), .A2(\SB1_4_4/i0_3 ), .A3(
        \SB1_4_4/i1_7 ), .ZN(n6241) );
  NAND3_X1 U842 ( .A1(\SB1_4_6/i0[9] ), .A2(\SB1_4_6/i1_5 ), .A3(
        \SB1_4_6/i0[6] ), .ZN(n6655) );
  NAND3_X1 U843 ( .A1(\SB1_4_26/i0[6] ), .A2(\SB1_4_26/i0_3 ), .A3(
        \SB1_4_26/i0[10] ), .ZN(n4079) );
  NAND2_X1 U845 ( .A1(n7003), .A2(n4186), .ZN(n5585) );
  NAND3_X1 U861 ( .A1(\SB1_4_6/i0[9] ), .A2(\RI1[4][155] ), .A3(
        \SB1_4_6/i0[8] ), .ZN(n6952) );
  NAND3_X1 U862 ( .A1(\SB1_4_23/i0[9] ), .A2(\SB1_4_23/i0_4 ), .A3(
        \SB1_4_23/i0[6] ), .ZN(n3242) );
  NAND3_X1 U868 ( .A1(\SB1_4_18/i0_3 ), .A2(\SB1_4_18/i0[9] ), .A3(
        \SB1_4_18/i0[10] ), .ZN(n7431) );
  NAND3_X1 U871 ( .A1(\SB1_4_23/i0[8] ), .A2(\SB1_4_23/i0_4 ), .A3(
        \SB1_4_23/i1_7 ), .ZN(n7203) );
  NAND3_X1 U873 ( .A1(\SB1_4_9/i0_0 ), .A2(\SB1_4_9/i1_5 ), .A3(\SB1_4_9/i0_4 ), .ZN(n2538) );
  NAND3_X1 U877 ( .A1(\SB1_4_1/i0[9] ), .A2(\SB1_4_1/i0[8] ), .A3(
        \SB1_4_1/i0_3 ), .ZN(n6160) );
  NAND2_X1 U878 ( .A1(\SB1_4_17/i3[0] ), .A2(\SB1_4_17/i0_0 ), .ZN(n3796) );
  NAND3_X1 U880 ( .A1(\SB1_4_24/i0[9] ), .A2(\SB1_4_24/i0_4 ), .A3(
        \SB1_4_24/i0[6] ), .ZN(n6871) );
  NAND3_X1 U881 ( .A1(\SB1_4_0/i0[8] ), .A2(\SB1_4_0/i1_7 ), .A3(\RI1[4][191] ), .ZN(\SB1_4_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U885 ( .A1(\SB1_4_14/i0_4 ), .A2(\SB1_4_14/i1_5 ), .A3(
        \SB1_4_14/i1[9] ), .ZN(n5990) );
  NAND3_X1 U889 ( .A1(\SB1_4_16/i0[10] ), .A2(\SB1_4_16/i1_5 ), .A3(
        \SB1_4_16/i1[9] ), .ZN(\SB1_4_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U892 ( .A1(\SB1_4_21/i0[10] ), .A2(\SB1_4_21/i1[9] ), .A3(
        \SB1_4_21/i1_5 ), .ZN(n6670) );
  NAND3_X1 U901 ( .A1(\SB1_4_17/i3[0] ), .A2(\SB1_4_17/i0[8] ), .A3(
        \SB1_4_17/i1_5 ), .ZN(n6349) );
  NAND3_X1 U902 ( .A1(\SB1_4_25/i0_0 ), .A2(\SB1_4_25/i0[9] ), .A3(
        \SB1_4_25/i0[8] ), .ZN(n6665) );
  NAND3_X1 U905 ( .A1(\SB1_4_9/i0[8] ), .A2(\SB1_4_9/i3[0] ), .A3(
        \SB1_4_9/i1_5 ), .ZN(n6726) );
  NAND3_X1 U907 ( .A1(\SB1_4_21/i0[10] ), .A2(\SB1_4_21/i0_3 ), .A3(
        \SB1_4_21/i0[9] ), .ZN(n7058) );
  NAND3_X1 U916 ( .A1(\SB1_4_29/i3[0] ), .A2(\SB1_4_29/i0_0 ), .A3(
        \SB1_4_29/i1_7 ), .ZN(n7127) );
  NAND3_X1 U917 ( .A1(\SB1_4_17/i0[8] ), .A2(\SB1_4_17/i0_4 ), .A3(
        \SB1_4_17/i1_7 ), .ZN(n6948) );
  NAND3_X1 U918 ( .A1(\SB1_4_1/i3[0] ), .A2(\SB1_4_1/i0[8] ), .A3(
        \SB1_4_1/i1_5 ), .ZN(n6238) );
  NAND3_X1 U920 ( .A1(\SB1_4_31/i0[9] ), .A2(\RI1[4][5] ), .A3(
        \SB1_4_31/i0[8] ), .ZN(\SB1_4_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U925 ( .A1(\SB1_4_10/i1_5 ), .A2(\SB1_4_10/i0_0 ), .A3(
        \SB1_4_10/i0_4 ), .ZN(n7146) );
  NAND3_X1 U926 ( .A1(\SB1_4_17/i0[9] ), .A2(\SB1_4_17/i0[6] ), .A3(
        \SB1_4_17/i0_4 ), .ZN(n6469) );
  NAND3_X1 U928 ( .A1(\SB1_4_16/i0_4 ), .A2(\SB1_4_16/i1_5 ), .A3(
        \SB1_4_16/i0_0 ), .ZN(n3451) );
  INV_X1 U929 ( .I(\MC_ARK_ARC_1_3/buf_output[49] ), .ZN(\SB1_4_23/i1_7 ) );
  BUF_X2 U934 ( .I(\MC_ARK_ARC_1_3/buf_output[124] ), .Z(\SB1_4_11/i0_4 ) );
  BUF_X1 U938 ( .I(\SB1_4_22/i1[9] ), .Z(n6774) );
  INV_X4 U939 ( .I(n5530), .ZN(\RI1[4][26] ) );
  INV_X1 U940 ( .I(\MC_ARK_ARC_1_3/buf_output[150] ), .ZN(\SB1_4_6/i3[0] ) );
  INV_X4 U941 ( .I(n7105), .ZN(\RI1[4][17] ) );
  NAND3_X1 U944 ( .A1(\SB2_3_11/i0_3 ), .A2(\SB2_3_11/i0[6] ), .A3(
        \SB2_3_11/i1[9] ), .ZN(n3810) );
  NAND3_X1 U945 ( .A1(\SB2_3_13/i0_3 ), .A2(\SB2_3_13/i0[9] ), .A3(
        \SB2_3_13/i0[10] ), .ZN(\SB2_3_13/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U947 ( .A1(\SB2_3_2/i0[10] ), .A2(\SB2_3_2/i0_3 ), .A3(
        \SB2_3_2/i0[9] ), .ZN(n7077) );
  NAND3_X1 U950 ( .A1(\SB2_3_14/i0[8] ), .A2(\SB2_3_14/i3[0] ), .A3(
        \SB2_3_14/i1_5 ), .ZN(\SB2_3_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U951 ( .A1(\SB2_3_21/i0[10] ), .A2(\SB2_3_21/i1[9] ), .A3(
        \SB2_3_21/i1_7 ), .ZN(n6920) );
  NAND3_X1 U954 ( .A1(\SB2_3_26/i3[0] ), .A2(\SB2_3_26/i1_5 ), .A3(
        \SB2_3_26/i0[8] ), .ZN(\SB2_3_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U964 ( .A1(\SB2_3_21/i0[8] ), .A2(\SB2_3_21/i3[0] ), .A3(
        \SB2_3_21/i1_5 ), .ZN(\SB2_3_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U967 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0[10] ), .A3(
        \SB2_3_17/i0_4 ), .ZN(n3817) );
  NAND3_X1 U971 ( .A1(\SB2_3_0/i0_4 ), .A2(\SB2_3_0/i1_5 ), .A3(\SB2_3_0/i0_0 ), .ZN(n7341) );
  NAND3_X1 U973 ( .A1(\SB2_3_11/i0_4 ), .A2(\SB2_3_11/i0_0 ), .A3(
        \SB2_3_11/i0_3 ), .ZN(n5606) );
  NAND3_X1 U984 ( .A1(\SB2_3_28/i1[9] ), .A2(\SB1_3_29/buf_output[4] ), .A3(
        \SB2_3_28/i1_5 ), .ZN(n5232) );
  NAND3_X1 U986 ( .A1(\SB2_3_28/i0[9] ), .A2(\SB2_3_28/i0[6] ), .A3(
        \SB1_3_29/buf_output[4] ), .ZN(
        \SB2_3_28/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U987 ( .A1(\SB2_3_17/i0_4 ), .A2(\SB2_3_17/i0_0 ), .A3(
        \SB2_3_17/i1_5 ), .ZN(n4151) );
  NAND3_X1 U990 ( .A1(\SB2_3_29/i0_3 ), .A2(\SB2_3_29/i0_0 ), .A3(
        \SB2_3_29/i0_4 ), .ZN(n6700) );
  NAND3_X1 U994 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0_0 ), .A3(
        \SB2_3_17/i0_4 ), .ZN(n5749) );
  NAND3_X1 U995 ( .A1(\SB2_3_28/i0_0 ), .A2(\SB2_3_28/i0_3 ), .A3(
        \SB1_3_29/buf_output[4] ), .ZN(n7037) );
  NAND3_X1 U997 ( .A1(\SB2_3_31/i0_0 ), .A2(\SB2_3_31/i0[9] ), .A3(
        \SB2_3_31/i0[8] ), .ZN(\SB2_3_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1003 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB1_3_20/buf_output[4] ), .A3(
        \SB2_3_19/i1[9] ), .ZN(\SB2_3_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1004 ( .A1(\SB2_3_28/i0_3 ), .A2(\SB2_3_28/i0[9] ), .A3(
        \SB2_3_28/i0[8] ), .ZN(n7558) );
  NAND3_X1 U1007 ( .A1(\SB2_3_19/i0[7] ), .A2(\SB2_3_19/i0_3 ), .A3(
        \SB2_3_19/i0_0 ), .ZN(n2232) );
  NAND3_X1 U1010 ( .A1(\SB2_3_12/i0_3 ), .A2(n592), .A3(\SB2_3_12/i0_0 ), .ZN(
        \SB2_3_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1016 ( .A1(\SB2_3_3/i0[10] ), .A2(\SB2_3_3/i0_3 ), .A3(
        \SB2_3_3/i0_4 ), .ZN(\SB2_3_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1019 ( .A1(\SB2_3_11/i0[10] ), .A2(\SB2_3_11/i0_3 ), .A3(
        \SB2_3_11/i0[6] ), .ZN(n1698) );
  NAND3_X1 U1020 ( .A1(\SB2_3_29/i0[10] ), .A2(\SB2_3_29/i1_5 ), .A3(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1021 ( .A1(\SB2_3_3/i0[7] ), .A2(\SB2_3_3/i0_3 ), .A3(
        \SB2_3_3/i0_0 ), .ZN(n6044) );
  NAND3_X1 U1023 ( .A1(\SB2_3_21/i0[6] ), .A2(\SB2_3_21/i1_5 ), .A3(
        \SB2_3_21/i0[9] ), .ZN(\SB2_3_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1024 ( .A1(\RI3[3][70] ), .A2(\SB2_3_20/i1_7 ), .A3(
        \SB2_3_20/i0[8] ), .ZN(\SB2_3_20/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 U1026 ( .A1(\SB2_3_28/i0_0 ), .A2(\SB2_3_28/i3[0] ), .ZN(n6167) );
  NAND3_X1 U1028 ( .A1(\SB2_3_29/i0_3 ), .A2(\SB2_3_29/i1[9] ), .A3(n6552), 
        .ZN(n6163) );
  NAND3_X1 U1029 ( .A1(\SB2_3_29/i0_0 ), .A2(\SB2_3_29/i1_7 ), .A3(
        \SB2_3_29/i3[0] ), .ZN(n5460) );
  NAND3_X1 U1031 ( .A1(\SB2_3_23/i0_0 ), .A2(\SB2_3_23/i3[0] ), .A3(
        \SB2_3_23/i1_7 ), .ZN(n7232) );
  NAND3_X1 U1032 ( .A1(\SB2_3_17/i0[9] ), .A2(\SB2_3_17/i0[10] ), .A3(
        \SB2_3_17/i0_3 ), .ZN(n6174) );
  NAND3_X1 U1038 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0[10] ), .A3(
        \SB2_3_0/i0[9] ), .ZN(n5977) );
  NAND3_X1 U1042 ( .A1(\SB2_3_9/i0[10] ), .A2(\SB2_3_9/i0_3 ), .A3(
        \SB2_3_9/i0[9] ), .ZN(n7265) );
  NAND3_X1 U1047 ( .A1(\SB2_3_24/i0_4 ), .A2(\SB2_3_24/i0[8] ), .A3(
        \SB2_3_24/i1_7 ), .ZN(n6940) );
  NAND3_X1 U1049 ( .A1(\SB2_3_17/i0_0 ), .A2(\SB2_3_17/i3[0] ), .A3(
        \SB2_3_17/i1_7 ), .ZN(\SB2_3_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1050 ( .A1(\SB2_3_9/i0_0 ), .A2(\SB2_3_9/i0[9] ), .A3(
        \SB2_3_9/i0[8] ), .ZN(n7061) );
  NAND3_X1 U1051 ( .A1(\SB2_3_28/i1_7 ), .A2(\SB1_3_29/buf_output[4] ), .A3(
        \SB2_3_28/i0[8] ), .ZN(n1182) );
  NAND3_X1 U1052 ( .A1(\SB2_3_22/i0_0 ), .A2(\SB2_3_22/i3[0] ), .A3(
        \SB2_3_22/i1_7 ), .ZN(\SB2_3_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1053 ( .A1(\SB2_3_23/i0_0 ), .A2(\SB2_3_23/i0[10] ), .A3(
        \SB2_3_23/i0[6] ), .ZN(n7128) );
  INV_X1 U1056 ( .I(\SB1_3_25/buf_output[1] ), .ZN(\SB2_3_21/i1_7 ) );
  INV_X1 U1057 ( .I(\SB1_3_9/buf_output[1] ), .ZN(\SB2_3_5/i1_7 ) );
  INV_X1 U1059 ( .I(\SB1_3_12/buf_output[1] ), .ZN(\SB2_3_8/i1_7 ) );
  AND2_X1 U1070 ( .A1(n4892), .A2(n3044), .Z(n6274) );
  NAND3_X1 U1071 ( .A1(\SB2_3_13/i0[10] ), .A2(\SB2_3_13/i1_5 ), .A3(
        \SB2_3_13/i1[9] ), .ZN(\SB2_3_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1075 ( .A1(\SB2_3_18/i0[6] ), .A2(\SB2_3_18/i0_4 ), .A3(
        \SB2_3_18/i0[9] ), .ZN(n6122) );
  NAND3_X1 U1076 ( .A1(\SB2_3_23/i0[9] ), .A2(\SB2_3_23/i0_4 ), .A3(
        \SB2_3_23/i0[6] ), .ZN(n7017) );
  NAND3_X1 U1077 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB2_3_7/i0[6] ), .A3(
        \SB2_3_7/i0[10] ), .ZN(n7255) );
  INV_X1 U1081 ( .I(\SB1_3_26/buf_output[2] ), .ZN(\SB2_3_23/i1[9] ) );
  BUF_X2 U1084 ( .I(\SB1_3_28/buf_output[1] ), .Z(\SB2_3_24/i0[6] ) );
  NAND2_X1 U1091 ( .A1(\SB2_3_21/i0_0 ), .A2(\SB2_3_21/i3[0] ), .ZN(n7012) );
  CLKBUF_X2 U1093 ( .I(\SB1_3_26/buf_output[0] ), .Z(\SB2_3_21/i0[9] ) );
  NAND3_X1 U1099 ( .A1(\SB1_3_13/i0[6] ), .A2(\SB1_3_13/i1_5 ), .A3(
        \SB1_3_13/i0[9] ), .ZN(\SB1_3_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1106 ( .A1(\SB1_3_12/i0[9] ), .A2(\SB1_3_12/i0[8] ), .A3(
        \SB1_3_12/i0_3 ), .ZN(n3246) );
  NAND3_X1 U1108 ( .A1(\SB1_3_5/i0[6] ), .A2(\SB1_3_5/i1_5 ), .A3(
        \SB1_3_5/i0[9] ), .ZN(\SB1_3_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1110 ( .A1(\SB1_3_31/i0_0 ), .A2(\SB1_3_31/i1_5 ), .A3(
        \SB1_3_31/i0_4 ), .ZN(\SB1_3_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1111 ( .A1(\SB1_3_1/i0[9] ), .A2(\SB1_3_1/i0[6] ), .A3(
        \SB1_3_1/i0_4 ), .ZN(n5191) );
  NAND3_X1 U1113 ( .A1(\SB1_3_12/i0[10] ), .A2(\SB1_3_12/i1[9] ), .A3(
        \SB1_3_12/i1_5 ), .ZN(\SB1_3_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1114 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i1[9] ), .A3(
        \SB1_3_17/i1_5 ), .ZN(n5927) );
  NAND3_X1 U1115 ( .A1(\SB1_3_11/i0[8] ), .A2(\SB1_3_11/i1_5 ), .A3(
        \SB1_3_11/i3[0] ), .ZN(n7423) );
  NAND3_X1 U1116 ( .A1(\SB1_3_17/i0[10] ), .A2(\SB1_3_17/i0_3 ), .A3(
        \SB1_3_17/i0[9] ), .ZN(\SB1_3_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1117 ( .A1(\SB1_3_20/i0_3 ), .A2(\SB1_3_20/i0[9] ), .A3(
        \SB1_3_20/i0[8] ), .ZN(n7325) );
  NAND3_X1 U1125 ( .A1(\SB1_3_4/i0[6] ), .A2(\SB1_3_4/i0[9] ), .A3(
        \SB1_3_4/i0_4 ), .ZN(n1361) );
  NAND2_X1 U1134 ( .A1(\SB1_3_25/i0[9] ), .A2(\SB1_3_25/i0[10] ), .ZN(n7188)
         );
  NAND2_X1 U1135 ( .A1(\SB1_3_28/i0[9] ), .A2(\SB1_3_28/i0[10] ), .ZN(n6994)
         );
  NAND3_X1 U1138 ( .A1(\SB1_3_28/i0_0 ), .A2(\SB1_3_28/i0_4 ), .A3(
        \SB1_3_28/i1_5 ), .ZN(n2675) );
  NAND3_X1 U1146 ( .A1(\SB1_3_15/i0[6] ), .A2(\SB1_3_15/i0_3 ), .A3(n5431), 
        .ZN(n5549) );
  NAND3_X1 U1147 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i0[6] ), .A3(
        \SB1_3_26/i1[9] ), .ZN(\SB1_3_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1152 ( .A1(\SB1_3_11/i0[9] ), .A2(\SB1_3_11/i0_3 ), .A3(
        \SB1_3_11/i0[8] ), .ZN(n7185) );
  NAND3_X1 U1157 ( .A1(\SB1_3_3/i0[9] ), .A2(\SB1_3_3/i0_4 ), .A3(
        \SB1_3_3/i0[6] ), .ZN(n6709) );
  NAND3_X1 U1158 ( .A1(\SB1_3_31/i0_0 ), .A2(\SB1_3_31/i1_7 ), .A3(
        \SB1_3_31/i3[0] ), .ZN(n6575) );
  NAND3_X1 U1159 ( .A1(\SB1_3_16/i3[0] ), .A2(\SB1_3_16/i0[8] ), .A3(
        \SB1_3_16/i1_5 ), .ZN(n4639) );
  NAND3_X1 U1163 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i0_0 ), .A3(
        \SB1_3_17/i1_5 ), .ZN(n5716) );
  NAND3_X1 U1167 ( .A1(\SB1_3_25/i0[9] ), .A2(\SB1_3_25/i0_3 ), .A3(
        \SB1_3_25/i0[10] ), .ZN(\SB1_3_25/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1169 ( .A1(\SB1_3_6/i0_4 ), .A2(\SB1_3_6/i0_0 ), .A3(
        \SB1_3_6/i1_5 ), .ZN(n3068) );
  NAND3_X1 U1181 ( .A1(\SB1_3_21/i0_0 ), .A2(\SB1_3_21/i0[10] ), .A3(
        \SB1_3_21/i0[6] ), .ZN(\SB1_3_21/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1182 ( .A1(\SB1_3_8/i0[9] ), .A2(\SB1_3_8/i0_0 ), .A3(
        \SB1_3_8/i0[8] ), .ZN(n5614) );
  BUF_X2 U1188 ( .I(\MC_ARK_ARC_1_2/buf_output[48] ), .Z(\SB1_3_23/i0[9] ) );
  NAND3_X1 U1192 ( .A1(\SB1_3_1/i0[9] ), .A2(\SB1_3_1/i0_3 ), .A3(
        \SB1_3_1/i0[10] ), .ZN(n6869) );
  CLKBUF_X2 U1200 ( .I(\MC_ARK_ARC_1_2/buf_output[19] ), .Z(\SB1_3_28/i0[6] )
         );
  NAND3_X1 U1202 ( .A1(\SB1_3_18/i0[10] ), .A2(\SB1_3_18/i1_5 ), .A3(
        \SB1_3_18/i1[9] ), .ZN(\SB1_3_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1227 ( .A1(\SB1_3_8/i1_5 ), .A2(\SB1_3_8/i0[8] ), .A3(
        \SB1_3_8/i3[0] ), .ZN(\SB1_3_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1232 ( .A1(\SB1_3_0/i0[10] ), .A2(\SB1_3_0/i0_3 ), .A3(
        \SB1_3_0/i0_4 ), .ZN(n6796) );
  NAND2_X1 U1233 ( .A1(\SB1_3_21/i0_0 ), .A2(\SB1_3_21/i3[0] ), .ZN(n5745) );
  NAND3_X1 U1238 ( .A1(\SB1_3_29/i0[10] ), .A2(\SB1_3_29/i1[9] ), .A3(
        \SB1_3_29/i1_7 ), .ZN(n4601) );
  BUF_X2 U1239 ( .I(\MC_ARK_ARC_1_2/buf_output[152] ), .Z(\SB1_3_6/i0_0 ) );
  BUF_X2 U1248 ( .I(\SB1_3_15/i1[9] ), .Z(n5431) );
  NAND3_X1 U1251 ( .A1(\SB2_2_2/i0_3 ), .A2(\SB2_2_2/i0_0 ), .A3(
        \SB2_2_2/i0_4 ), .ZN(\SB2_2_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1254 ( .A1(\SB2_2_31/i0[9] ), .A2(\SB2_2_31/i0_3 ), .A3(
        \SB2_2_31/i0[10] ), .ZN(\SB2_2_31/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1255 ( .A1(\SB2_2_21/i0_0 ), .A2(\SB1_2_22/buf_output[4] ), .A3(
        \SB2_2_21/i1_5 ), .ZN(n7223) );
  NAND3_X1 U1257 ( .A1(\SB2_2_5/i0_3 ), .A2(\SB2_2_5/i0_0 ), .A3(
        \SB2_2_5/i0_4 ), .ZN(\SB2_2_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1276 ( .A1(\SB2_2_13/i0_0 ), .A2(\SB2_2_13/i3[0] ), .A3(
        \SB2_2_13/i1_7 ), .ZN(\SB2_2_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1279 ( .A1(\SB2_2_21/i0[9] ), .A2(\SB1_2_22/buf_output[4] ), .A3(
        \SB2_2_21/i0[6] ), .ZN(n7374) );
  NAND3_X1 U1280 ( .A1(\SB2_2_14/i0[10] ), .A2(\SB2_2_14/i1[9] ), .A3(
        \SB2_2_14/i1_7 ), .ZN(n882) );
  NAND3_X1 U1282 ( .A1(\SB2_2_5/i0[9] ), .A2(\SB2_2_5/i0[6] ), .A3(
        \SB2_2_5/i1_5 ), .ZN(n5799) );
  NAND3_X1 U1293 ( .A1(\SB2_2_2/i0_4 ), .A2(n6267), .A3(\SB2_2_2/i1_5 ), .ZN(
        \SB2_2_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1295 ( .A1(\SB2_2_12/i0_4 ), .A2(\SB2_2_12/i0[8] ), .A3(
        \SB2_2_12/i1_7 ), .ZN(n6536) );
  NAND3_X1 U1304 ( .A1(\SB2_2_8/i0_4 ), .A2(\SB2_2_8/i1_7 ), .A3(
        \SB2_2_8/i0[8] ), .ZN(n7391) );
  NAND3_X1 U1305 ( .A1(\SB2_2_13/i0[9] ), .A2(\SB2_2_13/i0[8] ), .A3(
        \SB2_2_13/i0_3 ), .ZN(n6471) );
  NAND3_X1 U1319 ( .A1(\SB2_2_19/i0[10] ), .A2(\SB2_2_19/i1_7 ), .A3(
        \SB2_2_19/i1[9] ), .ZN(n3943) );
  NAND3_X1 U1324 ( .A1(\SB2_2_17/i0[10] ), .A2(\SB2_2_17/i0_0 ), .A3(
        \SB2_2_17/i0[6] ), .ZN(\SB2_2_17/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1325 ( .A1(\SB2_2_5/i1[9] ), .A2(\SB2_2_5/i0_3 ), .A3(
        \SB2_2_5/i0[6] ), .ZN(\SB2_2_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1327 ( .A1(\SB2_2_21/i0_3 ), .A2(\SB2_2_21/i0[10] ), .A3(
        \SB2_2_21/i0[6] ), .ZN(n7220) );
  NAND3_X1 U1333 ( .A1(\SB2_2_18/i0[6] ), .A2(\SB2_2_18/i0_0 ), .A3(
        \SB2_2_18/i0[10] ), .ZN(\SB2_2_18/Component_Function_5/NAND4_in[1] )
         );
  INV_X1 U1334 ( .I(\SB1_2_12/buf_output[1] ), .ZN(\SB2_2_8/i1_7 ) );
  NAND2_X1 U1335 ( .A1(\SB2_2_21/i0[9] ), .A2(\SB2_2_21/i0[10] ), .ZN(
        \SB2_2_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U1347 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0[10] ), .A3(
        \SB2_2_28/i0[9] ), .ZN(n7539) );
  NAND3_X1 U1352 ( .A1(\SB2_2_8/i0[6] ), .A2(\SB2_2_8/i0[10] ), .A3(
        \SB2_2_8/i0_3 ), .ZN(n7101) );
  NAND3_X1 U1353 ( .A1(\SB2_2_9/i0[6] ), .A2(\SB1_2_14/buf_output[0] ), .A3(
        \SB2_2_9/i1_5 ), .ZN(\SB2_2_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1362 ( .A1(\SB2_2_4/i0_0 ), .A2(\SB2_2_4/i0[9] ), .A3(
        \SB2_2_4/i0[8] ), .ZN(n5453) );
  NAND3_X1 U1386 ( .A1(\SB2_2_20/i1_7 ), .A2(\SB2_2_20/i0[8] ), .A3(
        \SB2_2_20/i0_4 ), .ZN(\SB2_2_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1392 ( .A1(\SB2_2_29/i0[8] ), .A2(\SB2_2_29/i1_5 ), .A3(
        \SB2_2_29/i3[0] ), .ZN(n6177) );
  NAND3_X1 U1393 ( .A1(\SB2_2_14/i0[6] ), .A2(\SB2_2_14/i0[10] ), .A3(
        \SB2_2_14/i0_0 ), .ZN(\SB2_2_14/Component_Function_5/NAND4_in[1] ) );
  INV_X1 U1394 ( .I(\SB1_2_0/buf_output[3] ), .ZN(\SB2_2_30/i0[8] ) );
  NAND3_X1 U1405 ( .A1(\SB1_2_26/i0_3 ), .A2(\SB1_2_26/i0[8] ), .A3(
        \SB1_2_26/i1_7 ), .ZN(\SB1_2_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1406 ( .A1(\SB1_2_0/i1_5 ), .A2(\SB1_2_0/i1[9] ), .A3(
        \SB1_2_0/i0_4 ), .ZN(n7020) );
  NAND3_X1 U1409 ( .A1(\SB1_2_4/i0[10] ), .A2(\SB1_2_4/i1[9] ), .A3(
        \SB1_2_4/i1_7 ), .ZN(n6956) );
  NAND3_X1 U1418 ( .A1(\SB1_2_5/i0_0 ), .A2(\SB1_2_5/i0_3 ), .A3(
        \SB1_2_5/i0[7] ), .ZN(n7346) );
  NAND3_X1 U1419 ( .A1(\SB1_2_29/i0[10] ), .A2(\SB1_2_29/i0[9] ), .A3(
        \RI1[2][17] ), .ZN(\SB1_2_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1421 ( .A1(n3839), .A2(\SB1_2_29/i0_4 ), .A3(\SB1_2_29/i1[9] ), 
        .ZN(n5454) );
  NAND2_X1 U1424 ( .A1(n4077), .A2(n7199), .ZN(n7200) );
  NAND3_X1 U1426 ( .A1(\SB1_2_21/i0[9] ), .A2(\SB1_2_21/i0_4 ), .A3(
        \SB1_2_21/i0[6] ), .ZN(n5128) );
  NAND3_X1 U1429 ( .A1(\SB1_2_2/i0_3 ), .A2(\SB1_2_2/i0_4 ), .A3(
        \SB1_2_2/i1[9] ), .ZN(\SB1_2_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1434 ( .A1(\SB1_2_10/i0[6] ), .A2(\SB1_2_10/i1_5 ), .A3(
        \SB1_2_10/i0[9] ), .ZN(n6907) );
  NAND3_X1 U1435 ( .A1(\SB1_2_3/i0_4 ), .A2(\SB1_2_3/i0_3 ), .A3(
        \SB1_2_3/i0_0 ), .ZN(\SB1_2_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1438 ( .A1(\SB1_2_7/i0[10] ), .A2(\RI1[2][149] ), .A3(
        \SB1_2_7/i0_4 ), .ZN(n2243) );
  NAND2_X1 U1444 ( .A1(\SB1_2_26/i0[9] ), .A2(\SB1_2_26/i0[10] ), .ZN(
        \SB1_2_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U1449 ( .A1(\SB1_2_2/i0_3 ), .A2(\SB1_2_2/i0[6] ), .A3(
        \SB1_2_2/i1[9] ), .ZN(n2725) );
  NAND3_X1 U1451 ( .A1(\SB1_2_5/i0[6] ), .A2(\SB1_2_5/i1_5 ), .A3(
        \SB1_2_5/i0[9] ), .ZN(n6732) );
  NAND3_X1 U1453 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i0_4 ), .A3(
        \SB1_2_18/i1[9] ), .ZN(\SB1_2_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1454 ( .A1(\SB1_2_15/i1_5 ), .A2(\SB1_2_15/i1[9] ), .A3(
        \SB1_2_15/i0[10] ), .ZN(\SB1_2_15/Component_Function_2/NAND4_in[0] )
         );
  NAND3_X1 U1456 ( .A1(\SB1_2_14/i0[9] ), .A2(\SB1_2_14/i0[6] ), .A3(
        \SB1_2_14/i1_5 ), .ZN(\SB1_2_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1460 ( .A1(\SB1_2_4/i0_3 ), .A2(\SB1_2_4/i1_7 ), .A3(
        \SB1_2_4/i0[8] ), .ZN(\SB1_2_4/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1465 ( .A1(\SB1_2_13/i0[10] ), .A2(\SB1_2_13/i1[9] ), .A3(
        \SB1_2_13/i1_7 ), .ZN(n1573) );
  NAND3_X1 U1466 ( .A1(\SB1_2_28/i0[8] ), .A2(\SB1_2_28/i1_5 ), .A3(
        \SB1_2_28/i3[0] ), .ZN(n3455) );
  NAND3_X1 U1468 ( .A1(\SB1_2_8/i0[10] ), .A2(\SB1_2_8/i1[9] ), .A3(
        \SB1_2_8/i1_7 ), .ZN(\SB1_2_8/Component_Function_3/NAND4_in[2] ) );
  OAI21_X1 U1474 ( .A1(\SB1_2_10/i0_4 ), .A2(\SB1_2_10/i0_3 ), .B(n6909), .ZN(
        n6908) );
  NAND3_X1 U1480 ( .A1(\SB1_2_18/i0[10] ), .A2(\SB1_2_18/i1[9] ), .A3(
        \SB1_2_18/i1_7 ), .ZN(n6053) );
  NAND3_X1 U1481 ( .A1(\SB1_2_9/i0[8] ), .A2(\SB1_2_9/i3[0] ), .A3(
        \SB1_2_9/i1_5 ), .ZN(n5474) );
  NAND3_X1 U1482 ( .A1(\SB1_2_26/i0_3 ), .A2(\SB1_2_26/i0_0 ), .A3(
        \SB1_2_26/i0[7] ), .ZN(n5207) );
  NAND3_X1 U1488 ( .A1(\SB1_2_12/i0[6] ), .A2(\SB1_2_12/i0[8] ), .A3(
        \SB1_2_12/i0[7] ), .ZN(\SB1_2_12/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1489 ( .A1(\SB1_2_17/i0[6] ), .A2(\SB1_2_17/i0[8] ), .A3(
        \SB1_2_17/i0[7] ), .ZN(n6400) );
  NAND3_X1 U1490 ( .A1(\SB1_2_24/i0[9] ), .A2(\SB1_2_24/i0[6] ), .A3(
        \SB1_2_24/i1_5 ), .ZN(\SB1_2_24/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U1497 ( .A1(\SB1_2_27/i0[9] ), .A2(\SB1_2_27/i0[10] ), .ZN(n7116)
         );
  NAND3_X1 U1501 ( .A1(\SB1_2_16/i0_3 ), .A2(\SB1_2_16/i0_0 ), .A3(
        \SB1_2_16/i0[7] ), .ZN(n5808) );
  NAND3_X1 U1503 ( .A1(\SB1_2_26/i0[6] ), .A2(\SB1_2_26/i0[8] ), .A3(
        \SB1_2_26/i0[7] ), .ZN(\SB1_2_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1504 ( .A1(\SB1_2_23/i0_0 ), .A2(\SB1_2_23/i0[7] ), .A3(
        \SB1_2_23/i0_3 ), .ZN(n5935) );
  NAND3_X1 U1505 ( .A1(\SB1_2_6/i0_4 ), .A2(\SB1_2_6/i1[9] ), .A3(
        \SB1_2_6/i1_5 ), .ZN(n6310) );
  NAND3_X1 U1511 ( .A1(\SB1_2_12/i1_5 ), .A2(\RI1[2][116] ), .A3(
        \SB1_2_12/i0_4 ), .ZN(n2438) );
  NAND3_X1 U1512 ( .A1(\SB1_2_15/i0_0 ), .A2(\RI1[2][101] ), .A3(
        \SB1_2_15/i0_4 ), .ZN(n6693) );
  NAND3_X1 U1513 ( .A1(\SB1_2_9/i0_4 ), .A2(\SB1_2_9/i0[8] ), .A3(
        \SB1_2_9/i1_7 ), .ZN(n7163) );
  NAND3_X1 U1518 ( .A1(\SB1_2_8/i0[10] ), .A2(\SB1_2_8/i0_3 ), .A3(
        \SB1_2_8/i0_4 ), .ZN(n5873) );
  NAND3_X1 U1520 ( .A1(\SB1_2_26/i0_3 ), .A2(\SB1_2_26/i0[10] ), .A3(
        \SB1_2_26/i0[9] ), .ZN(n7358) );
  NAND3_X1 U1533 ( .A1(\SB1_2_4/i0[10] ), .A2(\SB1_2_4/i0_0 ), .A3(
        \SB1_2_4/i0[6] ), .ZN(n3575) );
  NAND2_X1 U1534 ( .A1(\SB1_2_9/i0_0 ), .A2(\SB1_2_9/i3[0] ), .ZN(n5551) );
  NAND3_X1 U1535 ( .A1(\SB1_2_30/i0[10] ), .A2(\SB1_2_30/i0[9] ), .A3(
        \SB1_2_30/i0_3 ), .ZN(n7302) );
  NAND3_X1 U1537 ( .A1(\SB1_2_16/i0_3 ), .A2(\SB1_2_16/i0[6] ), .A3(
        \SB1_2_16/i1[9] ), .ZN(\SB1_2_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1539 ( .A1(\SB1_2_30/i0[6] ), .A2(\SB1_2_30/i0_4 ), .A3(
        \SB1_2_30/i0[9] ), .ZN(n7347) );
  NAND3_X1 U1543 ( .A1(\SB1_2_22/i0[9] ), .A2(\SB1_2_22/i0[8] ), .A3(
        \RI1[2][59] ), .ZN(n7464) );
  NAND3_X1 U1544 ( .A1(\SB1_2_29/i0_4 ), .A2(\SB1_2_29/i0[8] ), .A3(
        \SB1_2_29/i1_7 ), .ZN(n3212) );
  NAND3_X1 U1545 ( .A1(\SB1_2_18/i1_7 ), .A2(\SB1_2_18/i0[8] ), .A3(
        \SB1_2_18/i0_4 ), .ZN(\SB1_2_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1546 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i1_7 ), .A3(
        \SB1_2_18/i0[8] ), .ZN(\SB1_2_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1549 ( .A1(\SB1_2_25/i0[10] ), .A2(\SB1_2_25/i1[9] ), .A3(
        \SB1_2_25/i1_7 ), .ZN(n7237) );
  NAND3_X1 U1553 ( .A1(\SB1_2_8/i0[10] ), .A2(\SB1_2_8/i1[9] ), .A3(
        \SB1_2_8/i1_5 ), .ZN(n4926) );
  NAND3_X1 U1557 ( .A1(\SB1_2_11/i0[10] ), .A2(\SB1_2_11/i0[6] ), .A3(
        \SB1_2_11/i0_3 ), .ZN(n5791) );
  NAND3_X1 U1562 ( .A1(\SB1_2_30/i0_0 ), .A2(\SB1_2_30/i0_3 ), .A3(
        \SB1_2_30/i0[7] ), .ZN(n7400) );
  NAND3_X1 U1564 ( .A1(\SB1_2_1/i0[9] ), .A2(\SB1_2_1/i0[10] ), .A3(
        \SB1_2_1/i0_3 ), .ZN(n7193) );
  INV_X1 U1565 ( .I(\RI1[2][149] ), .ZN(n7286) );
  NAND3_X1 U1567 ( .A1(\SB2_1_7/i0_4 ), .A2(\SB2_1_7/i0_0 ), .A3(
        \SB2_1_7/i1_5 ), .ZN(\SB2_1_7/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1568 ( .A1(\SB2_1_26/i0_0 ), .A2(\SB2_1_26/i0_4 ), .A3(
        \SB2_1_26/i1_5 ), .ZN(n7190) );
  NAND3_X1 U1572 ( .A1(\SB2_1_0/i0[6] ), .A2(\SB2_1_0/i1_5 ), .A3(
        \SB2_1_0/i0[9] ), .ZN(\SB2_1_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1574 ( .A1(\SB2_1_16/i0_4 ), .A2(\SB2_1_16/i0[8] ), .A3(
        \SB2_1_16/i1_7 ), .ZN(n7360) );
  NAND3_X1 U1581 ( .A1(\SB2_1_30/i0[10] ), .A2(\SB2_1_30/i1_7 ), .A3(
        \SB2_1_30/i1[9] ), .ZN(\SB2_1_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1583 ( .A1(\SB2_1_17/i3[0] ), .A2(n3990), .A3(\SB2_1_17/i0[8] ), 
        .ZN(n6569) );
  NAND3_X1 U1587 ( .A1(\SB2_1_19/i0_4 ), .A2(\SB2_1_19/i0[8] ), .A3(
        \SB2_1_19/i1_7 ), .ZN(n7533) );
  NAND3_X1 U1591 ( .A1(\SB2_1_6/i3[0] ), .A2(\SB2_1_6/i1_5 ), .A3(
        \SB2_1_6/i0[8] ), .ZN(n6729) );
  NAND2_X1 U1594 ( .A1(\SB2_1_24/i0[10] ), .A2(\SB2_1_24/i0[9] ), .ZN(n6987)
         );
  NAND3_X1 U1615 ( .A1(\SB2_1_21/i0_0 ), .A2(\SB2_1_21/i0_3 ), .A3(
        \SB2_1_21/i0[7] ), .ZN(n1465) );
  NAND3_X1 U1619 ( .A1(\SB2_1_28/i0_4 ), .A2(\SB2_1_28/i0[8] ), .A3(
        \SB2_1_28/i1_7 ), .ZN(n6803) );
  NAND3_X1 U1622 ( .A1(\SB2_1_27/i1[9] ), .A2(\SB2_1_27/i0_4 ), .A3(
        \SB2_1_27/i1_5 ), .ZN(\SB2_1_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1628 ( .A1(\SB2_1_10/i0_4 ), .A2(\SB2_1_10/i0_0 ), .A3(
        \SB2_1_10/i1_5 ), .ZN(n6683) );
  NAND3_X1 U1634 ( .A1(\SB2_1_11/i0[6] ), .A2(\SB2_1_11/i1_5 ), .A3(
        \SB2_1_11/i0[9] ), .ZN(n7318) );
  NAND2_X1 U1636 ( .A1(\SB2_1_19/i0[9] ), .A2(\SB2_1_19/i0[10] ), .ZN(n5862)
         );
  NAND3_X1 U1637 ( .A1(\SB2_1_24/i0_4 ), .A2(\SB2_1_24/i0[9] ), .A3(
        \SB2_1_24/i0[6] ), .ZN(\SB2_1_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1640 ( .A1(\SB2_1_22/i0[10] ), .A2(\SB2_1_22/i1_7 ), .A3(
        \SB2_1_22/i1[9] ), .ZN(\SB2_1_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1641 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i0_0 ), .A3(
        \SB2_1_15/i0[7] ), .ZN(n7365) );
  NAND3_X1 U1645 ( .A1(\SB2_1_2/i0[7] ), .A2(\SB2_1_2/i0_0 ), .A3(
        \SB2_1_2/i0_3 ), .ZN(n5783) );
  NAND3_X1 U1646 ( .A1(\SB2_1_15/i0[10] ), .A2(\SB2_1_15/i0_3 ), .A3(
        \SB2_1_15/i0[9] ), .ZN(n7252) );
  CLKBUF_X2 U1647 ( .I(\SB1_1_11/buf_output[1] ), .Z(\SB2_1_7/i0[6] ) );
  NAND2_X1 U1649 ( .A1(n1666), .A2(n6517), .ZN(n4840) );
  NAND3_X1 U1650 ( .A1(\SB2_1_1/i0_4 ), .A2(\SB2_1_1/i0_0 ), .A3(
        \SB2_1_1/i1_5 ), .ZN(\SB2_1_1/Component_Function_2/NAND4_in[3] ) );
  INV_X1 U1653 ( .I(\SB1_1_15/buf_output[1] ), .ZN(\SB2_1_11/i1_7 ) );
  NAND3_X1 U1667 ( .A1(\SB2_1_2/i0[9] ), .A2(\SB2_1_2/i0_4 ), .A3(
        \SB2_1_2/i0[6] ), .ZN(n5781) );
  NAND2_X1 U1673 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i0[6] ), .ZN(n6517) );
  NAND3_X1 U1677 ( .A1(\SB1_1_9/i1[9] ), .A2(\SB1_1_9/i0_3 ), .A3(
        \SB1_1_9/i0[6] ), .ZN(\SB1_1_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1683 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i1[9] ), .A3(
        \SB1_1_10/i0_4 ), .ZN(n2589) );
  NAND3_X1 U1691 ( .A1(\SB1_1_29/i0[10] ), .A2(\SB1_1_29/i0_3 ), .A3(
        \SB1_1_29/i0[9] ), .ZN(n7491) );
  NAND3_X1 U1696 ( .A1(\SB1_1_3/i0_4 ), .A2(\SB1_1_3/i0_3 ), .A3(
        \SB1_1_3/i1[9] ), .ZN(n5754) );
  NAND3_X1 U1706 ( .A1(\SB1_1_29/i0_0 ), .A2(\SB1_1_29/i0[8] ), .A3(
        \SB1_1_29/i0[9] ), .ZN(\SB1_1_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1707 ( .A1(\SB1_1_29/i0_0 ), .A2(\SB1_1_29/i1_7 ), .A3(
        \SB1_1_29/i3[0] ), .ZN(\SB1_1_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1709 ( .A1(\SB1_1_10/i0[6] ), .A2(\SB1_1_10/i0[9] ), .A3(
        \SB1_1_10/i0_4 ), .ZN(n5715) );
  NAND3_X1 U1713 ( .A1(\SB1_1_18/i0[9] ), .A2(\SB1_1_18/i0[6] ), .A3(
        \SB1_1_18/i1_5 ), .ZN(\SB1_1_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1714 ( .A1(\SB1_1_8/i0[10] ), .A2(\SB1_1_8/i0_3 ), .A3(
        \SB1_1_8/i0[9] ), .ZN(n5746) );
  NAND3_X1 U1718 ( .A1(\SB1_1_30/i3[0] ), .A2(\SB1_1_30/i0[8] ), .A3(
        \SB1_1_30/i1_5 ), .ZN(n4231) );
  NAND3_X1 U1720 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i0[6] ), .A3(
        \SB1_1_10/i1[9] ), .ZN(n6718) );
  NAND3_X1 U1728 ( .A1(\SB1_1_5/i0[10] ), .A2(\SB1_1_5/i1[9] ), .A3(
        \SB1_1_5/i1_7 ), .ZN(\SB1_1_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1730 ( .A1(\SB1_1_13/i0[10] ), .A2(\SB1_1_13/i0_0 ), .A3(
        \SB1_1_13/i0[6] ), .ZN(\SB1_1_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1739 ( .A1(\SB1_1_27/i0_4 ), .A2(\SB1_1_27/i0_3 ), .A3(
        \SB1_1_27/i1[9] ), .ZN(n6585) );
  NAND3_X1 U1741 ( .A1(\SB1_1_15/i0[8] ), .A2(\SB1_1_15/i3[0] ), .A3(
        \SB1_1_15/i1_5 ), .ZN(n2877) );
  NAND3_X1 U1742 ( .A1(\SB1_1_28/i0_3 ), .A2(\SB1_1_28/i0_0 ), .A3(
        \SB1_1_28/i0[7] ), .ZN(n2430) );
  NAND3_X1 U1745 ( .A1(\SB1_1_5/i0[9] ), .A2(\SB1_1_5/i0_4 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[157] ), .ZN(n6620) );
  NAND3_X1 U1746 ( .A1(\SB1_1_28/i0[8] ), .A2(\SB1_1_28/i1_5 ), .A3(
        \SB1_1_28/i3[0] ), .ZN(n6437) );
  NAND3_X1 U1752 ( .A1(\SB1_1_17/i0_4 ), .A2(\SB1_1_17/i1[9] ), .A3(
        \SB1_1_17/i1_5 ), .ZN(n7481) );
  NAND2_X1 U1756 ( .A1(\SB1_1_30/Component_Function_4/NAND4_in[1] ), .A2(n1922), .ZN(n6673) );
  NAND2_X1 U1770 ( .A1(\SB1_1_6/i0_0 ), .A2(\SB1_1_6/i3[0] ), .ZN(n6937) );
  NAND3_X1 U1774 ( .A1(\SB1_1_4/i0[10] ), .A2(\SB1_1_4/i1[9] ), .A3(
        \SB1_1_4/i1_5 ), .ZN(n6067) );
  NAND3_X1 U1778 ( .A1(\SB1_1_9/i0[10] ), .A2(\SB1_1_9/i1[9] ), .A3(
        \SB1_1_9/i1_5 ), .ZN(n6986) );
  NAND3_X1 U1782 ( .A1(\SB1_1_16/i0_0 ), .A2(\SB1_1_16/i1_5 ), .A3(
        \SB1_1_16/i0_4 ), .ZN(n5709) );
  NAND3_X1 U1783 ( .A1(\SB1_1_14/i0[8] ), .A2(\SB1_1_14/i0[9] ), .A3(
        \SB1_1_14/i0_0 ), .ZN(\SB1_1_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1785 ( .A1(\SB1_1_8/i0[8] ), .A2(\SB1_1_8/i3[0] ), .A3(
        \SB1_1_8/i1_5 ), .ZN(n6664) );
  NAND3_X1 U1789 ( .A1(\SB1_1_28/i0[8] ), .A2(\SB1_1_28/i0[6] ), .A3(
        \SB1_1_28/i0[7] ), .ZN(n6542) );
  NAND3_X1 U1790 ( .A1(\SB1_1_18/i0[8] ), .A2(\SB1_1_18/i3[0] ), .A3(
        \SB1_1_18/i1_5 ), .ZN(\SB1_1_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1791 ( .A1(\SB1_1_25/i0[8] ), .A2(\SB1_1_25/i1_5 ), .A3(
        \SB1_1_25/i3[0] ), .ZN(n5809) );
  NAND3_X1 U1805 ( .A1(\SB1_1_27/i0_4 ), .A2(\SB1_1_27/i1_7 ), .A3(
        \SB1_1_27/i0[8] ), .ZN(n6740) );
  NAND2_X1 U1808 ( .A1(\SB1_1_1/i0_0 ), .A2(\SB1_1_1/i3[0] ), .ZN(n6022) );
  NAND3_X1 U1809 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0_0 ), .A3(
        \SB1_1_6/i0_4 ), .ZN(n7228) );
  NAND3_X1 U1811 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i0[9] ), .A3(
        \SB1_1_0/i0[8] ), .ZN(n6979) );
  BUF_X2 U1816 ( .I(\MC_ARK_ARC_1_0/buf_output[0] ), .Z(\SB1_1_31/i0[9] ) );
  NAND3_X1 U1817 ( .A1(\SB1_1_0/i0[10] ), .A2(\SB1_1_0/i0_3 ), .A3(
        \SB1_1_0/i0[9] ), .ZN(\SB1_1_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1832 ( .A1(\SB1_1_30/i0_0 ), .A2(\SB1_1_30/i0[8] ), .A3(
        \SB1_1_30/i0[9] ), .ZN(n6880) );
  NAND3_X1 U1835 ( .A1(\SB1_1_3/i0[8] ), .A2(\SB1_1_3/i3[0] ), .A3(
        \SB1_1_3/i1_5 ), .ZN(n6480) );
  NAND3_X1 U1839 ( .A1(\SB1_1_5/i0[6] ), .A2(\SB1_1_5/i1_5 ), .A3(
        \SB1_1_5/i0[9] ), .ZN(\SB1_1_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1840 ( .A1(\SB2_0_30/i0_3 ), .A2(\SB2_0_30/i0_4 ), .A3(
        \SB2_0_30/i0[10] ), .ZN(n5858) );
  NAND3_X1 U1841 ( .A1(\SB2_0_15/i0_3 ), .A2(\RI3[0][100] ), .A3(
        \SB1_0_18/buf_output[2] ), .ZN(n7181) );
  NAND3_X1 U1844 ( .A1(\SB2_0_15/i0_3 ), .A2(\SB2_0_15/i0[6] ), .A3(n1508), 
        .ZN(n6205) );
  NAND3_X1 U1847 ( .A1(\SB2_0_14/i0_3 ), .A2(\SB2_0_14/i0_4 ), .A3(
        \SB2_0_14/i1[9] ), .ZN(\SB2_0_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1851 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0[9] ), .A3(
        \SB2_0_4/i0[8] ), .ZN(\SB2_0_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1857 ( .A1(\RI3[0][52] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i0[10] ), .ZN(\SB2_0_23/Component_Function_0/NAND4_in[2] )
         );
  NAND3_X1 U1863 ( .A1(\SB2_0_0/i0[9] ), .A2(\SB2_0_0/i0[6] ), .A3(
        \SB2_0_0/i1_5 ), .ZN(n6034) );
  NAND3_X1 U1867 ( .A1(\SB2_0_15/i0[9] ), .A2(\SB2_0_15/i0_3 ), .A3(
        \SB2_0_15/i0[10] ), .ZN(n7180) );
  NAND3_X1 U1868 ( .A1(\SB2_0_0/i0[6] ), .A2(\RI3[0][190] ), .A3(
        \SB2_0_0/i0[9] ), .ZN(n5604) );
  NAND3_X1 U1869 ( .A1(\SB2_0_13/i0_0 ), .A2(\SB2_0_13/i0[10] ), .A3(
        \SB2_0_13/i0[6] ), .ZN(\SB2_0_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1876 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0[10] ), .A3(
        \SB2_0_4/i0[9] ), .ZN(n6256) );
  NAND3_X1 U1879 ( .A1(\SB2_0_6/i0[10] ), .A2(\SB2_0_6/i0_0 ), .A3(
        \SB2_0_6/i0[6] ), .ZN(n6990) );
  NAND3_X1 U1882 ( .A1(\SB2_0_26/i0_3 ), .A2(\SB2_0_26/i0_4 ), .A3(
        \SB2_0_26/i1[9] ), .ZN(\SB2_0_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1888 ( .A1(\SB2_0_10/i0[10] ), .A2(\SB2_0_10/i0[6] ), .A3(
        \SB2_0_10/i0_3 ), .ZN(n6031) );
  NAND3_X1 U1896 ( .A1(\RI3[0][52] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i0_0 ), .ZN(\SB2_0_23/Component_Function_3/NAND4_in[1] ) );
  OAI21_X1 U1897 ( .A1(n5434), .A2(n1508), .B(\SB2_0_15/i0_3 ), .ZN(n5188) );
  NAND3_X1 U1898 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i0_0 ), .A3(
        \SB2_0_28/i0_4 ), .ZN(\SB2_0_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1900 ( .A1(\SB2_0_30/i0_3 ), .A2(\SB2_0_30/i0[8] ), .A3(
        \SB2_0_30/i0[9] ), .ZN(n7508) );
  NAND3_X1 U1901 ( .A1(\SB2_0_21/i0[6] ), .A2(\SB2_0_21/i0[9] ), .A3(
        \SB2_0_21/i0_4 ), .ZN(\SB2_0_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1902 ( .A1(\SB2_0_27/i0_0 ), .A2(\SB2_0_27/i1_5 ), .A3(
        \RI3[0][28] ), .ZN(n748) );
  NAND3_X1 U1903 ( .A1(\SB2_0_7/i0_0 ), .A2(\SB2_0_7/i3[0] ), .A3(
        \SB2_0_7/i1_7 ), .ZN(\SB2_0_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1905 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i0[6] ), .A3(
        \SB2_0_25/i0[10] ), .ZN(\SB2_0_25/Component_Function_2/NAND4_in[1] )
         );
  INV_X1 U1906 ( .I(\SB1_0_1/buf_output[5] ), .ZN(\SB2_0_1/i1_5 ) );
  INV_X1 U1909 ( .I(\SB1_0_25/buf_output[0] ), .ZN(\SB2_0_20/i3[0] ) );
  INV_X2 U1913 ( .I(\SB2_0_15/i0[7] ), .ZN(\RI3[0][100] ) );
  INV_X2 U1923 ( .I(\RI3[0][141] ), .ZN(\SB2_0_8/i0[8] ) );
  INV_X2 U1926 ( .I(n6651), .ZN(n594) );
  NAND2_X1 U1928 ( .A1(\SB1_0_5/i0[9] ), .A2(\SB1_0_5/i0[10] ), .ZN(
        \SB1_0_5/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U1929 ( .A1(n2609), .A2(\SB1_0_15/Component_Function_4/NAND4_in[1] ), .ZN(n7160) );
  NAND3_X1 U1933 ( .A1(n5433), .A2(\SB1_0_28/i0[10] ), .A3(\SB1_0_28/i0_3 ), 
        .ZN(\SB1_0_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1934 ( .A1(\SB1_0_9/i1[9] ), .A2(\SB1_0_9/i0_3 ), .A3(
        \SB1_0_9/i0[6] ), .ZN(\SB1_0_9/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U1938 ( .A1(\SB1_0_14/i0_0 ), .A2(\SB1_0_14/i3[0] ), .ZN(n6068) );
  NAND3_X1 U1940 ( .A1(\SB1_0_30/i0[6] ), .A2(\SB1_0_30/i1[9] ), .A3(
        \SB1_0_30/i0_3 ), .ZN(n6085) );
  NAND3_X1 U1944 ( .A1(\SB1_0_31/i0[10] ), .A2(\SB1_0_31/i1_5 ), .A3(
        \SB1_0_31/i1[9] ), .ZN(\SB1_0_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1945 ( .A1(n5433), .A2(\SB1_0_28/i0[8] ), .A3(\SB1_0_28/i1_7 ), 
        .ZN(\SB1_0_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1946 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0_4 ), .A3(
        \SB1_0_15/i1[9] ), .ZN(n7156) );
  NAND3_X1 U1952 ( .A1(\SB1_0_17/i0[10] ), .A2(\SB1_0_17/i1_7 ), .A3(
        \SB1_0_17/i1[9] ), .ZN(n6576) );
  NAND3_X1 U1958 ( .A1(\SB1_0_5/i0[10] ), .A2(\SB1_0_5/i0_4 ), .A3(
        \SB1_0_5/i0_3 ), .ZN(n7161) );
  NAND3_X1 U1977 ( .A1(\SB1_0_14/i0_4 ), .A2(\SB1_0_14/i1_5 ), .A3(
        \SB1_0_14/i0_0 ), .ZN(n4917) );
  NAND3_X1 U1981 ( .A1(\SB1_0_30/i0_4 ), .A2(\SB1_0_30/i0_0 ), .A3(
        \SB1_0_30/i1_5 ), .ZN(n7515) );
  BUF_X2 U1992 ( .I(n241), .Z(\SB1_0_11/i0[6] ) );
  NAND2_X1 U1997 ( .A1(\SB1_0_25/i1_5 ), .A2(n7269), .ZN(n7268) );
  NAND3_X1 U1998 ( .A1(n5433), .A2(\SB1_0_28/i0_0 ), .A3(\SB1_0_28/i0_3 ), 
        .ZN(\SB1_0_28/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U2010 ( .I(n285), .ZN(\SB1_0_15/i3[0] ) );
  NAND2_X2 U2015 ( .A1(\SB2_2_18/i0_3 ), .A2(\SB2_2_18/i1[9] ), .ZN(
        \SB2_2_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U2018 ( .A1(\SB2_3_21/i0[6] ), .A2(\SB2_3_21/i0_3 ), .A3(
        \SB2_3_21/i0[10] ), .ZN(n6853) );
  NAND3_X2 U2020 ( .A1(\SB1_4_19/i0[7] ), .A2(\SB1_4_19/i0_3 ), .A3(
        \SB1_4_19/i0_0 ), .ZN(\SB1_4_19/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 U2029 ( .I(\MC_ARK_ARC_1_1/buf_output[85] ), .Z(\SB1_2_17/i0[6] ) );
  BUF_X4 U2030 ( .I(\SB1_3_25/buf_output[1] ), .Z(\SB2_3_21/i0[6] ) );
  NAND3_X2 U2046 ( .A1(\SB1_2_10/buf_output[1] ), .A2(\SB2_2_6/i0_4 ), .A3(
        \SB2_2_6/i0[9] ), .ZN(n7060) );
  NAND3_X2 U2047 ( .A1(\SB2_4_2/i0[9] ), .A2(\SB2_4_2/i1_5 ), .A3(
        \SB2_4_2/i0[6] ), .ZN(n5703) );
  NAND3_X2 U2049 ( .A1(\SB1_4_19/i0_0 ), .A2(\SB1_4_19/i0_4 ), .A3(
        \SB1_4_19/i0_3 ), .ZN(n934) );
  INV_X2 U2066 ( .I(\SB1_2_26/buf_output[0] ), .ZN(\SB2_2_21/i3[0] ) );
  NAND3_X2 U2068 ( .A1(\SB1_4_19/i0_3 ), .A2(\SB1_4_19/i1[9] ), .A3(
        \SB1_4_19/i0_4 ), .ZN(n2467) );
  BUF_X2 U2069 ( .I(\SB1_3_8/buf_output[2] ), .Z(\SB2_3_5/i0_0 ) );
  BUF_X8 U2097 ( .I(\RI1[5][11] ), .Z(\SB3_30/i0_3 ) );
  NAND3_X2 U2105 ( .A1(\SB3_13/i1_5 ), .A2(\SB3_13/i1[9] ), .A3(\SB3_13/i0_4 ), 
        .ZN(n6954) );
  BUF_X4 U2107 ( .I(n278), .Z(\SB1_0_19/i0_0 ) );
  INV_X8 U2120 ( .I(\RI1[2][59] ), .ZN(\SB1_2_22/i1_5 ) );
  NAND3_X2 U2121 ( .A1(\SB1_3_12/i1[9] ), .A2(\SB1_3_12/i0_3 ), .A3(
        \SB1_3_12/i0[6] ), .ZN(\SB1_3_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U2123 ( .A1(\SB2_4_9/i0_3 ), .A2(\SB2_4_9/i0_4 ), .A3(
        \SB2_4_9/i1[9] ), .ZN(n5140) );
  NAND3_X2 U2127 ( .A1(\SB1_0_13/i0_3 ), .A2(\SB1_0_13/i0[10] ), .A3(
        \SB1_0_13/i0[9] ), .ZN(n3358) );
  NAND3_X2 U2130 ( .A1(\SB1_4_14/i3[0] ), .A2(\SB1_4_14/i1_5 ), .A3(
        \SB1_4_14/i0[8] ), .ZN(n4493) );
  NAND3_X2 U2131 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i0_4 ), .A3(
        \SB1_3_10/i1[9] ), .ZN(n2309) );
  BUF_X2 U2137 ( .I(\MC_ARK_ARC_1_2/buf_output[128] ), .Z(\SB1_3_10/i0_0 ) );
  INV_X2 U2143 ( .I(\MC_ARK_ARC_1_2/buf_output[188] ), .ZN(\SB1_3_0/i1[9] ) );
  NAND2_X2 U2145 ( .A1(\SB1_0_19/i0_3 ), .A2(\SB1_0_19/i0[7] ), .ZN(n3434) );
  BUF_X4 U2151 ( .I(\SB1_3_23/buf_output[0] ), .Z(\SB2_3_18/i0[9] ) );
  NAND2_X2 U2160 ( .A1(\SB4_6/i0_3 ), .A2(\SB4_6/i1[9] ), .ZN(
        \SB4_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U2169 ( .A1(\SB2_4_23/i0[8] ), .A2(\SB2_4_23/i0[7] ), .A3(
        \SB2_4_23/i0[6] ), .ZN(\SB2_4_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X2 U2172 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i1[9] ), .ZN(
        \SB1_0_23/Component_Function_1/NAND4_in[0] ) );
  INV_X2 U2176 ( .I(\MC_ARK_ARC_1_0/buf_output[123] ), .ZN(\SB1_1_11/i0[8] )
         );
  NAND3_X2 U2178 ( .A1(\SB2_1_3/i0_4 ), .A2(\SB2_1_3/i0_3 ), .A3(
        \SB2_1_3/i1[9] ), .ZN(n4305) );
  NAND3_X2 U2179 ( .A1(\SB2_0_18/i0[9] ), .A2(\SB2_0_18/i0_0 ), .A3(
        \SB2_0_18/i0[8] ), .ZN(\SB2_0_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U2182 ( .A1(\SB3_13/i1_5 ), .A2(\SB3_13/i0[6] ), .A3(\SB3_13/i0[9] ), .ZN(\SB3_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U2184 ( .A1(\SB2_1_31/i0_0 ), .A2(\SB2_1_31/i3[0] ), .A3(
        \SB2_1_31/i1_7 ), .ZN(\SB2_1_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U2188 ( .A1(\SB2_1_13/i0_3 ), .A2(\SB2_1_13/i0[8] ), .A3(
        \SB2_1_13/i0[9] ), .ZN(\SB2_1_13/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X2 U2194 ( .I(\MC_ARK_ARC_1_4/buf_output[132] ), .Z(\SB3_9/i0[9] ) );
  CLKBUF_X2 U2197 ( .I(\SB3_6/buf_output[5] ), .Z(n6057) );
  CLKBUF_X4 U2201 ( .I(\SB2_3_22/buf_output[1] ), .Z(\RI5[3][79] ) );
  NAND3_X1 U2203 ( .A1(\SB1_4_15/i0[8] ), .A2(\SB1_4_15/i0[7] ), .A3(
        \SB1_4_15/i0[6] ), .ZN(\SB1_4_15/Component_Function_0/NAND4_in[1] ) );
  INV_X2 U2210 ( .I(\SB1_4_15/i0_4 ), .ZN(\SB1_4_15/i0[7] ) );
  NAND4_X1 U2212 ( .A1(n4284), .A2(n1916), .A3(
        \SB4_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_13/Component_Function_3/NAND4_in[3] ), .ZN(n5750) );
  CLKBUF_X4 U2220 ( .I(\SB1_4_8/buf_output[4] ), .Z(\RI3[4][148] ) );
  INV_X1 U2225 ( .I(\SB1_4_7/buf_output[5] ), .ZN(\SB2_4_7/i1_5 ) );
  CLKBUF_X4 U2231 ( .I(\SB1_4_7/buf_output[5] ), .Z(\SB2_4_7/i0_3 ) );
  BUF_X2 U2233 ( .I(\MC_ARK_ARC_1_2/buf_output[25] ), .Z(\SB1_3_27/i0[6] ) );
  NAND3_X1 U2238 ( .A1(\SB1_4_24/i0_0 ), .A2(\SB1_4_24/i3[0] ), .A3(
        \SB1_4_24/i1_7 ), .ZN(n7559) );
  NAND3_X1 U2239 ( .A1(\SB1_4_11/i0_4 ), .A2(\SB1_4_11/i0_0 ), .A3(
        \SB1_4_11/i1_5 ), .ZN(n4053) );
  NAND3_X1 U2240 ( .A1(\SB1_4_11/i0[9] ), .A2(\SB1_4_11/i0[6] ), .A3(
        \SB1_4_11/i0_4 ), .ZN(n6821) );
  NAND3_X1 U2246 ( .A1(\SB1_4_11/i1[9] ), .A2(\SB1_4_11/i0_4 ), .A3(
        \SB1_4_11/i1_5 ), .ZN(n2009) );
  NAND3_X1 U2247 ( .A1(\SB3_10/i0_3 ), .A2(\SB3_10/i1[9] ), .A3(\SB3_10/i0_4 ), 
        .ZN(n5366) );
  NAND3_X1 U2249 ( .A1(\SB3_10/i0_4 ), .A2(\SB3_10/i0[6] ), .A3(\SB3_10/i0[9] ), .ZN(n5519) );
  NAND3_X1 U2258 ( .A1(\SB3_10/i0[8] ), .A2(\SB3_10/i0_4 ), .A3(\SB3_10/i1_7 ), 
        .ZN(\SB3_10/Component_Function_1/NAND4_in[3] ) );
  BUF_X2 U2260 ( .I(\SB3_19/buf_output[0] ), .Z(\SB4_14/i0[9] ) );
  NAND3_X1 U2261 ( .A1(\SB2_1_18/i0_0 ), .A2(\SB2_1_18/i0_4 ), .A3(
        \SB2_1_18/i1_5 ), .ZN(\SB2_1_18/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2268 ( .A1(\SB2_1_18/i0_0 ), .A2(\SB2_1_18/i0_3 ), .A3(
        \SB2_1_18/i0_4 ), .ZN(\SB2_1_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2271 ( .A1(\SB2_1_18/i0[6] ), .A2(\SB2_1_18/i0_0 ), .A3(
        \SB2_1_18/i0[10] ), .ZN(n5336) );
  NAND2_X1 U2273 ( .A1(\SB2_1_18/i0_0 ), .A2(\SB2_1_18/i3[0] ), .ZN(n1400) );
  NAND3_X1 U2274 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB2_1_18/i0_0 ), .A3(
        \SB2_1_18/i0[7] ), .ZN(n1659) );
  NAND3_X1 U2280 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB2_1_18/i0_4 ), .A3(
        \SB2_1_18/i1[9] ), .ZN(n2185) );
  NAND3_X1 U2281 ( .A1(\SB2_1_18/i1[9] ), .A2(\SB2_1_18/i0_3 ), .A3(
        \SB2_1_18/i0[6] ), .ZN(\SB2_1_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2283 ( .A1(\SB2_1_18/i1[9] ), .A2(\SB2_1_18/i1_5 ), .A3(
        \SB2_1_18/i0_4 ), .ZN(\SB2_1_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2294 ( .A1(\SB2_1_18/i0[10] ), .A2(\SB2_1_18/i1_7 ), .A3(
        \SB2_1_18/i1[9] ), .ZN(n3101) );
  NAND3_X1 U2295 ( .A1(\SB2_1_18/i0[10] ), .A2(\SB2_1_18/i1_5 ), .A3(
        \SB2_1_18/i1[9] ), .ZN(\SB2_1_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2298 ( .A1(\SB1_4_21/i0[9] ), .A2(\SB1_4_21/i0[8] ), .A3(
        \SB1_4_21/i0_0 ), .ZN(n3233) );
  NAND3_X1 U2300 ( .A1(\SB1_4_21/i0_0 ), .A2(\SB1_4_21/i0[6] ), .A3(
        \SB1_4_21/i0[10] ), .ZN(\SB1_4_21/Component_Function_5/NAND4_in[1] )
         );
  INV_X1 U2302 ( .I(\MC_ARK_ARC_1_4/buf_output[15] ), .ZN(\SB3_29/i0[8] ) );
  BUF_X2 U2306 ( .I(\MC_ARK_ARC_1_4/buf_output[15] ), .Z(\SB3_29/i0[10] ) );
  NAND3_X1 U2310 ( .A1(\SB4_3/i0[10] ), .A2(\SB4_3/i0_4 ), .A3(\SB4_3/i0_3 ), 
        .ZN(\SB4_3/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U2319 ( .I(\SB3_3/buf_output[5] ), .Z(\SB4_3/i0_3 ) );
  INV_X1 U2322 ( .I(\MC_ARK_ARC_1_2/buf_output[43] ), .ZN(\SB1_3_24/i1_7 ) );
  BUF_X2 U2327 ( .I(\MC_ARK_ARC_1_2/buf_output[43] ), .Z(\SB1_3_24/i0[6] ) );
  INV_X1 U2332 ( .I(\MC_ARK_ARC_1_3/buf_output[13] ), .ZN(\SB1_4_29/i1_7 ) );
  BUF_X2 U2335 ( .I(\MC_ARK_ARC_1_3/buf_output[13] ), .Z(\SB1_4_29/i0[6] ) );
  NAND3_X1 U2337 ( .A1(\SB3_4/i1_7 ), .A2(\SB3_4/i0[8] ), .A3(\SB3_4/i0_4 ), 
        .ZN(\SB3_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2338 ( .A1(\SB2_0_10/i0[10] ), .A2(\SB2_0_10/i1[9] ), .A3(
        \SB2_0_10/i1_7 ), .ZN(\SB2_0_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2339 ( .A1(\SB2_0_10/i0[10] ), .A2(\SB2_0_10/i1[9] ), .A3(
        \SB2_0_10/i1_5 ), .ZN(\SB2_0_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2340 ( .A1(\SB2_0_10/i1[9] ), .A2(\SB2_0_10/i0_3 ), .A3(
        \SB2_0_10/i0_4 ), .ZN(n3583) );
  NAND3_X1 U2342 ( .A1(\SB2_0_10/i1[9] ), .A2(\SB2_0_10/i0_3 ), .A3(
        \SB2_0_10/i0[6] ), .ZN(\SB2_0_10/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U2349 ( .I(n1501), .ZN(\SB2_0_10/i1[9] ) );
  NAND3_X1 U2353 ( .A1(\SB3_11/i0_3 ), .A2(\SB3_11/i0[9] ), .A3(
        \SB3_11/i0[10] ), .ZN(\SB3_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2355 ( .A1(\SB3_11/i0[10] ), .A2(\SB3_11/i0_4 ), .A3(\SB3_11/i0_3 ), .ZN(\SB3_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2361 ( .A1(\SB3_11/i0_3 ), .A2(\SB3_11/i0_4 ), .A3(\SB3_11/i0_0 ), 
        .ZN(\SB3_11/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U2364 ( .A1(\SB3_11/i0_3 ), .A2(\SB3_11/i1[9] ), .ZN(
        \SB3_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2366 ( .A1(\SB2_4_9/i0[6] ), .A2(\SB2_4_9/i0_3 ), .A3(
        \SB2_4_9/i0[10] ), .ZN(n4635) );
  NAND3_X1 U2369 ( .A1(\SB2_4_9/i0_0 ), .A2(\SB2_4_9/i0_3 ), .A3(
        \SB2_4_9/i0_4 ), .ZN(n4255) );
  CLKBUF_X4 U2372 ( .I(\SB2_4_10/buf_output[4] ), .Z(\RI5[4][136] ) );
  NAND3_X1 U2374 ( .A1(\SB4_1/i0[9] ), .A2(\SB4_1/i0_0 ), .A3(\SB4_1/i0[8] ), 
        .ZN(\SB4_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2381 ( .A1(\SB2_4_8/i1_5 ), .A2(\SB2_4_8/i0[8] ), .A3(
        \SB2_4_8/i3[0] ), .ZN(\SB2_4_8/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X4 U2382 ( .I(\MC_ARK_ARC_1_4/buf_output[154] ), .Z(\SB3_6/i0_4 ) );
  NAND3_X1 U2384 ( .A1(\SB4_4/i0_0 ), .A2(\SB4_4/i3[0] ), .A3(\SB4_4/i1_7 ), 
        .ZN(\SB4_4/Component_Function_4/NAND4_in[1] ) );
  CLKBUF_X4 U2390 ( .I(\SB3_24/buf_output[5] ), .Z(\SB4_24/i0_3 ) );
  CLKBUF_X4 U2393 ( .I(\MC_ARK_ARC_1_4/buf_output[3] ), .Z(\SB3_31/i0[10] ) );
  NAND3_X1 U2397 ( .A1(\SB2_4_28/i1_5 ), .A2(n4000), .A3(\SB2_4_28/i3[0] ), 
        .ZN(\SB2_4_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2399 ( .A1(\SB2_4_28/i1_5 ), .A2(\SB2_4_28/i0[6] ), .A3(
        \SB2_4_28/i0[9] ), .ZN(\SB2_4_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2401 ( .A1(\SB2_4_28/i0_0 ), .A2(\SB2_4_28/i0_4 ), .A3(
        \SB2_4_28/i1_5 ), .ZN(n5806) );
  NAND3_X1 U2415 ( .A1(\SB2_3_22/i0_3 ), .A2(\SB2_3_22/i1[9] ), .A3(
        \RI3[3][58] ), .ZN(\SB2_3_22/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2427 ( .A1(\SB2_3_22/i1[9] ), .A2(\SB2_3_22/i1_7 ), .A3(
        \SB2_3_22/i0[10] ), .ZN(\SB2_3_22/Component_Function_3/NAND4_in[2] )
         );
  NAND2_X1 U2433 ( .A1(\SB2_3_22/i0_3 ), .A2(\SB2_3_22/i1[9] ), .ZN(
        \SB2_3_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2441 ( .A1(\SB2_3_22/i1_5 ), .A2(\SB2_3_22/i0[10] ), .A3(
        \SB2_3_22/i1[9] ), .ZN(\SB2_3_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2445 ( .A1(\SB2_3_22/i1[9] ), .A2(\SB2_3_22/i0_3 ), .A3(
        \SB2_3_22/i0[6] ), .ZN(\SB2_3_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2446 ( .A1(\SB2_3_22/i1[9] ), .A2(\SB2_3_22/i1_5 ), .A3(
        \RI3[3][58] ), .ZN(\SB2_3_22/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U2448 ( .I(\SB2_4_8/buf_output[2] ), .Z(\RI5[4][158] ) );
  NAND3_X1 U2450 ( .A1(\SB1_4_22/i0[9] ), .A2(\SB1_4_22/i0[8] ), .A3(
        \RI1[4][59] ), .ZN(\SB1_4_22/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 U2463 ( .A1(n6774), .A2(\RI1[4][59] ), .ZN(
        \SB1_4_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2464 ( .A1(\SB1_4_22/i0_4 ), .A2(\SB1_4_22/i0_0 ), .A3(
        \RI1[4][59] ), .ZN(n3563) );
  NAND3_X1 U2465 ( .A1(\RI1[4][59] ), .A2(\SB1_4_22/i0[10] ), .A3(
        \SB1_4_22/i0_4 ), .ZN(\SB1_4_22/Component_Function_0/NAND4_in[2] ) );
  INV_X1 U2470 ( .I(\MC_ARK_ARC_1_3/buf_output[43] ), .ZN(\SB1_4_24/i1_7 ) );
  BUF_X2 U2478 ( .I(\MC_ARK_ARC_1_3/buf_output[43] ), .Z(\SB1_4_24/i0[6] ) );
  NAND3_X1 U2480 ( .A1(\SB3_5/i0[9] ), .A2(\SB3_5/i0[6] ), .A3(\SB3_5/i0_4 ), 
        .ZN(\SB3_5/Component_Function_5/NAND4_in[3] ) );
  CLKBUF_X4 U2481 ( .I(\SB3_29/buf_output[5] ), .Z(\SB4_29/i0_3 ) );
  NAND3_X1 U2483 ( .A1(\SB2_3_3/i0[7] ), .A2(\SB2_3_3/i0[8] ), .A3(
        \SB2_3_3/i0[6] ), .ZN(\SB2_3_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 U2484 ( .A1(\SB3_28/i0_0 ), .A2(\SB3_28/i3[0] ), .ZN(
        \SB3_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2487 ( .A1(\SB3_28/i0[10] ), .A2(\SB3_28/i0_0 ), .A3(
        \SB3_28/i0[6] ), .ZN(\SB3_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2491 ( .A1(\SB3_28/i1_5 ), .A2(\SB3_28/i0_0 ), .A3(\SB3_28/i0_4 ), 
        .ZN(\SB3_28/Component_Function_2/NAND4_in[3] ) );
  CLKBUF_X4 U2498 ( .I(\MC_ARK_ARC_1_4/buf_output[20] ), .Z(\SB3_28/i0_0 ) );
  NAND3_X1 U2499 ( .A1(\SB4_3/i0[9] ), .A2(\SB4_3/i0[6] ), .A3(\SB4_3/i0_4 ), 
        .ZN(\SB4_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2500 ( .A1(\SB4_3/i0_3 ), .A2(\SB4_3/i0[6] ), .A3(\SB4_3/i1[9] ), 
        .ZN(n7258) );
  NAND3_X1 U2502 ( .A1(\SB4_3/i0[6] ), .A2(\SB4_3/i0_3 ), .A3(\SB4_3/i0[10] ), 
        .ZN(n2728) );
  CLKBUF_X2 U2505 ( .I(\SB3_7/buf_output[1] ), .Z(\SB4_3/i0[6] ) );
  NAND3_X1 U2507 ( .A1(\SB2_4_15/i1_5 ), .A2(\SB2_4_15/i0[8] ), .A3(
        \SB2_4_15/i3[0] ), .ZN(\SB2_4_15/Component_Function_3/NAND4_in[3] ) );
  BUF_X2 U2508 ( .I(\MC_ARK_ARC_1_4/buf_output[82] ), .Z(\SB3_18/i0_4 ) );
  INV_X1 U2510 ( .I(\SB1_3_10/buf_output[3] ), .ZN(\SB2_3_8/i0[8] ) );
  BUF_X2 U2515 ( .I(\SB1_3_10/buf_output[3] ), .Z(\SB2_3_8/i0[10] ) );
  NAND3_X1 U2516 ( .A1(\SB1_3_10/i0[6] ), .A2(\SB1_3_10/i1[9] ), .A3(
        \SB1_3_10/i0_3 ), .ZN(\SB1_3_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2518 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i0[10] ), .A3(
        \SB1_3_10/i0[6] ), .ZN(\SB1_3_10/Component_Function_2/NAND4_in[1] ) );
  INV_X1 U2521 ( .I(\MC_ARK_ARC_1_4/buf_output[73] ), .ZN(\SB3_19/i1_7 ) );
  BUF_X2 U2524 ( .I(\MC_ARK_ARC_1_4/buf_output[73] ), .Z(\SB3_19/i0[6] ) );
  INV_X1 U2525 ( .I(\MC_ARK_ARC_1_4/buf_output[48] ), .ZN(\SB3_23/i3[0] ) );
  BUF_X2 U2526 ( .I(\MC_ARK_ARC_1_4/buf_output[48] ), .Z(\SB3_23/i0[9] ) );
  NAND3_X1 U2528 ( .A1(\SB1_4_24/i0_0 ), .A2(\SB1_4_24/i0_3 ), .A3(
        \SB1_4_24/i0_4 ), .ZN(\SB1_4_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2529 ( .A1(\SB1_4_24/i0[6] ), .A2(\SB1_4_24/i0[10] ), .A3(
        \SB1_4_24/i0_3 ), .ZN(n6096) );
  NAND3_X1 U2532 ( .A1(\SB1_4_24/i0_0 ), .A2(\SB1_4_24/i0[7] ), .A3(
        \SB1_4_24/i0_3 ), .ZN(n4764) );
  NAND2_X1 U2533 ( .A1(\SB1_4_24/i0_3 ), .A2(\SB1_4_24/i1[9] ), .ZN(
        \SB1_4_24/Component_Function_1/NAND4_in[0] ) );
  CLKBUF_X4 U2534 ( .I(\SB3_2/buf_output[5] ), .Z(\SB4_2/i0_3 ) );
  INV_X1 U2535 ( .I(\SB3_0/buf_output[3] ), .ZN(\SB4_30/i0[8] ) );
  CLKBUF_X2 U2536 ( .I(\SB3_0/buf_output[3] ), .Z(\SB4_30/i0[10] ) );
  NAND3_X1 U2539 ( .A1(\SB3_21/i0_3 ), .A2(\SB3_21/i0_4 ), .A3(\SB3_21/i1[9] ), 
        .ZN(n6820) );
  BUF_X4 U2540 ( .I(\MC_ARK_ARC_1_4/buf_output[65] ), .Z(\SB3_21/i0_3 ) );
  BUF_X2 U2541 ( .I(\MC_ARK_ARC_1_4/buf_output[21] ), .Z(\SB3_28/i0[10] ) );
  INV_X1 U2544 ( .I(\MC_ARK_ARC_1_4/buf_output[21] ), .ZN(\SB3_28/i0[8] ) );
  NAND3_X1 U2545 ( .A1(\RI1[4][17] ), .A2(\SB1_4_29/i1[9] ), .A3(
        \SB1_4_29/i0[6] ), .ZN(\SB1_4_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2549 ( .A1(\RI1[4][17] ), .A2(\SB1_4_29/i0[10] ), .A3(
        \SB1_4_29/i0[6] ), .ZN(\SB1_4_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2550 ( .A1(\SB1_4_29/i0[10] ), .A2(\SB1_4_29/i0[9] ), .A3(
        \RI1[4][17] ), .ZN(n7527) );
  NAND3_X1 U2551 ( .A1(\SB1_4_29/i0_4 ), .A2(\RI1[4][17] ), .A3(
        \SB1_4_29/i1[9] ), .ZN(n6682) );
  NAND3_X1 U2552 ( .A1(\SB1_4_29/i0[8] ), .A2(\SB1_4_29/i0[9] ), .A3(
        \RI1[4][17] ), .ZN(n4156) );
  NAND3_X1 U2557 ( .A1(\SB1_4_29/i0[8] ), .A2(\RI1[4][17] ), .A3(
        \SB1_4_29/i1_7 ), .ZN(n5826) );
  NAND3_X1 U2558 ( .A1(\RI1[4][17] ), .A2(\SB1_4_29/i0[7] ), .A3(
        \SB1_4_29/i0_0 ), .ZN(n2787) );
  NAND3_X1 U2559 ( .A1(\SB1_4_29/i0_0 ), .A2(\RI1[4][17] ), .A3(
        \SB1_4_29/i0_4 ), .ZN(\SB1_4_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2565 ( .A1(\SB4_22/i0[6] ), .A2(\SB4_22/i0_4 ), .A3(\SB4_22/i0[9] ), .ZN(n5961) );
  CLKBUF_X4 U2566 ( .I(\MC_ARK_ARC_1_4/buf_output[88] ), .Z(\SB3_17/i0_4 ) );
  INV_X1 U2567 ( .I(\MC_ARK_ARC_1_4/buf_output[1] ), .ZN(\SB3_31/i1_7 ) );
  BUF_X2 U2569 ( .I(\MC_ARK_ARC_1_4/buf_output[1] ), .Z(\SB3_31/i0[6] ) );
  NAND3_X1 U2571 ( .A1(\SB4_19/i0_3 ), .A2(\SB4_19/i0[8] ), .A3(\SB4_19/i0[9] ), .ZN(\SB4_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2574 ( .A1(\SB1_4_23/i0[9] ), .A2(\SB1_4_23/i0[10] ), .A3(
        \SB1_4_23/i0_3 ), .ZN(\SB1_4_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2580 ( .A1(\SB1_4_23/i0[10] ), .A2(\SB1_4_23/i1_7 ), .A3(
        \SB1_4_23/i1[9] ), .ZN(n3376) );
  NAND3_X1 U2582 ( .A1(\SB1_4_23/i0_0 ), .A2(\SB1_4_23/i0[6] ), .A3(
        \SB1_4_23/i0[10] ), .ZN(\SB1_4_23/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U2592 ( .A1(\SB1_4_23/i1_5 ), .A2(\SB1_4_23/i0[10] ), .A3(
        \SB1_4_23/i1[9] ), .ZN(\SB1_4_23/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U2596 ( .I(\MC_ARK_ARC_1_2/buf_output[170] ), .ZN(\SB1_3_3/i1[9] ) );
  BUF_X2 U2601 ( .I(\MC_ARK_ARC_1_2/buf_output[170] ), .Z(\SB1_3_3/i0_0 ) );
  BUF_X2 U2603 ( .I(\MC_ARK_ARC_1_4/buf_output[163] ), .Z(\SB3_4/i0[6] ) );
  CLKBUF_X4 U2604 ( .I(\SB2_4_22/buf_output[3] ), .Z(\RI5[4][69] ) );
  INV_X1 U2608 ( .I(\MC_ARK_ARC_1_3/buf_output[181] ), .ZN(\SB1_4_1/i1_7 ) );
  BUF_X2 U2609 ( .I(\MC_ARK_ARC_1_3/buf_output[181] ), .Z(\SB1_4_1/i0[6] ) );
  NAND3_X1 U2610 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i1_5 ), .A3(\SB4_10/i0_4 ), 
        .ZN(n6747) );
  NAND3_X1 U2612 ( .A1(\SB3_5/i0_0 ), .A2(\SB3_5/i0[6] ), .A3(\SB3_5/i0[10] ), 
        .ZN(\SB3_5/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X2 U2613 ( .I(\SB3_10/buf_output[0] ), .Z(\SB4_5/i0[9] ) );
  NAND2_X1 U2616 ( .A1(\SB2_4_19/i0_0 ), .A2(\SB2_4_19/i3[0] ), .ZN(
        \SB2_4_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2622 ( .A1(\SB2_4_19/i0[10] ), .A2(\SB2_4_19/i0_0 ), .A3(
        \SB2_4_19/i0[6] ), .ZN(\SB2_4_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2623 ( .A1(\SB2_4_19/i3[0] ), .A2(\SB2_4_19/i0_0 ), .A3(
        \SB2_4_19/i1_7 ), .ZN(\SB2_4_19/Component_Function_4/NAND4_in[1] ) );
  CLKBUF_X2 U2626 ( .I(\SB3_13/buf_output[0] ), .Z(\SB4_8/i0[9] ) );
  NAND2_X1 U2627 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i3[0] ), .ZN(
        \SB4_13/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U2632 ( .I(\SB3_31/buf_output[5] ), .Z(\SB4_31/i0_3 ) );
  NAND3_X1 U2633 ( .A1(\SB2_4_19/i1_5 ), .A2(\SB2_4_19/i0[10] ), .A3(
        \SB2_4_19/i1[9] ), .ZN(\SB2_4_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2644 ( .A1(\SB2_4_19/i0[10] ), .A2(\SB2_4_19/i1_7 ), .A3(
        \SB2_4_19/i1[9] ), .ZN(n7221) );
  NAND3_X1 U2645 ( .A1(\SB2_4_19/i0_4 ), .A2(\SB2_4_19/i1[9] ), .A3(
        \SB2_4_19/i1_5 ), .ZN(n4141) );
  NAND3_X1 U2648 ( .A1(\SB2_4_19/i1[9] ), .A2(\SB2_4_19/i0_3 ), .A3(
        \SB2_4_19/i0[6] ), .ZN(\SB2_4_19/Component_Function_3/NAND4_in[0] ) );
  INV_X1 U2649 ( .I(\MC_ARK_ARC_1_4/buf_output[159] ), .ZN(\SB3_5/i0[8] ) );
  BUF_X2 U2654 ( .I(\MC_ARK_ARC_1_4/buf_output[159] ), .Z(\SB3_5/i0[10] ) );
  NAND3_X1 U2659 ( .A1(\SB1_4_18/i1_7 ), .A2(\SB1_4_18/i0[8] ), .A3(
        \SB1_4_18/i0_4 ), .ZN(\SB1_4_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2660 ( .A1(\SB1_4_18/i0[9] ), .A2(\SB1_4_18/i0_0 ), .A3(
        \SB1_4_18/i0[8] ), .ZN(\SB1_4_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2664 ( .A1(\SB1_4_18/i0[8] ), .A2(\SB1_4_18/i1_5 ), .A3(
        \SB1_4_18/i3[0] ), .ZN(n6904) );
  NAND3_X1 U2666 ( .A1(\SB1_4_18/i0_3 ), .A2(\SB1_4_18/i1_7 ), .A3(
        \SB1_4_18/i0[8] ), .ZN(\SB1_4_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2674 ( .A1(\SB1_4_18/i0_3 ), .A2(\SB1_4_18/i0[9] ), .A3(
        \SB1_4_18/i0[8] ), .ZN(n3306) );
  NAND3_X1 U2675 ( .A1(\SB4_12/i1_5 ), .A2(\SB4_12/i0[6] ), .A3(\SB4_12/i0[9] ), .ZN(\SB4_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2676 ( .A1(\SB4_12/i0_3 ), .A2(\SB4_12/i0[8] ), .A3(\SB4_12/i0[9] ), .ZN(\SB4_12/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U2677 ( .I(\SB3_17/buf_output[0] ), .Z(\SB4_12/i0[9] ) );
  NAND3_X1 U2679 ( .A1(\SB4_8/i0_4 ), .A2(\SB4_8/i0_3 ), .A3(n3996), .ZN(n4858) );
  NAND3_X1 U2680 ( .A1(\SB1_1_31/i0[10] ), .A2(\SB1_1_31/i1[9] ), .A3(
        \SB1_1_31/i1_7 ), .ZN(n2519) );
  NAND3_X1 U2685 ( .A1(\SB1_1_31/i0[10] ), .A2(\SB1_1_31/i1[9] ), .A3(
        \SB1_1_31/i1_5 ), .ZN(\SB1_1_31/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U2686 ( .A1(\SB1_1_31/i0[10] ), .A2(\SB1_1_31/i0[9] ), .ZN(
        \SB1_1_31/Component_Function_0/NAND4_in[0] ) );
  INV_X1 U2687 ( .I(\MC_ARK_ARC_1_4/buf_output[133] ), .ZN(\SB3_9/i1_7 ) );
  BUF_X2 U2688 ( .I(\MC_ARK_ARC_1_4/buf_output[133] ), .Z(\SB3_9/i0[6] ) );
  NAND3_X1 U2689 ( .A1(\SB4_24/i0_4 ), .A2(\SB4_24/i0[6] ), .A3(\SB4_24/i0[9] ), .ZN(n6413) );
  NAND3_X1 U2692 ( .A1(\SB4_24/i0_4 ), .A2(\SB4_24/i1[9] ), .A3(\SB4_24/i1_5 ), 
        .ZN(n997) );
  NAND3_X1 U2694 ( .A1(\SB4_24/i1[9] ), .A2(\SB4_24/i0_4 ), .A3(\SB4_24/i0_3 ), 
        .ZN(\SB4_24/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2696 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i0[6] ), .A3(
        \SB4_22/i0[10] ), .ZN(\SB4_22/Component_Function_5/NAND4_in[1] ) );
  INV_X1 U2699 ( .I(\MC_ARK_ARC_1_1/buf_output[127] ), .ZN(\SB1_2_10/i1_7 ) );
  INV_X1 U2700 ( .I(\MC_ARK_ARC_1_4/buf_output[69] ), .ZN(\SB3_20/i0[8] ) );
  BUF_X2 U2702 ( .I(\MC_ARK_ARC_1_4/buf_output[69] ), .Z(\SB3_20/i0[10] ) );
  NAND3_X1 U2704 ( .A1(\SB3_28/i0[7] ), .A2(\SB3_28/i0_3 ), .A3(\SB3_28/i0_0 ), 
        .ZN(\SB3_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2709 ( .A1(\SB3_28/i1[9] ), .A2(\SB3_28/i0_3 ), .A3(\SB3_28/i0[6] ), .ZN(\SB3_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2710 ( .A1(\SB3_28/i0_3 ), .A2(\SB3_28/i1_7 ), .A3(\SB3_28/i0[8] ), 
        .ZN(\SB3_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2713 ( .A1(\SB3_28/i0_3 ), .A2(\SB3_28/i0[10] ), .A3(
        \SB3_28/i0[6] ), .ZN(\SB3_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2714 ( .A1(\SB3_28/i0_0 ), .A2(\SB3_28/i0_3 ), .A3(\SB3_28/i0_4 ), 
        .ZN(\SB3_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2719 ( .A1(\SB3_28/i0_3 ), .A2(\SB3_28/i1[9] ), .A3(\SB3_28/i0_4 ), 
        .ZN(n5235) );
  NAND3_X1 U2722 ( .A1(\SB3_20/i0[6] ), .A2(\SB3_20/i0[9] ), .A3(\SB3_20/i1_5 ), .ZN(n6491) );
  NAND3_X1 U2723 ( .A1(\SB3_9/i1_5 ), .A2(\SB3_9/i0[8] ), .A3(\SB3_9/i3[0] ), 
        .ZN(\SB3_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2724 ( .A1(\SB3_9/i0[8] ), .A2(\SB3_9/i0[7] ), .A3(\SB3_9/i0[6] ), 
        .ZN(\SB3_9/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2735 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i0_4 ), .A3(n4002), .ZN(
        n3754) );
  NAND3_X1 U2738 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i3[0] ), .A3(\SB4_13/i1_7 ), 
        .ZN(n1216) );
  NAND3_X1 U2739 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i0_3 ), .A3(\SB4_13/i0[7] ), 
        .ZN(n2697) );
  CLKBUF_X4 U2743 ( .I(\SB3_16/buf_output[2] ), .Z(\SB4_13/i0_0 ) );
  NAND3_X1 U2744 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i0[6] ), .A3(
        \SB2_3_4/i1[9] ), .ZN(\SB2_3_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2746 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i0_0 ), .A3(
        \SB2_3_4/i0_4 ), .ZN(n7234) );
  NAND3_X1 U2751 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i0[8] ), .A3(
        \SB2_3_4/i0[9] ), .ZN(\SB2_3_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2753 ( .A1(\SB2_3_4/i0[10] ), .A2(\SB2_3_4/i0_3 ), .A3(
        \SB2_3_4/i0_4 ), .ZN(n6117) );
  NAND3_X1 U2754 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i1[9] ), .A3(
        \SB2_3_4/i0_4 ), .ZN(n5392) );
  CLKBUF_X4 U2758 ( .I(\SB2_4_29/buf_output[2] ), .Z(\RI5[4][32] ) );
  NAND3_X1 U2771 ( .A1(\SB1_4_8/i0_0 ), .A2(\SB1_4_8/i0[6] ), .A3(
        \SB1_4_8/i0[10] ), .ZN(\SB1_4_8/Component_Function_5/NAND4_in[1] ) );
  INV_X1 U2773 ( .I(\MC_ARK_ARC_1_4/buf_output[37] ), .ZN(\SB3_25/i1_7 ) );
  BUF_X2 U2774 ( .I(\MC_ARK_ARC_1_4/buf_output[37] ), .Z(\SB3_25/i0[6] ) );
  CLKBUF_X4 U2775 ( .I(\RI5[4][175] ), .Z(n3165) );
  CLKBUF_X4 U2776 ( .I(\SB3_29/buf_output[4] ), .Z(\SB4_28/i0_4 ) );
  NAND3_X1 U2777 ( .A1(\SB3_24/i0_0 ), .A2(\SB3_24/i0[7] ), .A3(\SB3_24/i0_3 ), 
        .ZN(\SB3_24/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U2785 ( .A1(\SB3_24/i0_0 ), .A2(\SB3_24/i3[0] ), .ZN(
        \SB3_24/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U2786 ( .I(\SB3_11/buf_output[5] ), .Z(\SB4_11/i0_3 ) );
  NAND3_X1 U2788 ( .A1(\SB3_24/i0_0 ), .A2(\SB3_24/i1_5 ), .A3(\SB3_24/i0_4 ), 
        .ZN(\SB3_24/Component_Function_2/NAND4_in[3] ) );
  INV_X1 U2794 ( .I(\MC_ARK_ARC_1_4/buf_output[44] ), .ZN(\SB3_24/i1[9] ) );
  BUF_X2 U2799 ( .I(\MC_ARK_ARC_1_4/buf_output[44] ), .Z(\SB3_24/i0_0 ) );
  INV_X1 U2804 ( .I(\MC_ARK_ARC_1_2/buf_output[114] ), .ZN(\SB1_3_12/i3[0] )
         );
  BUF_X2 U2809 ( .I(\MC_ARK_ARC_1_2/buf_output[114] ), .Z(\SB1_3_12/i0[9] ) );
  INV_X1 U2813 ( .I(\SB1_2_26/buf_output[1] ), .ZN(\SB2_2_22/i1_7 ) );
  BUF_X2 U2814 ( .I(\SB1_2_26/buf_output[1] ), .Z(\SB2_2_22/i0[6] ) );
  INV_X1 U2816 ( .I(\SB1_1_31/buf_output[3] ), .ZN(\SB2_1_29/i0[8] ) );
  BUF_X2 U2820 ( .I(\SB1_1_31/buf_output[3] ), .Z(\SB2_1_29/i0[10] ) );
  NAND3_X1 U2822 ( .A1(\SB4_23/i0[6] ), .A2(\SB4_23/i0_4 ), .A3(\SB4_23/i0[9] ), .ZN(n649) );
  NAND3_X1 U2824 ( .A1(\SB4_23/i0[6] ), .A2(\SB4_23/i0[10] ), .A3(
        \SB4_23/i0_3 ), .ZN(n2129) );
  NAND3_X1 U2826 ( .A1(\SB4_23/i0[6] ), .A2(\SB4_23/i0_3 ), .A3(\SB4_23/i1[9] ), .ZN(n2141) );
  CLKBUF_X2 U2831 ( .I(\SB3_27/buf_output[1] ), .Z(\SB4_23/i0[6] ) );
  NAND3_X1 U2833 ( .A1(\SB2_4_23/i0_3 ), .A2(\SB2_4_23/i0[10] ), .A3(
        \SB2_4_23/i0[6] ), .ZN(\SB2_4_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2836 ( .A1(\SB2_4_23/i0[10] ), .A2(\SB2_4_23/i0_0 ), .A3(
        \SB2_4_23/i0[6] ), .ZN(\SB2_4_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2837 ( .A1(\SB2_4_23/i0[10] ), .A2(\SB2_4_23/i1_7 ), .A3(
        \SB2_4_23/i1[9] ), .ZN(\SB2_4_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2838 ( .A1(\SB3_15/i0_0 ), .A2(\SB3_15/i0_4 ), .A3(\SB3_15/i1_5 ), 
        .ZN(n6863) );
  NAND3_X1 U2841 ( .A1(\SB3_15/i0_0 ), .A2(\SB3_15/i0[10] ), .A3(
        \SB3_15/i0[6] ), .ZN(n6943) );
  NAND3_X1 U2843 ( .A1(\SB3_15/i0_0 ), .A2(\SB3_15/i0_3 ), .A3(\SB3_15/i0[7] ), 
        .ZN(n6063) );
  NAND2_X1 U2844 ( .A1(\SB3_15/i3[0] ), .A2(\SB3_15/i0_0 ), .ZN(n3476) );
  BUF_X2 U2845 ( .I(\SB3_0/buf_output[0] ), .Z(\SB4_27/i0[9] ) );
  NAND3_X1 U2847 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i0_4 ), .A3(
        \SB2_3_23/i0[10] ), .ZN(n4485) );
  NAND3_X1 U2849 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i0[8] ), .A3(
        \SB2_3_23/i0[9] ), .ZN(\SB2_3_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2850 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i0[10] ), .A3(
        \SB2_3_23/i0[6] ), .ZN(n6510) );
  NAND3_X1 U2852 ( .A1(\SB2_3_23/i0_0 ), .A2(\SB2_3_23/i0_3 ), .A3(
        \SB2_3_23/i0[7] ), .ZN(n6983) );
  NAND3_X1 U2855 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i1[9] ), .A3(
        \SB2_3_23/i0[6] ), .ZN(n4476) );
  NAND3_X1 U2856 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i0_4 ), .A3(
        \SB1_2_18/i1_5 ), .ZN(n1817) );
  NAND3_X1 U2857 ( .A1(\SB1_2_18/i0[8] ), .A2(\SB1_2_18/i1_5 ), .A3(
        \SB1_2_18/i3[0] ), .ZN(n7455) );
  INV_X1 U2860 ( .I(\MC_ARK_ARC_1_1/buf_output[85] ), .ZN(\SB1_2_17/i1_7 ) );
  INV_X1 U2862 ( .I(\MC_ARK_ARC_1_4/buf_output[98] ), .ZN(\SB3_15/i1[9] ) );
  BUF_X2 U2864 ( .I(\MC_ARK_ARC_1_4/buf_output[98] ), .Z(\SB3_15/i0_0 ) );
  INV_X1 U2865 ( .I(\MC_ARK_ARC_1_4/buf_output[150] ), .ZN(\SB3_6/i3[0] ) );
  BUF_X2 U2874 ( .I(\MC_ARK_ARC_1_4/buf_output[150] ), .Z(\SB3_6/i0[9] ) );
  NAND3_X1 U2880 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i0[10] ), .A3(
        \SB2_1_26/i0_4 ), .ZN(n2046) );
  NAND3_X1 U2886 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i1_7 ), .A3(
        \SB2_1_26/i0[8] ), .ZN(\SB2_1_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2887 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i1[9] ), .A3(
        \SB2_1_26/i0_4 ), .ZN(\SB2_1_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2891 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i0[10] ), .A3(
        \SB2_1_26/i0[6] ), .ZN(\SB2_1_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2896 ( .A1(\SB2_1_26/i1[9] ), .A2(\SB2_1_26/i0_3 ), .A3(
        \SB2_1_26/i0[6] ), .ZN(\SB2_1_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2897 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i0_0 ), .A3(
        \SB2_1_26/i0_4 ), .ZN(\SB2_1_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2903 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i0[9] ), .A3(
        \SB2_1_26/i0[10] ), .ZN(n2047) );
  NAND2_X1 U2904 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i1[9] ), .ZN(
        \SB2_1_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2905 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i0_0 ), .A3(
        \SB2_1_26/i0[7] ), .ZN(n5496) );
  CLKBUF_X4 U2908 ( .I(\SB2_1_26/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[50] ) );
  NAND2_X1 U2913 ( .A1(\SB1_2_22/i0[8] ), .A2(n7143), .ZN(n4565) );
  NAND3_X1 U2914 ( .A1(\SB1_4_8/i0[9] ), .A2(\SB1_4_8/i0_3 ), .A3(
        \SB1_4_8/i0[8] ), .ZN(n7204) );
  NAND3_X1 U2919 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i0[6] ), .A3(
        \SB4_30/i0_3 ), .ZN(n5598) );
  OR3_X1 U2929 ( .A1(\MC_ARK_ARC_1_3/buf_output[138] ), .A2(
        \MC_ARK_ARC_1_3/buf_output[143] ), .A3(\RI1[4][141] ), .Z(n3013) );
  INV_X1 U2933 ( .I(\MC_ARK_ARC_1_4/buf_output[152] ), .ZN(\SB3_6/i1[9] ) );
  BUF_X2 U2935 ( .I(\MC_ARK_ARC_1_4/buf_output[152] ), .Z(\SB3_6/i0_0 ) );
  INV_X1 U2940 ( .I(\MC_ARK_ARC_1_4/buf_output[187] ), .ZN(\SB3_0/i1_7 ) );
  BUF_X2 U2941 ( .I(\MC_ARK_ARC_1_4/buf_output[187] ), .Z(\SB3_0/i0[6] ) );
  INV_X1 U2942 ( .I(\SB3_7/buf_output[2] ), .ZN(\SB4_4/i1[9] ) );
  BUF_X2 U2943 ( .I(\SB3_7/buf_output[2] ), .Z(\SB4_4/i0_0 ) );
  NAND3_X1 U2945 ( .A1(\SB4_8/i0[9] ), .A2(\SB4_8/i0_0 ), .A3(\SB4_8/i0[8] ), 
        .ZN(\SB4_8/Component_Function_4/NAND4_in[0] ) );
  BUF_X2 U2946 ( .I(\RI3[2][97] ), .Z(\SB2_2_15/i0[6] ) );
  INV_X1 U2949 ( .I(\RI3[2][97] ), .ZN(\SB2_2_15/i1_7 ) );
  INV_X1 U2951 ( .I(\SB3_17/buf_output[2] ), .ZN(\SB4_14/i1[9] ) );
  BUF_X2 U2952 ( .I(\SB3_17/buf_output[2] ), .Z(\SB4_14/i0_0 ) );
  BUF_X2 U2955 ( .I(\MC_ARK_ARC_1_1/buf_output[55] ), .Z(\SB1_2_22/i0[6] ) );
  INV_X1 U2960 ( .I(\MC_ARK_ARC_1_1/buf_output[55] ), .ZN(\SB1_2_22/i1_7 ) );
  INV_X1 U2962 ( .I(\MC_ARK_ARC_1_3/buf_output[42] ), .ZN(\SB1_4_24/i3[0] ) );
  BUF_X2 U2963 ( .I(\MC_ARK_ARC_1_3/buf_output[42] ), .Z(\SB1_4_24/i0[9] ) );
  INV_X1 U2964 ( .I(\SB3_20/buf_output[3] ), .ZN(\SB4_18/i0[8] ) );
  BUF_X2 U2966 ( .I(\SB3_20/buf_output[3] ), .Z(\SB4_18/i0[10] ) );
  INV_X1 U2968 ( .I(\MC_ARK_ARC_1_3/buf_output[158] ), .ZN(\SB1_4_5/i1[9] ) );
  BUF_X2 U2969 ( .I(\MC_ARK_ARC_1_3/buf_output[158] ), .Z(\SB1_4_5/i0_0 ) );
  CLKBUF_X2 U2972 ( .I(Key[83]), .Z(n86) );
  NAND2_X1 U2977 ( .A1(\SB4_8/i0[9] ), .A2(\SB4_8/i0[10] ), .ZN(n903) );
  CLKBUF_X4 U2983 ( .I(\SB3_8/buf_output[5] ), .Z(\SB4_8/i0_3 ) );
  CLKBUF_X4 U2984 ( .I(\SB1_3_25/buf_output[5] ), .Z(\SB2_3_25/i0_3 ) );
  NAND3_X1 U2986 ( .A1(\SB1_4_28/i0_3 ), .A2(\SB1_4_28/i0[8] ), .A3(
        \SB1_4_28/i0[9] ), .ZN(\SB1_4_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2990 ( .A1(\SB1_4_28/i1_5 ), .A2(\SB1_4_28/i0[8] ), .A3(
        \SB1_4_28/i3[0] ), .ZN(n3255) );
  INV_X1 U2991 ( .I(\RI3[5][128] ), .ZN(\SB4_10/i1[9] ) );
  BUF_X2 U2994 ( .I(\RI3[5][128] ), .Z(\SB4_10/i0_0 ) );
  NAND3_X1 U2998 ( .A1(\SB1_4_11/i0_3 ), .A2(\SB1_4_11/i1[9] ), .A3(
        \SB1_4_11/i0_4 ), .ZN(n5068) );
  NAND3_X1 U2999 ( .A1(\SB1_4_11/i0[7] ), .A2(\SB1_4_11/i0_3 ), .A3(
        \SB1_4_11/i0_0 ), .ZN(\SB1_4_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3000 ( .A1(\SB1_4_11/i0[9] ), .A2(\SB1_4_11/i0_3 ), .A3(
        \SB1_4_11/i0[10] ), .ZN(\SB1_4_11/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U3001 ( .A1(\SB1_4_11/i0_3 ), .A2(\SB1_4_11/i0[10] ), .A3(
        \SB1_4_11/i0[6] ), .ZN(\SB1_4_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3002 ( .A1(\SB1_4_11/i0_3 ), .A2(\SB1_4_11/i0[8] ), .A3(
        \SB1_4_11/i0[9] ), .ZN(\SB1_4_11/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 U3003 ( .A1(\SB1_4_11/i0_3 ), .A2(\SB1_4_11/i1[9] ), .ZN(
        \SB1_4_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3004 ( .A1(\SB1_4_11/i1[9] ), .A2(\SB1_4_11/i0_3 ), .A3(
        \SB1_4_11/i0[6] ), .ZN(\SB1_4_11/Component_Function_3/NAND4_in[0] ) );
  INV_X1 U3005 ( .I(\MC_ARK_ARC_1_4/buf_output[45] ), .ZN(\SB3_24/i0[8] ) );
  BUF_X2 U3007 ( .I(\MC_ARK_ARC_1_4/buf_output[45] ), .Z(\SB3_24/i0[10] ) );
  NAND3_X1 U3008 ( .A1(\SB1_4_14/i0_0 ), .A2(\SB1_4_14/i1_7 ), .A3(
        \SB1_4_14/i3[0] ), .ZN(\SB1_4_14/Component_Function_4/NAND4_in[1] ) );
  BUF_X2 U3013 ( .I(\SB1_0_13/buf_output[0] ), .Z(\SB2_0_8/i0[9] ) );
  NAND3_X1 U3015 ( .A1(\SB1_4_19/i0[6] ), .A2(\SB1_4_19/i0_3 ), .A3(
        \SB1_4_19/i0[10] ), .ZN(\SB1_4_19/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X1 U3016 ( .A1(\SB1_4_19/i0[9] ), .A2(\SB1_4_19/i0[10] ), .A3(
        \SB1_4_19/i0_3 ), .ZN(\SB1_4_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3021 ( .A1(\SB1_4_19/i0[10] ), .A2(\SB1_4_19/i0_4 ), .A3(
        \SB1_4_19/i0_3 ), .ZN(\SB1_4_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3022 ( .A1(\SB1_4_19/i0_3 ), .A2(\SB1_4_19/i1_7 ), .A3(
        \SB1_4_19/i0[8] ), .ZN(\SB1_4_19/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X4 U3025 ( .I(\SB1_3_21/buf_output[5] ), .Z(\SB2_3_21/i0_3 ) );
  BUF_X2 U3026 ( .I(\MC_ARK_ARC_1_2/buf_output[91] ), .Z(\SB1_3_16/i0[6] ) );
  INV_X1 U3027 ( .I(\MC_ARK_ARC_1_2/buf_output[91] ), .ZN(\SB1_3_16/i1_7 ) );
  CLKBUF_X4 U3034 ( .I(\SB2_1_31/i0_4 ), .Z(n5429) );
  AND2_X1 U3035 ( .A1(\SB1_1_0/Component_Function_4/NAND4_in[2] ), .A2(n3591), 
        .Z(n5426) );
  NAND3_X1 U3036 ( .A1(\SB3_9/i1[9] ), .A2(\SB3_9/i0[10] ), .A3(\SB3_9/i1_5 ), 
        .ZN(n5608) );
  NAND3_X1 U3037 ( .A1(\SB3_9/i1[9] ), .A2(\SB3_9/i1_7 ), .A3(\SB3_9/i0[10] ), 
        .ZN(\SB3_9/Component_Function_3/NAND4_in[2] ) );
  INV_X1 U3039 ( .I(\MC_ARK_ARC_1_2/buf_output[181] ), .ZN(\SB1_3_1/i1_7 ) );
  INV_X1 U3041 ( .I(\MC_ARK_ARC_1_2/buf_output[55] ), .ZN(\SB1_3_22/i1_7 ) );
  CLKBUF_X4 U3056 ( .I(n354), .Z(\SB1_0_13/i0_4 ) );
  INV_X1 U3058 ( .I(\MC_ARK_ARC_1_3/buf_output[36] ), .ZN(\SB1_4_25/i3[0] ) );
  CLKBUF_X4 U3061 ( .I(\SB1_2_22/buf_output[3] ), .Z(\SB2_2_20/i0[10] ) );
  NAND3_X1 U3062 ( .A1(\SB1_2_4/i1_5 ), .A2(\SB1_2_4/i0[6] ), .A3(
        \SB1_2_4/i0[9] ), .ZN(\SB1_2_4/Component_Function_1/NAND4_in[2] ) );
  INV_X1 U3064 ( .I(\MC_ARK_ARC_1_1/buf_output[71] ), .ZN(\SB1_2_20/i1_5 ) );
  INV_X1 U3065 ( .I(\SB1_3_10/buf_output[5] ), .ZN(\SB2_3_10/i1_5 ) );
  BUF_X2 U3067 ( .I(\SB1_2_13/buf_output[1] ), .Z(\SB2_2_9/i0[6] ) );
  INV_X1 U3071 ( .I(\SB1_2_13/buf_output[1] ), .ZN(\SB2_2_9/i1_7 ) );
  NAND3_X1 U3075 ( .A1(\SB2_3_29/i0_0 ), .A2(\SB2_3_29/i0_4 ), .A3(
        \SB2_3_29/i1_5 ), .ZN(n1876) );
  INV_X1 U3077 ( .I(\MC_ARK_ARC_1_3/buf_output[73] ), .ZN(\SB1_4_19/i1_7 ) );
  BUF_X2 U3078 ( .I(\MC_ARK_ARC_1_3/buf_output[73] ), .Z(\SB1_4_19/i0[6] ) );
  INV_X1 U3081 ( .I(\MC_ARK_ARC_1_3/buf_output[102] ), .ZN(\SB1_4_14/i3[0] )
         );
  BUF_X2 U3082 ( .I(\MC_ARK_ARC_1_0/buf_output[102] ), .Z(\SB1_1_14/i0[9] ) );
  CLKBUF_X4 U3084 ( .I(\SB1_2_15/buf_output[2] ), .Z(\SB2_2_12/i0_0 ) );
  CLKBUF_X4 U3086 ( .I(\SB2_2_2/buf_output[3] ), .Z(\RI5[2][189] ) );
  INV_X1 U3089 ( .I(\SB1_2_29/buf_output[1] ), .ZN(\SB2_2_25/i1_7 ) );
  INV_X1 U3095 ( .I(\SB1_4_19/buf_output[0] ), .ZN(\SB2_4_14/i3[0] ) );
  BUF_X2 U3097 ( .I(\SB1_4_19/buf_output[0] ), .Z(\SB2_4_14/i0[9] ) );
  INV_X1 U3100 ( .I(\MC_ARK_ARC_1_2/buf_output[18] ), .ZN(\SB1_3_28/i3[0] ) );
  NAND3_X1 U3102 ( .A1(n1495), .A2(\SB4_14/i0[8] ), .A3(\SB4_14/i3[0] ), .ZN(
        \SB4_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3108 ( .A1(\SB1_3_3/i0_4 ), .A2(\SB1_3_3/i1[9] ), .A3(
        \SB1_3_3/i1_5 ), .ZN(n5811) );
  NAND3_X1 U3109 ( .A1(\SB1_3_3/i0[10] ), .A2(\SB1_3_3/i1[9] ), .A3(
        \SB1_3_3/i1_7 ), .ZN(\SB1_3_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3112 ( .A1(\SB1_3_3/i0_3 ), .A2(\SB1_3_3/i1[9] ), .A3(
        \SB1_3_3/i0_4 ), .ZN(\SB1_3_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3114 ( .A1(\SB1_3_3/i0[10] ), .A2(\SB1_3_3/i1[9] ), .A3(
        \SB1_3_3/i1_5 ), .ZN(n6541) );
  NAND3_X1 U3117 ( .A1(\SB2_3_11/i0_3 ), .A2(\SB2_3_11/i0[8] ), .A3(
        \SB2_3_11/i0[9] ), .ZN(\SB2_3_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3118 ( .A1(\SB1_3_1/i0_3 ), .A2(\SB1_3_1/i0[8] ), .A3(
        \SB1_3_1/i1_7 ), .ZN(\SB1_3_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3119 ( .A1(\SB1_3_1/i0_0 ), .A2(\SB1_3_1/i0_3 ), .A3(
        \SB1_3_1/i0_4 ), .ZN(\SB1_3_1/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 U3125 ( .I(\SB2_1_11/buf_output[3] ), .Z(\RI5[1][135] ) );
  NAND2_X1 U3126 ( .A1(\SB2_0_14/i3[0] ), .A2(\SB2_0_14/i0_0 ), .ZN(
        \SB2_0_14/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U3128 ( .I(\MC_ARK_ARC_1_1/buf_output[90] ), .ZN(\SB1_2_16/i3[0] ) );
  NAND3_X1 U3132 ( .A1(n5431), .A2(\SB1_3_15/i1_7 ), .A3(\SB1_3_15/i0[10] ), 
        .ZN(\SB1_3_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3133 ( .A1(\SB1_3_15/i0_3 ), .A2(\SB1_3_15/i0[10] ), .A3(
        \SB1_3_15/i0[6] ), .ZN(\SB1_3_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3134 ( .A1(\SB1_3_15/i0[10] ), .A2(\SB1_3_15/i0_4 ), .A3(
        \SB1_3_15/i0_3 ), .ZN(\SB1_3_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3135 ( .A1(\SB1_3_15/i0[9] ), .A2(\SB1_3_15/i0[10] ), .A3(
        \SB1_3_15/i0_3 ), .ZN(\SB1_3_15/Component_Function_4/NAND4_in[2] ) );
  CLKBUF_X4 U3138 ( .I(\SB1_2_31/buf_output[3] ), .Z(\SB2_2_29/i0[10] ) );
  BUF_X4 U3139 ( .I(\MC_ARK_ARC_1_3/buf_output[15] ), .Z(\SB1_4_29/i0[10] ) );
  CLKBUF_X4 U3140 ( .I(\SB2_0_14/buf_output[3] ), .Z(\RI5[0][117] ) );
  INV_X1 U3141 ( .I(\MC_ARK_ARC_1_1/buf_output[95] ), .ZN(\SB1_2_16/i1_5 ) );
  INV_X1 U3142 ( .I(n345), .ZN(\SB1_0_17/i0[8] ) );
  BUF_X2 U3143 ( .I(n345), .Z(\SB1_0_17/i0[10] ) );
  BUF_X2 U3147 ( .I(n352), .Z(\SB1_0_14/i0_4 ) );
  CLKBUF_X4 U3151 ( .I(\SB1_2_10/buf_output[3] ), .Z(\SB2_2_8/i0[10] ) );
  NAND3_X1 U3152 ( .A1(\SB1_1_26/i1[9] ), .A2(\SB1_1_26/i0_4 ), .A3(
        \SB1_1_26/i0_3 ), .ZN(\SB1_1_26/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U3160 ( .I(\RI1[1][179] ), .ZN(\SB1_1_2/i1_5 ) );
  NAND3_X1 U3161 ( .A1(\SB4_4/i1_5 ), .A2(\SB4_4/i0[8] ), .A3(\SB4_4/i3[0] ), 
        .ZN(\SB4_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3162 ( .A1(\SB4_4/i0[10] ), .A2(\SB4_4/i1_5 ), .A3(\SB4_4/i1[9] ), 
        .ZN(n6188) );
  BUF_X2 U3164 ( .I(\MC_ARK_ARC_1_4/buf_output[49] ), .Z(\SB3_23/i0[6] ) );
  BUF_X4 U3168 ( .I(\SB1_1_23/buf_output[2] ), .Z(\SB2_1_20/i0_0 ) );
  NAND3_X1 U3170 ( .A1(\SB2_3_4/i0_0 ), .A2(\SB2_3_4/i0_3 ), .A3(n5683), .ZN(
        n6116) );
  NAND3_X1 U3171 ( .A1(\SB2_3_4/i0_0 ), .A2(\SB2_3_4/i0_4 ), .A3(
        \SB2_3_4/i1_5 ), .ZN(n1875) );
  NAND2_X1 U3172 ( .A1(\SB2_1_3/i0_3 ), .A2(\SB2_1_3/i1[9] ), .ZN(
        \SB2_1_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3179 ( .A1(\SB2_1_2/i0[10] ), .A2(\SB2_1_2/i0_3 ), .A3(
        \SB2_1_2/i0[9] ), .ZN(n2427) );
  NAND3_X1 U3180 ( .A1(\SB2_1_2/i0[10] ), .A2(\SB2_1_2/i0[6] ), .A3(
        \SB2_1_2/i0_3 ), .ZN(n3452) );
  BUF_X4 U3181 ( .I(\MC_ARK_ARC_1_1/buf_output[172] ), .Z(\SB1_2_3/i0_4 ) );
  CLKBUF_X4 U3192 ( .I(\MC_ARK_ARC_1_1/buf_output[164] ), .Z(\SB1_2_4/i0_0 )
         );
  INV_X1 U3204 ( .I(\SB1_4_16/buf_output[1] ), .ZN(\SB2_4_12/i1_7 ) );
  OR3_X2 U3205 ( .A1(\RI3[0][77] ), .A2(\SB1_0_21/buf_output[3] ), .A3(
        \RI3[0][72] ), .Z(\SB2_0_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3207 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i0[6] ), .A3(
        \SB2_1_25/i1[9] ), .ZN(\SB2_1_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3208 ( .A1(\SB2_1_25/i0[9] ), .A2(\SB2_1_25/i0_3 ), .A3(n3995), 
        .ZN(n4622) );
  CLKBUF_X4 U3217 ( .I(\MC_ARK_ARC_1_3/buf_output[116] ), .Z(\SB1_4_12/i0_0 )
         );
  INV_X1 U3223 ( .I(\MC_ARK_ARC_1_4/buf_output[19] ), .ZN(\SB3_28/i1_7 ) );
  NAND3_X1 U3225 ( .A1(\SB1_1_17/i0_3 ), .A2(\SB1_1_17/i0[8] ), .A3(
        \SB1_1_17/i1_7 ), .ZN(\SB1_1_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U3229 ( .A1(\SB1_1_17/i0_3 ), .A2(\SB1_1_17/i1[9] ), .ZN(
        \SB1_1_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3236 ( .A1(\SB1_1_17/i0[7] ), .A2(\SB1_1_17/i0_3 ), .A3(
        \SB1_1_17/i0_0 ), .ZN(\SB1_1_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3245 ( .A1(\SB1_1_17/i0_0 ), .A2(\SB1_1_17/i0_3 ), .A3(
        \SB1_1_17/i0_4 ), .ZN(\SB1_1_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3255 ( .A1(\SB1_1_17/i0_3 ), .A2(\SB1_1_17/i1[9] ), .A3(
        \SB1_1_17/i0[6] ), .ZN(n1723) );
  INV_X1 U3258 ( .I(\SB1_2_9/buf_output[1] ), .ZN(\SB2_2_5/i1_7 ) );
  CLKBUF_X4 U3260 ( .I(\SB2_3_0/buf_output[3] ), .Z(\RI5[3][9] ) );
  INV_X1 U3261 ( .I(\MC_ARK_ARC_1_4/buf_output[191] ), .ZN(\SB3_0/i1_5 ) );
  CLKBUF_X4 U3263 ( .I(\MC_ARK_ARC_1_4/buf_output[191] ), .Z(\SB3_0/i0_3 ) );
  INV_X1 U3266 ( .I(\MC_ARK_ARC_1_3/buf_output[115] ), .ZN(\SB1_4_12/i1_7 ) );
  BUF_X4 U3267 ( .I(\SB2_2_25/buf_output[3] ), .Z(\RI5[2][51] ) );
  NAND3_X1 U3268 ( .A1(\SB1_0_25/i1[9] ), .A2(\SB1_0_25/i0_3 ), .A3(
        \SB1_0_25/i0[6] ), .ZN(\SB1_0_25/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U3270 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i1[9] ), .ZN(
        \SB1_0_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3271 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0[10] ), .A3(
        \SB1_0_25/i0[9] ), .ZN(n6616) );
  NAND3_X1 U3274 ( .A1(\SB1_0_25/i0[10] ), .A2(\SB1_0_25/i0_3 ), .A3(
        \SB1_0_25/i0_4 ), .ZN(n5270) );
  NAND3_X1 U3280 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0_0 ), .A3(
        \SB1_0_25/i0[7] ), .ZN(n5269) );
  NAND3_X1 U3287 ( .A1(\SB2_1_13/i0[7] ), .A2(\SB2_1_13/i0_3 ), .A3(
        \SB2_1_13/i0_0 ), .ZN(\SB2_1_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3288 ( .A1(\SB2_1_13/i0_3 ), .A2(\SB2_1_13/i0[10] ), .A3(
        \SB2_1_13/i0_4 ), .ZN(\SB2_1_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3289 ( .A1(\SB2_1_13/i0[6] ), .A2(\SB2_1_13/i0_3 ), .A3(
        \SB2_1_13/i1[9] ), .ZN(n6966) );
  NAND3_X1 U3296 ( .A1(\SB2_1_13/i0[6] ), .A2(\SB2_1_13/i0_3 ), .A3(
        \SB2_1_13/i0[10] ), .ZN(n7267) );
  NAND3_X1 U3299 ( .A1(\SB2_1_13/i0_4 ), .A2(\SB2_1_13/i1[9] ), .A3(
        \SB2_1_13/i0_3 ), .ZN(n2570) );
  NAND3_X1 U3301 ( .A1(\SB2_1_13/i0_0 ), .A2(\SB2_1_13/i0_3 ), .A3(n2156), 
        .ZN(\SB2_1_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3302 ( .A1(\SB2_1_13/i0_3 ), .A2(\SB2_1_13/i0[10] ), .A3(
        \SB2_1_13/i0[9] ), .ZN(n6677) );
  CLKBUF_X4 U3305 ( .I(\SB4_30/i0_0 ), .Z(n5427) );
  NAND3_X2 U3307 ( .A1(\SB1_4_26/i0[10] ), .A2(\SB1_4_26/i1[9] ), .A3(
        \SB1_4_26/i1_7 ), .ZN(n1795) );
  BUF_X4 U3308 ( .I(\SB2_4_14/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[117] ) );
  NAND3_X1 U3309 ( .A1(\SB2_2_15/i0[10] ), .A2(\SB2_2_15/i1_5 ), .A3(
        \SB2_2_15/i1[9] ), .ZN(\SB2_2_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3315 ( .A1(\SB2_2_21/i0_3 ), .A2(\SB2_2_21/i1_7 ), .A3(
        \SB2_2_21/i0[8] ), .ZN(\SB2_2_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U3316 ( .A1(\SB2_2_21/i0_3 ), .A2(\SB2_2_21/i1[9] ), .ZN(
        \SB2_2_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3322 ( .A1(\SB2_2_21/i0[9] ), .A2(\SB2_2_21/i0_3 ), .A3(
        \SB2_2_21/i0[8] ), .ZN(n1052) );
  NAND3_X1 U3323 ( .A1(\SB2_2_21/i0[9] ), .A2(\SB2_2_21/i0_3 ), .A3(
        \SB2_2_21/i0[10] ), .ZN(n6040) );
  NAND3_X1 U3324 ( .A1(\SB2_2_21/i0_0 ), .A2(n7225), .A3(\SB2_2_21/i0_3 ), 
        .ZN(n4473) );
  NAND3_X1 U3328 ( .A1(\SB2_2_21/i0_0 ), .A2(\SB2_2_21/i0_3 ), .A3(
        \SB1_2_22/buf_output[4] ), .ZN(
        \SB2_2_21/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U3329 ( .I(\MC_ARK_ARC_1_1/buf_output[179] ), .ZN(\SB1_2_2/i1_5 ) );
  CLKBUF_X4 U3331 ( .I(\MC_ARK_ARC_1_1/buf_output[179] ), .Z(\SB1_2_2/i0_3 )
         );
  NAND3_X1 U3332 ( .A1(\SB1_4_30/i0_4 ), .A2(\SB1_4_30/i1[9] ), .A3(n3993), 
        .ZN(\SB1_4_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3334 ( .A1(\SB1_3_0/i0[8] ), .A2(\SB1_3_0/i1_5 ), .A3(
        \SB1_3_0/i3[0] ), .ZN(n6538) );
  BUF_X4 U3336 ( .I(n339), .Z(\SB1_0_20/i0[10] ) );
  INV_X1 U3349 ( .I(\SB1_4_25/buf_output[1] ), .ZN(\SB2_4_21/i1_7 ) );
  INV_X1 U3350 ( .I(\SB1_4_13/buf_output[5] ), .ZN(\SB2_4_13/i1_5 ) );
  NAND3_X1 U3357 ( .A1(\SB1_1_17/i1_7 ), .A2(\SB1_1_17/i0[8] ), .A3(
        \SB1_1_17/i0_4 ), .ZN(\SB1_1_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3360 ( .A1(\SB1_1_17/i3[0] ), .A2(\SB1_1_17/i0[8] ), .A3(
        \SB1_1_17/i1_5 ), .ZN(n6703) );
  INV_X1 U3363 ( .I(\RI1[3][191] ), .ZN(\SB1_3_0/i1_5 ) );
  CLKBUF_X4 U3365 ( .I(\RI1[3][191] ), .Z(\SB1_3_0/i0_3 ) );
  BUF_X4 U3368 ( .I(\MC_ARK_ARC_1_3/buf_output[182] ), .Z(\SB1_4_1/i0_0 ) );
  INV_X1 U3369 ( .I(\MC_ARK_ARC_1_1/buf_output[61] ), .ZN(\SB1_2_21/i1_7 ) );
  NAND2_X1 U3370 ( .A1(\SB1_4_26/i0_3 ), .A2(\SB1_4_26/i1[9] ), .ZN(
        \SB1_4_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3371 ( .A1(\SB1_4_26/i1[9] ), .A2(\SB1_4_26/i0_3 ), .A3(
        \SB1_4_26/i0[6] ), .ZN(\SB1_4_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3372 ( .A1(\SB1_4_26/i1[9] ), .A2(\SB1_4_26/i0_4 ), .A3(
        \SB1_4_26/i0_3 ), .ZN(\SB1_4_26/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U3373 ( .I(\MC_ARK_ARC_1_0/buf_output[114] ), .ZN(\SB1_1_12/i3[0] )
         );
  BUF_X2 U3374 ( .I(\MC_ARK_ARC_1_1/buf_output[121] ), .Z(\SB1_2_11/i0[6] ) );
  INV_X1 U3375 ( .I(\MC_ARK_ARC_1_1/buf_output[121] ), .ZN(\SB1_2_11/i1_7 ) );
  INV_X1 U3377 ( .I(\SB1_2_13/buf_output[5] ), .ZN(\SB2_2_13/i1_5 ) );
  CLKBUF_X4 U3378 ( .I(\SB1_2_13/buf_output[5] ), .Z(\SB2_2_13/i0_3 ) );
  NAND3_X1 U3379 ( .A1(\SB3_16/i1[9] ), .A2(\SB3_16/i0_3 ), .A3(\SB3_16/i0[6] ), .ZN(\SB3_16/Component_Function_3/NAND4_in[0] ) );
  INV_X1 U3391 ( .I(\MC_ARK_ARC_1_1/buf_output[123] ), .ZN(\SB1_2_11/i0[8] )
         );
  BUF_X2 U3392 ( .I(\MC_ARK_ARC_1_1/buf_output[123] ), .Z(\SB1_2_11/i0[10] )
         );
  CLKBUF_X4 U3394 ( .I(\SB1_2_27/buf_output[3] ), .Z(\SB2_2_25/i0[10] ) );
  CLKBUF_X4 U3395 ( .I(\SB1_1_22/buf_output[3] ), .Z(\SB2_1_20/i0[10] ) );
  BUF_X4 U3396 ( .I(\MC_ARK_ARC_1_0/buf_output[86] ), .Z(\SB1_1_17/i0_0 ) );
  INV_X1 U3399 ( .I(n361), .ZN(\SB1_0_9/i0[8] ) );
  BUF_X2 U3406 ( .I(n361), .Z(\SB1_0_9/i0[10] ) );
  NAND3_X1 U3408 ( .A1(\SB2_4_28/i0_3 ), .A2(\SB2_4_28/i0_4 ), .A3(
        \SB2_4_28/i0[10] ), .ZN(n2124) );
  NAND3_X1 U3410 ( .A1(\SB2_4_28/i0[10] ), .A2(\SB2_4_28/i1_5 ), .A3(
        \SB2_4_28/i1[9] ), .ZN(\SB2_4_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3411 ( .A1(\SB2_4_28/i0[10] ), .A2(\SB2_4_28/i1[9] ), .A3(
        \SB2_4_28/i1_7 ), .ZN(\SB2_4_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3412 ( .A1(\SB2_4_28/i0_3 ), .A2(\SB2_4_28/i0[10] ), .A3(
        \SB2_4_28/i0[6] ), .ZN(\SB2_4_28/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U3417 ( .I(\MC_ARK_ARC_1_2/buf_output[145] ), .Z(\SB1_3_7/i0[6] ) );
  NAND3_X1 U3426 ( .A1(\RI1[2][116] ), .A2(\SB1_2_12/i0[10] ), .A3(
        \SB1_2_12/i0[6] ), .ZN(\SB1_2_12/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X4 U3428 ( .I(\MC_ARK_ARC_1_1/buf_output[15] ), .Z(\SB1_2_29/i0[10] )
         );
  NAND3_X1 U3430 ( .A1(\SB1_4_16/i0[10] ), .A2(\SB1_4_16/i0_0 ), .A3(
        \SB1_4_16/i0[6] ), .ZN(\SB1_4_16/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3432 ( .A1(\SB1_4_16/i1_5 ), .A2(\SB1_4_16/i0[9] ), .A3(
        \SB1_4_16/i0[6] ), .ZN(n6611) );
  CLKBUF_X2 U3433 ( .I(\MC_ARK_ARC_1_3/buf_output[91] ), .Z(\SB1_4_16/i0[6] )
         );
  INV_X1 U3438 ( .I(n357), .ZN(\SB1_0_11/i0[8] ) );
  NAND3_X1 U3446 ( .A1(\SB2_4_14/i1_5 ), .A2(\SB2_4_14/i0[8] ), .A3(
        \SB2_4_14/i3[0] ), .ZN(\SB2_4_14/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U3447 ( .I(\MC_ARK_ARC_1_4/buf_output[153] ), .ZN(\SB3_6/i0[8] ) );
  CLKBUF_X12 U3449 ( .I(\MC_ARK_ARC_1_4/buf_output[153] ), .Z(\SB3_6/i0[10] )
         );
  NAND3_X1 U3451 ( .A1(\SB2_3_8/i0_0 ), .A2(\SB2_3_8/i0_4 ), .A3(
        \SB2_3_8/i1_5 ), .ZN(n1371) );
  NAND3_X1 U3452 ( .A1(\SB2_3_8/i0[9] ), .A2(\SB2_3_8/i0[6] ), .A3(
        \SB2_3_8/i1_5 ), .ZN(n4512) );
  NAND3_X1 U3456 ( .A1(\SB2_3_8/i1[9] ), .A2(\SB2_3_8/i1_5 ), .A3(
        \SB2_3_8/i0_4 ), .ZN(\SB2_3_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U3460 ( .A1(\SB2_3_9/i0[9] ), .A2(\SB2_3_9/i0[6] ), .A3(
        \SB1_3_10/buf_output[4] ), .ZN(
        \SB2_3_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U3463 ( .A1(\SB1_3_3/i1_5 ), .A2(\SB1_3_3/i0_0 ), .A3(
        \SB1_3_3/i0_4 ), .ZN(\SB1_3_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3464 ( .A1(\SB1_3_6/i0_3 ), .A2(\SB1_3_6/i0[10] ), .A3(
        \SB1_3_6/i0[9] ), .ZN(n1562) );
  NAND3_X1 U3475 ( .A1(\SB1_3_6/i0[7] ), .A2(\SB1_3_6/i0_0 ), .A3(
        \SB1_3_6/i0_3 ), .ZN(\SB1_3_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3476 ( .A1(\SB1_3_6/i0_3 ), .A2(\SB1_3_6/i0[9] ), .A3(
        \SB1_3_6/i0[8] ), .ZN(n1772) );
  NAND3_X1 U3482 ( .A1(\SB1_3_6/i0[10] ), .A2(\SB1_3_6/i0_3 ), .A3(
        \SB1_3_6/i0_4 ), .ZN(n3662) );
  NAND3_X1 U3483 ( .A1(\SB1_3_6/i0_0 ), .A2(\SB1_3_6/i0_3 ), .A3(
        \SB1_3_6/i0_4 ), .ZN(\SB1_3_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3484 ( .A1(\SB1_3_6/i0_3 ), .A2(\SB1_3_6/i0[10] ), .A3(
        \SB1_3_6/i0[6] ), .ZN(\SB1_3_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3487 ( .A1(n1102), .A2(\SB2_2_18/i0[8] ), .A3(\SB2_2_18/i0[6] ), 
        .ZN(n2708) );
  BUF_X4 U3489 ( .I(\SB1_3_5/buf_output[2] ), .Z(\SB2_3_2/i0_0 ) );
  CLKBUF_X4 U3490 ( .I(\MC_ARK_ARC_1_1/buf_output[83] ), .Z(\SB1_2_18/i0_3 )
         );
  INV_X1 U3492 ( .I(\MC_ARK_ARC_1_1/buf_output[83] ), .ZN(\SB1_2_18/i1_5 ) );
  NAND3_X1 U3501 ( .A1(\SB1_0_16/i1_5 ), .A2(\SB1_0_16/i0_0 ), .A3(
        \SB1_0_16/i0_4 ), .ZN(\SB1_0_16/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 U3503 ( .I(\MC_ARK_ARC_1_1/buf_output[86] ), .Z(\SB1_2_17/i0_0 ) );
  CLKBUF_X4 U3504 ( .I(n312), .Z(\SB1_0_2/i0_0 ) );
  INV_X1 U3509 ( .I(\RI1[5][173] ), .ZN(\SB3_3/i1_5 ) );
  NAND3_X2 U3515 ( .A1(\SB1_1_23/i0[7] ), .A2(\SB1_1_23/i0_3 ), .A3(
        \SB1_1_23/i0_0 ), .ZN(\SB1_1_23/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 U3518 ( .I(\SB1_0_13/i0[8] ), .Z(n5428) );
  INV_X1 U3520 ( .I(\MC_ARK_ARC_1_1/buf_output[181] ), .ZN(\SB1_2_1/i1_7 ) );
  BUF_X2 U3521 ( .I(\MC_ARK_ARC_1_1/buf_output[181] ), .Z(\SB1_2_1/i0[6] ) );
  NAND3_X1 U3522 ( .A1(\SB1_2_22/i0[9] ), .A2(\SB1_2_22/i0[10] ), .A3(
        \RI1[2][59] ), .ZN(\SB1_2_22/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3526 ( .A1(\SB1_2_22/i0[10] ), .A2(\SB1_2_22/i0_4 ), .A3(
        \RI1[2][59] ), .ZN(\SB1_2_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3530 ( .A1(\SB1_2_22/i0[6] ), .A2(\RI1[2][59] ), .A3(
        \SB1_2_22/i1[9] ), .ZN(n6941) );
  NOR2_X1 U3539 ( .A1(\RI1[2][59] ), .A2(n6938), .ZN(n7143) );
  NAND3_X1 U3547 ( .A1(\SB1_4_21/i0_3 ), .A2(\SB1_4_21/i1[9] ), .A3(
        \SB1_4_21/i0_4 ), .ZN(n3110) );
  NAND3_X1 U3562 ( .A1(\SB1_4_21/i1[9] ), .A2(\SB1_4_21/i1_7 ), .A3(
        \SB1_4_21/i0[10] ), .ZN(\SB1_4_21/Component_Function_3/NAND4_in[2] )
         );
  NAND2_X1 U3563 ( .A1(\SB1_4_21/i0_3 ), .A2(\SB1_4_21/i1[9] ), .ZN(
        \SB1_4_21/Component_Function_1/NAND4_in[0] ) );
  BUF_X2 U3566 ( .I(\SB2_1_31/i0_4 ), .Z(n5430) );
  NAND3_X1 U3577 ( .A1(\SB2_0_1/i1_5 ), .A2(\SB2_0_1/i0[10] ), .A3(
        \SB2_0_1/i1[9] ), .ZN(\SB2_0_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3579 ( .A1(\SB2_0_1/i0_4 ), .A2(\SB2_0_1/i1_5 ), .A3(
        \SB2_0_1/i1[9] ), .ZN(\SB2_0_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3580 ( .A1(\SB2_0_1/i1[9] ), .A2(\SB2_0_1/i0_3 ), .A3(
        \SB2_0_1/i0[6] ), .ZN(\SB2_0_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3588 ( .A1(\SB2_0_1/i1[9] ), .A2(\SB2_0_1/i0_4 ), .A3(
        \SB2_0_1/i0_3 ), .ZN(\SB2_0_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3591 ( .A1(\SB2_3_21/i0_3 ), .A2(\SB2_3_21/i0[9] ), .A3(
        \SB2_3_21/i0[8] ), .ZN(\SB2_3_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3594 ( .A1(\SB2_3_21/i0_3 ), .A2(\SB2_3_21/i0[8] ), .A3(
        \SB2_3_21/i1_7 ), .ZN(\SB2_3_21/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3598 ( .A1(\SB2_3_21/i0[10] ), .A2(\SB2_3_21/i0[9] ), .A3(
        \SB2_3_21/i0_3 ), .ZN(\SB2_3_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3599 ( .A1(\SB2_3_21/i0[10] ), .A2(\SB2_3_21/i0_3 ), .A3(
        \RI3[3][64] ), .ZN(n6386) );
  NAND3_X1 U3601 ( .A1(\SB2_3_21/i0_0 ), .A2(\SB2_3_21/i0_3 ), .A3(
        \RI3[3][64] ), .ZN(\SB2_3_21/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 U3602 ( .I(\MC_ARK_ARC_1_3/buf_output[157] ), .Z(\SB1_4_5/i0[6] ) );
  NAND3_X1 U3605 ( .A1(\RI1[4][41] ), .A2(\SB1_4_25/i0[8] ), .A3(
        \SB1_4_25/i1_7 ), .ZN(\SB1_4_25/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X4 U3610 ( .I(\MC_ARK_ARC_1_2/buf_output[83] ), .Z(\SB1_3_18/i0_3 )
         );
  NAND3_X1 U3618 ( .A1(\SB1_3_21/i1[9] ), .A2(\SB1_3_21/i1_7 ), .A3(
        \SB1_3_21/i0[10] ), .ZN(\SB1_3_21/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U3620 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0[9] ), .A3(
        \SB1_3_21/i0[10] ), .ZN(n4710) );
  NAND3_X1 U3622 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB2_3_19/i0[6] ), .A3(
        \SB2_3_19/i1[9] ), .ZN(\SB2_3_19/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U3623 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB2_3_19/i1[9] ), .ZN(
        \SB2_3_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3624 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB2_3_19/i0_0 ), .A3(
        \SB1_3_20/buf_output[4] ), .ZN(n5148) );
  CLKBUF_X4 U3625 ( .I(\SB2_4_16/buf_output[3] ), .Z(\RI5[4][105] ) );
  INV_X1 U3626 ( .I(n222), .ZN(\SB1_0_30/i1_7 ) );
  BUF_X4 U3634 ( .I(\MC_ARK_ARC_1_2/buf_output[56] ), .Z(\SB1_3_22/i0_0 ) );
  INV_X1 U3638 ( .I(\MC_ARK_ARC_1_0/buf_output[185] ), .ZN(\SB1_1_1/i1_5 ) );
  CLKBUF_X4 U3647 ( .I(\RI3[0][101] ), .Z(\SB2_0_15/i0_3 ) );
  INV_X1 U3650 ( .I(\RI3[0][101] ), .ZN(\SB2_0_15/i1_5 ) );
  INV_X1 U3653 ( .I(\SB1_3_22/buf_output[1] ), .ZN(\SB2_3_18/i1_7 ) );
  AND3_X2 U3654 ( .A1(\MC_ARK_ARC_1_3/buf_output[73] ), .A2(
        \MC_ARK_ARC_1_3/buf_output[72] ), .A3(\MC_ARK_ARC_1_3/buf_output[76] ), 
        .Z(n3397) );
  INV_X1 U3655 ( .I(\MC_ARK_ARC_1_3/buf_output[72] ), .ZN(\SB1_4_19/i3[0] ) );
  BUF_X2 U3656 ( .I(\MC_ARK_ARC_1_3/buf_output[72] ), .Z(\SB1_4_19/i0[9] ) );
  INV_X1 U3658 ( .I(\SB1_2_18/buf_output[0] ), .ZN(\SB2_2_13/i3[0] ) );
  CLKBUF_X4 U3661 ( .I(\MC_ARK_ARC_1_1/buf_output[167] ), .Z(\SB1_2_4/i0_3 )
         );
  INV_X1 U3662 ( .I(\MC_ARK_ARC_1_1/buf_output[167] ), .ZN(\SB1_2_4/i1_5 ) );
  INV_X1 U3667 ( .I(\SB1_4_17/buf_output[5] ), .ZN(\SB2_4_17/i1_5 ) );
  CLKBUF_X4 U3683 ( .I(\SB1_4_17/buf_output[5] ), .Z(\SB2_4_17/i0_3 ) );
  BUF_X2 U3686 ( .I(\MC_ARK_ARC_1_4/buf_output[32] ), .Z(\SB3_26/i0_0 ) );
  CLKBUF_X4 U3689 ( .I(\SB1_4_24/buf_output[2] ), .Z(\SB2_4_21/i0_0 ) );
  CLKBUF_X4 U3706 ( .I(\MC_ARK_ARC_1_2/buf_output[134] ), .Z(\SB1_3_9/i0_0 )
         );
  INV_X1 U3708 ( .I(\SB1_3_12/buf_output[5] ), .ZN(\SB2_3_12/i1_5 ) );
  CLKBUF_X4 U3709 ( .I(\SB1_3_12/buf_output[5] ), .Z(\SB2_3_12/i0_3 ) );
  INV_X1 U3714 ( .I(\MC_ARK_ARC_1_2/buf_output[187] ), .ZN(\SB1_3_0/i1_7 ) );
  INV_X1 U3715 ( .I(\RI1[3][165] ), .ZN(\SB1_3_4/i0[8] ) );
  BUF_X2 U3719 ( .I(\RI1[3][165] ), .Z(\SB1_3_4/i0[10] ) );
  NAND3_X1 U3723 ( .A1(\SB1_2_1/i0[10] ), .A2(\SB1_2_1/i1[9] ), .A3(
        \SB1_2_1/i1_7 ), .ZN(n4959) );
  NAND3_X1 U3724 ( .A1(\SB1_2_1/i0[10] ), .A2(\SB1_2_1/i1_5 ), .A3(
        \SB1_2_1/i1[9] ), .ZN(n6052) );
  CLKBUF_X4 U3734 ( .I(\MC_ARK_ARC_1_2/buf_output[99] ), .Z(\SB1_3_15/i0[10] )
         );
  CLKBUF_X4 U3739 ( .I(n384), .Z(\SB1_0_28/i0_3 ) );
  INV_X1 U3740 ( .I(n384), .ZN(\SB1_0_28/i1_5 ) );
  CLKBUF_X4 U3741 ( .I(\MC_ARK_ARC_1_3/buf_output[92] ), .Z(\SB1_4_16/i0_0 )
         );
  INV_X1 U3742 ( .I(\MC_ARK_ARC_1_3/buf_output[132] ), .ZN(\SB1_4_9/i3[0] ) );
  INV_X1 U3743 ( .I(\MC_ARK_ARC_1_1/buf_output[113] ), .ZN(\SB1_2_13/i1_5 ) );
  CLKBUF_X4 U3745 ( .I(\MC_ARK_ARC_1_1/buf_output[113] ), .Z(\SB1_2_13/i0_3 )
         );
  CLKBUF_X4 U3748 ( .I(\MC_ARK_ARC_1_4/buf_output[39] ), .Z(\SB3_25/i0[10] )
         );
  NAND3_X1 U3755 ( .A1(\SB1_3_26/i0[10] ), .A2(\SB1_3_26/i0_3 ), .A3(
        \SB1_3_26/i0_4 ), .ZN(\SB1_3_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3756 ( .A1(\SB1_3_26/i0[10] ), .A2(\SB1_3_26/i0_3 ), .A3(
        \SB1_3_26/i0[6] ), .ZN(\SB1_3_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3760 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i0[9] ), .A3(
        \SB1_3_26/i0[10] ), .ZN(n7238) );
  NAND3_X1 U3766 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i0[9] ), .A3(
        \SB1_3_26/i0[8] ), .ZN(n6864) );
  NAND3_X1 U3768 ( .A1(\SB1_3_26/i0_0 ), .A2(\SB1_3_26/i0_3 ), .A3(
        \SB1_3_26/i0[7] ), .ZN(n6104) );
  NAND3_X1 U3776 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i0_4 ), .A3(
        \SB1_3_26/i1[9] ), .ZN(\SB1_3_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3778 ( .A1(\SB1_3_26/i0_4 ), .A2(\SB1_3_26/i0_3 ), .A3(
        \SB1_3_26/i0_0 ), .ZN(n7259) );
  NAND3_X1 U3780 ( .A1(\SB1_2_1/i0_0 ), .A2(\SB1_2_1/i0[6] ), .A3(
        \SB1_2_1/i0[10] ), .ZN(\SB1_2_1/Component_Function_5/NAND4_in[1] ) );
  INV_X1 U3781 ( .I(\MC_ARK_ARC_1_4/buf_output[32] ), .ZN(\SB3_26/i1[9] ) );
  BUF_X4 U3784 ( .I(\SB2_3_24/buf_output[3] ), .Z(\RI5[3][57] ) );
  NAND3_X1 U3790 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[7] ), .A3(
        \SB1_3_31/i0_0 ), .ZN(n4842) );
  NAND3_X1 U3791 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[10] ), .A3(
        \SB1_3_31/i0_4 ), .ZN(\SB1_3_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3793 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i1[9] ), .A3(
        \SB1_3_31/i0_4 ), .ZN(\SB1_3_31/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3794 ( .A1(\SB1_3_31/i0_3 ), .A2(n5441), .A3(\SB1_3_31/i1_7 ), 
        .ZN(n1577) );
  NAND3_X1 U3795 ( .A1(\SB1_3_31/i0[10] ), .A2(\SB1_3_31/i0_3 ), .A3(
        \SB1_3_31/i0[9] ), .ZN(n2653) );
  NAND3_X1 U3797 ( .A1(\SB1_3_31/i0[9] ), .A2(\SB1_3_31/i0_3 ), .A3(n5441), 
        .ZN(\SB1_3_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3802 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[10] ), .A3(
        \SB1_3_31/i0[6] ), .ZN(n4924) );
  NAND3_X1 U3804 ( .A1(\SB2_3_5/i0_0 ), .A2(\SB2_3_5/i0_4 ), .A3(
        \SB2_3_5/i0_3 ), .ZN(\SB2_3_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3805 ( .A1(\SB2_3_5/i1[9] ), .A2(\SB2_3_5/i0_4 ), .A3(
        \SB2_3_5/i0_3 ), .ZN(\SB2_3_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3807 ( .A1(\SB2_3_5/i0_0 ), .A2(\SB2_3_5/i0_4 ), .A3(
        \SB2_3_5/i1_5 ), .ZN(n7224) );
  INV_X1 U3811 ( .I(\SB2_3_5/i0_4 ), .ZN(\SB2_3_5/i0[7] ) );
  INV_X1 U3812 ( .I(\MC_ARK_ARC_1_3/buf_output[0] ), .ZN(\SB1_4_31/i3[0] ) );
  INV_X1 U3815 ( .I(\MC_ARK_ARC_1_3/buf_output[84] ), .ZN(\SB1_4_17/i3[0] ) );
  BUF_X2 U3816 ( .I(\MC_ARK_ARC_1_3/buf_output[84] ), .Z(\SB1_4_17/i0[9] ) );
  NAND3_X1 U3820 ( .A1(\SB3_13/i0_0 ), .A2(\SB3_13/i0_4 ), .A3(\RI1[5][113] ), 
        .ZN(n6638) );
  INV_X2 U3821 ( .I(\RI1[5][113] ), .ZN(\SB3_13/i1_5 ) );
  NAND3_X1 U3822 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0_4 ), .A3(
        \SB2_1_24/i1[9] ), .ZN(n3152) );
  NAND2_X1 U3823 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i1[9] ), .ZN(
        \SB2_1_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3827 ( .A1(\SB2_1_24/i0[10] ), .A2(\SB2_1_24/i1[9] ), .A3(
        \SB2_1_24/i1_7 ), .ZN(\SB2_1_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3833 ( .A1(\SB2_1_24/i1[9] ), .A2(\SB2_1_24/i1_5 ), .A3(
        \SB2_1_24/i0_4 ), .ZN(\SB2_1_24/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U3834 ( .I(\SB2_3_21/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[80] ) );
  CLKBUF_X4 U3836 ( .I(\MC_ARK_ARC_1_1/buf_output[158] ), .Z(\SB1_2_5/i0_0 )
         );
  AND2_X2 U3852 ( .A1(\MC_ARK_ARC_1_3/buf_output[94] ), .A2(
        \MC_ARK_ARC_1_3/buf_output[95] ), .Z(n6846) );
  NAND3_X1 U3856 ( .A1(\SB2_3_25/i0_3 ), .A2(\SB2_3_25/i1_7 ), .A3(
        \SB2_3_25/i0[8] ), .ZN(\SB2_3_25/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3864 ( .A1(\SB2_3_25/i0_3 ), .A2(n5432), .A3(\SB2_3_25/i0[10] ), 
        .ZN(\SB2_3_25/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U3866 ( .A1(\SB2_3_25/i0_3 ), .A2(\SB2_3_25/i1[9] ), .ZN(
        \SB2_3_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3868 ( .A1(\SB2_3_25/i1[9] ), .A2(\SB2_3_25/i0_3 ), .A3(
        \SB2_3_25/i0[6] ), .ZN(\SB2_3_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3872 ( .A1(\SB2_3_25/i0_0 ), .A2(\SB2_3_25/i0_3 ), .A3(
        \SB2_3_25/i0[7] ), .ZN(n1796) );
  NAND3_X1 U3876 ( .A1(\SB2_3_25/i0_4 ), .A2(\SB2_3_25/i0_3 ), .A3(
        \SB2_3_25/i1[9] ), .ZN(\SB2_3_25/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U3877 ( .I(\MC_ARK_ARC_1_2/buf_output[0] ), .ZN(\SB1_3_31/i3[0] ) );
  INV_X1 U3879 ( .I(\SB1_1_24/buf_output[0] ), .ZN(\SB2_1_19/i3[0] ) );
  CLKBUF_X4 U3880 ( .I(\MC_ARK_ARC_1_3/buf_output[81] ), .Z(\SB1_4_18/i0[10] )
         );
  BUF_X2 U3882 ( .I(\MC_ARK_ARC_1_1/buf_output[81] ), .Z(\SB1_2_18/i0[10] ) );
  CLKBUF_X4 U3883 ( .I(\MC_ARK_ARC_1_2/buf_output[81] ), .Z(\SB1_3_18/i0[10] )
         );
  NAND3_X2 U3885 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \SB2_3_20/i0[9] ), .ZN(n2424) );
  NAND3_X1 U3886 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i1_7 ), .A3(
        \SB2_1_6/i0[8] ), .ZN(\SB2_1_6/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3891 ( .A1(\SB2_1_6/i0[10] ), .A2(\SB2_1_6/i0_3 ), .A3(
        \SB2_1_6/i0[9] ), .ZN(\SB2_1_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3892 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0[10] ), .A3(
        \SB2_1_6/i0_4 ), .ZN(n5144) );
  NAND3_X1 U3893 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0_0 ), .A3(
        \SB2_1_6/i0_4 ), .ZN(n5210) );
  NAND3_X1 U3896 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0_4 ), .A3(
        \SB2_1_6/i1[9] ), .ZN(n2435) );
  NAND3_X1 U3898 ( .A1(\SB2_1_6/i1[9] ), .A2(\SB2_1_6/i0_3 ), .A3(
        \SB2_1_6/i0[6] ), .ZN(\SB2_1_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U3901 ( .A1(\SB1_0_3/i0_0 ), .A2(\SB1_0_3/i0[6] ), .A3(
        \SB1_0_3/i0[10] ), .ZN(\SB1_0_3/Component_Function_5/NAND4_in[1] ) );
  INV_X1 U3904 ( .I(\MC_ARK_ARC_1_2/buf_output[63] ), .ZN(\SB1_3_21/i0[8] ) );
  BUF_X2 U3906 ( .I(\MC_ARK_ARC_1_2/buf_output[63] ), .Z(\SB1_3_21/i0[10] ) );
  BUF_X4 U3907 ( .I(\MC_ARK_ARC_1_4/buf_output[189] ), .Z(\SB3_0/i0[10] ) );
  INV_X1 U3910 ( .I(\MC_ARK_ARC_1_1/buf_output[153] ), .ZN(\SB1_2_6/i0[8] ) );
  BUF_X2 U3911 ( .I(\MC_ARK_ARC_1_1/buf_output[153] ), .Z(\SB1_2_6/i0[10] ) );
  NAND3_X1 U3912 ( .A1(\SB1_3_4/i0[10] ), .A2(\SB1_3_4/i1[9] ), .A3(
        \SB1_3_4/i1_7 ), .ZN(n2968) );
  NAND3_X1 U3915 ( .A1(\SB1_3_4/i1_5 ), .A2(\SB1_3_4/i0[10] ), .A3(
        \SB1_3_4/i1[9] ), .ZN(\SB1_3_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3921 ( .A1(\SB1_3_4/i1_5 ), .A2(\SB1_3_4/i1[9] ), .A3(
        \SB1_3_4/i0_4 ), .ZN(n1411) );
  BUF_X4 U3922 ( .I(\MC_ARK_ARC_1_1/buf_output[170] ), .Z(\SB1_2_3/i0_0 ) );
  CLKBUF_X4 U3925 ( .I(\SB2_2_0/buf_output[5] ), .Z(\RI5[2][191] ) );
  CLKBUF_X4 U3929 ( .I(\SB2_3_28/buf_output[2] ), .Z(\RI5[3][38] ) );
  NAND3_X1 U3932 ( .A1(\SB1_2_23/i0_4 ), .A2(\SB1_2_23/i1_7 ), .A3(
        \SB1_2_23/i0[8] ), .ZN(n1915) );
  NAND3_X1 U3935 ( .A1(\SB1_2_23/i0_3 ), .A2(\SB1_2_23/i1_7 ), .A3(
        \SB1_2_23/i0[8] ), .ZN(\SB1_2_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3936 ( .A1(\SB1_2_23/i0[8] ), .A2(\SB1_2_23/i3[0] ), .A3(
        \SB1_2_23/i1_5 ), .ZN(n1335) );
  INV_X1 U3939 ( .I(\MC_ARK_ARC_1_0/buf_output[150] ), .ZN(\SB1_1_6/i3[0] ) );
  BUF_X2 U3940 ( .I(\MC_ARK_ARC_1_0/buf_output[150] ), .Z(\SB1_1_6/i0[9] ) );
  BUF_X2 U3945 ( .I(n237), .Z(\SB1_0_15/i0[6] ) );
  INV_X1 U3946 ( .I(n237), .ZN(\SB1_0_15/i1_7 ) );
  INV_X1 U3962 ( .I(\SB1_2_10/buf_output[0] ), .ZN(\SB2_2_5/i3[0] ) );
  INV_X1 U3970 ( .I(\MC_ARK_ARC_1_0/buf_output[66] ), .ZN(\SB1_1_20/i3[0] ) );
  CLKBUF_X4 U3975 ( .I(n284), .Z(\SB1_0_16/i0_0 ) );
  INV_X1 U3977 ( .I(\MC_ARK_ARC_1_0/buf_output[156] ), .ZN(\SB1_1_5/i3[0] ) );
  NAND3_X1 U3979 ( .A1(\RI1[2][17] ), .A2(\SB1_2_29/i0_0 ), .A3(
        \SB1_2_29/i0_4 ), .ZN(\SB1_2_29/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U3981 ( .I(\MC_ARK_ARC_1_3/buf_output[87] ), .Z(\SB1_4_17/i0[10] )
         );
  INV_X1 U3982 ( .I(\MC_ARK_ARC_1_1/buf_output[173] ), .ZN(\SB1_2_3/i1_5 ) );
  CLKBUF_X4 U3984 ( .I(n396), .Z(\SB1_0_16/i0_3 ) );
  INV_X1 U3986 ( .I(n396), .ZN(\SB1_0_16/i1_5 ) );
  INV_X1 U3990 ( .I(\MC_ARK_ARC_1_1/buf_output[157] ), .ZN(\SB1_2_5/i1_7 ) );
  BUF_X4 U3991 ( .I(\MC_ARK_ARC_1_1/buf_output[157] ), .Z(\SB1_2_5/i0[6] ) );
  INV_X1 U3992 ( .I(\MC_ARK_ARC_1_1/buf_output[141] ), .ZN(\SB1_2_8/i0[8] ) );
  CLKBUF_X4 U3994 ( .I(\SB3_17/buf_output[4] ), .Z(\SB4_16/i0_4 ) );
  CLKBUF_X4 U3997 ( .I(\SB3_30/buf_output[5] ), .Z(\SB4_30/i0_3 ) );
  CLKBUF_X4 U4005 ( .I(\SB3_26/buf_output[2] ), .Z(\SB4_23/i0_0 ) );
  BUF_X2 U4006 ( .I(\SB3_22/buf_output[2] ), .Z(\SB4_19/i0_0 ) );
  BUF_X2 U4007 ( .I(\SB3_15/buf_output[0] ), .Z(\SB4_10/i0[9] ) );
  CLKBUF_X4 U4008 ( .I(\SB3_12/buf_output[5] ), .Z(\SB4_12/i0_3 ) );
  CLKBUF_X4 U4009 ( .I(\SB3_26/buf_output[5] ), .Z(\SB4_26/i0_3 ) );
  CLKBUF_X4 U4010 ( .I(\SB3_19/buf_output[2] ), .Z(\SB4_16/i0_0 ) );
  BUF_X2 U4012 ( .I(\SB3_4/buf_output[0] ), .Z(\SB4_31/i0[9] ) );
  CLKBUF_X4 U4017 ( .I(\SB3_9/buf_output[0] ), .Z(\SB4_4/i0[9] ) );
  CLKBUF_X4 U4018 ( .I(\MC_ARK_ARC_1_4/buf_output[0] ), .Z(\SB3_31/i0[9] ) );
  CLKBUF_X8 U4019 ( .I(\RI1[5][185] ), .Z(\SB3_1/i0_3 ) );
  NAND3_X2 U4021 ( .A1(\SB3_9/i0_3 ), .A2(\SB3_9/i1[9] ), .A3(\SB3_9/i0_4 ), 
        .ZN(n3038) );
  CLKBUF_X4 U4022 ( .I(\RI1[5][137] ), .Z(\SB3_9/i0_3 ) );
  CLKBUF_X4 U4023 ( .I(\MC_ARK_ARC_1_4/buf_output[181] ), .Z(\SB3_1/i0[6] ) );
  CLKBUF_X4 U4026 ( .I(\MC_ARK_ARC_1_4/buf_output[115] ), .Z(\SB3_12/i0[6] )
         );
  CLKBUF_X4 U4027 ( .I(\MC_ARK_ARC_1_4/buf_output[91] ), .Z(\SB3_16/i0[6] ) );
  BUF_X4 U4030 ( .I(n6271), .Z(\SB3_7/i0_3 ) );
  CLKBUF_X4 U4032 ( .I(\SB2_4_25/buf_output[1] ), .Z(\RI5[4][61] ) );
  CLKBUF_X4 U4037 ( .I(\SB2_4_27/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[39] ) );
  CLKBUF_X4 U4041 ( .I(\SB2_4_1/buf_output[2] ), .Z(\RI5[4][8] ) );
  CLKBUF_X4 U4043 ( .I(\SB1_4_19/buf_output[3] ), .Z(\SB2_4_17/i0[10] ) );
  CLKBUF_X4 U4049 ( .I(\SB1_4_31/buf_output[3] ), .Z(\SB2_4_29/i0[10] ) );
  CLKBUF_X4 U4051 ( .I(\SB1_4_14/buf_output[2] ), .Z(\SB2_4_11/i0_0 ) );
  BUF_X2 U4057 ( .I(\SB1_4_19/buf_output[1] ), .Z(\SB2_4_15/i0[6] ) );
  BUF_X4 U4063 ( .I(\SB1_4_10/buf_output[5] ), .Z(\SB2_4_10/i0_3 ) );
  INV_X1 U4067 ( .I(\SB1_4_30/Component_Function_5/NAND4_in[3] ), .ZN(n6961)
         );
  CLKBUF_X4 U4071 ( .I(\MC_ARK_ARC_1_3/buf_output[49] ), .Z(\SB1_4_23/i0[6] )
         );
  BUF_X4 U4072 ( .I(\MC_ARK_ARC_1_3/buf_output[59] ), .Z(\RI1[4][59] ) );
  BUF_X4 U4074 ( .I(\SB2_3_1/buf_output[4] ), .Z(\RI5[3][190] ) );
  CLKBUF_X4 U4076 ( .I(\SB2_3_21/buf_output[3] ), .Z(\RI5[3][75] ) );
  CLKBUF_X4 U4077 ( .I(\SB2_3_12/buf_output[1] ), .Z(\RI5[3][139] ) );
  BUF_X4 U4078 ( .I(\SB2_3_2/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[184] ) );
  CLKBUF_X4 U4079 ( .I(\SB2_3_4/buf_output[5] ), .Z(\RI5[3][167] ) );
  BUF_X4 U4081 ( .I(\SB2_3_27/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[29] ) );
  BUF_X4 U4087 ( .I(\SB2_3_23/buf_output[2] ), .Z(\RI5[3][68] ) );
  CLKBUF_X2 U4092 ( .I(n4677), .Z(n7586) );
  CLKBUF_X2 U4101 ( .I(\SB2_3_4/i0[7] ), .Z(n5683) );
  BUF_X2 U4103 ( .I(\SB1_3_2/buf_output[0] ), .Z(\SB2_3_29/i0[9] ) );
  CLKBUF_X4 U4104 ( .I(\SB1_3_12/buf_output[1] ), .Z(\SB2_3_8/i0[6] ) );
  NAND2_X1 U4108 ( .A1(\SB1_3_21/Component_Function_4/NAND4_in[3] ), .A2(n7261), .ZN(n5272) );
  BUF_X4 U4114 ( .I(\SB1_3_30/buf_output[0] ), .Z(n5432) );
  NAND3_X2 U4116 ( .A1(\SB1_3_29/i0_0 ), .A2(\SB1_3_29/i0[9] ), .A3(
        \SB1_3_29/i0[8] ), .ZN(n4912) );
  NAND2_X1 U4117 ( .A1(\SB1_3_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_4/NAND4_in[1] ), .ZN(n5932) );
  CLKBUF_X4 U4122 ( .I(\MC_ARK_ARC_1_2/buf_output[24] ), .Z(\SB1_3_27/i0[9] )
         );
  BUF_X2 U4132 ( .I(\MC_ARK_ARC_1_2/buf_output[169] ), .Z(\SB1_3_3/i0[6] ) );
  BUF_X2 U4133 ( .I(\MC_ARK_ARC_1_2/buf_output[126] ), .Z(\SB1_3_10/i0[9] ) );
  BUF_X4 U4134 ( .I(\SB2_2_27/buf_output[3] ), .Z(\RI5[2][39] ) );
  BUF_X4 U4137 ( .I(\SB2_2_30/buf_output[1] ), .Z(\RI5[2][31] ) );
  BUF_X2 U4139 ( .I(\SB1_2_2/buf_output[0] ), .Z(\SB2_2_29/i0[9] ) );
  BUF_X4 U4142 ( .I(\SB1_2_15/buf_output[5] ), .Z(\SB2_2_15/i0_3 ) );
  CLKBUF_X4 U4146 ( .I(\SB1_2_11/buf_output[1] ), .Z(\SB2_2_7/i0[6] ) );
  NAND2_X1 U4147 ( .A1(n7286), .A2(n7285), .ZN(n7284) );
  BUF_X2 U4148 ( .I(\MC_ARK_ARC_1_1/buf_output[174] ), .Z(\SB1_2_2/i0[9] ) );
  CLKBUF_X4 U4149 ( .I(\MC_ARK_ARC_1_1/buf_output[63] ), .Z(\SB1_2_21/i0[10] )
         );
  BUF_X4 U4150 ( .I(\SB2_1_6/buf_output[0] ), .Z(\RI5[1][180] ) );
  CLKBUF_X2 U4152 ( .I(\SB2_1_19/i0[7] ), .Z(n5883) );
  CLKBUF_X4 U4153 ( .I(\SB1_1_17/buf_output[3] ), .Z(\SB2_1_15/i0[10] ) );
  BUF_X2 U4157 ( .I(\SB1_1_2/buf_output[0] ), .Z(\SB2_1_29/i0[9] ) );
  CLKBUF_X2 U4159 ( .I(\SB1_1_29/buf_output[4] ), .Z(n5855) );
  NAND2_X1 U4164 ( .A1(\SB1_1_20/Component_Function_4/NAND4_in[0] ), .A2(n7273), .ZN(n2459) );
  CLKBUF_X4 U4166 ( .I(\MC_ARK_ARC_1_0/buf_output[26] ), .Z(\SB1_1_27/i0_0 )
         );
  BUF_X4 U4170 ( .I(\RI5[0][121] ), .Z(n7134) );
  CLKBUF_X4 U4171 ( .I(\SB2_0_15/buf_output[2] ), .Z(\RI5[0][116] ) );
  BUF_X4 U4172 ( .I(\SB2_0_10/buf_output[1] ), .Z(\RI5[0][151] ) );
  BUF_X4 U4175 ( .I(\SB2_0_12/buf_output[4] ), .Z(\RI5[0][124] ) );
  BUF_X4 U4177 ( .I(\SB2_0_5/buf_output[0] ), .Z(\RI5[0][186] ) );
  BUF_X4 U4179 ( .I(\SB2_0_29/buf_output[2] ), .Z(\RI5[0][32] ) );
  INV_X1 U4182 ( .I(n5857), .ZN(n5856) );
  CLKBUF_X2 U4185 ( .I(\SB1_0_25/buf_output[1] ), .Z(n5959) );
  NAND2_X1 U4186 ( .A1(\SB1_0_16/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_16/Component_Function_4/NAND4_in[3] ), .ZN(n6648) );
  NAND2_X1 U4189 ( .A1(n3877), .A2(\SB1_0_16/Component_Function_4/NAND4_in[0] ), .ZN(n6649) );
  BUF_X2 U4191 ( .I(n287), .Z(\SB1_0_14/i0[9] ) );
  CLKBUF_X4 U4195 ( .I(n324), .Z(n5433) );
  INV_X1 U4198 ( .I(n342), .ZN(\SB1_0_19/i0[7] ) );
  NAND3_X1 U4199 ( .A1(\SB1_0_16/i0[9] ), .A2(\SB1_0_16/i0_0 ), .A3(
        \SB1_0_16/i0[8] ), .ZN(\SB1_0_16/Component_Function_4/NAND4_in[0] ) );
  INV_X1 U4200 ( .I(n227), .ZN(\SB1_0_25/i1_7 ) );
  INV_X1 U4203 ( .I(\SB1_0_10/i0_4 ), .ZN(\SB1_0_10/i0[7] ) );
  CLKBUF_X4 U4208 ( .I(n232), .Z(\SB1_0_20/i0[6] ) );
  CLKBUF_X2 U4209 ( .I(n318), .Z(\SB1_0_31/i0_4 ) );
  CLKBUF_X4 U4210 ( .I(n285), .Z(\SB1_0_15/i0[9] ) );
  CLKBUF_X4 U4212 ( .I(n335), .Z(\SB1_0_22/i0[10] ) );
  NAND3_X1 U4213 ( .A1(n5433), .A2(\SB1_0_28/i1_5 ), .A3(\SB1_0_28/i1[9] ), 
        .ZN(n3505) );
  NAND3_X1 U4216 ( .A1(\SB1_0_27/i0_3 ), .A2(\SB1_0_27/i0_4 ), .A3(
        \SB1_0_27/i1[9] ), .ZN(\SB1_0_27/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U4217 ( .A1(\SB1_0_19/i0_3 ), .A2(\SB1_0_19/i1[9] ), .ZN(n3644) );
  NAND3_X1 U4220 ( .A1(\SB1_0_19/i0[10] ), .A2(\SB1_0_19/i0_3 ), .A3(
        \SB1_0_19/i0[9] ), .ZN(n3293) );
  NAND3_X1 U4223 ( .A1(\SB1_0_5/i0[6] ), .A2(\SB1_0_5/i0[9] ), .A3(
        \SB1_0_5/i1_5 ), .ZN(n4577) );
  NAND3_X1 U4225 ( .A1(\SB1_0_1/i0[7] ), .A2(\SB1_0_1/i0_3 ), .A3(
        \SB1_0_1/i0_0 ), .ZN(\SB1_0_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4226 ( .A1(\SB1_0_28/i1_5 ), .A2(\SB1_0_28/i0[8] ), .A3(
        \SB1_0_28/i3[0] ), .ZN(\SB1_0_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4230 ( .A1(\SB1_0_3/i0[10] ), .A2(\SB1_0_3/i0_4 ), .A3(
        \SB1_0_3/i0_3 ), .ZN(\SB1_0_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4238 ( .A1(\SB1_0_27/i0[10] ), .A2(\SB1_0_27/i1[9] ), .A3(
        \SB1_0_27/i1_7 ), .ZN(\SB1_0_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4239 ( .A1(\SB1_0_24/i0[9] ), .A2(\SB1_0_24/i0_0 ), .A3(
        \SB1_0_24/i0[8] ), .ZN(\SB1_0_24/Component_Function_4/NAND4_in[0] ) );
  CLKBUF_X2 U4240 ( .I(n239), .Z(\SB1_0_13/i0[6] ) );
  NAND3_X1 U4243 ( .A1(\SB2_0_21/i1_5 ), .A2(\SB2_0_21/i0[6] ), .A3(
        \SB2_0_21/i0[9] ), .ZN(\SB2_0_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4244 ( .A1(\SB2_0_7/i1[9] ), .A2(\RI3[0][148] ), .A3(
        \SB2_0_7/i0_3 ), .ZN(n5357) );
  NAND3_X1 U4248 ( .A1(\SB2_0_13/i1_5 ), .A2(\SB2_0_13/i0_0 ), .A3(
        \RI3[0][112] ), .ZN(\SB2_0_13/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 U4249 ( .A1(\SB2_0_23/i0_3 ), .A2(\SB2_0_23/i1[9] ), .ZN(n6072) );
  CLKBUF_X4 U4253 ( .I(\SB1_0_1/buf_output[4] ), .Z(\RI3[0][190] ) );
  CLKBUF_X4 U4257 ( .I(\RI3[0][87] ), .Z(\SB2_0_17/i0[10] ) );
  CLKBUF_X4 U4261 ( .I(\SB1_0_3/buf_output[0] ), .Z(\SB2_0_30/i0[9] ) );
  NAND3_X1 U4262 ( .A1(\SB2_0_27/i3[0] ), .A2(\SB2_0_27/i0_0 ), .A3(
        \SB2_0_27/i1_7 ), .ZN(\SB2_0_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4263 ( .A1(\SB2_0_14/i1_7 ), .A2(\SB2_0_14/i0_4 ), .A3(
        \SB2_0_14/i0[8] ), .ZN(\SB2_0_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4264 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i0_0 ), .A3(n2978), 
        .ZN(n6791) );
  NAND3_X1 U4266 ( .A1(\SB2_0_26/i0_3 ), .A2(\SB2_0_26/i1_7 ), .A3(
        \SB2_0_26/i0[8] ), .ZN(\SB2_0_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4270 ( .A1(\SB2_0_26/i3[0] ), .A2(\SB2_0_26/i0_0 ), .A3(
        \SB2_0_26/i1_7 ), .ZN(\SB2_0_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4271 ( .A1(\SB2_0_0/i1_5 ), .A2(\SB2_0_0/i0_0 ), .A3(\RI3[0][190] ), .ZN(\SB2_0_0/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4274 ( .A1(\SB2_0_27/i1_5 ), .A2(\SB2_0_27/i0[10] ), .A3(
        \SB2_0_27/i1[9] ), .ZN(\SB2_0_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4275 ( .A1(n6282), .A2(\SB2_0_5/i0[8] ), .A3(\SB2_0_5/i3[0] ), 
        .ZN(\SB2_0_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4276 ( .A1(\SB2_0_19/i0_0 ), .A2(\SB2_0_19/i1_7 ), .A3(
        \SB2_0_19/i3[0] ), .ZN(n4817) );
  NAND3_X1 U4278 ( .A1(\SB1_1_20/i0[10] ), .A2(\SB1_1_20/i0[9] ), .A3(
        \SB1_1_20/i0_3 ), .ZN(n2645) );
  CLKBUF_X4 U4280 ( .I(\MC_ARK_ARC_1_0/buf_output[9] ), .Z(\SB1_1_30/i0[10] )
         );
  NAND3_X1 U4283 ( .A1(\SB1_1_8/i1_5 ), .A2(\SB1_1_8/i0[6] ), .A3(
        \SB1_1_8/i0[9] ), .ZN(\SB1_1_8/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 U4286 ( .I(\MC_ARK_ARC_1_0/buf_output[40] ), .Z(\SB1_1_25/i0_4 )
         );
  CLKBUF_X4 U4294 ( .I(\MC_ARK_ARC_1_0/buf_output[97] ), .Z(\SB1_1_15/i0[6] )
         );
  BUF_X2 U4296 ( .I(\MC_ARK_ARC_1_0/buf_output[48] ), .Z(\SB1_1_23/i0[9] ) );
  CLKBUF_X4 U4305 ( .I(\MC_ARK_ARC_1_0/buf_output[53] ), .Z(\SB1_1_23/i0_3 )
         );
  INV_X1 U4308 ( .I(\MC_ARK_ARC_1_0/buf_output[102] ), .ZN(\SB1_1_14/i3[0] )
         );
  CLKBUF_X4 U4310 ( .I(\MC_ARK_ARC_1_0/buf_output[158] ), .Z(\SB1_1_5/i0_0 )
         );
  BUF_X2 U4315 ( .I(\MC_ARK_ARC_1_0/buf_output[121] ), .Z(\SB1_1_11/i0[6] ) );
  NAND3_X1 U4319 ( .A1(\SB1_1_8/i1[9] ), .A2(\SB1_1_8/i1_5 ), .A3(
        \SB1_1_8/i0_4 ), .ZN(\SB1_1_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4320 ( .A1(\SB1_1_31/i0_4 ), .A2(\SB1_1_31/i1[9] ), .A3(
        \SB1_1_31/i1_5 ), .ZN(n7555) );
  NAND3_X1 U4321 ( .A1(\SB1_1_13/i0[10] ), .A2(\SB1_1_13/i1_7 ), .A3(
        \SB1_1_13/i1[9] ), .ZN(n7456) );
  NAND3_X1 U4329 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i1[9] ), .A3(
        \SB1_1_6/i0_4 ), .ZN(\SB1_1_6/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4330 ( .A1(\SB1_1_24/i0[9] ), .A2(\SB1_1_24/i0[8] ), .A3(
        \RI1[1][47] ), .ZN(n6697) );
  NAND3_X1 U4332 ( .A1(\SB1_1_12/i1[9] ), .A2(\SB1_1_12/i0_3 ), .A3(
        \SB1_1_12/i0[6] ), .ZN(\SB1_1_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4334 ( .A1(\SB1_1_1/i0[10] ), .A2(\SB1_1_1/i0[9] ), .A3(
        \SB1_1_1/i0_3 ), .ZN(n647) );
  NAND3_X1 U4337 ( .A1(\SB1_1_28/i0[9] ), .A2(\SB1_1_28/i0[10] ), .A3(
        \SB1_1_28/i0_3 ), .ZN(\SB1_1_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4342 ( .A1(\SB1_1_27/i0[9] ), .A2(\SB1_1_27/i0_0 ), .A3(
        \SB1_1_27/i0[8] ), .ZN(\SB1_1_27/Component_Function_4/NAND4_in[0] ) );
  CLKBUF_X8 U4343 ( .I(\RI1[1][149] ), .Z(\SB1_1_7/i0_3 ) );
  NAND3_X1 U4347 ( .A1(\SB1_1_5/i3[0] ), .A2(\SB1_1_5/i0[8] ), .A3(
        \SB1_1_5/i1_5 ), .ZN(n7453) );
  CLKBUF_X4 U4348 ( .I(\MC_ARK_ARC_1_0/buf_output[188] ), .Z(\SB1_1_0/i0_0 )
         );
  NAND3_X1 U4349 ( .A1(\SB1_1_13/i1[9] ), .A2(\SB1_1_13/i1_5 ), .A3(
        \SB1_1_13/i0_4 ), .ZN(\SB1_1_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4353 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i1[9] ), .A3(
        \SB2_1_1/i1_5 ), .ZN(n5001) );
  CLKBUF_X4 U4356 ( .I(\SB1_1_16/buf_output[0] ), .Z(\SB2_1_11/i0[9] ) );
  CLKBUF_X4 U4360 ( .I(\SB1_1_28/buf_output[3] ), .Z(\SB2_1_26/i0[10] ) );
  NAND3_X1 U4363 ( .A1(\SB2_1_25/i0[9] ), .A2(\SB2_1_25/i1_5 ), .A3(
        \SB2_1_25/i0[6] ), .ZN(\SB2_1_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4364 ( .A1(\SB2_1_1/i0_4 ), .A2(\SB2_1_1/i1_7 ), .A3(
        \SB2_1_1/i0[8] ), .ZN(\SB2_1_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4369 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i0_4 ), .A3(
        \SB2_1_1/i0_3 ), .ZN(\SB2_1_1/Component_Function_0/NAND4_in[2] ) );
  INV_X2 U4370 ( .I(\SB2_1_22/i0[7] ), .ZN(\SB2_1_22/i0_4 ) );
  CLKBUF_X4 U4371 ( .I(\SB1_1_25/buf_output[3] ), .Z(\SB2_1_23/i0[10] ) );
  CLKBUF_X4 U4372 ( .I(\SB1_1_5/buf_output[0] ), .Z(\SB2_1_0/i0[9] ) );
  CLKBUF_X4 U4376 ( .I(\SB1_1_31/buf_output[1] ), .Z(\SB2_1_27/i0[6] ) );
  NAND3_X1 U4377 ( .A1(\SB1_1_27/buf_output[3] ), .A2(\SB2_1_25/i1_5 ), .A3(
        \SB2_1_25/i1[9] ), .ZN(\SB2_1_25/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U4383 ( .A1(\SB1_1_27/buf_output[3] ), .A2(\SB2_1_25/i0[9] ), .ZN(
        \SB2_1_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U4384 ( .A1(\SB2_1_9/i1_5 ), .A2(\SB2_1_9/i0_0 ), .A3(
        \SB2_1_9/i0_4 ), .ZN(\SB2_1_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4385 ( .A1(\SB2_1_30/i1_5 ), .A2(\SB2_1_30/i0_4 ), .A3(
        \SB2_1_30/i1[9] ), .ZN(n3086) );
  NAND2_X1 U4386 ( .A1(\SB2_1_15/i0_0 ), .A2(\SB2_1_15/i3[0] ), .ZN(
        \SB2_1_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4392 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i0[10] ), .A3(
        \SB2_1_14/i0[9] ), .ZN(n1991) );
  NAND3_X1 U4395 ( .A1(\SB2_1_18/i0[8] ), .A2(\SB2_1_18/i0[7] ), .A3(
        \SB2_1_18/i0[6] ), .ZN(\SB2_1_18/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U4396 ( .A1(\SB2_1_7/i0_4 ), .A2(\SB2_1_7/i1[9] ), .A3(
        \SB2_1_7/i1_5 ), .ZN(\SB2_1_7/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U4399 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i1[9] ), .ZN(
        \SB2_1_15/Component_Function_1/NAND4_in[0] ) );
  CLKBUF_X2 U4400 ( .I(\RI5[1][8] ), .Z(n3168) );
  CLKBUF_X4 U4401 ( .I(\SB2_1_17/buf_output[5] ), .Z(\RI5[1][89] ) );
  CLKBUF_X4 U4404 ( .I(\SB2_1_27/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[44] ) );
  CLKBUF_X4 U4405 ( .I(\SB2_1_18/buf_output[3] ), .Z(\RI5[1][93] ) );
  INV_X2 U4406 ( .I(\SB1_2_18/i0_4 ), .ZN(\SB1_2_18/i0[7] ) );
  INV_X1 U4407 ( .I(\MC_ARK_ARC_1_1/buf_output[138] ), .ZN(\SB1_2_8/i3[0] ) );
  CLKBUF_X4 U4408 ( .I(\MC_ARK_ARC_1_1/buf_output[110] ), .Z(\SB1_2_13/i0_0 )
         );
  INV_X1 U4409 ( .I(\MC_ARK_ARC_1_1/buf_output[60] ), .ZN(\SB1_2_21/i3[0] ) );
  INV_X1 U4410 ( .I(\MC_ARK_ARC_1_1/buf_output[115] ), .ZN(\SB1_2_12/i1_7 ) );
  CLKBUF_X4 U4416 ( .I(\MC_ARK_ARC_1_1/buf_output[148] ), .Z(\SB1_2_7/i0_4 )
         );
  NAND3_X1 U4417 ( .A1(\SB1_2_21/i1_7 ), .A2(\SB1_2_21/i0[8] ), .A3(
        \SB1_2_21/i0_4 ), .ZN(\SB1_2_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4421 ( .A1(\SB1_2_25/i0[8] ), .A2(\SB1_2_25/i3[0] ), .A3(
        \SB1_2_25/i1_5 ), .ZN(n2203) );
  CLKBUF_X4 U4423 ( .I(\MC_ARK_ARC_1_1/buf_output[118] ), .Z(\SB1_2_12/i0_4 )
         );
  NAND3_X1 U4427 ( .A1(\SB1_2_1/i0_4 ), .A2(\SB1_2_1/i0[8] ), .A3(
        \SB1_2_1/i1_7 ), .ZN(n6467) );
  NAND3_X1 U4428 ( .A1(\SB1_2_31/i0_0 ), .A2(\SB1_2_31/i0_3 ), .A3(
        \SB1_2_31/i0_4 ), .ZN(\SB1_2_31/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U4429 ( .A1(\SB1_2_16/i0_3 ), .A2(\SB1_2_16/i1[9] ), .ZN(
        \SB1_2_16/Component_Function_1/NAND4_in[0] ) );
  CLKBUF_X4 U4432 ( .I(\MC_ARK_ARC_1_1/buf_output[93] ), .Z(\SB1_2_16/i0[10] )
         );
  NAND3_X1 U4433 ( .A1(\SB1_2_22/i0_4 ), .A2(\SB1_2_22/i0[8] ), .A3(
        \SB1_2_22/i1_7 ), .ZN(n6058) );
  NAND3_X1 U4440 ( .A1(\SB1_2_11/i0[8] ), .A2(\SB1_2_11/i0_3 ), .A3(
        \SB1_2_11/i1_7 ), .ZN(\SB1_2_11/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4441 ( .A1(\SB1_2_7/i0_4 ), .A2(\SB1_2_7/i1[9] ), .A3(
        \RI1[2][149] ), .ZN(n7112) );
  NAND3_X1 U4449 ( .A1(\SB1_2_1/i0[8] ), .A2(\SB1_2_1/i0[7] ), .A3(
        \SB1_2_1/i0[6] ), .ZN(\SB1_2_1/Component_Function_0/NAND4_in[1] ) );
  CLKBUF_X4 U4451 ( .I(\MC_ARK_ARC_1_1/buf_output[189] ), .Z(\SB1_2_0/i0[10] )
         );
  NAND3_X1 U4456 ( .A1(\SB1_2_10/i1[9] ), .A2(\SB1_2_10/i0_4 ), .A3(
        \SB1_2_10/i1_5 ), .ZN(n2004) );
  NAND3_X1 U4459 ( .A1(\SB1_2_18/i0[7] ), .A2(\SB1_2_18/i0_0 ), .A3(
        \SB1_2_18/i0_3 ), .ZN(n5129) );
  CLKBUF_X4 U4460 ( .I(\MC_ARK_ARC_1_1/buf_output[39] ), .Z(\SB1_2_25/i0[10] )
         );
  NAND3_X1 U4461 ( .A1(\SB1_2_5/i1_7 ), .A2(\SB1_2_5/i0[8] ), .A3(
        \SB1_2_5/i0_4 ), .ZN(\SB1_2_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4464 ( .A1(\SB1_2_11/i0[8] ), .A2(\SB1_2_11/i0[7] ), .A3(
        \SB1_2_11/i0[6] ), .ZN(\SB1_2_11/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U4466 ( .A1(\SB1_2_31/i1_7 ), .A2(\SB1_2_31/i0[8] ), .A3(
        \SB1_2_31/i0_4 ), .ZN(\SB1_2_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4468 ( .A1(\SB1_2_5/i0_0 ), .A2(\SB1_2_5/i0[8] ), .A3(
        \SB1_2_5/i0[9] ), .ZN(n2991) );
  NAND2_X1 U4471 ( .A1(n2604), .A2(\SB1_2_22/Component_Function_4/NAND4_in[2] ), .ZN(n4546) );
  NAND2_X1 U4472 ( .A1(\SB1_2_19/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_2_19/Component_Function_4/NAND4_in[1] ), .ZN(n6866) );
  NAND3_X1 U4473 ( .A1(\SB1_2_27/i0[8] ), .A2(\SB1_2_27/i3[0] ), .A3(
        \SB1_2_27/i1_5 ), .ZN(n6187) );
  NAND3_X1 U4474 ( .A1(\SB1_2_0/i0_4 ), .A2(\SB1_2_0/i0[9] ), .A3(
        \SB1_2_0/i0[6] ), .ZN(n6250) );
  INV_X1 U4475 ( .I(\SB1_2_1/buf_output[1] ), .ZN(\SB2_2_29/i1_7 ) );
  CLKBUF_X4 U4477 ( .I(\SB1_2_19/buf_output[3] ), .Z(\SB2_2_17/i0[10] ) );
  CLKBUF_X4 U4479 ( .I(\SB1_2_11/buf_output[2] ), .Z(\SB2_2_8/i0_0 ) );
  INV_X1 U4480 ( .I(\SB1_2_22/buf_output[1] ), .ZN(\SB2_2_18/i1_7 ) );
  CLKBUF_X4 U4481 ( .I(\SB1_2_9/buf_output[3] ), .Z(\SB2_2_7/i0[10] ) );
  CLKBUF_X4 U4485 ( .I(\SB1_2_27/buf_output[2] ), .Z(\SB2_2_24/i0_0 ) );
  CLKBUF_X4 U4488 ( .I(\SB1_2_9/buf_output[5] ), .Z(\SB2_2_9/i0_3 ) );
  INV_X1 U4490 ( .I(\SB1_2_5/buf_output[1] ), .ZN(\SB2_2_1/i1_7 ) );
  INV_X1 U4495 ( .I(\SB1_2_10/buf_output[1] ), .ZN(\SB2_2_6/i1_7 ) );
  CLKBUF_X4 U4499 ( .I(\SB1_2_0/buf_output[0] ), .Z(\SB2_2_27/i0[9] ) );
  NAND3_X1 U4501 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0[9] ), .A3(
        \SB2_2_14/i0[10] ), .ZN(\SB2_2_14/Component_Function_4/NAND4_in[2] )
         );
  CLKBUF_X4 U4504 ( .I(\SB1_2_14/buf_output[1] ), .Z(\SB2_2_10/i0[6] ) );
  NAND3_X1 U4505 ( .A1(\SB2_2_29/i1_5 ), .A2(\SB2_2_29/i0[6] ), .A3(
        \SB2_2_29/i0[9] ), .ZN(\SB2_2_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4506 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0[7] ), .A3(
        \SB2_2_16/i0_0 ), .ZN(n1983) );
  NAND3_X1 U4507 ( .A1(\SB2_2_18/i0_3 ), .A2(\SB2_2_18/i0[10] ), .A3(
        \SB2_2_18/i0[9] ), .ZN(n5331) );
  NAND3_X1 U4508 ( .A1(\SB2_2_19/i0_0 ), .A2(\SB2_2_19/i0[10] ), .A3(
        \SB2_2_19/i0[6] ), .ZN(\SB2_2_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4510 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i0_0 ), .A3(
        \SB2_2_17/i0[7] ), .ZN(n7034) );
  NAND3_X1 U4515 ( .A1(\SB2_2_28/i0_0 ), .A2(\SB2_2_28/i0_3 ), .A3(
        \SB2_2_28/i0[7] ), .ZN(n1970) );
  NAND3_X1 U4516 ( .A1(\SB2_2_8/i0_0 ), .A2(\SB2_2_8/i0_3 ), .A3(
        \SB2_2_8/i0[7] ), .ZN(n4469) );
  CLKBUF_X4 U4517 ( .I(\SB1_2_30/buf_output[0] ), .Z(\SB2_2_25/i0[9] ) );
  NAND2_X1 U4519 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i1[9] ), .ZN(
        \SB2_2_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U4520 ( .A1(\SB2_2_25/i0_4 ), .A2(\SB2_2_25/i0[8] ), .A3(
        \SB2_2_25/i1_7 ), .ZN(n6186) );
  NAND3_X1 U4521 ( .A1(\SB2_2_6/i0[10] ), .A2(\SB2_2_6/i0_3 ), .A3(
        \SB2_2_6/i0[9] ), .ZN(n6348) );
  NAND3_X1 U4522 ( .A1(\SB2_2_13/i0[8] ), .A2(\SB2_2_13/i3[0] ), .A3(
        \SB2_2_13/i1_5 ), .ZN(n7092) );
  CLKBUF_X4 U4523 ( .I(\SB1_2_24/buf_output[3] ), .Z(\SB2_2_22/i0[10] ) );
  NAND2_X1 U4524 ( .A1(\SB2_2_22/i0[10] ), .A2(\SB2_2_22/i0[9] ), .ZN(
        \SB2_2_22/Component_Function_0/NAND4_in[0] ) );
  CLKBUF_X4 U4527 ( .I(\SB2_2_11/buf_output[1] ), .Z(\RI5[2][145] ) );
  INV_X2 U4528 ( .I(\SB1_3_6/i0_4 ), .ZN(\SB1_3_6/i0[7] ) );
  INV_X2 U4530 ( .I(\SB1_3_20/i0_4 ), .ZN(\SB1_3_20/i0[7] ) );
  INV_X1 U4531 ( .I(\MC_ARK_ARC_1_2/buf_output[67] ), .ZN(\SB1_3_20/i1_7 ) );
  INV_X1 U4532 ( .I(\MC_ARK_ARC_1_2/buf_output[133] ), .ZN(\SB1_3_9/i1_7 ) );
  CLKBUF_X4 U4535 ( .I(\MC_ARK_ARC_1_2/buf_output[146] ), .Z(\SB1_3_7/i0_0 )
         );
  CLKBUF_X2 U4536 ( .I(\MC_ARK_ARC_1_2/buf_output[121] ), .Z(\SB1_3_11/i0[6] )
         );
  INV_X1 U4537 ( .I(\MC_ARK_ARC_1_2/buf_output[47] ), .ZN(\SB1_3_24/i1_5 ) );
  NAND3_X1 U4539 ( .A1(\SB1_3_14/i0[10] ), .A2(\RI1[3][107] ), .A3(
        \SB1_3_14/i0[9] ), .ZN(n2202) );
  NAND3_X1 U4540 ( .A1(\SB1_3_9/i1_5 ), .A2(\SB1_3_9/i0_0 ), .A3(
        \SB1_3_9/i0_4 ), .ZN(\SB1_3_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4543 ( .A1(\SB1_3_2/i1_5 ), .A2(\SB1_3_2/i0[6] ), .A3(
        \SB1_3_2/i0[9] ), .ZN(\SB1_3_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4544 ( .A1(\SB1_3_9/i0_0 ), .A2(\SB1_3_9/i0_3 ), .A3(
        \SB1_3_9/i0_4 ), .ZN(\SB1_3_9/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U4545 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i1[9] ), .ZN(
        \SB1_3_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U4548 ( .A1(\SB1_3_28/i0[10] ), .A2(\SB1_3_28/i0_4 ), .A3(
        \SB1_3_28/i0_3 ), .ZN(\SB1_3_28/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 U4549 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i1[9] ), .ZN(
        \SB1_3_21/Component_Function_1/NAND4_in[0] ) );
  CLKBUF_X4 U4550 ( .I(\MC_ARK_ARC_1_2/buf_output[93] ), .Z(\SB1_3_16/i0[10] )
         );
  NAND3_X1 U4551 ( .A1(\SB1_3_18/i0[7] ), .A2(\SB1_3_18/i0_3 ), .A3(
        \SB1_3_18/i0_0 ), .ZN(\SB1_3_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4552 ( .A1(\SB1_3_0/i0[9] ), .A2(\SB1_3_0/i1_5 ), .A3(
        \SB1_3_0/i0[6] ), .ZN(n6801) );
  NAND2_X1 U4553 ( .A1(\SB1_3_26/i0_0 ), .A2(\SB1_3_26/i3[0] ), .ZN(
        \SB1_3_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4554 ( .A1(\SB1_3_9/i0_3 ), .A2(\SB1_3_9/i1_7 ), .A3(
        \SB1_3_9/i0[8] ), .ZN(\SB1_3_9/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4556 ( .A1(\SB1_3_24/i0[7] ), .A2(\SB1_3_24/i0_3 ), .A3(
        \SB1_3_24/i0_0 ), .ZN(\SB1_3_24/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U4557 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i3[0] ), .ZN(
        \SB1_3_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4558 ( .A1(\SB1_3_9/i0_0 ), .A2(\SB1_3_9/i0[10] ), .A3(
        \SB1_3_9/i0[6] ), .ZN(n5253) );
  NAND3_X1 U4563 ( .A1(\SB1_3_5/i0[8] ), .A2(\SB1_3_5/i3[0] ), .A3(
        \SB1_3_5/i1_5 ), .ZN(n3879) );
  NAND3_X1 U4564 ( .A1(\SB1_3_23/i0[10] ), .A2(\SB1_3_23/i0_3 ), .A3(
        \SB1_3_23/i0[9] ), .ZN(n3187) );
  NAND3_X1 U4565 ( .A1(\SB1_3_1/i0[8] ), .A2(\SB1_3_1/i3[0] ), .A3(
        \SB1_3_1/i1_5 ), .ZN(\SB1_3_1/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X4 U4568 ( .I(\MC_ARK_ARC_1_2/buf_output[186] ), .Z(\SB1_3_0/i0[9] )
         );
  NAND3_X1 U4569 ( .A1(\SB1_3_13/i0[10] ), .A2(\SB1_3_13/i1[9] ), .A3(
        \SB1_3_13/i1_5 ), .ZN(n4634) );
  NAND3_X1 U4572 ( .A1(\SB1_3_26/i1[9] ), .A2(\SB1_3_26/i1_5 ), .A3(
        \SB1_3_26/i0_4 ), .ZN(\SB1_3_26/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U4577 ( .I(\SB1_3_7/buf_output[0] ), .Z(\SB2_3_2/i0[9] ) );
  CLKBUF_X4 U4578 ( .I(\SB1_3_23/buf_output[2] ), .Z(\SB2_3_20/i0_0 ) );
  CLKBUF_X1 U4579 ( .I(n1427), .Z(n6716) );
  INV_X1 U4580 ( .I(\SB1_3_20/buf_output[4] ), .ZN(\SB2_3_19/i0[7] ) );
  INV_X1 U4581 ( .I(\SB1_3_16/buf_output[1] ), .ZN(\SB2_3_12/i1_7 ) );
  CLKBUF_X4 U4582 ( .I(\SB1_3_0/buf_output[1] ), .Z(\SB2_3_28/i0[6] ) );
  NAND3_X1 U4583 ( .A1(n5432), .A2(\SB2_3_25/i1_5 ), .A3(\SB2_3_25/i0[6] ), 
        .ZN(\SB2_3_25/Component_Function_1/NAND4_in[2] ) );
  INV_X1 U4585 ( .I(\SB1_3_9/buf_output[0] ), .ZN(\SB2_3_4/i3[0] ) );
  CLKBUF_X4 U4589 ( .I(\SB1_3_7/buf_output[2] ), .Z(\SB2_3_4/i0_0 ) );
  NAND3_X1 U4591 ( .A1(\SB2_3_23/i1_5 ), .A2(\SB2_3_23/i0[6] ), .A3(
        \SB2_3_23/i0[9] ), .ZN(\SB2_3_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4593 ( .A1(\SB2_3_8/i0[10] ), .A2(\SB2_3_8/i0_3 ), .A3(
        \SB2_3_8/i0[9] ), .ZN(\SB2_3_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4595 ( .A1(\SB2_3_14/i0_0 ), .A2(\SB2_3_14/i0_3 ), .A3(
        \SB2_3_14/i0[7] ), .ZN(n5009) );
  CLKBUF_X4 U4596 ( .I(\SB1_3_5/buf_output[3] ), .Z(\SB2_3_3/i0[10] ) );
  NAND3_X1 U4597 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i0[10] ), .A3(
        \SB2_3_27/i0_4 ), .ZN(\SB2_3_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4598 ( .A1(\SB2_3_14/i0_3 ), .A2(\SB2_3_14/i1_7 ), .A3(
        \SB2_3_14/i0[8] ), .ZN(\SB2_3_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4599 ( .A1(\SB2_3_3/i1[9] ), .A2(\SB2_3_3/i1_5 ), .A3(
        \SB2_3_3/i0_4 ), .ZN(\SB2_3_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4602 ( .A1(\SB2_3_17/i0_4 ), .A2(\SB2_3_17/i1_7 ), .A3(
        \SB2_3_17/i0[8] ), .ZN(n6200) );
  NAND2_X1 U4604 ( .A1(\SB2_3_8/i0_0 ), .A2(\SB2_3_8/i3[0] ), .ZN(
        \SB2_3_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4607 ( .A1(\SB2_3_19/i1[9] ), .A2(\SB1_3_20/buf_output[4] ), .A3(
        \SB2_3_19/i1_5 ), .ZN(n2823) );
  NAND3_X1 U4609 ( .A1(\SB2_3_0/i1[9] ), .A2(\SB2_3_0/i1_5 ), .A3(
        \SB2_3_0/i0_4 ), .ZN(\SB2_3_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4611 ( .A1(\SB2_3_8/i0_3 ), .A2(\SB2_3_8/i0_0 ), .A3(
        \SB2_3_8/i0_4 ), .ZN(\SB2_3_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4615 ( .A1(\SB2_3_12/i1[9] ), .A2(\SB2_3_12/i1_5 ), .A3(n592), 
        .ZN(\SB2_3_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4618 ( .A1(\SB2_3_15/i0[9] ), .A2(\SB2_3_15/i0[6] ), .A3(
        \SB2_3_15/i1_5 ), .ZN(n3914) );
  NAND2_X1 U4620 ( .A1(n5432), .A2(\SB2_3_25/i0[10] ), .ZN(n6373) );
  NAND3_X1 U4621 ( .A1(\SB2_3_24/i0[6] ), .A2(\SB2_3_24/i1_5 ), .A3(
        \SB2_3_24/i0[9] ), .ZN(\SB2_3_24/Component_Function_1/NAND4_in[2] ) );
  INV_X1 U4623 ( .I(n194), .ZN(n516) );
  NAND3_X1 U4628 ( .A1(\SB2_3_21/i0_0 ), .A2(\RI3[3][64] ), .A3(
        \SB2_3_21/i1_5 ), .ZN(n7013) );
  CLKBUF_X4 U4630 ( .I(\SB2_3_24/buf_output[1] ), .Z(\RI5[3][67] ) );
  INV_X1 U4631 ( .I(\MC_ARK_ARC_1_3/buf_output[61] ), .ZN(\SB1_4_21/i1_7 ) );
  INV_X4 U4636 ( .I(\RI1[4][131] ), .ZN(\SB1_4_10/i1_5 ) );
  NAND3_X1 U4638 ( .A1(\SB1_4_2/i0_4 ), .A2(\SB1_4_2/i1_5 ), .A3(
        \SB1_4_2/i1[9] ), .ZN(n5994) );
  CLKBUF_X4 U4640 ( .I(\MC_ARK_ARC_1_3/buf_output[74] ), .Z(\SB1_4_19/i0_0 )
         );
  CLKBUF_X4 U4642 ( .I(\MC_ARK_ARC_1_3/buf_output[93] ), .Z(\SB1_4_16/i0[10] )
         );
  CLKBUF_X4 U4643 ( .I(\MC_ARK_ARC_1_3/buf_output[136] ), .Z(\SB1_4_9/i0_4 )
         );
  CLKBUF_X4 U4648 ( .I(\MC_ARK_ARC_1_3/buf_output[148] ), .Z(\SB1_4_7/i0_4 )
         );
  CLKBUF_X4 U4649 ( .I(\MC_ARK_ARC_1_3/buf_output[111] ), .Z(\SB1_4_13/i0[10] ) );
  INV_X1 U4650 ( .I(\RI1[4][53] ), .ZN(\SB1_4_23/i1_5 ) );
  NAND2_X1 U4655 ( .A1(\SB1_4_6/i1[9] ), .A2(\RI1[4][155] ), .ZN(n5605) );
  NAND2_X1 U4656 ( .A1(\SB1_4_1/i0[10] ), .A2(\SB1_4_1/i0[9] ), .ZN(
        \SB1_4_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U4657 ( .A1(\SB1_4_26/i1_5 ), .A2(\SB1_4_26/i0[8] ), .A3(
        \SB1_4_26/i3[0] ), .ZN(\SB1_4_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4663 ( .A1(\SB1_4_15/i0[9] ), .A2(\SB1_4_15/i0[8] ), .A3(
        \SB1_4_15/i0_3 ), .ZN(n5400) );
  NAND3_X1 U4665 ( .A1(\SB1_4_10/i1_5 ), .A2(\SB1_4_10/i3[0] ), .A3(
        \SB1_4_10/i0[8] ), .ZN(n4246) );
  NAND2_X1 U4666 ( .A1(\SB1_4_31/i0_0 ), .A2(\SB1_4_31/i3[0] ), .ZN(
        \SB1_4_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4667 ( .A1(\SB1_4_22/i0[10] ), .A2(\SB1_4_22/i1[9] ), .A3(
        \SB1_4_22/i1_7 ), .ZN(\SB1_4_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4670 ( .A1(\SB1_4_21/i0[8] ), .A2(\SB1_4_21/i0[7] ), .A3(
        \SB1_4_21/i0[6] ), .ZN(\SB1_4_21/Component_Function_0/NAND4_in[1] ) );
  INV_X1 U4672 ( .I(\MC_ARK_ARC_1_3/buf_output[19] ), .ZN(\SB1_4_28/i1_7 ) );
  NAND3_X1 U4680 ( .A1(\SB1_4_1/i1_7 ), .A2(\SB1_4_1/i0[8] ), .A3(
        \SB1_4_1/i0_4 ), .ZN(\SB1_4_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4683 ( .A1(\SB1_4_2/i1_5 ), .A2(\SB1_4_2/i0[6] ), .A3(
        \SB1_4_2/i0[9] ), .ZN(\SB1_4_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4690 ( .A1(\SB1_4_30/i1_7 ), .A2(\SB1_4_30/i0[8] ), .A3(
        \SB1_4_30/i0_4 ), .ZN(\SB1_4_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4691 ( .A1(\SB1_4_26/i0_3 ), .A2(\SB1_4_26/i1_7 ), .A3(
        \SB1_4_26/i0[8] ), .ZN(\SB1_4_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4693 ( .A1(\SB1_4_15/i0[7] ), .A2(\SB1_4_15/i0_3 ), .A3(
        \SB1_4_15/i0_0 ), .ZN(\SB1_4_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4697 ( .A1(n6774), .A2(\SB1_4_22/i1_5 ), .A3(\SB1_4_22/i0_4 ), 
        .ZN(\SB1_4_22/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U4698 ( .I(\SB1_4_6/buf_output[4] ), .ZN(\SB2_4_5/i0[7] ) );
  CLKBUF_X4 U4700 ( .I(\SB1_4_10/buf_output[2] ), .Z(\SB2_4_7/i0_0 ) );
  CLKBUF_X4 U4701 ( .I(\SB1_4_31/buf_output[2] ), .Z(\SB2_4_28/i0_0 ) );
  CLKBUF_X4 U4702 ( .I(\SB1_4_20/buf_output[3] ), .Z(\SB2_4_18/i0[10] ) );
  CLKBUF_X4 U4704 ( .I(\SB1_4_0/buf_output[4] ), .Z(\SB2_4_31/i0_4 ) );
  CLKBUF_X4 U4705 ( .I(\SB1_4_29/buf_output[3] ), .Z(\SB2_4_27/i0[10] ) );
  CLKBUF_X4 U4708 ( .I(\SB1_4_15/buf_output[3] ), .Z(\SB2_4_13/i0[10] ) );
  NAND3_X1 U4709 ( .A1(\SB2_4_15/i0_3 ), .A2(\SB2_4_15/i0[10] ), .A3(
        \SB2_4_15/i0[9] ), .ZN(n1849) );
  NAND2_X1 U4712 ( .A1(\SB2_4_19/i0[10] ), .A2(\SB2_4_19/i0[9] ), .ZN(
        \SB2_4_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U4715 ( .A1(\SB2_4_7/i1_7 ), .A2(\SB2_4_7/i0[8] ), .A3(
        \RI3[4][148] ), .ZN(\SB2_4_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4716 ( .A1(\SB2_4_4/i1_5 ), .A2(\SB2_4_4/i0[6] ), .A3(
        \SB2_4_4/i0[9] ), .ZN(\SB2_4_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4717 ( .A1(\SB2_4_12/i3[0] ), .A2(\SB2_4_12/i0_0 ), .A3(
        \SB2_4_12/i1_7 ), .ZN(\SB2_4_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4718 ( .A1(\SB2_4_14/i0_4 ), .A2(\SB2_4_14/i1[9] ), .A3(
        \SB2_4_14/i1_5 ), .ZN(n7486) );
  NAND3_X1 U4719 ( .A1(\SB2_4_9/i0_0 ), .A2(\SB2_4_9/i0_3 ), .A3(
        \SB2_4_9/i0[7] ), .ZN(n4355) );
  NAND3_X1 U4722 ( .A1(\SB2_4_27/i0_3 ), .A2(\SB2_4_27/i0_0 ), .A3(
        \SB2_4_27/i0[7] ), .ZN(n7069) );
  NAND3_X1 U4723 ( .A1(\SB2_4_7/i0_3 ), .A2(\SB2_4_7/i0_0 ), .A3(
        \SB2_4_7/i0[7] ), .ZN(n6571) );
  NAND3_X1 U4724 ( .A1(\SB2_4_7/i0_3 ), .A2(\SB2_4_7/i0[10] ), .A3(
        \SB2_4_7/i0[9] ), .ZN(n6627) );
  NAND3_X1 U4725 ( .A1(\SB2_4_28/i0_0 ), .A2(n4000), .A3(\SB2_4_28/i0[9] ), 
        .ZN(n7198) );
  NAND3_X1 U4730 ( .A1(\SB2_4_6/i1[9] ), .A2(\SB2_4_6/i1_7 ), .A3(
        \SB2_4_6/i0[10] ), .ZN(\SB2_4_6/Component_Function_3/NAND4_in[2] ) );
  CLKBUF_X4 U4732 ( .I(\SB2_4_9/buf_output[3] ), .Z(\RI5[4][147] ) );
  INV_X1 U4734 ( .I(n41), .ZN(n564) );
  INV_X1 U4739 ( .I(n121), .ZN(n515) );
  INV_X1 U4741 ( .I(n67), .ZN(n531) );
  INV_X1 U4742 ( .I(n26), .ZN(n526) );
  INV_X1 U4746 ( .I(\MC_ARK_ARC_1_4/buf_output[114] ), .ZN(\SB3_12/i3[0] ) );
  CLKBUF_X4 U4747 ( .I(\MC_ARK_ARC_1_4/buf_output[116] ), .Z(\SB3_12/i0_0 ) );
  CLKBUF_X4 U4748 ( .I(\MC_ARK_ARC_1_4/buf_output[90] ), .Z(\SB3_16/i0[9] ) );
  CLKBUF_X4 U4752 ( .I(\MC_ARK_ARC_1_4/buf_output[68] ), .Z(\SB3_20/i0_0 ) );
  CLKBUF_X2 U4754 ( .I(\MC_ARK_ARC_1_4/buf_output[174] ), .Z(\SB3_2/i0[9] ) );
  NAND3_X1 U4755 ( .A1(\SB3_19/i0[6] ), .A2(\SB3_19/i1_5 ), .A3(\SB3_19/i0[9] ), .ZN(\SB3_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4758 ( .A1(\SB3_11/i1[9] ), .A2(\SB3_11/i0_4 ), .A3(\SB3_11/i1_5 ), 
        .ZN(n2215) );
  NAND3_X1 U4759 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i1[9] ), .A3(\SB3_2/i0[6] ), 
        .ZN(\SB3_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4760 ( .A1(\SB3_28/i0_3 ), .A2(\SB3_28/i0[9] ), .A3(
        \SB3_28/i0[10] ), .ZN(n6823) );
  NAND3_X1 U4761 ( .A1(\SB3_31/i0[9] ), .A2(\SB3_31/i0[6] ), .A3(\SB3_31/i1_5 ), .ZN(\SB3_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4765 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i1[9] ), .A3(\SB3_31/i0[6] ), .ZN(\SB3_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U4766 ( .A1(\SB3_7/i0[8] ), .A2(\SB3_7/i1_5 ), .A3(\SB3_7/i3[0] ), 
        .ZN(\SB3_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4770 ( .A1(\SB3_2/i0[9] ), .A2(\SB3_2/i0[6] ), .A3(\SB3_2/i1_5 ), 
        .ZN(n2597) );
  NAND3_X1 U4771 ( .A1(\SB3_31/i0[6] ), .A2(\SB3_31/i0[9] ), .A3(\SB3_31/i0_4 ), .ZN(n4751) );
  NAND3_X1 U4774 ( .A1(\SB3_25/i0_4 ), .A2(\SB3_25/i1[9] ), .A3(\SB3_25/i1_5 ), 
        .ZN(n998) );
  CLKBUF_X4 U4777 ( .I(\MC_ARK_ARC_1_4/buf_output[10] ), .Z(\SB3_30/i0_4 ) );
  NAND3_X1 U4778 ( .A1(\SB3_20/i0_3 ), .A2(\SB3_20/i0[10] ), .A3(
        \SB3_20/i0[9] ), .ZN(n4759) );
  NAND3_X1 U4779 ( .A1(\SB3_7/i0[7] ), .A2(\SB3_7/i0_3 ), .A3(\SB3_7/i0_0 ), 
        .ZN(\SB3_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4788 ( .A1(\SB3_2/i0_0 ), .A2(\SB3_2/i0[6] ), .A3(\SB3_2/i0[10] ), 
        .ZN(\SB3_2/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4790 ( .A1(\SB3_20/i0_0 ), .A2(\SB3_20/i0[6] ), .A3(
        \SB3_20/i0[10] ), .ZN(\SB3_20/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X4 U4793 ( .I(\MC_ARK_ARC_1_4/buf_output[108] ), .Z(\SB3_13/i0[9] )
         );
  CLKBUF_X4 U4794 ( .I(\MC_ARK_ARC_1_4/buf_output[105] ), .Z(\SB3_14/i0[10] )
         );
  NAND3_X1 U4796 ( .A1(\SB3_11/i0_3 ), .A2(\SB3_11/i0_0 ), .A3(\SB3_11/i0[7] ), 
        .ZN(n6514) );
  NAND3_X1 U4797 ( .A1(\SB3_6/i0_0 ), .A2(\SB3_6/i0[6] ), .A3(\SB3_6/i0[10] ), 
        .ZN(\SB3_6/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4798 ( .A1(\SB3_4/i0[10] ), .A2(\SB3_4/i0_3 ), .A3(\SB3_4/i0[6] ), 
        .ZN(n1846) );
  NAND3_X1 U4799 ( .A1(\SB3_26/i1_5 ), .A2(\SB3_26/i0[6] ), .A3(\SB3_26/i0[9] ), .ZN(\SB3_26/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 U4800 ( .I(\SB3_21/buf_output[0] ), .Z(\SB4_16/i0[9] ) );
  CLKBUF_X4 U4805 ( .I(\SB3_5/buf_output[5] ), .Z(\SB4_5/i0_3 ) );
  CLKBUF_X4 U4807 ( .I(\SB3_25/buf_output[0] ), .Z(\SB4_20/i0[9] ) );
  NAND3_X1 U4808 ( .A1(\SB4_7/i0_0 ), .A2(\SB4_7/i0_3 ), .A3(\SB4_7/i0_4 ), 
        .ZN(n4862) );
  NAND3_X1 U4809 ( .A1(\SB4_15/i0[7] ), .A2(\SB4_15/i0_3 ), .A3(\SB4_15/i0_0 ), 
        .ZN(\SB4_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4812 ( .A1(\SB4_12/i0[8] ), .A2(\SB4_12/i0[7] ), .A3(
        \SB4_12/i0[6] ), .ZN(\SB4_12/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U4814 ( .A1(\SB4_26/i0_3 ), .A2(\SB4_26/i0[10] ), .A3(
        \SB4_26/i0[6] ), .ZN(n5168) );
  NAND2_X1 U4817 ( .A1(\SB4_3/i0[10] ), .A2(\SB4_3/i0[9] ), .ZN(
        \SB4_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U4819 ( .A1(\SB4_5/i0_0 ), .A2(\SB4_5/i0_3 ), .A3(\SB4_5/i0_4 ), 
        .ZN(\SB4_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4823 ( .A1(\SB4_31/i0[10] ), .A2(\SB4_31/i0_4 ), .A3(\SB4_31/i0_3 ), .ZN(\SB4_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4826 ( .A1(\SB4_31/i0_3 ), .A2(\SB4_31/i0[10] ), .A3(
        \SB4_31/i0[9] ), .ZN(n3732) );
  NAND3_X1 U4829 ( .A1(\SB4_20/i0_4 ), .A2(\SB4_20/i1[9] ), .A3(\SB4_20/i1_5 ), 
        .ZN(n6393) );
  NAND3_X1 U4831 ( .A1(\SB4_27/i0[10] ), .A2(\SB4_27/i1[9] ), .A3(
        \SB4_27/i1_7 ), .ZN(\SB4_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4833 ( .A1(n1494), .A2(\SB4_24/i0[7] ), .A3(\SB4_24/i0[6] ), .ZN(
        n7531) );
  NAND2_X1 U4834 ( .A1(\SB4_24/i0_0 ), .A2(\SB4_24/i3[0] ), .ZN(
        \SB4_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4836 ( .A1(\SB4_13/i0[9] ), .A2(\SB4_13/i0[6] ), .A3(\SB4_13/i0_4 ), .ZN(n792) );
  NAND3_X1 U4841 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i0_4 ), .A3(\SB4_30/i0_3 ), .ZN(n6212) );
  NAND3_X1 U4849 ( .A1(\SB4_31/i0_3 ), .A2(\SB4_31/i0_4 ), .A3(\SB4_31/i0_0 ), 
        .ZN(n3374) );
  NOR2_X1 U4852 ( .A1(\RI3[0][97] ), .A2(\RI3[0][99] ), .ZN(n5434) );
  AND2_X1 U4855 ( .A1(\SB1_0_10/i0[6] ), .A2(\SB1_0_10/i0_3 ), .Z(n5435) );
  AND2_X1 U4857 ( .A1(\SB1_0_10/i1_5 ), .A2(\SB1_0_10/i1[9] ), .Z(n5436) );
  OR2_X1 U4858 ( .A1(n4398), .A2(\SB2_3_8/i0_3 ), .Z(n5437) );
  AND2_X1 U4862 ( .A1(n6710), .A2(\SB1_2_27/Component_Function_4/NAND4_in[1] ), 
        .Z(n5439) );
  AND4_X2 U4865 ( .A1(n2533), .A2(n4830), .A3(
        \SB1_3_20/Component_Function_5/NAND4_in[0] ), .A4(n4020), .Z(n5440) );
  INV_X2 U4868 ( .I(n2592), .ZN(\SB2_0_1/i0[9] ) );
  XNOR2_X1 U4869 ( .A1(\MC_ARK_ARC_1_2/temp5[3] ), .A2(
        \MC_ARK_ARC_1_2/temp6[3] ), .ZN(n5441) );
  AND4_X2 U4871 ( .A1(\SB3_1/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_1/Component_Function_5/NAND4_in[2] ), .A3(n2627), .A4(
        \SB3_1/Component_Function_5/NAND4_in[0] ), .Z(n5442) );
  AND4_X2 U4873 ( .A1(\SB1_4_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_4_27/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_4_27/Component_Function_2/NAND4_in[1] ), .A4(n3069), .Z(n5443) );
  OR2_X2 U4877 ( .A1(n7200), .A2(n4838), .Z(n5444) );
  INV_X1 U4878 ( .I(\SB3_22/buf_output[2] ), .ZN(\SB4_19/i1[9] ) );
  NAND4_X2 U4879 ( .A1(n5253), .A2(n6736), .A3(
        \SB1_3_9/Component_Function_5/NAND4_in[2] ), .A4(n5445), .ZN(
        \SB1_3_9/buf_output[5] ) );
  NAND2_X2 U4880 ( .A1(\SB1_3_9/i0_0 ), .A2(\SB1_3_9/i3[0] ), .ZN(n5445) );
  NAND4_X2 U4881 ( .A1(\SB3_16/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_16/Component_Function_5/NAND4_in[1] ), .A3(n5848), .A4(
        \SB3_16/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_16/buf_output[5] ) );
  XOR2_X1 U4883 ( .A1(\MC_ARK_ARC_1_2/temp5[132] ), .A2(
        \MC_ARK_ARC_1_2/temp6[132] ), .Z(\MC_ARK_ARC_1_2/buf_output[132] ) );
  XOR2_X1 U4884 ( .A1(\MC_ARK_ARC_1_2/temp1[132] ), .A2(
        \MC_ARK_ARC_1_2/temp2[132] ), .Z(\MC_ARK_ARC_1_2/temp5[132] ) );
  XOR2_X1 U4886 ( .A1(n6501), .A2(n6500), .Z(\MC_ARK_ARC_1_2/buf_output[175] )
         );
  INV_X1 U4888 ( .I(\SB1_3_26/buf_output[1] ), .ZN(\SB2_3_22/i1_7 ) );
  NAND4_X2 U4891 ( .A1(\SB1_3_26/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_26/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_3_26/Component_Function_1/NAND4_in[0] ), .A4(n4729), .ZN(
        \SB1_3_26/buf_output[1] ) );
  INV_X1 U4895 ( .I(\SB3_31/buf_output[2] ), .ZN(\SB4_28/i1[9] ) );
  NAND4_X2 U4898 ( .A1(\SB3_31/Component_Function_2/NAND4_in[1] ), .A2(n6692), 
        .A3(\SB3_31/Component_Function_2/NAND4_in[2] ), .A4(n6417), .ZN(
        \SB3_31/buf_output[2] ) );
  XOR2_X1 U4900 ( .A1(\MC_ARK_ARC_1_2/temp1[19] ), .A2(
        \MC_ARK_ARC_1_2/temp2[19] ), .Z(\MC_ARK_ARC_1_2/temp5[19] ) );
  XOR2_X1 U4906 ( .A1(\MC_ARK_ARC_1_3/temp4[13] ), .A2(n5446), .Z(
        \MC_ARK_ARC_1_3/temp6[13] ) );
  XOR2_X1 U4907 ( .A1(\RI5[3][79] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[115] ), 
        .Z(n5446) );
  NAND4_X2 U4909 ( .A1(\SB1_4_29/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_4_29/Component_Function_1/NAND4_in[3] ), .A3(n5826), .A4(
        \SB1_4_29/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_4_29/buf_output[1] ) );
  NAND4_X2 U4910 ( .A1(\SB3_17/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_17/Component_Function_0/NAND4_in[1] ), .A3(n3782), .A4(
        \SB3_17/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_17/buf_output[0] ) );
  XOR2_X1 U4911 ( .A1(\MC_ARK_ARC_1_1/temp1[188] ), .A2(n5447), .Z(n7028) );
  XOR2_X1 U4913 ( .A1(\RI5[1][134] ), .A2(\RI5[1][158] ), .Z(n5447) );
  NAND3_X1 U4914 ( .A1(\SB4_12/i3[0] ), .A2(\SB4_12/i0[8] ), .A3(\SB4_12/i1_5 ), .ZN(n1255) );
  BUF_X4 U4916 ( .I(\MC_ARK_ARC_1_3/buf_output[39] ), .Z(\SB1_4_25/i0[10] ) );
  CLKBUF_X4 U4917 ( .I(\SB1_4_25/buf_output[3] ), .Z(\SB2_4_23/i0[10] ) );
  NAND3_X2 U4921 ( .A1(\SB2_2_25/i0[6] ), .A2(\SB2_2_25/i0[10] ), .A3(
        \SB2_2_25/i0_0 ), .ZN(\SB2_2_25/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U4922 ( .A1(\SB1_3_20/i0_0 ), .A2(\SB1_3_20/i0_3 ), .A3(
        \SB1_3_20/i0_4 ), .ZN(n5554) );
  XOR2_X1 U4923 ( .A1(\RI5[4][41] ), .A2(\RI5[4][65] ), .Z(n5542) );
  NAND3_X2 U4924 ( .A1(\SB2_4_14/i0[9] ), .A2(\SB2_4_14/i0_4 ), .A3(
        \SB2_4_14/i0[6] ), .ZN(n7167) );
  NAND2_X2 U4926 ( .A1(n5831), .A2(n7091), .ZN(\SB2_3_7/i0_4 ) );
  XOR2_X1 U4928 ( .A1(\RI5[0][50] ), .A2(\RI5[0][98] ), .Z(n4402) );
  XOR2_X1 U4929 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[143] ), .A2(\RI5[3][11] ), 
        .Z(n6074) );
  NAND4_X2 U4930 ( .A1(n5024), .A2(n3135), .A3(
        \SB2_4_20/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_4_20/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_4_20/buf_output[5] ) );
  NAND3_X2 U4933 ( .A1(\SB2_4_22/i0_0 ), .A2(\SB2_4_22/i0[10] ), .A3(
        \SB2_4_22/i0[6] ), .ZN(\SB2_4_22/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U4935 ( .A1(\SB1_2_11/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_11/Component_Function_1/NAND4_in[0] ), .A3(n3276), .A4(
        \SB1_2_11/Component_Function_1/NAND4_in[1] ), .ZN(
        \SB1_2_11/buf_output[1] ) );
  NAND4_X2 U4936 ( .A1(\SB2_2_4/Component_Function_3/NAND4_in[2] ), .A2(n6622), 
        .A3(\SB2_2_4/Component_Function_3/NAND4_in[3] ), .A4(n5448), .ZN(
        \SB2_2_4/buf_output[3] ) );
  NAND3_X2 U4937 ( .A1(\SB2_2_4/i0_0 ), .A2(\SB2_2_4/i0_3 ), .A3(
        \SB2_2_4/i0_4 ), .ZN(n5448) );
  NAND3_X2 U4938 ( .A1(\SB3_9/i0_0 ), .A2(\SB3_9/i1_5 ), .A3(\SB3_9/i0_4 ), 
        .ZN(n7338) );
  NAND3_X1 U4940 ( .A1(\SB2_4_25/i0_4 ), .A2(\SB2_4_25/i1_5 ), .A3(
        \SB2_4_25/i1[9] ), .ZN(n744) );
  XOR2_X1 U4941 ( .A1(n3701), .A2(n5449), .Z(n2976) );
  XOR2_X1 U4942 ( .A1(\RI5[4][38] ), .A2(\RI5[4][8] ), .Z(n5449) );
  BUF_X2 U4943 ( .I(\SB2_0_31/i3[0] ), .Z(n5450) );
  XOR2_X1 U4946 ( .A1(n5451), .A2(n166), .Z(Ciphertext[68]) );
  NAND4_X2 U4947 ( .A1(n6707), .A2(\SB4_20/Component_Function_2/NAND4_in[0] ), 
        .A3(n1457), .A4(n4863), .ZN(n5451) );
  XOR2_X1 U4950 ( .A1(n5452), .A2(\MC_ARK_ARC_1_3/temp4[31] ), .Z(
        \MC_ARK_ARC_1_3/temp6[31] ) );
  XOR2_X1 U4953 ( .A1(\RI5[3][97] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[133] ), 
        .Z(n5452) );
  NAND4_X2 U4959 ( .A1(\SB2_2_4/Component_Function_4/NAND4_in[1] ), .A2(n5413), 
        .A3(\SB2_2_4/Component_Function_4/NAND4_in[2] ), .A4(n5453), .ZN(
        \SB2_2_4/buf_output[4] ) );
  NAND4_X2 U4961 ( .A1(\SB1_2_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_4/NAND4_in[2] ), .A4(n5454), .ZN(
        \SB1_2_29/buf_output[4] ) );
  NAND4_X2 U4963 ( .A1(\SB2_4_14/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_4_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_14/Component_Function_1/NAND4_in[2] ), .A4(n5455), .ZN(
        \SB2_4_14/buf_output[1] ) );
  NAND2_X1 U4967 ( .A1(\SB2_4_14/i0_3 ), .A2(\SB2_4_14/i1[9] ), .ZN(n5455) );
  INV_X1 U4971 ( .I(\RI3[0][131] ), .ZN(\SB2_0_10/i1_5 ) );
  NAND3_X2 U4978 ( .A1(n4803), .A2(\SB1_0_10/Component_Function_5/NAND4_in[1] ), .A3(n3357), .ZN(\RI3[0][131] ) );
  NAND4_X2 U4982 ( .A1(n3041), .A2(\SB2_4_13/Component_Function_5/NAND4_in[0] ), .A3(n5457), .A4(n5456), .ZN(\SB2_4_13/buf_output[5] ) );
  NAND3_X2 U4985 ( .A1(\SB2_4_13/i0_0 ), .A2(\SB2_4_13/i0[10] ), .A3(
        \SB2_4_13/i0[6] ), .ZN(n5456) );
  NAND3_X1 U4986 ( .A1(\SB2_4_13/i0[9] ), .A2(\SB1_4_14/buf_output[4] ), .A3(
        \SB2_4_13/i0[6] ), .ZN(n5457) );
  INV_X1 U4988 ( .I(\SB3_10/buf_output[5] ), .ZN(\SB4_10/i1_5 ) );
  NAND4_X2 U4993 ( .A1(\SB3_10/Component_Function_5/NAND4_in[1] ), .A2(n5366), 
        .A3(n5519), .A4(\SB3_10/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_10/buf_output[5] ) );
  XOR2_X1 U4994 ( .A1(n5459), .A2(n5458), .Z(n6626) );
  XOR2_X1 U4995 ( .A1(\RI5[2][173] ), .A2(n529), .Z(n5458) );
  XOR2_X1 U5000 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[23] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[179] ), .Z(n5459) );
  NAND4_X2 U5009 ( .A1(\SB2_3_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_29/Component_Function_4/NAND4_in[3] ), .A3(n4027), .A4(n5460), 
        .ZN(\SB2_3_29/buf_output[4] ) );
  XOR2_X1 U5012 ( .A1(n5461), .A2(n220), .Z(Ciphertext[100]) );
  NAND4_X2 U5014 ( .A1(n2824), .A2(n7526), .A3(
        \SB4_15/Component_Function_4/NAND4_in[0] ), .A4(
        \SB4_15/Component_Function_4/NAND4_in[3] ), .ZN(n5461) );
  XOR2_X1 U5015 ( .A1(\MC_ARK_ARC_1_4/temp6[127] ), .A2(n5462), .Z(
        \MC_ARK_ARC_1_4/buf_output[127] ) );
  XOR2_X1 U5017 ( .A1(\MC_ARK_ARC_1_4/temp1[127] ), .A2(n2332), .Z(n5462) );
  NAND3_X1 U5018 ( .A1(\SB2_0_8/i0[10] ), .A2(\RI3[0][142] ), .A3(
        \SB2_0_8/i0_3 ), .ZN(\SB2_0_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U5019 ( .A1(\SB2_4_6/i0_3 ), .A2(\SB2_4_6/i1_7 ), .A3(
        \SB2_4_6/i0[8] ), .ZN(\SB2_4_6/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U5020 ( .A1(\SB2_3_10/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_3_10/Component_Function_3/NAND4_in[0] ), .A3(n2405), .A4(n5463), 
        .ZN(\SB2_3_10/buf_output[3] ) );
  NAND3_X2 U5024 ( .A1(n851), .A2(\SB2_3_10/i0_3 ), .A3(\SB2_3_10/i0_0 ), .ZN(
        n5463) );
  XOR2_X1 U5025 ( .A1(\MC_ARK_ARC_1_2/temp3[152] ), .A2(n5464), .Z(n3388) );
  XOR2_X1 U5028 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), .A2(\RI5[2][152] ), 
        .Z(n5464) );
  NAND4_X2 U5029 ( .A1(n2570), .A2(\SB2_1_13/Component_Function_5/NAND4_in[0] ), .A3(n6447), .A4(n5465), .ZN(\SB2_1_13/buf_output[5] ) );
  NAND3_X2 U5031 ( .A1(\SB2_1_13/i0_4 ), .A2(\SB2_1_13/i0[6] ), .A3(
        \SB2_1_13/i0[9] ), .ZN(n5465) );
  XOR2_X1 U5037 ( .A1(n5467), .A2(n5466), .Z(\MC_ARK_ARC_1_0/buf_output[81] )
         );
  XOR2_X1 U5039 ( .A1(\MC_ARK_ARC_1_0/temp3[81] ), .A2(
        \MC_ARK_ARC_1_0/temp4[81] ), .Z(n5466) );
  XOR2_X1 U5040 ( .A1(\MC_ARK_ARC_1_0/temp2[81] ), .A2(n2487), .Z(n5467) );
  XOR2_X1 U5045 ( .A1(\MC_ARK_ARC_1_1/temp2[119] ), .A2(n5468), .Z(
        \MC_ARK_ARC_1_1/temp5[119] ) );
  XOR2_X1 U5046 ( .A1(\RI5[1][119] ), .A2(\RI5[1][113] ), .Z(n5468) );
  XOR2_X1 U5049 ( .A1(n5502), .A2(\MC_ARK_ARC_1_0/temp1[88] ), .Z(
        \MC_ARK_ARC_1_0/temp5[88] ) );
  XOR2_X1 U5050 ( .A1(\RI5[0][34] ), .A2(\SB2_0_31/buf_output[4] ), .Z(n5898)
         );
  XOR2_X1 U5051 ( .A1(\MC_ARK_ARC_1_4/temp1[175] ), .A2(
        \MC_ARK_ARC_1_4/temp2[175] ), .Z(\MC_ARK_ARC_1_4/temp5[175] ) );
  NAND3_X2 U5056 ( .A1(\SB2_0_2/i0[10] ), .A2(\SB2_0_2/i1_7 ), .A3(
        \SB2_0_2/i1[9] ), .ZN(\SB2_0_2/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U5057 ( .A1(n2534), .A2(n5469), .Z(n3274) );
  XOR2_X1 U5067 ( .A1(\RI5[0][189] ), .A2(\RI5[0][21] ), .Z(n5469) );
  NAND4_X2 U5068 ( .A1(n3102), .A2(n2410), .A3(n3602), .A4(n5470), .ZN(
        \SB2_4_16/buf_output[5] ) );
  NAND3_X2 U5074 ( .A1(\SB2_4_16/i0_0 ), .A2(\SB2_4_16/i0[10] ), .A3(
        \SB2_4_16/i0[6] ), .ZN(n5470) );
  XOR2_X1 U5082 ( .A1(n5472), .A2(n5471), .Z(n5907) );
  XOR2_X1 U5084 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[92] ), .A2(n485), .Z(n5471) );
  XOR2_X1 U5085 ( .A1(\RI5[2][134] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[98] ), 
        .Z(n5472) );
  XOR2_X1 U5090 ( .A1(n5473), .A2(n2776), .Z(\MC_ARK_ARC_1_0/buf_output[102] )
         );
  XOR2_X1 U5093 ( .A1(n5866), .A2(n1927), .Z(n5473) );
  NAND4_X2 U5094 ( .A1(\SB1_2_9/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_9/Component_Function_3/NAND4_in[0] ), .A3(n6999), .A4(n5474), 
        .ZN(\SB1_2_9/buf_output[3] ) );
  INV_X2 U5095 ( .I(\SB1_3_20/buf_output[3] ), .ZN(\SB2_3_18/i0[8] ) );
  NAND4_X2 U5098 ( .A1(\SB1_3_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_20/Component_Function_3/NAND4_in[2] ), .A3(n5554), .A4(
        \SB1_3_20/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_20/buf_output[3] ) );
  NAND4_X2 U5099 ( .A1(n2993), .A2(\SB2_4_14/Component_Function_5/NAND4_in[0] ), .A3(n7167), .A4(n5475), .ZN(\SB2_4_14/buf_output[5] ) );
  NAND3_X2 U5109 ( .A1(\SB2_4_14/i0[10] ), .A2(\SB2_4_14/i0[6] ), .A3(
        \SB2_4_14/i0_0 ), .ZN(n5475) );
  XOR2_X1 U5110 ( .A1(n5477), .A2(n5476), .Z(n2480) );
  XOR2_X1 U5111 ( .A1(\RI5[0][20] ), .A2(\RI5[0][164] ), .Z(n5476) );
  XOR2_X1 U5112 ( .A1(\RI5[0][26] ), .A2(\RI5[0][188] ), .Z(n5477) );
  NAND4_X2 U5113 ( .A1(n4565), .A2(n6941), .A3(n4121), .A4(n5478), .ZN(
        \SB1_2_22/buf_output[3] ) );
  NAND3_X2 U5114 ( .A1(\SB1_2_22/i1_7 ), .A2(\SB1_2_22/i0[10] ), .A3(
        \SB1_2_22/i1[9] ), .ZN(n5478) );
  NAND4_X2 U5117 ( .A1(n5235), .A2(\SB3_28/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB3_28/Component_Function_5/NAND4_in[0] ), .A4(n5479), .ZN(
        \SB3_28/buf_output[5] ) );
  INV_X2 U5118 ( .I(\MC_ARK_ARC_1_3/buf_output[93] ), .ZN(\SB1_4_16/i0[8] ) );
  INV_X8 U5120 ( .I(n5480), .ZN(\RI1[4][155] ) );
  INV_X2 U5121 ( .I(\MC_ARK_ARC_1_3/buf_output[155] ), .ZN(n5480) );
  INV_X4 U5125 ( .I(n5481), .ZN(\SB1_0_27/i1[9] ) );
  BUF_X2 U5126 ( .I(n262), .Z(n5481) );
  NAND3_X2 U5127 ( .A1(\SB2_0_29/i0_3 ), .A2(\SB2_0_29/i0[8] ), .A3(
        \SB2_0_29/i1_7 ), .ZN(\SB2_0_29/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U5129 ( .A1(n5482), .A2(n85), .Z(Ciphertext[9]) );
  NAND4_X2 U5133 ( .A1(n3769), .A2(\SB4_30/Component_Function_3/NAND4_in[2] ), 
        .A3(n5546), .A4(\SB4_30/Component_Function_3/NAND4_in[3] ), .ZN(n5482)
         );
  XOR2_X1 U5137 ( .A1(\MC_ARK_ARC_1_1/temp4[179] ), .A2(n6760), .Z(n5915) );
  NAND4_X2 U5138 ( .A1(\SB3_7/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_7/Component_Function_4/NAND4_in[0] ), .A3(n5720), .A4(n4190), 
        .ZN(\SB3_7/buf_output[4] ) );
  NAND4_X2 U5139 ( .A1(\SB2_0_13/Component_Function_3/NAND4_in[0] ), .A2(n1835), .A3(n5552), .A4(\SB2_0_13/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_0_13/buf_output[3] ) );
  NAND4_X2 U5140 ( .A1(n3287), .A2(\SB2_1_10/Component_Function_5/NAND4_in[1] ), .A3(n2059), .A4(\SB2_1_10/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_10/buf_output[5] ) );
  NAND4_X1 U5145 ( .A1(\SB1_0_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_1/NAND4_in[1] ), .A3(n6553), .A4(
        \SB1_0_27/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_0_27/buf_output[1] ) );
  XOR2_X1 U5146 ( .A1(\RI5[0][123] ), .A2(\RI5[0][99] ), .Z(n4183) );
  CLKBUF_X12 U5149 ( .I(\MC_ARK_ARC_1_4/buf_output[122] ), .Z(n6243) );
  NAND4_X2 U5150 ( .A1(\SB3_3/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_3/Component_Function_2/NAND4_in[3] ), .A3(n4966), .A4(n5483), 
        .ZN(\SB3_3/buf_output[2] ) );
  NAND3_X2 U5156 ( .A1(\SB3_3/i0[10] ), .A2(\SB3_3/i0[6] ), .A3(\SB3_3/i0_3 ), 
        .ZN(n5483) );
  NAND4_X2 U5158 ( .A1(\SB2_2_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_12/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_12/Component_Function_5/NAND4_in[0] ), .A4(n5484), .ZN(
        \SB2_2_12/buf_output[5] ) );
  NAND3_X2 U5162 ( .A1(\SB2_2_12/i0[6] ), .A2(\SB2_2_12/i0_4 ), .A3(
        \SB2_2_12/i0[9] ), .ZN(n5484) );
  XOR2_X1 U5166 ( .A1(n5485), .A2(n136), .Z(Ciphertext[146]) );
  NAND4_X2 U5169 ( .A1(n5367), .A2(n7066), .A3(n5730), .A4(
        \SB4_7/Component_Function_2/NAND4_in[2] ), .ZN(n5485) );
  XOR2_X1 U5170 ( .A1(n5487), .A2(n5486), .Z(n4687) );
  XOR2_X1 U5171 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[183] ), .A2(n540), .Z(
        n5486) );
  XOR2_X1 U5173 ( .A1(\RI5[2][117] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[147] ), 
        .Z(n5487) );
  XOR2_X1 U5174 ( .A1(\MC_ARK_ARC_1_1/temp6[107] ), .A2(n961), .Z(
        \MC_ARK_ARC_1_1/buf_output[107] ) );
  XOR2_X1 U5177 ( .A1(n6456), .A2(n6455), .Z(\MC_ARK_ARC_1_1/temp6[107] ) );
  XOR2_X1 U5178 ( .A1(\RI5[0][73] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[97] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[127] ) );
  NAND4_X2 U5181 ( .A1(\SB2_3_5/Component_Function_5/NAND4_in[2] ), .A2(n2955), 
        .A3(\SB2_3_5/Component_Function_5/NAND4_in[0] ), .A4(n5488), .ZN(
        \SB2_3_5/buf_output[5] ) );
  NAND3_X2 U5189 ( .A1(\SB2_3_5/i0[6] ), .A2(\SB2_3_5/i0[10] ), .A3(
        \SB2_3_5/i0_0 ), .ZN(n5488) );
  NAND3_X1 U5193 ( .A1(\SB3_4/i0_3 ), .A2(\MC_ARK_ARC_1_4/buf_output[162] ), 
        .A3(\SB3_4/i0[8] ), .ZN(\SB3_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U5203 ( .A1(n590), .A2(\SB2_1_0/i1[9] ), .A3(\SB2_1_0/i1_5 ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[3] ) );
  INV_X2 U5205 ( .I(\SB1_0_21/buf_output[2] ), .ZN(\SB2_0_18/i1[9] ) );
  NAND4_X2 U5209 ( .A1(\SB1_0_21/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_21/Component_Function_2/NAND4_in[2] ), .A3(n4406), .A4(n5122), 
        .ZN(\SB1_0_21/buf_output[2] ) );
  NAND4_X2 U5217 ( .A1(n2894), .A2(\SB2_4_27/Component_Function_5/NAND4_in[0] ), .A3(n5107), .A4(n5489), .ZN(\SB2_4_27/buf_output[5] ) );
  NAND3_X2 U5225 ( .A1(\SB2_4_27/i0[6] ), .A2(\SB2_4_27/i0[10] ), .A3(
        \SB2_4_27/i0_0 ), .ZN(n5489) );
  XOR2_X1 U5230 ( .A1(n5490), .A2(n52), .Z(Ciphertext[180]) );
  NAND4_X2 U5233 ( .A1(\SB4_1/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_1/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_1/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_1/Component_Function_0/NAND4_in[0] ), .ZN(n5490) );
  NAND3_X1 U5235 ( .A1(\SB4_31/i0_3 ), .A2(\SB4_31/i0[8] ), .A3(\SB4_31/i0[9] ), .ZN(n5254) );
  XOR2_X1 U5238 ( .A1(n5492), .A2(n5491), .Z(n6213) );
  XOR2_X1 U5243 ( .A1(\RI5[2][59] ), .A2(n149), .Z(n5491) );
  XOR2_X1 U5244 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[23] ), .A2(\RI5[2][17] ), 
        .Z(n5492) );
  NAND4_X2 U5246 ( .A1(\SB2_2_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_22/Component_Function_5/NAND4_in[1] ), .A3(n5147), .A4(n5493), 
        .ZN(\SB2_2_22/buf_output[5] ) );
  NAND3_X2 U5247 ( .A1(\SB2_2_22/i0[6] ), .A2(\SB2_2_22/i0[9] ), .A3(
        \SB2_2_22/i0_4 ), .ZN(n5493) );
  NAND4_X2 U5248 ( .A1(\SB2_4_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_11/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_4_11/Component_Function_2/NAND4_in[1] ), .A4(n5494), .ZN(
        \SB2_4_11/buf_output[2] ) );
  NAND3_X2 U5249 ( .A1(\SB2_4_11/i0_4 ), .A2(\SB2_4_11/i0_0 ), .A3(
        \SB2_4_11/i1_5 ), .ZN(n5494) );
  XOR2_X1 U5253 ( .A1(n5495), .A2(n58), .Z(Ciphertext[3]) );
  NAND4_X2 U5257 ( .A1(n7550), .A2(\SB4_31/Component_Function_3/NAND4_in[2] ), 
        .A3(n7248), .A4(n3374), .ZN(n5495) );
  INV_X2 U5261 ( .I(\SB1_4_24/buf_output[2] ), .ZN(\SB2_4_21/i1[9] ) );
  NAND4_X2 U5264 ( .A1(\SB1_4_24/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_4_24/Component_Function_2/NAND4_in[3] ), .A3(n6096), .A4(
        \SB1_4_24/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_4_24/buf_output[2] ) );
  NAND4_X2 U5265 ( .A1(\SB2_1_26/Component_Function_0/NAND4_in[1] ), .A2(n6306), .A3(n2046), .A4(n5496), .ZN(\SB2_1_26/buf_output[0] ) );
  NAND4_X2 U5268 ( .A1(\SB2_3_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_14/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_14/Component_Function_5/NAND4_in[0] ), .A4(n5497), .ZN(
        \SB2_3_14/buf_output[5] ) );
  NAND3_X2 U5270 ( .A1(\SB2_3_14/i0[10] ), .A2(\SB2_3_14/i0[6] ), .A3(
        \SB2_3_14/i0_0 ), .ZN(n5497) );
  XOR2_X1 U5275 ( .A1(n5498), .A2(n29), .Z(Ciphertext[0]) );
  NAND4_X2 U5280 ( .A1(\SB4_31/Component_Function_0/NAND4_in[1] ), .A2(n7404), 
        .A3(\SB4_31/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_31/Component_Function_0/NAND4_in[2] ), .ZN(n5498) );
  NAND4_X2 U5283 ( .A1(\SB1_0_30/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_30/Component_Function_3/NAND4_in[2] ), .A3(n6085), .A4(n5499), 
        .ZN(\RI3[0][21] ) );
  NAND3_X1 U5284 ( .A1(\SB1_0_30/i0_4 ), .A2(\SB1_0_30/i0_0 ), .A3(
        \SB1_0_30/i0_3 ), .ZN(n5499) );
  XOR2_X1 U5293 ( .A1(n5500), .A2(n194), .Z(Ciphertext[185]) );
  NAND4_X2 U5294 ( .A1(\SB4_1/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_1/Component_Function_5/NAND4_in[1] ), .A3(n4682), .A4(
        \SB4_1/Component_Function_5/NAND4_in[0] ), .ZN(n5500) );
  XOR2_X1 U5295 ( .A1(n5501), .A2(n69), .Z(Ciphertext[184]) );
  NAND4_X2 U5296 ( .A1(\SB4_1/Component_Function_4/NAND4_in[3] ), .A2(n2562), 
        .A3(n4919), .A4(\SB4_1/Component_Function_4/NAND4_in[0] ), .ZN(n5501)
         );
  XOR2_X1 U5302 ( .A1(\RI5[0][58] ), .A2(\RI5[0][34] ), .Z(n5502) );
  XOR2_X1 U5306 ( .A1(\RI5[0][14] ), .A2(\SB2_0_26/buf_output[2] ), .Z(n6554)
         );
  XOR2_X1 U5307 ( .A1(n5503), .A2(n205), .Z(Ciphertext[188]) );
  NAND4_X2 U5311 ( .A1(\SB4_0/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_0/Component_Function_2/NAND4_in[0] ), .A3(
        \SB4_0/Component_Function_2/NAND4_in[1] ), .A4(n6007), .ZN(n5503) );
  XOR2_X1 U5312 ( .A1(n5505), .A2(n5504), .Z(\MC_ARK_ARC_1_4/buf_output[163] )
         );
  XOR2_X1 U5315 ( .A1(\MC_ARK_ARC_1_4/temp1[163] ), .A2(
        \MC_ARK_ARC_1_4/temp4[163] ), .Z(n5504) );
  XOR2_X1 U5325 ( .A1(\MC_ARK_ARC_1_4/temp2[163] ), .A2(
        \MC_ARK_ARC_1_4/temp3[163] ), .Z(n5505) );
  NAND4_X2 U5328 ( .A1(\SB1_2_19/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_19/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_2_19/Component_Function_1/NAND4_in[0] ), .A4(n5506), .ZN(
        \RI3[2][97] ) );
  NAND3_X2 U5330 ( .A1(\SB1_2_19/i0_3 ), .A2(\SB1_2_19/i0[8] ), .A3(
        \SB1_2_19/i1_7 ), .ZN(n5506) );
  NAND4_X2 U5337 ( .A1(\SB2_0_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_23/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_23/Component_Function_3/NAND4_in[1] ), .A4(n5507), .ZN(
        \SB2_0_23/buf_output[3] ) );
  NAND3_X2 U5339 ( .A1(\SB2_0_23/i3[0] ), .A2(\SB2_0_23/i0[8] ), .A3(
        \SB2_0_23/i1_5 ), .ZN(n5507) );
  XOR2_X1 U5344 ( .A1(n5508), .A2(n175), .Z(Ciphertext[176]) );
  NAND4_X2 U5348 ( .A1(\SB4_2/Component_Function_2/NAND4_in[0] ), .A2(n5888), 
        .A3(\SB4_2/Component_Function_2/NAND4_in[3] ), .A4(
        \SB4_2/Component_Function_2/NAND4_in[1] ), .ZN(n5508) );
  XOR2_X1 U5349 ( .A1(\RI5[1][12] ), .A2(\RI5[1][18] ), .Z(
        \MC_ARK_ARC_1_1/temp1[18] ) );
  XOR2_X1 U5350 ( .A1(n5591), .A2(n5509), .Z(\MC_ARK_ARC_1_2/buf_output[158] )
         );
  XOR2_X1 U5355 ( .A1(\MC_ARK_ARC_1_2/temp4[158] ), .A2(n5667), .Z(n5509) );
  XOR2_X1 U5357 ( .A1(n6560), .A2(n5510), .Z(\MC_ARK_ARC_1_0/buf_output[27] )
         );
  XOR2_X1 U5358 ( .A1(\MC_ARK_ARC_1_0/temp4[27] ), .A2(n6588), .Z(n5510) );
  XOR2_X1 U5360 ( .A1(\MC_ARK_ARC_1_2/temp2[56] ), .A2(n5511), .Z(n6361) );
  XOR2_X1 U5364 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[122] ), .A2(\RI5[2][158] ), 
        .Z(n5511) );
  XOR2_X1 U5365 ( .A1(n3096), .A2(n5321), .Z(\MC_ARK_ARC_1_1/buf_output[176] )
         );
  XOR2_X1 U5366 ( .A1(\MC_ARK_ARC_1_1/temp3[176] ), .A2(
        \MC_ARK_ARC_1_1/temp4[176] ), .Z(n3096) );
  NAND3_X2 U5368 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0[10] ), .A3(
        \SB2_1_23/i0_4 ), .ZN(n4454) );
  NAND4_X2 U5369 ( .A1(\SB2_3_27/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_27/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_3_27/Component_Function_1/NAND4_in[1] ), .A4(n5512), .ZN(
        \SB2_3_27/buf_output[1] ) );
  NAND2_X2 U5370 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i1[9] ), .ZN(n5512) );
  INV_X2 U5372 ( .I(\SB1_1_21/buf_output[2] ), .ZN(\SB2_1_18/i1[9] ) );
  NAND4_X2 U5373 ( .A1(n3083), .A2(\SB1_1_21/Component_Function_2/NAND4_in[1] ), .A3(\SB1_1_21/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_21/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_1_21/buf_output[2] ) );
  NAND4_X2 U5375 ( .A1(\SB3_2/Component_Function_3/NAND4_in[0] ), .A2(n1080), 
        .A3(n6915), .A4(n5513), .ZN(\SB3_2/buf_output[3] ) );
  NAND3_X2 U5378 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i0_0 ), .A3(\SB3_2/i0_4 ), 
        .ZN(n5513) );
  XOR2_X1 U5380 ( .A1(\MC_ARK_ARC_1_1/temp1[140] ), .A2(
        \MC_ARK_ARC_1_1/temp2[140] ), .Z(n5723) );
  NAND3_X2 U5384 ( .A1(\SB1_2_22/i0_4 ), .A2(\SB1_2_22/i1[9] ), .A3(
        \RI1[2][59] ), .ZN(\SB1_2_22/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U5388 ( .A1(\SB2_2_15/i0[9] ), .A2(\SB2_2_15/i0_3 ), .A3(
        \SB2_2_15/i0[8] ), .ZN(\SB2_2_15/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U5389 ( .A1(\SB1_3_26/Component_Function_2/NAND4_in[1] ), .A2(n6864), .A3(\SB1_3_26/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_3_26/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_3_26/buf_output[2] ) );
  NAND4_X2 U5391 ( .A1(\SB1_1_18/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_18/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_1_18/Component_Function_2/NAND4_in[0] ), .A4(n887), .ZN(
        \SB1_1_18/buf_output[2] ) );
  NAND3_X2 U5392 ( .A1(\SB1_3_30/i0[10] ), .A2(\SB1_3_30/i1[9] ), .A3(
        \SB1_3_30/i1_5 ), .ZN(n6296) );
  NAND3_X1 U5393 ( .A1(\SB2_1_23/i0[6] ), .A2(\SB1_1_28/buf_output[0] ), .A3(
        \SB2_1_23/i1_5 ), .ZN(\SB2_1_23/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U5397 ( .A1(\RI5[3][161] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[5] ), 
        .Z(n2831) );
  XOR2_X1 U5398 ( .A1(\RI5[2][116] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[164] ), 
        .Z(n3951) );
  NAND4_X2 U5399 ( .A1(\SB1_4_2/Component_Function_5/NAND4_in[2] ), .A2(n4431), 
        .A3(n5550), .A4(\SB1_4_2/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_4_2/buf_output[5] ) );
  XOR2_X1 U5413 ( .A1(\RI5[0][26] ), .A2(\RI5[0][50] ), .Z(n2702) );
  NAND4_X2 U5414 ( .A1(\SB2_2_26/Component_Function_5/NAND4_in[2] ), .A2(n6614), .A3(n5553), .A4(\SB2_2_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_26/buf_output[5] ) );
  XOR2_X1 U5415 ( .A1(\MC_ARK_ARC_1_1/temp6[164] ), .A2(n5514), .Z(
        \MC_ARK_ARC_1_1/buf_output[164] ) );
  XOR2_X1 U5417 ( .A1(\MC_ARK_ARC_1_1/temp1[164] ), .A2(
        \MC_ARK_ARC_1_1/temp2[164] ), .Z(n5514) );
  NAND4_X2 U5418 ( .A1(\SB1_3_12/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_12/Component_Function_3/NAND4_in[0] ), .A3(n6678), .A4(
        \SB1_3_12/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_12/buf_output[3] ) );
  NAND4_X2 U5424 ( .A1(\SB1_4_12/Component_Function_2/NAND4_in[0] ), .A2(n4205), .A3(n1483), .A4(\SB1_4_12/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB1_4_12/buf_output[2] ) );
  NAND3_X2 U5426 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0_4 ), .A3(
        \SB2_2_12/i1[9] ), .ZN(\SB2_2_12/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U5451 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[58] ), .A2(\RI5[1][82] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[112] ) );
  NAND3_X2 U5457 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i0_4 ), .A3(
        \SB2_1_15/i1[9] ), .ZN(\SB2_1_15/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U5459 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[58] ), .A2(\RI5[1][52] ), 
        .Z(n5884) );
  NAND4_X2 U5460 ( .A1(\SB1_3_27/Component_Function_5/NAND4_in[1] ), .A2(n4538), .A3(\SB1_3_27/Component_Function_5/NAND4_in[0] ), .A4(n6434), .ZN(
        \SB1_3_27/buf_output[5] ) );
  NAND4_X2 U5462 ( .A1(\SB1_1_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_8/Component_Function_4/NAND4_in[1] ), .A3(n5746), .A4(
        \SB1_1_8/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_8/buf_output[4] ) );
  NAND4_X2 U5463 ( .A1(n6250), .A2(\SB1_2_0/Component_Function_5/NAND4_in[2] ), 
        .A3(\SB1_2_0/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_2_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_0/buf_output[5] ) );
  XOR2_X1 U5464 ( .A1(n5896), .A2(n5515), .Z(\MC_ARK_ARC_1_1/temp5[101] ) );
  XOR2_X1 U5465 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[71] ), .A2(\RI5[1][47] ), 
        .Z(n5515) );
  NAND4_X2 U5467 ( .A1(n7101), .A2(\SB2_2_8/Component_Function_2/NAND4_in[0] ), 
        .A3(n4651), .A4(n4028), .ZN(\SB2_2_8/buf_output[2] ) );
  XOR2_X1 U5471 ( .A1(\RI5[0][50] ), .A2(\RI5[0][188] ), .Z(n816) );
  XOR2_X1 U5474 ( .A1(\RI5[0][53] ), .A2(\RI5[0][17] ), .Z(
        \MC_ARK_ARC_1_0/temp3[143] ) );
  NAND3_X2 U5478 ( .A1(\SB1_2_10/i0[6] ), .A2(\SB1_2_10/i0[10] ), .A3(
        \SB1_2_10/i0_0 ), .ZN(\SB1_2_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U5479 ( .A1(\SB1_0_28/i0[10] ), .A2(\SB1_0_28/i1[9] ), .A3(
        \SB1_0_28/i1_7 ), .ZN(n2540) );
  XOR2_X1 U5480 ( .A1(\MC_ARK_ARC_1_1/temp6[65] ), .A2(
        \MC_ARK_ARC_1_1/temp5[65] ), .Z(\MC_ARK_ARC_1_1/buf_output[65] ) );
  XOR2_X1 U5485 ( .A1(n2891), .A2(n6623), .Z(\MC_ARK_ARC_1_1/buf_output[112] )
         );
  XOR2_X1 U5488 ( .A1(\SB2_3_11/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[99] ), .Z(n5748) );
  XOR2_X1 U5493 ( .A1(\MC_ARK_ARC_1_0/temp6[37] ), .A2(
        \MC_ARK_ARC_1_0/temp5[37] ), .Z(\MC_ARK_ARC_1_0/buf_output[37] ) );
  XOR2_X1 U5494 ( .A1(\RI5[0][165] ), .A2(\SB2_0_12/buf_output[3] ), .Z(n4893)
         );
  NAND3_X2 U5497 ( .A1(\SB2_0_6/i0_4 ), .A2(\SB2_0_6/i0_0 ), .A3(
        \SB2_0_6/i0_3 ), .ZN(\SB2_0_6/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U5499 ( .A1(n2600), .A2(\SB2_0_16/Component_Function_4/NAND4_in[3] ), .A3(\SB2_0_16/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_0_16/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB2_0_16/buf_output[4] ) );
  NAND3_X2 U5501 ( .A1(\SB1_0_26/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_26/Component_Function_5/NAND4_in[2] ), .A3(n5516), .ZN(
        \RI3[0][35] ) );
  AOI22_X2 U5509 ( .A1(\SB1_0_26/i0_0 ), .A2(\SB1_0_26/i3[0] ), .B1(
        \SB1_0_26/i0_4 ), .B2(n5517), .ZN(n5516) );
  AND2_X1 U5510 ( .A1(n226), .A2(n263), .Z(n5517) );
  XOR2_X1 U5518 ( .A1(\MC_ARK_ARC_1_1/temp2[68] ), .A2(n5518), .Z(
        \MC_ARK_ARC_1_1/temp5[68] ) );
  XOR2_X1 U5519 ( .A1(\RI5[1][68] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .Z(n5518) );
  XOR2_X1 U5520 ( .A1(\MC_ARK_ARC_1_4/temp2[130] ), .A2(n5520), .Z(n6397) );
  XOR2_X1 U5523 ( .A1(\RI5[4][130] ), .A2(\RI5[4][124] ), .Z(n5520) );
  NAND4_X2 U5524 ( .A1(\SB1_2_20/Component_Function_3/NAND4_in[1] ), .A2(n3626), .A3(\SB1_2_20/Component_Function_3/NAND4_in[0] ), .A4(n5521), .ZN(
        \SB1_2_20/buf_output[3] ) );
  NAND3_X2 U5525 ( .A1(\SB1_2_20/i0[10] ), .A2(\SB1_2_20/i1[9] ), .A3(
        \SB1_2_20/i1_7 ), .ZN(n5521) );
  XOR2_X1 U5526 ( .A1(n5523), .A2(n5522), .Z(\MC_ARK_ARC_1_1/buf_output[141] )
         );
  XOR2_X1 U5528 ( .A1(n1126), .A2(\MC_ARK_ARC_1_1/temp4[141] ), .Z(n5522) );
  XOR2_X1 U5530 ( .A1(\MC_ARK_ARC_1_1/temp2[141] ), .A2(
        \MC_ARK_ARC_1_1/temp3[141] ), .Z(n5523) );
  NAND4_X2 U5532 ( .A1(\SB2_2_24/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_2_24/Component_Function_3/NAND4_in[3] ), .A3(n5525), .A4(n5524), 
        .ZN(\SB2_2_24/buf_output[3] ) );
  NAND3_X2 U5533 ( .A1(\SB2_2_24/i0[10] ), .A2(\SB2_2_24/i1[9] ), .A3(
        \SB2_2_24/i1_7 ), .ZN(n5524) );
  NAND3_X2 U5535 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i1[9] ), .A3(
        \SB2_2_24/i0[6] ), .ZN(n5525) );
  XOR2_X1 U5536 ( .A1(\MC_ARK_ARC_1_2/temp5[3] ), .A2(
        \MC_ARK_ARC_1_2/temp6[3] ), .Z(\MC_ARK_ARC_1_2/buf_output[3] ) );
  XOR2_X1 U5537 ( .A1(\MC_ARK_ARC_1_2/temp2[3] ), .A2(n6887), .Z(
        \MC_ARK_ARC_1_2/temp5[3] ) );
  NAND3_X2 U5538 ( .A1(\SB2_0_26/i0_0 ), .A2(\SB2_0_26/i1_5 ), .A3(
        \SB2_0_26/i0_4 ), .ZN(\SB2_0_26/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 U5540 ( .I(\SB2_3_25/buf_output[5] ), .Z(\RI5[3][41] ) );
  NAND3_X2 U5555 ( .A1(n6432), .A2(\SB2_1_16/i0_4 ), .A3(\SB2_1_16/i1_5 ), 
        .ZN(\SB2_1_16/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U5556 ( .A1(\SB1_2_3/Component_Function_5/NAND4_in[2] ), .A2(n2595), 
        .A3(\SB1_2_3/Component_Function_5/NAND4_in[0] ), .A4(n5394), .ZN(
        \SB1_2_3/buf_output[5] ) );
  XOR2_X1 U5557 ( .A1(n5526), .A2(n7392), .Z(\MC_ARK_ARC_1_4/buf_output[74] )
         );
  XOR2_X1 U5558 ( .A1(n7314), .A2(n7315), .Z(n5526) );
  XOR2_X1 U5559 ( .A1(\RI5[0][148] ), .A2(\RI5[0][142] ), .Z(
        \MC_ARK_ARC_1_0/temp1[148] ) );
  INV_X2 U5560 ( .I(\SB1_3_28/buf_output[2] ), .ZN(\SB2_3_25/i1[9] ) );
  NAND4_X2 U5561 ( .A1(n4977), .A2(\SB1_3_28/Component_Function_2/NAND4_in[2] ), .A3(n2675), .A4(\SB1_3_28/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_3_28/buf_output[2] ) );
  XOR2_X1 U5562 ( .A1(n5527), .A2(\MC_ARK_ARC_1_3/temp3[36] ), .Z(n4659) );
  XOR2_X1 U5564 ( .A1(\RI5[3][30] ), .A2(\RI5[3][36] ), .Z(n5527) );
  NAND4_X2 U5565 ( .A1(\SB2_1_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_5/Component_Function_2/NAND4_in[3] ), .A3(n4441), .A4(n5528), 
        .ZN(\SB2_1_5/buf_output[2] ) );
  NAND3_X1 U5567 ( .A1(\SB2_1_5/i0[10] ), .A2(\SB2_1_5/i0[6] ), .A3(
        \SB1_1_5/buf_output[5] ), .ZN(n5528) );
  NAND3_X1 U5568 ( .A1(\SB2_0_3/i0_0 ), .A2(\SB2_0_3/i3[0] ), .A3(
        \SB2_0_3/i1_7 ), .ZN(\SB2_0_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U5570 ( .A1(\SB1_1_19/i0_0 ), .A2(\SB1_1_19/i0_4 ), .A3(
        \SB1_1_19/i1_5 ), .ZN(\SB1_1_19/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U5573 ( .A1(\MC_ARK_ARC_1_1/temp5[64] ), .A2(n5529), .Z(
        \MC_ARK_ARC_1_1/buf_output[64] ) );
  XOR2_X1 U5574 ( .A1(\MC_ARK_ARC_1_1/temp4[64] ), .A2(
        \MC_ARK_ARC_1_1/temp3[64] ), .Z(n5529) );
  NAND3_X2 U5578 ( .A1(\SB2_4_11/i0_0 ), .A2(\SB2_4_11/i0_3 ), .A3(
        \SB2_4_11/i0_4 ), .ZN(n7114) );
  INV_X2 U5579 ( .I(\MC_ARK_ARC_1_3/buf_output[26] ), .ZN(n5530) );
  NAND4_X2 U5580 ( .A1(n5258), .A2(n2977), .A3(
        \SB4_0/Component_Function_3/NAND4_in[3] ), .A4(n6065), .ZN(n5534) );
  NAND3_X2 U5582 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i0[9] ), .A3(
        \SB2_3_24/i0[8] ), .ZN(\SB2_3_24/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U5583 ( .A1(\SB1_4_27/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_4_27/Component_Function_5/NAND4_in[1] ), .A3(n4587), .A4(
        \SB1_4_27/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_4_27/buf_output[5] ) );
  NAND4_X2 U5586 ( .A1(\SB1_1_8/Component_Function_5/NAND4_in[1] ), .A2(n4588), 
        .A3(\SB1_1_8/Component_Function_5/NAND4_in[0] ), .A4(n5177), .ZN(
        \SB1_1_8/buf_output[5] ) );
  XOR2_X1 U5589 ( .A1(\MC_ARK_ARC_1_3/temp1[119] ), .A2(n5531), .Z(n1947) );
  XOR2_X1 U5595 ( .A1(\RI5[3][65] ), .A2(\RI5[3][89] ), .Z(n5531) );
  NAND3_X1 U5596 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i0[8] ), .A3(
        \SB1_0_20/i0[9] ), .ZN(\SB1_0_20/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U5597 ( .A1(\MC_ARK_ARC_1_3/temp6[31] ), .A2(n5532), .Z(
        \MC_ARK_ARC_1_3/buf_output[31] ) );
  XOR2_X1 U5602 ( .A1(n5668), .A2(\MC_ARK_ARC_1_3/temp1[31] ), .Z(n5532) );
  NAND3_X2 U5603 ( .A1(\SB2_4_26/i0_3 ), .A2(\SB2_4_26/i0[9] ), .A3(
        \SB2_4_26/i0[8] ), .ZN(n6102) );
  XOR2_X1 U5604 ( .A1(n5533), .A2(n135), .Z(Ciphertext[91]) );
  NAND4_X2 U5606 ( .A1(\SB4_16/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_16/Component_Function_1/NAND4_in[1] ), .A3(n6045), .A4(
        \SB4_16/Component_Function_1/NAND4_in[0] ), .ZN(n5533) );
  XOR2_X1 U5610 ( .A1(n5534), .A2(n151), .Z(Ciphertext[189]) );
  XOR2_X1 U5611 ( .A1(n5828), .A2(n5535), .Z(n7350) );
  XOR2_X1 U5613 ( .A1(\RI5[4][179] ), .A2(\RI5[4][59] ), .Z(n5535) );
  INV_X1 U5615 ( .I(\SB3_2/buf_output[3] ), .ZN(\SB4_0/i0[8] ) );
  NAND4_X2 U5617 ( .A1(\SB2_4_11/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_11/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_4_11/Component_Function_0/NAND4_in[0] ), .A4(n5536), .ZN(
        \SB2_4_11/buf_output[0] ) );
  NAND3_X1 U5619 ( .A1(\SB2_4_11/i0_3 ), .A2(\SB2_4_11/i0_0 ), .A3(
        \SB2_4_11/i0[7] ), .ZN(n5536) );
  XOR2_X1 U5620 ( .A1(n5537), .A2(n46), .Z(Ciphertext[174]) );
  NAND4_X2 U5623 ( .A1(\SB4_2/Component_Function_0/NAND4_in[3] ), .A2(n5250), 
        .A3(\SB4_2/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_2/Component_Function_0/NAND4_in[0] ), .ZN(n5537) );
  XOR2_X1 U5625 ( .A1(\MC_ARK_ARC_1_4/temp5[114] ), .A2(n5538), .Z(
        \MC_ARK_ARC_1_4/buf_output[114] ) );
  XOR2_X1 U5627 ( .A1(\MC_ARK_ARC_1_4/temp4[114] ), .A2(
        \MC_ARK_ARC_1_4/temp3[114] ), .Z(n5538) );
  NAND3_X2 U5629 ( .A1(\RI3[0][82] ), .A2(\SB2_0_18/i0[8] ), .A3(
        \SB2_0_18/i1_7 ), .ZN(n7316) );
  XOR2_X1 U5631 ( .A1(\SB2_3_29/buf_output[3] ), .A2(\RI5[3][93] ), .Z(n7043)
         );
  INV_X2 U5633 ( .I(\RI3[0][3] ), .ZN(\SB2_0_31/i0[8] ) );
  NAND4_X2 U5637 ( .A1(\SB1_0_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_1/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_1/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_0_1/Component_Function_3/NAND4_in[1] ), .ZN(\RI3[0][3] ) );
  NAND4_X2 U5639 ( .A1(n6729), .A2(n5210), .A3(
        \SB2_1_6/Component_Function_3/NAND4_in[0] ), .A4(
        \SB2_1_6/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_1_6/buf_output[3] ) );
  NAND3_X1 U5640 ( .A1(\SB4_23/i0[6] ), .A2(\SB4_23/i0[9] ), .A3(\SB4_23/i1_5 ), .ZN(\SB4_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U5645 ( .A1(\SB3_31/i0[9] ), .A2(\SB3_31/i0[8] ), .A3(\SB3_31/i0_3 ), .ZN(\SB3_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U5646 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i0_3 ), .A3(\SB4_12/i0[7] ), 
        .ZN(\SB4_12/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U5651 ( .A1(n7552), .A2(\MC_ARK_ARC_1_0/temp2[47] ), .Z(n1569) );
  NAND3_X2 U5652 ( .A1(\SB1_1_8/i0_3 ), .A2(\SB1_1_8/i0[6] ), .A3(
        \SB1_1_8/i1[9] ), .ZN(\SB1_1_8/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U5654 ( .A1(n5539), .A2(\MC_ARK_ARC_1_3/temp4[95] ), .Z(n2845) );
  XOR2_X1 U5656 ( .A1(\RI5[3][95] ), .A2(\RI5[3][89] ), .Z(n5539) );
  NAND3_X2 U5659 ( .A1(\SB2_4_26/i0_3 ), .A2(\SB2_4_26/i1[9] ), .A3(
        \SB2_4_26/i0_4 ), .ZN(n1744) );
  BUF_X4 U5660 ( .I(\MC_ARK_ARC_1_4/buf_output[101] ), .Z(\SB3_15/i0_3 ) );
  BUF_X4 U5662 ( .I(\SB2_1_21/buf_output[3] ), .Z(\RI5[1][75] ) );
  NAND4_X2 U5664 ( .A1(n1403), .A2(\SB4_27/Component_Function_2/NAND4_in[0] ), 
        .A3(n4486), .A4(n5540), .ZN(n5657) );
  NAND3_X1 U5670 ( .A1(\SB4_27/i0_4 ), .A2(\SB4_27/i0_0 ), .A3(\SB4_27/i1_5 ), 
        .ZN(n5540) );
  XOR2_X1 U5671 ( .A1(n861), .A2(\MC_ARK_ARC_1_0/temp6[143] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[143] ) );
  NAND3_X1 U5677 ( .A1(\SB3_24/i0[9] ), .A2(\SB3_24/i0_4 ), .A3(
        \MC_ARK_ARC_1_4/buf_output[43] ), .ZN(
        \SB3_24/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 U5678 ( .I(\SB2_4_4/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[167] ) );
  XOR2_X1 U5679 ( .A1(n5880), .A2(n7468), .Z(n6317) );
  XOR2_X1 U5680 ( .A1(\MC_ARK_ARC_1_4/temp6[28] ), .A2(
        \MC_ARK_ARC_1_4/temp5[28] ), .Z(\MC_ARK_ARC_1_4/buf_output[28] ) );
  XOR2_X1 U5683 ( .A1(\MC_ARK_ARC_1_3/temp5[153] ), .A2(
        \MC_ARK_ARC_1_3/temp6[153] ), .Z(n3968) );
  XOR2_X1 U5685 ( .A1(n4274), .A2(\MC_ARK_ARC_1_3/temp4[153] ), .Z(
        \MC_ARK_ARC_1_3/temp6[153] ) );
  NAND3_X2 U5686 ( .A1(\SB2_1_21/i0[10] ), .A2(\SB2_1_21/i1_7 ), .A3(
        \SB2_1_21/i1[9] ), .ZN(\SB2_1_21/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U5687 ( .A1(n5542), .A2(n5541), .Z(n1720) );
  XOR2_X1 U5688 ( .A1(\RI5[4][95] ), .A2(\RI5[4][89] ), .Z(n5541) );
  NAND4_X2 U5690 ( .A1(n7189), .A2(\SB4_24/Component_Function_3/NAND4_in[1] ), 
        .A3(\SB4_24/Component_Function_3/NAND4_in[3] ), .A4(n6108), .ZN(n5701)
         );
  INV_X2 U5691 ( .I(\SB1_4_20/buf_output[2] ), .ZN(\SB2_4_17/i1[9] ) );
  NAND4_X2 U5692 ( .A1(\SB1_4_20/Component_Function_2/NAND4_in[2] ), .A2(n6485), .A3(n7119), .A4(n2034), .ZN(\SB1_4_20/buf_output[2] ) );
  XOR2_X1 U5693 ( .A1(\RI5[4][40] ), .A2(\RI5[4][46] ), .Z(
        \MC_ARK_ARC_1_4/temp1[46] ) );
  NAND3_X2 U5694 ( .A1(\SB1_0_1/i0[6] ), .A2(\SB1_0_1/i1_5 ), .A3(
        \SB1_0_1/i0[9] ), .ZN(\SB1_0_1/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U5695 ( .A1(\MC_ARK_ARC_1_1/temp2[165] ), .A2(n3319), .Z(n4044) );
  NAND4_X2 U5700 ( .A1(n2199), .A2(\SB1_4_26/Component_Function_5/NAND4_in[2] ), .A3(\SB1_4_26/Component_Function_5/NAND4_in[0] ), .A4(n5543), .ZN(
        \SB1_4_26/buf_output[5] ) );
  NAND3_X2 U5701 ( .A1(\SB1_4_26/i0[10] ), .A2(\SB1_4_26/i0[6] ), .A3(
        \SB1_4_26/i0_0 ), .ZN(n5543) );
  XOR2_X1 U5703 ( .A1(\MC_ARK_ARC_1_4/temp2[94] ), .A2(
        \MC_ARK_ARC_1_4/temp1[94] ), .Z(\MC_ARK_ARC_1_4/temp5[94] ) );
  NAND3_X1 U5704 ( .A1(\SB4_30/i0_4 ), .A2(\SB4_30/i0_3 ), .A3(n5427), .ZN(
        n5546) );
  NAND4_X2 U5705 ( .A1(\SB3_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_1/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_1/Component_Function_2/NAND4_in[1] ), .A4(n4293), .ZN(
        \SB4_30/i0_0 ) );
  NAND4_X2 U5708 ( .A1(n1537), .A2(\SB1_3_15/Component_Function_5/NAND4_in[2] ), .A3(n3637), .A4(\SB1_3_15/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_15/buf_output[5] ) );
  XOR2_X1 U5710 ( .A1(n5544), .A2(n72), .Z(Ciphertext[177]) );
  NAND4_X2 U5714 ( .A1(n7514), .A2(\SB4_2/Component_Function_3/NAND4_in[3] ), 
        .A3(n4222), .A4(\SB4_2/Component_Function_3/NAND4_in[2] ), .ZN(n5544)
         );
  NAND4_X2 U5719 ( .A1(n2454), .A2(n4819), .A3(
        \SB1_2_24/Component_Function_5/NAND4_in[0] ), .A4(n5545), .ZN(
        \SB1_2_24/buf_output[5] ) );
  NAND3_X2 U5721 ( .A1(\SB1_2_24/i0[6] ), .A2(\SB1_2_24/i0[10] ), .A3(
        \SB1_2_24/i0_0 ), .ZN(n5545) );
  NAND3_X2 U5722 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0[6] ), .A3(
        \SB2_3_15/i1[9] ), .ZN(\SB2_3_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U5725 ( .A1(\SB1_0_1/i0[6] ), .A2(\SB1_0_1/i0[8] ), .A3(
        \SB1_0_1/i0[7] ), .ZN(\SB1_0_1/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U5726 ( .A1(\SB4_12/Component_Function_5/NAND4_in[2] ), .A2(n7442), 
        .A3(\SB4_12/Component_Function_5/NAND4_in[3] ), .A4(n5547), .ZN(n6190)
         );
  XOR2_X1 U5727 ( .A1(\RI5[3][92] ), .A2(\RI5[3][98] ), .Z(
        \MC_ARK_ARC_1_3/temp1[98] ) );
  XOR2_X1 U5728 ( .A1(\MC_ARK_ARC_1_3/temp6[188] ), .A2(
        \MC_ARK_ARC_1_3/temp5[188] ), .Z(\MC_ARK_ARC_1_3/buf_output[188] ) );
  XOR2_X1 U5729 ( .A1(n4304), .A2(\MC_ARK_ARC_1_3/temp4[188] ), .Z(
        \MC_ARK_ARC_1_3/temp6[188] ) );
  XOR2_X1 U5734 ( .A1(n5548), .A2(n17), .Z(Ciphertext[123]) );
  NAND4_X2 U5736 ( .A1(\SB4_11/Component_Function_3/NAND4_in[1] ), .A2(n1790), 
        .A3(n6546), .A4(n5729), .ZN(n5548) );
  XOR2_X1 U5737 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), .A2(\RI5[3][85] ), 
        .Z(n2128) );
  AND3_X1 U5738 ( .A1(\MC_ARK_ARC_1_4/buf_output[67] ), .A2(
        \MC_ARK_ARC_1_4/buf_output[66] ), .A3(\MC_ARK_ARC_1_4/buf_output[70] ), 
        .Z(n5670) );
  NAND3_X2 U5739 ( .A1(n5669), .A2(n4913), .A3(
        \SB3_20/Component_Function_5/NAND4_in[1] ), .ZN(\SB3_20/buf_output[5] ) );
  NAND4_X2 U5740 ( .A1(n2516), .A2(\SB1_3_15/Component_Function_3/NAND4_in[2] ), .A3(\SB1_3_15/Component_Function_3/NAND4_in[1] ), .A4(n5549), .ZN(
        \SB1_3_15/buf_output[3] ) );
  NAND3_X2 U5744 ( .A1(\SB1_2_21/i0[9] ), .A2(\SB1_2_21/i0[8] ), .A3(
        \SB1_2_21/i0_3 ), .ZN(n6338) );
  NAND3_X2 U5748 ( .A1(\SB1_4_2/i0_0 ), .A2(\SB1_4_2/i0[10] ), .A3(
        \SB1_4_2/i0[6] ), .ZN(n5550) );
  NAND4_X2 U5749 ( .A1(n4466), .A2(\SB1_2_9/Component_Function_5/NAND4_in[2] ), 
        .A3(n5837), .A4(n5551), .ZN(\SB1_2_9/buf_output[5] ) );
  NAND3_X2 U5751 ( .A1(\SB2_0_13/i0_3 ), .A2(\RI3[0][112] ), .A3(
        \SB2_0_13/i0_0 ), .ZN(n5552) );
  NAND3_X2 U5752 ( .A1(\SB2_2_26/i0_0 ), .A2(\SB2_2_26/i0[6] ), .A3(
        \SB2_2_26/i0[10] ), .ZN(n5553) );
  XOR2_X1 U5755 ( .A1(\MC_ARK_ARC_1_2/temp2[119] ), .A2(n5555), .Z(n5759) );
  XOR2_X1 U5760 ( .A1(\RI5[2][119] ), .A2(\RI5[2][113] ), .Z(n5555) );
  NAND4_X2 U5761 ( .A1(\SB2_4_14/Component_Function_2/NAND4_in[0] ), .A2(n6654), .A3(\SB2_4_14/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_4_14/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_4_14/buf_output[2] ) );
  XOR2_X1 U5764 ( .A1(n1608), .A2(n5556), .Z(n2197) );
  XOR2_X1 U5768 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[164] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[158] ), .Z(n5556) );
  NAND4_X2 U5769 ( .A1(n2045), .A2(\SB1_3_18/Component_Function_5/NAND4_in[0] ), .A3(\SB1_3_18/Component_Function_5/NAND4_in[1] ), .A4(n5557), .ZN(
        \SB1_3_18/buf_output[5] ) );
  NAND3_X2 U5770 ( .A1(\SB1_3_18/i0_3 ), .A2(\SB1_3_18/i1[9] ), .A3(
        \SB1_3_18/i0_4 ), .ZN(n5557) );
  XOR2_X1 U5775 ( .A1(n1480), .A2(n4979), .Z(\MC_ARK_ARC_1_3/buf_output[117] )
         );
  XOR2_X1 U5776 ( .A1(n727), .A2(\MC_ARK_ARC_1_3/temp4[117] ), .Z(n1480) );
  NAND3_X2 U5780 ( .A1(\SB2_2_9/i0[10] ), .A2(\SB2_2_9/i0_3 ), .A3(
        \SB2_2_9/i0[6] ), .ZN(n6032) );
  NAND4_X2 U5782 ( .A1(\SB2_2_10/Component_Function_5/NAND4_in[2] ), .A2(n4245), .A3(\SB2_2_10/Component_Function_5/NAND4_in[1] ), .A4(n5558), .ZN(
        \SB2_2_10/buf_output[5] ) );
  NAND3_X2 U5784 ( .A1(\SB2_2_10/i0[6] ), .A2(\SB2_2_10/i0_4 ), .A3(
        \SB2_2_10/i0[9] ), .ZN(n5558) );
  XOR2_X1 U5787 ( .A1(n5559), .A2(n12), .Z(Ciphertext[4]) );
  NAND4_X2 U5790 ( .A1(\SB4_31/Component_Function_4/NAND4_in[3] ), .A2(n2233), 
        .A3(n5634), .A4(n3732), .ZN(n5559) );
  NAND4_X2 U5791 ( .A1(n5189), .A2(\SB1_2_11/Component_Function_3/NAND4_in[1] ), .A3(n6298), .A4(\SB1_2_11/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB1_2_11/buf_output[3] ) );
  NAND4_X2 U5798 ( .A1(n6821), .A2(\SB1_4_11/Component_Function_5/NAND4_in[1] ), .A3(n5068), .A4(\SB1_4_11/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_4_11/buf_output[5] ) );
  NAND4_X2 U5800 ( .A1(n6944), .A2(n1551), .A3(n932), .A4(
        \SB2_1_10/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_10/buf_output[3] ) );
  NAND3_X2 U5801 ( .A1(\SB1_0_13/i0_3 ), .A2(n5428), .A3(\SB1_0_13/i1_7 ), 
        .ZN(\SB1_0_13/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U5802 ( .A1(n5560), .A2(n6725), .Z(n5625) );
  XOR2_X1 U5803 ( .A1(\RI5[3][57] ), .A2(\RI5[3][63] ), .Z(n5560) );
  XOR2_X1 U5806 ( .A1(\MC_ARK_ARC_1_1/temp6[35] ), .A2(n5561), .Z(
        \MC_ARK_ARC_1_1/buf_output[35] ) );
  XOR2_X1 U5808 ( .A1(n6151), .A2(n6436), .Z(n5561) );
  XOR2_X1 U5810 ( .A1(\RI5[0][138] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[36] ) );
  XOR2_X1 U5812 ( .A1(n6969), .A2(n5562), .Z(n3886) );
  XOR2_X1 U5814 ( .A1(\RI5[1][51] ), .A2(\RI5[1][159] ), .Z(n5562) );
  NAND4_X2 U5815 ( .A1(\SB2_2_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_14/Component_Function_2/NAND4_in[1] ), .A3(n5151), .A4(n5563), 
        .ZN(\SB2_2_14/buf_output[2] ) );
  NAND3_X2 U5817 ( .A1(\SB2_2_14/i0[10] ), .A2(\SB2_2_14/i1[9] ), .A3(
        \SB2_2_14/i1_5 ), .ZN(n5563) );
  XOR2_X1 U5818 ( .A1(\MC_ARK_ARC_1_0/temp2[117] ), .A2(n5564), .Z(n2509) );
  XOR2_X1 U5819 ( .A1(\RI5[0][117] ), .A2(\RI5[0][111] ), .Z(n5564) );
  NAND3_X2 U5822 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i0_4 ), .A3(
        \SB2_3_1/i1[9] ), .ZN(n1623) );
  XOR2_X1 U5836 ( .A1(n5565), .A2(n106), .Z(Ciphertext[46]) );
  NAND4_X2 U5837 ( .A1(\SB4_24/Component_Function_4/NAND4_in[0] ), .A2(n5026), 
        .A3(n997), .A4(n2744), .ZN(n5565) );
  XOR2_X1 U5838 ( .A1(n5567), .A2(n5566), .Z(n6938) );
  XOR2_X1 U5842 ( .A1(\MC_ARK_ARC_1_1/temp1[54] ), .A2(
        \MC_ARK_ARC_1_1/temp4[54] ), .Z(n5566) );
  XOR2_X1 U5843 ( .A1(\MC_ARK_ARC_1_1/temp2[54] ), .A2(
        \MC_ARK_ARC_1_1/temp3[54] ), .Z(n5567) );
  XOR2_X1 U5844 ( .A1(\MC_ARK_ARC_1_3/temp5[122] ), .A2(n5568), .Z(
        \MC_ARK_ARC_1_3/buf_output[122] ) );
  XOR2_X1 U5847 ( .A1(\MC_ARK_ARC_1_3/temp3[122] ), .A2(
        \MC_ARK_ARC_1_3/temp4[122] ), .Z(n5568) );
  INV_X2 U5853 ( .I(\SB1_3_27/buf_output[2] ), .ZN(\SB2_3_24/i1[9] ) );
  NAND4_X2 U5854 ( .A1(\SB1_3_27/Component_Function_2/NAND4_in[1] ), .A2(n4615), .A3(\SB1_3_27/Component_Function_2/NAND4_in[0] ), .A4(n3580), .ZN(
        \SB1_3_27/buf_output[2] ) );
  INV_X2 U5856 ( .I(\SB1_3_19/buf_output[2] ), .ZN(\SB2_3_16/i1[9] ) );
  NAND4_X2 U5857 ( .A1(\SB1_3_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_2/NAND4_in[3] ), .A3(n5106), .A4(n4911), 
        .ZN(\SB1_3_19/buf_output[2] ) );
  XOR2_X1 U5860 ( .A1(n5569), .A2(n177), .Z(Ciphertext[116]) );
  NAND4_X2 U5864 ( .A1(\SB4_12/Component_Function_2/NAND4_in[0] ), .A2(n2749), 
        .A3(\SB4_12/Component_Function_2/NAND4_in[2] ), .A4(n4051), .ZN(n5569)
         );
  NAND3_X2 U5865 ( .A1(\SB3_12/i0[10] ), .A2(\SB3_12/i0[6] ), .A3(
        \SB3_12/i0_0 ), .ZN(\SB3_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U5868 ( .A1(\SB2_4_8/i0_3 ), .A2(\SB2_4_8/i0_0 ), .A3(n3183), .ZN(
        n5576) );
  NAND4_X2 U5869 ( .A1(\SB2_0_7/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_7/Component_Function_2/NAND4_in[2] ), .A3(n3460), .A4(n5570), 
        .ZN(\SB2_0_7/buf_output[2] ) );
  NAND3_X2 U5870 ( .A1(\SB2_0_7/i0[10] ), .A2(\SB2_0_7/i1_5 ), .A3(
        \SB2_0_7/i1[9] ), .ZN(n5570) );
  NAND3_X2 U5872 ( .A1(n6746), .A2(\SB2_3_13/i1_5 ), .A3(\SB2_3_13/i0_0 ), 
        .ZN(n6070) );
  NAND4_X2 U5874 ( .A1(\SB2_4_9/Component_Function_2/NAND4_in[2] ), .A2(n1799), 
        .A3(n4635), .A4(n5571), .ZN(\SB2_4_9/buf_output[2] ) );
  NAND3_X1 U5875 ( .A1(\SB2_4_9/i0[10] ), .A2(\SB2_4_9/i1_5 ), .A3(
        \SB2_4_9/i1[9] ), .ZN(n5571) );
  XOR2_X1 U5879 ( .A1(n5572), .A2(n67), .Z(Ciphertext[120]) );
  NAND4_X2 U5881 ( .A1(\SB4_11/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_11/Component_Function_0/NAND4_in[2] ), .A3(n1911), .A4(
        \SB4_11/Component_Function_0/NAND4_in[0] ), .ZN(n5572) );
  INV_X1 U5882 ( .I(\SB3_1/buf_output[3] ), .ZN(\SB4_31/i0[8] ) );
  NAND4_X2 U5884 ( .A1(\SB3_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_1/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_1/Component_Function_3/NAND4_in[2] ), .A4(n2062), .ZN(
        \SB3_1/buf_output[3] ) );
  INV_X2 U5886 ( .I(\SB1_2_1/buf_output[2] ), .ZN(\SB2_2_30/i1[9] ) );
  NAND4_X2 U5887 ( .A1(\SB1_2_1/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_1/Component_Function_2/NAND4_in[1] ), .A3(n6052), .A4(n6860), 
        .ZN(\SB1_2_1/buf_output[2] ) );
  INV_X2 U5889 ( .I(\SB1_3_27/buf_output[3] ), .ZN(\SB2_3_25/i0[8] ) );
  NAND4_X2 U5890 ( .A1(\SB1_3_27/Component_Function_3/NAND4_in[0] ), .A2(n3887), .A3(n2763), .A4(n5886), .ZN(\SB1_3_27/buf_output[3] ) );
  XOR2_X1 U5891 ( .A1(\MC_ARK_ARC_1_2/temp2[58] ), .A2(n5573), .Z(
        \MC_ARK_ARC_1_2/temp5[58] ) );
  XOR2_X1 U5893 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[52] ), .A2(\RI5[2][58] ), 
        .Z(n5573) );
  XOR2_X1 U5897 ( .A1(n6826), .A2(n5574), .Z(n4608) );
  XOR2_X1 U5906 ( .A1(\RI5[0][125] ), .A2(\SB2_0_26/buf_output[5] ), .Z(n5574)
         );
  NAND4_X2 U5913 ( .A1(\SB2_4_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_4_8/Component_Function_2/NAND4_in[2] ), .A4(n5575), .ZN(
        \SB2_4_8/buf_output[2] ) );
  NAND3_X1 U5914 ( .A1(\SB2_4_8/i0_0 ), .A2(\SB2_4_8/i1_5 ), .A3(n3183), .ZN(
        n5575) );
  NAND4_X2 U5915 ( .A1(\SB2_4_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_8/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_4_8/Component_Function_3/NAND4_in[3] ), .A4(n5576), .ZN(
        \SB2_4_8/buf_output[3] ) );
  BUF_X4 U5917 ( .I(\MC_ARK_ARC_1_3/buf_output[76] ), .Z(\SB1_4_19/i0_4 ) );
  XOR2_X1 U5918 ( .A1(\RI5[3][22] ), .A2(\SB2_3_25/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/temp2[76] ) );
  XOR2_X1 U5921 ( .A1(n5577), .A2(\MC_ARK_ARC_1_1/temp2[81] ), .Z(n5579) );
  XOR2_X1 U5922 ( .A1(\SB2_1_21/buf_output[3] ), .A2(\RI5[1][81] ), .Z(n5577)
         );
  XOR2_X1 U5924 ( .A1(n5894), .A2(\MC_ARK_ARC_1_2/temp6[62] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[62] ) );
  NAND3_X1 U5928 ( .A1(\SB1_1_3/i0[6] ), .A2(\SB1_1_3/i0_3 ), .A3(
        \SB1_1_3/i1[9] ), .ZN(\SB1_1_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U5932 ( .A1(\SB1_0_24/i0[10] ), .A2(\SB1_0_24/i1[9] ), .A3(
        \SB1_0_24/i1_5 ), .ZN(n5023) );
  NAND4_X2 U5934 ( .A1(\SB1_1_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_16/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_1_16/Component_Function_2/NAND4_in[1] ), .A4(n5709), .ZN(
        \SB1_1_16/buf_output[2] ) );
  NAND4_X2 U5940 ( .A1(\SB2_3_25/Component_Function_2/NAND4_in[0] ), .A2(n7018), .A3(\SB2_3_25/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_25/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_3_25/buf_output[2] ) );
  NAND4_X2 U5945 ( .A1(n2291), .A2(\SB1_1_2/Component_Function_3/NAND4_in[1] ), 
        .A3(\SB1_1_2/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_1_2/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB1_1_2/buf_output[3] ) );
  NAND3_X2 U5947 ( .A1(\SB2_4_27/i0[6] ), .A2(\SB2_4_27/i0_4 ), .A3(
        \SB2_4_27/i0[9] ), .ZN(n5107) );
  NAND3_X2 U5948 ( .A1(\SB1_2_17/i0[10] ), .A2(\SB1_2_17/i1[9] ), .A3(
        \SB1_2_17/i1_5 ), .ZN(n6528) );
  XOR2_X1 U5951 ( .A1(\MC_ARK_ARC_1_2/temp6[61] ), .A2(
        \MC_ARK_ARC_1_2/temp5[61] ), .Z(\MC_ARK_ARC_1_2/buf_output[61] ) );
  INV_X4 U5952 ( .I(n5630), .ZN(\RI3[0][77] ) );
  NAND4_X2 U5953 ( .A1(n2431), .A2(n2180), .A3(
        \SB2_0_13/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_13/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_13/buf_output[5] ) );
  XOR2_X1 U5955 ( .A1(\MC_ARK_ARC_1_2/temp5[183] ), .A2(n1104), .Z(n6276) );
  XOR2_X1 U5958 ( .A1(n1296), .A2(\MC_ARK_ARC_1_2/temp4[183] ), .Z(n1104) );
  XOR2_X1 U5960 ( .A1(n1401), .A2(n5578), .Z(\MC_ARK_ARC_1_4/temp5[105] ) );
  XOR2_X1 U5968 ( .A1(\RI5[4][105] ), .A2(\RI5[4][99] ), .Z(n5578) );
  XOR2_X1 U5969 ( .A1(n666), .A2(n5579), .Z(\MC_ARK_ARC_1_1/buf_output[81] )
         );
  INV_X2 U5970 ( .I(\SB1_1_28/buf_output[3] ), .ZN(\SB2_1_26/i0[8] ) );
  NAND4_X2 U5979 ( .A1(\SB1_1_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_28/Component_Function_3/NAND4_in[1] ), .A3(n1717), .A4(n6437), 
        .ZN(\SB1_1_28/buf_output[3] ) );
  NAND3_X1 U5981 ( .A1(\SB3_27/i0_4 ), .A2(\SB3_27/i1_5 ), .A3(\SB3_27/i1[9] ), 
        .ZN(n4229) );
  XOR2_X1 U5982 ( .A1(n5581), .A2(n5580), .Z(\MC_ARK_ARC_1_3/buf_output[81] )
         );
  XOR2_X1 U5987 ( .A1(n6637), .A2(n6543), .Z(n5580) );
  XOR2_X1 U5992 ( .A1(n4248), .A2(n6544), .Z(n5581) );
  XOR2_X1 U5993 ( .A1(\MC_ARK_ARC_1_2/temp6[128] ), .A2(n5582), .Z(
        \MC_ARK_ARC_1_2/buf_output[128] ) );
  XOR2_X1 U5998 ( .A1(n6523), .A2(\MC_ARK_ARC_1_2/temp2[128] ), .Z(n5582) );
  NAND3_X1 U6001 ( .A1(\SB4_30/i0_3 ), .A2(\SB4_30/i0[7] ), .A3(n5427), .ZN(
        \SB4_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U6002 ( .A1(\SB2_4_5/i0_0 ), .A2(\SB1_4_6/buf_output[4] ), .A3(
        \SB2_4_5/i1_5 ), .ZN(\SB2_4_5/Component_Function_2/NAND4_in[3] ) );
  INV_X2 U6003 ( .I(\SB1_2_17/buf_output[2] ), .ZN(\SB2_2_14/i1[9] ) );
  NAND4_X2 U6004 ( .A1(\SB1_2_17/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_17/Component_Function_2/NAND4_in[2] ), .A3(n633), .A4(n6528), 
        .ZN(\SB1_2_17/buf_output[2] ) );
  XOR2_X1 U6005 ( .A1(n885), .A2(n5583), .Z(n5591) );
  XOR2_X1 U6006 ( .A1(\RI5[2][128] ), .A2(\RI5[2][104] ), .Z(n5583) );
  NAND4_X2 U6007 ( .A1(\SB2_1_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_2/NAND4_in[2] ), .A4(n5584), .ZN(
        \SB2_1_12/buf_output[2] ) );
  NAND3_X2 U6011 ( .A1(\SB2_1_12/i0_0 ), .A2(\SB2_1_12/i0_4 ), .A3(
        \SB2_1_12/i1_5 ), .ZN(n5584) );
  NOR2_X2 U6012 ( .A1(n7004), .A2(n5585), .ZN(n7587) );
  NAND3_X2 U6016 ( .A1(\SB2_0_13/i0_3 ), .A2(\SB2_0_13/i0[9] ), .A3(
        \SB2_0_13/i0[8] ), .ZN(\SB2_0_13/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U6019 ( .A1(n1994), .A2(n5586), .Z(n7312) );
  XOR2_X1 U6023 ( .A1(\RI5[0][128] ), .A2(\RI5[0][134] ), .Z(n5586) );
  NAND4_X2 U6024 ( .A1(\SB1_1_14/Component_Function_5/NAND4_in[2] ), .A2(n4786), .A3(\SB1_1_14/Component_Function_5/NAND4_in[0] ), .A4(n2723), .ZN(
        \SB1_1_14/buf_output[5] ) );
  NAND4_X2 U6026 ( .A1(\SB2_2_28/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_28/Component_Function_2/NAND4_in[0] ), .A3(n3075), .A4(
        \SB2_2_28/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_2_28/buf_output[2] ) );
  NAND4_X2 U6036 ( .A1(\SB2_0_16/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_16/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_16/Component_Function_3/NAND4_in[0] ), .A4(n5007), .ZN(
        \SB2_0_16/buf_output[3] ) );
  NAND4_X2 U6037 ( .A1(\SB2_3_0/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_0/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_3_0/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_3_0/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_0/buf_output[1] ) );
  NAND3_X2 U6038 ( .A1(\SB2_0_12/i0_0 ), .A2(\RI3[0][118] ), .A3(\RI3[0][119] ), .ZN(\SB2_0_12/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U6039 ( .A1(\MC_ARK_ARC_1_3/temp6[93] ), .A2(
        \MC_ARK_ARC_1_3/temp5[93] ), .Z(\MC_ARK_ARC_1_3/buf_output[93] ) );
  NAND3_X2 U6041 ( .A1(\SB1_3_0/i0[10] ), .A2(\SB1_3_0/i0_0 ), .A3(
        \SB1_3_0/i0[6] ), .ZN(\SB1_3_0/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U6042 ( .A1(n5588), .A2(n5587), .Z(n6988) );
  XOR2_X1 U6043 ( .A1(\SB2_0_11/buf_output[3] ), .A2(\RI5[0][81] ), .Z(n5587)
         );
  XOR2_X1 U6046 ( .A1(\RI5[0][129] ), .A2(\RI5[0][105] ), .Z(n5588) );
  NAND3_X2 U6051 ( .A1(\SB1_3_23/i0[10] ), .A2(\SB1_3_23/i0[6] ), .A3(
        \SB1_3_23/i0_0 ), .ZN(\SB1_3_23/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U6056 ( .A1(\SB1_0_4/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_4/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_0_4/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_4/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][0] ) );
  XOR2_X1 U6057 ( .A1(\SB2_0_0/buf_output[3] ), .A2(\RI5[0][3] ), .Z(n5637) );
  INV_X8 U6061 ( .I(\RI1[4][155] ), .ZN(\SB1_4_6/i1_5 ) );
  NAND4_X2 U6066 ( .A1(\SB2_1_26/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_26/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_26/Component_Function_5/NAND4_in[0] ), .A4(n5589), .ZN(
        \SB2_1_26/buf_output[5] ) );
  NAND3_X2 U6067 ( .A1(\SB2_1_26/i0[6] ), .A2(\SB2_1_26/i0_4 ), .A3(
        \SB2_1_26/i0[9] ), .ZN(n5589) );
  NAND4_X2 U6068 ( .A1(\SB1_0_4/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_4/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_5/NAND4_in[0] ), .A4(n5590), .ZN(
        \RI3[0][167] ) );
  NAND3_X2 U6069 ( .A1(\SB1_0_4/i0_4 ), .A2(\SB1_0_4/i0[6] ), .A3(
        \SB1_0_4/i0[9] ), .ZN(n5590) );
  INV_X2 U6070 ( .I(\SB3_9/buf_output[2] ), .ZN(\SB4_6/i1[9] ) );
  NAND4_X2 U6071 ( .A1(\SB3_9/Component_Function_2/NAND4_in[2] ), .A2(n7338), 
        .A3(n5608), .A4(n5912), .ZN(\SB3_9/buf_output[2] ) );
  NAND3_X2 U6073 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i0[8] ), .A3(
        \SB2_1_28/i1_7 ), .ZN(\SB2_1_28/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U6077 ( .A1(\SB2_0_15/Component_Function_5/NAND4_in[0] ), .A2(n7082), .A3(n7083), .A4(n5592), .ZN(\SB2_0_15/buf_output[5] ) );
  NAND3_X2 U6081 ( .A1(\SB2_0_15/i0_3 ), .A2(\RI3[0][100] ), .A3(n1508), .ZN(
        n5592) );
  XOR2_X1 U6082 ( .A1(n5594), .A2(n5593), .Z(n5004) );
  XOR2_X1 U6085 ( .A1(\RI5[0][125] ), .A2(n189), .Z(n5593) );
  XOR2_X1 U6087 ( .A1(\RI5[0][161] ), .A2(\RI5[0][95] ), .Z(n5594) );
  XOR2_X1 U6088 ( .A1(n5596), .A2(n5595), .Z(n7524) );
  XOR2_X1 U6092 ( .A1(\RI5[0][131] ), .A2(n200), .Z(n5595) );
  XOR2_X1 U6095 ( .A1(\RI5[0][101] ), .A2(\RI5[0][167] ), .Z(n5596) );
  NAND4_X2 U6100 ( .A1(\SB4_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_2/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_2/Component_Function_5/NAND4_in[0] ), .A4(n5597), .ZN(n7466) );
  NAND3_X1 U6104 ( .A1(\SB4_2/i0[10] ), .A2(\SB4_2/i0[6] ), .A3(\SB4_2/i0_0 ), 
        .ZN(n5597) );
  NAND4_X2 U6106 ( .A1(n6171), .A2(\SB4_30/Component_Function_2/NAND4_in[0] ), 
        .A3(n6233), .A4(n5598), .ZN(n5953) );
  XOR2_X1 U6107 ( .A1(n5599), .A2(n91), .Z(Ciphertext[47]) );
  NAND4_X2 U6110 ( .A1(\SB4_24/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_24/Component_Function_5/NAND4_in[2] ), .A3(n6413), .A4(
        \SB4_24/Component_Function_5/NAND4_in[0] ), .ZN(n5599) );
  NAND4_X2 U6111 ( .A1(n6011), .A2(\SB4_22/Component_Function_3/NAND4_in[3] ), 
        .A3(n7036), .A4(n5600), .ZN(n5672) );
  NAND3_X1 U6117 ( .A1(\SB4_22/i0[10] ), .A2(\SB4_22/i1_7 ), .A3(
        \SB4_22/i1[9] ), .ZN(n5600) );
  NAND4_X2 U6123 ( .A1(\SB1_3_22/Component_Function_5/NAND4_in[3] ), .A2(n7294), .A3(n895), .A4(n5601), .ZN(\SB1_3_22/buf_output[5] ) );
  NAND3_X2 U6124 ( .A1(\SB1_3_22/i0[10] ), .A2(\SB1_3_22/i0[6] ), .A3(
        \SB1_3_22/i0_0 ), .ZN(n5601) );
  XOR2_X1 U6130 ( .A1(n6319), .A2(n5602), .Z(n855) );
  XOR2_X1 U6131 ( .A1(\RI5[0][123] ), .A2(\RI5[0][69] ), .Z(n5602) );
  XOR2_X1 U6132 ( .A1(\MC_ARK_ARC_1_4/temp6[108] ), .A2(n5603), .Z(
        \MC_ARK_ARC_1_4/buf_output[108] ) );
  XOR2_X1 U6137 ( .A1(\MC_ARK_ARC_1_4/temp2[108] ), .A2(n7308), .Z(n5603) );
  NAND4_X2 U6138 ( .A1(n1518), .A2(\SB2_0_0/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_0_0/Component_Function_5/NAND4_in[0] ), .A4(n5604), .ZN(
        \SB2_0_0/buf_output[5] ) );
  NAND4_X2 U6144 ( .A1(\SB1_3_3/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_3/Component_Function_5/NAND4_in[2] ), .A3(n6709), .A4(
        \SB1_3_3/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_3/buf_output[5] ) );
  NAND4_X2 U6150 ( .A1(n6655), .A2(\SB1_4_6/Component_Function_1/NAND4_in[1] ), 
        .A3(n3153), .A4(n5605), .ZN(\SB1_4_6/buf_output[1] ) );
  NAND4_X2 U6152 ( .A1(\SB1_1_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_20/Component_Function_5/NAND4_in[2] ), .A3(n7513), .A4(
        \SB1_1_20/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_20/buf_output[5] ) );
  NAND4_X2 U6158 ( .A1(n5239), .A2(\SB2_3_11/Component_Function_3/NAND4_in[3] ), .A3(n3810), .A4(n5606), .ZN(\SB2_3_11/buf_output[3] ) );
  XOR2_X1 U6164 ( .A1(n5607), .A2(n27), .Z(Ciphertext[49]) );
  NAND4_X2 U6165 ( .A1(\SB4_23/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_23/Component_Function_1/NAND4_in[3] ), .A4(
        \SB4_23/Component_Function_1/NAND4_in[0] ), .ZN(n5607) );
  NAND4_X2 U6173 ( .A1(\SB2_4_8/Component_Function_4/NAND4_in[0] ), .A2(n2655), 
        .A3(\SB2_4_8/Component_Function_4/NAND4_in[3] ), .A4(n5609), .ZN(
        \SB2_4_8/buf_output[4] ) );
  NAND3_X1 U6174 ( .A1(\SB2_4_8/i0_0 ), .A2(\SB2_4_8/i3[0] ), .A3(
        \SB2_4_8/i1_7 ), .ZN(n5609) );
  BUF_X4 U6176 ( .I(\SB3_23/buf_output[5] ), .Z(\SB4_23/i0_3 ) );
  NAND4_X2 U6180 ( .A1(\SB1_4_13/Component_Function_5/NAND4_in[1] ), .A2(n6953), .A3(\SB1_4_13/Component_Function_5/NAND4_in[0] ), .A4(n5610), .ZN(
        \SB1_4_13/buf_output[5] ) );
  NAND3_X2 U6181 ( .A1(\SB1_4_13/i0[9] ), .A2(\SB1_4_13/i0_4 ), .A3(
        \SB1_4_13/i0[6] ), .ZN(n5610) );
  XOR2_X1 U6182 ( .A1(\RI5[2][116] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[122] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[122] ) );
  XOR2_X1 U6190 ( .A1(\RI5[4][180] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[12] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[42] ) );
  XOR2_X1 U6191 ( .A1(n5611), .A2(n48), .Z(Ciphertext[181]) );
  NAND4_X2 U6193 ( .A1(\SB4_1/Component_Function_1/NAND4_in[2] ), .A2(n4735), 
        .A3(\SB4_1/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_1/Component_Function_1/NAND4_in[0] ), .ZN(n5611) );
  XOR2_X1 U6195 ( .A1(n5613), .A2(n5612), .Z(\MC_ARK_ARC_1_0/temp6[56] ) );
  XOR2_X1 U6196 ( .A1(\RI5[0][122] ), .A2(n24), .Z(n5612) );
  XOR2_X1 U6201 ( .A1(\RI5[0][92] ), .A2(\RI5[0][158] ), .Z(n5613) );
  XOR2_X1 U6202 ( .A1(\SB2_0_10/buf_output[3] ), .A2(\RI5[0][165] ), .Z(n3648)
         );
  AND2_X1 U6211 ( .A1(n6547), .A2(n5614), .Z(n5831) );
  XOR2_X1 U6212 ( .A1(n6594), .A2(n5615), .Z(n4359) );
  XOR2_X1 U6214 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[15] ), .A2(\RI5[3][153] ), 
        .Z(n5615) );
  XOR2_X1 U6222 ( .A1(\MC_ARK_ARC_1_0/temp2[0] ), .A2(n5616), .Z(
        \MC_ARK_ARC_1_0/temp5[0] ) );
  XOR2_X1 U6224 ( .A1(\RI5[0][0] ), .A2(\RI5[0][186] ), .Z(n5616) );
  XOR2_X1 U6226 ( .A1(n5618), .A2(n5617), .Z(\MC_ARK_ARC_1_1/temp5[129] ) );
  XOR2_X1 U6227 ( .A1(\RI5[1][129] ), .A2(\RI5[1][99] ), .Z(n5617) );
  XOR2_X1 U6234 ( .A1(\RI5[1][75] ), .A2(\RI5[1][123] ), .Z(n5618) );
  NAND4_X2 U6235 ( .A1(\SB2_1_16/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_16/Component_Function_0/NAND4_in[3] ), .A3(n4647), .A4(n5619), 
        .ZN(\SB2_1_16/buf_output[0] ) );
  NAND2_X2 U6236 ( .A1(\SB2_1_16/i0[9] ), .A2(\SB2_1_16/i0[10] ), .ZN(n5619)
         );
  NAND4_X2 U6237 ( .A1(\SB1_3_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_14/Component_Function_2/NAND4_in[3] ), .A3(n5014), .A4(n5620), 
        .ZN(\SB1_3_14/buf_output[2] ) );
  NAND3_X2 U6240 ( .A1(\SB1_3_14/i0[9] ), .A2(\RI1[3][107] ), .A3(
        \SB1_3_14/i0[8] ), .ZN(n5620) );
  NAND3_X2 U6243 ( .A1(\SB2_3_11/i0[6] ), .A2(\SB2_3_11/i0[10] ), .A3(
        \SB2_3_11/i0_0 ), .ZN(n5706) );
  XOR2_X1 U6249 ( .A1(n5622), .A2(n5621), .Z(\MC_ARK_ARC_1_1/buf_output[172] )
         );
  XOR2_X1 U6250 ( .A1(\MC_ARK_ARC_1_1/temp4[172] ), .A2(n3202), .Z(n5621) );
  XOR2_X1 U6254 ( .A1(n3203), .A2(n6080), .Z(n5622) );
  XOR2_X1 U6255 ( .A1(n5624), .A2(n5623), .Z(\MC_ARK_ARC_1_0/buf_output[20] )
         );
  XOR2_X1 U6257 ( .A1(n5854), .A2(n7241), .Z(n5623) );
  XOR2_X1 U6262 ( .A1(n2601), .A2(n7242), .Z(n5624) );
  NAND3_X2 U6264 ( .A1(\SB2_0_25/i0[10] ), .A2(\SB2_0_25/i1_5 ), .A3(
        \SB2_0_25/i1[9] ), .ZN(\SB2_0_25/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U6265 ( .A1(\SB3_30/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_30/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_30/Component_Function_2/NAND4_in[0] ), .A4(
        \SB3_30/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_30/buf_output[2] ) );
  INV_X2 U6268 ( .I(\SB1_3_15/buf_output[2] ), .ZN(\SB2_3_12/i1[9] ) );
  NAND4_X2 U6273 ( .A1(\SB1_3_15/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_3_15/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_3_15/buf_output[2] ) );
  INV_X2 U6274 ( .I(\SB1_3_1/buf_output[2] ), .ZN(\SB2_3_30/i1[9] ) );
  NAND4_X2 U6275 ( .A1(n2724), .A2(n6587), .A3(
        \SB1_3_1/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_3_1/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_3_1/buf_output[2] ) );
  NAND4_X2 U6276 ( .A1(\SB1_3_1/Component_Function_5/NAND4_in[2] ), .A2(n5191), 
        .A3(n5816), .A4(\SB1_3_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_1/buf_output[5] ) );
  XOR2_X1 U6281 ( .A1(n4225), .A2(\MC_ARK_ARC_1_3/temp1[117] ), .Z(n4979) );
  BUF_X4 U6284 ( .I(\SB2_1_31/buf_output[1] ), .Z(\RI5[1][25] ) );
  XOR2_X1 U6287 ( .A1(n5625), .A2(n4686), .Z(\MC_ARK_ARC_1_3/buf_output[63] )
         );
  XOR2_X1 U6293 ( .A1(\MC_ARK_ARC_1_2/temp1[87] ), .A2(n5626), .Z(n3064) );
  XOR2_X1 U6296 ( .A1(\RI5[2][57] ), .A2(\RI5[2][33] ), .Z(n5626) );
  INV_X1 U6297 ( .I(\SB1_1_31/buf_output[5] ), .ZN(\SB2_1_31/i1_5 ) );
  NAND4_X2 U6298 ( .A1(\SB1_1_31/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_31/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_1_31/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_1_31/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_1_31/buf_output[5] ) );
  NAND3_X2 U6306 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0_0 ), .A3(
        \SB2_3_15/i0[7] ), .ZN(\SB2_3_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U6309 ( .A1(\SB3_6/i1_5 ), .A2(\SB3_6/i0_0 ), .A3(\SB3_6/i0_4 ), 
        .ZN(n7026) );
  NAND4_X2 U6318 ( .A1(\SB1_1_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_30/Component_Function_3/NAND4_in[1] ), .A3(n5132), .A4(n4231), 
        .ZN(\SB1_1_30/buf_output[3] ) );
  NAND4_X2 U6323 ( .A1(n4477), .A2(n4591), .A3(
        \SB1_3_12/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_3_12/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_12/buf_output[5] ) );
  NAND3_X2 U6324 ( .A1(\SB2_2_10/i0[10] ), .A2(\SB2_2_10/i1[9] ), .A3(
        \SB2_2_10/i1_7 ), .ZN(n821) );
  NAND4_X2 U6326 ( .A1(n2285), .A2(n3681), .A3(n5094), .A4(
        \SB2_4_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_4_18/buf_output[5] ) );
  NAND4_X2 U6331 ( .A1(n6859), .A2(\SB2_1_28/Component_Function_3/NAND4_in[0] ), .A3(n6858), .A4(\SB2_1_28/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_1_28/buf_output[3] ) );
  NAND4_X2 U6332 ( .A1(\SB2_0_28/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_28/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_0_28/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_28/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_28/buf_output[2] ) );
  XOR2_X1 U6335 ( .A1(n2073), .A2(n3597), .Z(\MC_ARK_ARC_1_0/buf_output[66] )
         );
  NAND4_X2 U6336 ( .A1(\SB1_3_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_3/NAND4_in[2] ), .A4(n5627), .ZN(
        \SB1_3_19/buf_output[3] ) );
  NAND3_X2 U6337 ( .A1(\SB1_3_19/i0[8] ), .A2(\SB1_3_19/i1_5 ), .A3(
        \SB1_3_19/i3[0] ), .ZN(n5627) );
  NOR2_X2 U6338 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  NAND2_X2 U6345 ( .A1(\SB1_0_19/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_0_19/Component_Function_5/NAND4_in[0] ), .ZN(n5628) );
  NAND2_X2 U6348 ( .A1(\SB1_0_19/Component_Function_5/NAND4_in[1] ), .A2(n3900), .ZN(n5629) );
  BUF_X4 U6350 ( .I(\SB3_12/buf_output[1] ), .Z(\SB4_8/i0[6] ) );
  XOR2_X1 U6351 ( .A1(\RI5[1][116] ), .A2(\RI5[1][140] ), .Z(n6300) );
  NAND3_X2 U6352 ( .A1(\SB1_4_25/i0[9] ), .A2(\SB1_4_25/i0[8] ), .A3(
        \RI1[4][41] ), .ZN(n5631) );
  XOR2_X1 U6358 ( .A1(n3087), .A2(\MC_ARK_ARC_1_1/temp5[170] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[170] ) );
  XOR2_X1 U6360 ( .A1(n7394), .A2(\MC_ARK_ARC_1_2/temp2[138] ), .Z(
        \MC_ARK_ARC_1_2/temp5[138] ) );
  NAND3_X1 U6361 ( .A1(\SB1_0_15/i0_0 ), .A2(\SB1_0_15/i0_3 ), .A3(n350), .ZN(
        \SB1_0_15/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U6365 ( .A1(\SB2_0_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_25/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_25/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_0_25/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_25/buf_output[3] ) );
  BUF_X4 U6368 ( .I(\SB1_4_25/buf_output[2] ), .Z(\SB2_4_22/i0_0 ) );
  XOR2_X1 U6369 ( .A1(n6303), .A2(\MC_ARK_ARC_1_0/temp6[56] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[56] ) );
  NAND3_X2 U6372 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0_0 ), .A3(
        \SB2_2_22/i0[7] ), .ZN(n6905) );
  NAND4_X2 U6377 ( .A1(\SB1_4_25/Component_Function_2/NAND4_in[1] ), .A2(n890), 
        .A3(n6525), .A4(n5631), .ZN(\SB1_4_25/buf_output[2] ) );
  XOR2_X1 U6378 ( .A1(n5633), .A2(n5632), .Z(\MC_ARK_ARC_1_3/buf_output[176] )
         );
  XOR2_X1 U6380 ( .A1(\MC_ARK_ARC_1_3/temp1[176] ), .A2(n3703), .Z(n5632) );
  XOR2_X1 U6382 ( .A1(\MC_ARK_ARC_1_3/temp2[176] ), .A2(n3704), .Z(n5633) );
  NAND3_X1 U6383 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i1_7 ), .A3(\SB4_31/i3[0] ), 
        .ZN(n5634) );
  NAND4_X2 U6387 ( .A1(n4153), .A2(\SB2_4_29/Component_Function_3/NAND4_in[0] ), .A3(\SB2_4_29/Component_Function_3/NAND4_in[1] ), .A4(n5635), .ZN(
        \SB2_4_29/buf_output[3] ) );
  NAND3_X2 U6388 ( .A1(\SB2_4_29/i0[10] ), .A2(\SB2_4_29/i1[9] ), .A3(
        \SB2_4_29/i1_7 ), .ZN(n5635) );
  XOR2_X1 U6390 ( .A1(n5636), .A2(n155), .Z(Ciphertext[2]) );
  NAND4_X2 U6391 ( .A1(n2649), .A2(n3375), .A3(
        \SB4_31/Component_Function_2/NAND4_in[0] ), .A4(n5254), .ZN(n5636) );
  XOR2_X1 U6392 ( .A1(\MC_ARK_ARC_1_0/temp2[9] ), .A2(n5637), .Z(n1893) );
  XOR2_X1 U6393 ( .A1(n6488), .A2(n5638), .Z(n3025) );
  XOR2_X1 U6394 ( .A1(n575), .A2(\MC_ARK_ARC_1_3/buf_datainput[99] ), .Z(n5638) );
  NAND3_X1 U6396 ( .A1(\SB1_0_11/i0[10] ), .A2(\SB1_0_11/i1[9] ), .A3(
        \SB1_0_11/i1_7 ), .ZN(n5059) );
  NAND3_X2 U6397 ( .A1(\SB1_2_11/i1_5 ), .A2(\SB1_2_11/i1[9] ), .A3(
        \SB1_2_11/i0_4 ), .ZN(n1244) );
  XOR2_X1 U6399 ( .A1(n5640), .A2(n5639), .Z(\MC_ARK_ARC_1_4/temp5[179] ) );
  XOR2_X1 U6400 ( .A1(\RI5[4][179] ), .A2(\RI5[4][125] ), .Z(n5639) );
  XOR2_X1 U6402 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[173] ), .A2(\RI5[4][149] ), 
        .Z(n5640) );
  XOR2_X1 U6403 ( .A1(n2091), .A2(n5641), .Z(\MC_ARK_ARC_1_4/temp5[27] ) );
  XOR2_X1 U6404 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[27] ), .A2(\RI5[4][21] ), 
        .Z(n5641) );
  XOR2_X1 U6405 ( .A1(n5643), .A2(n5642), .Z(\MC_ARK_ARC_1_2/temp5[99] ) );
  XOR2_X1 U6408 ( .A1(\SB2_2_18/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[99] ), .Z(n5642) );
  XOR2_X1 U6410 ( .A1(\RI5[2][69] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .Z(n5643) );
  NAND4_X2 U6411 ( .A1(\SB4_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_19/Component_Function_0/NAND4_in[3] ), .A3(n4315), .A4(n5644), 
        .ZN(n7133) );
  NAND3_X1 U6412 ( .A1(\SB4_19/i0[6] ), .A2(\SB4_19/i0[8] ), .A3(
        \SB4_19/i0[7] ), .ZN(n5644) );
  NAND4_X2 U6413 ( .A1(\SB2_3_13/Component_Function_3/NAND4_in[2] ), .A2(n5179), .A3(\SB2_3_13/Component_Function_3/NAND4_in[3] ), .A4(n5645), .ZN(
        \RI5[3][123] ) );
  NAND3_X2 U6424 ( .A1(n6746), .A2(\SB2_3_13/i0_3 ), .A3(\SB2_3_13/i0_0 ), 
        .ZN(n5645) );
  NAND3_X1 U6426 ( .A1(\SB1_1_30/i0[8] ), .A2(\SB1_1_30/i1_7 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[10] ), .ZN(n1718) );
  NAND2_X1 U6428 ( .A1(\SB1_4_29/i3[0] ), .A2(n6531), .ZN(
        \SB1_4_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U6430 ( .A1(\SB1_3_7/i0[6] ), .A2(\SB1_3_7/i0[8] ), .A3(
        \SB1_3_7/i0[7] ), .ZN(\SB1_3_7/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U6431 ( .A1(\MC_ARK_ARC_1_0/temp2[19] ), .A2(
        \MC_ARK_ARC_1_0/temp1[19] ), .Z(\MC_ARK_ARC_1_0/temp5[19] ) );
  NAND4_X2 U6434 ( .A1(\SB2_1_12/Component_Function_3/NAND4_in[3] ), .A2(n5298), .A3(\SB2_1_12/Component_Function_3/NAND4_in[0] ), .A4(n5646), .ZN(
        \SB2_1_12/buf_output[3] ) );
  NAND3_X2 U6436 ( .A1(\SB2_1_12/i0_0 ), .A2(\SB2_1_12/i0_4 ), .A3(
        \SB2_1_12/i0_3 ), .ZN(n5646) );
  NAND4_X2 U6437 ( .A1(\SB2_4_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_4/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_4_4/Component_Function_2/NAND4_in[1] ), .A4(n5647), .ZN(
        \SB2_4_4/buf_output[2] ) );
  NAND3_X2 U6438 ( .A1(\SB2_4_4/i0_0 ), .A2(\SB2_4_4/i0_4 ), .A3(
        \SB2_4_4/i1_5 ), .ZN(n5647) );
  NAND3_X2 U6442 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0[8] ), .A3(\SB4_16/i0[9] ), .ZN(\SB4_16/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U6443 ( .A1(n5649), .A2(n5648), .Z(n5389) );
  XOR2_X1 U6448 ( .A1(\RI5[2][177] ), .A2(\RI5[2][39] ), .Z(n5648) );
  XOR2_X1 U6449 ( .A1(\RI5[2][9] ), .A2(\RI5[2][33] ), .Z(n5649) );
  XOR2_X1 U6450 ( .A1(\MC_ARK_ARC_1_4/temp5[46] ), .A2(n5650), .Z(
        \MC_ARK_ARC_1_4/buf_output[46] ) );
  XOR2_X1 U6457 ( .A1(\MC_ARK_ARC_1_4/temp4[46] ), .A2(
        \MC_ARK_ARC_1_4/temp3[46] ), .Z(n5650) );
  XOR2_X1 U6458 ( .A1(\MC_ARK_ARC_1_4/temp2[6] ), .A2(n5651), .Z(n3830) );
  XOR2_X1 U6460 ( .A1(\RI5[4][0] ), .A2(\RI5[4][6] ), .Z(n5651) );
  NAND4_X2 U6461 ( .A1(\SB2_4_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_19/Component_Function_0/NAND4_in[1] ), .A3(n6600), .A4(
        \SB2_4_19/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_4_19/buf_output[0] ) );
  XOR2_X1 U6463 ( .A1(\MC_ARK_ARC_1_3/temp1[146] ), .A2(n5652), .Z(
        \MC_ARK_ARC_1_3/temp5[146] ) );
  XOR2_X1 U6467 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), .A2(\RI5[3][92] ), 
        .Z(n5652) );
  NAND3_X1 U6471 ( .A1(\SB4_8/i0[9] ), .A2(\SB4_8/i0_4 ), .A3(\SB4_8/i0[6] ), 
        .ZN(\SB4_8/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U6474 ( .A1(n5653), .A2(n184), .Z(Ciphertext[52]) );
  NAND4_X2 U6475 ( .A1(\SB4_23/Component_Function_4/NAND4_in[3] ), .A2(n2695), 
        .A3(n2775), .A4(n5252), .ZN(n5653) );
  NAND4_X2 U6481 ( .A1(\SB3_13/Component_Function_0/NAND4_in[2] ), .A2(n1806), 
        .A3(\SB3_13/Component_Function_0/NAND4_in[0] ), .A4(
        \SB3_13/Component_Function_0/NAND4_in[1] ), .ZN(\SB3_13/buf_output[0] ) );
  NAND3_X2 U6482 ( .A1(\SB1_1_12/i0[9] ), .A2(\SB1_1_12/i0_4 ), .A3(
        \SB1_1_12/i0[6] ), .ZN(n7330) );
  NAND4_X2 U6492 ( .A1(\SB2_4_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_28/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_4_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_4_28/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_4_28/buf_output[3] ) );
  NAND4_X2 U6493 ( .A1(n2349), .A2(n6257), .A3(
        \SB2_4_29/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_4_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_4_29/buf_output[5] ) );
  NAND3_X2 U6496 ( .A1(\SB3_0/i0[9] ), .A2(\SB3_0/i0[8] ), .A3(\SB3_0/i0_3 ), 
        .ZN(n2556) );
  XOR2_X1 U6498 ( .A1(n7121), .A2(n7122), .Z(n6019) );
  NAND3_X1 U6502 ( .A1(\SB2_4_29/i0[10] ), .A2(\SB2_4_29/i0[6] ), .A3(
        \SB2_4_29/i0_3 ), .ZN(\SB2_4_29/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U6505 ( .A1(\SB1_3_23/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_23/Component_Function_2/NAND4_in[3] ), .A3(n5803), .A4(
        \SB1_3_23/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_3_23/buf_output[2] ) );
  NAND4_X2 U6506 ( .A1(\SB1_2_16/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_16/Component_Function_3/NAND4_in[0] ), .A3(n1270), .A4(n3812), 
        .ZN(\SB1_2_16/buf_output[3] ) );
  NAND4_X2 U6507 ( .A1(n935), .A2(n6911), .A3(
        \SB2_4_25/Component_Function_2/NAND4_in[0] ), .A4(n746), .ZN(
        \SB2_4_25/buf_output[2] ) );
  NAND4_X2 U6508 ( .A1(\SB2_0_8/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_0_8/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_0_8/Component_Function_4/NAND4_in[1] ), .A4(n7401), .ZN(
        \SB2_0_8/buf_output[4] ) );
  INV_X1 U6509 ( .I(\SB3_30/buf_output[2] ), .ZN(\SB4_27/i1[9] ) );
  NAND4_X2 U6512 ( .A1(\SB2_4_31/Component_Function_5/NAND4_in[1] ), .A2(n5655), .A3(\SB2_4_31/Component_Function_5/NAND4_in[0] ), .A4(n5654), .ZN(
        \SB2_4_31/buf_output[5] ) );
  NAND3_X2 U6513 ( .A1(\SB2_4_31/i0_4 ), .A2(\SB2_4_31/i0[6] ), .A3(
        \SB2_4_31/i0[9] ), .ZN(n5654) );
  NAND3_X2 U6515 ( .A1(\SB2_4_31/i0_3 ), .A2(\SB2_4_31/i0_4 ), .A3(
        \SB2_4_31/i1[9] ), .ZN(n5655) );
  NAND4_X2 U6518 ( .A1(\SB2_1_28/Component_Function_1/NAND4_in[0] ), .A2(n6803), .A3(\SB2_1_28/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_1_28/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_28/buf_output[1] ) );
  NAND4_X2 U6520 ( .A1(\SB3_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_4/Component_Function_3/NAND4_in[3] ), .A4(n5656), .ZN(
        \SB3_4/buf_output[3] ) );
  NAND3_X1 U6522 ( .A1(\SB3_4/i0[10] ), .A2(\SB3_4/i1_7 ), .A3(\SB3_4/i1[9] ), 
        .ZN(n5656) );
  XOR2_X1 U6525 ( .A1(n5657), .A2(n36), .Z(Ciphertext[26]) );
  XOR2_X1 U6530 ( .A1(n2803), .A2(n5658), .Z(\MC_ARK_ARC_1_2/buf_output[89] )
         );
  XOR2_X1 U6535 ( .A1(n7320), .A2(n6083), .Z(n5658) );
  NAND4_X2 U6536 ( .A1(n2821), .A2(\SB2_1_9/Component_Function_5/NAND4_in[0] ), 
        .A3(n5717), .A4(\SB2_1_9/Component_Function_5/NAND4_in[1] ), .ZN(
        \SB2_1_9/buf_output[5] ) );
  NAND3_X1 U6539 ( .A1(\SB1_4_15/i0_0 ), .A2(\SB1_4_15/i3[0] ), .A3(
        \SB1_4_15/i1_7 ), .ZN(\SB1_4_15/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U6546 ( .A1(n6659), .A2(\SB1_4_7/Component_Function_5/NAND4_in[3] ), 
        .A3(n5819), .A4(n6201), .ZN(\SB1_4_7/buf_output[5] ) );
  XOR2_X1 U6548 ( .A1(n5660), .A2(n5659), .Z(\MC_ARK_ARC_1_4/temp5[125] ) );
  XOR2_X1 U6549 ( .A1(\RI5[4][125] ), .A2(\RI5[4][119] ), .Z(n5659) );
  XOR2_X1 U6550 ( .A1(\RI5[4][95] ), .A2(\RI5[4][71] ), .Z(n5660) );
  XOR2_X1 U6552 ( .A1(n4894), .A2(n7233), .Z(\MC_ARK_ARC_1_4/buf_output[123] )
         );
  XOR2_X1 U6556 ( .A1(\MC_ARK_ARC_1_4/temp4[123] ), .A2(
        \MC_ARK_ARC_1_4/temp3[123] ), .Z(n4894) );
  NAND4_X2 U6564 ( .A1(\SB2_2_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_0/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_0/Component_Function_2/NAND4_in[1] ), .A4(n5661), .ZN(
        \SB2_2_0/buf_output[2] ) );
  NAND3_X2 U6565 ( .A1(\SB2_2_0/i0_0 ), .A2(\SB2_2_0/i1_5 ), .A3(n5444), .ZN(
        n5661) );
  XOR2_X1 U6568 ( .A1(\MC_ARK_ARC_1_2/temp1[93] ), .A2(n5662), .Z(n2371) );
  XOR2_X1 U6573 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[63] ), .A2(\RI5[2][39] ), 
        .Z(n5662) );
  XOR2_X1 U6576 ( .A1(\MC_ARK_ARC_1_4/temp4[189] ), .A2(n5663), .Z(n905) );
  XOR2_X1 U6577 ( .A1(\SB2_4_23/buf_output[3] ), .A2(\RI5[4][99] ), .Z(n5663)
         );
  XOR2_X1 U6578 ( .A1(n5664), .A2(n147), .Z(Ciphertext[98]) );
  NAND4_X2 U6579 ( .A1(\SB4_15/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_15/Component_Function_2/NAND4_in[0] ), .A3(n3880), .A4(
        \SB4_15/Component_Function_2/NAND4_in[1] ), .ZN(n5664) );
  NAND3_X2 U6580 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0[10] ), .A3(
        \SB2_3_26/i0[6] ), .ZN(\SB2_3_26/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U6582 ( .A1(n5666), .A2(n5665), .Z(\MC_ARK_ARC_1_3/buf_output[41] )
         );
  XOR2_X1 U6583 ( .A1(n6074), .A2(\MC_ARK_ARC_1_3/temp4[41] ), .Z(n5665) );
  XOR2_X1 U6584 ( .A1(n6075), .A2(n2193), .Z(n5666) );
  XOR2_X1 U6586 ( .A1(\RI5[2][158] ), .A2(\RI5[2][152] ), .Z(n5667) );
  NAND2_X1 U6587 ( .A1(\SB1_0_25/Component_Function_4/NAND4_in[3] ), .A2(n6616), .ZN(n931) );
  NAND4_X2 U6588 ( .A1(\SB2_0_8/Component_Function_5/NAND4_in[1] ), .A2(n2096), 
        .A3(\SB2_0_8/Component_Function_5/NAND4_in[0] ), .A4(n2097), .ZN(
        \SB2_0_8/buf_output[5] ) );
  NAND4_X2 U6589 ( .A1(n5754), .A2(\SB1_1_3/Component_Function_5/NAND4_in[1] ), 
        .A3(n7575), .A4(\SB1_1_3/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_3/buf_output[5] ) );
  XOR2_X1 U6591 ( .A1(\RI5[3][169] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[1] ), 
        .Z(n5668) );
  NAND3_X2 U6592 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i0_3 ), .A3(n590), .ZN(
        \SB2_1_0/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U6595 ( .A1(\MC_ARK_ARC_1_3/temp4[147] ), .A2(n5671), .Z(n6518) );
  XOR2_X1 U6598 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[147] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[141] ), .Z(n5671) );
  XOR2_X1 U6599 ( .A1(n5672), .A2(n63), .Z(Ciphertext[57]) );
  XOR2_X1 U6605 ( .A1(\MC_ARK_ARC_1_4/temp2[118] ), .A2(n5673), .Z(n3439) );
  XOR2_X1 U6610 ( .A1(\RI5[4][112] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[118] ), 
        .Z(n5673) );
  NAND3_X2 U6611 ( .A1(\SB1_3_16/i0_4 ), .A2(\SB1_3_16/i0[8] ), .A3(
        \SB1_3_16/i1_7 ), .ZN(n6304) );
  XOR2_X1 U6612 ( .A1(n5674), .A2(n132), .Z(Ciphertext[58]) );
  NAND4_X2 U6616 ( .A1(\SB4_22/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_22/Component_Function_4/NAND4_in[3] ), .A3(
        \SB4_22/Component_Function_4/NAND4_in[0] ), .A4(n3213), .ZN(n5674) );
  NAND3_X1 U6617 ( .A1(\SB1_2_13/i0[10] ), .A2(\SB1_2_13/i1[9] ), .A3(
        \SB1_2_13/i1_5 ), .ZN(\SB1_2_13/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U6619 ( .A1(n5675), .A2(\MC_ARK_ARC_1_2/temp4[80] ), .Z(
        \MC_ARK_ARC_1_2/temp6[80] ) );
  XOR2_X1 U6621 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), .A2(\RI5[2][182] ), 
        .Z(n5675) );
  NAND4_X2 U6622 ( .A1(\SB2_2_10/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_10/Component_Function_2/NAND4_in[1] ), .A3(n4192), .A4(n5676), 
        .ZN(\SB2_2_10/buf_output[2] ) );
  NAND3_X2 U6624 ( .A1(\SB2_2_10/i0_0 ), .A2(\SB2_2_10/i0_4 ), .A3(n589), .ZN(
        n5676) );
  XOR2_X1 U6626 ( .A1(n5677), .A2(n123), .Z(Ciphertext[59]) );
  NAND4_X2 U6627 ( .A1(\SB4_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_22/Component_Function_5/NAND4_in[1] ), .A3(n5961), .A4(
        \SB4_22/Component_Function_5/NAND4_in[0] ), .ZN(n5677) );
  NAND4_X2 U6629 ( .A1(\SB4_4/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_4/Component_Function_0/NAND4_in[1] ), .A3(n2684), .A4(n5678), 
        .ZN(n5686) );
  NAND3_X1 U6630 ( .A1(\SB4_4/i0_0 ), .A2(\SB4_4/i0_3 ), .A3(\SB4_4/i0[7] ), 
        .ZN(n5678) );
  XOR2_X1 U6632 ( .A1(n5679), .A2(n137), .Z(Ciphertext[122]) );
  NAND4_X2 U6634 ( .A1(n3023), .A2(n1696), .A3(n5260), .A4(
        \SB4_11/Component_Function_2/NAND4_in[2] ), .ZN(n5679) );
  XOR2_X1 U6635 ( .A1(n3464), .A2(n5680), .Z(n3491) );
  XOR2_X1 U6637 ( .A1(\RI5[3][175] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[7] ), 
        .Z(n5680) );
  XOR2_X1 U6639 ( .A1(n5681), .A2(\MC_ARK_ARC_1_0/temp4[107] ), .Z(n5983) );
  XOR2_X1 U6640 ( .A1(\RI5[0][17] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[173] ), 
        .Z(n5681) );
  NAND4_X2 U6642 ( .A1(\SB1_1_14/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_14/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_1_14/Component_Function_3/NAND4_in[2] ), .A4(n2712), .ZN(
        \SB1_1_14/buf_output[3] ) );
  INV_X2 U6643 ( .I(\SB1_3_3/buf_output[2] ), .ZN(\SB2_3_0/i1[9] ) );
  NAND4_X2 U6644 ( .A1(n7280), .A2(\SB1_3_3/Component_Function_2/NAND4_in[2] ), 
        .A3(n6541), .A4(\SB1_3_3/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_3_3/buf_output[2] ) );
  XOR2_X1 U6648 ( .A1(n6446), .A2(n5682), .Z(n3076) );
  XOR2_X1 U6649 ( .A1(\RI5[2][9] ), .A2(\RI5[2][33] ), .Z(n5682) );
  NAND4_X2 U6655 ( .A1(n2963), .A2(\SB2_1_19/Component_Function_5/NAND4_in[3] ), .A3(\SB2_1_19/Component_Function_5/NAND4_in[0] ), .A4(n5684), .ZN(
        \SB2_1_19/buf_output[5] ) );
  NAND3_X2 U6659 ( .A1(\SB2_1_19/i0[6] ), .A2(\SB2_1_19/i0_0 ), .A3(
        \SB2_1_19/i0[10] ), .ZN(n5684) );
  NAND4_X2 U6660 ( .A1(\SB1_0_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_0/NAND4_in[0] ), .A4(n5685), .ZN(
        \SB1_0_28/buf_output[0] ) );
  NAND3_X1 U6661 ( .A1(\SB1_0_28/i0[7] ), .A2(\SB1_0_28/i0_0 ), .A3(
        \SB1_0_28/i0_3 ), .ZN(n5685) );
  XOR2_X1 U6665 ( .A1(n5686), .A2(n2), .Z(Ciphertext[162]) );
  XOR2_X1 U6666 ( .A1(n5687), .A2(n209), .Z(Ciphertext[167]) );
  NAND4_X2 U6670 ( .A1(\SB4_4/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_4/Component_Function_5/NAND4_in[2] ), .A3(n5173), .A4(
        \SB4_4/Component_Function_5/NAND4_in[0] ), .ZN(n5687) );
  XOR2_X1 U6671 ( .A1(n4291), .A2(n5688), .Z(\MC_ARK_ARC_1_0/buf_output[99] )
         );
  XOR2_X1 U6672 ( .A1(n1713), .A2(n4204), .Z(n5688) );
  NAND4_X2 U6673 ( .A1(\SB3_6/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_6/Component_Function_3/NAND4_in[3] ), .A3(n6055), .A4(n5689), 
        .ZN(\SB3_6/buf_output[3] ) );
  NAND3_X1 U6681 ( .A1(\SB3_6/i0[6] ), .A2(\SB3_6/i1[9] ), .A3(\SB3_6/i0_3 ), 
        .ZN(n5689) );
  NAND4_X2 U6682 ( .A1(n4676), .A2(\SB2_4_22/Component_Function_2/NAND4_in[0] ), .A3(n7219), .A4(n3098), .ZN(\SB2_4_22/buf_output[2] ) );
  INV_X1 U6683 ( .I(\SB3_0/buf_output[1] ), .ZN(\SB4_28/i1_7 ) );
  NAND4_X2 U6684 ( .A1(\SB3_0/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_0/Component_Function_1/NAND4_in[1] ), .A3(n2769), .A4(n1575), 
        .ZN(\SB3_0/buf_output[1] ) );
  XOR2_X1 U6689 ( .A1(n5690), .A2(\MC_ARK_ARC_1_4/temp5[151] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[151] ) );
  XOR2_X1 U6690 ( .A1(\MC_ARK_ARC_1_4/temp4[151] ), .A2(
        \MC_ARK_ARC_1_4/temp3[151] ), .Z(n5690) );
  XOR2_X1 U6695 ( .A1(\MC_ARK_ARC_1_4/temp6[10] ), .A2(n5691), .Z(
        \MC_ARK_ARC_1_4/buf_output[10] ) );
  XOR2_X1 U6699 ( .A1(\MC_ARK_ARC_1_4/temp2[10] ), .A2(
        \MC_ARK_ARC_1_4/temp1[10] ), .Z(n5691) );
  INV_X2 U6704 ( .I(\SB1_3_26/buf_output[3] ), .ZN(\SB2_3_24/i0[8] ) );
  NAND4_X2 U6708 ( .A1(\SB1_3_26/Component_Function_3/NAND4_in[2] ), .A2(n7259), .A3(\SB1_3_26/Component_Function_3/NAND4_in[0] ), .A4(n3365), .ZN(
        \SB1_3_26/buf_output[3] ) );
  AND2_X1 U6712 ( .A1(n1562), .A2(n874), .Z(n572) );
  NAND4_X2 U6719 ( .A1(\SB1_2_18/Component_Function_3/NAND4_in[1] ), .A2(n6053), .A3(n7455), .A4(\SB1_2_18/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB1_2_18/buf_output[3] ) );
  XOR2_X1 U6725 ( .A1(n5693), .A2(n5692), .Z(n7349) );
  XOR2_X1 U6730 ( .A1(\RI5[4][113] ), .A2(n52), .Z(n5692) );
  XOR2_X1 U6733 ( .A1(\RI5[4][107] ), .A2(\RI5[4][83] ), .Z(n5693) );
  XOR2_X1 U6741 ( .A1(n5695), .A2(n5694), .Z(\MC_ARK_ARC_1_0/temp6[47] ) );
  XOR2_X1 U6746 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[113] ), .A2(n217), .Z(
        n5694) );
  XOR2_X1 U6747 ( .A1(\SB2_0_18/buf_output[5] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[149] ), .Z(n5695) );
  NAND3_X1 U6751 ( .A1(\SB1_0_21/i0_0 ), .A2(\SB1_0_21/i0_3 ), .A3(
        \SB1_0_21/i0[7] ), .ZN(\SB1_0_21/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U6755 ( .A1(\SB2_0_24/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_0_24/Component_Function_2/NAND4_in[0] ), .A3(n5800), .A4(
        \SB2_0_24/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_24/buf_output[2] ) );
  NAND3_X2 U6756 ( .A1(\SB1_1_7/i0[10] ), .A2(\SB1_1_7/i0_0 ), .A3(
        \SB1_1_7/i0[6] ), .ZN(\SB1_1_7/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U6758 ( .A1(\SB1_0_3/i0_4 ), .A2(\SB1_0_3/i1[9] ), .A3(
        \SB1_0_3/i0_3 ), .ZN(\SB1_0_3/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U6760 ( .A1(\SB1_1_9/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_9/Component_Function_3/NAND4_in[0] ), .A3(n2157), .A4(
        \SB1_1_9/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_1_9/buf_output[3] ) );
  NAND3_X2 U6763 ( .A1(\SB1_4_14/i0[6] ), .A2(\SB1_4_14/i0[10] ), .A3(
        \SB1_4_14/i0_3 ), .ZN(n6879) );
  NAND4_X2 U6765 ( .A1(\SB1_1_6/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_1_6/Component_Function_5/NAND4_in[2] ), .A3(n5740), .A4(n6937), 
        .ZN(\SB1_1_6/buf_output[5] ) );
  NAND4_X2 U6766 ( .A1(\SB2_1_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_14/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_14/Component_Function_2/NAND4_in[1] ), .A4(n1082), .ZN(
        \SB2_1_14/buf_output[2] ) );
  NAND3_X1 U6767 ( .A1(\SB1_2_18/i0[10] ), .A2(\SB1_2_18/i1[9] ), .A3(
        \SB1_2_18/i1_5 ), .ZN(n3554) );
  NAND3_X2 U6770 ( .A1(\SB2_1_25/i0_4 ), .A2(\SB2_1_25/i0_3 ), .A3(
        \SB2_1_25/i0_0 ), .ZN(\SB2_1_25/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 U6771 ( .I(\SB1_4_22/buf_output[5] ), .Z(\SB2_4_22/i0_3 ) );
  NAND3_X2 U6772 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0_4 ), .A3(
        \SB2_2_20/i1[9] ), .ZN(\SB2_2_20/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U6774 ( .A1(\RI5[1][116] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[146] ), 
        .Z(n6490) );
  NAND4_X2 U6779 ( .A1(\SB2_0_8/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_8/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_8/Component_Function_3/NAND4_in[1] ), .A4(n4571), .ZN(
        \SB2_0_8/buf_output[3] ) );
  XOR2_X1 U6780 ( .A1(n5697), .A2(n5696), .Z(\MC_ARK_ARC_1_3/buf_output[14] )
         );
  XOR2_X1 U6783 ( .A1(\MC_ARK_ARC_1_3/temp1[14] ), .A2(
        \MC_ARK_ARC_1_3/temp4[14] ), .Z(n5696) );
  XOR2_X1 U6784 ( .A1(\MC_ARK_ARC_1_3/temp3[14] ), .A2(
        \MC_ARK_ARC_1_3/temp2[14] ), .Z(n5697) );
  NAND4_X2 U6787 ( .A1(\SB2_0_23/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_23/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_23/Component_Function_2/NAND4_in[3] ), .A4(n5698), .ZN(
        \SB2_0_23/buf_output[2] ) );
  NAND3_X2 U6797 ( .A1(\SB2_0_23/i0[10] ), .A2(\SB2_0_23/i1[9] ), .A3(
        \SB2_0_23/i1_5 ), .ZN(n5698) );
  XOR2_X1 U6803 ( .A1(\MC_ARK_ARC_1_1/temp1[111] ), .A2(n5699), .Z(
        \MC_ARK_ARC_1_1/temp5[111] ) );
  XOR2_X1 U6804 ( .A1(\RI5[1][57] ), .A2(\RI5[1][81] ), .Z(n5699) );
  XOR2_X1 U6805 ( .A1(\MC_ARK_ARC_1_3/temp1[28] ), .A2(n5700), .Z(n6464) );
  XOR2_X1 U6811 ( .A1(\RI5[3][166] ), .A2(\RI5[3][190] ), .Z(n5700) );
  XOR2_X1 U6812 ( .A1(n5701), .A2(n15), .Z(Ciphertext[45]) );
  NAND4_X2 U6814 ( .A1(\SB2_0_6/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_0_6/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_6/Component_Function_4/NAND4_in[2] ), .A4(n5702), .ZN(
        \SB2_0_6/buf_output[4] ) );
  NAND2_X2 U6821 ( .A1(n5856), .A2(\SB2_0_6/i0_4 ), .ZN(n5702) );
  NAND4_X2 U6822 ( .A1(\SB2_4_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_4_2/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_4_2/Component_Function_1/NAND4_in[0] ), .A4(n5703), .ZN(
        \SB2_4_2/buf_output[1] ) );
  NAND4_X2 U6823 ( .A1(\SB2_3_23/Component_Function_2/NAND4_in[0] ), .A2(n1389), .A3(\SB2_3_23/Component_Function_2/NAND4_in[2] ), .A4(n6510), .ZN(
        \SB2_3_23/buf_output[2] ) );
  NAND3_X2 U6824 ( .A1(\SB1_3_23/i0[10] ), .A2(\SB1_3_23/i1[9] ), .A3(
        \SB1_3_23/i1_5 ), .ZN(n5803) );
  XOR2_X1 U6825 ( .A1(n5705), .A2(n5704), .Z(\MC_ARK_ARC_1_1/temp6[66] ) );
  XOR2_X1 U6826 ( .A1(\RI5[1][132] ), .A2(n560), .Z(n5704) );
  XOR2_X1 U6827 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[168] ), .A2(\RI5[1][102] ), 
        .Z(n5705) );
  XOR2_X1 U6830 ( .A1(n6389), .A2(n6388), .Z(n961) );
  NAND3_X2 U6832 ( .A1(\SB2_1_19/i0[6] ), .A2(\SB2_1_19/i0[9] ), .A3(
        \SB2_1_19/i0_4 ), .ZN(\SB2_1_19/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U6833 ( .A1(\SB2_3_11/Component_Function_5/NAND4_in[3] ), .A2(n2514), .A3(\SB2_3_11/Component_Function_5/NAND4_in[0] ), .A4(n5706), .ZN(
        \SB2_3_11/buf_output[5] ) );
  INV_X1 U6835 ( .I(\SB3_19/buf_output[1] ), .ZN(\SB4_15/i1_7 ) );
  NAND4_X2 U6836 ( .A1(\SB3_19/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_19/Component_Function_1/NAND4_in[1] ), .A3(n6779), .A4(
        \SB3_19/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_19/buf_output[1] ) );
  NAND4_X2 U6838 ( .A1(\SB1_4_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_7/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_4_7/Component_Function_0/NAND4_in[1] ), .A4(n5707), .ZN(
        \SB1_4_7/buf_output[0] ) );
  NAND3_X2 U6839 ( .A1(\SB1_4_7/i0_0 ), .A2(\SB1_4_7/i0_3 ), .A3(
        \SB1_4_7/i0[7] ), .ZN(n5707) );
  INV_X1 U6843 ( .I(\SB3_12/buf_output[3] ), .ZN(\SB4_10/i0[8] ) );
  NAND4_X2 U6852 ( .A1(n3480), .A2(\SB3_12/Component_Function_3/NAND4_in[3] ), 
        .A3(\SB3_12/Component_Function_3/NAND4_in[0] ), .A4(n5753), .ZN(
        \SB3_12/buf_output[3] ) );
  XOR2_X1 U6858 ( .A1(n5708), .A2(\MC_ARK_ARC_1_0/temp5[112] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[112] ) );
  XOR2_X1 U6859 ( .A1(\MC_ARK_ARC_1_0/temp4[112] ), .A2(
        \MC_ARK_ARC_1_0/temp3[112] ), .Z(n5708) );
  NAND2_X2 U6860 ( .A1(\SB1_0_18/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_18/Component_Function_4/NAND4_in[2] ), .ZN(n6493) );
  XOR2_X1 U6862 ( .A1(n3226), .A2(\MC_ARK_ARC_1_4/temp4[21] ), .Z(n4812) );
  INV_X2 U6868 ( .I(\SB3_15/buf_output[2] ), .ZN(\SB4_12/i1[9] ) );
  NAND4_X2 U6869 ( .A1(\SB3_15/Component_Function_2/NAND4_in[1] ), .A2(n6863), 
        .A3(n5718), .A4(\SB3_15/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB3_15/buf_output[2] ) );
  NAND4_X2 U6870 ( .A1(\SB1_1_8/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_8/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_8/Component_Function_0/NAND4_in[0] ), .A4(n5710), .ZN(
        \SB1_1_8/buf_output[0] ) );
  NAND3_X2 U6873 ( .A1(\SB1_1_8/i0[10] ), .A2(\SB1_1_8/i0_3 ), .A3(
        \SB1_1_8/i0_4 ), .ZN(n5710) );
  XOR2_X1 U6874 ( .A1(\MC_ARK_ARC_1_0/temp2[87] ), .A2(n5711), .Z(n6176) );
  XOR2_X1 U6878 ( .A1(\SB2_0_19/buf_output[3] ), .A2(\RI5[0][81] ), .Z(n5711)
         );
  XOR2_X1 U6881 ( .A1(n6322), .A2(n5712), .Z(n6453) );
  XOR2_X1 U6882 ( .A1(\RI5[1][173] ), .A2(\RI5[1][47] ), .Z(n5712) );
  NAND4_X2 U6883 ( .A1(\SB2_3_15/Component_Function_3/NAND4_in[3] ), .A2(n6685), .A3(\SB2_3_15/Component_Function_3/NAND4_in[0] ), .A4(n714), .ZN(
        \SB2_3_15/buf_output[3] ) );
  NAND3_X1 U6885 ( .A1(\SB1_4_13/i0_0 ), .A2(\SB1_4_13/i3[0] ), .A3(
        \SB1_4_13/i1_7 ), .ZN(\SB1_4_13/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U6889 ( .A1(n1029), .A2(n3067), .A3(n4288), .A4(n5713), .ZN(n5737)
         );
  NAND3_X2 U6890 ( .A1(\SB4_29/i0_4 ), .A2(\SB4_29/i0_0 ), .A3(\SB4_29/i0_3 ), 
        .ZN(n5713) );
  XOR2_X1 U6893 ( .A1(n5714), .A2(n4160), .Z(\MC_ARK_ARC_1_0/buf_output[92] )
         );
  XOR2_X1 U6894 ( .A1(n595), .A2(n5283), .Z(n5714) );
  XOR2_X1 U6895 ( .A1(\RI5[0][51] ), .A2(\RI5[0][57] ), .Z(
        \MC_ARK_ARC_1_0/temp1[57] ) );
  XOR2_X1 U6897 ( .A1(\RI5[3][121] ), .A2(\RI5[3][85] ), .Z(n5909) );
  NAND4_X2 U6909 ( .A1(\SB1_1_10/Component_Function_5/NAND4_in[1] ), .A2(n2589), .A3(\SB1_1_10/Component_Function_5/NAND4_in[0] ), .A4(n5715), .ZN(
        \SB1_1_10/buf_output[5] ) );
  NAND4_X2 U6914 ( .A1(\SB1_3_17/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_3_17/Component_Function_2/NAND4_in[1] ), .A3(n5215), .A4(n5716), 
        .ZN(\SB1_3_17/buf_output[2] ) );
  NAND3_X2 U6915 ( .A1(\SB2_1_27/i0[6] ), .A2(\SB2_1_27/i0[10] ), .A3(
        \SB2_1_27/i0_3 ), .ZN(\SB2_1_27/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U6916 ( .A1(n5346), .A2(\SB4_8/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB4_8/Component_Function_5/NAND4_in[0] ), .A4(n4858), .ZN(n7051)
         );
  XOR2_X1 U6919 ( .A1(\MC_ARK_ARC_1_4/temp4[125] ), .A2(
        \MC_ARK_ARC_1_4/temp3[125] ), .Z(\MC_ARK_ARC_1_4/temp6[125] ) );
  NAND4_X2 U6920 ( .A1(\SB2_0_8/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_0_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_8/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_0_8/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_0_8/buf_output[0] ) );
  NAND4_X2 U6922 ( .A1(\SB3_30/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_30/Component_Function_4/NAND4_in[3] ), .A3(n3749), .A4(
        \SB3_30/Component_Function_4/NAND4_in[0] ), .ZN(\SB3_30/buf_output[4] ) );
  INV_X2 U6924 ( .I(\SB1_2_29/buf_output[2] ), .ZN(\SB2_2_26/i1[9] ) );
  NAND4_X2 U6926 ( .A1(\SB1_2_29/Component_Function_2/NAND4_in[0] ), .A2(n3949), .A3(\SB1_2_29/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_2_29/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_2_29/buf_output[2] ) );
  NAND3_X2 U6927 ( .A1(\SB1_3_23/i0[8] ), .A2(\SB1_3_23/i1_5 ), .A3(
        \SB1_3_23/i3[0] ), .ZN(n6947) );
  NAND3_X2 U6928 ( .A1(\SB4_29/i0_4 ), .A2(\SB4_29/i0[10] ), .A3(\SB4_29/i0_3 ), .ZN(n7379) );
  NAND4_X2 U6935 ( .A1(\SB2_0_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_8/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_8/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_8/buf_output[2] ) );
  NAND3_X1 U6941 ( .A1(\SB2_4_17/i0[9] ), .A2(\SB2_4_17/i0[6] ), .A3(
        \SB1_4_18/buf_output[4] ), .ZN(n1016) );
  NAND3_X2 U6946 ( .A1(\SB2_1_9/i0[9] ), .A2(\SB2_1_9/i0_4 ), .A3(
        \SB2_1_9/i0[6] ), .ZN(n5717) );
  NAND3_X2 U6948 ( .A1(\SB3_15/i0[9] ), .A2(\SB3_15/i0_3 ), .A3(\SB3_15/i0[8] ), .ZN(n5718) );
  XOR2_X1 U6950 ( .A1(n5719), .A2(n55), .Z(Ciphertext[12]) );
  NAND4_X2 U6952 ( .A1(\SB4_29/Component_Function_0/NAND4_in[1] ), .A2(n5349), 
        .A3(n7379), .A4(\SB4_29/Component_Function_0/NAND4_in[0] ), .ZN(n5719)
         );
  NAND3_X1 U6954 ( .A1(\SB3_7/i0_0 ), .A2(\SB3_7/i3[0] ), .A3(\SB3_7/i1_7 ), 
        .ZN(n5720) );
  INV_X2 U6955 ( .I(\RI3[0][111] ), .ZN(\SB2_0_13/i0[8] ) );
  NAND4_X2 U6956 ( .A1(\SB1_0_15/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_15/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_15/Component_Function_3/NAND4_in[1] ), .A4(n6965), .ZN(
        \RI3[0][111] ) );
  INV_X1 U6958 ( .I(\SB3_23/buf_output[2] ), .ZN(\SB4_20/i1[9] ) );
  NAND4_X2 U6959 ( .A1(\SB3_23/Component_Function_2/NAND4_in[1] ), .A2(n5728), 
        .A3(n5859), .A4(\SB3_23/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB3_23/buf_output[2] ) );
  NAND4_X2 U6965 ( .A1(\SB1_3_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_7/Component_Function_5/NAND4_in[1] ), .A3(n7250), .A4(n4585), 
        .ZN(\SB1_3_7/buf_output[5] ) );
  XOR2_X1 U6966 ( .A1(\MC_ARK_ARC_1_3/temp5[58] ), .A2(n5721), .Z(
        \MC_ARK_ARC_1_3/buf_output[58] ) );
  XOR2_X1 U6972 ( .A1(\MC_ARK_ARC_1_3/temp3[58] ), .A2(
        \MC_ARK_ARC_1_3/temp4[58] ), .Z(n5721) );
  XOR2_X1 U6974 ( .A1(\SB2_1_17/buf_output[5] ), .A2(\RI5[1][53] ), .Z(n6760)
         );
  XOR2_X1 U6976 ( .A1(\MC_ARK_ARC_1_0/temp3[188] ), .A2(n5722), .Z(n4822) );
  XOR2_X1 U6977 ( .A1(\RI5[0][158] ), .A2(\RI5[0][134] ), .Z(n5722) );
  XOR2_X1 U6978 ( .A1(\RI5[0][168] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[102] ), 
        .Z(n1927) );
  NAND3_X1 U6983 ( .A1(\SB2_2_3/i0_4 ), .A2(\SB2_2_3/i1_7 ), .A3(n3991), .ZN(
        \SB2_2_3/Component_Function_1/NAND4_in[3] ) );
  NOR2_X2 U6984 ( .A1(n6113), .A2(n6112), .ZN(n3991) );
  XOR2_X1 U6987 ( .A1(\MC_ARK_ARC_1_1/temp6[140] ), .A2(n5723), .Z(
        \MC_ARK_ARC_1_1/buf_output[140] ) );
  NAND4_X2 U6992 ( .A1(\SB1_0_16/Component_Function_2/NAND4_in[1] ), .A2(n864), 
        .A3(\SB1_0_16/Component_Function_2/NAND4_in[3] ), .A4(n5724), .ZN(
        \RI3[0][110] ) );
  NAND3_X2 U6993 ( .A1(\SB1_0_16/i0[10] ), .A2(\SB1_0_16/i1[9] ), .A3(
        \SB1_0_16/i1_5 ), .ZN(n5724) );
  NAND3_X1 U6997 ( .A1(\SB3_11/i1[9] ), .A2(\SB3_11/i0_4 ), .A3(\SB3_11/i0_3 ), 
        .ZN(\SB3_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U6998 ( .A1(\SB2_1_19/i0[10] ), .A2(\SB2_1_19/i1_5 ), .A3(
        \SB2_1_19/i1[9] ), .ZN(\SB2_1_19/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U7009 ( .I(\SB2_2_13/buf_output[3] ), .Z(\RI5[2][123] ) );
  XOR2_X1 U7010 ( .A1(n3307), .A2(n5725), .Z(\MC_ARK_ARC_1_2/buf_output[9] )
         );
  XOR2_X1 U7011 ( .A1(\MC_ARK_ARC_1_2/temp4[9] ), .A2(n5825), .Z(n5725) );
  NAND3_X1 U7012 ( .A1(\SB1_2_16/i0_3 ), .A2(\SB1_2_16/i0_0 ), .A3(
        \SB1_2_16/i0_4 ), .ZN(\SB1_2_16/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U7013 ( .A1(\SB2_4_5/Component_Function_0/NAND4_in[1] ), .A2(n5726), 
        .A3(\SB2_4_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_4_5/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_4_5/buf_output[0] ) );
  NAND3_X2 U7015 ( .A1(\SB2_4_5/i0[7] ), .A2(\SB2_4_5/i0_0 ), .A3(
        \SB2_4_5/i0_3 ), .ZN(n5726) );
  XOR2_X1 U7017 ( .A1(\MC_ARK_ARC_1_3/temp5[158] ), .A2(n5727), .Z(
        \MC_ARK_ARC_1_3/buf_output[158] ) );
  XOR2_X1 U7021 ( .A1(\MC_ARK_ARC_1_3/temp4[158] ), .A2(
        \MC_ARK_ARC_1_3/temp3[158] ), .Z(n5727) );
  NAND3_X1 U7025 ( .A1(\SB4_11/i0_3 ), .A2(\SB4_11/i1[9] ), .A3(\SB4_11/i0[6] ), .ZN(n5729) );
  NAND3_X1 U7031 ( .A1(\SB4_7/i0[6] ), .A2(\SB4_7/i0_3 ), .A3(
        \SB3_9/buf_output[3] ), .ZN(n5730) );
  NAND4_X2 U7033 ( .A1(\SB2_2_28/Component_Function_4/NAND4_in[3] ), .A2(n7539), .A3(\SB2_2_28/Component_Function_4/NAND4_in[0] ), .A4(n5731), .ZN(
        \SB2_2_28/buf_output[4] ) );
  NAND3_X1 U7034 ( .A1(\SB2_2_28/i0_0 ), .A2(\SB2_2_28/i3[0] ), .A3(
        \SB2_2_28/i1_7 ), .ZN(n5731) );
  NAND4_X2 U7035 ( .A1(\SB1_1_2/Component_Function_5/NAND4_in[2] ), .A2(n836), 
        .A3(\SB1_1_2/Component_Function_5/NAND4_in[0] ), .A4(n5732), .ZN(
        \SB1_1_2/buf_output[5] ) );
  NAND3_X2 U7038 ( .A1(\SB1_1_2/i0_4 ), .A2(\SB1_1_2/i0[9] ), .A3(
        \SB1_1_2/i0[6] ), .ZN(n5732) );
  XOR2_X1 U7039 ( .A1(\SB2_2_14/buf_output[3] ), .A2(\RI5[2][111] ), .Z(
        \MC_ARK_ARC_1_2/temp1[117] ) );
  XOR2_X1 U7040 ( .A1(\MC_ARK_ARC_1_0/temp2[66] ), .A2(n5733), .Z(n2073) );
  XOR2_X1 U7042 ( .A1(\RI5[0][60] ), .A2(\RI5[0][66] ), .Z(n5733) );
  NAND4_X2 U7047 ( .A1(\SB2_2_15/Component_Function_3/NAND4_in[3] ), .A2(n1802), .A3(\SB2_2_15/Component_Function_3/NAND4_in[1] ), .A4(n5734), .ZN(
        \SB2_2_15/buf_output[3] ) );
  NAND3_X2 U7049 ( .A1(\SB2_2_15/i0[6] ), .A2(\SB2_2_15/i0_3 ), .A3(
        \SB2_2_15/i1[9] ), .ZN(n5734) );
  XOR2_X1 U7050 ( .A1(n5735), .A2(n21), .Z(Ciphertext[70]) );
  NAND4_X2 U7051 ( .A1(n3607), .A2(n2698), .A3(
        \SB4_20/Component_Function_4/NAND4_in[2] ), .A4(n6393), .ZN(n5735) );
  XOR2_X1 U7052 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[50] ), .A2(
        \SB2_1_22/buf_output[2] ), .Z(n4630) );
  XOR2_X1 U7056 ( .A1(n5736), .A2(n96), .Z(Ciphertext[187]) );
  NAND4_X2 U7059 ( .A1(\SB4_0/Component_Function_1/NAND4_in[1] ), .A2(n3046), 
        .A3(n4818), .A4(\SB4_0/Component_Function_1/NAND4_in[0] ), .ZN(n5736)
         );
  XOR2_X1 U7060 ( .A1(n5737), .A2(n208), .Z(Ciphertext[15]) );
  NAND4_X2 U7061 ( .A1(\SB1_1_23/Component_Function_3/NAND4_in[0] ), .A2(n2401), .A3(\SB1_1_23/Component_Function_3/NAND4_in[1] ), .A4(n4199), .ZN(
        \SB1_1_23/buf_output[3] ) );
  XOR2_X1 U7062 ( .A1(n3458), .A2(\MC_ARK_ARC_1_0/temp6[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[5] ) );
  XOR2_X1 U7072 ( .A1(\MC_ARK_ARC_1_0/temp2[5] ), .A2(
        \MC_ARK_ARC_1_0/temp1[5] ), .Z(n3458) );
  NAND3_X2 U7074 ( .A1(\SB2_1_21/i0_3 ), .A2(\SB2_1_21/i0[9] ), .A3(
        \SB2_1_21/i0[8] ), .ZN(\SB2_1_21/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U7077 ( .A1(n3651), .A2(n5738), .Z(\MC_ARK_ARC_1_4/temp5[122] ) );
  XOR2_X1 U7078 ( .A1(\RI5[4][116] ), .A2(\RI5[4][122] ), .Z(n5738) );
  XOR2_X1 U7080 ( .A1(\MC_ARK_ARC_1_4/temp2[123] ), .A2(
        \MC_ARK_ARC_1_4/temp1[123] ), .Z(n7233) );
  INV_X2 U7081 ( .I(\SB1_2_19/buf_output[2] ), .ZN(\SB2_2_16/i1[9] ) );
  NAND4_X2 U7084 ( .A1(\SB1_2_19/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_19/Component_Function_2/NAND4_in[2] ), .A3(n6893), .A4(n3016), 
        .ZN(\SB1_2_19/buf_output[2] ) );
  XOR2_X1 U7093 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[80] ), .A2(\RI5[3][104] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[134] ) );
  NAND3_X2 U7094 ( .A1(\SB1_4_19/i1_7 ), .A2(\SB1_4_19/i0[10] ), .A3(
        \SB1_4_19/i1[9] ), .ZN(n2039) );
  NAND3_X2 U7095 ( .A1(\SB4_29/i0_4 ), .A2(\SB4_29/i1_7 ), .A3(\SB4_29/i0[8] ), 
        .ZN(\SB4_29/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U7096 ( .A1(\SB1_2_27/Component_Function_2/NAND4_in[1] ), .A2(n4103), .A3(n4306), .A4(n5739), .ZN(\SB1_2_27/buf_output[2] ) );
  NAND3_X2 U7097 ( .A1(\SB1_2_27/i0_0 ), .A2(\SB1_2_27/i0_4 ), .A3(
        \SB1_2_27/i1_5 ), .ZN(n5739) );
  NAND3_X2 U7098 ( .A1(\SB1_1_6/i0[10] ), .A2(\SB1_1_6/i0_0 ), .A3(
        \SB1_1_6/i0[6] ), .ZN(n5740) );
  XOR2_X1 U7100 ( .A1(n5741), .A2(n183), .Z(Ciphertext[44]) );
  NAND4_X2 U7102 ( .A1(n2745), .A2(n3807), .A3(n897), .A4(n6431), .ZN(n5741)
         );
  XOR2_X1 U7104 ( .A1(n2375), .A2(n5742), .Z(\MC_ARK_ARC_1_1/buf_output[182] )
         );
  XOR2_X1 U7122 ( .A1(\MC_ARK_ARC_1_1/temp3[182] ), .A2(
        \MC_ARK_ARC_1_1/temp4[182] ), .Z(n5742) );
  XOR2_X1 U7125 ( .A1(n5744), .A2(n5743), .Z(\MC_ARK_ARC_1_1/buf_output[45] )
         );
  XOR2_X1 U7128 ( .A1(\MC_ARK_ARC_1_1/temp3[45] ), .A2(n1574), .Z(n5743) );
  XOR2_X1 U7129 ( .A1(\MC_ARK_ARC_1_1/temp2[45] ), .A2(
        \MC_ARK_ARC_1_1/temp4[45] ), .Z(n5744) );
  NAND4_X2 U7134 ( .A1(\SB1_3_21/Component_Function_5/NAND4_in[2] ), .A2(n6854), .A3(\SB1_3_21/Component_Function_5/NAND4_in[1] ), .A4(n5745), .ZN(
        \SB1_3_21/buf_output[5] ) );
  NAND4_X2 U7140 ( .A1(n4351), .A2(n6059), .A3(n1224), .A4(n5747), .ZN(
        \SB2_1_7/buf_output[3] ) );
  NAND3_X2 U7143 ( .A1(\SB2_1_7/i0_4 ), .A2(\SB2_1_7/i0_0 ), .A3(
        \SB2_1_7/i0_3 ), .ZN(n5747) );
  XOR2_X1 U7145 ( .A1(\MC_ARK_ARC_1_3/temp4[33] ), .A2(n5748), .Z(n7130) );
  NAND4_X2 U7147 ( .A1(n7216), .A2(\SB2_3_17/Component_Function_3/NAND4_in[0] ), .A3(n1933), .A4(n5749), .ZN(\SB2_3_17/buf_output[3] ) );
  XOR2_X1 U7151 ( .A1(n5750), .A2(n75), .Z(Ciphertext[111]) );
  XOR2_X1 U7156 ( .A1(n5752), .A2(n5751), .Z(\MC_ARK_ARC_1_1/buf_output[50] )
         );
  XOR2_X1 U7160 ( .A1(\MC_ARK_ARC_1_1/temp3[50] ), .A2(n7168), .Z(n5751) );
  XOR2_X1 U7161 ( .A1(\MC_ARK_ARC_1_1/temp1[50] ), .A2(
        \MC_ARK_ARC_1_1/temp4[50] ), .Z(n5752) );
  INV_X2 U7163 ( .I(\SB3_19/buf_output[2] ), .ZN(\SB4_16/i1[9] ) );
  NAND4_X2 U7168 ( .A1(\SB3_19/Component_Function_2/NAND4_in[1] ), .A2(n5847), 
        .A3(\SB3_19/Component_Function_2/NAND4_in[3] ), .A4(n6387), .ZN(
        \SB3_19/buf_output[2] ) );
  NAND3_X2 U7169 ( .A1(\SB3_12/i0[10] ), .A2(\SB3_12/i1_7 ), .A3(
        \SB3_12/i1[9] ), .ZN(n5753) );
  NAND4_X2 U7175 ( .A1(\SB2_3_5/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_5/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_3_5/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_5/buf_output[1] ) );
  INV_X2 U7176 ( .I(\SB1_1_10/buf_output[3] ), .ZN(\SB2_1_8/i0[8] ) );
  NAND4_X2 U7184 ( .A1(\SB1_1_10/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_10/Component_Function_3/NAND4_in[2] ), .A3(n6718), .A4(n5309), 
        .ZN(\SB1_1_10/buf_output[3] ) );
  XOR2_X1 U7186 ( .A1(\MC_ARK_ARC_1_3/temp1[9] ), .A2(n5755), .Z(
        \MC_ARK_ARC_1_3/temp5[9] ) );
  XOR2_X1 U7191 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[147] ), .A2(\RI5[3][171] ), 
        .Z(n5755) );
  XOR2_X1 U7194 ( .A1(\RI5[4][95] ), .A2(\RI5[4][29] ), .Z(n3478) );
  NAND3_X1 U7200 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i0_4 ), .A3(
        \SB2_2_27/i1[9] ), .ZN(n4100) );
  INV_X2 U7206 ( .I(\SB1_4_4/buf_output[2] ), .ZN(\SB2_4_1/i1[9] ) );
  NAND4_X2 U7209 ( .A1(\SB1_4_4/Component_Function_2/NAND4_in[0] ), .A2(n2246), 
        .A3(n1428), .A4(\SB1_4_4/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_4_4/buf_output[2] ) );
  NAND4_X2 U7219 ( .A1(\SB1_2_19/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_19/Component_Function_5/NAND4_in[1] ), .A3(n4257), .A4(
        \SB1_2_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_19/buf_output[5] ) );
  XOR2_X1 U7220 ( .A1(n5756), .A2(n80), .Z(Ciphertext[5]) );
  NAND4_X2 U7221 ( .A1(\SB4_31/Component_Function_5/NAND4_in[1] ), .A2(n2881), 
        .A3(\SB4_31/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_31/Component_Function_5/NAND4_in[0] ), .ZN(n5756) );
  NAND4_X2 U7222 ( .A1(\SB3_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_20/Component_Function_3/NAND4_in[2] ), .A3(n7240), .A4(n5757), 
        .ZN(\SB3_20/buf_output[3] ) );
  NAND3_X2 U7223 ( .A1(\SB3_20/i0_4 ), .A2(\SB3_20/i0_0 ), .A3(\SB3_20/i0_3 ), 
        .ZN(n5757) );
  XOR2_X1 U7229 ( .A1(n2976), .A2(\MC_ARK_ARC_1_4/temp6[38] ), .Z(n6287) );
  XOR2_X1 U7233 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), .A2(\RI5[3][152] ), 
        .Z(n2209) );
  XOR2_X1 U7237 ( .A1(n5759), .A2(n5758), .Z(\MC_ARK_ARC_1_2/buf_output[119] )
         );
  XOR2_X1 U7238 ( .A1(n6006), .A2(\MC_ARK_ARC_1_2/temp4[119] ), .Z(n5758) );
  NAND4_X2 U7240 ( .A1(\SB2_0_15/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_15/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_0_15/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_0_15/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_15/buf_output[0] ) );
  INV_X2 U7241 ( .I(\SB1_3_11/buf_output[3] ), .ZN(\SB2_3_9/i0[8] ) );
  NAND4_X2 U7242 ( .A1(n2134), .A2(\SB1_3_11/Component_Function_3/NAND4_in[1] ), .A3(n6897), .A4(n7423), .ZN(\SB1_3_11/buf_output[3] ) );
  XOR2_X1 U7247 ( .A1(n5760), .A2(n152), .Z(Ciphertext[14]) );
  NAND4_X2 U7248 ( .A1(n852), .A2(n3763), .A3(
        \SB4_29/Component_Function_2/NAND4_in[0] ), .A4(
        \SB4_29/Component_Function_2/NAND4_in[2] ), .ZN(n5760) );
  NAND4_X2 U7255 ( .A1(\SB2_4_7/Component_Function_2/NAND4_in[0] ), .A2(n1712), 
        .A3(n5762), .A4(n5761), .ZN(\SB2_4_7/buf_output[2] ) );
  NAND3_X2 U7257 ( .A1(\RI3[4][148] ), .A2(\SB2_4_7/i0_0 ), .A3(\SB2_4_7/i1_5 ), .ZN(n5761) );
  NAND4_X2 U7258 ( .A1(n2101), .A2(\SB2_4_6/Component_Function_5/NAND4_in[0] ), 
        .A3(n7120), .A4(n5763), .ZN(\SB2_4_6/buf_output[5] ) );
  NAND3_X2 U7259 ( .A1(\SB2_4_6/i0[10] ), .A2(\SB2_4_6/i0[6] ), .A3(
        \SB2_4_6/i0_0 ), .ZN(n5763) );
  XOR2_X1 U7264 ( .A1(n5764), .A2(n162), .Z(Ciphertext[92]) );
  NAND4_X2 U7265 ( .A1(n1321), .A2(\SB4_16/Component_Function_2/NAND4_in[2] ), 
        .A3(n6133), .A4(n3188), .ZN(n5764) );
  XOR2_X1 U7268 ( .A1(\MC_ARK_ARC_1_4/temp5[171] ), .A2(n5765), .Z(
        \MC_ARK_ARC_1_4/buf_output[171] ) );
  XOR2_X1 U7271 ( .A1(\MC_ARK_ARC_1_4/temp3[171] ), .A2(
        \MC_ARK_ARC_1_4/temp4[171] ), .Z(n5765) );
  XOR2_X1 U7277 ( .A1(n5767), .A2(n5766), .Z(n5845) );
  XOR2_X1 U7280 ( .A1(\RI5[0][172] ), .A2(n117), .Z(n5766) );
  XOR2_X1 U7281 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[70] ), .A2(\RI5[0][100] ), 
        .Z(n5767) );
  XOR2_X1 U7282 ( .A1(n5769), .A2(n5768), .Z(\MC_ARK_ARC_1_2/buf_output[182] )
         );
  XOR2_X1 U7283 ( .A1(n5997), .A2(\MC_ARK_ARC_1_2/temp4[182] ), .Z(n5768) );
  XOR2_X1 U7286 ( .A1(\MC_ARK_ARC_1_2/temp1[182] ), .A2(
        \MC_ARK_ARC_1_2/temp3[182] ), .Z(n5769) );
  NAND3_X1 U7288 ( .A1(\SB4_0/i0_3 ), .A2(\SB4_0/i0[6] ), .A3(\SB4_0/i1[9] ), 
        .ZN(n2977) );
  XOR2_X1 U7290 ( .A1(n5770), .A2(n31), .Z(Ciphertext[182]) );
  NAND4_X2 U7291 ( .A1(n7030), .A2(n4224), .A3(
        \SB4_1/Component_Function_2/NAND4_in[0] ), .A4(n2558), .ZN(n5770) );
  XOR2_X1 U7293 ( .A1(\MC_ARK_ARC_1_2/temp5[27] ), .A2(
        \MC_ARK_ARC_1_2/temp6[27] ), .Z(\MC_ARK_ARC_1_2/buf_output[27] ) );
  XOR2_X1 U7302 ( .A1(n5772), .A2(n5771), .Z(n3862) );
  XOR2_X1 U7303 ( .A1(\RI5[0][11] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[113] ), 
        .Z(n5771) );
  XOR2_X1 U7308 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[77] ), .A2(\RI5[0][5] ), 
        .Z(n5772) );
  XOR2_X1 U7311 ( .A1(n5774), .A2(n5773), .Z(n3271) );
  XOR2_X1 U7318 ( .A1(\RI5[1][41] ), .A2(\RI5[1][161] ), .Z(n5773) );
  XOR2_X1 U7320 ( .A1(\RI5[1][65] ), .A2(\RI5[1][5] ), .Z(n5774) );
  NAND3_X1 U7321 ( .A1(\SB1_2_28/i0_0 ), .A2(\SB1_2_28/i0[7] ), .A3(
        \SB1_2_28/i0_3 ), .ZN(\SB1_2_28/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X8 U7323 ( .I(\RI3[0][93] ), .Z(n6976) );
  XOR2_X1 U7324 ( .A1(\MC_ARK_ARC_1_3/temp6[164] ), .A2(n2197), .Z(
        \MC_ARK_ARC_1_3/buf_output[164] ) );
  NAND3_X2 U7325 ( .A1(\SB2_2_31/i0[10] ), .A2(\SB2_2_31/i0_0 ), .A3(
        \SB2_2_31/i0[6] ), .ZN(n2071) );
  NAND4_X2 U7326 ( .A1(\SB1_2_1/Component_Function_3/NAND4_in[0] ), .A2(n4959), 
        .A3(n6093), .A4(n4958), .ZN(\SB1_2_1/buf_output[3] ) );
  XOR2_X1 U7327 ( .A1(n3499), .A2(n3424), .Z(n7451) );
  NAND4_X2 U7331 ( .A1(\SB2_0_19/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_0_19/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_19/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_0_19/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_0_19/buf_output[2] ) );
  NAND4_X2 U7333 ( .A1(\SB2_2_23/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_23/Component_Function_5/NAND4_in[3] ), .A3(n6159), .A4(
        \SB2_2_23/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_23/buf_output[5] ) );
  AND2_X1 U7334 ( .A1(n1836), .A2(n5317), .Z(n2890) );
  NAND4_X2 U7335 ( .A1(\SB1_4_18/Component_Function_3/NAND4_in[1] ), .A2(n2577), .A3(n6904), .A4(n5775), .ZN(\SB1_4_18/buf_output[3] ) );
  XOR2_X1 U7336 ( .A1(\SB2_1_22/buf_output[5] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[83] ), .Z(n4235) );
  BUF_X4 U7340 ( .I(\MC_ARK_ARC_1_4/buf_output[118] ), .Z(\SB3_12/i0_4 ) );
  NAND3_X2 U7341 ( .A1(\SB2_2_15/i0[6] ), .A2(\SB2_2_15/i0[10] ), .A3(
        \SB2_2_15/i0_0 ), .ZN(\SB2_2_15/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U7342 ( .A1(\SB1_4_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_19/Component_Function_4/NAND4_in[2] ), .A3(n6492), .A4(
        \SB1_4_19/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_4_19/buf_output[4] ) );
  NAND4_X2 U7343 ( .A1(\SB1_2_17/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_2_17/Component_Function_3/NAND4_in[0] ), .A3(n6795), .A4(
        \SB1_2_17/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_17/buf_output[3] ) );
  NAND3_X1 U7344 ( .A1(\SB2_1_18/i0_0 ), .A2(\SB2_1_18/i3[0] ), .A3(
        \SB2_1_18/i1_7 ), .ZN(\SB2_1_18/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U7348 ( .A1(\RI5[2][101] ), .A2(\RI5[2][155] ), .Z(n818) );
  XOR2_X1 U7357 ( .A1(\RI5[4][0] ), .A2(\RI5[4][186] ), .Z(
        \MC_ARK_ARC_1_4/temp1[0] ) );
  NAND3_X2 U7359 ( .A1(\SB1_3_28/i0_3 ), .A2(\SB1_3_28/i0[8] ), .A3(
        \SB1_3_28/i1_7 ), .ZN(\SB1_3_28/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U7360 ( .A1(n5776), .A2(\MC_ARK_ARC_1_0/temp6[139] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[139] ) );
  XOR2_X1 U7364 ( .A1(\MC_ARK_ARC_1_0/temp1[139] ), .A2(
        \MC_ARK_ARC_1_0/temp2[139] ), .Z(n5776) );
  NAND2_X2 U7365 ( .A1(n5423), .A2(n5777), .ZN(\SB2_3_13/i0_4 ) );
  AND2_X1 U7366 ( .A1(n2202), .A2(n2486), .Z(n5777) );
  XOR2_X1 U7369 ( .A1(\MC_ARK_ARC_1_1/temp2[114] ), .A2(n5778), .Z(
        \MC_ARK_ARC_1_1/temp5[114] ) );
  XOR2_X1 U7371 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[108] ), .A2(\RI5[1][114] ), 
        .Z(n5778) );
  NAND4_X2 U7372 ( .A1(\SB2_0_14/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_0_14/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_0_14/Component_Function_4/NAND4_in[0] ), .A4(n5779), .ZN(
        \SB2_0_14/buf_output[4] ) );
  NAND3_X1 U7379 ( .A1(\SB2_0_14/i0[10] ), .A2(\SB2_0_14/i0_3 ), .A3(
        \SB2_0_14/i0[9] ), .ZN(n5779) );
  NAND4_X2 U7381 ( .A1(n1075), .A2(\SB1_3_25/Component_Function_5/NAND4_in[3] ), .A3(\SB1_3_25/Component_Function_5/NAND4_in[0] ), .A4(n6412), .ZN(
        \SB1_3_25/buf_output[5] ) );
  INV_X2 U7382 ( .I(\SB1_4_18/buf_output[3] ), .ZN(\SB2_4_16/i0[8] ) );
  XOR2_X1 U7385 ( .A1(n5780), .A2(n28), .Z(Ciphertext[114]) );
  NAND4_X2 U7386 ( .A1(\SB4_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_12/Component_Function_0/NAND4_in[3] ), .A3(n5936), .A4(
        \SB4_12/Component_Function_0/NAND4_in[1] ), .ZN(n5780) );
  NAND3_X2 U7389 ( .A1(\SB2_0_21/i1[9] ), .A2(\SB2_0_21/i1_5 ), .A3(
        \SB2_0_21/i0[10] ), .ZN(\SB2_0_21/Component_Function_2/NAND4_in[0] )
         );
  NAND4_X2 U7396 ( .A1(n2240), .A2(\SB2_1_2/Component_Function_5/NAND4_in[2] ), 
        .A3(\SB2_1_2/Component_Function_5/NAND4_in[0] ), .A4(n5781), .ZN(
        \SB2_1_2/buf_output[5] ) );
  NAND4_X2 U7397 ( .A1(\SB1_1_24/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_1_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_24/Component_Function_1/NAND4_in[0] ), .A4(n5782), .ZN(
        \SB1_1_24/buf_output[1] ) );
  NAND3_X2 U7398 ( .A1(\SB1_1_24/i0_4 ), .A2(\SB1_1_24/i0[8] ), .A3(
        \SB1_1_24/i1_7 ), .ZN(n5782) );
  NAND3_X1 U7399 ( .A1(\SB3_5/i0[8] ), .A2(\SB3_5/i0_3 ), .A3(\SB3_5/i1_7 ), 
        .ZN(\SB3_5/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U7401 ( .A1(\SB2_1_2/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_2/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_2/Component_Function_0/NAND4_in[0] ), .A4(n5783), .ZN(
        \SB2_1_2/buf_output[0] ) );
  NAND3_X2 U7404 ( .A1(\SB2_0_14/i3[0] ), .A2(\SB2_0_14/i1_5 ), .A3(
        \SB2_0_14/i0[8] ), .ZN(\SB2_0_14/Component_Function_3/NAND4_in[3] ) );
  NAND2_X2 U7405 ( .A1(n4940), .A2(n5784), .ZN(n6548) );
  NAND3_X2 U7406 ( .A1(\SB2_4_15/i0[10] ), .A2(\SB2_4_15/i1_5 ), .A3(
        \SB2_4_15/i1[9] ), .ZN(n5784) );
  XOR2_X1 U7407 ( .A1(\MC_ARK_ARC_1_2/temp5[191] ), .A2(n5785), .Z(
        \RI1[3][191] ) );
  XOR2_X1 U7408 ( .A1(\MC_ARK_ARC_1_2/temp4[191] ), .A2(n6666), .Z(n5785) );
  NAND3_X2 U7411 ( .A1(\SB2_2_13/i0_0 ), .A2(\SB2_2_13/i1_5 ), .A3(
        \SB2_2_13/i0_4 ), .ZN(\SB2_2_13/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U7413 ( .A1(\SB3_7/Component_Function_2/NAND4_in[3] ), .A2(
        \SB3_7/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_7/Component_Function_2/NAND4_in[1] ), .A4(n5786), .ZN(
        \SB3_7/buf_output[2] ) );
  NAND3_X2 U7416 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i1[9] ), .A3(\SB3_7/i1_5 ), 
        .ZN(n5786) );
  XOR2_X1 U7418 ( .A1(\MC_ARK_ARC_1_3/temp6[78] ), .A2(n5787), .Z(
        \MC_ARK_ARC_1_3/buf_output[78] ) );
  XOR2_X1 U7419 ( .A1(\MC_ARK_ARC_1_3/temp1[78] ), .A2(
        \MC_ARK_ARC_1_3/temp2[78] ), .Z(n5787) );
  XOR2_X1 U7422 ( .A1(n5789), .A2(n5788), .Z(\MC_ARK_ARC_1_4/buf_output[93] )
         );
  XOR2_X1 U7425 ( .A1(\MC_ARK_ARC_1_4/temp4[93] ), .A2(n1049), .Z(n5788) );
  XOR2_X1 U7426 ( .A1(\MC_ARK_ARC_1_4/temp2[93] ), .A2(
        \MC_ARK_ARC_1_4/temp1[93] ), .Z(n5789) );
  NAND4_X2 U7429 ( .A1(\SB2_4_12/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_4_12/Component_Function_3/NAND4_in[0] ), .A3(n5127), .A4(
        \SB2_4_12/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_4_12/buf_output[3] ) );
  XOR2_X1 U7430 ( .A1(n5790), .A2(\MC_ARK_ARC_1_2/temp4[75] ), .Z(n4250) );
  XOR2_X1 U7436 ( .A1(\SB2_2_10/buf_output[3] ), .A2(\RI5[2][177] ), .Z(n5790)
         );
  NAND4_X2 U7438 ( .A1(\SB1_2_11/Component_Function_2/NAND4_in[0] ), .A2(n4777), .A3(n6494), .A4(n5791), .ZN(\SB1_2_11/buf_output[2] ) );
  XOR2_X1 U7442 ( .A1(\RI5[3][138] ), .A2(\RI5[3][162] ), .Z(
        \MC_ARK_ARC_1_3/temp2[0] ) );
  XOR2_X1 U7444 ( .A1(n5792), .A2(n179), .Z(Ciphertext[135]) );
  NAND4_X2 U7447 ( .A1(n2298), .A2(n7050), .A3(n7173), .A4(n3140), .ZN(n5792)
         );
  INV_X2 U7450 ( .I(\SB1_1_15/buf_output[2] ), .ZN(\SB2_1_12/i1[9] ) );
  NAND4_X2 U7451 ( .A1(\SB1_1_15/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_15/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_1_15/Component_Function_2/NAND4_in[0] ), .A4(n2455), .ZN(
        \SB1_1_15/buf_output[2] ) );
  NAND4_X2 U7452 ( .A1(n4672), .A2(n6923), .A3(
        \SB2_3_15/Component_Function_5/NAND4_in[0] ), .A4(n5793), .ZN(
        \SB2_3_15/buf_output[5] ) );
  NAND3_X2 U7453 ( .A1(\SB2_3_15/i0[10] ), .A2(\SB2_3_15/i0[6] ), .A3(
        \SB2_3_15/i0_0 ), .ZN(n5793) );
  NAND3_X2 U7454 ( .A1(\SB2_0_14/i0_3 ), .A2(\SB2_0_14/i0[8] ), .A3(
        \SB2_0_14/i0[9] ), .ZN(\SB2_0_14/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U7457 ( .A1(\SB2_4_23/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_23/Component_Function_0/NAND4_in[0] ), .A4(n5794), .ZN(
        \SB2_4_23/buf_output[0] ) );
  NAND3_X1 U7458 ( .A1(\SB2_4_23/i0_0 ), .A2(\SB2_4_23/i0_3 ), .A3(
        \SB2_4_23/i0[7] ), .ZN(n5794) );
  XOR2_X1 U7460 ( .A1(\MC_ARK_ARC_1_2/temp2[124] ), .A2(n5795), .Z(
        \MC_ARK_ARC_1_2/temp5[124] ) );
  XOR2_X1 U7461 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[124] ), .A2(\RI5[2][118] ), 
        .Z(n5795) );
  XOR2_X1 U7463 ( .A1(n5796), .A2(n134), .Z(Ciphertext[106]) );
  NAND4_X2 U7464 ( .A1(n7536), .A2(n7301), .A3(n2490), .A4(
        \SB4_14/Component_Function_4/NAND4_in[2] ), .ZN(n5796) );
  NAND3_X2 U7468 ( .A1(\SB2_2_22/i0[6] ), .A2(\SB2_2_22/i0_3 ), .A3(
        \SB2_2_22/i0[10] ), .ZN(n675) );
  XOR2_X1 U7469 ( .A1(n5797), .A2(n218), .Z(Ciphertext[160]) );
  NAND4_X2 U7470 ( .A1(\SB4_5/Component_Function_4/NAND4_in[1] ), .A2(
        \SB4_5/Component_Function_4/NAND4_in[0] ), .A3(n7387), .A4(n7006), 
        .ZN(n5797) );
  INV_X1 U7471 ( .I(\SB3_12/buf_output[2] ), .ZN(\SB4_9/i1[9] ) );
  NAND4_X2 U7476 ( .A1(n6996), .A2(\SB3_12/Component_Function_2/NAND4_in[0] ), 
        .A3(n6486), .A4(n1069), .ZN(\SB3_12/buf_output[2] ) );
  NAND4_X2 U7477 ( .A1(n3031), .A2(\SB2_2_5/Component_Function_5/NAND4_in[1] ), 
        .A3(n5798), .A4(\SB2_2_5/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_5/buf_output[5] ) );
  NAND3_X2 U7478 ( .A1(\SB2_2_5/i0[9] ), .A2(\SB2_2_5/i0[6] ), .A3(
        \SB2_2_5/i0_4 ), .ZN(n5798) );
  NAND4_X2 U7481 ( .A1(\SB2_2_5/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_5/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_2_5/Component_Function_1/NAND4_in[3] ), .A4(n5799), .ZN(
        \SB2_2_5/buf_output[1] ) );
  XOR2_X1 U7486 ( .A1(n6865), .A2(\MC_ARK_ARC_1_3/temp5[35] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[35] ) );
  NAND3_X1 U7487 ( .A1(\SB2_0_24/i0[6] ), .A2(\SB2_0_24/i0[10] ), .A3(
        \SB2_0_24/i0_3 ), .ZN(n5800) );
  XOR2_X1 U7489 ( .A1(n4048), .A2(n5801), .Z(n7022) );
  XOR2_X1 U7491 ( .A1(\RI5[2][51] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .Z(n5801) );
  NAND4_X2 U7492 ( .A1(\SB3_27/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_27/Component_Function_5/NAND4_in[1] ), .A3(n7335), .A4(
        \SB3_27/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_27/buf_output[5] ) );
  NAND4_X2 U7498 ( .A1(\SB2_4_10/Component_Function_5/NAND4_in[2] ), .A2(n1043), .A3(n7487), .A4(n5802), .ZN(\SB2_4_10/buf_output[5] ) );
  NAND2_X2 U7500 ( .A1(\SB2_4_10/i0_0 ), .A2(\SB2_4_10/i3[0] ), .ZN(n5802) );
  XOR2_X1 U7505 ( .A1(\MC_ARK_ARC_1_2/temp4[100] ), .A2(n5804), .Z(n2814) );
  XOR2_X1 U7506 ( .A1(\RI5[2][166] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[10] ), 
        .Z(n5804) );
  XOR2_X1 U7509 ( .A1(\SB2_3_13/buf_output[0] ), .A2(\SB2_3_19/buf_output[0] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[36] ) );
  XOR2_X1 U7510 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[157] ), .A2(\RI5[3][181] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[19] ) );
  XOR2_X1 U7512 ( .A1(\RI5[3][98] ), .A2(\RI5[3][134] ), .Z(
        \MC_ARK_ARC_1_3/temp3[32] ) );
  XOR2_X1 U7513 ( .A1(\MC_ARK_ARC_1_4/temp4[152] ), .A2(n5805), .Z(n3134) );
  XOR2_X1 U7515 ( .A1(\RI5[4][62] ), .A2(\RI5[4][26] ), .Z(n5805) );
  NAND4_X2 U7516 ( .A1(\SB2_4_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_4_28/Component_Function_2/NAND4_in[2] ), .A4(n5806), .ZN(
        \SB2_4_28/buf_output[2] ) );
  XOR2_X1 U7519 ( .A1(n5807), .A2(n143), .Z(Ciphertext[112]) );
  NAND4_X2 U7521 ( .A1(\SB4_13/Component_Function_4/NAND4_in[2] ), .A2(n1214), 
        .A3(\SB4_13/Component_Function_4/NAND4_in[3] ), .A4(n1216), .ZN(n5807)
         );
  NAND4_X2 U7523 ( .A1(\SB1_2_16/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_16/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_16/Component_Function_0/NAND4_in[1] ), .A4(n5808), .ZN(
        \SB1_2_16/buf_output[0] ) );
  XOR2_X1 U7524 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[177] ), .A2(\RI5[3][171] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[177] ) );
  NAND4_X2 U7526 ( .A1(\SB1_1_25/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_25/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_1_25/Component_Function_3/NAND4_in[0] ), .A4(n5809), .ZN(
        \SB1_1_25/buf_output[3] ) );
  XOR2_X1 U7527 ( .A1(\MC_ARK_ARC_1_2/temp6[125] ), .A2(n5810), .Z(
        \MC_ARK_ARC_1_2/buf_output[125] ) );
  XOR2_X1 U7532 ( .A1(\MC_ARK_ARC_1_2/temp1[125] ), .A2(n7435), .Z(n5810) );
  NAND3_X2 U7533 ( .A1(\SB2_0_27/i0_0 ), .A2(\SB2_0_27/i0[10] ), .A3(
        \SB2_0_27/i0[6] ), .ZN(n4487) );
  NAND3_X2 U7534 ( .A1(\SB1_4_27/i0_4 ), .A2(\RI1[4][26] ), .A3(
        \SB1_4_27/i1_5 ), .ZN(n3069) );
  NAND4_X2 U7537 ( .A1(\SB1_3_3/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_3/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_3_3/Component_Function_4/NAND4_in[2] ), .A4(n5811), .ZN(
        \SB1_3_3/buf_output[4] ) );
  XOR2_X1 U7538 ( .A1(n5813), .A2(n5812), .Z(n906) );
  XOR2_X1 U7541 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[135] ), .A2(\RI5[4][189] ), 
        .Z(n5812) );
  XOR2_X1 U7545 ( .A1(\RI5[4][159] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[183] ), 
        .Z(n5813) );
  NAND3_X2 U7551 ( .A1(\SB2_3_12/i0[9] ), .A2(\SB2_3_12/i0_3 ), .A3(
        \SB2_3_12/i0[8] ), .ZN(n7478) );
  NAND3_X2 U7552 ( .A1(\SB3_13/i1_5 ), .A2(\SB3_13/i0_0 ), .A3(\SB3_13/i0_4 ), 
        .ZN(n7064) );
  NAND3_X2 U7553 ( .A1(\SB1_2_30/i0_0 ), .A2(\SB1_2_30/i1_5 ), .A3(
        \SB1_2_30/i0_4 ), .ZN(n3963) );
  NAND3_X1 U7554 ( .A1(\SB1_2_20/i0_3 ), .A2(\MC_ARK_ARC_1_1/buf_output[66] ), 
        .A3(\SB1_2_20/i0[8] ), .ZN(\SB1_2_20/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U7557 ( .I(\SB2_3_0/buf_output[5] ), .Z(\RI5[3][191] ) );
  NAND3_X2 U7562 ( .A1(\SB2_3_9/i0_3 ), .A2(\SB2_3_9/i0[6] ), .A3(
        \SB2_3_9/i1[9] ), .ZN(\SB2_3_9/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U7564 ( .I(\SB1_4_21/buf_output[5] ), .Z(\SB2_4_21/i0_3 ) );
  NAND4_X2 U7568 ( .A1(n5851), .A2(n6433), .A3(n2844), .A4(n6032), .ZN(
        \SB2_2_9/buf_output[2] ) );
  XOR2_X1 U7573 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[176] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[170] ), .Z(\MC_ARK_ARC_1_3/temp1[176] )
         );
  XOR2_X1 U7574 ( .A1(\RI5[3][117] ), .A2(\RI5[3][93] ), .Z(n5948) );
  NOR2_X2 U7576 ( .A1(n5815), .A2(n5814), .ZN(n4002) );
  NAND2_X1 U7577 ( .A1(n4876), .A2(\SB3_13/Component_Function_5/NAND4_in[0] ), 
        .ZN(n5814) );
  NAND3_X1 U7578 ( .A1(\SB2_3_2/i0_4 ), .A2(\SB2_3_2/i0[9] ), .A3(
        \SB1_3_6/buf_output[1] ), .ZN(
        \SB2_3_2/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U7579 ( .A1(\SB1_3_1/i0[6] ), .A2(\SB1_3_1/i0[10] ), .A3(
        \SB1_3_1/i0_0 ), .ZN(n5816) );
  NAND4_X2 U7580 ( .A1(\SB1_3_14/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_14/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_14/Component_Function_5/NAND4_in[2] ), .A4(n5180), .ZN(
        \SB1_3_14/buf_output[5] ) );
  NAND4_X2 U7585 ( .A1(\SB1_1_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_3/NAND4_in[1] ), .A3(n5836), .A4(n6429), 
        .ZN(\SB1_1_29/buf_output[3] ) );
  XOR2_X1 U7586 ( .A1(\RI5[2][129] ), .A2(\RI5[2][153] ), .Z(n4025) );
  XOR2_X1 U7594 ( .A1(\RI5[4][80] ), .A2(\RI5[4][56] ), .Z(
        \MC_ARK_ARC_1_4/temp2[110] ) );
  XOR2_X1 U7596 ( .A1(\RI5[0][104] ), .A2(\RI5[0][110] ), .Z(
        \MC_ARK_ARC_1_0/temp1[110] ) );
  XOR2_X1 U7597 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[14] ), .A2(\RI5[2][80] ), 
        .Z(n7310) );
  XOR2_X1 U7601 ( .A1(n6317), .A2(n5817), .Z(\MC_ARK_ARC_1_4/buf_output[101] )
         );
  XOR2_X1 U7603 ( .A1(n7551), .A2(\MC_ARK_ARC_1_4/temp4[101] ), .Z(n5817) );
  NAND4_X2 U7612 ( .A1(\SB2_4_21/Component_Function_2/NAND4_in[2] ), .A2(n6539), .A3(\SB2_4_21/Component_Function_2/NAND4_in[0] ), .A4(n4159), .ZN(
        \SB2_4_21/buf_output[2] ) );
  NAND3_X2 U7614 ( .A1(\SB1_4_25/i0_3 ), .A2(\SB1_4_25/i0_0 ), .A3(
        \SB1_4_25/i0_4 ), .ZN(\SB1_4_25/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U7615 ( .A1(n5818), .A2(n204), .Z(Ciphertext[39]) );
  NAND4_X2 U7622 ( .A1(n2042), .A2(\SB4_25/Component_Function_3/NAND4_in[1] ), 
        .A3(n2840), .A4(\SB4_25/Component_Function_3/NAND4_in[3] ), .ZN(n5818)
         );
  NAND3_X2 U7628 ( .A1(\SB1_4_7/i0[10] ), .A2(\SB1_4_7/i0_0 ), .A3(
        \SB1_4_7/i0[6] ), .ZN(n5819) );
  NAND3_X2 U7629 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i0[6] ), .A3(
        \SB2_3_24/i1[9] ), .ZN(\SB2_3_24/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U7630 ( .I(\SB1_1_16/buf_output[5] ), .ZN(\SB2_1_16/i1_5 ) );
  NAND4_X2 U7632 ( .A1(\SB1_1_16/Component_Function_5/NAND4_in[2] ), .A2(n6041), .A3(n2764), .A4(\SB1_1_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_16/buf_output[5] ) );
  XOR2_X1 U7633 ( .A1(n5820), .A2(n116), .Z(Ciphertext[13]) );
  NAND4_X2 U7634 ( .A1(\SB4_29/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_29/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_29/Component_Function_1/NAND4_in[3] ), .A4(
        \SB4_29/Component_Function_1/NAND4_in[0] ), .ZN(n5820) );
  XOR2_X1 U7637 ( .A1(n5087), .A2(n5821), .Z(n5424) );
  XOR2_X1 U7638 ( .A1(n2759), .A2(n2760), .Z(n5821) );
  XOR2_X1 U7639 ( .A1(\RI5[0][83] ), .A2(\RI5[0][47] ), .Z(
        \MC_ARK_ARC_1_0/temp3[173] ) );
  NAND3_X1 U7643 ( .A1(\SB2_3_3/i0_3 ), .A2(\SB2_3_3/i0[10] ), .A3(
        \SB2_3_3/i0[9] ), .ZN(\SB2_3_3/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U7645 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), .A2(\RI5[2][5] ), 
        .Z(n3265) );
  INV_X2 U7646 ( .I(\SB1_2_9/buf_output[5] ), .ZN(\SB2_2_9/i1_5 ) );
  XOR2_X1 U7647 ( .A1(n5822), .A2(\MC_ARK_ARC_1_2/temp1[70] ), .Z(n1882) );
  XOR2_X1 U7652 ( .A1(\RI5[2][16] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[40] ), 
        .Z(n5822) );
  INV_X1 U7653 ( .I(\SB1_3_14/buf_output[1] ), .ZN(\SB2_3_10/i1_7 ) );
  NAND4_X2 U7655 ( .A1(\SB1_3_14/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_3_14/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_14/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_3_14/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_14/buf_output[1] ) );
  NAND4_X2 U7663 ( .A1(\SB2_4_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_0/Component_Function_3/NAND4_in[3] ), .A3(n4145), .A4(n5823), 
        .ZN(\SB2_4_0/buf_output[3] ) );
  NAND3_X2 U7670 ( .A1(\SB2_4_0/i0_4 ), .A2(\SB2_4_0/i0_3 ), .A3(
        \SB2_4_0/i0_0 ), .ZN(n5823) );
  NAND4_X2 U7675 ( .A1(\SB2_2_30/Component_Function_4/NAND4_in[1] ), .A2(n7567), .A3(\SB2_2_30/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_2_30/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_2_30/buf_output[4] ) );
  INV_X1 U7676 ( .I(\SB1_2_15/buf_output[5] ), .ZN(\SB2_2_15/i1_5 ) );
  NAND4_X2 U7679 ( .A1(\SB1_2_15/Component_Function_5/NAND4_in[3] ), .A2(n2833), .A3(n5940), .A4(\SB1_2_15/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_15/buf_output[5] ) );
  NAND3_X1 U7680 ( .A1(\SB1_1_2/i0[8] ), .A2(\SB1_1_2/i3[0] ), .A3(
        \SB1_1_2/i1_5 ), .ZN(\SB1_1_2/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U7681 ( .A1(\SB1_4_18/Component_Function_5/NAND4_in[2] ), .A2(n6123), .A3(\SB1_4_18/Component_Function_5/NAND4_in[0] ), .A4(n5824), .ZN(
        \SB1_4_18/buf_output[5] ) );
  NAND3_X2 U7683 ( .A1(\SB1_4_18/i0[6] ), .A2(\SB1_4_18/i0[9] ), .A3(
        \SB1_4_18/i0_4 ), .ZN(n5824) );
  NAND3_X2 U7686 ( .A1(\SB2_4_1/i0[10] ), .A2(n6277), .A3(\SB2_4_1/i1[9] ), 
        .ZN(\SB2_4_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U7688 ( .A1(\SB3_30/i0[10] ), .A2(\SB3_30/i1_7 ), .A3(
        \SB3_30/i1[9] ), .ZN(n2312) );
  XOR2_X1 U7689 ( .A1(\RI5[2][75] ), .A2(\RI5[2][111] ), .Z(n5825) );
  XOR2_X1 U7690 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[70] ), .A2(\RI5[0][106] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[4] ) );
  NAND3_X2 U7692 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0[9] ), .A3(
        \SB2_2_20/i0[10] ), .ZN(n681) );
  XOR2_X1 U7696 ( .A1(\MC_ARK_ARC_1_3/temp4[102] ), .A2(
        \MC_ARK_ARC_1_3/temp2[102] ), .Z(n604) );
  XOR2_X1 U7698 ( .A1(n2330), .A2(n5827), .Z(\MC_ARK_ARC_1_2/buf_output[40] )
         );
  XOR2_X1 U7700 ( .A1(\MC_ARK_ARC_1_2/temp4[40] ), .A2(
        \MC_ARK_ARC_1_2/temp3[40] ), .Z(n5827) );
  NAND3_X2 U7704 ( .A1(\SB1_2_21/i0[9] ), .A2(\SB1_2_21/i0_3 ), .A3(
        \SB1_2_21/i0[10] ), .ZN(n6579) );
  NAND3_X2 U7705 ( .A1(\SB2_0_1/i0[10] ), .A2(\SB2_0_1/i1[9] ), .A3(
        \SB2_0_1/i1_7 ), .ZN(\SB2_0_1/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U7706 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[23] ), .A2(\RI5[4][149] ), 
        .Z(n5828) );
  NAND4_X2 U7709 ( .A1(\SB3_13/Component_Function_1/NAND4_in[1] ), .A2(n5032), 
        .A3(n2399), .A4(\SB3_13/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB3_13/buf_output[1] ) );
  XOR2_X1 U7714 ( .A1(n4175), .A2(n5829), .Z(n4112) );
  XOR2_X1 U7715 ( .A1(\RI5[4][185] ), .A2(\RI5[4][191] ), .Z(n5829) );
  NAND3_X2 U7718 ( .A1(\SB2_4_1/i0[10] ), .A2(\SB2_4_1/i1_7 ), .A3(
        \SB2_4_1/i1[9] ), .ZN(n7426) );
  XOR2_X1 U7721 ( .A1(\MC_ARK_ARC_1_3/temp6[165] ), .A2(n5830), .Z(
        \MC_ARK_ARC_1_3/buf_output[165] ) );
  XOR2_X1 U7723 ( .A1(\MC_ARK_ARC_1_3/temp2[165] ), .A2(n3728), .Z(n5830) );
  NAND3_X2 U7725 ( .A1(\SB2_4_22/i0_4 ), .A2(\SB2_4_22/i0_3 ), .A3(
        \SB2_4_22/i1[9] ), .ZN(\SB2_4_22/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U7726 ( .A1(\SB1_4_16/Component_Function_5/NAND4_in[1] ), .A2(n3136), .A3(n6845), .A4(n4361), .ZN(\SB1_4_16/buf_output[5] ) );
  NAND4_X2 U7728 ( .A1(\SB2_3_15/Component_Function_0/NAND4_in[1] ), .A2(n6672), .A3(\SB2_3_15/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_15/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_15/buf_output[0] ) );
  BUF_X4 U7732 ( .I(\SB3_14/buf_output[4] ), .Z(\SB4_13/i0_4 ) );
  NAND3_X2 U7733 ( .A1(\SB2_0_21/i1[9] ), .A2(\SB2_0_21/i1_7 ), .A3(
        \SB2_0_21/i0[10] ), .ZN(n3253) );
  NAND4_X2 U7738 ( .A1(\SB2_4_27/Component_Function_3/NAND4_in[2] ), .A2(n1429), .A3(n5861), .A4(\SB2_4_27/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB2_4_27/buf_output[3] ) );
  XOR2_X1 U7739 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[29] ), .Z(n1236) );
  NAND3_X1 U7741 ( .A1(n320), .A2(\SB1_0_30/i1[9] ), .A3(\SB1_0_30/i0_3 ), 
        .ZN(\SB1_0_30/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7742 ( .A1(n4698), .A2(\MC_ARK_ARC_1_4/temp4[2] ), .Z(n3003) );
  NAND4_X2 U7744 ( .A1(\SB1_2_12/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_2_12/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_12/Component_Function_4/NAND4_in[1] ), .A4(n2915), .ZN(
        \SB1_2_12/buf_output[4] ) );
  XOR2_X1 U7745 ( .A1(n6578), .A2(n1090), .Z(n5165) );
  NAND3_X2 U7746 ( .A1(\SB2_4_23/i0_3 ), .A2(\SB2_4_23/i0[9] ), .A3(
        \SB2_4_23/i0[8] ), .ZN(\SB2_4_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U7750 ( .A1(\SB4_13/i0_0 ), .A2(\SB3_15/buf_output[3] ), .A3(
        \SB4_13/i0[6] ), .ZN(\SB4_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U7752 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i1_7 ), .A3(
        \SB4_28/i1[9] ), .ZN(\SB4_28/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U7757 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[77] ), .A2(\RI5[4][71] ), 
        .Z(\MC_ARK_ARC_1_4/temp1[77] ) );
  NAND3_X2 U7758 ( .A1(\SB2_3_6/i0[10] ), .A2(\SB2_3_6/i0_0 ), .A3(
        \SB2_3_6/i0[6] ), .ZN(n5401) );
  NAND3_X2 U7764 ( .A1(\SB2_2_24/i0[9] ), .A2(\SB2_2_24/i0_4 ), .A3(
        \SB2_2_24/i0[6] ), .ZN(n6343) );
  XOR2_X1 U7767 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[75] ), .A2(\RI5[0][81] ), 
        .Z(n2487) );
  NAND4_X2 U7768 ( .A1(\SB3_30/Component_Function_5/NAND4_in[1] ), .A2(n2585), 
        .A3(\SB3_30/Component_Function_5/NAND4_in[0] ), .A4(n5832), .ZN(
        \SB3_30/buf_output[5] ) );
  NAND3_X2 U7771 ( .A1(\SB3_30/i0[6] ), .A2(\SB3_30/i0[9] ), .A3(\SB3_30/i0_4 ), .ZN(n5832) );
  NAND3_X2 U7772 ( .A1(\SB3_19/i0[9] ), .A2(\SB3_19/i0_3 ), .A3(\SB3_19/i0[8] ), .ZN(n5847) );
  NAND4_X2 U7773 ( .A1(n1866), .A2(n5392), .A3(n7444), .A4(n3288), .ZN(
        \SB2_3_4/buf_output[5] ) );
  NAND4_X2 U7776 ( .A1(\SB1_4_22/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_4_22/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_4_22/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_4_22/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_4_22/buf_output[2] ) );
  XOR2_X1 U7778 ( .A1(\RI5[3][161] ), .A2(\RI5[3][137] ), .Z(n3073) );
  NAND4_X2 U7781 ( .A1(\SB3_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_16/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_2/NAND4_in[2] ), .A4(n6179), .ZN(
        \SB3_16/buf_output[2] ) );
  XOR2_X1 U7783 ( .A1(\RI5[3][61] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[37] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[91] ) );
  XOR2_X1 U7785 ( .A1(n1851), .A2(n5833), .Z(\MC_ARK_ARC_1_2/temp5[75] ) );
  XOR2_X1 U7786 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[45] ), .A2(\RI5[2][21] ), 
        .Z(n5833) );
  NAND3_X1 U7788 ( .A1(\SB2_2_26/i0_0 ), .A2(\SB2_2_26/i0_3 ), .A3(
        \SB2_2_26/i0[7] ), .ZN(n2322) );
  XOR2_X1 U7794 ( .A1(\MC_ARK_ARC_1_2/temp2[81] ), .A2(
        \MC_ARK_ARC_1_2/temp1[81] ), .Z(\MC_ARK_ARC_1_2/temp5[81] ) );
  NAND4_X2 U7795 ( .A1(\SB2_2_18/Component_Function_2/NAND4_in[0] ), .A2(n4174), .A3(\SB2_2_18/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_18/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_18/buf_output[2] ) );
  XOR2_X1 U7799 ( .A1(\MC_ARK_ARC_1_4/temp4[6] ), .A2(
        \MC_ARK_ARC_1_4/temp3[6] ), .Z(n796) );
  XOR2_X1 U7800 ( .A1(\RI5[3][110] ), .A2(\RI5[3][86] ), .Z(
        \MC_ARK_ARC_1_3/temp2[140] ) );
  XOR2_X1 U7801 ( .A1(n5834), .A2(\MC_ARK_ARC_1_3/temp4[24] ), .Z(
        \MC_ARK_ARC_1_3/temp6[24] ) );
  XOR2_X1 U7803 ( .A1(\RI5[3][126] ), .A2(\RI5[3][90] ), .Z(n5834) );
  NAND4_X2 U7805 ( .A1(\SB1_4_8/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_8/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_4_8/Component_Function_0/NAND4_in[1] ), .A4(n5835), .ZN(
        \SB1_4_8/buf_output[0] ) );
  NAND3_X1 U7811 ( .A1(\SB1_4_8/i0_0 ), .A2(\SB1_4_8/i0_3 ), .A3(
        \SB1_4_8/i0[7] ), .ZN(n5835) );
  NAND3_X2 U7813 ( .A1(\SB1_2_25/i0[10] ), .A2(\SB1_2_25/i0_0 ), .A3(
        \SB1_2_25/i0[6] ), .ZN(\SB1_2_25/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U7816 ( .A1(\RI5[3][161] ), .A2(\RI5[3][125] ), .Z(n4986) );
  NAND4_X2 U7819 ( .A1(\SB1_0_12/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_12/Component_Function_5/NAND4_in[0] ), .A3(n2414), .A4(n2413), 
        .ZN(\SB1_0_12/buf_output[5] ) );
  NAND3_X1 U7820 ( .A1(\SB2_2_0/i1[9] ), .A2(\SB1_2_0/buf_output[5] ), .A3(
        n5444), .ZN(\SB2_2_0/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U7824 ( .A1(\SB1_1_29/i0[8] ), .A2(\SB1_1_29/i1_5 ), .A3(
        \SB1_1_29/i3[0] ), .ZN(n5836) );
  NAND3_X2 U7825 ( .A1(\SB2_3_13/i0[6] ), .A2(\SB2_3_13/i0[9] ), .A3(
        \SB2_3_13/i0_4 ), .ZN(n6069) );
  NAND3_X2 U7827 ( .A1(\SB1_2_9/i0_0 ), .A2(\SB1_2_9/i0[10] ), .A3(
        \SB1_2_9/i0[6] ), .ZN(n5837) );
  XOR2_X1 U7829 ( .A1(\MC_ARK_ARC_1_0/temp3[86] ), .A2(n5838), .Z(n7570) );
  XOR2_X1 U7830 ( .A1(\RI5[0][56] ), .A2(\RI5[0][32] ), .Z(n5838) );
  XOR2_X1 U7840 ( .A1(\RI5[0][55] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[31] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[85] ) );
  NAND4_X2 U7841 ( .A1(\SB2_2_31/Component_Function_1/NAND4_in[1] ), .A2(n4366), .A3(\SB2_2_31/Component_Function_1/NAND4_in[0] ), .A4(n5839), .ZN(
        \SB2_2_31/buf_output[1] ) );
  NAND3_X2 U7844 ( .A1(\SB2_2_31/i0[9] ), .A2(\SB2_2_31/i1_5 ), .A3(
        \SB2_2_31/i0[6] ), .ZN(n5839) );
  NAND4_X2 U7848 ( .A1(n3517), .A2(n7321), .A3(n6828), .A4(n5840), .ZN(
        \SB2_4_11/buf_output[5] ) );
  NAND3_X2 U7849 ( .A1(\SB2_4_11/i0[9] ), .A2(\SB2_4_11/i0[6] ), .A3(
        \SB1_4_12/buf_output[4] ), .ZN(n5840) );
  XOR2_X1 U7853 ( .A1(n5841), .A2(n217), .Z(Ciphertext[118]) );
  NAND4_X2 U7855 ( .A1(n1726), .A2(n7522), .A3(
        \SB4_12/Component_Function_4/NAND4_in[1] ), .A4(
        \SB4_12/Component_Function_4/NAND4_in[3] ), .ZN(n5841) );
  NAND4_X2 U7856 ( .A1(\SB1_3_15/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_15/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_3_15/Component_Function_4/NAND4_in[0] ), .A4(n5842), .ZN(
        \SB1_3_15/buf_output[4] ) );
  NAND3_X1 U7857 ( .A1(\SB1_3_15/i0_4 ), .A2(n5431), .A3(\SB1_3_15/i1_5 ), 
        .ZN(n5842) );
  XOR2_X1 U7858 ( .A1(\MC_ARK_ARC_1_1/temp3[121] ), .A2(n5843), .Z(n5872) );
  XOR2_X1 U7861 ( .A1(\RI5[1][67] ), .A2(\RI5[1][121] ), .Z(n5843) );
  INV_X2 U7866 ( .I(\SB1_2_23/buf_output[2] ), .ZN(\SB2_2_20/i1[9] ) );
  NAND4_X2 U7868 ( .A1(\SB1_2_23/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_23/Component_Function_2/NAND4_in[1] ), .A3(n2403), .A4(
        \SB1_2_23/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_2_23/buf_output[2] ) );
  XOR2_X1 U7875 ( .A1(n2080), .A2(n5844), .Z(\MC_ARK_ARC_1_4/temp5[8] ) );
  XOR2_X1 U7877 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[170] ), .A2(\RI5[4][146] ), 
        .Z(n5844) );
  XOR2_X1 U7878 ( .A1(n7078), .A2(n7079), .Z(\MC_ARK_ARC_1_3/temp6[148] ) );
  NAND3_X2 U7879 ( .A1(\SB1_4_7/i0_4 ), .A2(\SB1_4_7/i0[9] ), .A3(
        \SB1_4_7/i0[6] ), .ZN(\SB1_4_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U7880 ( .A1(\SB1_4_16/i0_3 ), .A2(\SB1_4_16/i1[9] ), .A3(
        \SB1_4_16/i0[6] ), .ZN(n3236) );
  XOR2_X1 U7882 ( .A1(n3430), .A2(n5845), .Z(\MC_ARK_ARC_1_0/buf_output[34] )
         );
  NAND4_X2 U7890 ( .A1(\SB2_1_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_19/Component_Function_2/NAND4_in[1] ), .A3(n2733), .A4(n5846), 
        .ZN(\SB2_1_19/buf_output[2] ) );
  NAND3_X2 U7892 ( .A1(\SB2_1_19/i0[9] ), .A2(\SB2_1_19/i0_3 ), .A3(
        \SB2_1_19/i0[8] ), .ZN(n5846) );
  INV_X2 U7898 ( .I(\SB1_1_1/buf_output[2] ), .ZN(\SB2_1_30/i1[9] ) );
  NAND4_X2 U7899 ( .A1(\SB1_1_1/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_1/Component_Function_2/NAND4_in[0] ), .A3(n6005), .A4(
        \SB1_1_1/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_1_1/buf_output[2] ) );
  NAND3_X2 U7906 ( .A1(\SB3_16/i0_4 ), .A2(\SB3_16/i0_3 ), .A3(\SB3_16/i1[9] ), 
        .ZN(n5848) );
  XOR2_X1 U7908 ( .A1(\SB2_2_2/buf_output[3] ), .A2(\RI5[2][33] ), .Z(n4047)
         );
  XOR2_X1 U7909 ( .A1(n5849), .A2(n34), .Z(Ciphertext[142]) );
  NAND4_X2 U7911 ( .A1(\SB4_8/Component_Function_4/NAND4_in[1] ), .A2(
        \SB4_8/Component_Function_4/NAND4_in[2] ), .A3(
        \SB4_8/Component_Function_4/NAND4_in[0] ), .A4(n2969), .ZN(n5849) );
  NAND4_X2 U7917 ( .A1(\SB1_1_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_30/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_5/NAND4_in[0] ), .A4(n5850), .ZN(
        \SB1_1_30/buf_output[5] ) );
  NAND3_X2 U7928 ( .A1(\SB1_1_30/i0[9] ), .A2(\SB1_1_30/i0[6] ), .A3(
        \SB1_1_30/i0_4 ), .ZN(n5850) );
  NAND3_X2 U7930 ( .A1(\SB2_2_9/i0[10] ), .A2(\SB2_2_9/i1[9] ), .A3(
        \SB2_2_9/i1_5 ), .ZN(n5851) );
  NAND3_X2 U7937 ( .A1(\SB1_0_4/i0_3 ), .A2(\SB1_0_4/i1[9] ), .A3(
        \SB1_0_4/i0_4 ), .ZN(\SB1_0_4/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U7941 ( .A1(\SB1_0_28/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_0_28/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[0][38] ) );
  NAND3_X2 U7942 ( .A1(\SB2_0_18/i0[10] ), .A2(\SB2_0_18/i0_3 ), .A3(
        \SB2_0_18/i0[9] ), .ZN(n6835) );
  NAND4_X2 U7943 ( .A1(\SB1_1_0/Component_Function_5/NAND4_in[3] ), .A2(n6975), 
        .A3(n6522), .A4(\SB1_1_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_0/buf_output[5] ) );
  NAND4_X2 U7948 ( .A1(\SB1_0_3/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_0_3/Component_Function_2/NAND4_in[2] ), .A3(n5890), .A4(n7447), 
        .ZN(\RI3[0][188] ) );
  NAND2_X2 U7949 ( .A1(n3044), .A2(n4892), .ZN(\SB2_3_29/i0_4 ) );
  XOR2_X1 U7951 ( .A1(n6932), .A2(n3840), .Z(\MC_ARK_ARC_1_3/buf_output[27] )
         );
  XOR2_X1 U7953 ( .A1(\MC_ARK_ARC_1_3/temp1[27] ), .A2(
        \MC_ARK_ARC_1_3/temp3[27] ), .Z(n6932) );
  NAND4_X2 U7958 ( .A1(n3080), .A2(n6125), .A3(n6124), .A4(
        \SB2_1_30/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_30/buf_output[5] ) );
  NAND3_X2 U7961 ( .A1(\SB3_11/i0[9] ), .A2(\SB3_11/i0_3 ), .A3(\SB3_11/i0[8] ), .ZN(\SB3_11/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U7971 ( .A1(\SB4_8/Component_Function_3/NAND4_in[3] ), .A2(n2195), 
        .A3(\SB4_8/Component_Function_3/NAND4_in[1] ), .A4(
        \SB4_8/Component_Function_3/NAND4_in[0] ), .ZN(n6100) );
  XOR2_X1 U7972 ( .A1(n6735), .A2(n5852), .Z(n1263) );
  XOR2_X1 U7976 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[7] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[1] ), .Z(n5852) );
  NAND3_X1 U7979 ( .A1(\SB2_0_30/i0[8] ), .A2(\SB2_0_30/i1_7 ), .A3(
        \RI3[0][10] ), .ZN(\SB2_0_30/Component_Function_1/NAND4_in[3] ) );
  INV_X2 U7980 ( .I(\SB1_4_27/buf_output[3] ), .ZN(\SB2_4_25/i0[8] ) );
  NAND4_X2 U7981 ( .A1(\SB1_4_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_27/Component_Function_3/NAND4_in[2] ), .A3(n6800), .A4(
        \SB1_4_27/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB1_4_27/buf_output[3] ) );
  XOR2_X1 U7982 ( .A1(n6558), .A2(\MC_ARK_ARC_1_4/temp1[96] ), .Z(
        \MC_ARK_ARC_1_4/temp5[96] ) );
  XOR2_X1 U7991 ( .A1(n4606), .A2(n5853), .Z(\MC_ARK_ARC_1_0/buf_output[22] )
         );
  XOR2_X1 U7993 ( .A1(\MC_ARK_ARC_1_0/temp2[22] ), .A2(
        \MC_ARK_ARC_1_0/temp1[22] ), .Z(n5853) );
  XOR2_X1 U7995 ( .A1(\RI5[0][86] ), .A2(\RI5[0][122] ), .Z(n5854) );
  NAND3_X2 U8000 ( .A1(\SB2_0_20/i0_0 ), .A2(\SB2_0_20/i1_5 ), .A3(
        \SB1_0_21/buf_output[4] ), .ZN(
        \SB2_0_20/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 U8001 ( .A1(\SB2_0_6/i1[9] ), .A2(\SB2_0_6/i1_5 ), .ZN(n5857) );
  NAND4_X2 U8002 ( .A1(n1568), .A2(\SB2_0_30/Component_Function_0/NAND4_in[1] ), .A3(\SB2_0_30/Component_Function_0/NAND4_in[0] ), .A4(n5858), .ZN(
        \SB2_0_30/buf_output[0] ) );
  NAND3_X2 U8003 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i0[8] ), .A3(\SB3_23/i0[9] ), .ZN(n5859) );
  XOR2_X1 U8004 ( .A1(n5860), .A2(n47), .Z(Ciphertext[117]) );
  NAND4_X2 U8006 ( .A1(n2791), .A2(\SB4_12/Component_Function_3/NAND4_in[0] ), 
        .A3(n1255), .A4(\SB4_12/Component_Function_3/NAND4_in[1] ), .ZN(n5860)
         );
  NAND4_X2 U8010 ( .A1(\SB1_0_28/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_28/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_0_28/buf_output[1] ) );
  NAND4_X2 U8011 ( .A1(n1863), .A2(\SB1_1_22/Component_Function_3/NAND4_in[0] ), .A3(\SB1_1_22/Component_Function_3/NAND4_in[2] ), .A4(n7492), .ZN(
        \SB1_1_22/buf_output[3] ) );
  NAND4_X2 U8013 ( .A1(\SB1_4_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_28/Component_Function_4/NAND4_in[1] ), .A3(n2238), .A4(
        \SB1_4_28/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_4_28/buf_output[4] ) );
  NAND3_X2 U8015 ( .A1(\SB2_4_27/i0_4 ), .A2(\SB2_4_27/i0_3 ), .A3(
        \SB2_4_27/i0_0 ), .ZN(n5861) );
  NAND3_X2 U8018 ( .A1(\SB2_3_14/i0_0 ), .A2(\SB2_3_14/i1_5 ), .A3(
        \SB2_3_14/i0_4 ), .ZN(n6078) );
  NAND4_X2 U8021 ( .A1(\SB2_1_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_19/Component_Function_0/NAND4_in[1] ), .A3(n5289), .A4(n5862), 
        .ZN(\SB2_1_19/buf_output[0] ) );
  XOR2_X1 U8022 ( .A1(n5863), .A2(n78), .Z(Ciphertext[121]) );
  NAND4_X2 U8023 ( .A1(\SB4_11/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_11/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_11/Component_Function_1/NAND4_in[3] ), .A4(
        \SB4_11/Component_Function_1/NAND4_in[0] ), .ZN(n5863) );
  NAND3_X1 U8026 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i0_0 ), .A3(
        \SB2_0_28/i0[7] ), .ZN(\SB2_0_28/Component_Function_0/NAND4_in[3] ) );
  NOR2_X2 U8028 ( .A1(n5865), .A2(n5864), .ZN(n3996) );
  XOR2_X1 U8029 ( .A1(\RI5[0][12] ), .A2(\RI5[0][96] ), .Z(n5866) );
  NAND3_X1 U8030 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i0[10] ), .A3(
        \SB2_0_28/i0_4 ), .ZN(\SB2_0_28/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U8031 ( .A1(\MC_ARK_ARC_1_3/temp4[10] ), .A2(n5867), .Z(n7152) );
  XOR2_X1 U8032 ( .A1(\RI5[3][112] ), .A2(\RI5[3][76] ), .Z(n5867) );
  NAND3_X2 U8034 ( .A1(\SB1_2_24/i0[8] ), .A2(\SB1_2_24/i3[0] ), .A3(
        \SB1_2_24/i1_5 ), .ZN(n6475) );
  NAND4_X2 U8035 ( .A1(n1353), .A2(n1637), .A3(n4951), .A4(n5868), .ZN(
        \SB1_2_24/buf_output[2] ) );
  NAND3_X2 U8036 ( .A1(\SB1_2_24/i0_4 ), .A2(\SB1_2_24/i0_0 ), .A3(
        \SB1_2_24/i1_5 ), .ZN(n5868) );
  XOR2_X1 U8037 ( .A1(n5870), .A2(n5869), .Z(\MC_ARK_ARC_1_2/temp6[110] ) );
  XOR2_X1 U8043 ( .A1(\RI5[2][20] ), .A2(n413), .Z(n5869) );
  XOR2_X1 U8046 ( .A1(\RI5[2][176] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .Z(n5870) );
  XOR2_X1 U8048 ( .A1(n5872), .A2(n5871), .Z(\MC_ARK_ARC_1_1/buf_output[121] )
         );
  XOR2_X1 U8049 ( .A1(\MC_ARK_ARC_1_1/temp4[121] ), .A2(n6335), .Z(n5871) );
  NAND4_X2 U8052 ( .A1(\SB2_1_28/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_28/Component_Function_5/NAND4_in[1] ), .A3(n3684), .A4(
        \SB2_1_28/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_28/buf_output[5] ) );
  NAND4_X2 U8053 ( .A1(\SB1_2_8/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_8/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_8/Component_Function_0/NAND4_in[3] ), .A4(n5873), .ZN(
        \SB1_2_8/buf_output[0] ) );
  XOR2_X1 U8055 ( .A1(n5874), .A2(n172), .Z(Ciphertext[183]) );
  NAND4_X2 U8057 ( .A1(n7172), .A2(\SB4_1/Component_Function_3/NAND4_in[3] ), 
        .A3(n5065), .A4(\SB4_1/Component_Function_3/NAND4_in[0] ), .ZN(n5874)
         );
  NAND3_X2 U8061 ( .A1(\SB1_2_24/i1_7 ), .A2(\SB1_2_24/i0[8] ), .A3(
        \SB1_2_24/i0_4 ), .ZN(\SB1_2_24/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U8063 ( .A1(n5875), .A2(n3), .Z(Ciphertext[134]) );
  NAND4_X2 U8064 ( .A1(\SB4_9/Component_Function_2/NAND4_in[0] ), .A2(n5924), 
        .A3(n5025), .A4(n1447), .ZN(n5875) );
  BUF_X4 U8068 ( .I(\SB2_4_8/buf_output[3] ), .Z(\RI5[4][153] ) );
  XOR2_X1 U8076 ( .A1(n5876), .A2(n191), .Z(Ciphertext[82]) );
  NAND4_X2 U8084 ( .A1(\SB4_18/Component_Function_4/NAND4_in[3] ), .A2(n7416), 
        .A3(n7343), .A4(\SB4_18/Component_Function_4/NAND4_in[1] ), .ZN(n5876)
         );
  NAND4_X2 U8085 ( .A1(n1781), .A2(\SB3_12/Component_Function_4/NAND4_in[1] ), 
        .A3(\SB3_12/Component_Function_4/NAND4_in[0] ), .A4(n5877), .ZN(
        \SB3_12/buf_output[4] ) );
  NAND3_X1 U8086 ( .A1(\SB3_12/i0[10] ), .A2(\SB3_12/i0[9] ), .A3(
        \RI1[5][119] ), .ZN(n5877) );
  NAND3_X1 U8088 ( .A1(\SB1_4_8/i0_0 ), .A2(\SB1_4_8/i3[0] ), .A3(
        \SB1_4_8/i1_7 ), .ZN(\SB1_4_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U8091 ( .A1(\SB1_4_17/i0[9] ), .A2(\SB1_4_17/i0[8] ), .A3(
        \SB1_4_17/i0_3 ), .ZN(n7375) );
  XOR2_X1 U8095 ( .A1(n5878), .A2(n188), .Z(Ciphertext[190]) );
  NAND4_X2 U8096 ( .A1(\SB4_0/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_0/Component_Function_4/NAND4_in[0] ), .A3(n2707), .A4(n1801), 
        .ZN(n5878) );
  NAND3_X2 U8097 ( .A1(\SB1_4_6/i0[9] ), .A2(\SB1_4_6/i0_4 ), .A3(
        \SB1_4_6/i0[6] ), .ZN(\SB1_4_6/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U8099 ( .A1(\SB1_2_13/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_13/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_13/Component_Function_2/NAND4_in[2] ), .A4(n5879), .ZN(
        \SB1_2_13/buf_output[2] ) );
  NAND3_X1 U8101 ( .A1(\SB1_2_13/i0_0 ), .A2(\SB1_2_13/i1_5 ), .A3(
        \MC_ARK_ARC_1_1/buf_output[112] ), .ZN(n5879) );
  XOR2_X1 U8105 ( .A1(\RI5[4][161] ), .A2(\RI5[4][5] ), .Z(n7519) );
  XOR2_X1 U8112 ( .A1(\RI5[4][11] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[167] ), 
        .Z(n5880) );
  NAND3_X1 U8115 ( .A1(\SB1_2_19/i0[10] ), .A2(\SB1_2_19/i0_3 ), .A3(
        \SB1_2_19/i0[9] ), .ZN(n2369) );
  NAND3_X1 U8120 ( .A1(\SB1_4_6/buf_output[4] ), .A2(\SB2_4_5/i0[9] ), .A3(
        \SB2_4_5/i0[6] ), .ZN(n3002) );
  XOR2_X1 U8121 ( .A1(n5881), .A2(n40), .Z(Ciphertext[136]) );
  NAND4_X2 U8122 ( .A1(\SB4_9/Component_Function_4/NAND4_in[3] ), .A2(n2107), 
        .A3(n2941), .A4(n1068), .ZN(n5881) );
  XOR2_X1 U8127 ( .A1(n5882), .A2(n207), .Z(Ciphertext[152]) );
  NAND4_X2 U8128 ( .A1(\SB4_6/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_6/Component_Function_2/NAND4_in[0] ), .A3(
        \SB4_6/Component_Function_2/NAND4_in[3] ), .A4(n6017), .ZN(n5882) );
  BUF_X4 U8129 ( .I(\SB2_0_18/buf_output[1] ), .Z(\RI5[0][103] ) );
  NAND4_X2 U8130 ( .A1(\SB1_4_30/Component_Function_2/NAND4_in[0] ), .A2(n1344), .A3(n3562), .A4(n6789), .ZN(\SB1_4_30/buf_output[2] ) );
  NAND4_X2 U8131 ( .A1(\SB1_0_18/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_18/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_18/Component_Function_5/NAND4_in[0] ), .A4(n901), .ZN(
        \RI3[0][83] ) );
  NAND4_X2 U8132 ( .A1(n671), .A2(\SB1_2_17/Component_Function_5/NAND4_in[3] ), 
        .A3(n5905), .A4(\SB1_2_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_17/buf_output[5] ) );
  NAND3_X2 U8133 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0_4 ), .A3(
        \SB1_1_20/i1[9] ), .ZN(\SB1_1_20/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U8134 ( .A1(\SB1_1_14/i0[6] ), .A2(\SB1_1_14/i0_4 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[102] ), .ZN(n2723) );
  XOR2_X1 U8136 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[71] ), .A2(\RI5[1][95] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[125] ) );
  NAND3_X2 U8141 ( .A1(\SB2_4_27/i0_3 ), .A2(\SB2_4_27/i1[9] ), .A3(
        \SB2_4_27/i0_4 ), .ZN(n2894) );
  NAND4_X2 U8148 ( .A1(\SB2_0_1/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_1/Component_Function_0/NAND4_in[3] ), .A3(n7192), .A4(
        \SB2_0_1/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_1/buf_output[0] ) );
  XOR2_X1 U8160 ( .A1(\MC_ARK_ARC_1_1/temp2[58] ), .A2(n5884), .Z(
        \MC_ARK_ARC_1_1/temp5[58] ) );
  NAND4_X2 U8163 ( .A1(\SB2_0_16/Component_Function_2/NAND4_in[0] ), .A2(n5071), .A3(n6405), .A4(n5885), .ZN(\SB2_0_16/buf_output[2] ) );
  NAND3_X2 U8166 ( .A1(\SB2_0_16/i0_0 ), .A2(n594), .A3(\SB2_0_16/i1_5 ), .ZN(
        n5885) );
  NAND3_X2 U8167 ( .A1(\SB1_3_27/i0_3 ), .A2(\SB1_3_27/i0_0 ), .A3(
        \SB1_3_27/i0_4 ), .ZN(n5886) );
  XOR2_X1 U8170 ( .A1(n3457), .A2(n5887), .Z(n3326) );
  XOR2_X1 U8175 ( .A1(\RI5[1][92] ), .A2(\RI5[1][158] ), .Z(n5887) );
  NAND3_X2 U8176 ( .A1(\SB2_2_22/i1[9] ), .A2(\SB2_2_22/i0_3 ), .A3(
        \SB2_2_22/i0[6] ), .ZN(\SB2_2_22/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U8177 ( .A1(\RI5[1][26] ), .A2(\SB2_1_29/buf_output[2] ), .Z(n5954)
         );
  NAND3_X1 U8179 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i0[8] ), .A3(\SB4_2/i0[9] ), 
        .ZN(n5888) );
  NAND4_X2 U8183 ( .A1(\SB1_1_4/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_4/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_4/Component_Function_1/NAND4_in[0] ), .A4(n5889), .ZN(
        \SB1_1_4/buf_output[1] ) );
  NAND3_X2 U8185 ( .A1(\SB1_1_4/i0_4 ), .A2(\SB1_1_4/i0[8] ), .A3(
        \SB1_1_4/i1_7 ), .ZN(n5889) );
  NAND4_X2 U8188 ( .A1(n6044), .A2(\SB2_3_3/Component_Function_0/NAND4_in[1] ), 
        .A3(\SB2_3_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_3/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_3/buf_output[0] ) );
  NAND3_X2 U8192 ( .A1(\SB1_0_3/i0[10] ), .A2(\SB1_0_3/i1[9] ), .A3(
        \SB1_0_3/i1_5 ), .ZN(n5890) );
  NAND3_X2 U8195 ( .A1(\SB1_2_17/i0_4 ), .A2(\SB1_2_17/i0[9] ), .A3(
        \SB1_2_17/i0[6] ), .ZN(\SB1_2_17/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U8199 ( .A1(\MC_ARK_ARC_1_1/temp4[88] ), .A2(n5891), .Z(
        \MC_ARK_ARC_1_1/temp6[88] ) );
  XOR2_X1 U8203 ( .A1(\SB2_1_1/buf_output[4] ), .A2(\RI5[1][154] ), .Z(n5891)
         );
  NAND4_X2 U8204 ( .A1(\SB1_2_8/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_8/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_2_8/Component_Function_5/NAND4_in[0] ), .A4(n5892), .ZN(
        \SB1_2_8/buf_output[5] ) );
  NAND3_X2 U8205 ( .A1(\SB1_2_8/i0[9] ), .A2(\SB1_2_8/i0_4 ), .A3(
        \SB1_2_8/i0[6] ), .ZN(n5892) );
  XOR2_X1 U8206 ( .A1(n5893), .A2(n103), .Z(Ciphertext[178]) );
  NAND4_X2 U8207 ( .A1(n6918), .A2(\SB4_2/Component_Function_4/NAND4_in[3] ), 
        .A3(\SB4_2/Component_Function_4/NAND4_in[0] ), .A4(n2898), .ZN(n5893)
         );
  XOR2_X1 U8208 ( .A1(\MC_ARK_ARC_1_2/temp2[62] ), .A2(
        \MC_ARK_ARC_1_2/temp1[62] ), .Z(n5894) );
  XOR2_X1 U8214 ( .A1(n3009), .A2(n5105), .Z(\MC_ARK_ARC_1_1/buf_output[147] )
         );
  XOR2_X1 U8215 ( .A1(n5380), .A2(n4820), .Z(n3009) );
  NAND4_X2 U8227 ( .A1(n7227), .A2(\SB2_3_1/Component_Function_4/NAND4_in[0] ), 
        .A3(\SB2_3_1/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_1/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_3_1/buf_output[4] ) );
  NAND4_X2 U8228 ( .A1(\SB1_3_8/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_8/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_8/Component_Function_2/NAND4_in[2] ), .A4(n5895), .ZN(
        \SB1_3_8/buf_output[2] ) );
  NAND3_X2 U8236 ( .A1(\SB1_3_8/i0_0 ), .A2(\SB1_3_8/i1_5 ), .A3(
        \SB1_3_8/i0_4 ), .ZN(n5895) );
  INV_X2 U8237 ( .I(\SB1_4_29/buf_output[2] ), .ZN(\SB2_4_26/i1[9] ) );
  NAND4_X2 U8238 ( .A1(\SB1_4_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_4_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_4_29/Component_Function_2/NAND4_in[3] ), .A4(n4156), .ZN(
        \SB1_4_29/buf_output[2] ) );
  NAND3_X2 U8240 ( .A1(\SB2_0_21/i0_0 ), .A2(\SB2_0_21/i1_5 ), .A3(
        \SB2_0_21/i0_4 ), .ZN(n7433) );
  XOR2_X1 U8242 ( .A1(\RI5[1][101] ), .A2(\RI5[1][95] ), .Z(n5896) );
  XOR2_X1 U8243 ( .A1(\RI5[3][174] ), .A2(\SB2_3_3/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/temp2[36] ) );
  NAND4_X2 U8247 ( .A1(\SB1_3_18/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_18/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_3_18/Component_Function_2/NAND4_in[0] ), .A4(n5897), .ZN(
        \SB1_3_18/buf_output[2] ) );
  NAND3_X2 U8250 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i1_5 ), .A3(
        \SB1_3_18/i0_4 ), .ZN(n5897) );
  XOR2_X1 U8252 ( .A1(n7266), .A2(n5898), .Z(\MC_ARK_ARC_1_0/temp5[64] ) );
  NAND3_X2 U8260 ( .A1(n6686), .A2(\SB1_2_31/buf_output[0] ), .A3(
        \SB2_2_26/i0[6] ), .ZN(n6614) );
  NAND4_X2 U8263 ( .A1(\SB2_4_5/Component_Function_3/NAND4_in[2] ), .A2(n1937), 
        .A3(n7384), .A4(n5899), .ZN(\SB2_4_5/buf_output[3] ) );
  NAND3_X2 U8264 ( .A1(\SB2_4_5/i0_3 ), .A2(\SB2_4_5/i0[6] ), .A3(
        \SB2_4_5/i1[9] ), .ZN(n5899) );
  NAND4_X2 U8277 ( .A1(\SB2_3_8/Component_Function_2/NAND4_in[0] ), .A2(n1371), 
        .A3(\SB2_3_8/Component_Function_2/NAND4_in[2] ), .A4(n6562), .ZN(
        \SB2_3_8/buf_output[2] ) );
  NAND3_X2 U8279 ( .A1(\SB1_1_9/i0[10] ), .A2(\SB1_1_9/i1[9] ), .A3(
        \SB1_1_9/i1_7 ), .ZN(\SB1_1_9/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U8280 ( .A1(\MC_ARK_ARC_1_1/temp5[83] ), .A2(n5900), .Z(
        \MC_ARK_ARC_1_1/buf_output[83] ) );
  XOR2_X1 U8282 ( .A1(n3389), .A2(n3390), .Z(n5900) );
  XOR2_X1 U8285 ( .A1(n5902), .A2(n5901), .Z(\MC_ARK_ARC_1_1/temp5[62] ) );
  XOR2_X1 U8287 ( .A1(\RI5[1][56] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .Z(n5901) );
  XOR2_X1 U8292 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[32] ), .A2(n3167), .Z(
        n5902) );
  XOR2_X1 U8294 ( .A1(n5904), .A2(n5903), .Z(n4495) );
  XOR2_X1 U8305 ( .A1(\RI5[1][104] ), .A2(n71), .Z(n5903) );
  XOR2_X1 U8307 ( .A1(\RI5[1][170] ), .A2(\RI5[1][80] ), .Z(n5904) );
  NAND4_X2 U8309 ( .A1(n2435), .A2(\SB2_1_6/Component_Function_5/NAND4_in[0] ), 
        .A3(\SB2_1_6/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_6/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_1_6/buf_output[5] ) );
  NAND3_X2 U8311 ( .A1(\SB1_2_17/i0_0 ), .A2(\SB1_2_17/i0[6] ), .A3(
        \SB1_2_17/i0[10] ), .ZN(n5905) );
  NAND4_X2 U8314 ( .A1(\SB1_0_15/Component_Function_2/NAND4_in[0] ), .A2(n4049), .A3(\SB1_0_15/Component_Function_2/NAND4_in[2] ), .A4(n5906), .ZN(
        \RI3[0][116] ) );
  NAND3_X2 U8315 ( .A1(\SB1_0_15/i0_4 ), .A2(\SB1_0_15/i1_5 ), .A3(
        \SB1_0_15/i0_0 ), .ZN(n5906) );
  NAND4_X2 U8316 ( .A1(\SB1_3_6/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_3_6/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_3_6/Component_Function_0/NAND4_in[0] ), .A4(n3662), .ZN(
        \SB1_3_6/buf_output[0] ) );
  XOR2_X1 U8319 ( .A1(n5908), .A2(n5907), .Z(\MC_ARK_ARC_1_2/buf_output[98] )
         );
  XOR2_X1 U8322 ( .A1(\MC_ARK_ARC_1_2/temp3[98] ), .A2(
        \MC_ARK_ARC_1_2/temp2[98] ), .Z(n5908) );
  XOR2_X1 U8323 ( .A1(n5909), .A2(\MC_ARK_ARC_1_3/temp4[19] ), .Z(
        \MC_ARK_ARC_1_3/temp6[19] ) );
  XOR2_X1 U8330 ( .A1(\MC_ARK_ARC_1_1/temp2[110] ), .A2(
        \MC_ARK_ARC_1_1/temp1[110] ), .Z(n4665) );
  NAND3_X2 U8332 ( .A1(\SB2_0_21/i1[9] ), .A2(\SB2_0_21/i0_3 ), .A3(
        \SB2_0_21/i0_4 ), .ZN(\SB2_0_21/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U8335 ( .I(\SB3_9/buf_output[5] ), .Z(\SB4_9/i0_3 ) );
  XOR2_X1 U8341 ( .A1(n1576), .A2(\MC_ARK_ARC_1_0/temp6[24] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[24] ) );
  XOR2_X1 U8344 ( .A1(\RI5[0][90] ), .A2(\RI5[0][126] ), .Z(
        \MC_ARK_ARC_1_0/temp3[24] ) );
  NAND3_X2 U8346 ( .A1(n6585), .A2(n6379), .A3(
        \SB1_1_27/Component_Function_5/NAND4_in[1] ), .ZN(
        \SB1_1_27/buf_output[5] ) );
  XOR2_X1 U8350 ( .A1(n3683), .A2(n5910), .Z(\MC_ARK_ARC_1_1/buf_output[113] )
         );
  XOR2_X1 U8351 ( .A1(n4235), .A2(\MC_ARK_ARC_1_1/temp4[113] ), .Z(n5910) );
  NAND4_X2 U8354 ( .A1(\SB4_6/Component_Function_3/NAND4_in[2] ), .A2(
        \SB4_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_6/Component_Function_3/NAND4_in[3] ), .A4(n5911), .ZN(n6939) );
  NAND3_X2 U8356 ( .A1(\SB4_6/i0[6] ), .A2(\SB4_6/i0_3 ), .A3(\SB4_6/i1[9] ), 
        .ZN(n5911) );
  NAND3_X2 U8364 ( .A1(\SB3_9/i0[6] ), .A2(\SB3_9/i0[10] ), .A3(\SB3_9/i0_3 ), 
        .ZN(n5912) );
  NAND4_X2 U8372 ( .A1(\SB4_9/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_9/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_9/Component_Function_0/NAND4_in[1] ), .A4(n2308), .ZN(n6742) );
  NAND3_X1 U8373 ( .A1(n1498), .A2(\SB4_13/i3[0] ), .A3(n4002), .ZN(
        \SB4_13/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U8374 ( .A1(\SB3_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_4/NAND4_in[2] ), .A3(n2215), .A4(n5913), 
        .ZN(\SB3_11/buf_output[4] ) );
  NAND3_X1 U8378 ( .A1(\SB3_11/i0_0 ), .A2(\SB3_11/i1_7 ), .A3(\SB3_11/i3[0] ), 
        .ZN(n5913) );
  XOR2_X1 U8379 ( .A1(\MC_ARK_ARC_1_3/temp1[158] ), .A2(n5914), .Z(
        \MC_ARK_ARC_1_3/temp5[158] ) );
  XOR2_X1 U8385 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[128] ), .A2(\RI5[3][104] ), 
        .Z(n5914) );
  XOR2_X1 U8387 ( .A1(n7463), .A2(n5915), .Z(\MC_ARK_ARC_1_1/buf_output[179] )
         );
  XOR2_X1 U8390 ( .A1(n5916), .A2(n215), .Z(Ciphertext[43]) );
  NAND4_X2 U8393 ( .A1(\SB4_24/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_24/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_24/Component_Function_1/NAND4_in[2] ), .ZN(n5916) );
  XOR2_X1 U8394 ( .A1(\MC_ARK_ARC_1_3/temp4[62] ), .A2(n5917), .Z(n5947) );
  XOR2_X1 U8396 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[128] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[164] ), .Z(n5917) );
  XOR2_X1 U8398 ( .A1(n5918), .A2(n114), .Z(Ciphertext[32]) );
  NAND4_X2 U8401 ( .A1(n5421), .A2(\SB4_26/Component_Function_2/NAND4_in[0] ), 
        .A3(n967), .A4(n5168), .ZN(n5918) );
  NAND3_X1 U8403 ( .A1(\SB2_4_20/i0_4 ), .A2(\SB2_4_20/i1[9] ), .A3(
        \SB2_4_20/i1_5 ), .ZN(\SB2_4_20/Component_Function_4/NAND4_in[3] ) );
  NAND2_X2 U8406 ( .A1(n5104), .A2(n6724), .ZN(\SB2_4_20/i0_4 ) );
  XOR2_X1 U8407 ( .A1(n5919), .A2(n59), .Z(Ciphertext[158]) );
  NAND4_X2 U8412 ( .A1(n3398), .A2(n3541), .A3(n7029), .A4(
        \SB4_5/Component_Function_2/NAND4_in[2] ), .ZN(n5919) );
  NAND3_X1 U8414 ( .A1(\SB4_25/i0_0 ), .A2(n6266), .A3(\SB4_25/i0[8] ), .ZN(
        \SB4_25/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U8416 ( .A1(\SB1_4_28/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_4_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_28/Component_Function_1/NAND4_in[0] ), .A4(n5920), .ZN(
        \SB1_4_28/buf_output[1] ) );
  NAND3_X1 U8417 ( .A1(\SB1_4_28/i0[6] ), .A2(\SB1_4_28/i1_5 ), .A3(
        \SB1_4_28/i0[9] ), .ZN(n5920) );
  NAND3_X2 U8418 ( .A1(\SB2_4_24/i0[10] ), .A2(\SB2_4_24/i1_7 ), .A3(n5443), 
        .ZN(n7257) );
  XOR2_X1 U8422 ( .A1(n6756), .A2(n5921), .Z(\MC_ARK_ARC_1_4/buf_output[147] )
         );
  XOR2_X1 U8436 ( .A1(n6076), .A2(\MC_ARK_ARC_1_4/temp4[147] ), .Z(n5921) );
  NAND3_X2 U8437 ( .A1(\SB2_4_26/i1_5 ), .A2(\SB2_4_26/i0[8] ), .A3(
        \SB2_4_26/i3[0] ), .ZN(\SB2_4_26/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U8438 ( .A1(n5922), .A2(n128), .Z(Ciphertext[94]) );
  NAND4_X2 U8439 ( .A1(\SB4_16/Component_Function_4/NAND4_in[1] ), .A2(n2923), 
        .A3(\SB4_16/Component_Function_4/NAND4_in[0] ), .A4(n6484), .ZN(n5922)
         );
  NAND4_X2 U8441 ( .A1(n2902), .A2(\SB1_2_15/Component_Function_4/NAND4_in[0] ), .A3(n1821), .A4(n5923), .ZN(\SB1_2_15/buf_output[4] ) );
  NAND3_X1 U8443 ( .A1(\SB1_2_15/i0_0 ), .A2(\SB1_2_15/i3[0] ), .A3(
        \SB1_2_15/i1_7 ), .ZN(n5923) );
  NAND3_X1 U8445 ( .A1(\SB4_9/i0_0 ), .A2(n6272), .A3(\SB4_9/i1_5 ), .ZN(n5924) );
  NAND2_X2 U8448 ( .A1(n1303), .A2(n5925), .ZN(\RI5[4][109] ) );
  AND2_X1 U8450 ( .A1(\SB2_4_17/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_4_17/Component_Function_1/NAND4_in[0] ), .Z(n5925) );
  NAND4_X2 U8452 ( .A1(n3922), .A2(\SB2_4_12/Component_Function_2/NAND4_in[2] ), .A3(\SB2_4_12/Component_Function_2/NAND4_in[0] ), .A4(n5926), .ZN(
        \SB2_4_12/buf_output[2] ) );
  NAND3_X2 U8461 ( .A1(\SB2_4_12/i0[6] ), .A2(\SB2_4_12/i0_3 ), .A3(
        \SB2_4_12/i0[10] ), .ZN(n5926) );
  NAND4_X2 U8463 ( .A1(\SB1_3_17/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_17/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_3_17/Component_Function_4/NAND4_in[2] ), .A4(n5927), .ZN(
        \SB1_3_17/buf_output[4] ) );
  XOR2_X1 U8466 ( .A1(\MC_ARK_ARC_1_4/temp2[134] ), .A2(n5928), .Z(n7296) );
  XOR2_X1 U8467 ( .A1(\RI5[4][134] ), .A2(\RI5[4][128] ), .Z(n5928) );
  INV_X2 U8472 ( .I(\SB1_4_19/buf_output[3] ), .ZN(\SB2_4_17/i0[8] ) );
  NAND4_X2 U8473 ( .A1(\SB1_4_19/Component_Function_3/NAND4_in[0] ), .A2(n2039), .A3(n934), .A4(n1035), .ZN(\SB1_4_19/buf_output[3] ) );
  XOR2_X1 U8474 ( .A1(n5929), .A2(n154), .Z(Ciphertext[128]) );
  NAND4_X2 U8478 ( .A1(n3932), .A2(n5369), .A3(n3477), .A4(n6747), .ZN(n5929)
         );
  NAND3_X2 U8484 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i1[9] ), .A3(n5433), 
        .ZN(\SB1_0_28/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U8486 ( .A1(\SB1_1_9/Component_Function_5/NAND4_in[2] ), .A2(n1878), 
        .A3(\SB1_1_9/Component_Function_5/NAND4_in[0] ), .A4(n5930), .ZN(
        \SB1_1_9/buf_output[5] ) );
  NAND3_X2 U8490 ( .A1(\SB1_1_9/i0[6] ), .A2(\SB1_1_9/i0_4 ), .A3(
        \SB1_1_9/i0[9] ), .ZN(n5930) );
  XOR2_X1 U8493 ( .A1(\RI5[1][123] ), .A2(\RI5[1][93] ), .Z(n4036) );
  NAND4_X2 U8498 ( .A1(\SB1_1_4/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_4/Component_Function_2/NAND4_in[2] ), .A3(n6067), .A4(n5931), 
        .ZN(\SB1_1_4/buf_output[2] ) );
  NAND3_X2 U8501 ( .A1(\SB1_1_4/i0_4 ), .A2(\SB1_1_4/i0_0 ), .A3(
        \SB1_1_4/i1_5 ), .ZN(n5931) );
  NOR2_X2 U8504 ( .A1(n2599), .A2(n5932), .ZN(\SB2_3_4/i0[7] ) );
  XOR2_X1 U8505 ( .A1(\MC_ARK_ARC_1_2/temp2[159] ), .A2(n5933), .Z(
        \MC_ARK_ARC_1_2/temp5[159] ) );
  XOR2_X1 U8506 ( .A1(\RI5[2][159] ), .A2(\RI5[2][153] ), .Z(n5933) );
  XOR2_X1 U8508 ( .A1(\RI5[1][190] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[34] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[124] ) );
  XOR2_X1 U8509 ( .A1(\MC_ARK_ARC_1_1/temp6[124] ), .A2(n817), .Z(
        \MC_ARK_ARC_1_1/buf_output[124] ) );
  XOR2_X1 U8510 ( .A1(n7292), .A2(n5934), .Z(\MC_ARK_ARC_1_0/buf_output[41] )
         );
  XOR2_X1 U8514 ( .A1(\MC_ARK_ARC_1_0/temp3[41] ), .A2(
        \MC_ARK_ARC_1_0/temp1[41] ), .Z(n5934) );
  XOR2_X1 U8532 ( .A1(\MC_ARK_ARC_1_0/temp4[7] ), .A2(
        \MC_ARK_ARC_1_0/temp3[7] ), .Z(\MC_ARK_ARC_1_0/temp6[7] ) );
  XOR2_X1 U8535 ( .A1(\MC_ARK_ARC_1_0/temp3[172] ), .A2(
        \MC_ARK_ARC_1_0/temp2[172] ), .Z(n1641) );
  NAND4_X2 U8536 ( .A1(\SB1_2_23/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_0/NAND4_in[0] ), .A4(n5935), .ZN(
        \SB1_2_23/buf_output[0] ) );
  NAND2_X1 U8537 ( .A1(\SB4_12/i0[9] ), .A2(\SB4_12/i0[10] ), .ZN(n5936) );
  NAND3_X2 U8538 ( .A1(\SB1_1_14/i0[10] ), .A2(\SB1_1_14/i0_0 ), .A3(
        \SB1_1_14/i0[6] ), .ZN(n4786) );
  NAND3_X2 U8540 ( .A1(\SB2_0_17/i0_0 ), .A2(\SB2_0_17/i0_3 ), .A3(
        \RI3[0][88] ), .ZN(n7247) );
  NAND3_X2 U8541 ( .A1(\SB3_17/i0_3 ), .A2(\SB3_17/i0[7] ), .A3(\SB3_17/i0_0 ), 
        .ZN(n3782) );
  NAND3_X2 U8542 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0_4 ), .A3(\SB4_16/i0_3 ), 
        .ZN(n6912) );
  NAND4_X2 U8544 ( .A1(\SB2_3_10/Component_Function_2/NAND4_in[0] ), .A2(n7418), .A3(n3373), .A4(\SB2_3_10/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_3_10/buf_output[2] ) );
  XOR2_X1 U8550 ( .A1(\RI5[4][83] ), .A2(\RI5[4][89] ), .Z(n7103) );
  NAND3_X2 U8551 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0_4 ), .A3(
        \SB2_1_9/i1[9] ), .ZN(n2821) );
  XOR2_X1 U8552 ( .A1(\RI5[3][174] ), .A2(\RI5[3][168] ), .Z(
        \MC_ARK_ARC_1_3/temp1[174] ) );
  XOR2_X1 U8553 ( .A1(\RI5[2][158] ), .A2(\RI5[2][134] ), .Z(n3381) );
  XOR2_X1 U8563 ( .A1(n7451), .A2(n5937), .Z(\MC_ARK_ARC_1_1/buf_output[59] )
         );
  XOR2_X1 U8564 ( .A1(\MC_ARK_ARC_1_1/temp4[59] ), .A2(n4569), .Z(n5937) );
  XOR2_X1 U8567 ( .A1(\RI5[0][99] ), .A2(\RI5[0][105] ), .Z(
        \MC_ARK_ARC_1_0/temp1[105] ) );
  XOR2_X1 U8572 ( .A1(n5939), .A2(n5938), .Z(\MC_ARK_ARC_1_1/buf_output[167] )
         );
  XOR2_X1 U8575 ( .A1(n3543), .A2(n6439), .Z(n5938) );
  XOR2_X1 U8579 ( .A1(n3544), .A2(n3337), .Z(n5939) );
  NAND3_X2 U8586 ( .A1(\SB1_2_15/i0_0 ), .A2(\SB1_2_15/i0[10] ), .A3(
        \SB1_2_15/i0[6] ), .ZN(n5940) );
  NAND4_X2 U8591 ( .A1(\SB2_4_2/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_4_2/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_4_2/Component_Function_4/NAND4_in[3] ), .A4(n5941), .ZN(
        \SB2_4_2/buf_output[4] ) );
  XOR2_X1 U8595 ( .A1(n5943), .A2(n5942), .Z(\MC_ARK_ARC_1_2/buf_output[21] )
         );
  XOR2_X1 U8597 ( .A1(\MC_ARK_ARC_1_2/temp1[21] ), .A2(
        \MC_ARK_ARC_1_2/temp4[21] ), .Z(n5942) );
  XOR2_X1 U8599 ( .A1(\MC_ARK_ARC_1_2/temp3[21] ), .A2(
        \MC_ARK_ARC_1_2/temp2[21] ), .Z(n5943) );
  NAND3_X2 U8601 ( .A1(\SB3_13/i0_3 ), .A2(\SB3_13/i0[10] ), .A3(
        \SB3_13/i0[9] ), .ZN(n5229) );
  NAND3_X2 U8603 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i0_3 ), .A3(\SB4_12/i0_4 ), 
        .ZN(\SB4_12/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U8604 ( .A1(\SB1_4_21/Component_Function_5/NAND4_in[1] ), .A2(n3110), .A3(n2463), .A4(n5944), .ZN(\SB1_4_21/buf_output[5] ) );
  NAND2_X1 U8606 ( .A1(\SB1_4_21/i0_0 ), .A2(\SB1_4_21/i3[0] ), .ZN(n5944) );
  XOR2_X1 U8615 ( .A1(n5945), .A2(n66), .Z(Ciphertext[51]) );
  NAND4_X2 U8616 ( .A1(\SB4_23/Component_Function_3/NAND4_in[3] ), .A2(n3350), 
        .A3(n2141), .A4(\SB4_23/Component_Function_3/NAND4_in[1] ), .ZN(n5945)
         );
  XOR2_X1 U8619 ( .A1(n5947), .A2(n5946), .Z(\MC_ARK_ARC_1_3/buf_output[62] )
         );
  XOR2_X1 U8623 ( .A1(\MC_ARK_ARC_1_3/temp1[62] ), .A2(
        \MC_ARK_ARC_1_3/temp2[62] ), .Z(n5946) );
  NAND3_X2 U8624 ( .A1(\SB3_11/i1[9] ), .A2(\SB3_11/i0[10] ), .A3(
        \SB3_11/i1_7 ), .ZN(\SB3_11/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U8625 ( .A1(\MC_ARK_ARC_1_3/temp3[147] ), .A2(n5948), .Z(n6519) );
  INV_X1 U8631 ( .I(\SB3_28/buf_output[0] ), .ZN(\SB4_23/i3[0] ) );
  NAND4_X2 U8632 ( .A1(\SB3_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_0/NAND4_in[0] ), .A4(
        \SB3_28/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_28/buf_output[0] ) );
  XOR2_X1 U8633 ( .A1(n5949), .A2(n24), .Z(Ciphertext[133]) );
  NAND4_X2 U8634 ( .A1(\SB4_9/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_9/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_9/Component_Function_1/NAND4_in[0] ), .ZN(n5949) );
  XOR2_X1 U8636 ( .A1(n5951), .A2(n5950), .Z(\RI1[5][77] ) );
  XOR2_X1 U8638 ( .A1(\MC_ARK_ARC_1_4/temp1[77] ), .A2(
        \MC_ARK_ARC_1_4/temp4[77] ), .Z(n5950) );
  XOR2_X1 U8639 ( .A1(\MC_ARK_ARC_1_4/temp2[77] ), .A2(
        \MC_ARK_ARC_1_4/temp3[77] ), .Z(n5951) );
  INV_X2 U8640 ( .I(\SB1_2_20/buf_output[3] ), .ZN(\SB2_2_18/i0[8] ) );
  NAND3_X2 U8642 ( .A1(\SB2_3_24/i0[6] ), .A2(\SB2_3_24/i0_4 ), .A3(
        \SB2_3_24/i0[9] ), .ZN(\SB2_3_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U8645 ( .A1(\SB1_2_10/i0[10] ), .A2(\SB1_2_10/i0[9] ), .A3(
        \SB1_2_10/i0_3 ), .ZN(\SB1_2_10/Component_Function_4/NAND4_in[2] ) );
  INV_X2 U8648 ( .I(\SB1_4_15/buf_output[2] ), .ZN(\SB2_4_12/i1[9] ) );
  NAND4_X2 U8649 ( .A1(n1545), .A2(\SB1_4_15/Component_Function_2/NAND4_in[1] ), .A3(n3920), .A4(n5400), .ZN(\SB1_4_15/buf_output[2] ) );
  XOR2_X1 U8652 ( .A1(n6896), .A2(n5952), .Z(n4480) );
  XOR2_X1 U8653 ( .A1(\RI5[0][176] ), .A2(\RI5[0][8] ), .Z(n5952) );
  NAND4_X2 U8655 ( .A1(\SB1_3_31/Component_Function_2/NAND4_in[2] ), .A2(n4924), .A3(\SB1_3_31/Component_Function_2/NAND4_in[3] ), .A4(n4329), .ZN(
        \SB1_3_31/buf_output[2] ) );
  NAND4_X2 U8657 ( .A1(\SB3_28/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_28/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_28/Component_Function_2/NAND4_in[1] ), .A4(
        \SB3_28/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_28/buf_output[2] ) );
  XOR2_X1 U8658 ( .A1(n5953), .A2(n62), .Z(Ciphertext[8]) );
  XOR2_X1 U8660 ( .A1(\MC_ARK_ARC_1_1/temp2[32] ), .A2(n5954), .Z(n4357) );
  NAND4_X2 U8662 ( .A1(\SB1_4_12/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_4_12/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_4_12/Component_Function_3/NAND4_in[3] ), .A4(n5955), .ZN(
        \SB1_4_12/buf_output[3] ) );
  NAND3_X2 U8665 ( .A1(\SB1_4_12/i0[10] ), .A2(\SB1_4_12/i1_7 ), .A3(
        \SB1_4_12/i1[9] ), .ZN(n5955) );
  INV_X4 U8666 ( .I(n6612), .ZN(\SB2_1_29/i0_4 ) );
  XOR2_X1 U8668 ( .A1(\MC_ARK_ARC_1_3/temp5[169] ), .A2(
        \MC_ARK_ARC_1_3/temp6[169] ), .Z(\MC_ARK_ARC_1_3/buf_output[169] ) );
  NAND2_X1 U8671 ( .A1(n2311), .A2(n6880), .ZN(n7277) );
  NAND4_X2 U8672 ( .A1(\SB1_4_1/Component_Function_4/NAND4_in[0] ), .A2(n6094), 
        .A3(\SB1_4_1/Component_Function_4/NAND4_in[1] ), .A4(n5956), .ZN(
        \SB1_4_1/buf_output[4] ) );
  NAND3_X2 U8673 ( .A1(\SB1_4_1/i0[10] ), .A2(\SB1_4_1/i0[9] ), .A3(
        \SB1_4_1/i0_3 ), .ZN(n5956) );
  XOR2_X1 U8678 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[35] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[71] ), .Z(\MC_ARK_ARC_1_0/temp3[161] )
         );
  NAND4_X2 U8679 ( .A1(\SB2_0_24/Component_Function_5/NAND4_in[3] ), .A2(n4169), .A3(n6144), .A4(n5957), .ZN(\SB2_0_24/buf_output[5] ) );
  NAND2_X2 U8680 ( .A1(\SB2_0_24/i0_0 ), .A2(\SB2_0_24/i3[0] ), .ZN(n5957) );
  NAND4_X2 U8681 ( .A1(\SB3_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_10/Component_Function_3/NAND4_in[3] ), .A3(
        \SB3_10/Component_Function_3/NAND4_in[2] ), .A4(n5958), .ZN(
        \SB3_10/buf_output[3] ) );
  NAND3_X1 U8682 ( .A1(\SB3_10/i0_3 ), .A2(\SB3_10/i0_4 ), .A3(\SB3_10/i0_0 ), 
        .ZN(n5958) );
  XOR2_X1 U8684 ( .A1(\RI5[4][101] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[77] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[131] ) );
  XOR2_X1 U8692 ( .A1(n642), .A2(n5960), .Z(n5034) );
  XOR2_X1 U8693 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[45] ), .A2(\RI5[4][21] ), 
        .Z(n5960) );
  XOR2_X1 U8707 ( .A1(\RI5[0][26] ), .A2(\RI5[0][32] ), .Z(
        \MC_ARK_ARC_1_0/temp1[32] ) );
  XOR2_X1 U8710 ( .A1(\RI5[0][116] ), .A2(\RI5[0][140] ), .Z(
        \MC_ARK_ARC_1_0/temp2[170] ) );
  XOR2_X1 U8712 ( .A1(\MC_ARK_ARC_1_3/temp1[21] ), .A2(n5962), .Z(
        \MC_ARK_ARC_1_3/temp5[21] ) );
  XOR2_X1 U8713 ( .A1(\SB2_3_3/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[159] ), .Z(n5962) );
  XOR2_X1 U8715 ( .A1(\MC_ARK_ARC_1_3/temp2[99] ), .A2(n5963), .Z(
        \MC_ARK_ARC_1_3/temp5[99] ) );
  XOR2_X1 U8719 ( .A1(\RI5[3][93] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[99] ), 
        .Z(n5963) );
  XOR2_X1 U8723 ( .A1(\MC_ARK_ARC_1_3/temp2[40] ), .A2(
        \MC_ARK_ARC_1_3/temp1[40] ), .Z(\MC_ARK_ARC_1_3/temp5[40] ) );
  XOR2_X1 U8724 ( .A1(n1131), .A2(n3093), .Z(\MC_ARK_ARC_1_3/buf_output[189] )
         );
  NAND3_X2 U8726 ( .A1(\SB1_3_14/i0[6] ), .A2(\SB1_3_14/i0[10] ), .A3(
        \RI1[3][107] ), .ZN(n5014) );
  NAND3_X1 U8727 ( .A1(\SB4_27/i0_4 ), .A2(\SB4_27/i1_5 ), .A3(\SB4_27/i1[9] ), 
        .ZN(n2217) );
  XOR2_X1 U8735 ( .A1(\RI5[2][62] ), .A2(\RI5[2][86] ), .Z(
        \MC_ARK_ARC_1_2/temp2[116] ) );
  XOR2_X1 U8738 ( .A1(\MC_ARK_ARC_1_2/temp2[103] ), .A2(
        \MC_ARK_ARC_1_2/temp1[103] ), .Z(n6595) );
  NAND4_X2 U8739 ( .A1(n6809), .A2(\SB2_4_16/Component_Function_3/NAND4_in[0] ), .A3(\SB2_4_16/Component_Function_3/NAND4_in[3] ), .A4(n920), .ZN(
        \SB2_4_16/buf_output[3] ) );
  NAND4_X2 U8741 ( .A1(\SB1_1_31/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_31/Component_Function_1/NAND4_in[0] ), .A3(n3712), .A4(
        \SB1_1_31/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_1_31/buf_output[1] ) );
  INV_X2 U8743 ( .I(\SB1_4_19/buf_output[5] ), .ZN(\SB2_4_19/i1_5 ) );
  NAND3_X2 U8744 ( .A1(n3396), .A2(n2467), .A3(
        \SB1_4_19/Component_Function_5/NAND4_in[1] ), .ZN(
        \SB1_4_19/buf_output[5] ) );
  NAND4_X2 U8746 ( .A1(\SB2_2_23/Component_Function_2/NAND4_in[0] ), .A2(n6342), .A3(\SB2_2_23/Component_Function_2/NAND4_in[2] ), .A4(n5964), .ZN(
        \SB2_2_23/buf_output[2] ) );
  NAND3_X2 U8747 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0[10] ), .A3(
        \SB2_2_23/i0[6] ), .ZN(n5964) );
  XOR2_X1 U8748 ( .A1(\SB2_3_31/buf_output[4] ), .A2(\RI5[3][166] ), .Z(n599)
         );
  XOR2_X1 U8751 ( .A1(n5965), .A2(n198), .Z(Ciphertext[165]) );
  NAND4_X2 U8752 ( .A1(n5209), .A2(n3783), .A3(
        \SB4_4/Component_Function_3/NAND4_in[1] ), .A4(
        \SB4_4/Component_Function_3/NAND4_in[3] ), .ZN(n5965) );
  NAND4_X2 U8754 ( .A1(n5011), .A2(\SB2_3_5/Component_Function_4/NAND4_in[0] ), 
        .A3(\SB2_3_5/Component_Function_4/NAND4_in[1] ), .A4(n5966), .ZN(
        \SB2_3_5/buf_output[4] ) );
  NAND3_X1 U8756 ( .A1(\SB2_3_5/i0_3 ), .A2(\SB2_3_5/i0[10] ), .A3(
        \SB2_3_5/i0[9] ), .ZN(n5966) );
  NAND4_X2 U8757 ( .A1(n2043), .A2(n6921), .A3(
        \SB1_3_5/Component_Function_5/NAND4_in[0] ), .A4(n5967), .ZN(
        \SB1_3_5/buf_output[5] ) );
  NAND3_X2 U8761 ( .A1(\SB1_3_5/i0[6] ), .A2(\SB1_3_5/i0[10] ), .A3(
        \SB1_3_5/i0_0 ), .ZN(n5967) );
  XOR2_X1 U8764 ( .A1(\RI5[1][161] ), .A2(\RI5[1][167] ), .Z(n6439) );
  NAND4_X2 U8766 ( .A1(\SB2_1_25/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_1_25/Component_Function_5/NAND4_in[3] ), .A3(n3436), .A4(n5968), 
        .ZN(\SB2_1_25/buf_output[5] ) );
  NAND3_X2 U8767 ( .A1(\SB2_1_25/i0_4 ), .A2(\SB2_1_25/i0_3 ), .A3(
        \SB2_1_25/i1[9] ), .ZN(n5968) );
  XOR2_X1 U8772 ( .A1(n5970), .A2(n5969), .Z(\MC_ARK_ARC_1_2/temp6[153] ) );
  XOR2_X1 U8773 ( .A1(\RI5[2][27] ), .A2(n82), .Z(n5969) );
  XOR2_X1 U8776 ( .A1(\RI5[2][189] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[63] ), 
        .Z(n5970) );
  XOR2_X1 U8777 ( .A1(\MC_ARK_ARC_1_4/temp2[131] ), .A2(n5971), .Z(
        \MC_ARK_ARC_1_4/temp5[131] ) );
  XOR2_X1 U8780 ( .A1(\RI5[4][131] ), .A2(\RI5[4][125] ), .Z(n5971) );
  XOR2_X1 U8782 ( .A1(n6804), .A2(n5972), .Z(\MC_ARK_ARC_1_0/temp5[59] ) );
  XOR2_X1 U8783 ( .A1(\RI5[0][53] ), .A2(\RI5[0][29] ), .Z(n5972) );
  XOR2_X1 U8790 ( .A1(n5973), .A2(n200), .Z(Ciphertext[148]) );
  NAND4_X2 U8795 ( .A1(n2506), .A2(\SB4_7/Component_Function_4/NAND4_in[1] ), 
        .A3(n6222), .A4(n2673), .ZN(n5973) );
  XOR2_X1 U8797 ( .A1(n4930), .A2(n5974), .Z(\MC_ARK_ARC_1_3/buf_output[124] )
         );
  XOR2_X1 U8798 ( .A1(\MC_ARK_ARC_1_3/temp1[124] ), .A2(
        \MC_ARK_ARC_1_3/temp2[124] ), .Z(n5974) );
  BUF_X4 U8799 ( .I(\MC_ARK_ARC_1_3/buf_output[190] ), .Z(\SB1_4_0/i0_4 ) );
  NAND4_X2 U8801 ( .A1(\SB2_3_24/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_24/Component_Function_3/NAND4_in[0] ), .A3(n3924), .A4(n5975), 
        .ZN(\SB2_3_24/buf_output[3] ) );
  NAND3_X2 U8802 ( .A1(\SB2_3_24/i0[10] ), .A2(\SB2_3_24/i1[9] ), .A3(
        \SB2_3_24/i1_7 ), .ZN(n5975) );
  NAND4_X2 U8803 ( .A1(\SB1_1_10/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_10/Component_Function_2/NAND4_in[0] ), .A3(n7454), .A4(n5976), 
        .ZN(\SB1_1_10/buf_output[2] ) );
  NAND3_X2 U8805 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i0[9] ), .A3(
        \SB1_1_10/i0[8] ), .ZN(n5976) );
  XOR2_X1 U8806 ( .A1(\RI5[1][87] ), .A2(\RI5[1][81] ), .Z(
        \MC_ARK_ARC_1_1/temp1[87] ) );
  NAND4_X2 U8807 ( .A1(\SB2_3_0/Component_Function_4/NAND4_in[3] ), .A2(n7288), 
        .A3(n7072), .A4(n5977), .ZN(\SB2_3_0/buf_output[4] ) );
  AOI21_X2 U8808 ( .A1(\SB2_4_12/i0_0 ), .A2(\SB2_4_12/i3[0] ), .B(n5978), 
        .ZN(n5403) );
  INV_X1 U8811 ( .I(n5979), .ZN(n5978) );
  NAND3_X1 U8817 ( .A1(\SB1_4_16/buf_output[1] ), .A2(\SB1_4_13/buf_output[4] ), .A3(\SB1_4_17/buf_output[0] ), .ZN(n5979) );
  INV_X2 U8821 ( .I(\SB3_30/buf_output[3] ), .ZN(\SB4_28/i0[8] ) );
  NAND4_X2 U8822 ( .A1(\SB3_30/Component_Function_3/NAND4_in[1] ), .A2(n2312), 
        .A3(\SB3_30/Component_Function_3/NAND4_in[0] ), .A4(n6970), .ZN(
        \SB3_30/buf_output[3] ) );
  XOR2_X1 U8824 ( .A1(\MC_ARK_ARC_1_1/temp2[125] ), .A2(n5980), .Z(
        \MC_ARK_ARC_1_1/temp5[125] ) );
  XOR2_X1 U8825 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[125] ), .A2(\RI5[1][119] ), 
        .Z(n5980) );
  NAND4_X2 U8827 ( .A1(n7341), .A2(\SB2_3_0/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB2_3_0/Component_Function_2/NAND4_in[2] ), .A4(n5981), .ZN(
        \SB2_3_0/buf_output[2] ) );
  NAND3_X2 U8834 ( .A1(\SB2_3_0/i0[10] ), .A2(\SB2_3_0/i1_5 ), .A3(
        \SB2_3_0/i1[9] ), .ZN(n5981) );
  NAND4_X2 U8838 ( .A1(n5128), .A2(n2981), .A3(
        \SB1_2_21/Component_Function_5/NAND4_in[0] ), .A4(n5982), .ZN(
        \SB1_2_21/buf_output[5] ) );
  NAND3_X2 U8845 ( .A1(\SB1_2_21/i0[6] ), .A2(\SB1_2_21/i0[10] ), .A3(
        \SB1_2_21/i0_0 ), .ZN(n5982) );
  NAND3_X1 U8851 ( .A1(\SB2_4_31/i0_3 ), .A2(\SB2_4_31/i0[10] ), .A3(
        \SB2_4_31/i0[9] ), .ZN(n3689) );
  NAND3_X2 U8852 ( .A1(\SB2_3_11/i0_3 ), .A2(\SB2_3_11/i0_4 ), .A3(
        \SB2_3_11/i1[9] ), .ZN(n2514) );
  XOR2_X1 U8854 ( .A1(n5984), .A2(n5983), .Z(\MC_ARK_ARC_1_0/buf_output[107] )
         );
  XOR2_X1 U8857 ( .A1(n4086), .A2(n5182), .Z(n5984) );
  NAND3_X1 U8858 ( .A1(\SB2_4_25/i0_3 ), .A2(\SB2_4_25/i0_0 ), .A3(
        \SB2_4_25/i0[7] ), .ZN(n2606) );
  NAND4_X2 U8860 ( .A1(\SB1_0_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_3/Component_Function_3/NAND4_in[3] ), .A3(n6981), .A4(n833), 
        .ZN(\RI3[0][183] ) );
  XOR2_X1 U8864 ( .A1(n2440), .A2(n5985), .Z(n7162) );
  XOR2_X1 U8868 ( .A1(\SB2_0_2/buf_output[3] ), .A2(\RI5[0][183] ), .Z(n5985)
         );
  XOR2_X1 U8869 ( .A1(n5987), .A2(n5986), .Z(n2137) );
  XOR2_X1 U8874 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), .A2(n554), .Z(
        n5986) );
  XOR2_X1 U8875 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[110] ), .A2(\RI5[2][80] ), 
        .Z(n5987) );
  NAND3_X1 U8877 ( .A1(\SB1_3_24/i0[6] ), .A2(\SB1_3_24/i0_0 ), .A3(
        \SB1_3_24/i0[10] ), .ZN(\SB1_3_24/Component_Function_5/NAND4_in[1] )
         );
  NOR2_X2 U8878 ( .A1(n6231), .A2(n2546), .ZN(n2657) );
  XOR2_X1 U8879 ( .A1(\SB2_3_28/buf_output[2] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[62] ), .Z(n2837) );
  XOR2_X1 U8881 ( .A1(\SB2_4_27/buf_output[2] ), .A2(\RI5[4][14] ), .Z(n6526)
         );
  XOR2_X1 U8883 ( .A1(n3004), .A2(n5988), .Z(n6884) );
  XOR2_X1 U8884 ( .A1(\RI5[2][33] ), .A2(\RI5[2][27] ), .Z(n5988) );
  NAND2_X2 U8885 ( .A1(\SB1_1_8/i0[9] ), .A2(n5989), .ZN(n5177) );
  AND2_X1 U8887 ( .A1(\MC_ARK_ARC_1_0/buf_output[139] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[142] ), .Z(n5989) );
  NAND4_X2 U8890 ( .A1(\SB1_4_14/Component_Function_4/NAND4_in[0] ), .A2(n6778), .A3(\SB1_4_14/Component_Function_4/NAND4_in[1] ), .A4(n5990), .ZN(
        \SB1_4_14/buf_output[4] ) );
  NAND4_X2 U8900 ( .A1(\SB2_4_13/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_13/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_4_13/Component_Function_0/NAND4_in[0] ), .A4(n5991), .ZN(
        \SB2_4_13/buf_output[0] ) );
  NAND3_X1 U8903 ( .A1(\SB2_4_13/i0_4 ), .A2(\SB2_4_13/i0_3 ), .A3(
        \SB2_4_13/i0[10] ), .ZN(n5991) );
  INV_X2 U8909 ( .I(\SB1_2_14/buf_output[3] ), .ZN(\SB2_2_12/i0[8] ) );
  NAND4_X2 U8912 ( .A1(\SB1_2_14/Component_Function_3/NAND4_in[1] ), .A2(n7126), .A3(n3005), .A4(n7068), .ZN(\SB1_2_14/buf_output[3] ) );
  INV_X2 U8914 ( .I(\SB1_1_13/buf_output[2] ), .ZN(\SB2_1_10/i1[9] ) );
  NAND4_X2 U8922 ( .A1(\SB1_1_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_1_13/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_1_13/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_1_13/buf_output[2] ) );
  XOR2_X1 U8927 ( .A1(\MC_ARK_ARC_1_3/temp5[178] ), .A2(n5992), .Z(
        \MC_ARK_ARC_1_3/buf_output[178] ) );
  XOR2_X1 U8939 ( .A1(\MC_ARK_ARC_1_3/temp4[178] ), .A2(
        \MC_ARK_ARC_1_3/temp3[178] ), .Z(n5992) );
  XOR2_X1 U8948 ( .A1(\MC_ARK_ARC_1_3/temp6[106] ), .A2(n5993), .Z(
        \MC_ARK_ARC_1_3/buf_output[106] ) );
  XOR2_X1 U8950 ( .A1(\MC_ARK_ARC_1_3/temp2[106] ), .A2(
        \MC_ARK_ARC_1_3/temp1[106] ), .Z(n5993) );
  NAND2_X2 U8951 ( .A1(n5046), .A2(n5994), .ZN(n3512) );
  INV_X2 U8953 ( .I(\RI3[0][27] ), .ZN(\SB2_0_27/i0[8] ) );
  NAND4_X2 U8955 ( .A1(\SB1_0_29/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_29/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_0_29/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_0_29/Component_Function_3/NAND4_in[2] ), .ZN(\RI3[0][27] ) );
  XOR2_X1 U8964 ( .A1(\MC_ARK_ARC_1_3/temp1[26] ), .A2(n5995), .Z(
        \MC_ARK_ARC_1_3/temp5[26] ) );
  XOR2_X1 U8967 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[164] ), .A2(n1506), .Z(
        n5995) );
  XOR2_X1 U8968 ( .A1(n1952), .A2(n5996), .Z(\MC_ARK_ARC_1_1/buf_output[31] )
         );
  XOR2_X1 U8969 ( .A1(n7373), .A2(n6337), .Z(n5996) );
  INV_X2 U8970 ( .I(\SB1_3_14/buf_output[5] ), .ZN(\SB2_3_14/i1_5 ) );
  XOR2_X1 U8972 ( .A1(\RI5[2][128] ), .A2(\RI5[2][152] ), .Z(n5997) );
  XOR2_X1 U8974 ( .A1(\MC_ARK_ARC_1_2/temp5[19] ), .A2(n5998), .Z(
        \MC_ARK_ARC_1_2/buf_output[19] ) );
  XOR2_X1 U8975 ( .A1(\MC_ARK_ARC_1_2/temp3[19] ), .A2(
        \MC_ARK_ARC_1_2/temp4[19] ), .Z(n5998) );
  XOR2_X1 U8976 ( .A1(n6004), .A2(\MC_ARK_ARC_1_3/temp4[91] ), .Z(n5078) );
  NAND3_X1 U8981 ( .A1(\SB1_4_17/i0_3 ), .A2(\SB1_4_17/i0_4 ), .A3(
        \SB1_4_17/i1[9] ), .ZN(n5006) );
  XOR2_X1 U8984 ( .A1(n5295), .A2(n5999), .Z(\MC_ARK_ARC_1_3/temp5[7] ) );
  XOR2_X1 U8986 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[1] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[7] ), .Z(n5999) );
  NAND4_X2 U8988 ( .A1(\SB2_3_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_30/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_30/Component_Function_4/NAND4_in[1] ), .A4(n6000), .ZN(
        \SB2_3_30/buf_output[4] ) );
  NAND3_X1 U8989 ( .A1(\SB2_3_30/i0[10] ), .A2(\SB2_3_30/i0_3 ), .A3(
        \SB1_3_3/buf_output[0] ), .ZN(n6000) );
  NAND4_X2 U8992 ( .A1(\SB4_19/Component_Function_5/NAND4_in[1] ), .A2(n7132), 
        .A3(\SB4_19/Component_Function_5/NAND4_in[0] ), .A4(n6001), .ZN(n6936)
         );
  NAND3_X1 U8993 ( .A1(\SB4_19/i0[6] ), .A2(\SB4_19/i0_4 ), .A3(\SB4_19/i0[9] ), .ZN(n6001) );
  NAND3_X2 U8995 ( .A1(\SB2_1_11/i1[9] ), .A2(\SB2_1_11/i1_5 ), .A3(
        \SB2_1_11/i0_4 ), .ZN(\SB2_1_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U8996 ( .A1(\SB2_2_26/i0_3 ), .A2(\SB2_2_26/i1_7 ), .A3(
        \SB2_2_26/i0[8] ), .ZN(\SB2_2_26/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U8997 ( .A1(\RI5[0][47] ), .A2(\RI5[0][11] ), .Z(
        \MC_ARK_ARC_1_0/temp3[137] ) );
  NAND4_X2 U9000 ( .A1(\SB1_2_10/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_2_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_10/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_2_10/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[2][131] ) );
  XOR2_X1 U9002 ( .A1(n6002), .A2(\MC_ARK_ARC_1_3/temp4[131] ), .Z(n1826) );
  XOR2_X1 U9003 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[5] ), .A2(\RI5[3][41] ), 
        .Z(n6002) );
  NAND3_X2 U9005 ( .A1(\SB2_0_22/i0_3 ), .A2(\RI3[0][55] ), .A3(
        \SB2_0_22/i0[10] ), .ZN(\SB2_0_22/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U9006 ( .A1(\MC_ARK_ARC_1_4/temp4[29] ), .A2(n6003), .Z(n1356) );
  XOR2_X1 U9008 ( .A1(\RI5[4][95] ), .A2(\RI5[4][131] ), .Z(n6003) );
  XOR2_X1 U9009 ( .A1(\SB2_3_21/buf_output[1] ), .A2(\RI5[3][91] ), .Z(n6004)
         );
  NAND3_X2 U9010 ( .A1(\SB1_1_1/i0[10] ), .A2(\SB1_1_1/i0_3 ), .A3(
        \SB1_1_1/i0[6] ), .ZN(n6005) );
  XOR2_X1 U9016 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), .A2(\RI5[2][185] ), 
        .Z(n6006) );
  NAND3_X2 U9017 ( .A1(\SB4_0/i0_4 ), .A2(\SB4_0/i0_0 ), .A3(\SB4_0/i1_5 ), 
        .ZN(n6007) );
  XOR2_X1 U9018 ( .A1(n6009), .A2(n6008), .Z(\MC_ARK_ARC_1_4/temp6[33] ) );
  XOR2_X1 U9025 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[135] ), .A2(n468), .Z(
        n6008) );
  XOR2_X1 U9026 ( .A1(\RI5[4][69] ), .A2(\RI5[4][99] ), .Z(n6009) );
  BUF_X4 U9036 ( .I(\MC_ARK_ARC_1_4/buf_output[95] ), .Z(\SB3_16/i0_3 ) );
  NAND3_X2 U9042 ( .A1(\SB2_3_30/i0_4 ), .A2(\SB2_3_30/i0_0 ), .A3(
        \SB2_3_30/i1_5 ), .ZN(n6135) );
  INV_X1 U9043 ( .I(\SB1_4_22/buf_output[5] ), .ZN(\SB2_4_22/i1_5 ) );
  NAND4_X2 U9047 ( .A1(\SB1_4_22/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_4_22/Component_Function_5/NAND4_in[1] ), .A3(n6082), .A4(n1091), 
        .ZN(\SB1_4_22/buf_output[5] ) );
  XOR2_X1 U9049 ( .A1(\MC_ARK_ARC_1_0/temp2[110] ), .A2(n6010), .Z(n3301) );
  XOR2_X1 U9051 ( .A1(\RI5[0][20] ), .A2(\RI5[0][176] ), .Z(n6010) );
  NAND3_X1 U9052 ( .A1(\SB4_22/i0[6] ), .A2(\SB4_22/i0_3 ), .A3(\SB4_22/i1[9] ), .ZN(n6011) );
  NAND4_X2 U9057 ( .A1(\SB1_4_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_4_23/Component_Function_1/NAND4_in[0] ), .A3(n7203), .A4(n6012), 
        .ZN(\SB1_4_23/buf_output[1] ) );
  NAND3_X2 U9058 ( .A1(\SB1_4_23/i0[6] ), .A2(\SB1_4_23/i0[9] ), .A3(
        \SB1_4_23/i1_5 ), .ZN(n6012) );
  BUF_X2 U9060 ( .I(\SB3_1/buf_output[1] ), .Z(\SB4_29/i0[6] ) );
  NAND4_X2 U9063 ( .A1(\SB2_4_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_17/Component_Function_3/NAND4_in[3] ), .A3(n939), .A4(n6013), 
        .ZN(\SB2_4_17/buf_output[3] ) );
  NAND3_X2 U9064 ( .A1(\SB2_4_17/i0_4 ), .A2(\SB2_4_17/i0_3 ), .A3(
        \SB2_4_17/i0_0 ), .ZN(n6013) );
  NAND4_X2 U9066 ( .A1(\SB1_4_7/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_4_7/Component_Function_2/NAND4_in[2] ), .A3(n4062), .A4(n6014), 
        .ZN(\SB1_4_7/buf_output[2] ) );
  NAND3_X2 U9067 ( .A1(\SB1_4_7/i0_4 ), .A2(\SB1_4_7/i0_0 ), .A3(
        \SB1_4_7/i1_5 ), .ZN(n6014) );
  NAND4_X2 U9069 ( .A1(\SB1_2_1/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_1/Component_Function_0/NAND4_in[0] ), .A4(n6015), .ZN(
        \SB1_2_1/buf_output[0] ) );
  NAND3_X1 U9072 ( .A1(\SB1_2_1/i0_0 ), .A2(\SB1_2_1/i0_3 ), .A3(
        \SB1_2_1/i0[7] ), .ZN(n6015) );
  BUF_X4 U9075 ( .I(\SB1_4_12/buf_output[1] ), .Z(\SB2_4_8/i0[6] ) );
  NAND3_X2 U9077 ( .A1(\SB3_26/i0_0 ), .A2(\SB3_26/i1_5 ), .A3(\SB3_26/i0_4 ), 
        .ZN(n7293) );
  NAND3_X2 U9078 ( .A1(\SB2_1_13/i0_0 ), .A2(\SB2_1_13/i0[6] ), .A3(
        \SB2_1_13/i0[10] ), .ZN(n6447) );
  NAND4_X2 U9079 ( .A1(\SB2_3_2/Component_Function_2/NAND4_in[0] ), .A2(n1092), 
        .A3(n6114), .A4(n1925), .ZN(\SB2_3_2/buf_output[2] ) );
  NAND4_X2 U9080 ( .A1(\SB1_4_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_4_14/Component_Function_2/NAND4_in[2] ), .A3(n6879), .A4(n6220), 
        .ZN(\SB1_4_14/buf_output[2] ) );
  BUF_X4 U9082 ( .I(\MC_ARK_ARC_1_3/buf_output[80] ), .Z(\SB1_4_18/i0_0 ) );
  XOR2_X1 U9084 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[41] ), .A2(\RI5[0][65] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[95] ) );
  XOR2_X1 U9086 ( .A1(\RI5[3][2] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[158] ), 
        .Z(n6088) );
  NAND3_X2 U9088 ( .A1(\SB2_4_13/i0_4 ), .A2(\SB2_4_13/i0_3 ), .A3(
        \SB2_4_13/i1[9] ), .ZN(n3041) );
  XOR2_X1 U9090 ( .A1(\RI5[3][23] ), .A2(\RI5[3][179] ), .Z(
        \MC_ARK_ARC_1_3/temp3[113] ) );
  NAND4_X2 U9091 ( .A1(\SB2_4_18/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_4_18/Component_Function_0/NAND4_in[1] ), .A3(n6127), .A4(
        \SB2_4_18/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_4_18/buf_output[0] ) );
  XOR2_X1 U9093 ( .A1(\RI5[1][60] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[114] ) );
  NAND3_X1 U9094 ( .A1(\SB1_4_13/i0[10] ), .A2(\SB1_4_13/i0_3 ), .A3(
        \SB1_4_13/i0_4 ), .ZN(\SB1_4_13/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U9097 ( .A1(\RI5[3][134] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[170] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[68] ) );
  XOR2_X1 U9099 ( .A1(\RI5[2][125] ), .A2(\RI5[2][119] ), .Z(
        \MC_ARK_ARC_1_2/temp1[125] ) );
  XOR2_X1 U9101 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[14] ), .A2(\RI5[2][8] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[14] ) );
  BUF_X4 U9102 ( .I(\SB2_4_18/buf_output[1] ), .Z(\RI5[4][103] ) );
  INV_X1 U9108 ( .I(\SB3_5/buf_output[5] ), .ZN(\SB4_5/i1_5 ) );
  NAND4_X2 U9109 ( .A1(\SB3_5/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_5/Component_Function_5/NAND4_in[2] ), .A3(
        \SB3_5/Component_Function_5/NAND4_in[3] ), .A4(
        \SB3_5/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_5/buf_output[5] )
         );
  AND2_X1 U9111 ( .A1(n1196), .A2(n6504), .Z(n7523) );
  XOR2_X1 U9112 ( .A1(\MC_ARK_ARC_1_3/temp2[94] ), .A2(n6016), .Z(n4946) );
  XOR2_X1 U9115 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[94] ), .A2(\RI5[3][88] ), 
        .Z(n6016) );
  XOR2_X1 U9128 ( .A1(\RI5[1][29] ), .A2(\RI5[1][185] ), .Z(
        \MC_ARK_ARC_1_1/temp3[119] ) );
  INV_X2 U9136 ( .I(\SB1_1_30/buf_output[3] ), .ZN(\SB2_1_28/i0[8] ) );
  NAND3_X1 U9138 ( .A1(\SB3_25/i0[10] ), .A2(\SB3_25/i0_3 ), .A3(
        \SB3_25/i0[9] ), .ZN(n6064) );
  NAND3_X2 U9140 ( .A1(\SB4_6/i0[10] ), .A2(\SB4_6/i0[6] ), .A3(\SB4_6/i0_3 ), 
        .ZN(n6017) );
  AND2_X1 U9143 ( .A1(\SB2_0_31/i1_7 ), .A2(\SB2_0_31/i3[0] ), .Z(n6533) );
  NAND4_X2 U9144 ( .A1(n2364), .A2(\SB2_3_24/Component_Function_5/NAND4_in[3] ), .A3(\SB2_3_24/Component_Function_5/NAND4_in[0] ), .A4(n6018), .ZN(
        \SB2_3_24/buf_output[5] ) );
  NAND3_X2 U9145 ( .A1(\SB2_3_24/i0[10] ), .A2(\SB2_3_24/i0_0 ), .A3(
        \SB2_3_24/i0[6] ), .ZN(n6018) );
  XOR2_X1 U9146 ( .A1(n4474), .A2(n6019), .Z(\MC_ARK_ARC_1_1/buf_output[26] )
         );
  XOR2_X1 U9148 ( .A1(\MC_ARK_ARC_1_1/temp2[4] ), .A2(n6020), .Z(
        \MC_ARK_ARC_1_1/temp5[4] ) );
  XOR2_X1 U9149 ( .A1(\RI5[1][190] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[4] ), 
        .Z(n6020) );
  NAND4_X2 U9152 ( .A1(\SB2_2_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_30/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_30/Component_Function_2/NAND4_in[1] ), .A4(n6021), .ZN(
        \SB2_2_30/buf_output[2] ) );
  NAND3_X2 U9157 ( .A1(\SB2_2_30/i0_4 ), .A2(\SB2_2_30/i0_0 ), .A3(
        \SB2_2_30/i1_5 ), .ZN(n6021) );
  NAND4_X2 U9159 ( .A1(n4950), .A2(\SB1_1_1/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB1_1_1/Component_Function_5/NAND4_in[2] ), .A4(n6022), .ZN(
        \SB1_1_1/buf_output[5] ) );
  NAND3_X1 U9162 ( .A1(\SB1_2_31/i0_4 ), .A2(\SB1_2_31/i1[9] ), .A3(
        \SB1_2_31/i1_5 ), .ZN(\SB1_2_31/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U9163 ( .A1(\SB3_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_7/Component_Function_0/NAND4_in[3] ), .A3(
        \SB3_7/Component_Function_0/NAND4_in[0] ), .A4(n6023), .ZN(
        \SB3_7/buf_output[0] ) );
  NAND3_X1 U9166 ( .A1(\SB3_7/i0[6] ), .A2(\SB3_7/i0[8] ), .A3(\SB3_7/i0[7] ), 
        .ZN(n6023) );
  XOR2_X1 U9167 ( .A1(n6025), .A2(n6024), .Z(\MC_ARK_ARC_1_0/buf_output[131] )
         );
  XOR2_X1 U9169 ( .A1(\MC_ARK_ARC_1_0/temp1[131] ), .A2(
        \MC_ARK_ARC_1_0/temp4[131] ), .Z(n6024) );
  XOR2_X1 U9172 ( .A1(n2670), .A2(n5262), .Z(n6025) );
  XOR2_X1 U9173 ( .A1(n6026), .A2(n23), .Z(Ciphertext[40]) );
  NAND4_X2 U9174 ( .A1(\SB4_25/Component_Function_4/NAND4_in[1] ), .A2(
        \SB4_25/Component_Function_4/NAND4_in[3] ), .A3(
        \SB4_25/Component_Function_4/NAND4_in[0] ), .A4(n7566), .ZN(n6026) );
  XOR2_X1 U9175 ( .A1(n6028), .A2(n6027), .Z(\MC_ARK_ARC_1_1/buf_output[47] )
         );
  XOR2_X1 U9177 ( .A1(n6128), .A2(n4457), .Z(n6027) );
  XOR2_X1 U9181 ( .A1(\MC_ARK_ARC_1_1/temp2[47] ), .A2(n4458), .Z(n6028) );
  XOR2_X1 U9182 ( .A1(n1259), .A2(n6029), .Z(\MC_ARK_ARC_1_4/temp5[53] ) );
  XOR2_X1 U9184 ( .A1(\RI5[4][47] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[53] ), 
        .Z(n6029) );
  BUF_X4 U9188 ( .I(\RI3[0][95] ), .Z(\SB2_0_16/i0_3 ) );
  NAND4_X2 U9192 ( .A1(\SB1_1_5/Component_Function_5/NAND4_in[1] ), .A2(n4442), 
        .A3(n6620), .A4(\SB1_1_5/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_5/buf_output[5] ) );
  BUF_X4 U9200 ( .I(\SB2_4_29/buf_output[0] ), .Z(\RI5[4][42] ) );
  XOR2_X1 U9205 ( .A1(\MC_ARK_ARC_1_0/temp1[160] ), .A2(n6030), .Z(n7157) );
  XOR2_X1 U9207 ( .A1(\RI5[0][106] ), .A2(\RI5[0][130] ), .Z(n6030) );
  NAND4_X2 U9213 ( .A1(\SB2_0_10/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_0_10/Component_Function_2/NAND4_in[2] ), .A4(n6031), .ZN(
        \SB2_0_10/buf_output[2] ) );
  NAND3_X2 U9222 ( .A1(\SB1_1_24/i1[9] ), .A2(\RI1[1][47] ), .A3(
        \MC_ARK_ARC_1_0/buf_output[46] ), .ZN(n6474) );
  NAND3_X1 U9233 ( .A1(\SB1_4_3/i0_3 ), .A2(\SB1_4_3/i0_0 ), .A3(
        \SB1_4_3/i0_4 ), .ZN(\SB1_4_3/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U9242 ( .A1(\SB2_4_1/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_4_1/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_4_1/Component_Function_0/NAND4_in[0] ), .A4(n4302), .ZN(
        \SB2_4_1/buf_output[0] ) );
  XOR2_X1 U9244 ( .A1(n4613), .A2(n6033), .Z(n4191) );
  XOR2_X1 U9245 ( .A1(\RI5[4][140] ), .A2(\RI5[4][146] ), .Z(n6033) );
  XOR2_X1 U9250 ( .A1(n3874), .A2(n5362), .Z(n7503) );
  XOR2_X1 U9251 ( .A1(\SB2_0_31/buf_output[1] ), .A2(\RI5[0][19] ), .Z(
        \MC_ARK_ARC_1_0/temp1[25] ) );
  NAND4_X2 U9255 ( .A1(\SB2_0_0/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_0/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_0_0/Component_Function_1/NAND4_in[0] ), .A4(n6034), .ZN(
        \SB2_0_0/buf_output[1] ) );
  NAND4_X2 U9258 ( .A1(n7180), .A2(\SB2_0_15/Component_Function_4/NAND4_in[3] ), .A3(\SB2_0_15/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_0_15/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB2_0_15/buf_output[4] ) );
  NAND4_X2 U9262 ( .A1(\SB2_2_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_6/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_2_6/Component_Function_2/NAND4_in[1] ), .A4(n6035), .ZN(
        \SB2_2_6/buf_output[2] ) );
  NAND3_X2 U9270 ( .A1(\SB2_2_6/i0_3 ), .A2(\SB2_2_6/i0[9] ), .A3(
        \SB2_2_6/i0[8] ), .ZN(n6035) );
  BUF_X4 U9272 ( .I(\MC_ARK_ARC_1_3/buf_output[167] ), .Z(\SB1_4_4/i0_3 ) );
  XOR2_X1 U9275 ( .A1(n6036), .A2(n110), .Z(Ciphertext[87]) );
  NAND4_X2 U9277 ( .A1(\SB4_17/Component_Function_3/NAND4_in[2] ), .A2(
        \SB4_17/Component_Function_3/NAND4_in[0] ), .A3(n6935), .A4(
        \SB4_17/Component_Function_3/NAND4_in[1] ), .ZN(n6036) );
  NAND4_X2 U9279 ( .A1(n5100), .A2(\SB3_20/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB3_20/Component_Function_2/NAND4_in[0] ), .A4(n6037), .ZN(
        \SB3_20/buf_output[2] ) );
  NAND3_X2 U9289 ( .A1(\SB3_20/i0_4 ), .A2(\SB3_20/i0_0 ), .A3(\SB3_20/i1_5 ), 
        .ZN(n6037) );
  NAND4_X2 U9290 ( .A1(\SB3_28/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_28/Component_Function_1/NAND4_in[0] ), .A3(
        \SB3_28/Component_Function_1/NAND4_in[1] ), .A4(n6038), .ZN(
        \SB3_28/buf_output[1] ) );
  NAND3_X1 U9292 ( .A1(\SB3_28/i0[6] ), .A2(\SB3_28/i1_5 ), .A3(\SB3_28/i0[9] ), .ZN(n6038) );
  NAND4_X2 U9302 ( .A1(\SB1_4_20/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_4_20/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_4_20/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_4_20/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_4_20/buf_output[0] ) );
  XOR2_X1 U9303 ( .A1(\RI5[3][98] ), .A2(\RI5[3][122] ), .Z(
        \MC_ARK_ARC_1_3/temp2[152] ) );
  NAND4_X2 U9304 ( .A1(\SB2_3_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_24/Component_Function_2/NAND4_in[2] ), .A4(n6039), .ZN(
        \SB2_3_24/buf_output[2] ) );
  NAND3_X2 U9306 ( .A1(\SB2_3_24/i0_0 ), .A2(\SB2_3_24/i0_4 ), .A3(
        \SB2_3_24/i1_5 ), .ZN(n6039) );
  NAND4_X2 U9308 ( .A1(\SB2_2_21/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_21/Component_Function_4/NAND4_in[0] ), .A4(n6040), .ZN(
        \SB2_2_21/buf_output[4] ) );
  NAND3_X2 U9311 ( .A1(\SB1_1_16/i0_0 ), .A2(\SB1_1_16/i0[10] ), .A3(
        \SB1_1_16/i0[6] ), .ZN(n6041) );
  XOR2_X1 U9312 ( .A1(\MC_ARK_ARC_1_3/temp2[50] ), .A2(n6042), .Z(
        \MC_ARK_ARC_1_3/temp5[50] ) );
  XOR2_X1 U9314 ( .A1(\RI5[3][50] ), .A2(\RI5[3][44] ), .Z(n6042) );
  XOR2_X1 U9316 ( .A1(\RI5[4][101] ), .A2(\RI5[4][155] ), .Z(n2442) );
  XOR2_X1 U9317 ( .A1(\MC_ARK_ARC_1_1/temp1[77] ), .A2(n6043), .Z(
        \MC_ARK_ARC_1_1/temp5[77] ) );
  XOR2_X1 U9318 ( .A1(\RI5[1][47] ), .A2(\RI5[1][23] ), .Z(n6043) );
  NAND3_X1 U9319 ( .A1(\SB4_16/i0[6] ), .A2(\SB4_16/i0[9] ), .A3(\SB4_16/i1_5 ), .ZN(n6045) );
  NAND3_X2 U9321 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0[8] ), .A3(
        \SB2_3_26/i0[9] ), .ZN(\SB2_3_26/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U9322 ( .I(\MC_ARK_ARC_1_4/buf_output[122] ), .Z(\SB3_11/i0_0 ) );
  XOR2_X1 U9323 ( .A1(n6047), .A2(n6046), .Z(\MC_ARK_ARC_1_2/buf_output[29] )
         );
  XOR2_X1 U9324 ( .A1(\MC_ARK_ARC_1_2/temp3[29] ), .A2(
        \MC_ARK_ARC_1_2/temp4[29] ), .Z(n6046) );
  XOR2_X1 U9325 ( .A1(\MC_ARK_ARC_1_2/temp2[29] ), .A2(
        \MC_ARK_ARC_1_2/temp1[29] ), .Z(n6047) );
  BUF_X4 U9326 ( .I(n3970), .Z(\SB3_11/i0_3 ) );
  NAND3_X1 U9330 ( .A1(\SB2_2_28/i0_4 ), .A2(\SB2_2_28/i1_5 ), .A3(
        \SB2_2_28/i1[9] ), .ZN(\SB2_2_28/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U9331 ( .A1(\SB1_4_28/Component_Function_2/NAND4_in[1] ), .A2(n2172), .A3(\SB1_4_28/Component_Function_2/NAND4_in[2] ), .A4(n6048), .ZN(
        \SB1_4_28/buf_output[2] ) );
  NAND3_X2 U9332 ( .A1(\SB1_4_28/i0[10] ), .A2(\SB1_4_28/i1[9] ), .A3(
        \SB1_4_28/i1_5 ), .ZN(n6048) );
  XOR2_X1 U9335 ( .A1(\RI5[0][153] ), .A2(\RI5[0][147] ), .Z(n4182) );
  XOR2_X1 U9336 ( .A1(n6049), .A2(\MC_ARK_ARC_1_3/temp2[19] ), .Z(n1315) );
  XOR2_X1 U9338 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[19] ), .A2(\RI5[3][13] ), 
        .Z(n6049) );
  NAND4_X2 U9339 ( .A1(\SB1_2_31/Component_Function_2/NAND4_in[1] ), .A2(n1618), .A3(\SB1_2_31/Component_Function_2/NAND4_in[0] ), .A4(n6050), .ZN(
        \SB1_2_31/buf_output[2] ) );
  NAND3_X1 U9340 ( .A1(\SB1_2_31/i0[9] ), .A2(\SB1_2_31/i0[8] ), .A3(
        \SB1_2_31/i0_3 ), .ZN(n6050) );
  XOR2_X1 U9341 ( .A1(n7170), .A2(n6051), .Z(\MC_ARK_ARC_1_2/buf_output[22] )
         );
  XOR2_X1 U9342 ( .A1(\MC_ARK_ARC_1_2/temp3[22] ), .A2(
        \MC_ARK_ARC_1_2/temp4[22] ), .Z(n6051) );
  NAND4_X2 U9343 ( .A1(\SB1_1_12/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_12/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_1_12/Component_Function_3/NAND4_in[1] ), .A4(n6768), .ZN(
        \SB1_1_12/buf_output[3] ) );
  NAND4_X2 U9344 ( .A1(\SB2_0_15/Component_Function_2/NAND4_in[0] ), .A2(n7187), .A3(\SB2_0_15/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_15/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_15/buf_output[2] ) );
  NAND3_X1 U9348 ( .A1(\SB1_4_24/i0[6] ), .A2(\SB1_4_24/i1[9] ), .A3(
        \SB1_4_24/i0_3 ), .ZN(\SB1_4_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U9350 ( .A1(\SB2_2_25/i0[10] ), .A2(\SB2_2_25/i1_5 ), .A3(
        \SB2_2_25/i1[9] ), .ZN(\SB2_2_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U9351 ( .A1(\SB4_31/i0[10] ), .A2(\SB4_31/i1_7 ), .A3(
        \SB4_31/i1[9] ), .ZN(\SB4_31/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U9353 ( .A1(\SB1_0_30/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_30/Component_Function_5/NAND4_in[2] ), .A3(n6185), .A4(
        \SB1_0_30/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_30/buf_output[5] ) );
  BUF_X4 U9354 ( .I(\MC_ARK_ARC_1_2/buf_output[87] ), .Z(\SB1_3_17/i0[10] ) );
  NAND4_X2 U9355 ( .A1(\SB2_3_18/Component_Function_5/NAND4_in[2] ), .A2(n2932), .A3(n6122), .A4(\SB2_3_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_18/buf_output[5] ) );
  NAND3_X1 U9356 ( .A1(\SB1_4_23/i0_3 ), .A2(\SB1_4_23/i0[8] ), .A3(
        \SB1_4_23/i1_7 ), .ZN(\SB1_4_23/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U9360 ( .A1(\RI5[4][133] ), .A2(\RI5[4][109] ), .Z(
        \MC_ARK_ARC_1_4/temp2[163] ) );
  XOR2_X1 U9362 ( .A1(\RI5[3][51] ), .A2(\RI5[3][45] ), .Z(
        \MC_ARK_ARC_1_3/temp1[51] ) );
  NAND4_X2 U9363 ( .A1(\SB1_0_23/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_23/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_0_23/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_23/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[0][68] ) );
  NAND3_X2 U9366 ( .A1(\SB1_1_3/i0[10] ), .A2(\SB1_1_3/i1[9] ), .A3(
        \SB1_1_3/i1_7 ), .ZN(n6060) );
  XOR2_X1 U9367 ( .A1(\RI5[0][80] ), .A2(\RI5[0][44] ), .Z(
        \MC_ARK_ARC_1_0/temp3[170] ) );
  XOR2_X1 U9369 ( .A1(\RI5[3][83] ), .A2(\RI5[3][131] ), .Z(n1999) );
  XOR2_X1 U9371 ( .A1(n7477), .A2(\MC_ARK_ARC_1_3/temp6[43] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[43] ) );
  XOR2_X1 U9372 ( .A1(\MC_ARK_ARC_1_1/temp6[183] ), .A2(n4730), .Z(
        \MC_ARK_ARC_1_1/buf_output[183] ) );
  NAND3_X1 U9374 ( .A1(\SB1_4_24/i0[6] ), .A2(\SB1_4_24/i0_0 ), .A3(
        \SB1_4_24/i0[10] ), .ZN(\SB1_4_24/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U9384 ( .A1(\SB1_1_9/i0_4 ), .A2(\SB1_1_9/i1_7 ), .A3(
        \SB1_1_9/i0[8] ), .ZN(\SB1_1_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U9389 ( .A1(\SB3_11/i0[9] ), .A2(\SB3_11/i0[8] ), .A3(\SB3_11/i0_0 ), .ZN(\SB3_11/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U9393 ( .A1(n4967), .A2(\SB3_11/Component_Function_2/NAND4_in[0] ), 
        .A3(\SB3_11/Component_Function_2/NAND4_in[1] ), .A4(
        \SB3_11/Component_Function_2/NAND4_in[2] ), .ZN(\SB4_8/i0_0 ) );
  NAND4_X2 U9394 ( .A1(\SB1_4_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_13/Component_Function_3/NAND4_in[1] ), .A3(n4360), .A4(
        \SB1_4_13/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_4_13/buf_output[3] ) );
  INV_X2 U9395 ( .I(\SB1_2_28/buf_output[3] ), .ZN(\SB2_2_26/i0[8] ) );
  NAND4_X2 U9399 ( .A1(n7548), .A2(\SB1_2_28/Component_Function_3/NAND4_in[1] ), .A3(\SB1_2_28/Component_Function_3/NAND4_in[0] ), .A4(n3455), .ZN(
        \SB1_2_28/buf_output[3] ) );
  INV_X2 U9400 ( .I(\SB1_3_31/buf_output[2] ), .ZN(\SB2_3_28/i1[9] ) );
  XOR2_X1 U9404 ( .A1(\MC_ARK_ARC_1_1/temp6[21] ), .A2(n6054), .Z(
        \MC_ARK_ARC_1_1/buf_output[21] ) );
  XOR2_X1 U9405 ( .A1(n801), .A2(n3664), .Z(n6054) );
  BUF_X4 U9407 ( .I(\SB3_6/buf_output[5] ), .Z(\SB4_6/i0_3 ) );
  NAND3_X1 U9411 ( .A1(\SB3_6/i0[10] ), .A2(\SB3_6/i1[9] ), .A3(\SB3_6/i1_7 ), 
        .ZN(n6055) );
  XOR2_X1 U9412 ( .A1(\RI5[1][100] ), .A2(\SB2_1_22/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/temp3[190] ) );
  NAND4_X2 U9414 ( .A1(\SB1_0_25/Component_Function_2/NAND4_in[0] ), .A2(n2323), .A3(n3303), .A4(\SB1_0_25/Component_Function_2/NAND4_in[3] ), .ZN(
        \RI3[0][56] ) );
  XOR2_X1 U9415 ( .A1(\MC_ARK_ARC_1_2/temp5[108] ), .A2(n6056), .Z(
        \MC_ARK_ARC_1_2/buf_output[108] ) );
  XOR2_X1 U9426 ( .A1(\MC_ARK_ARC_1_2/temp4[108] ), .A2(
        \MC_ARK_ARC_1_2/temp3[108] ), .Z(n6056) );
  NAND3_X2 U9427 ( .A1(\SB1_2_11/i0[10] ), .A2(\SB1_2_11/i1[9] ), .A3(
        \SB1_2_11/i1_7 ), .ZN(n6298) );
  XOR2_X1 U9429 ( .A1(\RI5[0][38] ), .A2(\RI5[0][44] ), .Z(
        \MC_ARK_ARC_1_0/temp1[44] ) );
  NAND3_X2 U9432 ( .A1(\SB2_4_21/i0[6] ), .A2(\SB2_4_21/i0_4 ), .A3(
        \SB2_4_21/i0[9] ), .ZN(n6137) );
  NAND3_X1 U9436 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i1_7 ), .A3(\SB4_16/i3[0] ), 
        .ZN(\SB4_16/Component_Function_4/NAND4_in[1] ) );
  INV_X4 U9439 ( .I(n6057), .ZN(\SB4_6/i1_5 ) );
  XOR2_X1 U9441 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[89] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[65] ), .Z(\MC_ARK_ARC_1_2/temp2[119] )
         );
  NAND4_X2 U9442 ( .A1(\SB1_1_18/Component_Function_5/NAND4_in[1] ), .A2(n5053), .A3(n4852), .A4(\SB1_1_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_18/buf_output[5] ) );
  NAND4_X2 U9447 ( .A1(\SB1_3_31/Component_Function_5/NAND4_in[2] ), .A2(n4760), .A3(\SB1_3_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_3_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_31/buf_output[5] ) );
  NAND4_X2 U9448 ( .A1(\SB2_2_9/Component_Function_5/NAND4_in[3] ), .A2(n2126), 
        .A3(n6244), .A4(\SB2_2_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_9/buf_output[5] ) );
  XOR2_X1 U9454 ( .A1(\RI5[2][137] ), .A2(\RI5[2][101] ), .Z(
        \MC_ARK_ARC_1_2/temp3[35] ) );
  NAND4_X2 U9458 ( .A1(n3865), .A2(n4111), .A3(
        \SB1_2_18/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_2_18/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_2_18/buf_output[4] ) );
  XOR2_X1 U9459 ( .A1(\RI5[0][83] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[77] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[83] ) );
  NAND4_X2 U9460 ( .A1(\SB2_1_30/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_30/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_30/Component_Function_2/NAND4_in[2] ), .A4(n7554), .ZN(
        \SB2_1_30/buf_output[2] ) );
  NAND3_X1 U9463 ( .A1(\SB2_4_26/i0[9] ), .A2(\SB2_4_26/i1_5 ), .A3(
        \SB2_4_26/i0[6] ), .ZN(\SB2_4_26/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U9464 ( .A1(n3863), .A2(\SB1_2_22/Component_Function_1/NAND4_in[1] ), .A3(\SB1_2_22/Component_Function_1/NAND4_in[0] ), .A4(n6058), .ZN(
        \SB1_2_22/buf_output[1] ) );
  NAND3_X2 U9466 ( .A1(\SB2_1_7/i0[10] ), .A2(\SB2_1_7/i1_7 ), .A3(
        \SB2_1_7/i1[9] ), .ZN(n6059) );
  NAND4_X2 U9467 ( .A1(\SB1_1_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_3/Component_Function_3/NAND4_in[1] ), .A3(n6480), .A4(n6060), 
        .ZN(\SB1_1_3/buf_output[3] ) );
  NAND4_X2 U9468 ( .A1(\SB4_25/Component_Function_2/NAND4_in[3] ), .A2(n3716), 
        .A3(n2883), .A4(n6061), .ZN(n6073) );
  NAND3_X1 U9471 ( .A1(\SB4_25/i0_3 ), .A2(n6266), .A3(\SB4_25/i0[8] ), .ZN(
        n6061) );
  NAND4_X2 U9472 ( .A1(\SB2_4_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_17/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_4_17/Component_Function_4/NAND4_in[1] ), .A4(n6062), .ZN(
        \SB2_4_17/buf_output[4] ) );
  NAND3_X1 U9473 ( .A1(\SB2_4_17/i0[10] ), .A2(\SB2_4_17/i0_3 ), .A3(
        \SB2_4_17/i0[9] ), .ZN(n6062) );
  NAND3_X2 U9477 ( .A1(\SB2_2_30/i0[10] ), .A2(\SB2_2_30/i1_5 ), .A3(
        \SB2_2_30/i1[9] ), .ZN(\SB2_2_30/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U9481 ( .A1(\SB3_15/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_15/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_15/Component_Function_0/NAND4_in[1] ), .A4(n6063), .ZN(
        \SB3_15/buf_output[0] ) );
  NAND4_X2 U9483 ( .A1(\SB3_25/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_25/Component_Function_4/NAND4_in[0] ), .A3(n998), .A4(n6064), 
        .ZN(\SB3_25/buf_output[4] ) );
  NAND3_X2 U9485 ( .A1(\SB4_0/i0_4 ), .A2(\SB4_0/i0_3 ), .A3(\SB4_0/i0_0 ), 
        .ZN(n6065) );
  XOR2_X1 U9487 ( .A1(n6066), .A2(n189), .Z(Ciphertext[10]) );
  NAND4_X2 U9488 ( .A1(n1424), .A2(\SB4_30/Component_Function_4/NAND4_in[3] ), 
        .A3(n6202), .A4(\SB4_30/Component_Function_4/NAND4_in[1] ), .ZN(n6066)
         );
  NAND3_X2 U9489 ( .A1(\SB2_2_5/i0[10] ), .A2(\SB2_2_5/i0_3 ), .A3(
        \SB2_2_5/i0[6] ), .ZN(\SB2_2_5/Component_Function_2/NAND4_in[1] ) );
  INV_X1 U9490 ( .I(\SB3_25/buf_output[2] ), .ZN(\SB4_22/i1[9] ) );
  NAND4_X2 U9492 ( .A1(\SB3_25/Component_Function_2/NAND4_in[2] ), .A2(n7254), 
        .A3(\SB3_25/Component_Function_2/NAND4_in[0] ), .A4(
        \SB3_25/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_25/buf_output[2] ) );
  XOR2_X1 U9493 ( .A1(\RI5[0][135] ), .A2(\RI5[0][159] ), .Z(n2440) );
  XOR2_X1 U9496 ( .A1(\RI5[4][90] ), .A2(\RI5[4][126] ), .Z(
        \MC_ARK_ARC_1_4/temp3[24] ) );
  XOR2_X1 U9511 ( .A1(\RI5[0][111] ), .A2(\RI5[0][87] ), .Z(
        \MC_ARK_ARC_1_0/temp2[141] ) );
  NAND3_X2 U9512 ( .A1(\SB2_0_20/i0[10] ), .A2(\SB2_0_20/i1[9] ), .A3(
        \SB2_0_20/i1_7 ), .ZN(\SB2_0_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U9513 ( .A1(\SB1_4_22/i1_5 ), .A2(\SB1_4_22/i0[8] ), .A3(
        \SB1_4_22/i3[0] ), .ZN(n4301) );
  XOR2_X1 U9515 ( .A1(\RI5[2][69] ), .A2(\RI5[2][93] ), .Z(n1018) );
  NAND4_X2 U9522 ( .A1(\SB1_0_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_14/Component_Function_5/NAND4_in[1] ), .A3(n2483), .A4(n6068), 
        .ZN(\SB1_0_14/buf_output[5] ) );
  XOR2_X1 U9525 ( .A1(\SB2_0_19/buf_output[5] ), .A2(\RI5[0][53] ), .Z(n5182)
         );
  NAND4_X2 U9526 ( .A1(\SB2_3_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_5/NAND4_in[0] ), .A4(n6069), .ZN(
        \SB2_3_13/buf_output[5] ) );
  NAND4_X2 U9527 ( .A1(\SB2_3_13/Component_Function_2/NAND4_in[0] ), .A2(n6221), .A3(\SB2_3_13/Component_Function_2/NAND4_in[2] ), .A4(n6070), .ZN(
        \SB2_3_13/buf_output[2] ) );
  NAND4_X2 U9531 ( .A1(\SB1_2_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_13/Component_Function_4/NAND4_in[2] ), .A4(n6071), .ZN(
        \SB1_2_13/buf_output[4] ) );
  NAND3_X1 U9533 ( .A1(\SB1_2_13/i0_4 ), .A2(\SB1_2_13/i1[9] ), .A3(
        \SB1_2_13/i1_5 ), .ZN(n6071) );
  NAND4_X2 U9534 ( .A1(\SB1_3_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_16/Component_Function_5/NAND4_in[0] ), .A4(n1547), .ZN(
        \SB1_3_16/buf_output[5] ) );
  NAND3_X2 U9538 ( .A1(\SB1_3_16/i0_4 ), .A2(\SB1_3_16/i0[6] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[90] ), .ZN(n1547) );
  NAND3_X2 U9542 ( .A1(\SB2_4_19/i0_3 ), .A2(\SB2_4_19/i0[9] ), .A3(
        \SB2_4_19/i0[8] ), .ZN(n4616) );
  NAND4_X2 U9545 ( .A1(\SB2_0_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_23/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_0_23/Component_Function_1/NAND4_in[2] ), .A4(n6072), .ZN(
        \SB2_0_23/buf_output[1] ) );
  NAND4_X2 U9548 ( .A1(\SB4_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_20/Component_Function_3/NAND4_in[2] ), .A3(
        \SB4_20/Component_Function_3/NAND4_in[3] ), .A4(n6574), .ZN(n6997) );
  BUF_X2 U9552 ( .I(\SB3_2/buf_output[2] ), .Z(\SB4_31/i0_0 ) );
  XOR2_X1 U9560 ( .A1(n6073), .A2(n182), .Z(Ciphertext[38]) );
  NAND3_X2 U9564 ( .A1(\SB2_0_19/i0[8] ), .A2(\SB2_0_19/i0[9] ), .A3(
        \RI3[0][77] ), .ZN(\SB2_0_19/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U9566 ( .A1(\RI5[3][107] ), .A2(\RI5[3][179] ), .Z(n6075) );
  NAND4_X2 U9568 ( .A1(n4323), .A2(n3622), .A3(
        \SB1_3_17/Component_Function_1/NAND4_in[3] ), .A4(n4420), .ZN(
        \SB1_3_17/buf_output[1] ) );
  NAND4_X2 U9570 ( .A1(n3505), .A2(\SB1_0_28/Component_Function_4/NAND4_in[2] ), .A3(\SB1_0_28/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_0_28/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB1_0_28/buf_output[4] ) );
  XOR2_X1 U9571 ( .A1(\RI5[4][57] ), .A2(\RI5[4][21] ), .Z(n6076) );
  NAND4_X2 U9572 ( .A1(\SB1_1_27/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_27/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_27/Component_Function_0/NAND4_in[0] ), .A4(n6077), .ZN(
        \SB1_1_27/buf_output[0] ) );
  NAND3_X2 U9575 ( .A1(\SB1_1_27/i0_4 ), .A2(\SB1_1_27/i0[10] ), .A3(
        \SB1_1_27/i0_3 ), .ZN(n6077) );
  NAND4_X2 U9576 ( .A1(\SB2_3_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_14/Component_Function_2/NAND4_in[0] ), .A3(n1716), .A4(n6078), 
        .ZN(\SB2_3_14/buf_output[2] ) );
  XOR2_X1 U9582 ( .A1(n6079), .A2(\MC_ARK_ARC_1_1/temp1[44] ), .Z(n4490) );
  XOR2_X1 U9586 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[182] ), .A2(\RI5[1][14] ), 
        .Z(n6079) );
  XOR2_X1 U9587 ( .A1(\RI5[1][46] ), .A2(\RI5[1][82] ), .Z(n6080) );
  NAND4_X2 U9592 ( .A1(\SB2_0_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_4/NAND4_in[3] ), .A4(n6081), .ZN(
        \SB2_0_28/buf_output[4] ) );
  NAND3_X1 U9593 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i0[10] ), .A3(
        \SB2_0_28/i0[9] ), .ZN(n6081) );
  NAND3_X1 U9594 ( .A1(\SB1_4_22/i1[9] ), .A2(\RI1[4][59] ), .A3(
        \MC_ARK_ARC_1_3/buf_output[58] ), .ZN(n6082) );
  XOR2_X1 U9597 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[89] ), .A2(\RI5[2][83] ), 
        .Z(n6083) );
  NAND4_X2 U9601 ( .A1(\SB1_4_24/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_4_24/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_4_24/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_4_24/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_4_24/buf_output[1] ) );
  NAND4_X2 U9604 ( .A1(\SB1_0_13/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_0_13/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_0_13/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_2/NAND4_in[1] ), .ZN(n1501) );
  NAND3_X2 U9605 ( .A1(\SB1_0_13/i0[6] ), .A2(\SB1_0_13/i0_3 ), .A3(
        \SB1_0_13/i0[10] ), .ZN(\SB1_0_13/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U9610 ( .A1(n6084), .A2(n3491), .Z(\MC_ARK_ARC_1_3/buf_output[37] )
         );
  XOR2_X1 U9613 ( .A1(\MC_ARK_ARC_1_3/temp4[37] ), .A2(
        \MC_ARK_ARC_1_3/temp3[37] ), .Z(n6084) );
  NAND3_X1 U9614 ( .A1(\SB2_2_31/i0[6] ), .A2(\SB2_2_31/i0[8] ), .A3(
        \SB2_2_31/i0[7] ), .ZN(\SB2_2_31/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U9617 ( .A1(\RI5[0][188] ), .A2(\RI5[0][32] ), .Z(
        \MC_ARK_ARC_1_0/temp3[122] ) );
  XOR2_X1 U9618 ( .A1(n6086), .A2(n4), .Z(Ciphertext[74]) );
  NAND4_X2 U9620 ( .A1(\SB4_19/Component_Function_2/NAND4_in[3] ), .A2(n1030), 
        .A3(n7065), .A4(\SB4_19/Component_Function_2/NAND4_in[2] ), .ZN(n6086)
         );
  XOR2_X1 U9629 ( .A1(n2186), .A2(n3037), .Z(n6270) );
  XOR2_X1 U9632 ( .A1(n4031), .A2(n4032), .Z(n3037) );
  NAND3_X2 U9633 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0[10] ), .A3(
        \SB2_3_17/i0[6] ), .ZN(\SB2_3_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U9634 ( .A1(\SB2_3_13/i1_7 ), .A2(n6746), .A3(\SB2_3_13/i0[8] ), 
        .ZN(n6794) );
  XOR2_X1 U9641 ( .A1(\MC_ARK_ARC_1_0/temp1[49] ), .A2(
        \MC_ARK_ARC_1_0/temp2[49] ), .Z(n1161) );
  BUF_X4 U9643 ( .I(\SB1_4_31/buf_output[5] ), .Z(\SB2_4_31/i0_3 ) );
  NAND4_X2 U9650 ( .A1(\SB1_0_16/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_16/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_16/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_0_16/Component_Function_1/NAND4_in[2] ), .ZN(\RI3[0][115] ) );
  XOR2_X1 U9651 ( .A1(\RI5[4][20] ), .A2(\RI5[4][122] ), .Z(n6407) );
  NAND4_X2 U9661 ( .A1(\SB2_4_2/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_4_2/Component_Function_5/NAND4_in[0] ), .A3(n6753), .A4(n6087), 
        .ZN(\SB2_4_2/buf_output[5] ) );
  XOR2_X1 U9667 ( .A1(\MC_ARK_ARC_1_3/temp4[92] ), .A2(n6088), .Z(
        \MC_ARK_ARC_1_3/temp6[92] ) );
  NAND4_X2 U9668 ( .A1(\SB2_3_8/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_3_8/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_8/Component_Function_3/NAND4_in[1] ), .A4(n5437), .ZN(
        \SB2_3_8/buf_output[3] ) );
  INV_X2 U9670 ( .I(\SB1_1_10/buf_output[2] ), .ZN(\SB2_1_7/i1[9] ) );
  NAND4_X2 U9675 ( .A1(\SB1_2_17/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_17/Component_Function_1/NAND4_in[0] ), .A4(n6089), .ZN(
        \SB1_2_17/buf_output[1] ) );
  NAND3_X2 U9679 ( .A1(\SB1_2_17/i0_4 ), .A2(\SB1_2_17/i1_7 ), .A3(
        \SB1_2_17/i0[8] ), .ZN(n6089) );
  XOR2_X1 U9681 ( .A1(n6091), .A2(n6090), .Z(\MC_ARK_ARC_1_4/buf_output[19] )
         );
  XOR2_X1 U9691 ( .A1(\MC_ARK_ARC_1_4/temp3[19] ), .A2(n6157), .Z(n6090) );
  XOR2_X1 U9707 ( .A1(n4666), .A2(\MC_ARK_ARC_1_4/temp4[19] ), .Z(n6091) );
  INV_X2 U9712 ( .I(\RI3[0][152] ), .ZN(\SB2_0_6/i1[9] ) );
  NAND4_X2 U9715 ( .A1(\SB1_0_9/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_9/Component_Function_2/NAND4_in[0] ), .A3(n2432), .A4(
        \SB1_0_9/Component_Function_2/NAND4_in[2] ), .ZN(\RI3[0][152] ) );
  XOR2_X1 U9730 ( .A1(n3751), .A2(n6092), .Z(\MC_ARK_ARC_1_4/temp5[23] ) );
  XOR2_X1 U9732 ( .A1(\RI5[4][161] ), .A2(\RI5[4][185] ), .Z(n6092) );
  NAND3_X2 U9733 ( .A1(\SB1_2_1/i0_0 ), .A2(\SB1_2_1/i0_3 ), .A3(
        \SB1_2_1/i0_4 ), .ZN(n6093) );
  NAND3_X1 U9734 ( .A1(\SB1_4_1/i0_4 ), .A2(\SB1_4_1/i1[9] ), .A3(
        \SB1_4_1/i1_5 ), .ZN(n6094) );
  NAND4_X2 U9736 ( .A1(\SB2_4_8/Component_Function_5/NAND4_in[2] ), .A2(n7412), 
        .A3(n4692), .A4(n6095), .ZN(\SB2_4_8/buf_output[5] ) );
  NAND3_X2 U9751 ( .A1(\SB2_4_8/i0[9] ), .A2(\SB2_4_8/i0[6] ), .A3(n3183), 
        .ZN(n6095) );
  XOR2_X1 U9757 ( .A1(\MC_ARK_ARC_1_4/temp6[129] ), .A2(n6097), .Z(
        \MC_ARK_ARC_1_4/buf_output[129] ) );
  XOR2_X1 U9758 ( .A1(n4266), .A2(n4267), .Z(n6097) );
  NAND3_X2 U9765 ( .A1(\SB1_0_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_6/Component_Function_5/NAND4_in[1] ), .A3(n6098), .ZN(
        \RI3[0][155] ) );
  AOI22_X2 U9772 ( .A1(\SB1_0_6/i0_0 ), .A2(\SB1_0_6/i3[0] ), .B1(
        \SB1_0_6/i0[9] ), .B2(n6099), .ZN(n6098) );
  AND2_X1 U9773 ( .A1(n368), .A2(n246), .Z(n6099) );
  XOR2_X1 U9777 ( .A1(n6100), .A2(n104), .Z(Ciphertext[141]) );
  XOR2_X1 U9779 ( .A1(\MC_ARK_ARC_1_3/temp3[182] ), .A2(n6101), .Z(n3640) );
  XOR2_X1 U9783 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[182] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[176] ), .Z(n6101) );
  INV_X2 U9785 ( .I(\SB1_4_6/buf_output[2] ), .ZN(\SB2_4_3/i1[9] ) );
  NAND4_X2 U9791 ( .A1(n6952), .A2(n6423), .A3(n5079), .A4(n6721), .ZN(
        \SB1_4_6/buf_output[2] ) );
  NAND4_X2 U9793 ( .A1(\SB2_4_26/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_4_26/Component_Function_2/NAND4_in[0] ), .A3(n7151), .A4(n6102), 
        .ZN(\SB2_4_26/buf_output[2] ) );
  NAND4_X2 U9799 ( .A1(\SB3_6/Component_Function_5/NAND4_in[1] ), .A2(n6130), 
        .A3(\SB3_6/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_6/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_6/buf_output[5] )
         );
  XOR2_X1 U9801 ( .A1(\MC_ARK_ARC_1_2/temp2[179] ), .A2(n6103), .Z(n4007) );
  XOR2_X1 U9806 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[89] ), .A2(\RI5[2][53] ), 
        .Z(n6103) );
  NAND4_X2 U9809 ( .A1(\SB1_3_26/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_26/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_3_26/Component_Function_0/NAND4_in[1] ), .A4(n6104), .ZN(
        \SB1_3_26/buf_output[0] ) );
  XOR2_X1 U9811 ( .A1(n1356), .A2(n6105), .Z(\MC_ARK_ARC_1_4/buf_output[29] )
         );
  XOR2_X1 U9812 ( .A1(\MC_ARK_ARC_1_4/temp1[29] ), .A2(
        \MC_ARK_ARC_1_4/temp2[29] ), .Z(n6105) );
  XOR2_X1 U9815 ( .A1(n6106), .A2(n39), .Z(Ciphertext[150]) );
  NAND4_X2 U9819 ( .A1(\SB4_6/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_6/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_6/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_6/Component_Function_0/NAND4_in[2] ), .ZN(n6106) );
  NAND3_X2 U9820 ( .A1(\SB2_1_30/i0[6] ), .A2(\SB2_1_30/i0_3 ), .A3(
        \SB2_1_30/i0[10] ), .ZN(\SB2_1_30/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U9821 ( .A1(n4439), .A2(\MC_ARK_ARC_1_0/temp5[176] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[176] ) );
  XOR2_X1 U9827 ( .A1(\RI5[4][17] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[23] ), 
        .Z(n3751) );
  XOR2_X1 U9829 ( .A1(\RI5[4][179] ), .A2(\RI5[4][143] ), .Z(
        \MC_ARK_ARC_1_4/temp3[77] ) );
  XOR2_X1 U9830 ( .A1(n6148), .A2(n6107), .Z(\RI1[5][155] ) );
  XOR2_X1 U9833 ( .A1(n3088), .A2(\MC_ARK_ARC_1_4/temp4[155] ), .Z(n6107) );
  NAND3_X1 U9835 ( .A1(\SB4_24/i1_7 ), .A2(\SB4_24/i1[9] ), .A3(
        \SB3_26/buf_output[3] ), .ZN(n6108) );
  NAND3_X1 U9836 ( .A1(\SB2_1_30/i0[6] ), .A2(\SB2_1_30/i0[8] ), .A3(
        \SB2_1_30/i0[7] ), .ZN(\SB2_1_30/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U9839 ( .A1(\SB2_4_11/i0_0 ), .A2(\SB2_4_11/i0[10] ), .A3(
        \SB2_4_11/i0[6] ), .ZN(n6828) );
  NAND4_X2 U9840 ( .A1(\SB2_2_17/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_17/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_17/Component_Function_5/NAND4_in[0] ), .A4(n6109), .ZN(
        \SB2_2_17/buf_output[5] ) );
  NAND3_X2 U9846 ( .A1(\RI3[2][88] ), .A2(\SB2_2_17/i0[9] ), .A3(
        \SB2_2_17/i0[6] ), .ZN(n6109) );
  NAND3_X2 U9847 ( .A1(\SB4_6/i0[10] ), .A2(\SB4_6/i0_0 ), .A3(\SB4_6/i0[6] ), 
        .ZN(n7149) );
  XOR2_X1 U9850 ( .A1(\MC_ARK_ARC_1_4/temp5[159] ), .A2(n3148), .Z(
        \MC_ARK_ARC_1_4/buf_output[159] ) );
  NAND4_X2 U9851 ( .A1(\SB2_4_18/Component_Function_1/NAND4_in[1] ), .A2(n2316), .A3(n3765), .A4(\SB2_4_18/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_4_18/buf_output[1] ) );
  NAND4_X2 U9852 ( .A1(n6205), .A2(\SB2_0_15/Component_Function_3/NAND4_in[2] ), .A3(n7181), .A4(\SB2_0_15/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_15/buf_output[3] ) );
  NAND4_X2 U9855 ( .A1(\SB1_2_14/Component_Function_5/NAND4_in[1] ), .A2(n5156), .A3(n6421), .A4(\SB1_2_14/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_14/buf_output[5] ) );
  NAND3_X2 U9856 ( .A1(\SB1_1_4/i0[10] ), .A2(\SB1_1_4/i0[6] ), .A3(
        \SB1_1_4/i0_0 ), .ZN(n798) );
  XOR2_X1 U9858 ( .A1(\RI5[1][106] ), .A2(\RI5[1][100] ), .Z(
        \MC_ARK_ARC_1_1/temp1[106] ) );
  NAND4_X2 U9860 ( .A1(\SB1_1_29/Component_Function_4/NAND4_in[0] ), .A2(n7491), .A3(\SB1_1_29/Component_Function_4/NAND4_in[1] ), .A4(n3747), .ZN(
        \SB1_1_29/buf_output[4] ) );
  NAND4_X2 U9861 ( .A1(\SB2_1_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_28/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_1_28/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_1_28/buf_output[4] ) );
  XOR2_X1 U9862 ( .A1(n7323), .A2(\MC_ARK_ARC_1_1/temp1[82] ), .Z(n1818) );
  XOR2_X1 U9863 ( .A1(\RI5[4][33] ), .A2(\RI5[4][69] ), .Z(
        \MC_ARK_ARC_1_4/temp3[159] ) );
  NAND3_X2 U9867 ( .A1(\SB1_4_28/i0[6] ), .A2(\SB1_4_28/i0_4 ), .A3(
        \SB1_4_28/i0[9] ), .ZN(n6906) );
  XOR2_X1 U9869 ( .A1(\MC_ARK_ARC_1_0/temp1[12] ), .A2(n4207), .Z(
        \MC_ARK_ARC_1_0/temp5[12] ) );
  XOR2_X1 U9870 ( .A1(\RI5[4][28] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[64] ), 
        .Z(\MC_ARK_ARC_1_4/temp3[154] ) );
  NAND4_X2 U9871 ( .A1(\SB2_3_5/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_5/Component_Function_2/NAND4_in[0] ), .A3(n7224), .A4(n6110), 
        .ZN(\SB2_3_5/buf_output[2] ) );
  NAND3_X2 U9875 ( .A1(\SB2_3_5/i0_3 ), .A2(\SB2_3_5/i0[10] ), .A3(
        \SB2_3_5/i0[6] ), .ZN(n6110) );
  NAND3_X2 U9876 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i0[10] ), .A3(\SB3_5/i0[6] ), 
        .ZN(\SB3_5/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U9879 ( .A1(\SB2_4_26/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_26/Component_Function_0/NAND4_in[0] ), .A4(n6111), .ZN(
        \SB2_4_26/buf_output[0] ) );
  NAND3_X2 U9880 ( .A1(\SB2_4_26/i0_0 ), .A2(\SB2_4_26/i0_3 ), .A3(
        \SB2_4_26/i0[7] ), .ZN(n6111) );
  NAND2_X1 U9881 ( .A1(\SB1_2_5/Component_Function_3/NAND4_in[3] ), .A2(n4722), 
        .ZN(n6112) );
  NAND3_X2 U9882 ( .A1(\SB1_2_5/i0[6] ), .A2(\SB1_2_5/i0_3 ), .A3(
        \SB1_2_5/i1[9] ), .ZN(n4722) );
  NAND2_X1 U9883 ( .A1(\SB1_2_5/Component_Function_3/NAND4_in[1] ), .A2(n2041), 
        .ZN(n6113) );
  NAND3_X2 U9887 ( .A1(\SB1_3_31/i0[9] ), .A2(\SB1_3_31/i0_4 ), .A3(
        \SB1_3_31/i0[6] ), .ZN(n4760) );
  NAND3_X2 U9888 ( .A1(\SB2_1_10/i0[10] ), .A2(\SB2_1_10/i1_5 ), .A3(
        \SB2_1_10/i1[9] ), .ZN(\SB2_1_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U9889 ( .A1(\SB2_3_2/i0[6] ), .A2(\SB2_3_2/i0[10] ), .A3(
        \SB2_3_2/i0_3 ), .ZN(n6114) );
  NAND3_X2 U9890 ( .A1(\SB2_4_5/i0[10] ), .A2(\SB2_4_5/i0_3 ), .A3(
        \SB1_4_6/buf_output[4] ), .ZN(
        \SB2_4_5/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U9891 ( .A1(\MC_ARK_ARC_1_1/temp4[93] ), .A2(n6115), .Z(n3115) );
  XOR2_X1 U9892 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[3] ), .A2(\RI5[1][159] ), 
        .Z(n6115) );
  NAND4_X2 U9894 ( .A1(\SB2_3_4/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_4/Component_Function_0/NAND4_in[0] ), .A3(n6117), .A4(n6116), 
        .ZN(\SB2_3_4/buf_output[0] ) );
  NAND4_X2 U9897 ( .A1(\SB2_4_15/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_4_15/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_4_15/Component_Function_3/NAND4_in[0] ), .A4(n6118), .ZN(
        \SB2_4_15/buf_output[3] ) );
  NAND3_X2 U9898 ( .A1(\SB2_4_15/i0_0 ), .A2(\SB2_4_15/i0_3 ), .A3(
        \SB2_4_15/i0_4 ), .ZN(n6118) );
  NAND4_X2 U9902 ( .A1(\SB3_19/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_19/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_19/Component_Function_3/NAND4_in[3] ), .A4(
        \SB3_19/Component_Function_3/NAND4_in[1] ), .ZN(\SB4_17/i0[10] ) );
  NAND4_X2 U9904 ( .A1(\SB1_2_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_25/Component_Function_5/NAND4_in[0] ), .A4(n6119), .ZN(
        \SB1_2_25/buf_output[5] ) );
  NAND3_X2 U9905 ( .A1(\SB1_2_25/i0[6] ), .A2(\SB1_2_25/i0_4 ), .A3(
        \SB1_2_25/i0[9] ), .ZN(n6119) );
  INV_X2 U9908 ( .I(\RI3[0][188] ), .ZN(\SB2_0_0/i1[9] ) );
  XOR2_X1 U9910 ( .A1(n6120), .A2(\MC_ARK_ARC_1_1/temp6[37] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[37] ) );
  XOR2_X1 U9911 ( .A1(\MC_ARK_ARC_1_1/temp1[37] ), .A2(
        \MC_ARK_ARC_1_1/temp2[37] ), .Z(n6120) );
  XOR2_X1 U9915 ( .A1(n5078), .A2(n5077), .Z(\MC_ARK_ARC_1_3/buf_output[91] )
         );
  XOR2_X1 U9918 ( .A1(\MC_ARK_ARC_1_1/temp2[53] ), .A2(n6121), .Z(
        \MC_ARK_ARC_1_1/temp5[53] ) );
  XOR2_X1 U9919 ( .A1(\RI5[1][47] ), .A2(\RI5[1][53] ), .Z(n6121) );
  NAND3_X2 U9924 ( .A1(\SB1_4_18/i0[10] ), .A2(\SB1_4_18/i0_0 ), .A3(
        \SB1_4_18/i0[6] ), .ZN(n6123) );
  NAND3_X2 U9925 ( .A1(\SB2_1_30/i0[6] ), .A2(\SB2_1_30/i0[10] ), .A3(
        \SB2_1_30/i0_0 ), .ZN(n6124) );
  NAND3_X2 U9926 ( .A1(\SB2_1_30/i0[6] ), .A2(\SB2_1_30/i0_4 ), .A3(
        \SB2_1_30/i0[9] ), .ZN(n6125) );
  XOR2_X1 U9928 ( .A1(n3361), .A2(n6126), .Z(n4326) );
  XOR2_X1 U9929 ( .A1(\RI5[3][83] ), .A2(\RI5[3][119] ), .Z(n6126) );
  INV_X1 U9931 ( .I(\SB1_3_28/buf_output[1] ), .ZN(\SB2_3_24/i1_7 ) );
  NAND4_X2 U9932 ( .A1(\SB1_3_28/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_28/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_3_28/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_3_28/Component_Function_1/NAND4_in[1] ), .ZN(
        \SB1_3_28/buf_output[1] ) );
  XOR2_X1 U9934 ( .A1(\RI5[1][41] ), .A2(\RI5[1][47] ), .Z(n6128) );
  NAND4_X1 U9935 ( .A1(\SB4_6/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_6/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_6/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_6/Component_Function_1/NAND4_in[0] ), .ZN(n7147) );
  INV_X2 U9940 ( .I(\SB1_4_1/buf_output[3] ), .ZN(\SB2_4_31/i0[8] ) );
  NAND4_X2 U9941 ( .A1(\SB1_4_1/Component_Function_3/NAND4_in[0] ), .A2(n6238), 
        .A3(\SB1_4_1/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_4_1/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_4_1/buf_output[3] ) );
  NAND4_X2 U9944 ( .A1(n6949), .A2(\SB1_4_7/Component_Function_3/NAND4_in[1] ), 
        .A3(n7537), .A4(n6129), .ZN(\SB1_4_7/buf_output[3] ) );
  NAND3_X2 U9947 ( .A1(\SB3_6/i0[6] ), .A2(\SB3_6/i0_4 ), .A3(\SB3_6/i0[9] ), 
        .ZN(n6130) );
  XOR2_X1 U9951 ( .A1(n7305), .A2(n6131), .Z(\MC_ARK_ARC_1_1/buf_output[115] )
         );
  XOR2_X1 U9957 ( .A1(n3946), .A2(\MC_ARK_ARC_1_1/temp4[115] ), .Z(n6131) );
  INV_X2 U9958 ( .I(\RI3[0][116] ), .ZN(\SB2_0_12/i1[9] ) );
  NAND4_X2 U9963 ( .A1(\SB2_2_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_4/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_4/Component_Function_2/NAND4_in[1] ), .A4(n6132), .ZN(
        \SB2_2_4/buf_output[2] ) );
  NAND3_X2 U9965 ( .A1(\SB2_2_4/i0_0 ), .A2(\SB2_2_4/i0_4 ), .A3(
        \SB2_2_4/i1_5 ), .ZN(n6132) );
  NAND3_X1 U9969 ( .A1(\SB1_1_14/i0_3 ), .A2(\SB1_1_14/i0_0 ), .A3(
        \SB1_1_14/i0[7] ), .ZN(\SB1_1_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U9973 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0_4 ), .A3(\SB4_16/i1_5 ), 
        .ZN(n6133) );
  NAND4_X2 U9975 ( .A1(\SB1_4_20/Component_Function_5/NAND4_in[1] ), .A2(n5111), .A3(n6502), .A4(n6134), .ZN(\SB1_4_20/buf_output[5] ) );
  XOR2_X1 U9976 ( .A1(\RI5[4][19] ), .A2(\RI5[4][13] ), .Z(n4666) );
  NAND4_X2 U9978 ( .A1(\SB2_3_30/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_30/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_30/Component_Function_2/NAND4_in[1] ), .A4(n6135), .ZN(
        \SB2_3_30/buf_output[2] ) );
  NAND4_X2 U9980 ( .A1(\SB2_0_3/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_3/Component_Function_3/NAND4_in[0] ), .A3(n6184), .A4(n4465), 
        .ZN(\SB2_0_3/buf_output[3] ) );
  XOR2_X1 U9981 ( .A1(n6136), .A2(n169), .Z(Ciphertext[27]) );
  NAND4_X2 U9982 ( .A1(n5204), .A2(\SB4_27/Component_Function_3/NAND4_in[1] ), 
        .A3(\SB4_27/Component_Function_3/NAND4_in[3] ), .A4(
        \SB4_27/Component_Function_3/NAND4_in[2] ), .ZN(n6136) );
  NAND4_X2 U9983 ( .A1(\SB2_4_21/Component_Function_5/NAND4_in[1] ), .A2(n6137), .A3(\SB2_4_21/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_4_21/Component_Function_5/NAND4_in[2] ), .ZN(
        \SB2_4_21/buf_output[5] ) );
  XOR2_X1 U9990 ( .A1(\RI5[4][61] ), .A2(\RI5[4][85] ), .Z(
        \MC_ARK_ARC_1_4/temp2[115] ) );
  XOR2_X1 U9991 ( .A1(n7436), .A2(\MC_ARK_ARC_1_4/temp2[91] ), .Z(
        \MC_ARK_ARC_1_4/temp5[91] ) );
  XOR2_X1 U9995 ( .A1(n6138), .A2(n140), .Z(Ciphertext[20]) );
  NAND4_X2 U9996 ( .A1(n2015), .A2(n5304), .A3(n6751), .A4(
        \SB4_28/Component_Function_2/NAND4_in[2] ), .ZN(n6138) );
  INV_X4 U9997 ( .I(\SB2_2_4/i0[7] ), .ZN(\SB2_2_4/i0_4 ) );
  NAND3_X1 U10003 ( .A1(\SB2_2_4/i0_0 ), .A2(\SB2_2_4/i0_3 ), .A3(
        \SB2_2_4/i0[7] ), .ZN(n1600) );
  NOR2_X2 U10004 ( .A1(n5015), .A2(n4642), .ZN(\SB2_2_4/i0[7] ) );
  BUF_X4 U10005 ( .I(\SB3_28/buf_output[5] ), .Z(\SB4_28/i0_3 ) );
  NAND3_X2 U10010 ( .A1(n3991), .A2(n3994), .A3(\SB2_2_3/i3[0] ), .ZN(
        \SB2_2_3/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U10011 ( .A1(n6139), .A2(n1165), .Z(\MC_ARK_ARC_1_2/temp5[154] ) );
  XOR2_X1 U10012 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[124] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[100] ), .Z(n6139) );
  INV_X2 U10013 ( .I(\SB1_2_27/buf_output[3] ), .ZN(\SB2_2_25/i0[8] ) );
  NAND4_X2 U10014 ( .A1(\SB1_2_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_27/Component_Function_3/NAND4_in[2] ), .A4(n6187), .ZN(
        \SB1_2_27/buf_output[3] ) );
  NAND3_X1 U10015 ( .A1(\SB2_0_25/i0_0 ), .A2(\SB2_0_25/i0[9] ), .A3(
        \SB2_0_25/i0[8] ), .ZN(\SB2_0_25/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U10016 ( .A1(\SB1_2_21/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_2_21/Component_Function_2/NAND4_in[1] ), .A3(n6338), .A4(n6140), 
        .ZN(\SB1_2_21/buf_output[2] ) );
  NAND3_X1 U10017 ( .A1(\SB1_2_21/i0[10] ), .A2(\SB1_2_21/i1_5 ), .A3(
        \SB1_2_21/i1[9] ), .ZN(n6140) );
  XOR2_X1 U10018 ( .A1(n6141), .A2(n6669), .Z(n2375) );
  XOR2_X1 U10019 ( .A1(\RI5[1][128] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[152] ), .Z(n6141) );
  INV_X2 U10021 ( .I(\SB1_3_8/buf_output[2] ), .ZN(\SB2_3_5/i1[9] ) );
  XOR2_X1 U10025 ( .A1(n6142), .A2(n109), .Z(Ciphertext[93]) );
  NAND4_X2 U10027 ( .A1(\SB4_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_16/Component_Function_3/NAND4_in[3] ), .A3(n6912), .A4(n1453), 
        .ZN(n6142) );
  XOR2_X1 U10032 ( .A1(\MC_ARK_ARC_1_0/temp6[100] ), .A2(n6143), .Z(
        \MC_ARK_ARC_1_0/buf_output[100] ) );
  XOR2_X1 U10039 ( .A1(\MC_ARK_ARC_1_0/temp2[100] ), .A2(
        \MC_ARK_ARC_1_0/temp1[100] ), .Z(n6143) );
  NAND3_X2 U10040 ( .A1(\SB2_0_24/i0[6] ), .A2(\SB2_0_24/i0_0 ), .A3(
        \SB2_0_24/i0[10] ), .ZN(n6144) );
  NAND4_X2 U10042 ( .A1(\SB1_3_31/Component_Function_0/NAND4_in[1] ), .A2(
        n4842), .A3(\SB1_3_31/Component_Function_0/NAND4_in[2] ), .A4(n6145), 
        .ZN(\SB1_3_31/buf_output[0] ) );
  NAND2_X1 U10047 ( .A1(\SB1_3_31/i0[9] ), .A2(\SB1_3_31/i0[10] ), .ZN(n6145)
         );
  XOR2_X1 U10050 ( .A1(\MC_ARK_ARC_1_3/temp5[115] ), .A2(n6146), .Z(
        \MC_ARK_ARC_1_3/buf_output[115] ) );
  XOR2_X1 U10051 ( .A1(\MC_ARK_ARC_1_3/temp3[115] ), .A2(
        \MC_ARK_ARC_1_3/temp4[115] ), .Z(n6146) );
  NAND4_X2 U10055 ( .A1(\SB2_4_0/Component_Function_5/NAND4_in[2] ), .A2(n7108), .A3(n1262), .A4(n6147), .ZN(\SB2_4_0/buf_output[5] ) );
  NAND2_X2 U10056 ( .A1(\SB2_4_0/i0_0 ), .A2(\SB2_4_0/i3[0] ), .ZN(n6147) );
  BUF_X4 U10057 ( .I(\MC_ARK_ARC_1_0/buf_output[173] ), .Z(\SB1_1_3/i0_3 ) );
  XOR2_X1 U10060 ( .A1(\RI5[3][10] ), .A2(\RI5[3][40] ), .Z(n4767) );
  NAND3_X1 U10065 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i1[9] ), .A3(
        \SB2_3_31/i0[6] ), .ZN(\SB2_3_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10066 ( .A1(\SB1_0_16/i0[9] ), .A2(\SB1_0_16/i0[6] ), .A3(
        \SB1_0_16/i1_5 ), .ZN(\SB1_0_16/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U10068 ( .A1(n2442), .A2(\MC_ARK_ARC_1_4/temp3[155] ), .Z(n6148) );
  BUF_X2 U10071 ( .I(n283), .Z(n6149) );
  XOR2_X1 U10072 ( .A1(n6150), .A2(n122), .Z(Ciphertext[166]) );
  NAND4_X2 U10073 ( .A1(\SB4_4/Component_Function_4/NAND4_in[3] ), .A2(n3882), 
        .A3(\SB4_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB4_4/Component_Function_4/NAND4_in[1] ), .ZN(n6150) );
  NAND3_X2 U10076 ( .A1(\SB2_4_21/i0[6] ), .A2(\SB2_4_21/i0_0 ), .A3(
        \SB2_4_21/i0[10] ), .ZN(\SB2_4_21/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X2 U10077 ( .A1(\SB1_3_0/i0_3 ), .A2(\SB1_3_0/i0_4 ), .A3(
        \SB1_3_0/i1[9] ), .ZN(\SB1_3_0/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U10078 ( .A1(\SB2_1_8/i0_3 ), .A2(\SB2_1_8/i0[8] ), .A3(
        \SB2_1_8/i0[9] ), .ZN(\SB2_1_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U10080 ( .A1(\SB2_2_18/i0[10] ), .A2(\SB2_2_18/i1_7 ), .A3(
        \SB2_2_18/i1[9] ), .ZN(\SB2_2_18/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U10081 ( .A1(\SB2_2_5/buf_output[1] ), .A2(\RI5[2][187] ), .Z(n4705)
         );
  XOR2_X1 U10085 ( .A1(\RI5[1][65] ), .A2(\RI5[1][59] ), .Z(
        \MC_ARK_ARC_1_1/temp1[65] ) );
  NAND3_X2 U10089 ( .A1(\SB1_3_23/i0_4 ), .A2(\SB1_3_23/i0[6] ), .A3(
        \SB1_3_23/i0[9] ), .ZN(n4433) );
  NAND3_X2 U10090 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i1_7 ), .A3(
        \SB2_1_20/i1[9] ), .ZN(n4276) );
  XOR2_X1 U10091 ( .A1(\RI5[1][5] ), .A2(\RI5[1][173] ), .Z(n6151) );
  XOR2_X1 U10092 ( .A1(\MC_ARK_ARC_1_2/temp6[52] ), .A2(
        \MC_ARK_ARC_1_2/temp5[52] ), .Z(\MC_ARK_ARC_1_2/buf_output[52] ) );
  NAND3_X2 U10093 ( .A1(\SB2_4_10/i0[10] ), .A2(\SB2_4_10/i1[9] ), .A3(n6269), 
        .ZN(n6308) );
  XOR2_X1 U10095 ( .A1(\MC_ARK_ARC_1_1/temp5[135] ), .A2(
        \MC_ARK_ARC_1_1/temp6[135] ), .Z(\MC_ARK_ARC_1_1/buf_output[135] ) );
  NAND4_X2 U10097 ( .A1(\SB1_3_19/Component_Function_5/NAND4_in[3] ), .A2(
        n2502), .A3(\SB1_3_19/Component_Function_5/NAND4_in[0] ), .A4(n6152), 
        .ZN(\SB1_3_19/buf_output[5] ) );
  NAND3_X2 U10099 ( .A1(\SB1_3_19/i0[10] ), .A2(\SB1_3_19/i0_0 ), .A3(
        \SB1_3_19/i0[6] ), .ZN(n6152) );
  INV_X2 U10100 ( .I(\SB1_2_21/buf_output[2] ), .ZN(\SB2_2_18/i1[9] ) );
  NAND4_X2 U10105 ( .A1(n4536), .A2(\SB2_2_7/Component_Function_2/NAND4_in[0] ), .A3(n6843), .A4(n6153), .ZN(\SB2_2_7/buf_output[2] ) );
  NAND3_X2 U10106 ( .A1(\SB2_2_7/i0[10] ), .A2(\SB2_2_7/i0_3 ), .A3(
        \SB2_2_7/i0[6] ), .ZN(n6153) );
  BUF_X4 U10107 ( .I(\SB2_4_19/buf_output[2] ), .Z(\RI5[4][92] ) );
  XOR2_X1 U10108 ( .A1(\SB2_4_7/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[3] ), .Z(n1049) );
  XOR2_X1 U10113 ( .A1(\MC_ARK_ARC_1_3/temp1[185] ), .A2(n6154), .Z(n5082) );
  XOR2_X1 U10117 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), .A2(\RI5[3][131] ), .Z(n6154) );
  NAND3_X2 U10123 ( .A1(\SB2_4_27/i1[9] ), .A2(\SB2_4_27/i0_3 ), .A3(
        \SB2_4_27/i0[6] ), .ZN(\SB2_4_27/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U10128 ( .A1(n6155), .A2(n190), .Z(Ciphertext[103]) );
  NAND4_X2 U10131 ( .A1(\SB4_14/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_14/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_14/Component_Function_1/NAND4_in[2] ), .ZN(n6155) );
  INV_X1 U10132 ( .I(\SB3_16/buf_output[3] ), .ZN(\SB4_14/i0[8] ) );
  NAND4_X2 U10133 ( .A1(n4713), .A2(\SB3_16/Component_Function_3/NAND4_in[1] ), 
        .A3(n4773), .A4(\SB3_16/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB3_16/buf_output[3] ) );
  XOR2_X1 U10136 ( .A1(\MC_ARK_ARC_1_4/temp6[9] ), .A2(n6156), .Z(
        \MC_ARK_ARC_1_4/buf_output[9] ) );
  XOR2_X1 U10137 ( .A1(\MC_ARK_ARC_1_4/temp2[9] ), .A2(
        \MC_ARK_ARC_1_4/temp1[9] ), .Z(n6156) );
  NAND3_X1 U10139 ( .A1(\SB2_3_7/i0_4 ), .A2(\SB2_3_7/i1[9] ), .A3(
        \SB2_3_7/i1_5 ), .ZN(\SB2_3_7/Component_Function_4/NAND4_in[3] ) );
  INV_X2 U10144 ( .I(\SB1_4_7/buf_output[3] ), .ZN(\SB2_4_5/i0[8] ) );
  XOR2_X1 U10148 ( .A1(\RI5[4][181] ), .A2(\SB2_4_9/buf_output[1] ), .Z(n6157)
         );
  NAND3_X2 U10151 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i0[9] ), .A3(
        \SB2_2_17/i0[8] ), .ZN(n4029) );
  INV_X2 U10153 ( .I(\SB1_1_4/buf_output[3] ), .ZN(\SB2_1_2/i0[8] ) );
  NAND4_X2 U10155 ( .A1(\SB1_1_4/Component_Function_3/NAND4_in[1] ), .A2(n3487), .A3(\SB1_1_4/Component_Function_3/NAND4_in[0] ), .A4(n1693), .ZN(
        \SB1_1_4/buf_output[3] ) );
  NAND4_X2 U10161 ( .A1(\SB2_4_12/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_4_12/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_4_12/Component_Function_0/NAND4_in[2] ), .A4(n6158), .ZN(
        \SB2_4_12/buf_output[0] ) );
  NAND3_X2 U10167 ( .A1(\SB2_4_12/i0[7] ), .A2(\SB2_4_12/i0[6] ), .A3(
        \SB2_4_12/i0[8] ), .ZN(n6158) );
  NAND3_X2 U10168 ( .A1(\SB2_2_23/i0_0 ), .A2(\SB2_2_23/i0[10] ), .A3(
        \SB2_2_23/i0[6] ), .ZN(n6159) );
  NAND4_X2 U10169 ( .A1(\SB1_4_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_4_1/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_4_1/Component_Function_2/NAND4_in[3] ), .A4(n6160), .ZN(
        \SB1_4_1/buf_output[2] ) );
  XOR2_X1 U10173 ( .A1(n6161), .A2(n6594), .Z(\MC_ARK_ARC_1_3/temp5[39] ) );
  XOR2_X1 U10174 ( .A1(\RI5[3][33] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[39] ), 
        .Z(n6161) );
  XOR2_X1 U10175 ( .A1(\RI5[0][116] ), .A2(\RI5[0][20] ), .Z(n6499) );
  XOR2_X1 U10176 ( .A1(n6162), .A2(\MC_ARK_ARC_1_4/temp4[23] ), .Z(
        \MC_ARK_ARC_1_4/temp6[23] ) );
  XOR2_X1 U10178 ( .A1(\RI5[4][89] ), .A2(\RI5[4][125] ), .Z(n6162) );
  NAND4_X2 U10184 ( .A1(n2972), .A2(
        \SB2_3_29/Component_Function_3/NAND4_in[3] ), .A3(n6700), .A4(n6163), 
        .ZN(\SB2_3_29/buf_output[3] ) );
  NAND4_X2 U10185 ( .A1(\SB3_13/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_13/Component_Function_2/NAND4_in[0] ), .A3(n7064), .A4(n6164), 
        .ZN(\RI3[5][128] ) );
  NAND3_X2 U10186 ( .A1(\SB3_13/i0[9] ), .A2(\SB3_13/i0[8] ), .A3(
        \RI1[5][113] ), .ZN(n6164) );
  NAND2_X1 U10187 ( .A1(\SB1_4_6/i0[9] ), .A2(\SB1_4_6/i0[10] ), .ZN(
        \SB1_4_6/Component_Function_0/NAND4_in[0] ) );
  XOR2_X1 U10188 ( .A1(\RI5[0][103] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[139] ), .Z(\MC_ARK_ARC_1_0/temp3[37] ) );
  INV_X2 U10190 ( .I(\SB1_3_13/buf_output[2] ), .ZN(\SB2_3_10/i1[9] ) );
  NAND4_X2 U10191 ( .A1(\SB1_3_13/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_13/Component_Function_2/NAND4_in[2] ), .A3(n4634), .A4(n4808), 
        .ZN(\SB1_3_13/buf_output[2] ) );
  XOR2_X1 U10192 ( .A1(n940), .A2(n6165), .Z(\MC_ARK_ARC_1_2/buf_output[111] )
         );
  XOR2_X1 U10193 ( .A1(\MC_ARK_ARC_1_2/temp2[111] ), .A2(
        \MC_ARK_ARC_1_2/temp1[111] ), .Z(n6165) );
  NAND3_X2 U10195 ( .A1(n6686), .A2(\SB2_2_26/i0_3 ), .A3(\SB2_2_26/i0[10] ), 
        .ZN(n6602) );
  INV_X1 U10196 ( .I(\SB1_1_28/buf_output[1] ), .ZN(\SB2_1_24/i1_7 ) );
  NAND4_X2 U10197 ( .A1(\SB1_1_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_28/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_1_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_28/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_28/buf_output[1] ) );
  XOR2_X1 U10198 ( .A1(\MC_ARK_ARC_1_1/temp5[131] ), .A2(n6166), .Z(
        \MC_ARK_ARC_1_1/buf_output[131] ) );
  XOR2_X1 U10199 ( .A1(\MC_ARK_ARC_1_1/temp3[131] ), .A2(
        \MC_ARK_ARC_1_1/temp4[131] ), .Z(n6166) );
  NAND3_X1 U10200 ( .A1(\SB1_4_16/i0_3 ), .A2(\SB1_4_16/i0[9] ), .A3(
        \SB1_4_16/i0[10] ), .ZN(\SB1_4_16/Component_Function_4/NAND4_in[2] )
         );
  NAND4_X2 U10208 ( .A1(n4421), .A2(
        \SB2_3_28/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_28/Component_Function_5/NAND4_in[1] ), .A4(n6167), .ZN(
        \SB2_3_28/buf_output[5] ) );
  XOR2_X1 U10209 ( .A1(\MC_ARK_ARC_1_2/temp3[3] ), .A2(
        \MC_ARK_ARC_1_2/temp4[3] ), .Z(\MC_ARK_ARC_1_2/temp6[3] ) );
  NAND4_X2 U10211 ( .A1(\SB1_1_25/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_25/Component_Function_5/NAND4_in[2] ), .A3(n5383), .A4(n6168), 
        .ZN(\SB1_1_25/buf_output[5] ) );
  NAND3_X2 U10212 ( .A1(\SB1_1_25/i0[6] ), .A2(\SB1_1_25/i0[9] ), .A3(
        \SB1_1_25/i0_4 ), .ZN(n6168) );
  NAND4_X2 U10215 ( .A1(\SB2_4_16/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_4_16/Component_Function_4/NAND4_in[0] ), .A3(n7388), .A4(n6169), 
        .ZN(\SB2_4_16/buf_output[4] ) );
  NAND3_X1 U10217 ( .A1(\SB2_4_16/i0_0 ), .A2(\SB2_4_16/i1_7 ), .A3(
        \SB2_4_16/i3[0] ), .ZN(n6169) );
  NAND3_X2 U10218 ( .A1(\SB2_3_20/i0[6] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \SB2_3_20/i1[9] ), .ZN(\SB2_3_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U10224 ( .A1(\SB1_4_22/i0[6] ), .A2(\SB1_4_22/i0_4 ), .A3(
        \SB1_4_22/i0[9] ), .ZN(\SB1_4_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U10226 ( .A1(n1494), .A2(\SB4_24/i1_5 ), .A3(\SB4_24/i3[0] ), .ZN(
        \SB4_24/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U10228 ( .A1(n6170), .A2(\MC_ARK_ARC_1_4/temp1[133] ), .Z(
        \MC_ARK_ARC_1_4/temp5[133] ) );
  XOR2_X1 U10229 ( .A1(\RI5[4][79] ), .A2(\RI5[4][103] ), .Z(n6170) );
  NAND3_X1 U10230 ( .A1(\SB4_30/i0[9] ), .A2(\SB4_30/i0_3 ), .A3(
        \SB4_30/i0[8] ), .ZN(n6171) );
  NAND4_X2 U10238 ( .A1(n2630), .A2(
        \SB2_1_21/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_1_21/Component_Function_5/NAND4_in[0] ), .A4(n6172), .ZN(
        \SB2_1_21/buf_output[5] ) );
  NAND3_X2 U10239 ( .A1(\SB2_1_21/i0[6] ), .A2(\SB2_1_21/i0_0 ), .A3(
        \SB2_1_21/i0[10] ), .ZN(n6172) );
  NAND4_X2 U10240 ( .A1(\SB2_4_22/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_4_22/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_4_22/Component_Function_1/NAND4_in[0] ), .A4(n6173), .ZN(
        \SB2_4_22/buf_output[1] ) );
  NAND3_X1 U10244 ( .A1(\SB2_4_22/i0[9] ), .A2(\SB2_4_22/i0[6] ), .A3(
        \SB2_4_22/i1_5 ), .ZN(n6173) );
  NAND4_X2 U10247 ( .A1(\SB2_3_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_17/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_17/Component_Function_4/NAND4_in[1] ), .A4(n6174), .ZN(
        \SB2_3_17/buf_output[4] ) );
  NAND4_X2 U10250 ( .A1(n3127), .A2(
        \SB1_2_31/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_2_31/Component_Function_3/NAND4_in[1] ), .A4(n6175), .ZN(
        \SB1_2_31/buf_output[3] ) );
  NAND3_X1 U10252 ( .A1(\SB1_2_31/i0[8] ), .A2(\SB1_2_31/i3[0] ), .A3(
        \SB1_2_31/i1_5 ), .ZN(n6175) );
  NAND3_X2 U10255 ( .A1(\SB2_3_6/i0_3 ), .A2(\SB2_3_6/i0[8] ), .A3(
        \SB2_3_6/i1_7 ), .ZN(\SB2_3_6/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U10256 ( .A1(\MC_ARK_ARC_1_0/temp6[87] ), .A2(n6176), .Z(
        \MC_ARK_ARC_1_0/buf_output[87] ) );
  NAND4_X2 U10259 ( .A1(\SB2_2_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_29/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_2_29/Component_Function_3/NAND4_in[1] ), .A4(n6177), .ZN(
        \SB2_2_29/buf_output[3] ) );
  XOR2_X1 U10260 ( .A1(\MC_ARK_ARC_1_1/temp4[3] ), .A2(n6178), .Z(
        \MC_ARK_ARC_1_1/temp6[3] ) );
  XOR2_X1 U10262 ( .A1(\RI5[1][69] ), .A2(\RI5[1][105] ), .Z(n6178) );
  BUF_X2 U10268 ( .I(\MC_ARK_ARC_1_4/buf_output[78] ), .Z(\SB3_18/i0[9] ) );
  NAND3_X1 U10269 ( .A1(\SB3_16/i0_4 ), .A2(\SB3_16/i0_0 ), .A3(\SB3_16/i1_5 ), 
        .ZN(n6179) );
  XOR2_X1 U10270 ( .A1(\MC_ARK_ARC_1_0/temp6[82] ), .A2(n6180), .Z(
        \MC_ARK_ARC_1_0/buf_output[82] ) );
  XOR2_X1 U10274 ( .A1(\MC_ARK_ARC_1_0/temp2[82] ), .A2(
        \MC_ARK_ARC_1_0/temp1[82] ), .Z(n6180) );
  NAND3_X2 U10276 ( .A1(\SB3_6/i1_5 ), .A2(\SB3_6/i1[9] ), .A3(\SB3_6/i0_4 ), 
        .ZN(n7385) );
  NAND4_X2 U10279 ( .A1(\SB1_2_20/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_20/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_5/NAND4_in[0] ), .A4(n6181), .ZN(
        \SB1_2_20/buf_output[5] ) );
  NAND3_X2 U10287 ( .A1(\SB1_2_20/i0[9] ), .A2(\SB1_2_20/i0_4 ), .A3(
        \SB1_2_20/i0[6] ), .ZN(n6181) );
  NAND4_X2 U10288 ( .A1(\SB2_4_24/Component_Function_5/NAND4_in[2] ), .A2(n686), .A3(\SB2_4_24/Component_Function_5/NAND4_in[0] ), .A4(n6182), .ZN(
        \SB2_4_24/buf_output[5] ) );
  NAND3_X2 U10289 ( .A1(\SB2_4_24/i0_4 ), .A2(\SB2_4_24/i0[9] ), .A3(
        \SB2_4_24/i0[6] ), .ZN(n6182) );
  XOR2_X1 U10290 ( .A1(\RI5[3][6] ), .A2(\RI5[3][42] ), .Z(n1179) );
  XOR2_X1 U10291 ( .A1(\MC_ARK_ARC_1_4/temp1[153] ), .A2(
        \MC_ARK_ARC_1_4/temp2[153] ), .Z(n1656) );
  NAND3_X2 U10294 ( .A1(\SB1_2_25/i1[9] ), .A2(\SB1_2_25/i0_3 ), .A3(
        \SB1_2_25/i0[6] ), .ZN(\SB1_2_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U10295 ( .A1(\SB4_3/i0_0 ), .A2(\SB4_3/i0[8] ), .A3(\SB4_3/i0[9] ), 
        .ZN(\SB4_3/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U10296 ( .A1(\RI5[3][51] ), .A2(\RI5[3][117] ), .Z(n7113) );
  XOR2_X1 U10297 ( .A1(\RI5[0][29] ), .A2(\RI5[0][185] ), .Z(
        \MC_ARK_ARC_1_0/temp3[119] ) );
  XOR2_X1 U10298 ( .A1(n6731), .A2(\MC_ARK_ARC_1_3/temp6[113] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[113] ) );
  XOR2_X1 U10299 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[164] ), .A2(\RI5[2][8] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[98] ) );
  NAND4_X2 U10303 ( .A1(\SB1_4_23/Component_Function_5/NAND4_in[1] ), .A2(
        n3242), .A3(\SB1_4_23/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_4_23/Component_Function_5/NAND4_in[2] ), .ZN(
        \SB1_4_23/buf_output[5] ) );
  XOR2_X1 U10305 ( .A1(\RI5[3][9] ), .A2(\RI5[3][3] ), .Z(
        \MC_ARK_ARC_1_3/temp1[9] ) );
  XOR2_X1 U10306 ( .A1(\MC_ARK_ARC_1_2/temp5[187] ), .A2(n6183), .Z(
        \MC_ARK_ARC_1_2/buf_output[187] ) );
  XOR2_X1 U10307 ( .A1(\MC_ARK_ARC_1_2/temp3[187] ), .A2(
        \MC_ARK_ARC_1_2/temp4[187] ), .Z(n6183) );
  NAND3_X2 U10308 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0_0 ), .A3(
        \SB2_3_0/i0_4 ), .ZN(\SB2_3_0/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U10309 ( .A1(\MC_ARK_ARC_1_0/temp6[119] ), .A2(
        \MC_ARK_ARC_1_0/temp5[119] ), .Z(\MC_ARK_ARC_1_0/buf_output[119] ) );
  NAND4_X2 U10312 ( .A1(\SB1_4_29/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_29/Component_Function_0/NAND4_in[0] ), .A4(n2787), .ZN(
        \SB1_4_29/buf_output[0] ) );
  NAND4_X2 U10318 ( .A1(\SB2_0_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_26/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_0_26/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_26/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_26/buf_output[2] ) );
  NAND3_X1 U10319 ( .A1(\SB2_0_3/i0_3 ), .A2(\SB2_0_3/i0_0 ), .A3(
        \RI3[0][172] ), .ZN(n6184) );
  XOR2_X1 U10320 ( .A1(\RI5[0][133] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[139] ), .Z(\MC_ARK_ARC_1_0/temp1[139] ) );
  NAND3_X2 U10321 ( .A1(\SB3_6/i1_5 ), .A2(\SB3_6/i0[8] ), .A3(\SB3_6/i3[0] ), 
        .ZN(\SB3_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U10323 ( .A1(\SB1_0_30/i0[6] ), .A2(\SB1_0_30/i0_4 ), .A3(
        \SB1_0_30/i0[9] ), .ZN(n6185) );
  NAND4_X2 U10325 ( .A1(\SB2_2_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_25/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_25/Component_Function_1/NAND4_in[0] ), .A4(n6186), .ZN(
        \SB2_2_25/buf_output[1] ) );
  NAND4_X2 U10326 ( .A1(n1295), .A2(\SB4_4/Component_Function_2/NAND4_in[2] ), 
        .A3(n3780), .A4(n6188), .ZN(n6189) );
  XOR2_X1 U10329 ( .A1(n6189), .A2(n22), .Z(Ciphertext[164]) );
  XOR2_X1 U10330 ( .A1(\MC_ARK_ARC_1_4/temp5[133] ), .A2(
        \MC_ARK_ARC_1_4/temp6[133] ), .Z(\MC_ARK_ARC_1_4/buf_output[133] ) );
  XOR2_X1 U10332 ( .A1(n6190), .A2(n160), .Z(Ciphertext[119]) );
  NAND4_X2 U10333 ( .A1(\SB1_3_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_29/Component_Function_2/NAND4_in[2] ), .A4(n756), .ZN(
        \SB1_3_29/buf_output[2] ) );
  NAND3_X2 U10334 ( .A1(\SB2_3_26/i0_4 ), .A2(\SB2_3_26/i0_3 ), .A3(
        \SB2_3_26/i1[9] ), .ZN(\SB2_3_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U10336 ( .A1(\SB1_0_5/i0[6] ), .A2(\SB1_0_5/i0_3 ), .A3(
        \SB1_0_5/i1[9] ), .ZN(\SB1_0_5/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 U10341 ( .A1(n2398), .A2(n6191), .ZN(\SB2_1_2/i0_4 ) );
  AND2_X1 U10342 ( .A1(n4640), .A2(\SB1_1_3/Component_Function_4/NAND4_in[1] ), 
        .Z(n6191) );
  XOR2_X1 U10343 ( .A1(n6193), .A2(n6192), .Z(n6198) );
  XOR2_X1 U10347 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[32] ), .A2(n474), .Z(
        n6192) );
  XOR2_X1 U10348 ( .A1(\RI5[3][38] ), .A2(\RI5[3][74] ), .Z(n6193) );
  INV_X2 U10351 ( .I(\SB1_2_30/buf_output[2] ), .ZN(\SB2_2_27/i1[9] ) );
  NAND4_X2 U10354 ( .A1(n936), .A2(n4944), .A3(n4129), .A4(n3963), .ZN(
        \SB1_2_30/buf_output[2] ) );
  INV_X2 U10355 ( .I(\MC_ARK_ARC_1_0/buf_output[173] ), .ZN(\SB1_1_3/i1_5 ) );
  INV_X1 U10358 ( .I(n2287), .ZN(\SB2_3_8/i1_5 ) );
  NAND4_X2 U10360 ( .A1(n1271), .A2(\SB1_3_8/Component_Function_5/NAND4_in[1] ), .A3(n2306), .A4(n4392), .ZN(n2287) );
  NAND3_X2 U10361 ( .A1(\SB2_4_25/i0_3 ), .A2(\SB2_4_25/i1_7 ), .A3(
        \SB2_4_25/i0[8] ), .ZN(\SB2_4_25/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U10362 ( .A1(\MC_ARK_ARC_1_3/temp6[190] ), .A2(n6194), .Z(
        \MC_ARK_ARC_1_3/buf_output[190] ) );
  XOR2_X1 U10363 ( .A1(\MC_ARK_ARC_1_3/temp2[190] ), .A2(
        \MC_ARK_ARC_1_3/temp1[190] ), .Z(n6194) );
  NAND4_X2 U10364 ( .A1(n1415), .A2(
        \SB2_2_30/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_30/Component_Function_5/NAND4_in[0] ), .A4(n6195), .ZN(
        \SB2_2_30/buf_output[5] ) );
  NAND3_X2 U10366 ( .A1(\SB2_2_30/i0_0 ), .A2(\SB2_2_30/i0[10] ), .A3(
        \SB2_2_30/i0[6] ), .ZN(n6195) );
  XOR2_X1 U10368 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[179] ), .A2(\RI5[2][11] ), 
        .Z(n6252) );
  XOR2_X1 U10369 ( .A1(\MC_ARK_ARC_1_4/temp5[22] ), .A2(n6196), .Z(
        \MC_ARK_ARC_1_4/buf_output[22] ) );
  XOR2_X1 U10371 ( .A1(\MC_ARK_ARC_1_4/temp3[22] ), .A2(
        \MC_ARK_ARC_1_4/temp4[22] ), .Z(n6196) );
  NAND3_X2 U10372 ( .A1(n851), .A2(\SB2_3_10/i1_5 ), .A3(\SB2_3_10/i0_0 ), 
        .ZN(n7418) );
  BUF_X4 U10374 ( .I(\SB2_3_10/buf_output[2] ), .Z(\RI5[3][146] ) );
  NAND4_X2 U10376 ( .A1(\SB1_4_4/Component_Function_5/NAND4_in[1] ), .A2(n6872), .A3(\SB1_4_4/Component_Function_5/NAND4_in[0] ), .A4(n2056), .ZN(
        \SB1_4_4/buf_output[5] ) );
  XOR2_X1 U10378 ( .A1(\MC_ARK_ARC_1_2/temp6[109] ), .A2(n6420), .Z(
        \MC_ARK_ARC_1_2/buf_output[109] ) );
  NAND3_X2 U10381 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0_4 ), .A3(
        \SB1_1_22/i1[9] ), .ZN(\SB1_1_22/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U10382 ( .A1(n6198), .A2(n6197), .Z(\MC_ARK_ARC_1_3/buf_output[38] )
         );
  XOR2_X1 U10383 ( .A1(\MC_ARK_ARC_1_3/temp2[38] ), .A2(n4189), .Z(n6197) );
  NAND4_X2 U10384 ( .A1(n1454), .A2(
        \SB2_0_27/Component_Function_5/NAND4_in[2] ), .A3(n4335), .A4(n4487), 
        .ZN(\SB2_0_27/buf_output[5] ) );
  BUF_X4 U10385 ( .I(\SB1_4_27/buf_output[5] ), .Z(\SB2_4_27/i0_3 ) );
  XOR2_X1 U10387 ( .A1(\MC_ARK_ARC_1_1/temp5[8] ), .A2(n6362), .Z(
        \MC_ARK_ARC_1_1/buf_output[8] ) );
  XOR2_X1 U10388 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[58] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[34] ), .Z(\MC_ARK_ARC_1_1/temp2[88] ) );
  NAND3_X2 U10390 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0_4 ), .A3(
        \SB2_1_23/i0_0 ), .ZN(\SB2_1_23/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U10391 ( .A1(\RI5[1][179] ), .A2(\RI5[1][155] ), .Z(
        \MC_ARK_ARC_1_1/temp2[17] ) );
  NAND4_X2 U10398 ( .A1(\SB2_2_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_25/Component_Function_5/NAND4_in[1] ), .A3(n6629), .A4(
        \SB2_2_25/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_25/buf_output[5] ) );
  NAND3_X1 U10401 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i0_3 ), .A3(
        \SB4_11/i0[9] ), .ZN(n7535) );
  NAND4_X2 U10405 ( .A1(\SB1_4_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_24/Component_Function_3/NAND4_in[1] ), .A3(n6236), .A4(n6973), 
        .ZN(\SB1_4_24/buf_output[3] ) );
  XOR2_X1 U10410 ( .A1(n6199), .A2(\MC_ARK_ARC_1_1/temp3[63] ), .Z(n6226) );
  XOR2_X1 U10411 ( .A1(\RI5[1][63] ), .A2(\RI5[1][57] ), .Z(n6199) );
  NAND4_X2 U10412 ( .A1(\SB2_2_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_26/Component_Function_3/NAND4_in[2] ), .A3(n6603), .A4(n4873), 
        .ZN(\SB2_2_26/buf_output[3] ) );
  NAND4_X2 U10415 ( .A1(\SB2_4_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_27/Component_Function_4/NAND4_in[1] ), .A3(n7208), .A4(
        \SB2_4_27/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_4_27/buf_output[4] ) );
  NAND3_X1 U10417 ( .A1(\SB1_3_30/i0[8] ), .A2(\SB1_3_30/i3[0] ), .A3(
        \SB1_3_30/i1_5 ), .ZN(\SB1_3_30/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U10418 ( .A1(\RI5[4][34] ), .A2(\RI5[4][190] ), .Z(n4519) );
  NAND3_X1 U10419 ( .A1(\SB1_3_18/i0_4 ), .A2(\SB1_3_18/i1_5 ), .A3(
        \SB1_3_18/i1[9] ), .ZN(n6223) );
  XOR2_X1 U10425 ( .A1(n5034), .A2(n4310), .Z(\MC_ARK_ARC_1_4/buf_output[75] )
         );
  XOR2_X1 U10426 ( .A1(\RI5[3][92] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[128] ), 
        .Z(n1045) );
  NAND3_X2 U10427 ( .A1(\SB2_2_21/i0_3 ), .A2(\SB1_2_22/buf_output[4] ), .A3(
        \SB2_2_21/i0[10] ), .ZN(n6862) );
  NAND3_X2 U10429 ( .A1(\SB3_19/i0[10] ), .A2(\SB3_19/i1[9] ), .A3(
        \SB3_19/i1_5 ), .ZN(n6387) );
  XOR2_X1 U10430 ( .A1(n2204), .A2(\MC_ARK_ARC_1_3/temp1[163] ), .Z(n7494) );
  NAND4_X2 U10439 ( .A1(\SB2_2_17/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_17/Component_Function_1/NAND4_in[3] ), .A3(n6477), .A4(
        \SB2_2_17/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_2_17/buf_output[1] ) );
  NAND3_X2 U10441 ( .A1(\SB1_3_11/i0[9] ), .A2(\SB1_3_11/i0[10] ), .A3(
        \SB1_3_11/i0_3 ), .ZN(n1196) );
  NAND4_X2 U10442 ( .A1(\SB2_3_17/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_17/Component_Function_1/NAND4_in[0] ), .A4(n6200), .ZN(
        \SB2_3_17/buf_output[1] ) );
  NAND2_X2 U10443 ( .A1(\SB1_4_7/i0_0 ), .A2(\SB1_4_7/i3[0] ), .ZN(n6201) );
  BUF_X4 U10444 ( .I(\RI1[5][173] ), .Z(\SB3_3/i0_3 ) );
  NAND3_X1 U10445 ( .A1(\SB4_30/i0[9] ), .A2(\SB4_30/i0[10] ), .A3(
        \SB4_30/i0_3 ), .ZN(n6202) );
  XOR2_X1 U10446 ( .A1(\MC_ARK_ARC_1_3/temp2[132] ), .A2(n6203), .Z(n5175) );
  XOR2_X1 U10449 ( .A1(\RI5[3][132] ), .A2(\RI5[3][126] ), .Z(n6203) );
  NAND3_X1 U10450 ( .A1(\SB2_1_3/i1_5 ), .A2(\SB1_1_8/buf_output[0] ), .A3(
        \SB1_1_7/buf_output[1] ), .ZN(
        \SB2_1_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U10454 ( .A1(\SB2_2_17/i0_3 ), .A2(\RI3[2][88] ), .A3(
        \SB2_2_17/i0_0 ), .ZN(\SB2_2_17/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U10456 ( .A1(\SB3_30/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_30/Component_Function_1/NAND4_in[0] ), .A3(
        \SB3_30/Component_Function_1/NAND4_in[1] ), .A4(n6204), .ZN(
        \SB3_30/buf_output[1] ) );
  NAND3_X1 U10457 ( .A1(\SB1_4_31/i0_3 ), .A2(\SB1_4_31/i0[6] ), .A3(
        \SB1_4_31/i0[10] ), .ZN(\SB1_4_31/Component_Function_2/NAND4_in[1] )
         );
  NAND2_X2 U10459 ( .A1(\SB1_4_6/i3[0] ), .A2(\SB1_4_6/i0_0 ), .ZN(
        \SB1_4_6/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U10461 ( .I(\SB1_3_20/buf_output[2] ), .ZN(\SB2_3_17/i1[9] ) );
  NAND4_X2 U10464 ( .A1(\SB1_3_20/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_20/Component_Function_2/NAND4_in[3] ), .A3(n7325), .A4(
        \SB1_3_20/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_3_20/buf_output[2] ) );
  NAND3_X2 U10469 ( .A1(\SB4_21/i0[10] ), .A2(\SB4_21/i0_3 ), .A3(
        \SB4_21/i0[6] ), .ZN(\SB4_21/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U10473 ( .A1(n6206), .A2(\MC_ARK_ARC_1_4/temp3[56] ), .Z(n4798) );
  XOR2_X1 U10475 ( .A1(\RI5[4][56] ), .A2(\RI5[4][50] ), .Z(n6206) );
  NAND4_X2 U10478 ( .A1(\SB1_2_12/Component_Function_2/NAND4_in[0] ), .A2(
        n2438), .A3(\SB1_2_12/Component_Function_2/NAND4_in[2] ), .A4(n6207), 
        .ZN(\SB1_2_12/buf_output[2] ) );
  NAND3_X2 U10483 ( .A1(\SB1_2_12/i0[10] ), .A2(\SB1_2_12/i0[6] ), .A3(
        \RI1[2][119] ), .ZN(n6207) );
  NAND4_X2 U10485 ( .A1(n2092), .A2(\SB4_19/Component_Function_4/NAND4_in[3] ), 
        .A3(\SB4_19/Component_Function_4/NAND4_in[1] ), .A4(n6208), .ZN(n7319)
         );
  NAND3_X1 U10487 ( .A1(\SB4_19/i0_0 ), .A2(\SB4_19/i0[9] ), .A3(
        \SB4_19/i0[8] ), .ZN(n6208) );
  INV_X2 U10488 ( .I(\MC_ARK_ARC_1_3/buf_output[95] ), .ZN(\SB1_4_16/i1_5 ) );
  XOR2_X1 U10489 ( .A1(n4978), .A2(\MC_ARK_ARC_1_4/temp4[99] ), .Z(
        \MC_ARK_ARC_1_4/temp6[99] ) );
  NAND3_X2 U10495 ( .A1(\SB2_4_13/i1[9] ), .A2(\SB2_4_13/i0_3 ), .A3(
        \SB2_4_13/i0[6] ), .ZN(\SB2_4_13/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U10496 ( .I(\SB1_3_7/buf_output[2] ), .ZN(\SB2_3_4/i1[9] ) );
  NAND4_X2 U10497 ( .A1(\SB1_3_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_7/Component_Function_2/NAND4_in[2] ), .A4(n1247), .ZN(
        \SB1_3_7/buf_output[2] ) );
  XOR2_X1 U10500 ( .A1(n1104), .A2(\MC_ARK_ARC_1_2/temp5[183] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[183] ) );
  XOR2_X1 U10501 ( .A1(n4025), .A2(n4026), .Z(\MC_ARK_ARC_1_2/temp5[183] ) );
  NAND3_X2 U10504 ( .A1(\SB2_4_20/i1_5 ), .A2(\SB2_4_20/i0_0 ), .A3(
        \SB2_4_20/i0_4 ), .ZN(\SB2_4_20/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U10505 ( .A1(n1980), .A2(n6209), .Z(\MC_ARK_ARC_1_2/temp5[28] ) );
  XOR2_X1 U10510 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[28] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[22] ), .Z(n6209) );
  NAND4_X2 U10511 ( .A1(\SB2_3_12/Component_Function_2/NAND4_in[0] ), .A2(
        n7478), .A3(\SB2_3_12/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_3_12/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_3_12/buf_output[2] ) );
  XOR2_X1 U10513 ( .A1(\MC_ARK_ARC_1_0/temp5[93] ), .A2(n6210), .Z(
        \MC_ARK_ARC_1_0/buf_output[93] ) );
  XOR2_X1 U10518 ( .A1(\MC_ARK_ARC_1_0/temp4[93] ), .A2(
        \MC_ARK_ARC_1_0/temp3[93] ), .Z(n6210) );
  INV_X2 U10520 ( .I(\SB1_2_18/buf_output[2] ), .ZN(\SB2_2_15/i1[9] ) );
  NAND4_X2 U10521 ( .A1(n4390), .A2(n3554), .A3(
        \SB1_2_18/Component_Function_2/NAND4_in[2] ), .A4(n1817), .ZN(
        \SB1_2_18/buf_output[2] ) );
  NAND3_X2 U10522 ( .A1(\SB2_3_20/i0[9] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \SB2_3_20/i0[8] ), .ZN(\SB2_3_20/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U10523 ( .A1(\SB1_2_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_27/Component_Function_0/NAND4_in[1] ), .A3(n7116), .A4(n6211), 
        .ZN(\SB1_2_27/buf_output[0] ) );
  NAND3_X2 U10525 ( .A1(\SB1_2_27/i0_0 ), .A2(\SB1_2_27/i0_3 ), .A3(
        \SB1_2_27/i0[7] ), .ZN(n6211) );
  NAND4_X2 U10526 ( .A1(\SB4_30/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_30/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_30/Component_Function_0/NAND4_in[0] ), .A4(n6212), .ZN(n4765) );
  NAND3_X1 U10529 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i0[6] ), .A3(
        \SB2_0_11/i1[9] ), .ZN(\SB2_0_11/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U10531 ( .A1(n4120), .A2(n6213), .Z(\MC_ARK_ARC_1_2/buf_output[23] )
         );
  XOR2_X1 U10533 ( .A1(n745), .A2(n6214), .Z(n3574) );
  XOR2_X1 U10534 ( .A1(\RI5[1][191] ), .A2(\RI5[1][167] ), .Z(n6214) );
  NAND4_X2 U10536 ( .A1(\SB1_1_20/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_1_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_20/Component_Function_1/NAND4_in[0] ), .A4(n6215), .ZN(
        \SB1_1_20/buf_output[1] ) );
  NAND3_X1 U10537 ( .A1(\SB1_1_20/i0[8] ), .A2(\SB1_1_20/i0_4 ), .A3(
        \SB1_1_20/i1_7 ), .ZN(n6215) );
  XOR2_X1 U10540 ( .A1(\MC_ARK_ARC_1_0/temp5[69] ), .A2(n6216), .Z(
        \MC_ARK_ARC_1_0/buf_output[69] ) );
  XOR2_X1 U10543 ( .A1(\MC_ARK_ARC_1_0/temp3[69] ), .A2(
        \MC_ARK_ARC_1_0/temp4[69] ), .Z(n6216) );
  NAND4_X2 U10544 ( .A1(\SB2_1_16/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_16/Component_Function_2/NAND4_in[0] ), .A3(n5393), .A4(n6217), 
        .ZN(\SB2_1_16/buf_output[2] ) );
  NAND3_X2 U10547 ( .A1(\SB2_1_16/i0[6] ), .A2(\SB2_1_16/i0[10] ), .A3(
        \SB2_1_16/i0_3 ), .ZN(n6217) );
  NAND3_X2 U10550 ( .A1(\SB1_4_25/i1_7 ), .A2(\SB1_4_25/i0[10] ), .A3(
        \SB1_4_25/i1[9] ), .ZN(n7177) );
  BUF_X4 U10557 ( .I(\SB3_16/buf_output[5] ), .Z(\SB4_16/i0_3 ) );
  NAND4_X2 U10558 ( .A1(\SB2_0_9/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_9/Component_Function_5/NAND4_in[0] ), .A3(n1708), .A4(n6218), 
        .ZN(\SB2_0_9/buf_output[5] ) );
  NAND3_X2 U10559 ( .A1(\SB2_0_9/i0_4 ), .A2(\SB2_0_9/i0[9] ), .A3(
        \SB2_0_9/i0[6] ), .ZN(n6218) );
  XOR2_X1 U10560 ( .A1(n6219), .A2(n213), .Z(Ciphertext[172]) );
  NAND4_X2 U10562 ( .A1(n2789), .A2(n2417), .A3(n2026), .A4(
        \SB4_3/Component_Function_4/NAND4_in[0] ), .ZN(n6219) );
  NAND3_X2 U10563 ( .A1(\SB3_16/i0[10] ), .A2(\SB3_16/i0[6] ), .A3(
        \SB3_16/i0_0 ), .ZN(\SB3_16/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U10564 ( .A1(\SB2_3_13/i0[10] ), .A2(\SB2_3_13/i0_3 ), .A3(
        \SB2_3_13/i0[6] ), .ZN(n6221) );
  NAND3_X1 U10565 ( .A1(\SB4_7/i0[9] ), .A2(n3965), .A3(\SB4_7/i0_0 ), .ZN(
        n6222) );
  NAND4_X2 U10571 ( .A1(\SB1_3_18/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_3_18/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_3_18/Component_Function_4/NAND4_in[1] ), .A4(n6223), .ZN(
        \SB1_3_18/buf_output[4] ) );
  NAND3_X1 U10578 ( .A1(\SB3_12/i0_0 ), .A2(\RI1[5][119] ), .A3(\SB3_12/i0[7] ), .ZN(n2580) );
  INV_X2 U10579 ( .I(\MC_ARK_ARC_1_2/buf_output[93] ), .ZN(\SB1_3_16/i0[8] )
         );
  NAND4_X2 U10581 ( .A1(\SB2_0_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_17/Component_Function_2/NAND4_in[2] ), .A3(n3884), .A4(n6224), 
        .ZN(\SB2_0_17/buf_output[2] ) );
  NAND3_X2 U10586 ( .A1(\SB2_0_17/i0_0 ), .A2(\SB2_0_17/i1_5 ), .A3(
        \RI3[0][88] ), .ZN(n6224) );
  XOR2_X1 U10590 ( .A1(n6226), .A2(n6225), .Z(\MC_ARK_ARC_1_1/buf_output[63] )
         );
  XOR2_X1 U10593 ( .A1(\MC_ARK_ARC_1_1/temp2[63] ), .A2(
        \MC_ARK_ARC_1_1/temp4[63] ), .Z(n6225) );
  XOR2_X1 U10599 ( .A1(n6228), .A2(n6227), .Z(\MC_ARK_ARC_1_1/temp6[32] ) );
  XOR2_X1 U10600 ( .A1(\RI5[1][98] ), .A2(n509), .Z(n6227) );
  XOR2_X1 U10606 ( .A1(\RI5[1][68] ), .A2(\RI5[1][134] ), .Z(n6228) );
  INV_X1 U10607 ( .I(\SB1_0_5/buf_output[0] ), .ZN(\SB2_0_0/i3[0] ) );
  NAND4_X2 U10612 ( .A1(\SB1_0_5/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_0_5/Component_Function_0/NAND4_in[3] ), .A3(n7161), .A4(
        \SB1_0_5/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_5/buf_output[0] ) );
  NAND3_X2 U10613 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i1[9] ), .A3(
        \SB1_0_18/i0_4 ), .ZN(\SB1_0_18/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U10618 ( .A1(n6229), .A2(n4632), .Z(\MC_ARK_ARC_1_2/temp5[110] ) );
  XOR2_X1 U10619 ( .A1(\RI5[2][80] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .Z(n6229) );
  XOR2_X1 U10621 ( .A1(n6230), .A2(n142), .Z(Ciphertext[124]) );
  NAND4_X2 U10622 ( .A1(\SB4_11/Component_Function_4/NAND4_in[0] ), .A2(n1461), 
        .A3(n7535), .A4(n7324), .ZN(n6230) );
  NAND2_X1 U10623 ( .A1(\SB1_0_30/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_30/Component_Function_4/NAND4_in[0] ), .ZN(n6231) );
  NAND4_X2 U10626 ( .A1(\SB1_2_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_17/Component_Function_4/NAND4_in[2] ), .A4(n6232), .ZN(
        \SB1_2_17/buf_output[4] ) );
  NAND3_X2 U10628 ( .A1(\SB1_2_17/i0_4 ), .A2(\SB1_2_17/i1[9] ), .A3(
        \SB1_2_17/i1_5 ), .ZN(n6232) );
  NAND3_X1 U10629 ( .A1(\SB4_30/i0_4 ), .A2(n5427), .A3(\SB4_30/i1_5 ), .ZN(
        n6233) );
  BUF_X4 U10631 ( .I(\MC_ARK_ARC_1_3/buf_output[146] ), .Z(\SB1_4_7/i0_0 ) );
  NAND4_X2 U10632 ( .A1(\SB2_2_7/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_7/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_2_7/Component_Function_1/NAND4_in[2] ), .A4(n6234), .ZN(
        \SB2_2_7/buf_output[1] ) );
  NAND3_X2 U10633 ( .A1(\SB2_2_7/i0_4 ), .A2(\SB2_2_7/i1_7 ), .A3(
        \SB2_2_7/i0[8] ), .ZN(n6234) );
  XOR2_X1 U10634 ( .A1(\RI5[0][55] ), .A2(\RI5[0][79] ), .Z(
        \MC_ARK_ARC_1_0/temp2[109] ) );
  XOR2_X1 U10638 ( .A1(n6235), .A2(\MC_ARK_ARC_1_2/temp4[181] ), .Z(n5174) );
  XOR2_X1 U10641 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[55] ), .A2(\RI5[2][91] ), 
        .Z(n6235) );
  NAND3_X2 U10642 ( .A1(\SB1_4_24/i0[10] ), .A2(\SB1_4_24/i1_7 ), .A3(
        \SB1_4_24/i1[9] ), .ZN(n6236) );
  XOR2_X1 U10644 ( .A1(\SB2_1_16/buf_output[0] ), .A2(\RI5[1][156] ), .Z(
        \MC_ARK_ARC_1_1/temp3[54] ) );
  XOR2_X1 U10646 ( .A1(\MC_ARK_ARC_1_0/temp6[108] ), .A2(n6237), .Z(
        \MC_ARK_ARC_1_0/buf_output[108] ) );
  XOR2_X1 U10647 ( .A1(\MC_ARK_ARC_1_0/temp2[108] ), .A2(
        \MC_ARK_ARC_1_0/temp1[108] ), .Z(n6237) );
  BUF_X4 U10651 ( .I(\RI1[5][107] ), .Z(\SB3_14/i0_3 ) );
  NAND4_X2 U10652 ( .A1(\SB4_17/Component_Function_4/NAND4_in[0] ), .A2(n4931), 
        .A3(n2828), .A4(n6239), .ZN(n6251) );
  NAND3_X1 U10657 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i0[10] ), .A3(
        \SB4_17/i0[9] ), .ZN(n6239) );
  NAND3_X1 U10658 ( .A1(\SB1_3_2/i0[6] ), .A2(\SB1_3_2/i0[8] ), .A3(
        \SB1_3_2/i0[7] ), .ZN(\SB1_3_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U10659 ( .A1(\SB2_4_10/i0_4 ), .A2(\SB2_4_10/i1[9] ), .A3(n6269), 
        .ZN(\SB2_4_10/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U10664 ( .A1(\SB2_0_30/Component_Function_5/NAND4_in[1] ), .A2(
        n6240), .A3(\SB2_0_30/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_30/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_30/buf_output[5] ) );
  NAND3_X2 U10668 ( .A1(\SB2_0_30/i0_3 ), .A2(\SB2_0_30/i0_4 ), .A3(
        \SB2_0_30/i1[9] ), .ZN(n6240) );
  NAND4_X2 U10673 ( .A1(\SB1_4_4/Component_Function_1/NAND4_in[3] ), .A2(n7111), .A3(\SB1_4_4/Component_Function_1/NAND4_in[0] ), .A4(n6241), .ZN(
        \SB1_4_4/buf_output[1] ) );
  NAND4_X2 U10675 ( .A1(\SB1_2_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_4/Component_Function_4/NAND4_in[3] ), .A4(n6242), .ZN(
        \SB1_2_4/buf_output[4] ) );
  NAND3_X2 U10676 ( .A1(\SB1_2_4/i0[10] ), .A2(\SB1_2_4/i0_3 ), .A3(
        \SB1_2_4/i0[9] ), .ZN(n6242) );
  XOR2_X1 U10677 ( .A1(\RI5[3][171] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[15] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[105] ) );
  NAND4_X2 U10684 ( .A1(\SB2_3_6/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_6/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_6/Component_Function_2/NAND4_in[0] ), .A4(n4922), .ZN(
        \SB2_3_6/buf_output[2] ) );
  INV_X4 U10689 ( .I(n6243), .ZN(\SB3_11/i1[9] ) );
  NAND3_X2 U10690 ( .A1(\SB2_2_9/i0_0 ), .A2(\SB2_2_9/i0[10] ), .A3(
        \SB2_2_9/i0[6] ), .ZN(n6244) );
  NAND4_X2 U10691 ( .A1(\SB3_1/Component_Function_4/NAND4_in[3] ), .A2(n1800), 
        .A3(\SB3_1/Component_Function_4/NAND4_in[2] ), .A4(n6245), .ZN(
        \SB3_1/buf_output[4] ) );
  NAND3_X1 U10695 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i3[0] ), .A3(\SB3_1/i1_7 ), 
        .ZN(n6245) );
  NAND4_X2 U10696 ( .A1(\SB3_24/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_24/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_24/Component_Function_1/NAND4_in[0] ), .A4(n6246), .ZN(
        \SB3_24/buf_output[1] ) );
  NAND3_X1 U10697 ( .A1(\SB3_24/i0[8] ), .A2(\SB3_24/i1_7 ), .A3(\SB3_24/i0_4 ), .ZN(n6246) );
  NAND4_X2 U10698 ( .A1(\SB4_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB4_21/Component_Function_4/NAND4_in[3] ), .A3(n4352), .A4(n6247), 
        .ZN(n7507) );
  NAND3_X1 U10700 ( .A1(\SB4_21/i1_7 ), .A2(\SB4_21/i3[0] ), .A3(
        \SB3_24/buf_output[2] ), .ZN(n6247) );
  XOR2_X1 U10701 ( .A1(\MC_ARK_ARC_1_3/temp2[57] ), .A2(n6248), .Z(n6658) );
  XOR2_X1 U10705 ( .A1(\RI5[3][57] ), .A2(\RI5[3][51] ), .Z(n6248) );
  XOR2_X1 U10706 ( .A1(n4036), .A2(n6249), .Z(\MC_ARK_ARC_1_1/temp5[123] ) );
  XOR2_X1 U10707 ( .A1(\RI5[1][69] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[117] ), 
        .Z(n6249) );
  INV_X2 U10710 ( .I(\MC_ARK_ARC_1_4/buf_output[68] ), .ZN(\SB3_20/i1[9] ) );
  INV_X2 U10717 ( .I(\SB1_2_11/buf_output[2] ), .ZN(\SB2_2_8/i1[9] ) );
  BUF_X4 U10718 ( .I(\MC_ARK_ARC_1_4/buf_output[71] ), .Z(\SB3_20/i0_3 ) );
  BUF_X4 U10719 ( .I(\MC_ARK_ARC_1_2/buf_output[14] ), .Z(\SB1_3_29/i0_0 ) );
  XOR2_X1 U10720 ( .A1(n6251), .A2(n126), .Z(Ciphertext[88]) );
  NAND4_X2 U10721 ( .A1(\SB2_3_29/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_29/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_29/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_29/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_29/buf_output[0] ) );
  BUF_X4 U10724 ( .I(\SB2_2_17/buf_output[2] ), .Z(\RI5[2][104] ) );
  BUF_X4 U10727 ( .I(\SB3_20/buf_output[5] ), .Z(\SB4_20/i0_3 ) );
  XOR2_X1 U10728 ( .A1(n5183), .A2(n6252), .Z(n6315) );
  NAND3_X2 U10732 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i1_7 ), .A3(
        \SB4_16/i1[9] ), .ZN(n1453) );
  NAND4_X2 U10734 ( .A1(\SB3_18/Component_Function_3/NAND4_in[1] ), .A2(n5138), 
        .A3(n6706), .A4(n6253), .ZN(\SB3_18/buf_output[3] ) );
  NAND3_X2 U10735 ( .A1(\SB3_18/i0[10] ), .A2(\SB3_18/i1[9] ), .A3(
        \SB3_18/i1_7 ), .ZN(n6253) );
  NAND3_X2 U10737 ( .A1(\SB2_4_30/i0_0 ), .A2(\SB2_4_30/i0[10] ), .A3(
        \SB2_4_30/i0[6] ), .ZN(\SB2_4_30/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U10742 ( .A1(n6636), .A2(n6254), .Z(n5039) );
  XOR2_X1 U10746 ( .A1(\RI5[4][11] ), .A2(\RI5[4][5] ), .Z(n6254) );
  INV_X1 U10747 ( .I(\SB1_1_5/buf_output[1] ), .ZN(\SB2_1_1/i1_7 ) );
  NAND4_X2 U10749 ( .A1(\SB1_1_5/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_5/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_1_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_5/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_5/buf_output[1] ) );
  NAND4_X2 U10750 ( .A1(\SB2_4_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_21/Component_Function_0/NAND4_in[0] ), .A4(n6255), .ZN(
        \SB2_4_21/buf_output[0] ) );
  NAND3_X1 U10752 ( .A1(\SB2_4_21/i0_3 ), .A2(\SB2_4_21/i0_0 ), .A3(
        \SB2_4_21/i0[7] ), .ZN(n6255) );
  NAND3_X2 U10753 ( .A1(\SB2_4_27/i0_3 ), .A2(\SB2_4_27/i0[9] ), .A3(
        \SB2_4_27/i0[8] ), .ZN(\SB2_4_27/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U10754 ( .A1(n4612), .A2(\SB2_0_4/Component_Function_4/NAND4_in[1] ), .A3(n1381), .A4(n6256), .ZN(\SB2_0_4/buf_output[4] ) );
  NAND3_X2 U10757 ( .A1(\SB1_4_0/i0_3 ), .A2(\SB1_4_0/i0[10] ), .A3(
        \SB1_4_0/i0_4 ), .ZN(\SB1_4_0/Component_Function_0/NAND4_in[2] ) );
  INV_X2 U10758 ( .I(\SB1_4_9/buf_output[5] ), .ZN(\SB2_4_9/i1_5 ) );
  BUF_X4 U10761 ( .I(\SB2_4_15/buf_output[3] ), .Z(\RI5[4][111] ) );
  NAND4_X2 U10765 ( .A1(\SB2_0_4/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_4/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_0_4/Component_Function_0/NAND4_in[0] ), .A4(n6258), .ZN(
        \SB2_0_4/buf_output[0] ) );
  NAND3_X2 U10769 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0_0 ), .A3(
        \SB2_0_4/i0[7] ), .ZN(n6258) );
  NAND4_X2 U10770 ( .A1(\SB2_0_29/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_29/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_0_29/Component_Function_0/NAND4_in[3] ), .A4(n6259), .ZN(
        \SB2_0_29/buf_output[0] ) );
  NAND3_X1 U10771 ( .A1(\SB2_0_29/i0[10] ), .A2(\SB2_0_29/i0_3 ), .A3(
        \SB2_0_29/i0_4 ), .ZN(n6259) );
  NAND3_X2 U10772 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i1[9] ), .A3(
        \SB1_1_26/i1_7 ), .ZN(n2392) );
  NAND3_X2 U10773 ( .A1(\SB2_4_4/i0[8] ), .A2(\SB2_4_4/i3[0] ), .A3(
        \SB2_4_4/i1_5 ), .ZN(n1638) );
  NAND3_X2 U10775 ( .A1(\SB2_1_29/i0_0 ), .A2(\SB2_1_29/i0_4 ), .A3(
        \SB2_1_29/i1_5 ), .ZN(n5217) );
  XOR2_X1 U10776 ( .A1(\RI5[1][170] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[164] ), .Z(n4058) );
  NAND4_X2 U10777 ( .A1(\SB1_1_0/Component_Function_2/NAND4_in[1] ), .A2(n6979), .A3(\SB1_1_0/Component_Function_2/NAND4_in[3] ), .A4(n6260), .ZN(
        \SB1_1_0/buf_output[2] ) );
  NAND3_X2 U10778 ( .A1(\SB1_1_0/i0[10] ), .A2(\SB1_1_0/i1[9] ), .A3(
        \SB1_1_0/i1_5 ), .ZN(n6260) );
  INV_X2 U10782 ( .I(\SB1_4_31/buf_output[5] ), .ZN(\SB2_4_31/i1_5 ) );
  INV_X2 U10784 ( .I(\SB1_3_30/buf_output[2] ), .ZN(\SB2_3_27/i1[9] ) );
  NAND4_X2 U10787 ( .A1(\SB1_3_30/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_30/Component_Function_2/NAND4_in[3] ), .A3(n6296), .A4(
        \SB1_3_30/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_3_30/buf_output[2] ) );
  XOR2_X1 U10790 ( .A1(\MC_ARK_ARC_1_2/temp2[9] ), .A2(n6261), .Z(n3307) );
  XOR2_X1 U10794 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[3] ), .A2(\RI5[2][9] ), 
        .Z(n6261) );
  XOR2_X1 U10796 ( .A1(n5212), .A2(n6262), .Z(n5301) );
  XOR2_X1 U10797 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[173] ), .A2(\RI5[4][5] ), 
        .Z(n6262) );
  NAND4_X2 U10801 ( .A1(\SB2_4_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_4_30/Component_Function_5/NAND4_in[0] ), .A3(
        \SB2_4_30/Component_Function_5/NAND4_in[1] ), .A4(n6263), .ZN(
        \SB2_4_30/buf_output[5] ) );
  NAND3_X2 U10803 ( .A1(\SB2_4_30/i0[9] ), .A2(\SB1_4_31/buf_output[4] ), .A3(
        \SB2_4_30/i0[6] ), .ZN(n6263) );
  NAND4_X2 U10804 ( .A1(\SB2_3_3/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_3/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_3/Component_Function_4/NAND4_in[1] ), .A4(n6264), .ZN(
        \SB2_3_3/buf_output[4] ) );
  NAND3_X1 U10805 ( .A1(\SB2_3_3/i0_0 ), .A2(\SB2_3_3/i0[9] ), .A3(
        \SB2_3_3/i0[8] ), .ZN(n6264) );
  NAND3_X2 U10806 ( .A1(\SB3_19/i0[8] ), .A2(\SB3_19/i0[7] ), .A3(
        \SB3_19/i0[6] ), .ZN(\SB3_19/Component_Function_0/NAND4_in[1] ) );
  BUF_X2 U10808 ( .I(n2554), .Z(n6265) );
  BUF_X4 U10811 ( .I(\MC_ARK_ARC_1_0/buf_output[8] ), .Z(\SB1_1_30/i0_0 ) );
  INV_X2 U10814 ( .I(\MC_ARK_ARC_1_4/buf_output[105] ), .ZN(\SB3_14/i0[8] ) );
  INV_X2 U10816 ( .I(\MC_ARK_ARC_1_0/buf_output[8] ), .ZN(\SB1_1_30/i1[9] ) );
  NAND3_X2 U10818 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i1[9] ), .A3(
        \SB1_1_26/i1_5 ), .ZN(n6440) );
  BUF_X4 U10822 ( .I(\SB3_19/buf_output[1] ), .Z(\SB4_15/i0[6] ) );
  NAND4_X2 U10827 ( .A1(\SB2_4_31/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_4_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_4_31/Component_Function_3/NAND4_in[0] ), .A4(
        \SB2_4_31/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_4_31/buf_output[3] ) );
  NAND3_X2 U10828 ( .A1(\SB1_4_1/i0[10] ), .A2(\SB1_4_1/i0_0 ), .A3(
        \SB1_4_1/i0[6] ), .ZN(\SB1_4_1/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U10831 ( .A1(\SB4_18/i0[10] ), .A2(\SB4_18/i0_3 ), .A3(
        \SB4_18/i0[9] ), .ZN(n7343) );
  NAND3_X1 U10836 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i0[10] ), .A3(
        \SB4_12/i0[6] ), .ZN(n7442) );
  OR3_X2 U10837 ( .A1(\MC_ARK_ARC_1_4/buf_output[3] ), .A2(n3981), .A3(
        \MC_ARK_ARC_1_4/buf_output[0] ), .Z(n3137) );
  NAND3_X1 U10841 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i0[10] ), .A3(\SB3_0/i0[6] ), 
        .ZN(\SB3_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U10844 ( .A1(\SB3_0/i0_0 ), .A2(\SB3_0/i0[6] ), .A3(\SB3_0/i0[10] ), 
        .ZN(\SB3_0/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U10848 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0[10] ), .A3(
        \SB2_3_26/i0[9] ), .ZN(n4740) );
  NAND3_X1 U10853 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0[10] ), .A3(
        \SB2_3_26/i0_4 ), .ZN(\SB2_3_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U10856 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0_0 ), .A3(n4081), 
        .ZN(n3596) );
  NAND3_X1 U10861 ( .A1(\SB2_3_26/i1[9] ), .A2(\SB2_3_26/i0_3 ), .A3(
        \SB2_3_26/i0[6] ), .ZN(\SB2_3_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10862 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0_4 ), .A3(
        \SB2_3_26/i0_0 ), .ZN(\SB2_3_26/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U10863 ( .I(\MC_ARK_ARC_1_1/buf_output[21] ), .Z(\SB1_2_28/i0[10] ) );
  BUF_X2 U10865 ( .I(\SB1_2_14/buf_output[0] ), .Z(\SB2_2_9/i0[9] ) );
  NAND4_X2 U10871 ( .A1(\SB3_30/Component_Function_0/NAND4_in[1] ), .A2(
        \SB3_30/Component_Function_0/NAND4_in[3] ), .A3(
        \SB3_30/Component_Function_0/NAND4_in[0] ), .A4(n1183), .ZN(n6266) );
  NAND3_X2 U10872 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0[10] ), .A3(
        \SB3_30/i0_4 ), .ZN(n1183) );
  NAND3_X1 U10873 ( .A1(\SB3_24/i0[9] ), .A2(\SB3_24/i0_0 ), .A3(
        \SB3_24/i0[8] ), .ZN(\SB3_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U10879 ( .A1(\SB3_14/i0[8] ), .A2(\SB3_14/i0_3 ), .A3(
        \SB3_14/i0[9] ), .ZN(n6752) );
  NAND3_X1 U10880 ( .A1(\SB3_14/i0[8] ), .A2(\SB3_14/i1_5 ), .A3(
        \SB3_14/i3[0] ), .ZN(n7357) );
  NAND3_X1 U10881 ( .A1(\SB1_4_5/i0[10] ), .A2(\SB1_4_5/i0[6] ), .A3(
        \SB1_4_5/i0_0 ), .ZN(\SB1_4_5/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X4 U10882 ( .I(\SB3_7/buf_output[4] ), .Z(\SB4_6/i0_4 ) );
  CLKBUF_X4 U10887 ( .I(\SB1_4_3/buf_output[3] ), .Z(\SB2_4_1/i0[10] ) );
  BUF_X2 U10892 ( .I(\MC_ARK_ARC_1_4/buf_output[142] ), .Z(\SB3_8/i0_4 ) );
  NAND3_X1 U10893 ( .A1(\SB2_4_4/i0[9] ), .A2(\SB2_4_4/i0_0 ), .A3(
        \SB2_4_4/i0[8] ), .ZN(\SB2_4_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U10894 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i0[9] ), .A3(
        \SB4_29/i0_3 ), .ZN(n3724) );
  CLKBUF_X4 U10895 ( .I(\SB2_2_25/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[41] ) );
  CLKBUF_X4 U10897 ( .I(\SB1_1_17/buf_output[2] ), .Z(\SB2_1_14/i0_0 ) );
  AND4_X2 U10898 ( .A1(\SB1_2_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_5/Component_Function_2/NAND4_in[1] ), .A3(n2685), .A4(
        \SB1_2_5/Component_Function_2/NAND4_in[2] ), .Z(n6267) );
  NAND3_X1 U10904 ( .A1(\SB2_4_22/i0_0 ), .A2(\SB2_4_22/i0_3 ), .A3(
        \SB2_4_22/i0_4 ), .ZN(\SB2_4_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U10905 ( .A1(\SB3_21/i0_0 ), .A2(\SB3_21/i0_4 ), .A3(\SB3_21/i0_3 ), 
        .ZN(\SB3_21/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U10906 ( .I(\SB1_4_5/buf_output[4] ), .Z(\SB2_4_4/i0_4 ) );
  AND2_X1 U10907 ( .A1(\SB1_4_5/buf_output[4] ), .A2(\SB1_4_4/buf_output[5] ), 
        .Z(n3178) );
  NAND2_X1 U10908 ( .A1(\SB3_27/i0_3 ), .A2(\SB3_27/i1[9] ), .ZN(
        \SB3_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10909 ( .A1(\SB3_27/i0_3 ), .A2(\SB3_27/i0_4 ), .A3(\SB3_27/i1[9] ), .ZN(n7335) );
  AND4_X2 U10910 ( .A1(\SB1_4_24/Component_Function_5/NAND4_in[1] ), .A2(n6871), .A3(n4108), .A4(\SB1_4_24/Component_Function_5/NAND4_in[0] ), .Z(n6268) );
  NAND2_X1 U10911 ( .A1(\SB1_4_24/i0_0 ), .A2(\SB1_4_24/i3[0] ), .ZN(
        \SB1_4_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U10912 ( .A1(\SB2_4_1/i0_3 ), .A2(\SB2_4_1/i0_4 ), .A3(
        \SB2_4_1/i1[9] ), .ZN(\SB2_4_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U10914 ( .A1(\SB2_4_1/i1[9] ), .A2(n6277), .A3(\SB2_4_1/i0_4 ), 
        .ZN(n3717) );
  NAND3_X1 U10915 ( .A1(\SB2_4_1/i1[9] ), .A2(\SB2_4_1/i0_3 ), .A3(
        \SB2_4_1/i0[6] ), .ZN(\SB2_4_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10918 ( .A1(\SB2_3_17/i0[7] ), .A2(\SB2_3_17/i0_3 ), .A3(
        \SB2_3_17/i0_0 ), .ZN(\SB2_3_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U10920 ( .A1(\SB4_25/i0[10] ), .A2(\SB4_25/i0_3 ), .A3(
        \SB4_25/i0[6] ), .ZN(n2883) );
  CLKBUF_X4 U10922 ( .I(\SB3_13/buf_output[4] ), .Z(\SB4_12/i0_4 ) );
  NAND2_X1 U10923 ( .A1(\SB2_4_7/i0_0 ), .A2(\SB2_4_7/i3[0] ), .ZN(
        \SB2_4_7/Component_Function_5/NAND4_in[0] ) );
  AND4_X2 U10925 ( .A1(\SB1_4_10/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_4_10/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_4_10/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_4_10/Component_Function_5/NAND4_in[2] ), .Z(n6269) );
  NAND3_X2 U10928 ( .A1(\SB1_4_10/i0[9] ), .A2(\SB1_4_10/i0[6] ), .A3(
        \SB1_4_10/i0_4 ), .ZN(\SB1_4_10/Component_Function_5/NAND4_in[3] ) );
  CLKBUF_X4 U10931 ( .I(\SB1_4_13/buf_output[5] ), .Z(\SB2_4_13/i0_3 ) );
  NAND3_X1 U10932 ( .A1(\SB2_4_24/i0_4 ), .A2(\SB2_4_24/i1_7 ), .A3(
        \SB2_4_24/i0[8] ), .ZN(\SB2_4_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U10933 ( .A1(\SB1_4_24/i0_3 ), .A2(\SB1_4_24/i0[8] ), .A3(
        \SB1_4_24/i0[9] ), .ZN(\SB1_4_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U10934 ( .A1(\SB1_4_24/i0_3 ), .A2(\SB1_4_24/i1_7 ), .A3(
        \SB1_4_24/i0[8] ), .ZN(\SB1_4_24/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U10943 ( .A1(\SB1_4_24/i0_4 ), .A2(\MC_ARK_ARC_1_3/buf_output[47] ), 
        .A3(\SB1_4_24/i1[9] ), .ZN(n4108) );
  CLKBUF_X4 U10945 ( .I(\SB3_31/buf_output[3] ), .Z(\SB4_29/i0[10] ) );
  NAND3_X1 U10950 ( .A1(\SB2_4_2/i1_5 ), .A2(\SB2_4_2/i0_0 ), .A3(
        \SB2_4_2/i0_4 ), .ZN(\SB2_4_2/Component_Function_2/NAND4_in[3] ) );
  CLKBUF_X4 U10953 ( .I(\SB3_31/buf_output[0] ), .Z(\SB4_26/i0[9] ) );
  XOR2_X1 U10954 ( .A1(n3037), .A2(n2186), .Z(n6271) );
  CLKBUF_X4 U10959 ( .I(\MC_ARK_ARC_1_4/buf_output[110] ), .Z(\SB3_13/i0_0 )
         );
  CLKBUF_X4 U10960 ( .I(\SB1_3_31/buf_output[3] ), .Z(\SB2_3_29/i0[10] ) );
  NAND3_X1 U10965 ( .A1(\SB2_4_4/i0_4 ), .A2(\SB2_4_4/i1_7 ), .A3(
        \SB2_4_4/i0[8] ), .ZN(\SB2_4_4/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 U10966 ( .I(\SB1_2_8/buf_output[0] ), .Z(\SB2_2_3/i0[9] ) );
  CLKBUF_X4 U10970 ( .I(\MC_ARK_ARC_1_4/buf_output[27] ), .Z(\SB3_27/i0[10] )
         );
  CLKBUF_X4 U10972 ( .I(\MC_ARK_ARC_1_4/buf_output[140] ), .Z(\SB3_8/i0_0 ) );
  BUF_X2 U10973 ( .I(\RI3[5][73] ), .Z(\SB4_19/i0[6] ) );
  CLKBUF_X4 U10978 ( .I(\SB1_2_22/buf_output[2] ), .Z(\SB2_2_19/i0_0 ) );
  CLKBUF_X4 U10980 ( .I(\SB3_25/buf_output[5] ), .Z(\SB4_25/i0_3 ) );
  NAND4_X2 U10981 ( .A1(\SB3_10/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_10/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_10/Component_Function_4/NAND4_in[3] ), .A4(n5307), .ZN(n6272) );
  NAND3_X1 U10984 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i0[9] ), .A3(
        \SB4_12/i0[8] ), .ZN(n7522) );
  CLKBUF_X4 U10985 ( .I(\SB1_4_29/buf_output[2] ), .Z(\SB2_4_26/i0_0 ) );
  NAND3_X1 U10989 ( .A1(\SB2_3_20/i0_0 ), .A2(\SB2_3_20/i0_3 ), .A3(n6819), 
        .ZN(\SB2_3_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U10992 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \RI3[3][70] ), .ZN(n2532) );
  CLKBUF_X4 U10994 ( .I(\SB2_1_22/buf_output[5] ), .Z(\RI5[1][59] ) );
  INV_X1 U10995 ( .I(\MC_ARK_ARC_1_3/buf_output[167] ), .ZN(\SB1_4_4/i1_5 ) );
  CLKBUF_X4 U10996 ( .I(\SB3_15/buf_output[5] ), .Z(\SB4_15/i0_3 ) );
  INV_X1 U10999 ( .I(\MC_ARK_ARC_1_2/buf_output[95] ), .ZN(\SB1_3_16/i1_5 ) );
  CLKBUF_X4 U11002 ( .I(\MC_ARK_ARC_1_2/buf_output[95] ), .Z(\SB1_3_16/i0_3 )
         );
  CLKBUF_X4 U11003 ( .I(\SB2_0_4/buf_output[0] ), .Z(\RI5[0][0] ) );
  CLKBUF_X4 U11005 ( .I(\MC_ARK_ARC_1_0/buf_output[15] ), .Z(\SB1_1_29/i0[10] ) );
  CLKBUF_X4 U11007 ( .I(\SB3_1/buf_output[4] ), .Z(\SB4_0/i0_4 ) );
  BUF_X2 U11008 ( .I(\MC_ARK_ARC_1_4/buf_output[79] ), .Z(\SB3_18/i0[6] ) );
  INV_X1 U11009 ( .I(\MC_ARK_ARC_1_4/buf_output[79] ), .ZN(\SB3_18/i1_7 ) );
  CLKBUF_X4 U11012 ( .I(\SB3_27/buf_output[2] ), .Z(\SB4_24/i0_0 ) );
  NAND3_X1 U11013 ( .A1(\SB3_18/i1_5 ), .A2(\SB3_18/i0[6] ), .A3(
        \SB3_18/i0[9] ), .ZN(\SB3_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U11014 ( .A1(\SB3_18/i0[9] ), .A2(\SB3_18/i0[6] ), .A3(
        \SB3_18/i0_4 ), .ZN(\SB3_18/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U11023 ( .A1(\SB2_4_11/i0_3 ), .A2(\SB2_4_11/i0_4 ), .A3(
        \SB2_4_11/i1[9] ), .ZN(n3517) );
  NAND3_X1 U11027 ( .A1(\SB3_21/i0[10] ), .A2(\SB3_21/i0_4 ), .A3(
        \SB3_21/i0_3 ), .ZN(\SB3_21/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U11028 ( .I(\SB2_4_14/buf_output[1] ), .Z(\RI5[4][127] ) );
  CLKBUF_X4 U11029 ( .I(\MC_ARK_ARC_1_4/buf_output[117] ), .Z(\SB3_12/i0[10] )
         );
  BUF_X2 U11032 ( .I(\MC_ARK_ARC_1_2/buf_output[84] ), .Z(\SB1_3_17/i0[9] ) );
  INV_X1 U11035 ( .I(\MC_ARK_ARC_1_2/buf_output[84] ), .ZN(\SB1_3_17/i3[0] )
         );
  CLKBUF_X4 U11036 ( .I(\MC_ARK_ARC_1_3/buf_output[114] ), .Z(\SB1_4_12/i0[9] ) );
  NAND3_X1 U11039 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i0[8] ), .A3(
        \SB1_2_18/i0[9] ), .ZN(n3865) );
  NAND3_X1 U11040 ( .A1(\SB3_16/i0_0 ), .A2(\SB3_16/i0_3 ), .A3(\SB3_16/i0_4 ), 
        .ZN(\SB3_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11043 ( .A1(\SB1_4_12/i1_5 ), .A2(\SB1_4_12/i0[6] ), .A3(
        \SB1_4_12/i0[9] ), .ZN(n4824) );
  CLKBUF_X4 U11046 ( .I(\SB1_2_22/buf_output[0] ), .Z(\SB2_2_17/i0[9] ) );
  CLKBUF_X4 U11047 ( .I(\SB2_4_9/buf_output[2] ), .Z(\RI5[4][152] ) );
  NAND3_X1 U11049 ( .A1(\SB2_3_11/i0[10] ), .A2(\SB2_3_11/i0_3 ), .A3(
        \SB2_3_11/i0_4 ), .ZN(n4372) );
  NAND3_X1 U11056 ( .A1(\SB1_3_12/buf_output[4] ), .A2(\SB2_3_11/i0[6] ), .A3(
        \SB2_3_11/i0[9] ), .ZN(\SB2_3_11/Component_Function_5/NAND4_in[3] ) );
  INV_X1 U11057 ( .I(\MC_ARK_ARC_1_2/buf_output[139] ), .ZN(\SB1_3_8/i1_7 ) );
  BUF_X2 U11059 ( .I(\MC_ARK_ARC_1_2/buf_output[139] ), .Z(\SB1_3_8/i0[6] ) );
  NAND3_X1 U11062 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i0[9] ), .A3(n1493), .ZN(
        n7557) );
  NAND3_X1 U11064 ( .A1(\SB2_4_30/i1_5 ), .A2(\SB2_4_30/i0[6] ), .A3(
        \SB2_4_30/i0[9] ), .ZN(\SB2_4_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U11065 ( .A1(\SB2_4_19/i0[10] ), .A2(\SB2_4_19/i0_4 ), .A3(
        \SB2_4_19/i0_3 ), .ZN(\SB2_4_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11066 ( .A1(\SB2_4_19/i0[9] ), .A2(\SB2_4_19/i0[10] ), .A3(
        \SB2_4_19/i0_3 ), .ZN(\SB2_4_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U11071 ( .A1(\SB2_4_19/i0_3 ), .A2(\SB2_4_19/i0_0 ), .A3(
        \SB2_4_19/i0[7] ), .ZN(n6600) );
  NAND3_X1 U11074 ( .A1(\SB2_4_19/i0_0 ), .A2(\SB1_4_19/buf_output[5] ), .A3(
        \SB2_4_19/i0_4 ), .ZN(\SB2_4_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11077 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i0_4 ), .A3(\SB4_12/i1_5 ), 
        .ZN(n2749) );
  NAND3_X1 U11078 ( .A1(\SB2_4_19/i0_4 ), .A2(\SB2_4_19/i0_0 ), .A3(
        \SB2_4_19/i1_5 ), .ZN(\SB2_4_19/Component_Function_2/NAND4_in[3] ) );
  NAND4_X1 U11079 ( .A1(\SB4_10/Component_Function_3/NAND4_in[1] ), .A2(n2739), 
        .A3(n2921), .A4(\SB4_10/Component_Function_3/NAND4_in[3] ), .ZN(n7410)
         );
  NAND3_X1 U11080 ( .A1(\SB2_0_31/i0[7] ), .A2(\SB2_0_31/i0[8] ), .A3(
        \SB2_0_31/i0[6] ), .ZN(n1251) );
  NAND3_X1 U11087 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i0_3 ), .A3(
        \SB4_29/i0[6] ), .ZN(n3763) );
  CLKBUF_X4 U11090 ( .I(\SB2_4_6/buf_output[0] ), .Z(\RI5[4][180] ) );
  NAND3_X1 U11097 ( .A1(\SB4_1/i0[6] ), .A2(\SB4_1/i0[10] ), .A3(\SB4_1/i0_3 ), 
        .ZN(n4224) );
  NAND3_X1 U11099 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i0[9] ), .A3(\SB3_2/i0[8] ), 
        .ZN(n4910) );
  NAND3_X1 U11107 ( .A1(\SB1_3_3/i0_3 ), .A2(\SB1_3_3/i1_7 ), .A3(
        \SB1_3_3/i0[8] ), .ZN(\SB1_3_3/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U11108 ( .A1(\SB1_3_3/i0[10] ), .A2(\SB1_3_3/i0_3 ), .A3(
        \SB1_3_3/i0[9] ), .ZN(\SB1_3_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U11109 ( .A1(\SB1_3_3/i0[10] ), .A2(\SB1_3_3/i0_3 ), .A3(
        \SB1_3_3/i0[6] ), .ZN(n7280) );
  NAND3_X1 U11110 ( .A1(\SB2_3_23/i0[10] ), .A2(\SB2_3_23/i1_7 ), .A3(
        \SB2_3_23/i1[9] ), .ZN(n2995) );
  NAND2_X1 U11111 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i1[9] ), .ZN(n6881) );
  NAND3_X1 U11113 ( .A1(\SB2_3_23/i1_5 ), .A2(\SB2_3_23/i0[10] ), .A3(
        \SB2_3_23/i1[9] ), .ZN(\SB2_3_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U11114 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i0_4 ), .A3(
        \SB2_3_23/i1[9] ), .ZN(\SB2_3_23/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U11115 ( .I(n290), .Z(\SB1_0_13/i0_0 ) );
  NAND3_X1 U11117 ( .A1(\SB2_4_31/i1[9] ), .A2(\SB2_4_31/i1_7 ), .A3(
        \SB2_4_31/i0[10] ), .ZN(\SB2_4_31/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U11122 ( .A1(\SB1_1_13/i3[0] ), .A2(\SB1_1_13/i0_0 ), .A3(
        \SB1_1_13/i1_7 ), .ZN(\SB1_1_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U11123 ( .A1(\SB1_4_9/i0_0 ), .A2(\SB1_4_9/i0_3 ), .A3(
        \SB1_4_9/i0_4 ), .ZN(\SB1_4_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11125 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i1_7 ), .A3(\SB4_10/i3[0] ), .ZN(n4286) );
  NAND2_X1 U11127 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i3[0] ), .ZN(n2925) );
  CLKBUF_X4 U11128 ( .I(\MC_ARK_ARC_1_2/buf_output[166] ), .Z(\SB1_3_4/i0_4 )
         );
  NAND3_X1 U11129 ( .A1(\SB1_3_28/i0[10] ), .A2(\SB1_3_28/i0_3 ), .A3(
        \SB1_3_28/i0[6] ), .ZN(n4977) );
  NAND3_X1 U11130 ( .A1(\SB1_3_28/i0[9] ), .A2(\SB1_3_28/i0[6] ), .A3(
        \SB1_3_28/i0_4 ), .ZN(n7094) );
  NAND3_X1 U11134 ( .A1(\SB1_3_28/i0[8] ), .A2(\SB1_3_28/i0[7] ), .A3(
        \SB1_3_28/i0[6] ), .ZN(\SB1_3_28/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U11135 ( .A1(\SB1_3_28/i1_5 ), .A2(\SB1_3_28/i0[6] ), .A3(
        \SB1_3_28/i0[9] ), .ZN(\SB1_3_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U11138 ( .A1(\RI1[5][119] ), .A2(\SB3_12/i0[10] ), .A3(
        \SB3_12/i0_4 ), .ZN(n2581) );
  CLKBUF_X4 U11140 ( .I(\MC_ARK_ARC_1_4/buf_output[119] ), .Z(\RI1[5][119] )
         );
  INV_X1 U11145 ( .I(\SB3_15/buf_output[0] ), .ZN(\SB4_10/i3[0] ) );
  NAND3_X1 U11147 ( .A1(\SB3_20/i0[7] ), .A2(\SB3_20/i0_3 ), .A3(\SB3_20/i0_0 ), .ZN(\SB3_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U11148 ( .A1(\SB3_20/i0_4 ), .A2(\SB3_20/i0[10] ), .A3(
        \SB3_20/i0_3 ), .ZN(\SB3_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11152 ( .A1(\SB2_4_31/i0_4 ), .A2(\SB2_4_31/i1[9] ), .A3(
        \SB2_4_31/i1_5 ), .ZN(n2469) );
  NAND3_X1 U11153 ( .A1(\SB2_4_31/i1_5 ), .A2(\SB2_4_31/i0[10] ), .A3(
        \SB2_4_31/i1[9] ), .ZN(\SB2_4_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U11156 ( .A1(\SB2_4_31/i1_5 ), .A2(\SB2_4_31/i0_0 ), .A3(
        \SB1_4_0/buf_output[4] ), .ZN(
        \SB2_4_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U11158 ( .A1(\RI1[5][17] ), .A2(\SB3_29/i0[10] ), .A3(
        \SB3_29/i0[6] ), .ZN(\SB3_29/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 U11163 ( .I(\SB2_4_22/buf_output[2] ), .Z(\RI5[4][74] ) );
  NAND3_X1 U11165 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i0[9] ), .A3(\SB4_2/i0[10] ), 
        .ZN(n6918) );
  CLKBUF_X4 U11166 ( .I(\MC_ARK_ARC_1_4/buf_output[166] ), .Z(\SB3_4/i0_4 ) );
  NAND3_X1 U11170 ( .A1(\SB1_4_17/i0[9] ), .A2(\SB1_4_17/i0[10] ), .A3(
        \SB1_4_17/i0_3 ), .ZN(\SB1_4_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U11171 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i1_7 ), .A3(\SB4_14/i3[0] ), .ZN(n7301) );
  NAND3_X1 U11172 ( .A1(\SB3_3/i0_0 ), .A2(\SB3_3/i0_3 ), .A3(\SB3_3/i0[7] ), 
        .ZN(n6516) );
  NAND3_X2 U11174 ( .A1(\SB3_23/i1_5 ), .A2(\SB3_23/i0[8] ), .A3(
        \SB3_23/i3[0] ), .ZN(n7071) );
  NAND3_X1 U11177 ( .A1(\SB3_23/i1_5 ), .A2(\SB3_23/i0[6] ), .A3(
        \SB3_23/i0[9] ), .ZN(\SB3_23/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 U11178 ( .I(n1491), .Z(\SB1_4_10/i0[10] ) );
  CLKBUF_X4 U11184 ( .I(\MC_ARK_ARC_1_4/buf_output[83] ), .Z(\SB3_18/i0_3 ) );
  INV_X1 U11185 ( .I(\MC_ARK_ARC_1_4/buf_output[83] ), .ZN(\SB3_18/i1_5 ) );
  INV_X1 U11186 ( .I(\SB3_18/buf_output[0] ), .ZN(\SB4_13/i3[0] ) );
  BUF_X2 U11187 ( .I(\SB3_18/buf_output[0] ), .Z(\SB4_13/i0[9] ) );
  NAND2_X1 U11189 ( .A1(\SB4_21/i0[10] ), .A2(\SB4_21/i0[9] ), .ZN(
        \SB4_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U11192 ( .A1(\SB1_4_8/i0[9] ), .A2(\SB1_4_8/i0[10] ), .A3(
        \SB1_4_8/i0_3 ), .ZN(\SB1_4_8/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U11193 ( .A1(\SB1_4_8/i0_3 ), .A2(\SB1_4_8/i1[9] ), .ZN(
        \SB1_4_8/Component_Function_1/NAND4_in[0] ) );
  CLKBUF_X2 U11194 ( .I(Key[56]), .Z(n154) );
  CLKBUF_X4 U11195 ( .I(\MC_ARK_ARC_1_0/buf_output[62] ), .Z(\SB1_1_21/i0_0 )
         );
  CLKBUF_X4 U11196 ( .I(\MC_ARK_ARC_1_3/buf_output[48] ), .Z(\SB1_4_23/i0[9] )
         );
  NAND3_X1 U11197 ( .A1(\SB3_21/i0[6] ), .A2(\SB3_21/i1[9] ), .A3(
        \SB3_21/i0_3 ), .ZN(\SB3_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U11203 ( .A1(\SB2_4_27/i0[10] ), .A2(\SB2_4_27/i0_3 ), .A3(
        \SB2_4_27/i0_4 ), .ZN(\SB2_4_27/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U11204 ( .I(\SB2_2_22/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[79] ) );
  CLKBUF_X4 U11205 ( .I(\SB2_4_9/buf_output[5] ), .Z(\RI5[4][137] ) );
  INV_X1 U11209 ( .I(\MC_ARK_ARC_1_4/buf_output[95] ), .ZN(\SB3_16/i1_5 ) );
  NAND3_X1 U11212 ( .A1(\SB3_16/i1_5 ), .A2(\SB3_16/i0[6] ), .A3(
        \SB3_16/i0[9] ), .ZN(\SB3_16/Component_Function_1/NAND4_in[2] ) );
  INV_X1 U11216 ( .I(\MC_ARK_ARC_1_3/buf_output[23] ), .ZN(\SB1_4_28/i1_5 ) );
  CLKBUF_X4 U11220 ( .I(\MC_ARK_ARC_1_3/buf_output[23] ), .Z(\SB1_4_28/i0_3 )
         );
  BUF_X4 U11221 ( .I(\SB2_3_24/buf_output[4] ), .Z(\RI5[3][52] ) );
  AND4_X2 U11222 ( .A1(n2337), .A2(\SB3_19/Component_Function_5/NAND4_in[1] ), 
        .A3(n5411), .A4(\SB3_19/Component_Function_5/NAND4_in[0] ), .Z(n6273)
         );
  NAND3_X1 U11225 ( .A1(\SB3_6/i3[0] ), .A2(\SB3_6/i0_0 ), .A3(\SB3_6/i1_7 ), 
        .ZN(\SB3_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U11226 ( .A1(\SB2_1_29/i0[10] ), .A2(\SB2_1_29/i0_4 ), .A3(
        \SB2_1_29/i0_3 ), .ZN(\SB2_1_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11227 ( .A1(\SB2_1_29/i0_0 ), .A2(\SB2_1_29/i0_4 ), .A3(
        \SB2_1_29/i0_3 ), .ZN(\SB2_1_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11231 ( .A1(\SB2_1_29/i0[6] ), .A2(\SB2_1_29/i0[9] ), .A3(
        \SB2_1_29/i0_4 ), .ZN(n1582) );
  CLKBUF_X4 U11234 ( .I(\SB1_4_1/buf_output[3] ), .Z(\SB2_4_31/i0[10] ) );
  CLKBUF_X4 U11241 ( .I(\MC_ARK_ARC_1_1/buf_output[184] ), .Z(\SB1_2_1/i0_4 )
         );
  NAND3_X1 U11245 ( .A1(\SB2_4_20/i3[0] ), .A2(\SB2_4_20/i1_5 ), .A3(
        \SB2_4_20/i0[8] ), .ZN(n1208) );
  INV_X1 U11246 ( .I(\SB1_4_0/buf_output[1] ), .ZN(\SB2_4_28/i1_7 ) );
  CLKBUF_X4 U11248 ( .I(\SB2_1_29/buf_output[0] ), .Z(\RI5[1][42] ) );
  CLKBUF_X4 U11250 ( .I(\MC_ARK_ARC_1_3/buf_output[56] ), .Z(\SB1_4_22/i0_0 )
         );
  NAND3_X1 U11251 ( .A1(\SB2_4_31/i0_3 ), .A2(\SB2_4_31/i0[8] ), .A3(
        \SB2_4_31/i0[9] ), .ZN(\SB2_4_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11259 ( .A1(\SB2_4_31/i0[10] ), .A2(\SB2_4_31/i0_3 ), .A3(
        \SB2_4_31/i0[6] ), .ZN(\SB2_4_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U11260 ( .A1(\SB2_4_31/i0_3 ), .A2(\SB2_4_31/i0_0 ), .A3(
        \SB2_4_31/i0_4 ), .ZN(\SB2_4_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11266 ( .A1(\SB2_4_31/i0[10] ), .A2(\SB2_4_31/i0_4 ), .A3(
        \SB2_4_31/i0_3 ), .ZN(\SB2_4_31/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U11267 ( .I(\SB1_3_17/buf_output[2] ), .Z(\SB2_3_14/i0_0 ) );
  NAND3_X1 U11268 ( .A1(\SB4_6/i0[9] ), .A2(\SB4_6/i0[8] ), .A3(\SB4_6/i0_0 ), 
        .ZN(\SB4_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U11270 ( .A1(\SB4_6/i0_0 ), .A2(\SB4_6/i0_3 ), .A3(\SB4_6/i0_4 ), 
        .ZN(\SB4_6/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U11272 ( .I(\SB1_4_3/buf_output[1] ), .Z(\SB2_4_31/i0[6] ) );
  NAND3_X1 U11273 ( .A1(\SB2_2_5/i0_3 ), .A2(\SB2_2_5/i0[8] ), .A3(
        \SB2_2_5/i0[9] ), .ZN(\SB2_2_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11275 ( .A1(\SB2_2_5/i0_3 ), .A2(\SB2_2_5/i0[10] ), .A3(
        \SB2_2_5/i0_4 ), .ZN(\SB2_2_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11280 ( .A1(\SB2_2_5/i0_3 ), .A2(\SB2_2_5/i0[10] ), .A3(
        \SB2_2_5/i0[9] ), .ZN(n4280) );
  NAND3_X1 U11281 ( .A1(\SB2_2_5/i0_3 ), .A2(\SB2_2_5/i0[8] ), .A3(
        \SB2_2_5/i1_7 ), .ZN(\SB2_2_5/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U11284 ( .A1(n6932), .A2(n3840), .Z(n6275) );
  AND2_X2 U11285 ( .A1(n6811), .A2(\SB1_3_30/Component_Function_4/NAND4_in[1] ), .Z(n4892) );
  AND2_X2 U11286 ( .A1(\SB1_3_30/Component_Function_4/NAND4_in[0] ), .A2(n5187), .Z(n3044) );
  NAND3_X1 U11287 ( .A1(\SB1_3_24/i1[9] ), .A2(\SB1_3_24/i0_3 ), .A3(
        \SB1_3_24/i0[6] ), .ZN(\SB1_3_24/Component_Function_3/NAND4_in[0] ) );
  CLKBUF_X8 U11288 ( .I(\RI1[4][191] ), .Z(\SB1_4_0/i0_3 ) );
  INV_X1 U11292 ( .I(\MC_ARK_ARC_1_2/buf_output[48] ), .ZN(\SB1_3_23/i3[0] )
         );
  NAND3_X1 U11293 ( .A1(\SB3_1/i1_5 ), .A2(\SB3_1/i0[6] ), .A3(\SB3_1/i0[9] ), 
        .ZN(\SB3_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U11294 ( .A1(\SB3_21/i0_0 ), .A2(\SB3_21/i0_3 ), .A3(\SB3_21/i0[7] ), .ZN(n1112) );
  NAND2_X1 U11298 ( .A1(\SB3_21/i0_0 ), .A2(\SB3_21/i3[0] ), .ZN(
        \SB3_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U11303 ( .A1(\SB3_21/i0_4 ), .A2(\SB3_21/i0_0 ), .A3(n3182), .ZN(
        \SB3_21/Component_Function_2/NAND4_in[3] ) );
  CLKBUF_X4 U11304 ( .I(\SB3_21/buf_output[5] ), .Z(\SB4_21/i0_3 ) );
  CLKBUF_X4 U11305 ( .I(\SB1_4_8/buf_output[5] ), .Z(\SB2_4_8/i0_3 ) );
  CLKBUF_X4 U11310 ( .I(\MC_ARK_ARC_1_4/buf_output[188] ), .Z(\SB3_0/i0_0 ) );
  NAND3_X1 U11311 ( .A1(\SB4_9/i0[6] ), .A2(\SB4_9/i1[9] ), .A3(\SB4_9/i0_3 ), 
        .ZN(n7050) );
  CLKBUF_X4 U11317 ( .I(\SB1_4_28/buf_output[4] ), .Z(\SB2_4_27/i0_4 ) );
  CLKBUF_X4 U11319 ( .I(\MC_ARK_ARC_1_4/buf_output[171] ), .Z(\SB3_3/i0[10] )
         );
  NAND3_X1 U11321 ( .A1(\SB3_3/i0_0 ), .A2(\SB3_3/i0[6] ), .A3(\SB3_3/i0[10] ), 
        .ZN(\SB3_3/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 U11322 ( .A1(\SB3_3/i0[10] ), .A2(\SB3_3/i0[9] ), .ZN(
        \SB3_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U11327 ( .A1(\SB3_3/i0[10] ), .A2(\SB3_3/i0_4 ), .A3(\SB3_3/i0_3 ), 
        .ZN(\SB3_3/Component_Function_0/NAND4_in[2] ) );
  INV_X1 U11329 ( .I(\SB1_4_8/buf_output[1] ), .ZN(\SB2_4_4/i1_7 ) );
  NAND3_X2 U11330 ( .A1(\SB3_25/i0[10] ), .A2(\SB3_25/i0_4 ), .A3(
        \SB3_25/i0_3 ), .ZN(\SB3_25/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U11332 ( .I(\SB1_3_27/buf_output[3] ), .Z(\SB2_3_25/i0[10] ) );
  CLKBUF_X4 U11336 ( .I(\MC_ARK_ARC_1_4/buf_output[186] ), .Z(\SB3_0/i0[9] )
         );
  NAND2_X1 U11343 ( .A1(\SB4_12/i0_3 ), .A2(\SB4_12/i1[9] ), .ZN(
        \SB4_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U11346 ( .A1(\SB4_12/i0[10] ), .A2(\SB4_12/i0_4 ), .A3(
        \SB4_12/i0_3 ), .ZN(\SB4_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11350 ( .A1(\SB3_31/i0[9] ), .A2(\SB3_31/i0_0 ), .A3(
        \SB3_31/i0[8] ), .ZN(\SB3_31/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 U11355 ( .A1(\SB3_31/i0_0 ), .A2(\SB3_31/i3[0] ), .ZN(
        \SB3_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U11357 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i0_0 ), .A3(\SB3_31/i0_4 ), 
        .ZN(\SB3_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11358 ( .A1(\SB2_4_28/i0_3 ), .A2(\SB2_4_28/i1_7 ), .A3(n4000), 
        .ZN(\SB2_4_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U11363 ( .A1(\SB4_15/i0_3 ), .A2(\SB3_17/buf_output[3] ), .A3(
        \SB4_15/i0[9] ), .ZN(n7526) );
  AND4_X2 U11364 ( .A1(\SB1_4_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_4_1/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_4_1/Component_Function_5/NAND4_in[0] ), .A4(n6385), .Z(n6277) );
  CLKBUF_X8 U11365 ( .I(\RI1[5][113] ), .Z(\SB3_13/i0_3 ) );
  NAND3_X1 U11375 ( .A1(\SB1_0_30/i1[9] ), .A2(\SB1_0_30/i1_5 ), .A3(
        \SB1_0_30/i0_4 ), .ZN(\SB1_0_30/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U11376 ( .I(\SB1_3_14/buf_output[0] ), .Z(\SB2_3_9/i0[9] ) );
  NAND3_X1 U11379 ( .A1(\SB1_4_17/i1[9] ), .A2(\SB1_4_17/i1_5 ), .A3(
        \SB1_4_17/i0_4 ), .ZN(\SB1_4_17/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U11380 ( .A1(\SB1_4_17/i0_3 ), .A2(\SB1_4_17/i1[9] ), .ZN(
        \SB1_4_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U11381 ( .A1(\SB1_4_17/i0[10] ), .A2(\SB1_4_17/i1[9] ), .A3(
        \SB1_4_17/i1_7 ), .ZN(n1037) );
  NAND2_X1 U11382 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i1[9] ), .ZN(
        \SB3_23/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 U11383 ( .A1(\SB2_4_13/i0_3 ), .A2(\SB2_4_13/i1[9] ), .ZN(
        \SB2_4_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U11385 ( .A1(\SB2_4_13/i0_3 ), .A2(\SB2_4_13/i0[10] ), .A3(
        \SB2_4_13/i0[9] ), .ZN(n4240) );
  NAND3_X1 U11387 ( .A1(\SB2_4_13/i0[7] ), .A2(\SB2_4_13/i0_3 ), .A3(
        \SB2_4_13/i0_0 ), .ZN(\SB2_4_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U11389 ( .A1(\SB2_4_13/i0_3 ), .A2(\SB2_4_13/i0[10] ), .A3(
        \SB2_4_13/i0[6] ), .ZN(n7541) );
  CLKBUF_X4 U11391 ( .I(\SB3_8/buf_output[3] ), .Z(\SB4_6/i0[10] ) );
  NAND2_X1 U11392 ( .A1(\SB2_4_11/i0_0 ), .A2(\SB2_4_11/i3[0] ), .ZN(n7321) );
  NAND3_X1 U11393 ( .A1(\SB2_4_11/i0[9] ), .A2(\SB2_4_11/i0_0 ), .A3(
        \SB2_4_11/i0[8] ), .ZN(\SB2_4_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U11400 ( .A1(\SB2_4_27/i0[9] ), .A2(\SB2_4_27/i0_3 ), .A3(
        \SB2_4_27/i0[10] ), .ZN(n7208) );
  CLKBUF_X4 U11401 ( .I(\MC_ARK_ARC_1_3/buf_output[33] ), .Z(\SB1_4_26/i0[10] ) );
  CLKBUF_X4 U11403 ( .I(\MC_ARK_ARC_1_3/buf_output[31] ), .Z(\SB1_4_26/i0[6] )
         );
  CLKBUF_X4 U11406 ( .I(\SB1_2_17/buf_output[2] ), .Z(\SB2_2_14/i0_0 ) );
  NAND3_X1 U11407 ( .A1(\SB1_3_16/i0_3 ), .A2(\SB1_3_16/i0[8] ), .A3(n1500), 
        .ZN(n7164) );
  NAND3_X1 U11409 ( .A1(\SB1_3_16/i0_0 ), .A2(\SB1_3_16/i0[8] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[90] ), .ZN(n4813) );
  NAND3_X1 U11411 ( .A1(\SB1_3_16/i0_3 ), .A2(\SB1_3_16/i1_7 ), .A3(
        \SB1_3_16/i0[8] ), .ZN(\SB1_3_16/Component_Function_1/NAND4_in[1] ) );
  INV_X1 U11412 ( .I(\RI1[5][107] ), .ZN(\SB3_14/i1_5 ) );
  CLKBUF_X12 U11417 ( .I(n295), .Z(\SB1_0_10/i0[9] ) );
  BUF_X2 U11419 ( .I(\MC_ARK_ARC_1_2/buf_output[73] ), .Z(\SB1_3_19/i0[6] ) );
  INV_X1 U11425 ( .I(\MC_ARK_ARC_1_2/buf_output[73] ), .ZN(\SB1_3_19/i1_7 ) );
  CLKBUF_X4 U11426 ( .I(\MC_ARK_ARC_1_3/buf_output[58] ), .Z(\SB1_4_22/i0_4 )
         );
  INV_X1 U11430 ( .I(\MC_ARK_ARC_1_2/buf_output[24] ), .ZN(\SB1_3_27/i3[0] )
         );
  XOR2_X1 U11431 ( .A1(\MC_ARK_ARC_1_0/temp6[5] ), .A2(n3458), .Z(n6278) );
  XOR2_X1 U11433 ( .A1(n5321), .A2(n3096), .Z(n6279) );
  NAND3_X1 U11434 ( .A1(\SB1_2_4/i0[8] ), .A2(\SB1_2_4/i3[0] ), .A3(
        \SB1_2_4/i1_5 ), .ZN(n2564) );
  NAND3_X1 U11436 ( .A1(\SB1_2_4/i0[9] ), .A2(\SB1_2_4/i0_0 ), .A3(
        \SB1_2_4/i0[8] ), .ZN(\SB1_2_4/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 U11437 ( .A1(\SB2_1_11/i0_3 ), .A2(\SB2_1_11/i1[9] ), .ZN(
        \SB2_1_11/Component_Function_1/NAND4_in[0] ) );
  CLKBUF_X4 U11439 ( .I(\MC_ARK_ARC_1_0/buf_output[87] ), .Z(\SB1_1_17/i0[10] ) );
  BUF_X4 U11442 ( .I(\SB1_1_18/buf_output[2] ), .Z(\SB2_1_15/i0_0 ) );
  NAND4_X2 U11443 ( .A1(n1523), .A2(\SB1_3_2/Component_Function_5/NAND4_in[1] ), .A3(n3961), .A4(\SB1_3_2/Component_Function_5/NAND4_in[0] ), .ZN(n6280) );
  NAND3_X1 U11445 ( .A1(\SB1_3_2/i0[6] ), .A2(\SB1_3_2/i0_3 ), .A3(
        \SB1_3_2/i1[9] ), .ZN(\SB1_3_2/Component_Function_3/NAND4_in[0] ) );
  INV_X1 U11446 ( .I(\RI3[0][95] ), .ZN(\SB2_0_16/i1_5 ) );
  NAND3_X1 U11449 ( .A1(\SB2_1_2/i0[10] ), .A2(\SB2_1_2/i0_4 ), .A3(
        \SB2_1_2/i0_3 ), .ZN(\SB2_1_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11450 ( .A1(\SB1_2_24/i0[8] ), .A2(\SB1_2_24/i0[7] ), .A3(
        \SB1_2_24/i0[6] ), .ZN(\SB1_2_24/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U11451 ( .A1(\SB1_1_30/i0[8] ), .A2(\SB1_1_30/i0[7] ), .A3(
        \SB1_1_30/i0[6] ), .ZN(\SB1_1_30/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U11452 ( .A1(Key[158]), .A2(Plaintext[158]), .Z(n6281) );
  AND4_X2 U11453 ( .A1(\SB1_0_5/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_5/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_5/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_5/Component_Function_5/NAND4_in[3] ), .Z(n6282) );
  AND4_X2 U11457 ( .A1(\SB1_1_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_24/Component_Function_3/NAND4_in[3] ), .A3(n1833), .A4(n6368), 
        .Z(n6283) );
  AND4_X2 U11458 ( .A1(\SB2_1_22/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_22/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_22/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_1_22/Component_Function_2/NAND4_in[2] ), .Z(n6284) );
  INV_X4 U11459 ( .I(n6284), .ZN(\SB2_1_22/buf_output[2] ) );
  NAND3_X1 U11465 ( .A1(\SB1_2_25/i0[10] ), .A2(\SB1_2_25/i1[9] ), .A3(
        \SB1_2_25/i1_5 ), .ZN(\SB1_2_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U11468 ( .A1(\SB1_2_25/i0_4 ), .A2(\SB1_2_25/i1[9] ), .A3(
        \SB1_2_25/i1_5 ), .ZN(n7588) );
  NAND3_X1 U11469 ( .A1(\SB1_2_25/i1[9] ), .A2(\SB1_2_25/i0_4 ), .A3(
        \SB1_2_25/i0_3 ), .ZN(\SB1_2_25/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U11470 ( .I(\MC_ARK_ARC_1_1/buf_output[159] ), .Z(\SB1_2_5/i0[10] ) );
  XOR2_X1 U11472 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[164] ), .A2(\RI5[2][188] ), .Z(n6285) );
  BUF_X2 U11476 ( .I(\MC_ARK_ARC_1_4/buf_output[135] ), .Z(\SB3_9/i0[10] ) );
  INV_X1 U11477 ( .I(\MC_ARK_ARC_1_4/buf_output[135] ), .ZN(\SB3_9/i0[8] ) );
  XOR2_X1 U11479 ( .A1(n4894), .A2(n7233), .Z(n6286) );
  NAND3_X1 U11480 ( .A1(\SB4_9/i0[6] ), .A2(\SB4_9/i0[10] ), .A3(\SB4_9/i0_3 ), 
        .ZN(n5025) );
  BUF_X2 U11483 ( .I(\MC_ARK_ARC_1_0/buf_output[120] ), .Z(\SB1_1_11/i0[9] )
         );
  INV_X1 U11484 ( .I(\MC_ARK_ARC_1_0/buf_output[120] ), .ZN(\SB1_1_11/i3[0] )
         );
  CLKBUF_X4 U11490 ( .I(\MC_ARK_ARC_1_3/buf_output[20] ), .Z(\SB1_4_28/i0_0 )
         );
  INV_X1 U11492 ( .I(\SB3_11/buf_output[0] ), .ZN(\SB4_6/i3[0] ) );
  BUF_X2 U11493 ( .I(\SB3_11/buf_output[0] ), .Z(\SB4_6/i0[9] ) );
  CLKBUF_X4 U11498 ( .I(\MC_ARK_ARC_1_1/buf_output[143] ), .Z(\SB1_2_8/i0_3 )
         );
  INV_X1 U11503 ( .I(\MC_ARK_ARC_1_1/buf_output[143] ), .ZN(\SB1_2_8/i1_5 ) );
  NAND3_X2 U11506 ( .A1(\SB1_4_3/i0[9] ), .A2(\SB1_4_3/i0_4 ), .A3(
        \SB1_4_3/i0[6] ), .ZN(n2584) );
  BUF_X4 U11511 ( .I(\SB2_4_11/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_4/buf_datainput[135] ) );
  CLKBUF_X4 U11522 ( .I(\MC_ARK_ARC_1_0/buf_output[27] ), .Z(\SB1_1_27/i0[10] ) );
  CLKBUF_X4 U11523 ( .I(\MC_ARK_ARC_1_1/buf_output[92] ), .Z(\SB1_2_16/i0_0 )
         );
  INV_X1 U11525 ( .I(\SB3_13/buf_output[1] ), .ZN(\SB4_9/i1_7 ) );
  AND2_X2 U11530 ( .A1(\MC_ARK_ARC_1_4/buf_output[40] ), .A2(n6287), .Z(n774)
         );
  CLKBUF_X4 U11531 ( .I(\SB3_25/buf_output[4] ), .Z(\SB4_24/i0_4 ) );
  NAND4_X2 U11532 ( .A1(\SB1_0_25/Component_Function_2/NAND4_in[0] ), .A2(
        n2323), .A3(n3303), .A4(\SB1_0_25/Component_Function_2/NAND4_in[3] ), 
        .ZN(n6288) );
  XOR2_X1 U11542 ( .A1(\MC_ARK_ARC_1_1/temp6[107] ), .A2(n961), .Z(n6289) );
  CLKBUF_X4 U11546 ( .I(n280), .Z(n6290) );
  XOR2_X1 U11547 ( .A1(n3344), .A2(n3343), .Z(n6291) );
  XOR2_X1 U11551 ( .A1(n6292), .A2(\MC_ARK_ARC_1_4/temp4[68] ), .Z(
        \MC_ARK_ARC_1_4/temp6[68] ) );
  XOR2_X1 U11553 ( .A1(\RI5[4][134] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[170] ), .Z(n6292) );
  NAND4_X2 U11554 ( .A1(\SB2_4_7/Component_Function_5/NAND4_in[0] ), .A2(n4845), .A3(n988), .A4(n6293), .ZN(\SB2_4_7/buf_output[5] ) );
  NAND3_X2 U11555 ( .A1(\SB2_4_7/i0_0 ), .A2(\SB2_4_7/i0[10] ), .A3(
        \SB2_4_7/i0[6] ), .ZN(n6293) );
  NAND3_X1 U11558 ( .A1(\SB2_3_13/i0_0 ), .A2(\SB2_3_13/i0[10] ), .A3(
        \SB1_3_17/buf_output[1] ), .ZN(
        \SB2_3_13/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U11559 ( .A1(n6295), .A2(n6294), .Z(\MC_ARK_ARC_1_3/temp6[5] ) );
  XOR2_X1 U11561 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[71] ), .A2(n118), .Z(
        n6294) );
  XOR2_X1 U11562 ( .A1(\RI5[3][107] ), .A2(\RI5[3][41] ), .Z(n6295) );
  XOR2_X1 U11563 ( .A1(n6297), .A2(n4362), .Z(n2518) );
  XOR2_X1 U11565 ( .A1(\RI5[0][83] ), .A2(\RI5[0][107] ), .Z(n6297) );
  NAND4_X2 U11566 ( .A1(\SB2_2_6/Component_Function_5/NAND4_in[2] ), .A2(n4417), .A3(n7060), .A4(\SB2_2_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_6/buf_output[5] ) );
  XOR2_X1 U11567 ( .A1(n1339), .A2(n6299), .Z(n1764) );
  XOR2_X1 U11568 ( .A1(\RI5[4][56] ), .A2(\RI5[4][62] ), .Z(n6299) );
  XOR2_X1 U11578 ( .A1(n4058), .A2(n6300), .Z(\MC_ARK_ARC_1_1/temp5[170] ) );
  INV_X2 U11582 ( .I(\RI3[0][170] ), .ZN(\SB2_0_3/i1[9] ) );
  NAND4_X2 U11583 ( .A1(n1749), .A2(n2079), .A3(n2918), .A4(
        \SB1_0_6/Component_Function_2/NAND4_in[2] ), .ZN(\RI3[0][170] ) );
  NAND4_X2 U11588 ( .A1(\SB1_1_3/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_3/Component_Function_2/NAND4_in[0] ), .A3(n2021), .A4(n6301), 
        .ZN(\SB1_1_3/buf_output[2] ) );
  NAND3_X2 U11589 ( .A1(\SB1_1_3/i0_0 ), .A2(\SB1_1_3/i0_4 ), .A3(
        \SB1_1_3/i1_5 ), .ZN(n6301) );
  NAND3_X1 U11592 ( .A1(\SB4_21/i0_4 ), .A2(\SB3_24/buf_output[2] ), .A3(
        \SB4_21/i1_5 ), .ZN(\SB4_21/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U11593 ( .A1(n6302), .A2(n7369), .Z(\MC_ARK_ARC_1_1/buf_output[132] ) );
  XOR2_X1 U11595 ( .A1(\MC_ARK_ARC_1_1/temp4[132] ), .A2(
        \MC_ARK_ARC_1_1/temp3[132] ), .Z(n6302) );
  XOR2_X1 U11596 ( .A1(\MC_ARK_ARC_1_0/temp2[56] ), .A2(n7002), .Z(n6303) );
  NAND4_X2 U11598 ( .A1(\SB1_3_16/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_16/Component_Function_1/NAND4_in[0] ), .A4(n6304), .ZN(
        \SB1_3_16/buf_output[1] ) );
  XOR2_X1 U11599 ( .A1(\MC_ARK_ARC_1_2/temp6[185] ), .A2(n6305), .Z(
        \MC_ARK_ARC_1_2/buf_output[185] ) );
  XOR2_X1 U11602 ( .A1(\MC_ARK_ARC_1_2/temp2[185] ), .A2(
        \MC_ARK_ARC_1_2/temp1[185] ), .Z(n6305) );
  NAND2_X1 U11610 ( .A1(\SB2_1_26/i0[9] ), .A2(\SB2_1_26/i0[10] ), .ZN(n6306)
         );
  NAND3_X1 U11613 ( .A1(\SB1_1_5/i0_0 ), .A2(\SB1_1_5/i1_7 ), .A3(
        \SB1_1_5/i3[0] ), .ZN(\SB1_1_5/Component_Function_4/NAND4_in[1] ) );
  INV_X2 U11614 ( .I(\SB1_3_29/buf_output[2] ), .ZN(\SB2_3_26/i1[9] ) );
  NAND3_X1 U11618 ( .A1(\SB1_2_23/i0_3 ), .A2(\SB1_2_23/i0[9] ), .A3(
        \SB1_2_23/i0[8] ), .ZN(\SB1_2_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U11623 ( .A1(\SB2_2_9/i0[10] ), .A2(\SB2_2_9/i1[9] ), .A3(
        \SB2_2_9/i1_7 ), .ZN(\SB2_2_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U11624 ( .A1(\SB1_2_18/i0[10] ), .A2(\SB1_2_18/i0_0 ), .A3(
        \SB1_2_18/i0[6] ), .ZN(\SB1_2_18/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U11625 ( .A1(\SB1_0_10/i0[9] ), .A2(\SB1_0_10/i0[8] ), .A3(
        \SB1_0_10/i0_0 ), .ZN(\SB1_0_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U11626 ( .A1(\SB2_3_12/i3[0] ), .A2(\SB2_3_12/i1_5 ), .A3(
        \SB2_3_12/i0[8] ), .ZN(\SB2_3_12/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U11628 ( .A1(n6307), .A2(n185), .Z(Ciphertext[71]) );
  NAND4_X2 U11630 ( .A1(\SB4_20/Component_Function_5/NAND4_in[2] ), .A2(n2700), 
        .A3(\SB4_20/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_20/Component_Function_5/NAND4_in[0] ), .ZN(n6307) );
  XOR2_X1 U11631 ( .A1(\RI5[2][175] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .Z(n2305) );
  NAND4_X2 U11632 ( .A1(\SB1_4_10/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_4_10/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_4_10/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_4_10/Component_Function_5/NAND4_in[2] ), .ZN(
        \SB1_4_10/buf_output[5] ) );
  NAND4_X2 U11635 ( .A1(\SB1_1_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_28/Component_Function_0/NAND4_in[0] ), .A3(n6542), .A4(n2430), 
        .ZN(\SB1_1_28/buf_output[0] ) );
  NAND4_X2 U11636 ( .A1(\SB2_4_10/Component_Function_2/NAND4_in[3] ), .A2(n788), .A3(n6787), .A4(n6308), .ZN(\SB2_4_10/buf_output[2] ) );
  NAND4_X2 U11639 ( .A1(n3422), .A2(n6621), .A3(n6474), .A4(
        \SB1_1_24/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_24/buf_output[5] ) );
  XOR2_X1 U11642 ( .A1(\MC_ARK_ARC_1_2/temp5[20] ), .A2(n6309), .Z(
        \MC_ARK_ARC_1_2/buf_output[20] ) );
  XOR2_X1 U11643 ( .A1(n3775), .A2(n3774), .Z(n6309) );
  NAND4_X2 U11644 ( .A1(\SB1_2_6/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_6/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_6/Component_Function_4/NAND4_in[2] ), .A4(n6310), .ZN(
        \SB1_2_6/buf_output[4] ) );
  NAND3_X2 U11645 ( .A1(\SB1_3_11/i0[10] ), .A2(\SB1_3_11/i1[9] ), .A3(
        \SB1_3_11/i1_5 ), .ZN(n6557) );
  NAND4_X2 U11647 ( .A1(\SB2_0_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_9/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_0_9/Component_Function_2/NAND4_in[1] ), .A4(n5119), .ZN(
        \SB2_0_9/buf_output[2] ) );
  NAND4_X2 U11648 ( .A1(n2522), .A2(\SB4_3/Component_Function_5/NAND4_in[2] ), 
        .A3(\SB4_3/Component_Function_5/NAND4_in[3] ), .A4(n6311), .ZN(n6409)
         );
  NAND2_X2 U11649 ( .A1(\SB4_3/i0_0 ), .A2(\SB4_3/i3[0] ), .ZN(n6311) );
  XOR2_X1 U11651 ( .A1(\RI5[3][26] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[62] ), 
        .Z(n2013) );
  XOR2_X1 U11652 ( .A1(\MC_ARK_ARC_1_3/temp2[18] ), .A2(n6312), .Z(n4461) );
  XOR2_X1 U11653 ( .A1(\RI5[3][12] ), .A2(\RI5[3][18] ), .Z(n6312) );
  NAND4_X2 U11657 ( .A1(\SB1_3_4/Component_Function_4/NAND4_in[1] ), .A2(n1411), .A3(n2786), .A4(n6313), .ZN(\SB1_3_4/buf_output[4] ) );
  NAND3_X2 U11658 ( .A1(\SB1_3_4/i0[9] ), .A2(\SB1_3_4/i0_0 ), .A3(
        \SB1_3_4/i0[8] ), .ZN(n6313) );
  XOR2_X1 U11660 ( .A1(\RI5[4][137] ), .A2(\RI5[4][161] ), .Z(n4175) );
  NAND3_X1 U11664 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i0_3 ), .A3(
        \SB1_3_2/i0_4 ), .ZN(\SB1_3_2/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U11665 ( .A1(\MC_ARK_ARC_1_3/temp3[69] ), .A2(
        \MC_ARK_ARC_1_3/temp4[69] ), .Z(n7532) );
  NAND4_X2 U11666 ( .A1(\SB2_2_11/Component_Function_2/NAND4_in[0] ), .A2(
        n4549), .A3(\SB2_2_11/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_11/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_2_11/buf_output[2] ) );
  NAND4_X2 U11671 ( .A1(n641), .A2(n6348), .A3(
        \SB2_2_6/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_2_6/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_2_6/buf_output[4] ) );
  NAND4_X2 U11674 ( .A1(n3161), .A2(n6717), .A3(
        \SB2_1_23/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_23/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_23/buf_output[5] ) );
  XOR2_X1 U11678 ( .A1(n6314), .A2(\MC_ARK_ARC_1_2/temp6[162] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[162] ) );
  XOR2_X1 U11680 ( .A1(\MC_ARK_ARC_1_2/temp2[162] ), .A2(n5089), .Z(n6314) );
  XOR2_X1 U11681 ( .A1(n3953), .A2(n6315), .Z(\MC_ARK_ARC_1_2/buf_output[41] )
         );
  XOR2_X1 U11685 ( .A1(\RI5[2][117] ), .A2(\RI5[2][153] ), .Z(
        \MC_ARK_ARC_1_2/temp3[51] ) );
  NAND4_X2 U11686 ( .A1(n4448), .A2(n1650), .A3(n6635), .A4(n4038), .ZN(
        \SB2_2_8/buf_output[3] ) );
  NAND4_X2 U11692 ( .A1(\SB2_3_1/Component_Function_1/NAND4_in[1] ), .A2(n3674), .A3(\SB2_3_1/Component_Function_1/NAND4_in[0] ), .A4(n6316), .ZN(
        \SB2_3_1/buf_output[1] ) );
  NAND3_X1 U11693 ( .A1(\SB2_3_1/i0_4 ), .A2(\SB2_3_1/i1_7 ), .A3(
        \SB2_3_1/i0[8] ), .ZN(n6316) );
  NAND4_X2 U11695 ( .A1(\SB1_3_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_2/Component_Function_4/NAND4_in[3] ), .A4(n6318), .ZN(
        \SB1_3_2/buf_output[4] ) );
  NAND3_X1 U11697 ( .A1(\SB1_3_2/i0_3 ), .A2(\SB1_3_2/i0[10] ), .A3(
        \SB1_3_2/i0[9] ), .ZN(n6318) );
  XOR2_X1 U11698 ( .A1(\RI5[0][117] ), .A2(\RI5[0][93] ), .Z(n6319) );
  XOR2_X1 U11701 ( .A1(n7271), .A2(n6320), .Z(\MC_ARK_ARC_1_1/temp5[135] ) );
  XOR2_X1 U11702 ( .A1(\RI5[1][81] ), .A2(\RI5[1][105] ), .Z(n6320) );
  XOR2_X1 U11703 ( .A1(\MC_ARK_ARC_1_1/temp2[156] ), .A2(n6321), .Z(
        \MC_ARK_ARC_1_1/temp5[156] ) );
  XOR2_X1 U11704 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[150] ), .A2(\RI5[1][156] ), .Z(n6321) );
  XOR2_X1 U11708 ( .A1(\RI5[1][143] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[83] ), 
        .Z(n6322) );
  XOR2_X1 U11710 ( .A1(\MC_ARK_ARC_1_2/temp2[140] ), .A2(n6323), .Z(
        \MC_ARK_ARC_1_2/temp5[140] ) );
  XOR2_X1 U11711 ( .A1(\RI5[2][134] ), .A2(\RI5[2][140] ), .Z(n6323) );
  XOR2_X1 U11712 ( .A1(n6325), .A2(n6324), .Z(n3063) );
  XOR2_X1 U11713 ( .A1(\RI5[4][83] ), .A2(n53), .Z(n6324) );
  XOR2_X1 U11715 ( .A1(\RI5[4][17] ), .A2(\RI5[4][47] ), .Z(n6325) );
  NAND2_X2 U11717 ( .A1(n7155), .A2(n6326), .ZN(\RI5[3][91] ) );
  AND2_X1 U11718 ( .A1(\SB2_3_20/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_20/Component_Function_1/NAND4_in[3] ), .Z(n6326) );
  NAND4_X2 U11725 ( .A1(\SB1_2_11/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_2_11/Component_Function_4/NAND4_in[1] ), .A3(n1244), .A4(n6327), 
        .ZN(\SB1_2_11/buf_output[4] ) );
  NAND3_X2 U11726 ( .A1(\SB1_2_11/i0[9] ), .A2(\SB1_2_11/i0[8] ), .A3(
        \SB1_2_11/i0_0 ), .ZN(n6327) );
  XOR2_X1 U11729 ( .A1(n6329), .A2(n6328), .Z(\MC_ARK_ARC_1_4/temp6[92] ) );
  XOR2_X1 U11730 ( .A1(\SB2_4_8/buf_output[2] ), .A2(n522), .Z(n6328) );
  XOR2_X1 U11732 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[2] ), .A2(\RI5[4][128] ), 
        .Z(n6329) );
  NAND4_X2 U11736 ( .A1(\SB2_4_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_2/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_4_2/Component_Function_2/NAND4_in[1] ), .A4(n6330), .ZN(
        \SB2_4_2/buf_output[2] ) );
  NAND3_X2 U11738 ( .A1(\SB2_4_2/i0[9] ), .A2(\SB2_4_2/i0_3 ), .A3(
        \SB2_4_2/i0[8] ), .ZN(n6330) );
  NAND4_X2 U11741 ( .A1(n1375), .A2(n1662), .A3(
        \SB1_1_3/Component_Function_1/NAND4_in[0] ), .A4(n6331), .ZN(
        \SB1_1_3/buf_output[1] ) );
  NAND3_X2 U11744 ( .A1(\SB1_1_3/i0_3 ), .A2(\SB1_1_3/i0[8] ), .A3(
        \SB1_1_3/i1_7 ), .ZN(n6331) );
  XOR2_X1 U11745 ( .A1(n6419), .A2(n6332), .Z(\MC_ARK_ARC_1_4/temp5[152] ) );
  XOR2_X1 U11746 ( .A1(\SB2_4_9/buf_output[2] ), .A2(\RI5[4][146] ), .Z(n6332)
         );
  XOR2_X1 U11750 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[117] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_4/temp2[171] )
         );
  XOR2_X1 U11751 ( .A1(n6333), .A2(n125), .Z(Ciphertext[191]) );
  NAND4_X2 U11753 ( .A1(\SB4_0/Component_Function_5/NAND4_in[2] ), .A2(n3936), 
        .A3(\SB4_0/Component_Function_5/NAND4_in[0] ), .A4(
        \SB4_0/Component_Function_5/NAND4_in[3] ), .ZN(n6333) );
  XOR2_X1 U11756 ( .A1(\MC_ARK_ARC_1_2/temp2[146] ), .A2(n6334), .Z(n1546) );
  XOR2_X1 U11757 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), .A2(\RI5[2][140] ), .Z(n6334) );
  XOR2_X1 U11761 ( .A1(\RI5[1][91] ), .A2(\RI5[1][115] ), .Z(n6335) );
  XOR2_X1 U11762 ( .A1(\MC_ARK_ARC_1_2/temp4[101] ), .A2(n6336), .Z(n6450) );
  XOR2_X1 U11766 ( .A1(\RI5[2][167] ), .A2(\RI5[2][11] ), .Z(n6336) );
  XOR2_X1 U11768 ( .A1(\RI5[1][169] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .Z(n6337) );
  INV_X2 U11769 ( .I(\SB1_4_23/buf_output[2] ), .ZN(\SB2_4_20/i1[9] ) );
  NAND4_X2 U11770 ( .A1(\SB1_4_23/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_4_23/Component_Function_2/NAND4_in[3] ), .A3(n7016), .A4(
        \SB1_4_23/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_4_23/buf_output[2] ) );
  XOR2_X1 U11771 ( .A1(\MC_ARK_ARC_1_2/temp1[14] ), .A2(n6339), .Z(n7262) );
  XOR2_X1 U11777 ( .A1(\SB2_2_5/buf_output[2] ), .A2(\RI5[2][152] ), .Z(n6339)
         );
  XOR2_X1 U11778 ( .A1(\RI5[1][12] ), .A2(\RI5[1][180] ), .Z(n2687) );
  XOR2_X1 U11781 ( .A1(n6340), .A2(n4342), .Z(\MC_ARK_ARC_1_2/temp5[53] ) );
  XOR2_X1 U11782 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[23] ), .A2(\RI5[2][53] ), 
        .Z(n6340) );
  XOR2_X1 U11783 ( .A1(\MC_ARK_ARC_1_1/temp6[20] ), .A2(n6341), .Z(
        \MC_ARK_ARC_1_1/buf_output[20] ) );
  XOR2_X1 U11784 ( .A1(n4299), .A2(n3252), .Z(n6341) );
  NAND3_X2 U11785 ( .A1(n600), .A2(\SB2_2_23/i0_0 ), .A3(\SB2_2_23/i1_5 ), 
        .ZN(n6342) );
  NAND3_X1 U11788 ( .A1(\SB1_1_27/i1_7 ), .A2(\SB1_1_27/i0_0 ), .A3(
        \SB1_1_27/i3[0] ), .ZN(\SB1_1_27/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U11789 ( .A1(\SB2_2_24/Component_Function_5/NAND4_in[2] ), .A2(
        n1962), .A3(\SB2_2_24/Component_Function_5/NAND4_in[0] ), .A4(n6343), 
        .ZN(\SB2_2_24/buf_output[5] ) );
  XOR2_X1 U11791 ( .A1(\SB2_2_11/buf_output[5] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[89] ), .Z(\MC_ARK_ARC_1_2/temp3[23] ) );
  XOR2_X1 U11795 ( .A1(\MC_ARK_ARC_1_1/temp1[92] ), .A2(n6344), .Z(n6366) );
  XOR2_X1 U11800 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[62] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[38] ), .Z(n6344) );
  XOR2_X1 U11803 ( .A1(\RI5[2][176] ), .A2(\RI5[2][8] ), .Z(n2555) );
  XOR2_X1 U11804 ( .A1(\MC_ARK_ARC_1_1/temp5[96] ), .A2(n6345), .Z(
        \MC_ARK_ARC_1_1/buf_output[96] ) );
  XOR2_X1 U11809 ( .A1(\MC_ARK_ARC_1_1/temp3[96] ), .A2(
        \MC_ARK_ARC_1_1/temp4[96] ), .Z(n6345) );
  NAND3_X2 U11810 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0[8] ), .A3(
        \SB2_2_1/i0[9] ), .ZN(\SB2_2_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11814 ( .A1(\SB1_3_22/i0_0 ), .A2(\MC_ARK_ARC_1_2/buf_output[58] ), 
        .A3(\SB1_3_22/i1_5 ), .ZN(\SB1_3_22/Component_Function_2/NAND4_in[3] )
         );
  NAND3_X2 U11817 ( .A1(\SB1_1_5/i0_3 ), .A2(\SB1_1_5/i1[9] ), .A3(
        \SB1_1_5/i0_4 ), .ZN(n4442) );
  INV_X8 U11824 ( .I(n6346), .ZN(\RI1[2][59] ) );
  INV_X2 U11827 ( .I(\MC_ARK_ARC_1_1/buf_output[59] ), .ZN(n6346) );
  NAND3_X1 U11829 ( .A1(\SB4_21/i0_4 ), .A2(n3998), .A3(\SB4_21/i1_5 ), .ZN(
        \SB4_21/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U11830 ( .A1(n4213), .A2(n4451), .A3(n6682), .A4(
        \SB1_4_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_4_29/buf_output[5] ) );
  NAND4_X2 U11831 ( .A1(\SB1_3_29/Component_Function_3/NAND4_in[0] ), .A2(
        n4601), .A3(\SB1_3_29/Component_Function_3/NAND4_in[1] ), .A4(n3756), 
        .ZN(\SB1_3_29/buf_output[3] ) );
  NAND3_X1 U11832 ( .A1(\SB4_24/i0_4 ), .A2(\SB3_26/buf_output[3] ), .A3(
        \SB4_24/i0_3 ), .ZN(\SB4_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U11836 ( .A1(\SB2_3_27/i0[10] ), .A2(\SB2_3_27/i0[6] ), .A3(
        \SB2_3_27/i0_0 ), .ZN(\SB2_3_27/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U11837 ( .A1(\RI5[0][98] ), .A2(\RI5[0][62] ), .Z(
        \MC_ARK_ARC_1_0/temp3[188] ) );
  NAND2_X2 U11838 ( .A1(n5425), .A2(n6347), .ZN(\RI5[4][116] ) );
  XOR2_X1 U11840 ( .A1(\RI5[0][168] ), .A2(\RI5[0][144] ), .Z(
        \MC_ARK_ARC_1_0/temp2[6] ) );
  INV_X2 U11842 ( .I(\SB1_1_26/buf_output[2] ), .ZN(\SB2_1_23/i1[9] ) );
  NAND4_X2 U11844 ( .A1(n4614), .A2(
        \SB1_1_26/Component_Function_2/NAND4_in[2] ), .A3(n6440), .A4(n4816), 
        .ZN(\SB1_1_26/buf_output[2] ) );
  NAND4_X2 U11845 ( .A1(\SB1_4_17/Component_Function_3/NAND4_in[1] ), .A2(
        n1037), .A3(n5373), .A4(n6349), .ZN(\SB1_4_17/buf_output[3] ) );
  NAND4_X2 U11846 ( .A1(\SB1_3_2/Component_Function_3/NAND4_in[0] ), .A2(n4511), .A3(n3523), .A4(n6350), .ZN(\SB1_3_2/buf_output[3] ) );
  NAND3_X2 U11849 ( .A1(\SB1_3_2/i3[0] ), .A2(\SB1_3_2/i0[8] ), .A3(
        \SB1_3_2/i1_5 ), .ZN(n6350) );
  NAND4_X2 U11852 ( .A1(\SB1_2_26/Component_Function_4/NAND4_in[3] ), .A2(
        n7358), .A3(\SB1_2_26/Component_Function_4/NAND4_in[1] ), .A4(n6351), 
        .ZN(\SB1_2_26/buf_output[4] ) );
  NAND3_X2 U11854 ( .A1(\SB1_2_26/i0[9] ), .A2(\SB1_2_26/i0[8] ), .A3(
        \SB1_2_26/i0_0 ), .ZN(n6351) );
  XOR2_X1 U11858 ( .A1(n6352), .A2(\MC_ARK_ARC_1_1/temp1[28] ), .Z(
        \MC_ARK_ARC_1_1/temp5[28] ) );
  XOR2_X1 U11859 ( .A1(\RI5[1][166] ), .A2(\RI5[1][190] ), .Z(n6352) );
  XOR2_X1 U11861 ( .A1(\MC_ARK_ARC_1_3/temp4[150] ), .A2(n6353), .Z(
        \MC_ARK_ARC_1_3/temp6[150] ) );
  XOR2_X1 U11862 ( .A1(\RI5[3][60] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[24] ), 
        .Z(n6353) );
  XOR2_X1 U11864 ( .A1(\RI5[1][17] ), .A2(\RI5[1][185] ), .Z(
        \MC_ARK_ARC_1_1/temp2[47] ) );
  NAND4_X2 U11865 ( .A1(\SB2_1_25/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_25/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_25/Component_Function_4/NAND4_in[2] ), .A4(n6354), .ZN(
        \SB2_1_25/buf_output[4] ) );
  NAND3_X1 U11868 ( .A1(\SB2_1_25/i0_4 ), .A2(\SB2_1_25/i1[9] ), .A3(
        \SB2_1_25/i1_5 ), .ZN(n6354) );
  XOR2_X1 U11869 ( .A1(\MC_ARK_ARC_1_3/temp1[136] ), .A2(n6355), .Z(
        \MC_ARK_ARC_1_3/temp5[136] ) );
  XOR2_X1 U11870 ( .A1(\RI5[3][106] ), .A2(\RI5[3][82] ), .Z(n6355) );
  XOR2_X1 U11872 ( .A1(\MC_ARK_ARC_1_0/temp5[64] ), .A2(n6356), .Z(
        \MC_ARK_ARC_1_0/buf_output[64] ) );
  XOR2_X1 U11873 ( .A1(\MC_ARK_ARC_1_0/temp4[64] ), .A2(
        \MC_ARK_ARC_1_0/temp3[64] ), .Z(n6356) );
  NAND4_X2 U11876 ( .A1(n2105), .A2(
        \SB2_2_29/Component_Function_2/NAND4_in[0] ), .A3(n3864), .A4(n6357), 
        .ZN(\SB2_2_29/buf_output[2] ) );
  NAND3_X2 U11877 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0[6] ), .A3(
        \SB2_2_29/i0[10] ), .ZN(n6357) );
  NAND3_X2 U11879 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0[9] ), .A3(
        \SB2_3_15/i0[10] ), .ZN(n1995) );
  XOR2_X1 U11884 ( .A1(\MC_ARK_ARC_1_2/temp4[99] ), .A2(n6358), .Z(n7244) );
  XOR2_X1 U11885 ( .A1(\RI5[2][165] ), .A2(\RI5[2][9] ), .Z(n6358) );
  NAND4_X2 U11886 ( .A1(\SB1_2_4/Component_Function_5/NAND4_in[2] ), .A2(n3575), .A3(\SB1_2_4/Component_Function_5/NAND4_in[0] ), .A4(n6359), .ZN(
        \SB1_2_4/buf_output[5] ) );
  NAND3_X2 U11892 ( .A1(\SB1_2_4/i0[6] ), .A2(\SB1_2_4/i0[9] ), .A3(
        \SB1_2_4/i0_4 ), .ZN(n6359) );
  NAND4_X2 U11893 ( .A1(\SB2_1_3/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_3/Component_Function_0/NAND4_in[3] ), .A4(n6360), .ZN(
        \SB2_1_3/buf_output[0] ) );
  NAND2_X1 U11895 ( .A1(\SB2_1_3/i0[9] ), .A2(\SB2_1_3/i0[10] ), .ZN(n6360) );
  XOR2_X1 U11898 ( .A1(n5282), .A2(n6361), .Z(\MC_ARK_ARC_1_2/buf_output[56] )
         );
  XOR2_X1 U11900 ( .A1(\MC_ARK_ARC_1_1/temp4[8] ), .A2(
        \MC_ARK_ARC_1_1/temp3[8] ), .Z(n6362) );
  XOR2_X1 U11902 ( .A1(n6364), .A2(n6363), .Z(\MC_ARK_ARC_1_1/temp6[135] ) );
  XOR2_X1 U11906 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[45] ), .A2(n466), .Z(
        n6363) );
  XOR2_X1 U11907 ( .A1(\RI5[1][9] ), .A2(\RI5[1][171] ), .Z(n6364) );
  XOR2_X1 U11912 ( .A1(n3025), .A2(\MC_ARK_ARC_1_3/temp6[129] ), .Z(n1491) );
  XOR2_X1 U11913 ( .A1(\MC_ARK_ARC_1_3/temp4[129] ), .A2(
        \MC_ARK_ARC_1_3/temp3[129] ), .Z(\MC_ARK_ARC_1_3/temp6[129] ) );
  NAND3_X2 U11915 ( .A1(\SB1_4_27/i1[9] ), .A2(\SB1_4_27/i0_3 ), .A3(
        \SB1_4_27/i0_4 ), .ZN(\SB1_4_27/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U11916 ( .A1(n6365), .A2(n141), .Z(Ciphertext[99]) );
  NAND4_X2 U11917 ( .A1(n2027), .A2(\SB4_15/Component_Function_3/NAND4_in[3] ), 
        .A3(\SB4_15/Component_Function_3/NAND4_in[1] ), .A4(n2663), .ZN(n6365)
         );
  NAND3_X2 U11921 ( .A1(\SB1_0_21/i0[8] ), .A2(\SB1_0_21/i1_5 ), .A3(
        \SB1_0_21/i3[0] ), .ZN(\SB1_0_21/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U11925 ( .A1(n6366), .A2(\MC_ARK_ARC_1_1/temp6[92] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[92] ) );
  XOR2_X1 U11927 ( .A1(n6367), .A2(\MC_ARK_ARC_1_0/temp4[68] ), .Z(n1548) );
  XOR2_X1 U11928 ( .A1(\RI5[0][38] ), .A2(\RI5[0][14] ), .Z(n6367) );
  NAND4_X2 U11936 ( .A1(\SB1_1_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_24/Component_Function_3/NAND4_in[3] ), .A3(n1833), .A4(n6368), 
        .ZN(\SB1_1_24/buf_output[3] ) );
  NAND3_X2 U11939 ( .A1(\SB1_1_24/i0_4 ), .A2(\RI1[1][47] ), .A3(
        \SB1_1_24/i0_0 ), .ZN(n6368) );
  NAND3_X2 U11940 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB2_3_7/i0_4 ), .A3(
        \SB2_3_7/i0_0 ), .ZN(n7576) );
  NAND4_X2 U11941 ( .A1(\SB2_1_19/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_19/Component_Function_4/NAND4_in[0] ), .A3(n4200), .A4(
        \SB2_1_19/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_1_19/buf_output[4] ) );
  NAND4_X2 U11943 ( .A1(\SB2_2_14/Component_Function_5/NAND4_in[1] ), .A2(
        n3114), .A3(n3317), .A4(\SB2_2_14/Component_Function_5/NAND4_in[0] ), 
        .ZN(\SB2_2_14/buf_output[5] ) );
  XOR2_X1 U11944 ( .A1(\SB2_3_28/buf_output[1] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[37] ), .Z(\MC_ARK_ARC_1_3/temp1[43] ) );
  NAND4_X2 U11947 ( .A1(n4325), .A2(
        \SB2_0_14/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_0_14/Component_Function_3/NAND4_in[0] ), .A4(
        \SB2_0_14/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_14/buf_output[3] ) );
  XOR2_X1 U11950 ( .A1(\MC_ARK_ARC_1_4/temp5[92] ), .A2(
        \MC_ARK_ARC_1_4/temp6[92] ), .Z(\MC_ARK_ARC_1_4/buf_output[92] ) );
  NAND4_X2 U11952 ( .A1(\SB1_3_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_31/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_3_31/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_3_31/buf_output[3] ) );
  XOR2_X1 U11956 ( .A1(\MC_ARK_ARC_1_0/temp6[46] ), .A2(
        \MC_ARK_ARC_1_0/temp5[46] ), .Z(\MC_ARK_ARC_1_0/buf_output[46] ) );
  NAND4_X2 U11959 ( .A1(n2561), .A2(
        \SB2_4_15/Component_Function_5/NAND4_in[3] ), .A3(n6549), .A4(n6551), 
        .ZN(\SB2_4_15/buf_output[5] ) );
  XOR2_X1 U11960 ( .A1(n4534), .A2(n5375), .Z(\MC_ARK_ARC_1_2/buf_output[145] ) );
  INV_X8 U11965 ( .I(n6369), .ZN(\RI1[2][191] ) );
  INV_X2 U11969 ( .I(\MC_ARK_ARC_1_1/buf_output[191] ), .ZN(n6369) );
  NAND4_X2 U11971 ( .A1(\SB1_4_9/Component_Function_5/NAND4_in[1] ), .A2(n6788), .A3(n2897), .A4(\SB1_4_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_4_9/buf_output[5] ) );
  NAND3_X2 U11973 ( .A1(\SB1_2_17/i0_4 ), .A2(\SB1_2_17/i0_0 ), .A3(
        \SB1_2_17/i0_3 ), .ZN(n6795) );
  NAND3_X1 U11977 ( .A1(\SB2_0_16/i0[8] ), .A2(\SB2_0_16/i0_3 ), .A3(
        \SB2_0_16/i0[9] ), .ZN(n5071) );
  NAND4_X2 U11981 ( .A1(\SB2_2_16/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_2_16/Component_Function_3/NAND4_in[0] ), .A3(n6398), .A4(
        \SB2_2_16/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_16/buf_output[3] ) );
  XOR2_X1 U11983 ( .A1(\MC_ARK_ARC_1_3/temp2[155] ), .A2(n6534), .Z(n2109) );
  NAND4_X2 U11984 ( .A1(\SB2_1_10/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_10/Component_Function_0/NAND4_in[1] ), .A3(n775), .A4(
        \SB2_1_10/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_10/buf_output[0] ) );
  XOR2_X1 U11990 ( .A1(\MC_ARK_ARC_1_3/temp1[86] ), .A2(n3440), .Z(
        \MC_ARK_ARC_1_3/temp5[86] ) );
  NAND3_X1 U11992 ( .A1(\SB2_3_29/i0[8] ), .A2(\SB2_3_29/i1_7 ), .A3(
        \SB2_3_29/i0_4 ), .ZN(\SB2_3_29/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U12003 ( .A1(\RI5[1][156] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[0] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[90] ) );
  XOR2_X1 U12004 ( .A1(n3509), .A2(\MC_ARK_ARC_1_1/temp5[90] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[90] ) );
  XOR2_X1 U12005 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[77] ), .A2(\RI5[0][101] ), 
        .Z(n2670) );
  NAND4_X2 U12006 ( .A1(\SB2_4_26/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_4_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_4_26/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_4_26/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_4_26/buf_output[4] ) );
  XOR2_X1 U12013 ( .A1(\RI5[0][74] ), .A2(\RI5[0][104] ), .Z(n6657) );
  NAND3_X2 U12014 ( .A1(\SB1_3_7/i0[6] ), .A2(\SB1_3_7/i0[9] ), .A3(
        \SB1_3_7/i0_4 ), .ZN(n7250) );
  XOR2_X1 U12018 ( .A1(\RI5[3][75] ), .A2(\RI5[3][81] ), .Z(n6637) );
  XOR2_X1 U12024 ( .A1(\MC_ARK_ARC_1_4/temp3[130] ), .A2(
        \MC_ARK_ARC_1_4/temp4[130] ), .Z(n3051) );
  NAND4_X2 U12025 ( .A1(\SB1_1_10/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_10/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_1_10/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_1_10/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_1_10/buf_output[1] ) );
  NAND4_X2 U12026 ( .A1(\SB2_1_6/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_1_6/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_6/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_1_6/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_6/buf_output[1] ) );
  NAND4_X2 U12027 ( .A1(\SB3_10/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_10/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_2/NAND4_in[0] ), .A4(n6370), .ZN(
        \SB3_10/buf_output[2] ) );
  NAND3_X1 U12031 ( .A1(\SB3_10/i0_4 ), .A2(\SB3_10/i0_0 ), .A3(\SB3_10/i1_5 ), 
        .ZN(n6370) );
  NAND4_X2 U12037 ( .A1(\SB2_4_1/Component_Function_4/NAND4_in[1] ), .A2(n6384), .A3(\SB2_4_1/Component_Function_4/NAND4_in[0] ), .A4(n3717), .ZN(
        \SB2_4_1/buf_output[4] ) );
  NAND4_X2 U12038 ( .A1(n4079), .A2(
        \SB1_4_26/Component_Function_2/NAND4_in[0] ), .A3(n1261), .A4(n6371), 
        .ZN(\SB1_4_26/buf_output[2] ) );
  NAND3_X2 U12040 ( .A1(\SB1_4_26/i0[9] ), .A2(\SB1_4_26/i0_3 ), .A3(
        \SB1_4_26/i0[8] ), .ZN(n6371) );
  NAND4_X2 U12041 ( .A1(\SB2_2_16/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_16/Component_Function_4/NAND4_in[1] ), .A3(n1097), .A4(n6372), 
        .ZN(\SB2_2_16/buf_output[4] ) );
  NAND3_X2 U12047 ( .A1(\SB2_2_16/i0_4 ), .A2(\SB2_2_16/i1[9] ), .A3(
        \SB2_2_16/i1_5 ), .ZN(n6372) );
  NAND4_X2 U12049 ( .A1(\SB2_3_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_25/Component_Function_0/NAND4_in[1] ), .A3(n1796), .A4(n6373), 
        .ZN(\SB2_3_25/buf_output[0] ) );
  NAND4_X2 U12050 ( .A1(\SB2_3_6/Component_Function_5/NAND4_in[2] ), .A2(n5401), .A3(\SB2_3_6/Component_Function_5/NAND4_in[0] ), .A4(n6374), .ZN(
        \SB2_3_6/buf_output[5] ) );
  NAND3_X2 U12054 ( .A1(\SB2_3_6/i0[9] ), .A2(\SB2_3_6/i0[6] ), .A3(
        \SB2_3_6/i0_4 ), .ZN(n6374) );
  XOR2_X1 U12055 ( .A1(n6375), .A2(\MC_ARK_ARC_1_1/temp2[88] ), .Z(n1277) );
  XOR2_X1 U12057 ( .A1(\RI5[1][82] ), .A2(\RI5[1][88] ), .Z(n6375) );
  NAND2_X1 U12059 ( .A1(\SB1_3_10/i1[9] ), .A2(\SB1_3_10/i0_3 ), .ZN(
        \SB1_3_10/Component_Function_1/NAND4_in[0] ) );
  XOR2_X1 U12064 ( .A1(n6377), .A2(n6376), .Z(\MC_ARK_ARC_1_4/temp5[92] ) );
  XOR2_X1 U12067 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[86] ), .A2(\RI5[4][62] ), 
        .Z(n6376) );
  XOR2_X1 U12068 ( .A1(\RI5[4][38] ), .A2(\RI5[4][92] ), .Z(n6377) );
  XOR2_X1 U12070 ( .A1(n6378), .A2(n202), .Z(Ciphertext[50]) );
  NAND4_X2 U12072 ( .A1(\SB4_23/Component_Function_2/NAND4_in[0] ), .A2(n2129), 
        .A3(n2778), .A4(\SB4_23/Component_Function_2/NAND4_in[2] ), .ZN(n6378)
         );
  AOI22_X2 U12075 ( .A1(n6586), .A2(\SB1_1_27/i0[9] ), .B1(\SB1_1_27/i0_0 ), 
        .B2(\SB1_1_27/i3[0] ), .ZN(n6379) );
  XOR2_X1 U12078 ( .A1(\MC_ARK_ARC_1_1/temp2[78] ), .A2(n6380), .Z(
        \MC_ARK_ARC_1_1/temp5[78] ) );
  XOR2_X1 U12081 ( .A1(\RI5[1][78] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[72] ), 
        .Z(n6380) );
  NAND4_X2 U12082 ( .A1(n4543), .A2(\SB2_1_1/Component_Function_5/NAND4_in[0] ), .A3(n1963), .A4(n6381), .ZN(\SB2_1_1/buf_output[5] ) );
  NAND3_X2 U12085 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i0_0 ), .A3(
        \SB2_1_1/i0[6] ), .ZN(n6381) );
  XOR2_X1 U12089 ( .A1(n6382), .A2(\MC_ARK_ARC_1_0/temp1[25] ), .Z(
        \MC_ARK_ARC_1_0/temp5[25] ) );
  XOR2_X1 U12097 ( .A1(\RI5[0][163] ), .A2(\RI5[0][187] ), .Z(n6382) );
  NAND3_X2 U12101 ( .A1(\SB3_31/i0[6] ), .A2(\SB3_31/i0_3 ), .A3(
        \SB3_31/i0[10] ), .ZN(\SB3_31/Component_Function_2/NAND4_in[1] ) );
  NAND2_X2 U12103 ( .A1(n4579), .A2(n3802), .ZN(\RI3[0][141] ) );
  XOR2_X1 U12105 ( .A1(n6383), .A2(n16), .Z(Ciphertext[144]) );
  NAND4_X2 U12107 ( .A1(\SB4_7/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB4_7/Component_Function_0/NAND4_in[0] ), .ZN(n6383) );
  NAND3_X1 U12109 ( .A1(\SB2_4_1/i0[9] ), .A2(\SB2_4_1/i0_3 ), .A3(
        \SB2_4_1/i0[10] ), .ZN(n6384) );
  NAND4_X2 U12113 ( .A1(\SB1_4_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_4_1/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_4_1/Component_Function_5/NAND4_in[0] ), .A4(n6385), .ZN(
        \SB1_4_1/buf_output[5] ) );
  NAND3_X2 U12114 ( .A1(\SB1_4_1/i0[9] ), .A2(\SB1_4_1/i0_4 ), .A3(
        \SB1_4_1/i0[6] ), .ZN(n6385) );
  NAND4_X2 U12115 ( .A1(\SB2_3_21/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_21/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_21/Component_Function_0/NAND4_in[0] ), .A4(n6386), .ZN(
        \SB2_3_21/buf_output[0] ) );
  NAND3_X1 U12116 ( .A1(\SB1_4_1/i0[9] ), .A2(\SB1_4_1/i0[6] ), .A3(
        \SB1_4_1/i1_5 ), .ZN(\SB1_4_1/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U12117 ( .A1(\RI5[1][53] ), .A2(\RI5[1][107] ), .Z(n6388) );
  XOR2_X1 U12123 ( .A1(\RI5[1][77] ), .A2(\RI5[1][101] ), .Z(n6389) );
  AND3_X1 U12124 ( .A1(\SB1_1_15/buf_output[4] ), .A2(\SB1_1_19/buf_output[0] ), .A3(\SB1_1_18/buf_output[1] ), .Z(n6653) );
  XOR2_X1 U12125 ( .A1(\MC_ARK_ARC_1_2/temp4[87] ), .A2(n6390), .Z(n7472) );
  XOR2_X1 U12131 ( .A1(\RI5[2][153] ), .A2(\RI5[2][189] ), .Z(n6390) );
  XOR2_X1 U12133 ( .A1(\RI5[0][24] ), .A2(\RI5[0][48] ), .Z(
        \MC_ARK_ARC_1_0/temp2[78] ) );
  XOR2_X1 U12134 ( .A1(n6391), .A2(n206), .Z(Ciphertext[171]) );
  NAND4_X2 U12135 ( .A1(\SB4_3/Component_Function_3/NAND4_in[1] ), .A2(n4949), 
        .A3(\SB4_3/Component_Function_3/NAND4_in[3] ), .A4(n7258), .ZN(n6391)
         );
  XOR2_X1 U12138 ( .A1(n6392), .A2(n156), .Z(Ciphertext[168]) );
  NAND4_X2 U12139 ( .A1(\SB4_3/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB4_3/Component_Function_0/NAND4_in[0] ), .ZN(n6392) );
  NAND3_X2 U12140 ( .A1(\SB2_4_30/i0[10] ), .A2(\SB2_4_30/i1_5 ), .A3(
        \SB2_4_30/i1[9] ), .ZN(\SB2_4_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U12142 ( .A1(\SB1_4_3/i0_3 ), .A2(\SB1_4_3/i0[9] ), .A3(
        \SB1_4_3/i0[8] ), .ZN(n1571) );
  NAND4_X2 U12145 ( .A1(\SB2_2_17/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_2_17/Component_Function_2/NAND4_in[0] ), .A3(n4029), .A4(
        \SB2_2_17/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_17/buf_output[2] ) );
  XOR2_X1 U12150 ( .A1(n3428), .A2(\MC_ARK_ARC_1_3/temp3[180] ), .Z(n6535) );
  XOR2_X1 U12158 ( .A1(n6394), .A2(\MC_ARK_ARC_1_3/temp6[173] ), .Z(
        \RI1[4][173] ) );
  XOR2_X1 U12164 ( .A1(\MC_ARK_ARC_1_3/temp2[173] ), .A2(
        \MC_ARK_ARC_1_3/temp1[173] ), .Z(n6394) );
  NAND3_X1 U12169 ( .A1(\SB1_4_3/i0_3 ), .A2(\SB1_4_3/i0[10] ), .A3(
        \SB1_4_3/i0_4 ), .ZN(\SB1_4_3/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U12170 ( .A1(n6395), .A2(n1997), .Z(\MC_ARK_ARC_1_3/buf_output[67] )
         );
  XOR2_X1 U12173 ( .A1(\MC_ARK_ARC_1_3/temp1[67] ), .A2(
        \MC_ARK_ARC_1_3/temp4[67] ), .Z(n6395) );
  NAND4_X2 U12175 ( .A1(\SB2_4_20/Component_Function_4/NAND4_in[1] ), .A2(
        n1426), .A3(\SB2_4_20/Component_Function_4/NAND4_in[3] ), .A4(n6396), 
        .ZN(\SB2_4_20/buf_output[4] ) );
  NAND3_X2 U12176 ( .A1(\SB2_4_20/i0[9] ), .A2(\SB2_4_20/i0_3 ), .A3(
        \SB2_4_20/i0[10] ), .ZN(n6396) );
  XOR2_X1 U12182 ( .A1(n3051), .A2(n6397), .Z(\MC_ARK_ARC_1_4/buf_output[130] ) );
  NAND3_X2 U12185 ( .A1(\SB2_2_16/i0_4 ), .A2(\RI3[2][95] ), .A3(
        \SB2_2_16/i0_0 ), .ZN(n6398) );
  NAND4_X2 U12188 ( .A1(n2973), .A2(
        \SB2_3_17/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_17/Component_Function_5/NAND4_in[0] ), .A4(n6399), .ZN(
        \SB2_3_17/buf_output[5] ) );
  NAND3_X2 U12190 ( .A1(\SB2_3_17/i0_4 ), .A2(\SB2_3_17/i0[6] ), .A3(
        \SB2_3_17/i0[9] ), .ZN(n6399) );
  XOR2_X1 U12191 ( .A1(\SB2_3_5/buf_output[0] ), .A2(\RI5[3][162] ), .Z(n6722)
         );
  NAND4_X2 U12193 ( .A1(n7467), .A2(
        \SB1_2_17/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_17/Component_Function_0/NAND4_in[0] ), .A4(n6400), .ZN(
        \SB1_2_17/buf_output[0] ) );
  NAND4_X2 U12194 ( .A1(\SB2_0_25/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_25/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_25/Component_Function_4/NAND4_in[0] ), .A4(n6401), .ZN(
        \SB2_0_25/buf_output[4] ) );
  NAND3_X1 U12201 ( .A1(\SB2_0_25/i0_0 ), .A2(\SB2_0_25/i3[0] ), .A3(
        \SB2_0_25/i1_7 ), .ZN(n6401) );
  XOR2_X1 U12203 ( .A1(\MC_ARK_ARC_1_1/temp2[38] ), .A2(n6402), .Z(n6458) );
  XOR2_X1 U12204 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[32] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[38] ), .Z(n6402) );
  XOR2_X1 U12206 ( .A1(n6403), .A2(n139), .Z(Ciphertext[102]) );
  NAND4_X2 U12207 ( .A1(n4997), .A2(\SB4_14/Component_Function_0/NAND4_in[2] ), 
        .A3(\SB4_14/Component_Function_0/NAND4_in[3] ), .A4(
        \SB4_14/Component_Function_0/NAND4_in[0] ), .ZN(n6403) );
  NAND4_X2 U12209 ( .A1(\SB2_4_24/Component_Function_2/NAND4_in[1] ), .A2(
        n4167), .A3(\SB2_4_24/Component_Function_2/NAND4_in[3] ), .A4(n6404), 
        .ZN(\SB2_4_24/buf_output[2] ) );
  NAND3_X2 U12210 ( .A1(\SB2_4_24/i0[10] ), .A2(n5443), .A3(n6268), .ZN(n6404)
         );
  NAND3_X2 U12211 ( .A1(n6976), .A2(\SB2_0_16/i0_3 ), .A3(\SB2_0_16/i0[6] ), 
        .ZN(n6405) );
  XOR2_X1 U12212 ( .A1(n6407), .A2(n6406), .Z(n3224) );
  XOR2_X1 U12223 ( .A1(\RI5[4][14] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[86] ), 
        .Z(n6406) );
  XOR2_X1 U12225 ( .A1(n4446), .A2(n6408), .Z(\MC_ARK_ARC_1_0/temp5[2] ) );
  XOR2_X1 U12226 ( .A1(\RI5[0][140] ), .A2(\RI5[0][164] ), .Z(n6408) );
  INV_X1 U12228 ( .I(\SB1_0_8/buf_output[0] ), .ZN(\SB2_0_3/i3[0] ) );
  NAND4_X2 U12231 ( .A1(\SB1_0_8/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_8/Component_Function_0/NAND4_in[0] ), .A3(n7287), .A4(
        \SB1_0_8/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_0_8/buf_output[0] ) );
  XOR2_X1 U12233 ( .A1(n6409), .A2(n26), .Z(Ciphertext[173]) );
  XOR2_X1 U12234 ( .A1(\MC_ARK_ARC_1_2/temp5[90] ), .A2(
        \MC_ARK_ARC_1_2/temp6[90] ), .Z(n1500) );
  XOR2_X1 U12235 ( .A1(n7356), .A2(\MC_ARK_ARC_1_2/temp2[90] ), .Z(
        \MC_ARK_ARC_1_2/temp5[90] ) );
  XOR2_X1 U12236 ( .A1(n6410), .A2(n42), .Z(Ciphertext[170]) );
  NAND4_X2 U12237 ( .A1(n1828), .A2(n4953), .A3(
        \SB4_3/Component_Function_2/NAND4_in[2] ), .A4(n2728), .ZN(n6410) );
  NAND3_X1 U12238 ( .A1(\SB3_27/i0_3 ), .A2(\SB3_27/i0[6] ), .A3(
        \SB3_27/i1[9] ), .ZN(\SB3_27/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U12239 ( .A1(\SB1_3_2/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_2/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_2/Component_Function_2/NAND4_in[2] ), .A4(n6411), .ZN(
        \SB1_3_2/buf_output[2] ) );
  NAND3_X2 U12240 ( .A1(\SB1_3_2/i0_0 ), .A2(\SB1_3_2/i1_5 ), .A3(
        \SB1_3_2/i0_4 ), .ZN(n6411) );
  NAND3_X2 U12241 ( .A1(\SB1_3_25/i0_0 ), .A2(\SB1_3_25/i0[10] ), .A3(
        \SB1_3_25/i0[6] ), .ZN(n6412) );
  NAND4_X2 U12245 ( .A1(\SB1_2_10/Component_Function_2/NAND4_in[1] ), .A2(n958), .A3(n2296), .A4(n6414), .ZN(\SB1_2_10/buf_output[2] ) );
  NAND3_X2 U12247 ( .A1(\SB1_2_10/i0[10] ), .A2(\SB1_2_10/i1[9] ), .A3(
        \SB1_2_10/i1_5 ), .ZN(n6414) );
  XOR2_X1 U12250 ( .A1(n6416), .A2(n6415), .Z(\MC_ARK_ARC_1_1/temp6[102] ) );
  XOR2_X1 U12253 ( .A1(\RI5[1][12] ), .A2(n533), .Z(n6415) );
  XOR2_X1 U12254 ( .A1(\RI5[1][138] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[168] ), .Z(n6416) );
  NAND3_X2 U12257 ( .A1(\SB3_31/i0_0 ), .A2(\SB3_31/i1_5 ), .A3(\SB3_31/i0_4 ), 
        .ZN(n6417) );
  NAND4_X2 U12258 ( .A1(\SB2_3_9/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_9/Component_Function_5/NAND4_in[3] ), .A3(n6730), .A4(
        \SB2_3_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_9/buf_output[5] ) );
  XOR2_X1 U12260 ( .A1(n5320), .A2(n6418), .Z(\MC_ARK_ARC_1_3/temp5[153] ) );
  XOR2_X1 U12261 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[147] ), .A2(\RI5[3][153] ), .Z(n6418) );
  XOR2_X1 U12262 ( .A1(\RI5[4][122] ), .A2(\RI5[4][98] ), .Z(n6419) );
  XOR2_X1 U12269 ( .A1(\MC_ARK_ARC_1_2/temp2[109] ), .A2(
        \MC_ARK_ARC_1_2/temp1[109] ), .Z(n6420) );
  NAND3_X2 U12270 ( .A1(\SB1_2_14/i0_4 ), .A2(\SB1_2_14/i0[9] ), .A3(
        \SB1_2_14/i0[6] ), .ZN(n6421) );
  NAND4_X2 U12273 ( .A1(\SB2_1_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_8/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_8/Component_Function_3/NAND4_in[2] ), .A4(n6422), .ZN(
        \SB2_1_8/buf_output[3] ) );
  NAND3_X2 U12275 ( .A1(\SB2_1_8/i3[0] ), .A2(\SB2_1_8/i0[8] ), .A3(
        \SB2_1_8/i1_5 ), .ZN(n6422) );
  NAND3_X2 U12276 ( .A1(\SB1_4_6/i1_5 ), .A2(\SB1_4_6/i0[10] ), .A3(
        \SB1_4_6/i1[9] ), .ZN(n6423) );
  XOR2_X1 U12279 ( .A1(\MC_ARK_ARC_1_4/temp5[69] ), .A2(n6424), .Z(
        \MC_ARK_ARC_1_4/buf_output[69] ) );
  XOR2_X1 U12281 ( .A1(\MC_ARK_ARC_1_4/temp4[69] ), .A2(
        \MC_ARK_ARC_1_4/temp3[69] ), .Z(n6424) );
  XOR2_X1 U12283 ( .A1(n6425), .A2(\MC_ARK_ARC_1_2/temp1[134] ), .Z(
        \MC_ARK_ARC_1_2/temp5[134] ) );
  XOR2_X1 U12287 ( .A1(\RI5[2][104] ), .A2(\RI5[2][80] ), .Z(n6425) );
  NAND4_X2 U12288 ( .A1(\SB2_2_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_1/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_1/Component_Function_5/NAND4_in[0] ), .A4(n6426), .ZN(
        \SB2_2_1/buf_output[5] ) );
  NAND3_X2 U12294 ( .A1(\SB2_2_1/i0[6] ), .A2(\SB1_2_2/buf_output[4] ), .A3(
        \SB2_2_1/i0[9] ), .ZN(n6426) );
  NAND4_X2 U12295 ( .A1(\SB2_2_10/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_2_10/Component_Function_3/NAND4_in[1] ), .A3(n821), .A4(n6427), 
        .ZN(\SB2_2_10/buf_output[3] ) );
  NAND3_X2 U12296 ( .A1(\SB2_2_10/i0[6] ), .A2(\SB2_2_10/i0_3 ), .A3(
        \SB2_2_10/i1[9] ), .ZN(n6427) );
  XOR2_X1 U12301 ( .A1(n1579), .A2(n6428), .Z(\MC_ARK_ARC_1_0/buf_output[10] )
         );
  XOR2_X1 U12304 ( .A1(\MC_ARK_ARC_1_0/temp2[10] ), .A2(
        \MC_ARK_ARC_1_0/temp4[10] ), .Z(n6428) );
  XOR2_X1 U12305 ( .A1(\RI5[2][127] ), .A2(\RI5[2][163] ), .Z(
        \MC_ARK_ARC_1_2/temp3[61] ) );
  XOR2_X1 U12306 ( .A1(\MC_ARK_ARC_1_3/temp1[144] ), .A2(
        \MC_ARK_ARC_1_3/temp2[144] ), .Z(\MC_ARK_ARC_1_3/temp5[144] ) );
  NAND4_X2 U12311 ( .A1(\SB1_2_10/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_2_10/Component_Function_4/NAND4_in[0] ), .A3(n2004), .A4(
        \SB1_2_10/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_2_10/buf_output[4] ) );
  NAND3_X2 U12312 ( .A1(\SB1_1_29/i0[10] ), .A2(\SB1_1_29/i1[9] ), .A3(
        \SB1_1_29/i1_7 ), .ZN(n6429) );
  NAND3_X2 U12314 ( .A1(\SB3_27/i0_3 ), .A2(\SB3_27/i0[8] ), .A3(
        \SB3_27/i0[9] ), .ZN(n7512) );
  XOR2_X1 U12318 ( .A1(n6430), .A2(\MC_ARK_ARC_1_4/temp4[188] ), .Z(
        \MC_ARK_ARC_1_4/temp6[188] ) );
  XOR2_X1 U12320 ( .A1(\RI5[4][98] ), .A2(\RI5[4][62] ), .Z(n6430) );
  NAND3_X1 U12321 ( .A1(\SB4_24/i1[9] ), .A2(\SB4_24/i1_5 ), .A3(
        \SB3_26/buf_output[3] ), .ZN(n6431) );
  NAND3_X2 U12322 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0[6] ), .A3(
        \SB2_0_16/i1[9] ), .ZN(\SB2_0_16/Component_Function_3/NAND4_in[0] ) );
  BUF_X2 U12324 ( .I(\SB2_1_16/i1[9] ), .Z(n6432) );
  NAND3_X1 U12325 ( .A1(\SB4_25/i0[10] ), .A2(\SB4_25/i1_7 ), .A3(
        \SB4_25/i1[9] ), .ZN(n2840) );
  NAND3_X1 U12327 ( .A1(\SB1_1_11/i0[10] ), .A2(\SB1_1_11/i0[6] ), .A3(
        \SB1_1_11/i0_3 ), .ZN(\SB1_1_11/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U12328 ( .A1(\SB2_3_19/Component_Function_5/NAND4_in[2] ), .A2(
        n3193), .A3(\SB2_3_19/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_19/buf_output[5] ) );
  NAND4_X2 U12329 ( .A1(n2164), .A2(n6473), .A3(n7076), .A4(
        \SB2_3_30/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_30/buf_output[5] ) );
  NAND4_X2 U12331 ( .A1(\SB1_4_24/Component_Function_5/NAND4_in[1] ), .A2(
        n6871), .A3(n4108), .A4(\SB1_4_24/Component_Function_5/NAND4_in[0] ), 
        .ZN(\SB1_4_24/buf_output[5] ) );
  NAND4_X2 U12333 ( .A1(\SB2_2_13/Component_Function_2/NAND4_in[0] ), .A2(
        n6471), .A3(\SB2_2_13/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_2_13/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_13/buf_output[2] ) );
  NAND3_X1 U12341 ( .A1(\SB3_28/i1[9] ), .A2(\SB3_28/i0[10] ), .A3(
        \SB3_28/i1_5 ), .ZN(\SB3_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U12343 ( .A1(\SB1_3_7/i0_3 ), .A2(\SB1_3_7/i0[9] ), .A3(
        \SB1_3_7/i0[8] ), .ZN(\SB1_3_7/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U12345 ( .A1(\SB2_2_9/i0[9] ), .A2(\SB2_2_9/i0_3 ), .A3(
        \SB2_2_9/i0[8] ), .ZN(n6433) );
  NAND3_X2 U12346 ( .A1(\SB1_3_27/i0[9] ), .A2(\SB1_3_27/i0_4 ), .A3(
        \SB1_3_27/i0[6] ), .ZN(n6434) );
  NAND3_X2 U12347 ( .A1(\SB3_19/i0[6] ), .A2(\SB3_19/i0_4 ), .A3(
        \SB3_19/i0[9] ), .ZN(n5411) );
  NAND3_X2 U12352 ( .A1(\SB2_0_26/i0[8] ), .A2(\SB2_0_26/i0[9] ), .A3(
        \SB2_0_26/i0_3 ), .ZN(\SB2_0_26/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U12355 ( .A1(n6435), .A2(n25), .Z(Ciphertext[66]) );
  NAND4_X2 U12356 ( .A1(n3909), .A2(n6959), .A3(n6917), .A4(
        \SB4_20/Component_Function_0/NAND4_in[0] ), .ZN(n6435) );
  INV_X2 U12362 ( .I(\SB1_1_3/buf_output[3] ), .ZN(\SB2_1_1/i0[8] ) );
  XOR2_X1 U12363 ( .A1(\RI5[1][35] ), .A2(\RI5[1][29] ), .Z(n6436) );
  NAND3_X2 U12365 ( .A1(\SB3_11/i0[10] ), .A2(\SB3_11/i0_3 ), .A3(
        \SB3_11/i0[6] ), .ZN(\SB3_11/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U12366 ( .A1(\SB2_3_23/buf_output[0] ), .A2(\RI5[3][84] ), .Z(
        \MC_ARK_ARC_1_3/temp1[84] ) );
  XOR2_X1 U12371 ( .A1(\SB2_1_6/buf_output[2] ), .A2(\RI5[1][2] ), .Z(
        \MC_ARK_ARC_1_1/temp2[32] ) );
  XOR2_X1 U12372 ( .A1(\MC_ARK_ARC_1_0/temp4[71] ), .A2(n1550), .Z(n6831) );
  XOR2_X1 U12375 ( .A1(\MC_ARK_ARC_1_1/temp1[157] ), .A2(n6438), .Z(n4165) );
  XOR2_X1 U12377 ( .A1(\RI5[1][127] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[103] ), .Z(n6438) );
  XOR2_X1 U12378 ( .A1(\RI5[0][87] ), .A2(\RI5[0][63] ), .Z(
        \MC_ARK_ARC_1_0/temp2[117] ) );
  XOR2_X1 U12382 ( .A1(\MC_ARK_ARC_1_0/temp4[173] ), .A2(n6441), .Z(n7421) );
  XOR2_X1 U12383 ( .A1(\RI5[0][167] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[173] ), .Z(n6441) );
  NAND4_X2 U12384 ( .A1(n4631), .A2(
        \SB2_1_22/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_1_22/Component_Function_3/NAND4_in[0] ), .A4(n6442), .ZN(
        \SB2_1_22/buf_output[3] ) );
  NAND3_X2 U12385 ( .A1(\SB2_1_22/i0_0 ), .A2(\SB2_1_22/i0_3 ), .A3(
        \SB2_1_22/i0_4 ), .ZN(n6442) );
  NAND4_X2 U12390 ( .A1(\SB1_1_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_12/Component_Function_1/NAND4_in[2] ), .A4(n6443), .ZN(
        \SB1_1_12/buf_output[1] ) );
  NAND3_X2 U12391 ( .A1(\SB1_1_12/i0[8] ), .A2(\SB1_1_12/i0_4 ), .A3(
        \SB1_1_12/i1_7 ), .ZN(n6443) );
  XOR2_X1 U12392 ( .A1(n6445), .A2(\MC_ARK_ARC_1_3/temp1[102] ), .Z(n603) );
  NAND4_X2 U12396 ( .A1(\SB2_0_4/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_4/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_4/Component_Function_5/NAND4_in[0] ), .A4(n6444), .ZN(
        \SB2_0_4/buf_output[5] ) );
  NAND3_X2 U12401 ( .A1(\SB2_0_4/i0[6] ), .A2(\RI3[0][166] ), .A3(
        \SB2_0_4/i0[9] ), .ZN(n6444) );
  NAND2_X1 U12402 ( .A1(\SB1_2_1/Component_Function_4/NAND4_in[3] ), .A2(n7193), .ZN(n4838) );
  XOR2_X1 U12403 ( .A1(\RI5[3][168] ), .A2(\RI5[3][12] ), .Z(n6445) );
  XOR2_X1 U12414 ( .A1(\RI5[2][57] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[63] ), 
        .Z(n6446) );
  OR3_X1 U12417 ( .A1(\RI3[0][33] ), .A2(\SB2_0_26/i0[6] ), .A3(n3510), .Z(
        n4535) );
  XOR2_X1 U12421 ( .A1(n6448), .A2(n49), .Z(Ciphertext[85]) );
  NAND4_X2 U12422 ( .A1(\SB4_17/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_17/Component_Function_1/NAND4_in[0] ), .ZN(n6448) );
  XOR2_X1 U12427 ( .A1(n5288), .A2(\MC_ARK_ARC_1_1/temp4[122] ), .Z(n4745) );
  XOR2_X1 U12428 ( .A1(n2852), .A2(\MC_ARK_ARC_1_2/temp6[168] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[168] ) );
  XOR2_X1 U12429 ( .A1(n7135), .A2(n6449), .Z(\MC_ARK_ARC_1_2/buf_output[59] )
         );
  XOR2_X1 U12431 ( .A1(\MC_ARK_ARC_1_2/temp1[59] ), .A2(n845), .Z(n6449) );
  INV_X2 U12435 ( .I(\RI3[0][177] ), .ZN(\SB2_0_2/i0[8] ) );
  NAND4_X2 U12436 ( .A1(\SB1_0_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_4/Component_Function_3/NAND4_in[1] ), .A3(n2622), .A4(
        \SB1_0_4/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][177] ) );
  INV_X1 U12437 ( .I(\SB1_2_14/buf_output[0] ), .ZN(\SB2_2_9/i3[0] ) );
  NAND4_X2 U12438 ( .A1(\SB1_2_14/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_14/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_14/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_14/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_14/buf_output[0] ) );
  XOR2_X1 U12444 ( .A1(\MC_ARK_ARC_1_2/temp5[101] ), .A2(n6450), .Z(
        \RI1[3][101] ) );
  NAND4_X2 U12445 ( .A1(n3631), .A2(
        \SB1_1_22/Component_Function_2/NAND4_in[2] ), .A3(n7578), .A4(
        \SB1_1_22/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_1_22/buf_output[2] ) );
  NAND4_X2 U12446 ( .A1(\SB1_1_17/Component_Function_4/NAND4_in[1] ), .A2(
        n4394), .A3(\SB1_1_17/Component_Function_4/NAND4_in[0] ), .A4(n7481), 
        .ZN(\SB1_1_17/buf_output[4] ) );
  XOR2_X1 U12448 ( .A1(n7570), .A2(n7571), .Z(\MC_ARK_ARC_1_0/buf_output[86] )
         );
  INV_X2 U12450 ( .I(\SB1_2_22/buf_output[2] ), .ZN(\SB2_2_19/i1[9] ) );
  NAND4_X2 U12452 ( .A1(\SB1_2_22/Component_Function_2/NAND4_in[1] ), .A2(
        n7464), .A3(n6599), .A4(n4582), .ZN(\SB1_2_22/buf_output[2] ) );
  XOR2_X1 U12454 ( .A1(\RI5[3][111] ), .A2(\RI5[3][87] ), .Z(
        \MC_ARK_ARC_1_3/temp2[141] ) );
  XOR2_X1 U12461 ( .A1(n2082), .A2(n2083), .Z(\MC_ARK_ARC_1_2/buf_output[123] ) );
  CLKBUF_X8 U12463 ( .I(\SB2_3_13/i0_4 ), .Z(n6746) );
  AND2_X1 U12465 ( .A1(n6563), .A2(n5160), .Z(n5255) );
  XOR2_X1 U12470 ( .A1(\RI5[3][174] ), .A2(\RI5[3][138] ), .Z(
        \MC_ARK_ARC_1_3/temp3[72] ) );
  XOR2_X1 U12476 ( .A1(n3855), .A2(n2371), .Z(\MC_ARK_ARC_1_2/buf_output[93] )
         );
  NAND4_X2 U12478 ( .A1(n5092), .A2(
        \SB1_3_12/Component_Function_4/NAND4_in[3] ), .A3(n4599), .A4(
        \SB1_3_12/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_3_12/buf_output[4] ) );
  XOR2_X1 U12484 ( .A1(n2394), .A2(n4865), .Z(\RI1[4][141] ) );
  XOR2_X1 U12485 ( .A1(\RI5[0][69] ), .A2(\RI5[0][105] ), .Z(
        \MC_ARK_ARC_1_0/temp3[3] ) );
  XOR2_X1 U12493 ( .A1(\RI5[4][44] ), .A2(\RI5[4][68] ), .Z(
        \MC_ARK_ARC_1_4/temp2[98] ) );
  NAND3_X2 U12494 ( .A1(\SB2_0_25/i0_0 ), .A2(\SB2_0_25/i1_5 ), .A3(
        \SB2_0_25/i0_4 ), .ZN(\SB2_0_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U12495 ( .A1(\SB1_4_16/i1_5 ), .A2(\SB1_4_16/i0[8] ), .A3(
        \SB1_4_16/i3[0] ), .ZN(n4834) );
  XOR2_X1 U12501 ( .A1(n6874), .A2(n6964), .Z(\MC_ARK_ARC_1_4/buf_output[186] ) );
  NAND2_X1 U12502 ( .A1(\SB1_4_14/i0_0 ), .A2(\SB1_4_14/i3[0] ), .ZN(n6555) );
  NAND3_X1 U12506 ( .A1(\SB4_29/i0_0 ), .A2(\SB4_29/i0_3 ), .A3(\SB4_29/i0[7] ), .ZN(n5349) );
  XOR2_X1 U12517 ( .A1(n6451), .A2(n86), .Z(Ciphertext[107]) );
  NAND4_X2 U12519 ( .A1(\SB4_14/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_14/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_14/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_14/Component_Function_5/NAND4_in[0] ), .ZN(n6451) );
  NAND3_X2 U12520 ( .A1(\SB1_0_20/i0[6] ), .A2(\SB1_0_20/i0[10] ), .A3(
        \SB1_0_20/i0_0 ), .ZN(\SB1_0_20/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U12521 ( .A1(n6453), .A2(n6452), .Z(\MC_ARK_ARC_1_1/buf_output[173] ) );
  XOR2_X1 U12530 ( .A1(n7005), .A2(\MC_ARK_ARC_1_1/temp4[173] ), .Z(n6452) );
  NAND4_X2 U12531 ( .A1(\SB1_0_4/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_4/Component_Function_2/NAND4_in[2] ), .A3(n3690), .A4(n6454), 
        .ZN(\RI3[0][182] ) );
  NAND3_X2 U12532 ( .A1(\SB1_0_4/i0[10] ), .A2(\SB1_0_4/i1[9] ), .A3(
        \SB1_0_4/i1_5 ), .ZN(n6454) );
  XOR2_X1 U12533 ( .A1(\RI5[1][173] ), .A2(n17), .Z(n6455) );
  XOR2_X1 U12536 ( .A1(\RI5[1][143] ), .A2(\RI5[1][17] ), .Z(n6456) );
  XOR2_X1 U12539 ( .A1(\MC_ARK_ARC_1_3/temp2[104] ), .A2(n6457), .Z(
        \MC_ARK_ARC_1_3/temp5[104] ) );
  XOR2_X1 U12540 ( .A1(\RI5[3][98] ), .A2(\RI5[3][104] ), .Z(n6457) );
  XOR2_X1 U12542 ( .A1(n6458), .A2(n2885), .Z(\MC_ARK_ARC_1_1/buf_output[38] )
         );
  XOR2_X1 U12544 ( .A1(n6460), .A2(n6459), .Z(n2049) );
  XOR2_X1 U12545 ( .A1(\SB2_0_22/buf_output[2] ), .A2(n78), .Z(n6459) );
  XOR2_X1 U12547 ( .A1(\SB2_0_28/buf_output[2] ), .A2(\RI5[0][8] ), .Z(n6460)
         );
  XOR2_X1 U12548 ( .A1(n3408), .A2(n6461), .Z(n4346) );
  XOR2_X1 U12549 ( .A1(\RI5[1][161] ), .A2(\RI5[1][185] ), .Z(n6461) );
  XOR2_X1 U12550 ( .A1(n6462), .A2(\MC_ARK_ARC_1_2/temp5[161] ), .Z(
        \RI1[3][161] ) );
  XOR2_X1 U12551 ( .A1(\MC_ARK_ARC_1_2/temp3[161] ), .A2(
        \MC_ARK_ARC_1_2/temp4[161] ), .Z(n6462) );
  INV_X2 U12556 ( .I(\SB1_1_8/buf_output[3] ), .ZN(\SB2_1_6/i0[8] ) );
  NAND4_X2 U12557 ( .A1(\SB1_1_8/Component_Function_3/NAND4_in[1] ), .A2(n5133), .A3(\SB1_1_8/Component_Function_3/NAND4_in[0] ), .A4(n6664), .ZN(
        \SB1_1_8/buf_output[3] ) );
  XOR2_X1 U12560 ( .A1(\RI5[2][104] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[98] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[104] ) );
  XOR2_X1 U12561 ( .A1(\MC_ARK_ARC_1_1/temp1[87] ), .A2(n6463), .Z(
        \MC_ARK_ARC_1_1/temp5[87] ) );
  XOR2_X1 U12562 ( .A1(\RI5[1][57] ), .A2(\RI5[1][33] ), .Z(n6463) );
  XOR2_X1 U12565 ( .A1(n6464), .A2(\MC_ARK_ARC_1_3/temp6[28] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[28] ) );
  XOR2_X1 U12567 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[147] ), .A2(\RI5[2][153] ), .Z(\MC_ARK_ARC_1_2/temp1[153] ) );
  XOR2_X1 U12568 ( .A1(n1645), .A2(n6465), .Z(n5321) );
  XOR2_X1 U12578 ( .A1(\RI5[1][170] ), .A2(\RI5[1][176] ), .Z(n6465) );
  INV_X2 U12581 ( .I(\SB1_3_12/buf_output[2] ), .ZN(\SB2_3_9/i1[9] ) );
  NAND4_X2 U12582 ( .A1(n3246), .A2(
        \SB1_3_12/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_12/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_3_12/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_3_12/buf_output[2] ) );
  XOR2_X1 U12584 ( .A1(n6466), .A2(\MC_ARK_ARC_1_3/temp6[24] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[24] ) );
  XOR2_X1 U12588 ( .A1(\MC_ARK_ARC_1_3/temp1[24] ), .A2(n6722), .Z(n6466) );
  NAND3_X2 U12592 ( .A1(\SB2_0_23/i0[6] ), .A2(\SB2_0_23/i1_5 ), .A3(
        \SB2_0_23/i0[9] ), .ZN(\SB2_0_23/Component_Function_1/NAND4_in[2] ) );
  INV_X2 U12601 ( .I(\SB1_3_31/buf_output[3] ), .ZN(\SB2_3_29/i0[8] ) );
  NAND3_X1 U12602 ( .A1(\SB3_11/i0[8] ), .A2(\SB3_11/i0_4 ), .A3(\SB3_11/i1_7 ), .ZN(\SB3_11/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U12605 ( .I(\SB1_1_22/buf_output[5] ), .ZN(\SB2_1_22/i1_5 ) );
  NAND4_X2 U12606 ( .A1(\SB1_1_22/Component_Function_5/NAND4_in[2] ), .A2(
        n2531), .A3(n6507), .A4(\SB1_1_22/Component_Function_5/NAND4_in[0] ), 
        .ZN(\SB1_1_22/buf_output[5] ) );
  NAND4_X2 U12614 ( .A1(\SB1_2_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_1/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_1/Component_Function_1/NAND4_in[0] ), .A4(n6467), .ZN(
        \SB1_2_1/buf_output[1] ) );
  NAND3_X2 U12616 ( .A1(n7139), .A2(n3065), .A3(n6468), .ZN(
        \SB1_1_21/buf_output[5] ) );
  AOI22_X2 U12619 ( .A1(n2355), .A2(\SB1_1_21/i0[9] ), .B1(\SB1_1_21/i3[0] ), 
        .B2(\SB1_1_21/i0_0 ), .ZN(n6468) );
  NAND4_X2 U12620 ( .A1(n5006), .A2(
        \SB1_4_17/Component_Function_5/NAND4_in[1] ), .A3(n3796), .A4(n6469), 
        .ZN(\SB1_4_17/buf_output[5] ) );
  INV_X2 U12627 ( .I(\RI3[0][182] ), .ZN(\SB2_0_1/i1[9] ) );
  NAND4_X2 U12628 ( .A1(\SB2_0_26/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_26/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_0_26/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_0_26/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_0_26/buf_output[0] ) );
  NAND4_X2 U12629 ( .A1(\SB2_3_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_9/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_3_9/Component_Function_2/NAND4_in[1] ), .A4(n6470), .ZN(
        \SB2_3_9/buf_output[2] ) );
  NAND3_X2 U12630 ( .A1(\SB2_3_9/i0_0 ), .A2(\SB2_3_9/i1_5 ), .A3(
        \SB1_3_10/buf_output[4] ), .ZN(n6470) );
  NAND4_X2 U12638 ( .A1(\SB1_0_28/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_28/Component_Function_3/NAND4_in[0] ), .A3(n2540), .A4(
        \SB1_0_28/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_0_28/buf_output[3] ) );
  NAND3_X1 U12639 ( .A1(\SB1_0_29/i0_0 ), .A2(\SB1_0_29/i3[0] ), .A3(
        \SB1_0_29/i1_7 ), .ZN(\SB1_0_29/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U12642 ( .A1(\SB2_0_4/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_4/Component_Function_2/NAND4_in[0] ), .A3(n5248), .A4(n6472), 
        .ZN(\SB2_0_4/buf_output[2] ) );
  NAND3_X2 U12643 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0[10] ), .A3(
        \SB2_0_4/i0[6] ), .ZN(n6472) );
  NAND3_X2 U12644 ( .A1(\SB2_3_30/i0_0 ), .A2(\SB2_3_30/i0[6] ), .A3(
        \SB2_3_30/i0[10] ), .ZN(n6473) );
  XOR2_X1 U12645 ( .A1(\RI5[0][81] ), .A2(\RI5[0][45] ), .Z(
        \MC_ARK_ARC_1_0/temp3[171] ) );
  NAND4_X2 U12655 ( .A1(\SB2_0_26/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_26/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_26/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_26/buf_output[3] ) );
  XOR2_X1 U12656 ( .A1(n1423), .A2(\MC_ARK_ARC_1_0/temp5[179] ), .Z(
        \RI1[1][179] ) );
  XOR2_X1 U12657 ( .A1(n1733), .A2(\MC_ARK_ARC_1_0/temp2[61] ), .Z(
        \MC_ARK_ARC_1_0/temp5[61] ) );
  NAND3_X2 U12660 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i0_0 ), .A3(\SB4_28/i0_4 ), 
        .ZN(n7497) );
  NAND3_X1 U12665 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i0_3 ), .A3(
        \SB4_28/i0[6] ), .ZN(n2015) );
  NAND4_X2 U12666 ( .A1(\SB1_2_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_2_3/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_3/buf_output[3] ) );
  NAND4_X2 U12667 ( .A1(\SB3_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_6/Component_Function_2/NAND4_in[1] ), .A3(n7026), .A4(
        \SB3_6/Component_Function_2/NAND4_in[2] ), .ZN(\SB3_6/buf_output[2] )
         );
  XOR2_X1 U12669 ( .A1(n3736), .A2(n3224), .Z(\MC_ARK_ARC_1_4/buf_output[20] )
         );
  NAND4_X2 U12670 ( .A1(n5233), .A2(
        \SB2_1_21/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_21/Component_Function_2/NAND4_in[2] ), .A4(n2931), .ZN(
        \SB2_1_21/buf_output[2] ) );
  INV_X2 U12672 ( .I(\SB1_1_24/buf_output[2] ), .ZN(\SB2_1_21/i1[9] ) );
  NAND4_X2 U12679 ( .A1(n2380), .A2(
        \SB1_1_24/Component_Function_2/NAND4_in[1] ), .A3(n6696), .A4(n6697), 
        .ZN(\SB1_1_24/buf_output[2] ) );
  NAND3_X1 U12680 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i0_3 ), .A3(
        \SB4_28/i0[9] ), .ZN(\SB4_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U12681 ( .A1(\SB1_2_22/i0[10] ), .A2(\SB1_2_22/i0[6] ), .A3(
        \SB1_2_22/i0_0 ), .ZN(\SB1_2_22/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U12682 ( .A1(\SB1_2_24/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_24/Component_Function_3/NAND4_in[0] ), .A3(n1019), .A4(n6475), 
        .ZN(\SB1_2_24/buf_output[3] ) );
  NAND4_X2 U12685 ( .A1(\SB2_1_25/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_25/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_25/Component_Function_0/NAND4_in[0] ), .A4(n6476), .ZN(
        \SB2_1_25/buf_output[0] ) );
  NAND3_X1 U12687 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB1_1_27/buf_output[3] ), .A3(
        \SB1_1_26/buf_output[4] ), .ZN(n6476) );
  NAND3_X2 U12688 ( .A1(\SB1_2_3/i0_4 ), .A2(\SB1_2_3/i0[9] ), .A3(
        \SB1_2_3/i0[6] ), .ZN(n2595) );
  NAND2_X2 U12689 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i1[9] ), .ZN(n6477) );
  NAND3_X1 U12692 ( .A1(\SB3_4/i3[0] ), .A2(\SB3_4/i1_5 ), .A3(\SB3_4/i0[8] ), 
        .ZN(\SB3_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U12693 ( .A1(\SB2_0_18/i0_3 ), .A2(\SB2_0_18/i0_0 ), .A3(
        \RI3[0][82] ), .ZN(\SB2_0_18/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U12696 ( .A1(n6478), .A2(\MC_ARK_ARC_1_2/temp5[73] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[73] ) );
  XOR2_X1 U12697 ( .A1(\MC_ARK_ARC_1_2/temp4[73] ), .A2(
        \MC_ARK_ARC_1_2/temp3[73] ), .Z(n6478) );
  NAND3_X2 U12698 ( .A1(\SB1_0_18/i0[10] ), .A2(\SB1_0_18/i0[6] ), .A3(n6290), 
        .ZN(\SB1_0_18/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U12699 ( .A1(\MC_ARK_ARC_1_0/temp3[1] ), .A2(
        \MC_ARK_ARC_1_0/temp4[1] ), .Z(n6615) );
  INV_X2 U12701 ( .I(\SB1_1_0/buf_output[3] ), .ZN(\SB2_1_30/i0[8] ) );
  NAND4_X2 U12703 ( .A1(\SB1_1_0/Component_Function_3/NAND4_in[1] ), .A2(n4391), .A3(\SB1_1_0/Component_Function_3/NAND4_in[0] ), .A4(n2496), .ZN(
        \SB1_1_0/buf_output[3] ) );
  NAND4_X2 U12705 ( .A1(\SB1_4_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_4_14/Component_Function_5/NAND4_in[3] ), .A3(n6555), .A4(n6479), 
        .ZN(\SB1_4_14/buf_output[5] ) );
  NAND3_X2 U12707 ( .A1(\SB1_4_14/i0[6] ), .A2(\SB1_4_14/i0[10] ), .A3(
        \SB1_4_14/i0_0 ), .ZN(n6479) );
  XOR2_X1 U12710 ( .A1(\MC_ARK_ARC_1_0/temp4[51] ), .A2(n6481), .Z(
        \MC_ARK_ARC_1_0/temp6[51] ) );
  XOR2_X1 U12711 ( .A1(\RI5[0][117] ), .A2(\RI5[0][153] ), .Z(n6481) );
  AND2_X1 U12712 ( .A1(n3939), .A2(n910), .Z(n2843) );
  NAND4_X2 U12713 ( .A1(\SB1_0_18/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_18/Component_Function_3/NAND4_in[0] ), .A3(n7485), .A4(
        \SB1_0_18/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_0_18/buf_output[3] ) );
  AND2_X1 U12714 ( .A1(\SB1_0_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_18/Component_Function_1/NAND4_in[3] ), .Z(n2842) );
  NAND3_X2 U12715 ( .A1(\SB2_1_9/i0[10] ), .A2(\SB2_1_9/i0_0 ), .A3(
        \SB2_1_9/i0[6] ), .ZN(\SB2_1_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U12716 ( .A1(\SB2_4_6/i0_3 ), .A2(\SB2_4_6/i0_4 ), .A3(
        \SB2_4_6/i1[9] ), .ZN(n2101) );
  NOR2_X2 U12717 ( .A1(n6825), .A2(n6824), .ZN(n4662) );
  NAND3_X2 U12718 ( .A1(\SB2_1_2/i0[10] ), .A2(\SB2_1_2/i1_5 ), .A3(
        \SB2_1_2/i1[9] ), .ZN(n6601) );
  NAND2_X2 U12719 ( .A1(n1920), .A2(\SB1_0_2/Component_Function_3/NAND4_in[1] ), .ZN(n3363) );
  XOR2_X1 U12720 ( .A1(\RI5[0][103] ), .A2(\RI5[0][127] ), .Z(
        \MC_ARK_ARC_1_0/temp2[157] ) );
  XOR2_X1 U12721 ( .A1(n1506), .A2(\MC_ARK_ARC_1_3/buf_datainput[32] ), .Z(
        \MC_ARK_ARC_1_3/temp3[122] ) );
  NAND3_X1 U12722 ( .A1(\SB1_2_17/i0[6] ), .A2(\SB1_2_17/i0_3 ), .A3(
        \SB1_2_17/i0[10] ), .ZN(\SB1_2_17/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U12723 ( .A1(n6482), .A2(\MC_ARK_ARC_1_1/temp4[85] ), .Z(
        \MC_ARK_ARC_1_1/temp6[85] ) );
  XOR2_X1 U12724 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[151] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[187] ), .Z(n6482) );
  XOR2_X1 U12725 ( .A1(n6483), .A2(n150), .Z(Ciphertext[95]) );
  NAND4_X2 U12726 ( .A1(\SB4_16/Component_Function_5/NAND4_in[2] ), .A2(n1020), 
        .A3(n5037), .A4(\SB4_16/Component_Function_5/NAND4_in[3] ), .ZN(n6483)
         );
  NAND3_X2 U12727 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i0_3 ), .A3(
        \SB4_16/i0[9] ), .ZN(n6484) );
  NAND3_X1 U12728 ( .A1(\SB1_3_28/i0[10] ), .A2(\SB1_3_28/i1[9] ), .A3(
        \SB1_3_28/i1_7 ), .ZN(\SB1_3_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U12729 ( .A1(\SB3_12/i0[9] ), .A2(\RI1[5][119] ), .A3(
        \SB3_12/i0[8] ), .ZN(n6486) );
  XOR2_X1 U12730 ( .A1(n6487), .A2(\MC_ARK_ARC_1_3/temp5[140] ), .Z(
        \RI1[4][140] ) );
  XOR2_X1 U12731 ( .A1(\MC_ARK_ARC_1_3/temp3[140] ), .A2(
        \MC_ARK_ARC_1_3/temp4[140] ), .Z(n6487) );
  NAND4_X2 U12732 ( .A1(\SB1_1_28/Component_Function_5/NAND4_in[1] ), .A2(
        n3107), .A3(n6894), .A4(\SB1_1_28/Component_Function_5/NAND4_in[0] ), 
        .ZN(\SB1_1_28/buf_output[5] ) );
  XOR2_X1 U12733 ( .A1(\RI5[3][75] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[129] ), 
        .Z(n6488) );
  NAND4_X2 U12734 ( .A1(\SB2_1_28/Component_Function_2/NAND4_in[0] ), .A2(n942), .A3(\SB2_1_28/Component_Function_2/NAND4_in[1] ), .A4(n3329), .ZN(
        \SB2_1_28/buf_output[2] ) );
  XOR2_X1 U12735 ( .A1(n6490), .A2(n6489), .Z(n4345) );
  XOR2_X1 U12736 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[182] ), .A2(n29), .Z(
        n6489) );
  NAND3_X1 U12737 ( .A1(\SB4_29/i0_0 ), .A2(\SB4_29/i0[10] ), .A3(
        \SB4_29/i0[6] ), .ZN(\SB4_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U12738 ( .A1(\SB1_1_23/i0[9] ), .A2(\SB1_1_23/i0[8] ), .A3(
        \SB1_1_23/i0_3 ), .ZN(n1634) );
  NAND4_X2 U12739 ( .A1(\SB3_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_0/Component_Function_2/NAND4_in[1] ), .A3(n2556), .A4(n2676), 
        .ZN(\SB3_0/buf_output[2] ) );
  NAND4_X2 U12740 ( .A1(\SB2_4_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_7/Component_Function_4/NAND4_in[3] ), .A3(n6627), .A4(
        \SB2_4_7/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_4_7/buf_output[4] ) );
  XOR2_X1 U12741 ( .A1(\RI5[1][106] ), .A2(\RI5[1][112] ), .Z(
        \MC_ARK_ARC_1_1/temp1[112] ) );
  NAND3_X1 U12742 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB2_3_7/i0_4 ), .A3(
        \SB2_3_7/i0[10] ), .ZN(\SB2_3_7/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U12743 ( .A1(\SB3_20/Component_Function_1/NAND4_in[1] ), .A2(n3916), 
        .A3(\SB3_20/Component_Function_1/NAND4_in[0] ), .A4(n6491), .ZN(
        \SB3_20/buf_output[1] ) );
  INV_X2 U12744 ( .I(\SB1_2_26/buf_output[2] ), .ZN(\SB2_2_23/i1[9] ) );
  NAND4_X2 U12745 ( .A1(\SB1_2_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_26/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_2_26/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_26/buf_output[2] ) );
  NAND3_X2 U12746 ( .A1(\SB1_4_19/i0_0 ), .A2(\SB1_4_19/i1_7 ), .A3(
        \SB1_4_19/i3[0] ), .ZN(n6492) );
  NAND4_X2 U12747 ( .A1(\SB1_4_21/Component_Function_2/NAND4_in[1] ), .A2(
        n4376), .A3(n6670), .A4(n6684), .ZN(\SB1_4_21/buf_output[2] ) );
  NOR2_X2 U12748 ( .A1(n2326), .A2(n6493), .ZN(\SB2_0_17/i0[7] ) );
  NAND3_X2 U12749 ( .A1(\SB1_2_11/i1_5 ), .A2(\SB1_2_11/i0_4 ), .A3(
        \SB1_2_11/i0_0 ), .ZN(n6494) );
  XOR2_X1 U12750 ( .A1(n6495), .A2(\MC_ARK_ARC_1_2/temp4[140] ), .Z(
        \MC_ARK_ARC_1_2/temp6[140] ) );
  XOR2_X1 U12751 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[14] ), .A2(\RI5[2][50] ), 
        .Z(n6495) );
  NAND2_X1 U12752 ( .A1(\SB1_0_26/Component_Function_4/NAND4_in[1] ), .A2(
        n6496), .ZN(n2064) );
  NAND3_X1 U12753 ( .A1(\SB1_0_26/i0_0 ), .A2(\SB1_0_26/i0[9] ), .A3(
        \SB1_0_26/i0[8] ), .ZN(n6496) );
  NAND4_X2 U12754 ( .A1(\SB2_3_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_28/Component_Function_1/NAND4_in[0] ), .A3(n1182), .A4(n6497), 
        .ZN(\SB2_3_28/buf_output[1] ) );
  NAND3_X2 U12755 ( .A1(\SB2_3_28/i0[9] ), .A2(\SB2_3_28/i1_5 ), .A3(
        \SB2_3_28/i0[6] ), .ZN(n6497) );
  XOR2_X1 U12756 ( .A1(n6499), .A2(n6498), .Z(n7377) );
  XOR2_X1 U12757 ( .A1(\RI5[0][44] ), .A2(\RI5[0][152] ), .Z(n6498) );
  INV_X2 U12758 ( .I(\SB1_2_7/buf_output[2] ), .ZN(\SB2_2_4/i1[9] ) );
  NAND4_X2 U12759 ( .A1(\SB1_2_7/Component_Function_2/NAND4_in[0] ), .A2(n5101), .A3(\SB1_2_7/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_2_7/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_7/buf_output[2] ) );
  NAND3_X2 U12760 ( .A1(\SB2_2_15/i0[6] ), .A2(\SB2_2_15/i0[10] ), .A3(
        \SB2_2_15/i0_3 ), .ZN(\SB2_2_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U12761 ( .A1(\SB1_3_2/i0[6] ), .A2(\SB1_3_2/i0_4 ), .A3(
        \SB1_3_2/i0[9] ), .ZN(n3961) );
  NAND3_X2 U12762 ( .A1(\SB2_3_9/i0[9] ), .A2(\SB2_3_9/i0_3 ), .A3(
        \SB2_3_9/i0[8] ), .ZN(\SB2_3_9/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U12763 ( .A1(n7363), .A2(n7362), .Z(\MC_ARK_ARC_1_2/buf_output[104] ) );
  NAND3_X2 U12764 ( .A1(\SB1_2_0/i0[10] ), .A2(\SB1_2_0/i0_0 ), .A3(
        \SB1_2_0/i0[6] ), .ZN(\SB1_2_0/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U12765 ( .A1(n7348), .A2(\SB2_3_9/Component_Function_3/NAND4_in[0] ), .A3(\SB2_3_9/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_3_9/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_3_9/buf_output[3] ) );
  NAND3_X2 U12766 ( .A1(\SB2_3_24/i0[6] ), .A2(\SB2_3_24/i0_3 ), .A3(
        \SB2_3_24/i0[10] ), .ZN(\SB2_3_24/Component_Function_2/NAND4_in[1] )
         );
  NAND4_X2 U12767 ( .A1(n3940), .A2(
        \SB2_3_20/Component_Function_3/NAND4_in[0] ), .A3(n6810), .A4(
        \SB2_3_20/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_20/buf_output[3] ) );
  NAND4_X2 U12768 ( .A1(n1710), .A2(
        \SB1_2_26/Component_Function_5/NAND4_in[2] ), .A3(n6639), .A4(
        \SB1_2_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_26/buf_output[5] ) );
  NAND4_X2 U12769 ( .A1(\SB1_2_14/Component_Function_2/NAND4_in[0] ), .A2(
        n1855), .A3(n7201), .A4(n7202), .ZN(\SB1_2_14/buf_output[2] ) );
  NAND3_X1 U12770 ( .A1(\SB2_4_20/i0_3 ), .A2(\SB2_4_20/i0[10] ), .A3(
        \SB2_4_20/i0_4 ), .ZN(n1195) );
  NAND4_X2 U12771 ( .A1(\SB1_2_20/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_20/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_20/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_2_20/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_2_20/buf_output[0] ) );
  XOR2_X1 U12772 ( .A1(\RI5[4][96] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[120] ), 
        .Z(n3526) );
  XOR2_X1 U12773 ( .A1(n6503), .A2(\MC_ARK_ARC_1_1/temp3[55] ), .Z(n709) );
  XOR2_X1 U12774 ( .A1(\MC_ARK_ARC_1_2/temp3[175] ), .A2(
        \MC_ARK_ARC_1_2/temp1[175] ), .Z(n6500) );
  XOR2_X1 U12775 ( .A1(n1604), .A2(\MC_ARK_ARC_1_2/temp4[175] ), .Z(n6501) );
  XOR2_X1 U12776 ( .A1(\RI5[1][140] ), .A2(\RI5[1][176] ), .Z(
        \MC_ARK_ARC_1_1/temp3[74] ) );
  NAND4_X2 U12777 ( .A1(\SB2_1_31/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_1_31/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_31/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_1_31/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_31/buf_output[1] ) );
  NAND4_X2 U12778 ( .A1(\SB1_2_0/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_0/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_0/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_2_0/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_0/buf_output[1] ) );
  NAND4_X2 U12779 ( .A1(n4492), .A2(
        \SB2_2_15/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_15/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_2_15/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_15/buf_output[1] ) );
  NAND4_X2 U12780 ( .A1(\SB2_2_12/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_12/Component_Function_4/NAND4_in[0] ), .A3(n3688), .A4(
        \SB2_2_12/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_2_12/buf_output[4] ) );
  XOR2_X1 U12781 ( .A1(\SB2_1_31/buf_output[1] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[1] ), .Z(n6503) );
  NAND3_X2 U12782 ( .A1(\SB1_3_11/i0_4 ), .A2(\SB1_3_11/i1_5 ), .A3(
        \SB1_3_11/i1[9] ), .ZN(n6504) );
  XOR2_X1 U12783 ( .A1(\MC_ARK_ARC_1_4/temp4[116] ), .A2(n6505), .Z(n7085) );
  XOR2_X1 U12784 ( .A1(\RI5[4][116] ), .A2(\RI5[4][110] ), .Z(n6505) );
  NAND4_X2 U12785 ( .A1(n1133), .A2(
        \SB2_3_11/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_11/Component_Function_4/NAND4_in[1] ), .A4(n6506), .ZN(
        \SB2_3_11/buf_output[4] ) );
  NAND3_X1 U12786 ( .A1(\SB2_3_11/i0_4 ), .A2(\SB2_3_11/i1_5 ), .A3(
        \SB2_3_11/i1[9] ), .ZN(n6506) );
  NAND3_X2 U12787 ( .A1(\SB1_1_22/i0[6] ), .A2(\SB1_1_22/i0[10] ), .A3(
        \SB1_1_22/i0_0 ), .ZN(n6507) );
  XOR2_X1 U12788 ( .A1(\MC_ARK_ARC_1_2/temp1[139] ), .A2(n6508), .Z(
        \MC_ARK_ARC_1_2/temp5[139] ) );
  XOR2_X1 U12789 ( .A1(\RI5[2][109] ), .A2(\RI5[2][85] ), .Z(n6508) );
  NAND3_X1 U12790 ( .A1(\SB2_1_22/i0_0 ), .A2(\SB2_1_22/i0_4 ), .A3(
        \SB2_1_22/i1_5 ), .ZN(\SB2_1_22/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U12791 ( .A1(\MC_ARK_ARC_1_0/temp5[55] ), .A2(n6509), .Z(
        \MC_ARK_ARC_1_0/buf_output[55] ) );
  XOR2_X1 U12792 ( .A1(\MC_ARK_ARC_1_0/temp4[55] ), .A2(
        \MC_ARK_ARC_1_0/temp3[55] ), .Z(n6509) );
  NAND4_X2 U12793 ( .A1(\SB2_4_20/Component_Function_3/NAND4_in[0] ), .A2(
        n4900), .A3(\SB2_4_20/Component_Function_3/NAND4_in[2] ), .A4(n1208), 
        .ZN(\SB2_4_20/buf_output[3] ) );
  XOR2_X1 U12794 ( .A1(n6512), .A2(n6511), .Z(n1841) );
  XOR2_X1 U12795 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[140] ), .A2(n195), .Z(
        n6511) );
  XOR2_X1 U12796 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[170] ), .A2(\RI5[3][14] ), 
        .Z(n6512) );
  XOR2_X1 U12797 ( .A1(n6513), .A2(n98), .Z(Ciphertext[17]) );
  NAND4_X2 U12798 ( .A1(\SB4_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_29/Component_Function_5/NAND4_in[0] ), .A4(n2200), .ZN(n6513) );
  NAND4_X2 U12799 ( .A1(\SB3_11/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_0/NAND4_in[0] ), .A4(n6514), .ZN(
        \SB3_11/buf_output[0] ) );
  NAND4_X2 U12800 ( .A1(\SB4_17/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_17/Component_Function_0/NAND4_in[3] ), .A3(n5397), .A4(n6515), 
        .ZN(n6838) );
  NAND2_X1 U12801 ( .A1(\SB4_17/i0[9] ), .A2(\SB4_17/i0[10] ), .ZN(n6515) );
  NAND4_X2 U12802 ( .A1(\SB3_3/Component_Function_0/NAND4_in[1] ), .A2(
        \SB3_3/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_3/Component_Function_0/NAND4_in[0] ), .A4(n6516), .ZN(
        \SB3_3/buf_output[0] ) );
  XOR2_X1 U12803 ( .A1(n6518), .A2(n6519), .Z(\MC_ARK_ARC_1_3/buf_output[147] ) );
  NAND4_X2 U12804 ( .A1(\SB2_3_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_30/Component_Function_3/NAND4_in[3] ), .A3(n7063), .A4(n6520), 
        .ZN(\SB2_3_30/buf_output[3] ) );
  NAND3_X2 U12805 ( .A1(\SB2_3_30/i0[10] ), .A2(\SB2_3_30/i1[9] ), .A3(
        \SB2_3_30/i1_7 ), .ZN(n6520) );
  NAND4_X2 U12806 ( .A1(\SB1_2_14/Component_Function_1/NAND4_in[1] ), .A2(
        n5277), .A3(\SB1_2_14/Component_Function_1/NAND4_in[2] ), .A4(n6521), 
        .ZN(\SB1_2_14/buf_output[1] ) );
  NAND2_X2 U12807 ( .A1(\RI1[2][107] ), .A2(\SB1_2_14/i1[9] ), .ZN(n6521) );
  NAND3_X2 U12808 ( .A1(\SB1_1_0/i0[10] ), .A2(\SB1_1_0/i0_0 ), .A3(
        \SB1_1_0/i0[6] ), .ZN(n6522) );
  XOR2_X1 U12809 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[122] ), .A2(\RI5[2][128] ), .Z(n6523) );
  NAND3_X1 U12810 ( .A1(\SB1_3_24/i0_3 ), .A2(\SB1_3_24/i0_4 ), .A3(
        \SB1_3_24/i1[9] ), .ZN(\SB1_3_24/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U12811 ( .A1(\MC_ARK_ARC_1_2/temp1[15] ), .A2(n6524), .Z(
        \MC_ARK_ARC_1_2/temp5[15] ) );
  XOR2_X1 U12812 ( .A1(\RI5[2][153] ), .A2(\RI5[2][177] ), .Z(n6524) );
  NAND3_X2 U12813 ( .A1(\SB2_3_14/i0_3 ), .A2(\SB2_3_14/i0_0 ), .A3(
        \SB2_3_14/i0_4 ), .ZN(\SB2_3_14/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U12814 ( .A1(n7372), .A2(n4727), .ZN(n6597) );
  NAND3_X2 U12815 ( .A1(\SB1_1_8/i0[10] ), .A2(\SB1_1_8/i1_5 ), .A3(
        \SB1_1_8/i1[9] ), .ZN(\SB1_1_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U12816 ( .A1(\SB1_4_25/i1_5 ), .A2(\SB1_4_25/i1[9] ), .A3(
        \SB1_4_25/i0[10] ), .ZN(n6525) );
  INV_X2 U12817 ( .I(\SB1_1_4/buf_output[2] ), .ZN(\SB2_1_1/i1[9] ) );
  XOR2_X1 U12818 ( .A1(n6527), .A2(n6526), .Z(\MC_ARK_ARC_1_4/temp5[44] ) );
  XOR2_X1 U12819 ( .A1(\RI5[4][38] ), .A2(\RI5[4][182] ), .Z(n6527) );
  INV_X2 U12820 ( .I(\SB1_3_22/buf_output[2] ), .ZN(\SB2_3_19/i1[9] ) );
  NAND4_X2 U12821 ( .A1(\SB1_3_22/Component_Function_2/NAND4_in[1] ), .A2(
        n4334), .A3(\SB1_3_22/Component_Function_2/NAND4_in[3] ), .A4(n4347), 
        .ZN(\SB1_3_22/buf_output[2] ) );
  NAND3_X1 U12822 ( .A1(\SB1_3_10/i0_0 ), .A2(\SB1_3_10/i0[9] ), .A3(
        \SB1_3_10/i0[8] ), .ZN(\SB1_3_10/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U12823 ( .A1(\MC_ARK_ARC_1_4/temp4[27] ), .A2(
        \MC_ARK_ARC_1_4/temp3[27] ), .Z(n2142) );
  NAND4_X2 U12824 ( .A1(\SB1_0_13/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_13/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_3/NAND4_in[1] ), .ZN(\RI3[0][123] ) );
  NAND4_X2 U12825 ( .A1(\SB2_0_5/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_0_5/Component_Function_5/NAND4_in[1] ), .A3(n1771), .A4(
        \SB2_0_5/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_5/buf_output[5] ) );
  XOR2_X1 U12826 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[110] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[164] ), .Z(n4778) );
  NAND4_X2 U12827 ( .A1(\SB2_3_19/Component_Function_2/NAND4_in[0] ), .A2(
        n5075), .A3(\SB2_3_19/Component_Function_2/NAND4_in[2] ), .A4(n6529), 
        .ZN(\SB2_3_19/buf_output[2] ) );
  NAND3_X2 U12828 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB2_3_19/i0[10] ), .A3(
        \SB2_3_19/i0[6] ), .ZN(n6529) );
  NAND3_X1 U12829 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0[8] ), .A3(
        \SB1_0_25/i1_7 ), .ZN(\SB1_0_25/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U12830 ( .A1(n3394), .A2(n6530), .Z(\MC_ARK_ARC_1_3/buf_output[114] ) );
  XOR2_X1 U12831 ( .A1(n5353), .A2(n7279), .Z(n6530) );
  NAND2_X1 U12832 ( .A1(\SB4_23/i0[10] ), .A2(\SB4_23/i0[9] ), .ZN(
        \SB4_23/Component_Function_0/NAND4_in[0] ) );
  NAND2_X2 U12833 ( .A1(n3386), .A2(n3385), .ZN(\SB4_23/i0[10] ) );
  NOR2_X1 U12834 ( .A1(\RI1[4][17] ), .A2(\MC_ARK_ARC_1_3/buf_output[15] ), 
        .ZN(n6531) );
  XOR2_X1 U12835 ( .A1(n6532), .A2(n32), .Z(Ciphertext[61]) );
  NAND4_X2 U12836 ( .A1(\SB4_21/Component_Function_1/NAND4_in[1] ), .A2(n1254), 
        .A3(\SB4_21/Component_Function_1/NAND4_in[3] ), .A4(n1699), .ZN(n6532)
         );
  NAND2_X2 U12837 ( .A1(n2530), .A2(n7215), .ZN(\RI5[1][8] ) );
  NAND3_X1 U12838 ( .A1(\SB4_24/i0_4 ), .A2(\SB4_24/i0_0 ), .A3(\SB4_24/i1_5 ), 
        .ZN(n2745) );
  NAND2_X2 U12839 ( .A1(\SB2_0_31/i0_0 ), .A2(n6533), .ZN(
        \SB2_0_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U12840 ( .A1(\SB2_3_15/i0_4 ), .A2(\SB2_3_15/i0_3 ), .A3(
        \SB2_3_15/i0[10] ), .ZN(n6672) );
  NAND3_X2 U12841 ( .A1(\SB1_3_14/i1_5 ), .A2(\SB1_3_14/i0_0 ), .A3(
        \SB1_3_14/i0_4 ), .ZN(\SB1_3_14/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U12842 ( .A1(\RI5[3][149] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[155] ), .Z(n6534) );
  XOR2_X1 U12843 ( .A1(n7465), .A2(n6535), .Z(\MC_ARK_ARC_1_3/buf_output[180] ) );
  NAND3_X2 U12844 ( .A1(\SB2_3_7/i0[10] ), .A2(\SB2_3_7/i0_0 ), .A3(
        \SB2_3_7/i0[6] ), .ZN(\SB2_3_7/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U12845 ( .A1(\MC_ARK_ARC_1_2/temp5[135] ), .A2(n2227), .Z(
        \MC_ARK_ARC_1_2/buf_output[135] ) );
  INV_X2 U12846 ( .I(\SB1_4_14/buf_output[2] ), .ZN(\SB2_4_11/i1[9] ) );
  NAND4_X2 U12847 ( .A1(\SB2_2_12/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_2_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_12/Component_Function_1/NAND4_in[0] ), .A4(n6536), .ZN(
        \SB2_2_12/buf_output[1] ) );
  XOR2_X1 U12848 ( .A1(\MC_ARK_ARC_1_3/temp3[165] ), .A2(
        \MC_ARK_ARC_1_3/temp4[165] ), .Z(\MC_ARK_ARC_1_3/temp6[165] ) );
  XOR2_X1 U12849 ( .A1(\RI5[3][117] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_3/temp2[171] ) );
  XOR2_X1 U12850 ( .A1(n1719), .A2(n4988), .Z(\MC_ARK_ARC_1_2/buf_output[1] )
         );
  XOR2_X1 U12851 ( .A1(n7010), .A2(n2652), .Z(\MC_ARK_ARC_1_3/buf_output[73] )
         );
  XOR2_X1 U12852 ( .A1(\MC_ARK_ARC_1_4/temp1[181] ), .A2(
        \MC_ARK_ARC_1_4/temp2[181] ), .Z(n7153) );
  NAND2_X2 U12853 ( .A1(n5426), .A2(n6537), .ZN(\SB2_1_31/i0_4 ) );
  AND2_X1 U12854 ( .A1(\SB1_1_0/Component_Function_4/NAND4_in[3] ), .A2(n4996), 
        .Z(n6537) );
  NAND4_X2 U12855 ( .A1(\SB1_3_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_3/NAND4_in[2] ), .A3(n3697), .A4(n6538), 
        .ZN(\SB1_3_0/buf_output[3] ) );
  NAND3_X1 U12856 ( .A1(\SB2_4_21/i0[10] ), .A2(\SB2_4_21/i0_3 ), .A3(
        \SB1_4_25/buf_output[1] ), .ZN(n6539) );
  NAND4_X2 U12857 ( .A1(\SB1_2_11/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_11/Component_Function_5/NAND4_in[0] ), .A3(n2797), .A4(n6540), 
        .ZN(\SB1_2_11/buf_output[5] ) );
  NAND3_X2 U12858 ( .A1(\SB1_2_11/i0[9] ), .A2(\SB1_2_11/i0[6] ), .A3(
        \SB1_2_11/i0_4 ), .ZN(n6540) );
  NAND3_X2 U12859 ( .A1(\SB2_3_3/i0[10] ), .A2(\SB2_3_3/i1_5 ), .A3(
        \SB2_3_3/i1[9] ), .ZN(\SB2_3_3/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U12860 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[147] ), .A2(n516), .Z(
        n6543) );
  XOR2_X1 U12861 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[183] ), .A2(\RI5[3][117] ), .Z(n6544) );
  NAND3_X2 U12862 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0[10] ), .A3(
        \SB2_3_0/i0[6] ), .ZN(\SB2_3_0/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U12863 ( .A1(n6766), .A2(\SB2_2_2/Component_Function_2/NAND4_in[0] ), .A3(\SB2_2_2/Component_Function_2/NAND4_in[2] ), .A4(n6545), .ZN(
        \SB2_2_2/buf_output[2] ) );
  NAND3_X2 U12864 ( .A1(\SB2_2_2/i0_3 ), .A2(\SB2_2_2/i0[10] ), .A3(
        \SB2_2_2/i0[6] ), .ZN(n6545) );
  NAND4_X2 U12865 ( .A1(\SB1_2_1/Component_Function_5/NAND4_in[1] ), .A2(n3209), .A3(n6727), .A4(\SB1_2_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_1/buf_output[5] ) );
  NAND4_X2 U12866 ( .A1(\SB3_26/Component_Function_2/NAND4_in[0] ), .A2(n6926), 
        .A3(\SB3_26/Component_Function_2/NAND4_in[1] ), .A4(n7293), .ZN(
        \SB3_26/buf_output[2] ) );
  XOR2_X1 U12867 ( .A1(\MC_ARK_ARC_1_2/temp2[48] ), .A2(n6738), .Z(
        \MC_ARK_ARC_1_2/temp5[48] ) );
  NAND4_X2 U12868 ( .A1(\SB3_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_3/NAND4_in[3] ), .A4(
        \SB3_26/Component_Function_3/NAND4_in[2] ), .ZN(\SB3_26/buf_output[3] ) );
  NAND4_X2 U12869 ( .A1(n886), .A2(n2879), .A3(n7344), .A4(
        \SB3_26/Component_Function_5/NAND4_in[1] ), .ZN(\SB3_26/buf_output[5] ) );
  NAND3_X1 U12870 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i1_7 ), .A3(
        \SB4_11/i1[9] ), .ZN(n6546) );
  NAND3_X1 U12871 ( .A1(\SB1_3_8/i0_0 ), .A2(\SB1_3_8/i3[0] ), .A3(
        \SB1_3_8/i1_7 ), .ZN(n6547) );
  NAND4_X2 U12872 ( .A1(\SB2_3_16/Component_Function_5/NAND4_in[2] ), .A2(
        n4909), .A3(n4137), .A4(n4853), .ZN(\SB2_3_16/buf_output[5] ) );
  NAND3_X2 U12873 ( .A1(\SB2_0_7/i0[10] ), .A2(\SB2_0_7/i1[9] ), .A3(
        \SB2_0_7/i1_7 ), .ZN(\SB2_0_7/Component_Function_3/NAND4_in[2] ) );
  INV_X2 U12874 ( .I(n6548), .ZN(n5425) );
  NAND3_X2 U12875 ( .A1(\SB2_4_15/i0_0 ), .A2(\SB2_4_15/i0[10] ), .A3(
        \SB2_4_15/i0[6] ), .ZN(n6549) );
  INV_X2 U12876 ( .I(\SB1_4_23/buf_output[3] ), .ZN(\SB2_4_21/i0[8] ) );
  NAND4_X2 U12877 ( .A1(\SB1_4_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_4_23/Component_Function_3/NAND4_in[1] ), .A3(n6572), .A4(n3376), 
        .ZN(\SB1_4_23/buf_output[3] ) );
  XOR2_X1 U12878 ( .A1(n6550), .A2(n165), .Z(Ciphertext[101]) );
  NAND4_X2 U12879 ( .A1(\SB4_15/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_15/Component_Function_5/NAND4_in[3] ), .A3(n2664), .A4(
        \SB4_15/Component_Function_5/NAND4_in[0] ), .ZN(n6550) );
  NAND2_X1 U12880 ( .A1(\SB1_2_11/i1[9] ), .A2(\SB1_2_11/i0_3 ), .ZN(
        \SB1_2_11/Component_Function_1/NAND4_in[0] ) );
  NAND2_X2 U12881 ( .A1(\SB2_4_15/i0_0 ), .A2(\SB2_4_15/i3[0] ), .ZN(n6551) );
  BUF_X2 U12882 ( .I(\SB1_3_1/buf_output[1] ), .Z(n6552) );
  NAND3_X1 U12883 ( .A1(\SB1_0_27/i0_4 ), .A2(\SB1_0_27/i0[8] ), .A3(
        \SB1_0_27/i1_7 ), .ZN(n6553) );
  XOR2_X1 U12884 ( .A1(n6554), .A2(\MC_ARK_ARC_1_0/temp4[140] ), .Z(n3521) );
  NAND4_X2 U12885 ( .A1(\SB1_0_29/Component_Function_2/NAND4_in[0] ), .A2(
        n4621), .A3(\SB1_0_29/Component_Function_2/NAND4_in[2] ), .A4(n6556), 
        .ZN(\SB1_0_29/buf_output[2] ) );
  NAND3_X2 U12886 ( .A1(\SB1_0_29/i0_0 ), .A2(\SB1_0_29/i0_4 ), .A3(
        \SB1_0_29/i1_5 ), .ZN(n6556) );
  NAND3_X2 U12887 ( .A1(\SB2_3_8/i0_4 ), .A2(\SB2_3_8/i0_3 ), .A3(
        \SB2_3_8/i1[9] ), .ZN(\SB2_3_8/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U12888 ( .A1(\SB1_3_11/Component_Function_2/NAND4_in[1] ), .A2(
        n7185), .A3(\SB1_3_11/Component_Function_2/NAND4_in[3] ), .A4(n6557), 
        .ZN(\SB1_3_11/buf_output[2] ) );
  XOR2_X1 U12889 ( .A1(\RI5[4][66] ), .A2(\RI5[4][42] ), .Z(n6558) );
  NAND4_X2 U12890 ( .A1(\SB2_1_25/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_25/Component_Function_2/NAND4_in[0] ), .A3(n4622), .A4(n6559), 
        .ZN(\SB2_1_25/buf_output[2] ) );
  NAND3_X2 U12891 ( .A1(\SB2_1_25/i0_4 ), .A2(\SB2_1_25/i0_0 ), .A3(
        \SB2_1_25/i1_5 ), .ZN(n6559) );
  NAND3_X1 U12892 ( .A1(\SB3_6/i1_7 ), .A2(\SB3_6/i0[8] ), .A3(\SB3_6/i0_3 ), 
        .ZN(\SB3_6/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U12893 ( .A1(\SB2_4_25/Component_Function_4/NAND4_in[0] ), .A2(n744), .A3(n7044), .A4(\SB2_4_25/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_4_25/buf_output[4] ) );
  NAND3_X2 U12894 ( .A1(\SB1_4_25/i0_3 ), .A2(\SB1_4_25/i0[6] ), .A3(
        \SB1_4_25/i0[10] ), .ZN(\SB1_4_25/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U12895 ( .A1(\MC_ARK_ARC_1_0/temp3[27] ), .A2(n7415), .Z(n6560) );
  NAND4_X2 U12896 ( .A1(\SB2_4_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_3/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_4_3/Component_Function_3/NAND4_in[1] ), .A4(n6561), .ZN(
        \SB2_4_3/buf_output[3] ) );
  NAND3_X2 U12897 ( .A1(\SB2_4_3/i0[10] ), .A2(\SB2_4_3/i1_7 ), .A3(
        \SB2_4_3/i1[9] ), .ZN(n6561) );
  NAND3_X2 U12898 ( .A1(\SB2_3_8/i0[10] ), .A2(\SB2_3_8/i0[6] ), .A3(
        \SB2_3_8/i0_3 ), .ZN(n6562) );
  NAND4_X2 U12899 ( .A1(\SB2_2_13/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_2_13/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_13/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_2_13/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_13/buf_output[5] ) );
  NAND3_X1 U12900 ( .A1(\SB1_3_11/i0[9] ), .A2(\SB1_3_11/i0_0 ), .A3(
        \SB1_3_11/i0[8] ), .ZN(n6563) );
  XOR2_X1 U12901 ( .A1(n6565), .A2(n6564), .Z(n4419) );
  XOR2_X1 U12902 ( .A1(\RI5[3][65] ), .A2(n456), .Z(n6564) );
  XOR2_X1 U12903 ( .A1(\RI5[3][191] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[29] ), 
        .Z(n6565) );
  NAND4_X2 U12904 ( .A1(\SB1_4_29/Component_Function_3/NAND4_in[3] ), .A2(
        n4132), .A3(\SB1_4_29/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_4_29/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB1_4_29/buf_output[3] ) );
  NAND4_X2 U12905 ( .A1(\SB2_0_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_2/NAND4_in[3] ), .A4(n6566), .ZN(
        \SB2_0_29/buf_output[2] ) );
  NAND3_X2 U12906 ( .A1(\SB2_0_29/i0_3 ), .A2(\SB2_0_29/i0[9] ), .A3(
        \SB2_0_29/i0[8] ), .ZN(n6566) );
  NAND4_X2 U12907 ( .A1(\SB1_0_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_29/Component_Function_5/NAND4_in[0] ), .A4(n6567), .ZN(
        \SB1_0_29/buf_output[5] ) );
  NAND3_X1 U12908 ( .A1(\SB1_0_29/i0[6] ), .A2(\SB1_0_29/i0[9] ), .A3(n322), 
        .ZN(n6567) );
  NAND4_X2 U12909 ( .A1(\SB2_0_29/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_29/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_29/Component_Function_3/NAND4_in[1] ), .A4(n6568), .ZN(
        \SB2_0_29/buf_output[3] ) );
  NAND3_X2 U12910 ( .A1(\SB2_0_29/i0_3 ), .A2(\SB2_0_29/i0[6] ), .A3(
        \SB2_0_29/i1[9] ), .ZN(n6568) );
  NAND4_X2 U12911 ( .A1(\SB2_1_17/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_1_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_17/Component_Function_3/NAND4_in[0] ), .A4(n6569), .ZN(
        \SB2_1_17/buf_output[3] ) );
  XOR2_X1 U12912 ( .A1(\RI5[1][17] ), .A2(\RI5[1][41] ), .Z(
        \MC_ARK_ARC_1_1/temp2[71] ) );
  XOR2_X1 U12913 ( .A1(n7484), .A2(n6570), .Z(\MC_ARK_ARC_1_1/buf_output[33] )
         );
  XOR2_X1 U12914 ( .A1(\MC_ARK_ARC_1_1/temp3[33] ), .A2(
        \MC_ARK_ARC_1_1/temp4[33] ), .Z(n6570) );
  NAND4_X2 U12915 ( .A1(\SB2_4_7/Component_Function_0/NAND4_in[2] ), .A2(n1808), .A3(\SB2_4_7/Component_Function_0/NAND4_in[0] ), .A4(n6571), .ZN(
        \SB2_4_7/buf_output[0] ) );
  INV_X2 U12916 ( .I(\SB1_1_27/buf_output[2] ), .ZN(\SB2_1_24/i1[9] ) );
  NAND4_X2 U12917 ( .A1(n5350), .A2(n4554), .A3(
        \SB1_1_27/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_27/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_1_27/buf_output[2] ) );
  NAND3_X1 U12918 ( .A1(\SB1_4_23/i0[8] ), .A2(\SB1_4_23/i3[0] ), .A3(
        \SB1_4_23/i1_5 ), .ZN(n6572) );
  NAND4_X2 U12919 ( .A1(n2578), .A2(
        \SB2_3_15/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_3_15/Component_Function_2/NAND4_in[0] ), .A4(n6573), .ZN(
        \SB2_3_15/buf_output[2] ) );
  NAND3_X2 U12920 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0[6] ), .A3(
        \SB2_3_15/i0[10] ), .ZN(n6573) );
  NAND3_X2 U12921 ( .A1(\SB2_1_14/Component_Function_5/NAND4_in[2] ), .A2(
        n6652), .A3(\SB2_1_14/Component_Function_5/NAND4_in[1] ), .ZN(
        \SB2_1_14/buf_output[5] ) );
  NAND3_X1 U12922 ( .A1(\SB1_2_22/i0_0 ), .A2(\RI1[2][59] ), .A3(
        \MC_ARK_ARC_1_1/buf_output[58] ), .ZN(n4121) );
  NAND4_X2 U12923 ( .A1(n2653), .A2(
        \SB1_3_31/Component_Function_4/NAND4_in[0] ), .A3(n2984), .A4(n6575), 
        .ZN(\SB1_3_31/buf_output[4] ) );
  NAND4_X2 U12924 ( .A1(\SB1_0_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_17/Component_Function_3/NAND4_in[3] ), .A4(n6576), .ZN(
        \RI3[0][99] ) );
  XOR2_X1 U12925 ( .A1(\RI5[0][107] ), .A2(\RI5[0][101] ), .Z(n4086) );
  NAND4_X2 U12926 ( .A1(n2569), .A2(n1485), .A3(
        \SB1_0_17/Component_Function_2/NAND4_in[2] ), .A4(n6577), .ZN(
        \SB1_0_17/buf_output[2] ) );
  NAND3_X2 U12927 ( .A1(\SB1_0_17/i0[10] ), .A2(\SB1_0_17/i0_3 ), .A3(
        \SB1_0_17/i0[6] ), .ZN(n6577) );
  INV_X2 U12928 ( .I(\RI3[0][38] ), .ZN(\SB2_0_25/i1[9] ) );
  XOR2_X1 U12929 ( .A1(\RI5[1][26] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[152] ), 
        .Z(n6578) );
  NAND4_X2 U12930 ( .A1(\SB1_2_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_2_21/Component_Function_4/NAND4_in[1] ), .A4(n6579), .ZN(
        \SB1_2_21/buf_output[4] ) );
  NAND4_X2 U12931 ( .A1(\SB1_0_0/Component_Function_2/NAND4_in[0] ), .A2(n2772), .A3(n1552), .A4(n6580), .ZN(\SB1_0_0/buf_output[2] ) );
  NAND3_X1 U12932 ( .A1(\SB1_0_0/i0_3 ), .A2(n315), .A3(\SB1_0_0/i0[8] ), .ZN(
        n6580) );
  BUF_X4 U12933 ( .I(\SB2_2_26/i0_4 ), .Z(n6686) );
  NAND2_X1 U12934 ( .A1(\SB1_0_6/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_6/Component_Function_4/NAND4_in[3] ), .ZN(n6598) );
  NAND4_X2 U12935 ( .A1(n3131), .A2(n2071), .A3(
        \SB2_2_31/Component_Function_5/NAND4_in[0] ), .A4(n6581), .ZN(
        \SB2_2_31/buf_output[5] ) );
  NAND3_X2 U12936 ( .A1(\SB2_2_31/i0[9] ), .A2(\SB2_2_31/i0_4 ), .A3(
        \SB2_2_31/i0[6] ), .ZN(n6581) );
  NAND4_X2 U12937 ( .A1(n4100), .A2(n2175), .A3(
        \SB2_2_27/Component_Function_5/NAND4_in[0] ), .A4(n6582), .ZN(
        \SB2_2_27/buf_output[5] ) );
  NAND3_X2 U12938 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i0_0 ), .A3(
        \SB2_2_27/i0[6] ), .ZN(n6582) );
  NAND4_X2 U12939 ( .A1(\SB1_2_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_4/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_4/buf_output[1] ) );
  NAND3_X2 U12940 ( .A1(\SB2_1_27/i1[9] ), .A2(\SB2_1_27/i1_5 ), .A3(
        \SB2_1_27/i0[10] ), .ZN(\SB2_1_27/Component_Function_2/NAND4_in[0] )
         );
  XOR2_X1 U12941 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), .A2(\RI5[3][191] ), .Z(\MC_ARK_ARC_1_3/temp3[89] ) );
  NAND3_X2 U12942 ( .A1(\SB2_4_28/i0[6] ), .A2(\SB2_4_28/i0_4 ), .A3(
        \SB2_4_28/i0[9] ), .ZN(n4530) );
  XOR2_X1 U12943 ( .A1(\RI5[3][63] ), .A2(\RI5[3][33] ), .Z(n4118) );
  NAND4_X2 U12944 ( .A1(\SB1_0_30/Component_Function_2/NAND4_in[0] ), .A2(
        n7515), .A3(\SB1_0_30/Component_Function_2/NAND4_in[2] ), .A4(n6583), 
        .ZN(\SB1_0_30/buf_output[2] ) );
  NAND3_X2 U12945 ( .A1(\SB1_0_30/i0[6] ), .A2(\SB1_0_30/i0[10] ), .A3(
        \SB1_0_30/i0_3 ), .ZN(n6583) );
  INV_X2 U12946 ( .I(n6584), .ZN(\SB1_1_27/buf_output[3] ) );
  AND4_X1 U12947 ( .A1(\SB1_1_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_27/Component_Function_3/NAND4_in[3] ), .A4(n4067), .Z(n6584) );
  XOR2_X1 U12948 ( .A1(\MC_ARK_ARC_1_3/temp4[7] ), .A2(
        \MC_ARK_ARC_1_3/temp3[7] ), .Z(\MC_ARK_ARC_1_3/temp6[7] ) );
  XOR2_X1 U12949 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[89] ), .A2(\RI5[2][113] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[143] ) );
  NAND4_X2 U12950 ( .A1(\SB2_2_11/Component_Function_5/NAND4_in[3] ), .A2(
        n1766), .A3(n6617), .A4(n6775), .ZN(\SB2_2_11/buf_output[5] ) );
  NAND3_X2 U12951 ( .A1(\SB1_1_30/i0_0 ), .A2(\SB1_1_30/i1_5 ), .A3(
        \SB1_1_30/i0_4 ), .ZN(n3109) );
  NAND3_X1 U12952 ( .A1(\SB1_4_30/i0[6] ), .A2(\SB1_4_30/i0_3 ), .A3(
        \SB1_4_30/i1[9] ), .ZN(\SB1_4_30/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U12953 ( .A1(n2967), .A2(\SB1_4_0/Component_Function_3/NAND4_in[3] ), .A3(n4746), .A4(n4462), .ZN(\SB1_4_0/buf_output[3] ) );
  NAND4_X2 U12954 ( .A1(\SB2_3_29/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_29/Component_Function_1/NAND4_in[3] ), .A3(n4793), .A4(
        \SB2_3_29/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_29/buf_output[1] ) );
  AND2_X1 U12955 ( .A1(\MC_ARK_ARC_1_0/buf_output[25] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[28] ), .Z(n6586) );
  NAND3_X2 U12956 ( .A1(\SB1_3_1/i0[9] ), .A2(\SB1_3_1/i0[8] ), .A3(
        \SB1_3_1/i0_3 ), .ZN(n6587) );
  XOR2_X1 U12957 ( .A1(\RI5[0][165] ), .A2(\RI5[0][27] ), .Z(n6588) );
  NAND3_X1 U12958 ( .A1(\SB2_4_6/i0[8] ), .A2(\SB2_4_6/i1_7 ), .A3(
        \SB1_4_7/buf_output[4] ), .ZN(
        \SB2_4_6/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U12959 ( .A1(\SB3_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_1/Component_Function_1/NAND4_in[2] ), .A3(
        \SB3_1/Component_Function_1/NAND4_in[0] ), .A4(n6589), .ZN(
        \SB3_1/buf_output[1] ) );
  XOR2_X1 U12960 ( .A1(\MC_ARK_ARC_1_4/temp1[50] ), .A2(n6590), .Z(n6827) );
  XOR2_X1 U12961 ( .A1(\RI5[4][20] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[188] ), 
        .Z(n6590) );
  NAND3_X2 U12962 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0[10] ), .A3(
        \SB2_0_5/i0[9] ), .ZN(n1239) );
  XOR2_X1 U12963 ( .A1(n6592), .A2(n6591), .Z(\RI1[5][107] ) );
  XOR2_X1 U12964 ( .A1(n7419), .A2(\MC_ARK_ARC_1_4/temp4[107] ), .Z(n6591) );
  XOR2_X1 U12965 ( .A1(\MC_ARK_ARC_1_4/temp3[107] ), .A2(n7334), .Z(n6592) );
  XOR2_X1 U12966 ( .A1(n4075), .A2(n6593), .Z(n3683) );
  XOR2_X1 U12967 ( .A1(\RI5[1][179] ), .A2(\RI5[1][23] ), .Z(n6593) );
  XOR2_X1 U12968 ( .A1(\SB2_3_4/buf_output[3] ), .A2(\SB2_3_0/buf_output[3] ), 
        .Z(n6594) );
  NAND4_X2 U12969 ( .A1(\SB1_4_16/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_4_16/Component_Function_1/NAND4_in[0] ), .A3(n6611), .A4(
        \SB1_4_16/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_4_16/buf_output[1] ) );
  XOR2_X1 U12970 ( .A1(\MC_ARK_ARC_1_2/temp6[103] ), .A2(n6595), .Z(
        \MC_ARK_ARC_1_2/buf_output[103] ) );
  NAND4_X2 U12971 ( .A1(\SB2_2_26/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_26/Component_Function_2/NAND4_in[2] ), .A4(n6596), .ZN(
        \SB2_2_26/buf_output[2] ) );
  NAND3_X2 U12972 ( .A1(n6686), .A2(\SB2_2_26/i0_0 ), .A3(\SB2_2_26/i1_5 ), 
        .ZN(n6596) );
  INV_X1 U12973 ( .I(\SB1_2_27/buf_output[1] ), .ZN(\SB2_2_23/i1_7 ) );
  NAND4_X2 U12974 ( .A1(\SB1_2_27/Component_Function_1/NAND4_in[1] ), .A2(
        n7331), .A3(\SB1_2_27/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_2_27/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_27/buf_output[1] ) );
  NOR2_X2 U12975 ( .A1(n6598), .A2(n6597), .ZN(n2381) );
  NAND3_X2 U12976 ( .A1(\SB1_2_22/i1_5 ), .A2(\SB1_2_22/i1[9] ), .A3(
        \SB1_2_22/i0[10] ), .ZN(n6599) );
  INV_X2 U12977 ( .I(\SB1_2_30/buf_output[3] ), .ZN(\SB2_2_28/i0[8] ) );
  NAND4_X2 U12978 ( .A1(\SB1_2_30/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_30/Component_Function_3/NAND4_in[0] ), .A3(n7129), .A4(
        \SB1_2_30/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_30/buf_output[3] ) );
  INV_X2 U12979 ( .I(\SB1_1_2/buf_output[5] ), .ZN(\SB2_1_2/i1_5 ) );
  NAND4_X2 U12980 ( .A1(\SB2_3_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_28/Component_Function_3/NAND4_in[2] ), .A3(n5296), .A4(n7037), 
        .ZN(\SB2_3_28/buf_output[3] ) );
  NAND4_X2 U12981 ( .A1(\SB2_1_2/Component_Function_2/NAND4_in[2] ), .A2(n3452), .A3(\SB2_1_2/Component_Function_2/NAND4_in[3] ), .A4(n6601), .ZN(
        \SB2_1_2/buf_output[2] ) );
  NAND4_X2 U12982 ( .A1(\SB2_2_26/Component_Function_0/NAND4_in[1] ), .A2(
        n2322), .A3(\SB2_2_26/Component_Function_0/NAND4_in[0] ), .A4(n6602), 
        .ZN(\SB2_2_26/buf_output[0] ) );
  NAND3_X2 U12983 ( .A1(n6686), .A2(\SB2_2_26/i0_3 ), .A3(\SB2_2_26/i0_0 ), 
        .ZN(n6603) );
  NAND4_X2 U12984 ( .A1(n684), .A2(n2150), .A3(
        \SB1_3_6/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_3_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_6/buf_output[5] ) );
  XOR2_X1 U12985 ( .A1(n6605), .A2(n6604), .Z(n7148) );
  XOR2_X1 U12986 ( .A1(\RI5[0][155] ), .A2(n468), .Z(n6604) );
  XOR2_X1 U12987 ( .A1(\RI5[0][53] ), .A2(\RI5[0][179] ), .Z(n6605) );
  XOR2_X1 U12988 ( .A1(\MC_ARK_ARC_1_2/temp5[44] ), .A2(n2137), .Z(
        \MC_ARK_ARC_1_2/buf_output[44] ) );
  NAND4_X2 U12989 ( .A1(\SB2_1_15/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_15/Component_Function_5/NAND4_in[3] ), .A3(n6702), .A4(
        \SB2_1_15/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_15/buf_output[5] ) );
  XOR2_X1 U12990 ( .A1(\RI5[4][101] ), .A2(\RI5[4][71] ), .Z(n7468) );
  NAND4_X2 U12991 ( .A1(\SB2_0_6/Component_Function_5/NAND4_in[2] ), .A2(n2437), .A3(n6990), .A4(\SB2_0_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_6/buf_output[5] ) );
  XOR2_X1 U12992 ( .A1(n6606), .A2(\MC_ARK_ARC_1_2/temp6[153] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[153] ) );
  XOR2_X1 U12993 ( .A1(\MC_ARK_ARC_1_2/temp2[153] ), .A2(
        \MC_ARK_ARC_1_2/temp1[153] ), .Z(n6606) );
  NAND4_X2 U12994 ( .A1(\SB1_2_14/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_2_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_14/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_2_14/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_2_14/buf_output[4] ) );
  NAND4_X2 U12995 ( .A1(\SB1_1_11/Component_Function_2/NAND4_in[1] ), .A2(
        n4016), .A3(\SB1_1_11/Component_Function_2/NAND4_in[0] ), .A4(n6607), 
        .ZN(\SB1_1_11/buf_output[2] ) );
  NAND3_X2 U12996 ( .A1(\SB1_1_11/i0_0 ), .A2(\SB1_1_11/i1_5 ), .A3(
        \SB1_1_11/i0_4 ), .ZN(n6607) );
  NAND4_X2 U12997 ( .A1(\SB2_1_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_3/NAND4_in[2] ), .A3(n4470), .A4(n6608), 
        .ZN(\SB2_1_30/buf_output[3] ) );
  NAND3_X2 U12998 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i0_4 ), .A3(
        \SB2_1_30/i0_0 ), .ZN(n6608) );
  NAND3_X2 U12999 ( .A1(\SB1_0_16/i0[6] ), .A2(\SB1_0_16/i0_4 ), .A3(
        \SB1_0_16/i0[9] ), .ZN(n1862) );
  XOR2_X1 U13000 ( .A1(n6610), .A2(n6609), .Z(\MC_ARK_ARC_1_0/buf_output[14] )
         );
  XOR2_X1 U13001 ( .A1(\MC_ARK_ARC_1_0/temp4[14] ), .A2(
        \MC_ARK_ARC_1_0/temp2[14] ), .Z(n6609) );
  XOR2_X1 U13002 ( .A1(\MC_ARK_ARC_1_0/temp3[14] ), .A2(
        \MC_ARK_ARC_1_0/temp1[14] ), .Z(n6610) );
  XOR2_X1 U13003 ( .A1(\MC_ARK_ARC_1_0/temp3[127] ), .A2(
        \MC_ARK_ARC_1_0/temp4[127] ), .Z(\MC_ARK_ARC_1_0/temp6[127] ) );
  NOR2_X2 U13004 ( .A1(n7277), .A2(n6673), .ZN(n6612) );
  NAND3_X1 U13005 ( .A1(\SB2_4_5/i0[6] ), .A2(\SB2_4_5/i0[9] ), .A3(
        \SB2_4_5/i1_5 ), .ZN(\SB2_4_5/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U13006 ( .A1(\RI5[0][116] ), .A2(\RI5[0][122] ), .Z(
        \MC_ARK_ARC_1_0/temp1[122] ) );
  NAND4_X2 U13007 ( .A1(\SB1_2_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_26/Component_Function_1/NAND4_in[3] ), .A4(n6613), .ZN(
        \SB1_2_26/buf_output[1] ) );
  NAND3_X2 U13008 ( .A1(\SB1_2_26/i0[9] ), .A2(\SB1_2_26/i0[6] ), .A3(
        \SB1_2_26/i1_5 ), .ZN(n6613) );
  NAND3_X2 U13009 ( .A1(\SB1_4_7/i0_3 ), .A2(\SB1_4_7/i0[6] ), .A3(
        \SB1_4_7/i1[9] ), .ZN(n7537) );
  INV_X2 U13010 ( .I(\SB1_3_25/buf_output[2] ), .ZN(\SB2_3_22/i1[9] ) );
  NAND4_X2 U13011 ( .A1(\SB1_3_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_25/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_3_25/Component_Function_2/NAND4_in[1] ), .A4(n3866), .ZN(
        \SB1_3_25/buf_output[2] ) );
  XOR2_X1 U13012 ( .A1(\MC_ARK_ARC_1_3/temp2[114] ), .A2(n1077), .Z(n3394) );
  NAND2_X2 U13013 ( .A1(n7311), .A2(n5439), .ZN(\SB2_2_26/i0_4 ) );
  XOR2_X1 U13014 ( .A1(n2520), .A2(n6615), .Z(\MC_ARK_ARC_1_0/buf_output[1] )
         );
  NAND3_X2 U13015 ( .A1(\SB2_2_26/i0[8] ), .A2(n6686), .A3(\SB2_2_26/i1_7 ), 
        .ZN(n7414) );
  NAND3_X1 U13016 ( .A1(\SB1_3_17/i1_7 ), .A2(\SB1_3_17/i0_0 ), .A3(
        \SB1_3_17/i3[0] ), .ZN(\SB1_3_17/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U13017 ( .A1(\MC_ARK_ARC_1_3/temp5[8] ), .A2(
        \MC_ARK_ARC_1_3/temp6[8] ), .Z(\MC_ARK_ARC_1_3/buf_output[8] ) );
  NAND3_X1 U13018 ( .A1(\SB2_0_5/i0[9] ), .A2(\SB2_0_5/i0_4 ), .A3(
        \SB2_0_5/i0[6] ), .ZN(\SB2_0_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U13019 ( .A1(\SB2_2_11/i0[10] ), .A2(\SB2_2_11/i0_0 ), .A3(
        \SB2_2_11/i0[6] ), .ZN(n6617) );
  XOR2_X1 U13020 ( .A1(\RI5[2][113] ), .A2(\RI5[2][149] ), .Z(
        \MC_ARK_ARC_1_2/temp3[47] ) );
  XOR2_X1 U13021 ( .A1(n6618), .A2(n138), .Z(Ciphertext[140]) );
  NAND4_X2 U13022 ( .A1(\SB4_8/Component_Function_2/NAND4_in[2] ), .A2(n4378), 
        .A3(n4332), .A4(n1642), .ZN(n6618) );
  XOR2_X1 U13023 ( .A1(\MC_ARK_ARC_1_2/temp5[36] ), .A2(n6619), .Z(
        \MC_ARK_ARC_1_2/buf_output[36] ) );
  XOR2_X1 U13024 ( .A1(\MC_ARK_ARC_1_2/temp4[36] ), .A2(
        \MC_ARK_ARC_1_2/temp3[36] ), .Z(n6619) );
  XOR2_X1 U13025 ( .A1(\RI5[4][5] ), .A2(\RI5[4][191] ), .Z(n4367) );
  XOR2_X1 U13026 ( .A1(\RI5[1][25] ), .A2(\RI5[1][181] ), .Z(n7565) );
  NAND3_X2 U13027 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i0_0 ), .A3(
        \SB2_0_25/i0_4 ), .ZN(\SB2_0_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U13028 ( .A1(\SB1_1_24/i0[10] ), .A2(\SB1_1_24/i0[6] ), .A3(
        \SB1_1_24/i0_0 ), .ZN(n6621) );
  XOR2_X1 U13029 ( .A1(n1191), .A2(n4799), .Z(n7010) );
  NAND3_X2 U13030 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0[6] ), .A3(
        \SB2_2_4/i1[9] ), .ZN(n6622) );
  XOR2_X1 U13031 ( .A1(\MC_ARK_ARC_1_1/temp3[112] ), .A2(
        \MC_ARK_ARC_1_1/temp4[112] ), .Z(n6623) );
  NAND2_X2 U13032 ( .A1(n4840), .A2(\SB2_1_1/i0_3 ), .ZN(n7215) );
  NAND3_X1 U13033 ( .A1(\SB4_7/i1_7 ), .A2(\SB4_7/i3[0] ), .A3(\SB4_7/i0_0 ), 
        .ZN(\SB4_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U13034 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0_0 ), .A3(
        \SB1_0_25/i0_4 ), .ZN(\SB1_0_25/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U13035 ( .A1(n6624), .A2(n161), .Z(Ciphertext[147]) );
  NAND4_X2 U13036 ( .A1(n3006), .A2(\SB4_7/Component_Function_3/NAND4_in[0] ), 
        .A3(\SB4_7/Component_Function_3/NAND4_in[3] ), .A4(n4862), .ZN(n6624)
         );
  NAND3_X2 U13037 ( .A1(\SB2_0_29/i0_3 ), .A2(\SB2_0_29/i0_4 ), .A3(
        \SB2_0_29/i1[9] ), .ZN(\SB2_0_29/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U13038 ( .A1(\SB3_0/Component_Function_5/NAND4_in[1] ), .A2(n7145), 
        .A3(n3309), .A4(\SB3_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_0/buf_output[5] ) );
  NAND4_X2 U13039 ( .A1(\SB2_4_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_7/Component_Function_3/NAND4_in[2] ), .A3(n2228), .A4(n6625), 
        .ZN(\SB2_4_7/buf_output[3] ) );
  NAND3_X2 U13040 ( .A1(\SB2_4_7/i0_3 ), .A2(\SB2_4_7/i0_0 ), .A3(
        \RI3[4][148] ), .ZN(n6625) );
  NAND3_X2 U13041 ( .A1(\SB1_3_2/i0_0 ), .A2(\SB1_3_2/i0_3 ), .A3(
        \SB1_3_2/i0[7] ), .ZN(n6634) );
  XOR2_X1 U13042 ( .A1(n4007), .A2(n6626), .Z(\MC_ARK_ARC_1_2/buf_output[179] ) );
  NAND3_X1 U13043 ( .A1(\SB2_1_12/i0[6] ), .A2(\SB2_1_12/i0[9] ), .A3(
        \SB2_1_12/i1_5 ), .ZN(\SB2_1_12/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U13044 ( .A1(n5232), .A2(
        \SB2_3_28/Component_Function_4/NAND4_in[0] ), .A3(n3227), .A4(n6628), 
        .ZN(\SB2_3_28/buf_output[4] ) );
  NAND3_X1 U13045 ( .A1(\SB2_3_28/i0_3 ), .A2(\SB1_3_1/buf_output[0] ), .A3(
        \SB2_3_28/i0[10] ), .ZN(n6628) );
  NAND3_X1 U13046 ( .A1(\SB2_2_11/i0[6] ), .A2(\SB2_2_11/i1_5 ), .A3(
        \SB2_2_11/i0[9] ), .ZN(\SB2_2_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U13047 ( .A1(\SB2_2_25/i0[6] ), .A2(\SB2_2_25/i0_4 ), .A3(
        \SB2_2_25/i0[9] ), .ZN(n6629) );
  NAND4_X2 U13048 ( .A1(\SB2_3_27/Component_Function_3/NAND4_in[1] ), .A2(
        n1154), .A3(\SB2_3_27/Component_Function_3/NAND4_in[3] ), .A4(n6630), 
        .ZN(\SB2_3_27/buf_output[3] ) );
  NAND3_X2 U13049 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i0[6] ), .A3(
        \SB2_3_27/i1[9] ), .ZN(n6630) );
  INV_X2 U13050 ( .I(\SB1_3_16/buf_output[2] ), .ZN(\SB2_3_13/i1[9] ) );
  NAND4_X2 U13051 ( .A1(\SB1_3_16/Component_Function_2/NAND4_in[1] ), .A2(
        n3520), .A3(n7164), .A4(n7110), .ZN(\SB1_3_16/buf_output[2] ) );
  XOR2_X1 U13052 ( .A1(\MC_ARK_ARC_1_1/temp5[101] ), .A2(n1532), .Z(
        \MC_ARK_ARC_1_1/buf_output[101] ) );
  XOR2_X1 U13053 ( .A1(n2005), .A2(n6631), .Z(\MC_ARK_ARC_1_0/buf_output[28] )
         );
  XOR2_X1 U13054 ( .A1(\MC_ARK_ARC_1_0/temp1[28] ), .A2(
        \MC_ARK_ARC_1_0/temp2[28] ), .Z(n6631) );
  NAND3_X2 U13055 ( .A1(\SB2_3_8/i0[6] ), .A2(\SB2_3_8/i0_4 ), .A3(
        \SB2_3_8/i0[9] ), .ZN(n6882) );
  NAND4_X2 U13056 ( .A1(n1670), .A2(
        \SB1_3_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_12/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_3_12/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_12/buf_output[1] ) );
  XOR2_X1 U13057 ( .A1(n6633), .A2(n6632), .Z(\MC_ARK_ARC_1_4/temp5[68] ) );
  XOR2_X1 U13058 ( .A1(\RI5[4][62] ), .A2(\RI5[4][14] ), .Z(n6632) );
  XOR2_X1 U13059 ( .A1(\RI5[4][38] ), .A2(\RI5[4][68] ), .Z(n6633) );
  XOR2_X1 U13060 ( .A1(\RI5[2][123] ), .A2(\RI5[2][87] ), .Z(
        \MC_ARK_ARC_1_2/temp3[21] ) );
  NAND4_X2 U13061 ( .A1(\SB2_4_22/Component_Function_4/NAND4_in[3] ), .A2(
        n6797), .A3(n6739), .A4(\SB2_4_22/Component_Function_4/NAND4_in[1] ), 
        .ZN(\SB2_4_22/buf_output[4] ) );
  NAND4_X2 U13062 ( .A1(\SB1_3_2/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_3_2/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_3_2/Component_Function_0/NAND4_in[0] ), .A4(n6634), .ZN(
        \SB1_3_2/buf_output[0] ) );
  NAND3_X2 U13063 ( .A1(\SB2_2_8/i0[8] ), .A2(\SB2_2_8/i1_5 ), .A3(
        \SB2_2_8/i3[0] ), .ZN(n6635) );
  NAND3_X1 U13064 ( .A1(\SB1_2_10/i0[6] ), .A2(\SB1_2_10/i1[9] ), .A3(
        \SB1_2_10/i0_3 ), .ZN(\SB1_2_10/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U13065 ( .A1(\RI5[4][149] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[173] ), .Z(n6636) );
  XOR2_X1 U13066 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[50] ), .A2(\RI5[1][86] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[176] ) );
  NAND3_X1 U13067 ( .A1(\SB1_4_21/i0_4 ), .A2(\SB1_4_21/i0_0 ), .A3(
        \SB1_4_21/i1_5 ), .ZN(n6684) );
  NAND4_X2 U13068 ( .A1(n2579), .A2(\SB3_13/Component_Function_3/NAND4_in[0] ), 
        .A3(n736), .A4(n6638), .ZN(\SB3_13/buf_output[3] ) );
  NAND3_X2 U13069 ( .A1(\SB1_1_30/i0_0 ), .A2(\SB1_1_30/i0_4 ), .A3(
        \SB1_1_30/i0_3 ), .ZN(\SB1_1_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U13070 ( .A1(\SB1_2_26/i0[6] ), .A2(\SB1_2_26/i0_0 ), .A3(
        \SB1_2_26/i0[10] ), .ZN(n6639) );
  NAND4_X2 U13071 ( .A1(\SB2_4_21/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_4_21/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_4_21/Component_Function_4/NAND4_in[3] ), .A4(n6640), .ZN(
        \SB2_4_21/buf_output[4] ) );
  NAND3_X1 U13072 ( .A1(\SB2_4_21/i0[10] ), .A2(\SB2_4_21/i0_3 ), .A3(
        \SB2_4_21/i0[9] ), .ZN(n6640) );
  NAND4_X2 U13073 ( .A1(\SB1_3_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_6/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_3_6/Component_Function_1/NAND4_in[2] ), .A4(n6641), .ZN(
        \SB1_3_6/buf_output[1] ) );
  NAND3_X2 U13074 ( .A1(\SB1_3_6/i0_4 ), .A2(\SB1_3_6/i0[8] ), .A3(
        \SB1_3_6/i1_7 ), .ZN(n6641) );
  NAND4_X2 U13075 ( .A1(\SB3_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_11/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_5/NAND4_in[0] ), .A4(n6642), .ZN(
        \SB3_11/buf_output[5] ) );
  NAND3_X1 U13076 ( .A1(\SB3_11/i0_4 ), .A2(\SB3_11/i0[6] ), .A3(
        \MC_ARK_ARC_1_4/buf_output[120] ), .ZN(n6642) );
  XOR2_X1 U13077 ( .A1(n6643), .A2(n180), .Z(Ciphertext[105]) );
  XOR2_X1 U13078 ( .A1(n6644), .A2(\MC_ARK_ARC_1_1/temp1[86] ), .Z(n4070) );
  XOR2_X1 U13079 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[32] ), .A2(\RI5[1][56] ), 
        .Z(n6644) );
  NAND3_X2 U13080 ( .A1(\SB1_2_27/i0[9] ), .A2(\SB1_2_27/i0_4 ), .A3(
        \SB1_2_27/i0[6] ), .ZN(n911) );
  NAND4_X2 U13081 ( .A1(\SB2_2_15/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_2_15/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_15/Component_Function_5/NAND4_in[0] ), .A4(n6645), .ZN(
        \SB2_2_15/buf_output[5] ) );
  NAND3_X2 U13082 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i0_4 ), .A3(
        \SB2_2_15/i1[9] ), .ZN(n6645) );
  XOR2_X1 U13083 ( .A1(n6646), .A2(n3737), .Z(\MC_ARK_ARC_1_2/buf_output[163] ) );
  XOR2_X1 U13084 ( .A1(\MC_ARK_ARC_1_2/temp2[163] ), .A2(
        \MC_ARK_ARC_1_2/temp1[163] ), .Z(n6646) );
  NAND3_X2 U13085 ( .A1(\SB1_3_24/i0_3 ), .A2(\SB1_3_24/i0[8] ), .A3(
        \SB1_3_24/i0[9] ), .ZN(n6968) );
  NAND3_X2 U13086 ( .A1(\SB1_2_26/i0[8] ), .A2(\SB1_2_26/i3[0] ), .A3(
        \SB1_2_26/i1_5 ), .ZN(n1975) );
  NAND4_X2 U13087 ( .A1(\SB2_4_26/Component_Function_5/NAND4_in[0] ), .A2(
        n1744), .A3(\SB2_4_26/Component_Function_5/NAND4_in[1] ), .A4(n6647), 
        .ZN(\SB2_4_26/buf_output[5] ) );
  NAND3_X2 U13088 ( .A1(\SB2_4_26/i0[9] ), .A2(\SB2_4_26/i0[6] ), .A3(
        \SB2_4_26/i0_4 ), .ZN(n6647) );
  NAND3_X1 U13089 ( .A1(\SB1_4_31/i0_0 ), .A2(\RI1[4][5] ), .A3(
        \SB1_4_31/i0[7] ), .ZN(n4828) );
  NAND3_X1 U13090 ( .A1(\SB2_0_15/i0[6] ), .A2(\SB2_0_15/i0[8] ), .A3(
        \SB2_0_15/i0[7] ), .ZN(\SB2_0_15/Component_Function_0/NAND4_in[1] ) );
  NOR2_X2 U13091 ( .A1(n6649), .A2(n6648), .ZN(\SB2_0_15/i0[7] ) );
  XOR2_X1 U13092 ( .A1(n7158), .A2(\MC_ARK_ARC_1_0/temp1[156] ), .Z(
        \MC_ARK_ARC_1_0/temp5[156] ) );
  NAND3_X2 U13093 ( .A1(\SB2_0_22/i0_0 ), .A2(\SB2_0_22/i1_5 ), .A3(
        \RI3[0][58] ), .ZN(\SB2_0_22/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U13094 ( .A1(\SB2_2_8/i0[6] ), .A2(\SB2_2_8/i0_3 ), .A3(
        \SB2_2_8/i1[9] ), .ZN(n1650) );
  NAND3_X2 U13095 ( .A1(\SB2_0_17/i0[10] ), .A2(\SB2_0_17/i0[6] ), .A3(
        \SB2_0_17/i0_3 ), .ZN(n3884) );
  NAND4_X2 U13096 ( .A1(\SB2_1_13/Component_Function_3/NAND4_in[3] ), .A2(
        n6966), .A3(n2878), .A4(\SB2_1_13/Component_Function_3/NAND4_in[1] ), 
        .ZN(\SB2_1_13/buf_output[3] ) );
  NAND3_X2 U13097 ( .A1(\SB1_4_12/i0[8] ), .A2(\SB1_4_12/i0[9] ), .A3(
        \RI1[4][119] ), .ZN(n4205) );
  NAND4_X2 U13098 ( .A1(n4830), .A2(n4020), .A3(n2533), .A4(
        \SB1_3_20/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_20/buf_output[5] ) );
  NAND3_X2 U13099 ( .A1(\SB2_3_25/i0[8] ), .A2(\SB2_3_25/i3[0] ), .A3(
        \SB2_3_25/i1_5 ), .ZN(\SB2_3_25/Component_Function_3/NAND4_in[3] ) );
  INV_X2 U13100 ( .I(\SB1_2_10/buf_output[3] ), .ZN(\SB2_2_8/i0[8] ) );
  NAND4_X2 U13101 ( .A1(\SB1_2_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_10/Component_Function_3/NAND4_in[1] ), .A3(n6695), .A4(n1956), 
        .ZN(\SB1_2_10/buf_output[3] ) );
  XOR2_X1 U13102 ( .A1(\MC_ARK_ARC_1_3/temp6[132] ), .A2(n5175), .Z(
        \MC_ARK_ARC_1_3/buf_output[132] ) );
  XOR2_X1 U13103 ( .A1(\RI5[0][22] ), .A2(\RI5[0][28] ), .Z(
        \MC_ARK_ARC_1_0/temp1[28] ) );
  XOR2_X1 U13104 ( .A1(\RI5[0][117] ), .A2(\RI5[0][141] ), .Z(n3147) );
  XOR2_X1 U13105 ( .A1(n6650), .A2(\MC_ARK_ARC_1_2/temp4[32] ), .Z(n6808) );
  XOR2_X1 U13106 ( .A1(\RI5[2][32] ), .A2(\RI5[2][26] ), .Z(n6650) );
  NAND4_X2 U13107 ( .A1(\SB1_2_6/Component_Function_5/NAND4_in[3] ), .A2(n4264), .A3(n6663), .A4(\SB1_2_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_6/buf_output[5] ) );
  NAND4_X2 U13108 ( .A1(n6886), .A2(
        \SB2_2_12/Component_Function_3/NAND4_in[2] ), .A3(n5330), .A4(
        \SB2_2_12/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_12/buf_output[3] ) );
  NAND3_X2 U13109 ( .A1(\SB2_3_20/i0_0 ), .A2(\SB2_3_20/i0_3 ), .A3(
        \RI3[3][70] ), .ZN(n6810) );
  XOR2_X1 U13110 ( .A1(\RI5[2][170] ), .A2(\RI5[2][134] ), .Z(
        \MC_ARK_ARC_1_2/temp3[68] ) );
  NAND4_X2 U13111 ( .A1(\SB1_2_29/Component_Function_5/NAND4_in[1] ), .A2(
        n5035), .A3(n6892), .A4(\SB1_2_29/Component_Function_5/NAND4_in[0] ), 
        .ZN(\SB1_2_29/buf_output[5] ) );
  XOR2_X1 U13112 ( .A1(n1480), .A2(n4979), .Z(n3975) );
  NOR2_X2 U13113 ( .A1(n1319), .A2(n1317), .ZN(n6651) );
  AOI21_X2 U13114 ( .A1(\SB2_1_14/i3[0] ), .A2(\SB2_1_14/i0_0 ), .B(n6653), 
        .ZN(n6652) );
  NAND3_X2 U13115 ( .A1(\SB2_4_14/i0_3 ), .A2(\SB2_4_14/i0[10] ), .A3(
        \SB2_4_14/i0[6] ), .ZN(n6654) );
  XOR2_X1 U13116 ( .A1(n6657), .A2(n6656), .Z(n4479) );
  XOR2_X1 U13117 ( .A1(\RI5[0][140] ), .A2(n190), .Z(n6656) );
  XOR2_X1 U13118 ( .A1(n4687), .A2(\MC_ARK_ARC_1_2/temp5[81] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[81] ) );
  XOR2_X1 U13119 ( .A1(n6658), .A2(\MC_ARK_ARC_1_3/temp6[57] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[57] ) );
  NAND3_X2 U13120 ( .A1(\SB2_3_29/i0_4 ), .A2(n6552), .A3(
        \SB1_3_2/buf_output[0] ), .ZN(n2407) );
  NAND3_X2 U13121 ( .A1(\SB2_4_7/i0_3 ), .A2(\SB2_4_7/i1[9] ), .A3(
        \RI3[4][148] ), .ZN(n4845) );
  XOR2_X1 U13122 ( .A1(\MC_ARK_ARC_1_3/temp6[149] ), .A2(
        \MC_ARK_ARC_1_3/temp5[149] ), .Z(\MC_ARK_ARC_1_3/buf_output[149] ) );
  NAND3_X2 U13123 ( .A1(\SB1_4_7/i0_3 ), .A2(\SB1_4_7/i0_4 ), .A3(
        \SB1_4_7/i1[9] ), .ZN(n6659) );
  NAND4_X2 U13124 ( .A1(\SB2_3_28/Component_Function_2/NAND4_in[0] ), .A2(
        n7558), .A3(\SB2_3_28/Component_Function_2/NAND4_in[3] ), .A4(n6660), 
        .ZN(\SB2_3_28/buf_output[2] ) );
  NAND3_X2 U13125 ( .A1(\SB2_3_28/i0_3 ), .A2(\SB2_3_28/i0[10] ), .A3(
        \SB2_3_28/i0[6] ), .ZN(n6660) );
  XOR2_X1 U13126 ( .A1(n6661), .A2(\MC_ARK_ARC_1_0/temp4[125] ), .Z(n3123) );
  XOR2_X1 U13127 ( .A1(\RI5[0][191] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[35] ), 
        .Z(n6661) );
  XOR2_X1 U13128 ( .A1(\MC_ARK_ARC_1_3/temp1[51] ), .A2(n6662), .Z(
        \MC_ARK_ARC_1_3/temp5[51] ) );
  XOR2_X1 U13129 ( .A1(\RI5[3][189] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[21] ), 
        .Z(n6662) );
  NAND3_X2 U13130 ( .A1(\SB1_2_6/i0_0 ), .A2(\SB1_2_6/i0[10] ), .A3(
        \SB1_2_6/i0[6] ), .ZN(n6663) );
  NAND3_X2 U13131 ( .A1(\SB2_2_2/i0_3 ), .A2(n6267), .A3(\SB2_2_2/i0[6] ), 
        .ZN(\SB2_2_2/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U13132 ( .A1(n690), .A2(\SB1_4_25/Component_Function_4/NAND4_in[2] ), .A3(\SB1_4_25/Component_Function_4/NAND4_in[1] ), .A4(n6665), .ZN(
        \SB1_4_25/buf_output[4] ) );
  NAND3_X1 U13133 ( .A1(\SB2_0_8/i0_0 ), .A2(\SB2_0_8/i3[0] ), .A3(
        \SB2_0_8/i1_7 ), .ZN(\SB2_0_8/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U13134 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[65] ), .A2(\RI5[2][101] ), 
        .Z(n6666) );
  XOR2_X1 U13135 ( .A1(n6668), .A2(n6667), .Z(\MC_ARK_ARC_1_4/temp6[11] ) );
  XOR2_X1 U13136 ( .A1(\RI5[4][113] ), .A2(n438), .Z(n6667) );
  XOR2_X1 U13137 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[77] ), .A2(\RI5[4][47] ), 
        .Z(n6668) );
  XOR2_X1 U13138 ( .A1(\RI5[1][176] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[182] ), .Z(n6669) );
  NAND4_X2 U13139 ( .A1(\SB2_4_24/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_24/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_4_24/Component_Function_0/NAND4_in[0] ), .A4(n6671), .ZN(
        \SB2_4_24/buf_output[0] ) );
  NAND3_X1 U13140 ( .A1(\SB2_4_24/i0_3 ), .A2(\SB2_4_24/i0[10] ), .A3(
        \SB2_4_24/i0_4 ), .ZN(n6671) );
  NAND3_X2 U13141 ( .A1(\SB1_2_8/i0[10] ), .A2(\SB1_2_8/i0_0 ), .A3(
        \SB1_2_8/i0[6] ), .ZN(\SB1_2_8/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U13142 ( .A1(\RI5[3][58] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[184] ), 
        .Z(n7079) );
  NAND4_X2 U13143 ( .A1(\SB2_3_23/Component_Function_4/NAND4_in[3] ), .A2(
        n2996), .A3(\SB2_3_23/Component_Function_4/NAND4_in[0] ), .A4(n7232), 
        .ZN(\SB2_3_23/buf_output[4] ) );
  XOR2_X1 U13144 ( .A1(n6674), .A2(\MC_ARK_ARC_1_2/temp6[133] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[133] ) );
  XOR2_X1 U13145 ( .A1(\MC_ARK_ARC_1_2/temp1[133] ), .A2(n6929), .Z(n6674) );
  XOR2_X1 U13146 ( .A1(\MC_ARK_ARC_1_2/temp6[173] ), .A2(n6675), .Z(
        \MC_ARK_ARC_1_2/buf_output[173] ) );
  XOR2_X1 U13147 ( .A1(n7295), .A2(\MC_ARK_ARC_1_2/temp1[173] ), .Z(n6675) );
  NAND3_X1 U13148 ( .A1(\SB2_1_11/i0[10] ), .A2(\SB2_1_11/i0_3 ), .A3(
        \SB2_1_11/i0_4 ), .ZN(\SB2_1_11/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U13149 ( .A1(n6870), .A2(n6676), .Z(n7086) );
  XOR2_X1 U13150 ( .A1(\RI5[4][62] ), .A2(\RI5[4][26] ), .Z(n6676) );
  NAND4_X2 U13151 ( .A1(\SB2_1_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_13/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_1_13/Component_Function_4/NAND4_in[1] ), .A4(n6677), .ZN(
        \SB2_1_13/buf_output[4] ) );
  NAND3_X2 U13152 ( .A1(\SB1_4_27/i1[9] ), .A2(\SB1_4_27/i0[10] ), .A3(
        \SB1_4_27/i1_7 ), .ZN(\SB1_4_27/Component_Function_3/NAND4_in[2] ) );
  INV_X2 U13153 ( .I(\SB1_2_19/buf_output[3] ), .ZN(\SB2_2_17/i0[8] ) );
  NAND4_X2 U13154 ( .A1(\SB1_2_19/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_19/Component_Function_3/NAND4_in[0] ), .A3(n3852), .A4(n2086), 
        .ZN(\SB1_2_19/buf_output[3] ) );
  NAND3_X2 U13155 ( .A1(\SB1_3_12/i0[10] ), .A2(\SB1_3_12/i1_7 ), .A3(
        \SB1_3_12/i1[9] ), .ZN(n6678) );
  NAND4_X2 U13156 ( .A1(\SB1_3_30/Component_Function_0/NAND4_in[1] ), .A2(
        n7549), .A3(\SB1_3_30/Component_Function_0/NAND4_in[3] ), .A4(n6679), 
        .ZN(\SB1_3_30/buf_output[0] ) );
  NAND2_X2 U13157 ( .A1(\SB1_3_30/i0[10] ), .A2(\SB1_3_30/i0[9] ), .ZN(n6679)
         );
  XOR2_X1 U13158 ( .A1(n6680), .A2(\MC_ARK_ARC_1_3/temp4[45] ), .Z(n6972) );
  XOR2_X1 U13159 ( .A1(\RI5[3][111] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[147] ), .Z(n6680) );
  XOR2_X1 U13160 ( .A1(\RI5[1][140] ), .A2(\RI5[1][134] ), .Z(
        \MC_ARK_ARC_1_1/temp1[140] ) );
  XOR2_X1 U13161 ( .A1(n7579), .A2(n6681), .Z(\MC_ARK_ARC_1_2/buf_output[115] ) );
  XOR2_X1 U13162 ( .A1(n4872), .A2(\MC_ARK_ARC_1_2/temp4[115] ), .Z(n6681) );
  NAND3_X2 U13163 ( .A1(\SB1_1_11/i0[9] ), .A2(\SB1_1_11/i0_4 ), .A3(
        \SB1_1_11/i0[6] ), .ZN(\SB1_1_11/Component_Function_5/NAND4_in[3] ) );
  INV_X2 U13164 ( .I(\SB1_3_11/buf_output[2] ), .ZN(\SB2_3_8/i1[9] ) );
  NAND3_X2 U13165 ( .A1(\SB2_4_6/i0_4 ), .A2(\SB2_4_6/i0[6] ), .A3(
        \SB2_4_6/i0[9] ), .ZN(n7120) );
  NAND4_X2 U13166 ( .A1(\SB2_1_10/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_10/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_10/Component_Function_2/NAND4_in[2] ), .A4(n6683), .ZN(
        \SB2_1_10/buf_output[2] ) );
  NAND3_X2 U13167 ( .A1(\SB2_3_15/i0_4 ), .A2(\SB2_3_15/i0_3 ), .A3(
        \SB2_3_15/i0_0 ), .ZN(n6685) );
  NAND4_X2 U13168 ( .A1(\SB2_1_11/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_1_11/Component_Function_2/NAND4_in[0] ), .A3(n6951), .A4(
        \SB2_1_11/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_1_11/buf_output[2] ) );
  XOR2_X1 U13169 ( .A1(\MC_ARK_ARC_1_2/temp5[141] ), .A2(
        \MC_ARK_ARC_1_2/temp6[141] ), .Z(\MC_ARK_ARC_1_2/buf_output[141] ) );
  NAND4_X2 U13170 ( .A1(n857), .A2(\SB1_3_29/Component_Function_5/NAND4_in[2] ), .A3(n7546), .A4(\SB1_3_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_29/buf_output[5] ) );
  XOR2_X1 U13171 ( .A1(\SB2_1_22/buf_output[2] ), .A2(\RI5[1][140] ), .Z(n7024) );
  NAND4_X2 U13172 ( .A1(\SB1_1_11/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_11/Component_Function_5/NAND4_in[3] ), .A3(n4427), .A4(
        \SB1_1_11/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_11/buf_output[5] ) );
  XOR2_X1 U13173 ( .A1(n6687), .A2(\MC_ARK_ARC_1_3/temp2[56] ), .Z(n626) );
  XOR2_X1 U13174 ( .A1(\RI5[3][122] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[158] ), .Z(n6687) );
  XOR2_X1 U13175 ( .A1(\MC_ARK_ARC_1_3/temp5[86] ), .A2(n6688), .Z(
        \MC_ARK_ARC_1_3/buf_output[86] ) );
  XOR2_X1 U13176 ( .A1(\MC_ARK_ARC_1_3/temp4[86] ), .A2(
        \MC_ARK_ARC_1_3/temp3[86] ), .Z(n6688) );
  XOR2_X1 U13177 ( .A1(n6689), .A2(\MC_ARK_ARC_1_4/temp6[166] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[166] ) );
  XOR2_X1 U13178 ( .A1(\MC_ARK_ARC_1_4/temp1[166] ), .A2(
        \MC_ARK_ARC_1_4/temp2[166] ), .Z(n6689) );
  XOR2_X1 U13179 ( .A1(n5385), .A2(n6690), .Z(\MC_ARK_ARC_1_1/buf_output[137] ) );
  XOR2_X1 U13180 ( .A1(\MC_ARK_ARC_1_1/temp3[137] ), .A2(
        \MC_ARK_ARC_1_1/temp4[137] ), .Z(n6690) );
  XOR2_X1 U13181 ( .A1(\MC_ARK_ARC_1_4/temp1[2] ), .A2(n6691), .Z(n1930) );
  XOR2_X1 U13182 ( .A1(\RI5[4][164] ), .A2(\RI5[4][140] ), .Z(n6691) );
  NAND3_X2 U13183 ( .A1(\SB3_31/i0[10] ), .A2(\SB3_31/i1[9] ), .A3(
        \SB3_31/i1_5 ), .ZN(n6692) );
  NAND3_X2 U13184 ( .A1(\SB3_30/i1_5 ), .A2(\SB3_30/i0[8] ), .A3(
        \SB3_30/i3[0] ), .ZN(n6970) );
  NAND4_X2 U13185 ( .A1(n2012), .A2(
        \SB1_2_15/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_2_15/Component_Function_3/NAND4_in[0] ), .A4(n6693), .ZN(
        \SB1_2_15/buf_output[3] ) );
  INV_X2 U13186 ( .I(\SB1_3_30/buf_output[3] ), .ZN(\SB2_3_28/i0[8] ) );
  NAND4_X2 U13187 ( .A1(\SB1_3_30/Component_Function_3/NAND4_in[1] ), .A2(
        n5109), .A3(\SB1_3_30/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_3_30/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_30/buf_output[3] ) );
  NAND3_X1 U13188 ( .A1(\SB4_10/i0_0 ), .A2(\SB4_10/i0_4 ), .A3(\SB4_10/i0_3 ), 
        .ZN(\SB4_10/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U13189 ( .A1(\SB1_4_16/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_4_16/Component_Function_2/NAND4_in[0] ), .A3(n3451), .A4(n6694), 
        .ZN(\SB1_4_16/buf_output[2] ) );
  NAND3_X2 U13190 ( .A1(\SB1_4_16/i0_3 ), .A2(\SB1_4_16/i0[8] ), .A3(
        \SB1_4_16/i0[9] ), .ZN(n6694) );
  NAND3_X2 U13191 ( .A1(\SB1_2_10/i0[10] ), .A2(\SB1_2_10/i1[9] ), .A3(
        \SB1_2_10/i1_7 ), .ZN(n6695) );
  NAND3_X2 U13192 ( .A1(\SB1_1_24/i1_5 ), .A2(\SB1_1_24/i1[9] ), .A3(
        \SB1_1_24/i0[10] ), .ZN(n6696) );
  XOR2_X1 U13193 ( .A1(n626), .A2(n6698), .Z(\MC_ARK_ARC_1_3/buf_output[56] )
         );
  XOR2_X1 U13194 ( .A1(n6783), .A2(n6784), .Z(n6698) );
  XOR2_X1 U13195 ( .A1(\RI5[2][12] ), .A2(\RI5[2][6] ), .Z(
        \MC_ARK_ARC_1_2/temp1[12] ) );
  XOR2_X1 U13196 ( .A1(\MC_ARK_ARC_1_3/temp2[148] ), .A2(n6699), .Z(
        \MC_ARK_ARC_1_3/temp5[148] ) );
  XOR2_X1 U13197 ( .A1(\SB2_3_9/buf_output[4] ), .A2(\RI5[3][148] ), .Z(n6699)
         );
  AND2_X1 U13198 ( .A1(\MC_ARK_ARC_1_3/buf_output[24] ), .A2(
        \MC_ARK_ARC_1_3/buf_output[28] ), .Z(n6701) );
  NAND3_X2 U13199 ( .A1(\SB2_1_15/i0[10] ), .A2(\SB2_1_15/i0_0 ), .A3(
        \SB2_1_15/i0[6] ), .ZN(n6702) );
  XOR2_X1 U13200 ( .A1(\MC_ARK_ARC_1_2/temp1[13] ), .A2(
        \MC_ARK_ARC_1_2/temp2[13] ), .Z(n6910) );
  NAND4_X2 U13201 ( .A1(\SB1_1_17/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_17/Component_Function_3/NAND4_in[1] ), .A3(n1723), .A4(n6703), 
        .ZN(\SB1_1_17/buf_output[3] ) );
  XOR2_X1 U13202 ( .A1(n4017), .A2(n4800), .Z(\MC_ARK_ARC_1_2/buf_output[113] ) );
  XOR2_X1 U13203 ( .A1(n4259), .A2(\MC_ARK_ARC_1_2/temp4[113] ), .Z(n4017) );
  XOR2_X1 U13204 ( .A1(n1599), .A2(n6704), .Z(\MC_ARK_ARC_1_4/buf_output[7] )
         );
  XOR2_X1 U13205 ( .A1(\MC_ARK_ARC_1_4/temp2[7] ), .A2(
        \MC_ARK_ARC_1_4/temp1[7] ), .Z(n6704) );
  XOR2_X1 U13206 ( .A1(\MC_ARK_ARC_1_4/temp5[40] ), .A2(n6705), .Z(
        \MC_ARK_ARC_1_4/buf_output[40] ) );
  XOR2_X1 U13207 ( .A1(n3904), .A2(\MC_ARK_ARC_1_4/temp4[40] ), .Z(n6705) );
  NAND3_X2 U13208 ( .A1(\SB3_18/i0[6] ), .A2(\SB3_18/i1[9] ), .A3(
        \SB3_18/i0_3 ), .ZN(n6706) );
  NAND3_X1 U13209 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i0[6] ), .A3(
        \SB4_20/i0[10] ), .ZN(n6707) );
  NAND3_X2 U13210 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i1[9] ), .A3(
        \SB3_30/i0[6] ), .ZN(\SB3_30/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U13211 ( .A1(\RI5[0][93] ), .A2(\RI5[0][99] ), .Z(
        \MC_ARK_ARC_1_0/temp1[99] ) );
  NAND3_X2 U13212 ( .A1(\SB1_4_25/i0[6] ), .A2(\SB1_4_25/i0[9] ), .A3(
        \SB1_4_25/i0_4 ), .ZN(\SB1_4_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U13213 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i1[9] ), .A3(
        \SB2_1_4/i0_4 ), .ZN(\SB2_1_4/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U13214 ( .A1(n7094), .A2(
        \SB1_3_28/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_3_28/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_3_28/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_28/buf_output[5] ) );
  NAND4_X2 U13215 ( .A1(\SB2_4_19/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_4_19/Component_Function_5/NAND4_in[1] ), .A3(n3678), .A4(
        \SB2_4_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_4_19/buf_output[5] ) );
  NAND4_X2 U13216 ( .A1(\SB2_3_28/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_28/Component_Function_0/NAND4_in[3] ), .A3(n6711), .A4(
        \SB2_3_28/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_28/buf_output[0] ) );
  XOR2_X1 U13217 ( .A1(\MC_ARK_ARC_1_4/temp4[80] ), .A2(n6708), .Z(n6849) );
  XOR2_X1 U13218 ( .A1(\RI5[4][182] ), .A2(\RI5[4][146] ), .Z(n6708) );
  XOR2_X1 U13219 ( .A1(\MC_ARK_ARC_1_3/temp6[174] ), .A2(n3195), .Z(
        \MC_ARK_ARC_1_3/buf_output[174] ) );
  NAND3_X1 U13220 ( .A1(\SB4_20/i1_5 ), .A2(\SB4_20/i0[10] ), .A3(
        \SB4_20/i1[9] ), .ZN(\SB4_20/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U13221 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i0[9] ), .ZN(n2412) );
  XOR2_X1 U13222 ( .A1(n1449), .A2(n1448), .Z(\MC_ARK_ARC_1_2/temp6[143] ) );
  NAND3_X2 U13223 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i0[9] ), .A3(
        \SB1_3_8/i0[10] ), .ZN(n3475) );
  NAND3_X2 U13224 ( .A1(\SB1_2_27/i0[9] ), .A2(\SB1_2_27/i0[8] ), .A3(
        \SB1_2_27/i0_0 ), .ZN(n6710) );
  NAND3_X1 U13225 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i0[9] ), .A3(
        \SB4_20/i0[8] ), .ZN(n4863) );
  XOR2_X1 U13226 ( .A1(\MC_ARK_ARC_1_4/temp1[66] ), .A2(
        \MC_ARK_ARC_1_4/temp2[66] ), .Z(n3368) );
  NAND3_X2 U13227 ( .A1(\SB2_2_2/i0_4 ), .A2(\SB2_2_2/i0[6] ), .A3(
        \SB2_2_2/i0[9] ), .ZN(n6712) );
  NAND2_X2 U13228 ( .A1(\SB1_2_15/i0_0 ), .A2(\SB1_2_15/i3[0] ), .ZN(
        \SB1_2_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U13229 ( .A1(\SB2_3_28/i0_3 ), .A2(\SB1_3_29/buf_output[4] ), .A3(
        \SB2_3_28/i0[10] ), .ZN(n6711) );
  NAND4_X2 U13230 ( .A1(\SB2_2_2/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_2/Component_Function_0/NAND4_in[3] ), .A3(n4387), .A4(
        \SB2_2_2/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_2/buf_output[0] ) );
  XOR2_X1 U13231 ( .A1(\RI5[3][48] ), .A2(\RI5[3][84] ), .Z(n1205) );
  NAND3_X2 U13232 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i0[9] ), .A3(
        \SB4_28/i0[8] ), .ZN(\SB4_28/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U13233 ( .A1(\MC_ARK_ARC_1_1/temp2[98] ), .A2(n4344), .Z(n4150) );
  NAND4_X2 U13234 ( .A1(n1143), .A2(n6712), .A3(
        \SB2_2_2/Component_Function_5/NAND4_in[0] ), .A4(n4527), .ZN(
        \SB2_2_2/buf_output[5] ) );
  XOR2_X1 U13235 ( .A1(n2343), .A2(n6713), .Z(\MC_ARK_ARC_1_0/buf_output[152] ) );
  XOR2_X1 U13236 ( .A1(n5056), .A2(n5055), .Z(n6713) );
  NAND4_X2 U13237 ( .A1(\SB4_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_28/Component_Function_1/NAND4_in[3] ), .A3(n2379), .A4(n6714), 
        .ZN(n3630) );
  NAND2_X2 U13238 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i1[9] ), .ZN(n6714) );
  XOR2_X1 U13239 ( .A1(\MC_ARK_ARC_1_2/temp5[118] ), .A2(n6715), .Z(
        \MC_ARK_ARC_1_2/buf_output[118] ) );
  XOR2_X1 U13240 ( .A1(\MC_ARK_ARC_1_2/temp3[118] ), .A2(
        \MC_ARK_ARC_1_2/temp4[118] ), .Z(n6715) );
  NAND3_X2 U13241 ( .A1(\SB2_2_2/i0_0 ), .A2(\SB2_2_2/i1_5 ), .A3(
        \SB2_2_2/i0_4 ), .ZN(n6766) );
  NAND3_X2 U13242 ( .A1(\SB2_4_10/i0[10] ), .A2(\SB2_4_10/i0[6] ), .A3(
        \SB2_4_10/i0_3 ), .ZN(n6787) );
  XOR2_X1 U13243 ( .A1(\RI5[2][128] ), .A2(\RI5[2][2] ), .Z(n7355) );
  NAND3_X2 U13244 ( .A1(\SB2_1_23/i0[9] ), .A2(\SB2_1_23/i0_4 ), .A3(
        \SB2_1_23/i0[6] ), .ZN(n6717) );
  NAND3_X1 U13245 ( .A1(\SB1_3_22/i0_4 ), .A2(\SB1_3_22/i1[9] ), .A3(
        \SB1_3_22/i1_5 ), .ZN(n2674) );
  NAND3_X1 U13246 ( .A1(\SB3_12/i0[10] ), .A2(\SB3_12/i0[6] ), .A3(
        \RI1[5][119] ), .ZN(n6996) );
  NAND4_X2 U13247 ( .A1(n974), .A2(\SB2_0_0/Component_Function_2/NAND4_in[2] ), 
        .A3(\SB2_0_0/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_0_0/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_0/buf_output[2] ) );
  NAND4_X2 U13248 ( .A1(\SB2_1_8/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_8/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_8/Component_Function_1/NAND4_in[2] ), .A4(n6719), .ZN(
        \SB2_1_8/buf_output[1] ) );
  NAND3_X2 U13249 ( .A1(\SB2_1_8/i0_4 ), .A2(\SB2_1_8/i1_7 ), .A3(
        \SB2_1_8/i0[8] ), .ZN(n6719) );
  NOR2_X1 U13250 ( .A1(\MC_ARK_ARC_1_1/buf_output[127] ), .A2(
        \MC_ARK_ARC_1_1/buf_output[129] ), .ZN(n6909) );
  NAND3_X1 U13251 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i0[10] ), .A3(
        \SB2_3_1/i0_4 ), .ZN(\SB2_3_1/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U13252 ( .A1(\SB2_3_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_1/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_3_1/Component_Function_3/NAND4_in[3] ), .A4(n6720), .ZN(
        \SB2_3_1/buf_output[3] ) );
  NAND3_X2 U13253 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i0_0 ), .A3(
        \SB2_3_1/i0_4 ), .ZN(n6720) );
  NAND3_X2 U13254 ( .A1(\SB1_4_6/i1_5 ), .A2(\SB1_4_6/i0_0 ), .A3(
        \SB1_4_6/i0_4 ), .ZN(n6721) );
  NAND3_X2 U13255 ( .A1(\SB2_3_0/i0_4 ), .A2(\SB2_3_0/i0[6] ), .A3(
        \SB2_3_0/i0[9] ), .ZN(\SB2_3_0/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U13256 ( .A1(n4918), .A2(n1246), .A3(
        \SB2_4_23/Component_Function_4/NAND4_in[3] ), .A4(n6723), .ZN(
        \SB2_4_23/buf_output[4] ) );
  NAND3_X1 U13257 ( .A1(\SB2_4_23/i0_0 ), .A2(\SB2_4_23/i3[0] ), .A3(
        \SB2_4_23/i1_7 ), .ZN(n6723) );
  AND2_X1 U13258 ( .A1(n3233), .A2(\SB1_4_21/Component_Function_4/NAND4_in[1] ), .Z(n6724) );
  XOR2_X1 U13259 ( .A1(\RI5[3][33] ), .A2(\RI5[3][9] ), .Z(n6725) );
  NAND3_X1 U13260 ( .A1(\SB2_3_5/i0[7] ), .A2(\SB2_3_5/i0[6] ), .A3(
        \SB2_3_5/i0[8] ), .ZN(\SB2_3_5/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U13261 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[145] ), .A2(\RI5[1][121] ), .Z(\MC_ARK_ARC_1_1/temp2[175] ) );
  NAND4_X2 U13262 ( .A1(\SB1_4_9/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_4_9/Component_Function_3/NAND4_in[1] ), .A3(n1228), .A4(n6726), 
        .ZN(\SB1_4_9/buf_output[3] ) );
  NAND3_X2 U13263 ( .A1(\SB1_2_1/i0_3 ), .A2(\SB1_2_1/i0_4 ), .A3(
        \SB1_2_1/i1[9] ), .ZN(n6727) );
  XOR2_X1 U13264 ( .A1(n6728), .A2(\MC_ARK_ARC_1_4/temp6[117] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[117] ) );
  XOR2_X1 U13265 ( .A1(n2225), .A2(\MC_ARK_ARC_1_4/temp1[117] ), .Z(n6728) );
  NAND3_X2 U13266 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0[10] ), .A3(
        \SB2_3_0/i0_4 ), .ZN(\SB2_3_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U13267 ( .A1(\SB2_0_0/i0[10] ), .A2(\SB2_0_0/i0[6] ), .A3(
        \SB2_0_0/i0_3 ), .ZN(n974) );
  XOR2_X1 U13268 ( .A1(\RI5[0][161] ), .A2(\RI5[0][155] ), .Z(
        \MC_ARK_ARC_1_0/temp1[161] ) );
  NAND3_X2 U13269 ( .A1(\SB2_3_9/i0_0 ), .A2(\SB2_3_9/i0[10] ), .A3(
        \SB2_3_9/i0[6] ), .ZN(n6730) );
  XOR2_X1 U13270 ( .A1(n6980), .A2(n1647), .Z(\MC_ARK_ARC_1_0/buf_output[191] ) );
  NAND4_X2 U13271 ( .A1(\SB1_3_6/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_6/Component_Function_3/NAND4_in[0] ), .A3(n3053), .A4(n2163), 
        .ZN(\SB1_3_6/buf_output[3] ) );
  XOR2_X1 U13272 ( .A1(\MC_ARK_ARC_1_3/temp2[113] ), .A2(
        \MC_ARK_ARC_1_3/temp1[113] ), .Z(n6731) );
  XOR2_X1 U13273 ( .A1(\RI5[0][191] ), .A2(\RI5[0][167] ), .Z(
        \MC_ARK_ARC_1_0/temp2[29] ) );
  XOR2_X1 U13274 ( .A1(\RI5[1][129] ), .A2(\RI5[1][165] ), .Z(
        \MC_ARK_ARC_1_1/temp3[63] ) );
  NAND3_X2 U13275 ( .A1(\SB1_4_13/i0_3 ), .A2(\SB1_4_13/i0[9] ), .A3(
        \SB1_4_13/i0[8] ), .ZN(n7353) );
  NAND4_X2 U13276 ( .A1(\SB1_0_4/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_4/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_0_4/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_4/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][187] ) );
  NAND3_X1 U13277 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0_4 ), .A3(n6290), 
        .ZN(\SB1_0_18/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U13278 ( .A1(\SB1_3_31/Component_Function_1/NAND4_in[0] ), .A2(
        n1577), .A3(\SB1_3_31/Component_Function_1/NAND4_in[3] ), .A4(n4762), 
        .ZN(\SB1_3_31/buf_output[1] ) );
  INV_X2 U13279 ( .I(\RI3[0][81] ), .ZN(\SB2_0_18/i0[8] ) );
  NAND3_X2 U13280 ( .A1(n2946), .A2(n6895), .A3(
        \SB1_0_20/Component_Function_3/NAND4_in[1] ), .ZN(\RI3[0][81] ) );
  NAND3_X1 U13281 ( .A1(\SB1_2_30/i0[6] ), .A2(\SB1_2_30/i0[7] ), .A3(
        \SB1_2_30/i0[8] ), .ZN(\SB1_2_30/Component_Function_0/NAND4_in[1] ) );
  INV_X2 U13282 ( .I(\SB1_1_13/buf_output[3] ), .ZN(\SB2_1_11/i0[8] ) );
  NAND4_X2 U13283 ( .A1(\SB1_1_13/Component_Function_3/NAND4_in[0] ), .A2(
        n7456), .A3(\SB1_1_13/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_1_13/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_13/buf_output[3] ) );
  NAND4_X2 U13284 ( .A1(\SB1_2_5/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_5/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_2_5/Component_Function_1/NAND4_in[3] ), .A4(n6732), .ZN(
        \SB1_2_5/buf_output[1] ) );
  XOR2_X1 U13285 ( .A1(\MC_ARK_ARC_1_3/temp1[184] ), .A2(n6733), .Z(n6781) );
  XOR2_X1 U13286 ( .A1(\RI5[3][154] ), .A2(\RI5[3][130] ), .Z(n6733) );
  XOR2_X1 U13287 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[122] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[98] ), .Z(n2957) );
  XOR2_X1 U13288 ( .A1(n2980), .A2(n6734), .Z(\MC_ARK_ARC_1_4/buf_output[110] ) );
  XOR2_X1 U13289 ( .A1(\MC_ARK_ARC_1_4/temp3[110] ), .A2(
        \MC_ARK_ARC_1_4/temp4[110] ), .Z(n6734) );
  NAND3_X2 U13290 ( .A1(\SB2_4_18/i0[10] ), .A2(\SB2_4_18/i0_0 ), .A3(
        \SB2_4_18/i0[6] ), .ZN(n5094) );
  XOR2_X1 U13291 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[145] ), .A2(\RI5[1][169] ), .Z(n6735) );
  XOR2_X1 U13292 ( .A1(n4140), .A2(\MC_ARK_ARC_1_1/temp4[73] ), .Z(n3878) );
  NAND4_X2 U13293 ( .A1(\SB2_1_13/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_13/Component_Function_2/NAND4_in[0] ), .A3(n7267), .A4(n3660), 
        .ZN(\SB2_1_13/buf_output[2] ) );
  NAND3_X2 U13294 ( .A1(\SB1_3_9/i0[6] ), .A2(n3979), .A3(\SB1_3_9/i0_4 ), 
        .ZN(n6736) );
  BUF_X2 U13295 ( .I(\SB1_2_7/buf_output[5] ), .Z(n6737) );
  NAND3_X2 U13296 ( .A1(\SB2_0_0/i0_3 ), .A2(\SB2_0_0/i0[6] ), .A3(
        \SB2_0_0/i1[9] ), .ZN(\SB2_0_0/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U13297 ( .A1(\SB2_1_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_11/Component_Function_5/NAND4_in[1] ), .A3(n7469), .A4(
        \SB2_1_11/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_11/buf_output[5] ) );
  XOR2_X1 U13298 ( .A1(\RI5[2][42] ), .A2(\RI5[2][48] ), .Z(n6738) );
  XOR2_X1 U13299 ( .A1(\RI5[3][3] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[159] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[93] ) );
  INV_X2 U13300 ( .I(\SB3_14/buf_output[3] ), .ZN(\SB4_12/i0[8] ) );
  NAND4_X2 U13301 ( .A1(\SB3_14/Component_Function_3/NAND4_in[2] ), .A2(n4050), 
        .A3(\SB3_14/Component_Function_3/NAND4_in[1] ), .A4(n7357), .ZN(
        \SB3_14/buf_output[3] ) );
  XOR2_X1 U13302 ( .A1(\MC_ARK_ARC_1_3/temp3[76] ), .A2(
        \MC_ARK_ARC_1_3/temp4[76] ), .Z(\MC_ARK_ARC_1_3/temp6[76] ) );
  NAND3_X2 U13303 ( .A1(\SB2_4_22/i0_0 ), .A2(\SB2_4_22/i0[8] ), .A3(
        \SB2_4_22/i0[9] ), .ZN(n6739) );
  NAND3_X2 U13304 ( .A1(\SB2_4_24/i0_3 ), .A2(\SB2_4_24/i0[9] ), .A3(
        \SB2_4_24/i0[8] ), .ZN(n4167) );
  NAND4_X2 U13305 ( .A1(\SB1_1_27/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_1_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_27/Component_Function_1/NAND4_in[0] ), .A4(n6740), .ZN(
        \SB1_1_27/buf_output[1] ) );
  NAND3_X2 U13306 ( .A1(\SB3_6/i0_4 ), .A2(\SB3_6/i1[9] ), .A3(\SB3_6/i0_3 ), 
        .ZN(\SB3_6/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U13307 ( .A1(n3551), .A2(
        \SB1_4_19/Component_Function_2/NAND4_in[1] ), .A3(n7140), .A4(n6741), 
        .ZN(\SB1_4_19/buf_output[2] ) );
  NAND3_X2 U13308 ( .A1(\SB1_4_19/i0_0 ), .A2(\SB1_4_19/i0_4 ), .A3(
        \SB1_4_19/i1_5 ), .ZN(n6741) );
  NAND3_X1 U13309 ( .A1(\SB1_0_4/i0_3 ), .A2(\SB1_0_4/i1[9] ), .A3(
        \SB1_0_4/i0[6] ), .ZN(\SB1_0_4/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U13310 ( .A1(n6742), .A2(n79), .Z(Ciphertext[132]) );
  XOR2_X1 U13311 ( .A1(n6839), .A2(n6743), .Z(\MC_ARK_ARC_1_1/temp5[146] ) );
  XOR2_X1 U13312 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[146] ), .A2(\RI5[1][92] ), 
        .Z(n6743) );
  NAND3_X2 U13313 ( .A1(\SB1_3_27/i0[10] ), .A2(\SB1_3_27/i1[9] ), .A3(
        \SB1_3_27/i1_5 ), .ZN(\SB1_3_27/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U13314 ( .A1(\SB2_0_0/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_0/Component_Function_4/NAND4_in[0] ), .A4(n6744), .ZN(
        \SB2_0_0/buf_output[4] ) );
  NAND3_X2 U13315 ( .A1(\SB2_0_0/i0[10] ), .A2(\SB2_0_0/i0[9] ), .A3(
        \SB2_0_0/i0_3 ), .ZN(n6744) );
  XOR2_X1 U13316 ( .A1(\MC_ARK_ARC_1_3/temp6[72] ), .A2(n6745), .Z(
        \MC_ARK_ARC_1_3/buf_output[72] ) );
  XOR2_X1 U13317 ( .A1(\MC_ARK_ARC_1_3/temp2[72] ), .A2(
        \MC_ARK_ARC_1_3/temp1[72] ), .Z(n6745) );
  NAND3_X1 U13318 ( .A1(\SB1_0_4/i0_3 ), .A2(\SB1_0_4/i0[8] ), .A3(
        \SB1_0_4/i1_7 ), .ZN(\SB1_0_4/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U13319 ( .A1(n6748), .A2(n88), .Z(Ciphertext[126]) );
  NAND4_X2 U13320 ( .A1(n3157), .A2(n6816), .A3(n3158), .A4(
        \SB4_10/Component_Function_0/NAND4_in[0] ), .ZN(n6748) );
  NAND3_X1 U13321 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i0[9] ), .A3(
        \SB4_10/i0_3 ), .ZN(n5275) );
  XOR2_X1 U13322 ( .A1(n6749), .A2(n2855), .Z(\MC_ARK_ARC_1_4/buf_output[115] ) );
  XOR2_X1 U13323 ( .A1(\MC_ARK_ARC_1_4/temp2[115] ), .A2(
        \MC_ARK_ARC_1_4/temp1[115] ), .Z(n6749) );
  NAND4_X2 U13324 ( .A1(\SB3_29/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_29/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_3/NAND4_in[0] ), .A4(n6750), .ZN(
        \SB3_29/buf_output[3] ) );
  NAND3_X1 U13325 ( .A1(\SB3_29/i1_5 ), .A2(\SB3_29/i0[8] ), .A3(
        \SB3_29/i3[0] ), .ZN(n6750) );
  NAND4_X2 U13326 ( .A1(\SB3_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_14/Component_Function_2/NAND4_in[3] ), .A3(n4412), .A4(n6752), 
        .ZN(\SB3_14/buf_output[2] ) );
  NAND3_X1 U13327 ( .A1(\SB3_29/i0[10] ), .A2(\RI1[5][17] ), .A3(
        \SB3_29/i0[9] ), .ZN(\SB3_29/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U13328 ( .A1(\RI5[4][46] ), .A2(\RI5[4][10] ), .Z(
        \MC_ARK_ARC_1_4/temp3[136] ) );
  XOR2_X1 U13329 ( .A1(\RI5[2][159] ), .A2(\RI5[2][135] ), .Z(n3872) );
  NAND3_X2 U13330 ( .A1(\SB2_4_2/i0_3 ), .A2(\SB2_4_2/i0_4 ), .A3(
        \SB2_4_2/i1[9] ), .ZN(n6753) );
  XOR2_X1 U13331 ( .A1(\MC_ARK_ARC_1_3/temp5[44] ), .A2(n2077), .Z(
        \MC_ARK_ARC_1_3/buf_output[44] ) );
  XOR2_X1 U13332 ( .A1(\MC_ARK_ARC_1_0/temp5[149] ), .A2(n1203), .Z(n1482) );
  NAND4_X2 U13333 ( .A1(\SB2_4_22/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_4_22/Component_Function_3/NAND4_in[0] ), .A3(n7131), .A4(
        \SB2_4_22/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_4_22/buf_output[3] ) );
  NAND3_X2 U13334 ( .A1(\SB2_4_31/i0[7] ), .A2(\SB2_4_31/i0_3 ), .A3(
        \SB2_4_31/i0_0 ), .ZN(n3423) );
  XOR2_X1 U13335 ( .A1(\RI5[2][38] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[74] ), 
        .Z(n4846) );
  XOR2_X1 U13336 ( .A1(\MC_ARK_ARC_1_2/temp2[44] ), .A2(n6754), .Z(
        \MC_ARK_ARC_1_2/temp5[44] ) );
  XOR2_X1 U13337 ( .A1(\RI5[2][38] ), .A2(\RI5[2][44] ), .Z(n6754) );
  NAND4_X2 U13338 ( .A1(n2416), .A2(
        \SB2_2_22/Component_Function_0/NAND4_in[1] ), .A3(n6905), .A4(
        \SB2_2_22/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_22/buf_output[0] ) );
  NAND4_X2 U13339 ( .A1(n1420), .A2(
        \SB1_2_28/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_5/NAND4_in[0] ), .A4(n6755), .ZN(
        \SB1_2_28/buf_output[5] ) );
  NAND3_X2 U13340 ( .A1(\SB1_2_28/i0[9] ), .A2(\SB1_2_28/i0[6] ), .A3(
        \SB1_2_28/i0_4 ), .ZN(n6755) );
  XOR2_X1 U13341 ( .A1(\MC_ARK_ARC_1_3/temp6[1] ), .A2(n1705), .Z(
        \MC_ARK_ARC_1_3/buf_output[1] ) );
  INV_X2 U13342 ( .I(\SB1_3_24/buf_output[2] ), .ZN(\SB2_3_21/i1[9] ) );
  NAND4_X2 U13343 ( .A1(\SB1_3_24/Component_Function_2/NAND4_in[1] ), .A2(
        n3770), .A3(\SB1_3_24/Component_Function_2/NAND4_in[0] ), .A4(n6968), 
        .ZN(\SB1_3_24/buf_output[2] ) );
  XOR2_X1 U13344 ( .A1(n1672), .A2(\MC_ARK_ARC_1_4/temp1[147] ), .Z(n6756) );
  NAND4_X2 U13345 ( .A1(\SB3_16/Component_Function_4/NAND4_in[3] ), .A2(
        \SB3_16/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_16/Component_Function_4/NAND4_in[1] ), .A4(n6757), .ZN(
        \SB3_16/buf_output[4] ) );
  NAND3_X1 U13346 ( .A1(\SB3_16/i0[9] ), .A2(\SB3_16/i0_3 ), .A3(
        \SB3_16/i0[10] ), .ZN(n6757) );
  XOR2_X1 U13347 ( .A1(n6759), .A2(n6758), .Z(n6786) );
  XOR2_X1 U13348 ( .A1(\RI5[1][14] ), .A2(\SB2_1_22/buf_output[2] ), .Z(n6758)
         );
  XOR2_X1 U13349 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[50] ), .A2(\RI5[1][170] ), 
        .Z(n6759) );
  NAND3_X2 U13350 ( .A1(\SB2_1_23/i0[10] ), .A2(\SB2_1_23/i0_0 ), .A3(
        \SB2_1_23/i0[6] ), .ZN(\SB2_1_23/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U13351 ( .A1(n1958), .A2(
        \SB1_3_17/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_3_17/Component_Function_3/NAND4_in[3] ), .A4(n6761), .ZN(
        \SB1_3_17/buf_output[3] ) );
  NAND3_X2 U13352 ( .A1(\SB1_3_17/i0_3 ), .A2(\SB1_3_17/i0_4 ), .A3(
        \SB1_3_17/i0_0 ), .ZN(n6761) );
  XOR2_X1 U13353 ( .A1(n6763), .A2(n6762), .Z(n1596) );
  XOR2_X1 U13354 ( .A1(\RI5[1][143] ), .A2(\RI5[1][149] ), .Z(n6762) );
  XOR2_X1 U13355 ( .A1(\RI5[1][119] ), .A2(\RI5[1][95] ), .Z(n6763) );
  XOR2_X1 U13356 ( .A1(n6764), .A2(\MC_ARK_ARC_1_1/temp3[69] ), .Z(n2222) );
  XOR2_X1 U13357 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[15] ), .A2(\RI5[1][39] ), 
        .Z(n6764) );
  INV_X4 U13358 ( .I(n7587), .ZN(\SB1_4_6/buf_output[4] ) );
  NAND2_X1 U13359 ( .A1(\SB1_4_6/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_4_6/Component_Function_4/NAND4_in[0] ), .ZN(n7004) );
  XOR2_X1 U13360 ( .A1(\MC_ARK_ARC_1_0/temp2[95] ), .A2(n6765), .Z(n2318) );
  XOR2_X1 U13361 ( .A1(\RI5[0][95] ), .A2(\RI5[0][89] ), .Z(n6765) );
  NAND4_X2 U13362 ( .A1(\SB1_3_16/Component_Function_3/NAND4_in[1] ), .A2(
        n4732), .A3(n4639), .A4(n6767), .ZN(\SB1_3_16/buf_output[3] ) );
  NAND3_X2 U13363 ( .A1(\SB1_3_16/i0[10] ), .A2(\SB1_3_16/i1[9] ), .A3(
        \SB1_3_16/i1_7 ), .ZN(n6767) );
  NAND3_X2 U13364 ( .A1(\SB1_1_12/i0[8] ), .A2(\SB1_1_12/i1_5 ), .A3(
        \SB1_1_12/i3[0] ), .ZN(n6768) );
  XOR2_X1 U13365 ( .A1(n6770), .A2(n6769), .Z(n3953) );
  XOR2_X1 U13366 ( .A1(\RI5[2][77] ), .A2(n140), .Z(n6769) );
  XOR2_X1 U13367 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[41] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[35] ), .Z(n6770) );
  NAND4_X2 U13368 ( .A1(\SB2_1_29/Component_Function_5/NAND4_in[2] ), .A2(
        n1582), .A3(n6919), .A4(\SB2_1_29/Component_Function_5/NAND4_in[0] ), 
        .ZN(\SB2_1_29/buf_output[5] ) );
  NAND4_X2 U13369 ( .A1(\SB1_1_31/Component_Function_3/NAND4_in[0] ), .A2(
        n2519), .A3(\SB1_1_31/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_1_31/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_31/buf_output[3] ) );
  NAND3_X2 U13370 ( .A1(\SB1_4_19/i0[10] ), .A2(\SB1_4_19/i1_5 ), .A3(
        \SB1_4_19/i1[9] ), .ZN(n7140) );
  NAND3_X1 U13371 ( .A1(\SB3_7/i0_0 ), .A2(\SB3_7/i0[8] ), .A3(\SB3_7/i0[9] ), 
        .ZN(\SB3_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U13372 ( .A1(\SB2_0_22/i0_3 ), .A2(\RI3[0][55] ), .A3(
        \SB2_0_22/i1[9] ), .ZN(n3652) );
  NAND4_X2 U13373 ( .A1(n7585), .A2(\SB2_1_7/Component_Function_5/NAND4_in[2] ), .A3(\SB2_1_7/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_7/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_7/buf_output[5] ) );
  INV_X1 U13374 ( .I(\SB3_25/buf_output[5] ), .ZN(\SB4_25/i1_5 ) );
  NAND4_X2 U13375 ( .A1(\SB3_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_25/Component_Function_5/NAND4_in[1] ), .A3(n7429), .A4(
        \SB3_25/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_25/buf_output[5] ) );
  XOR2_X1 U13376 ( .A1(n2278), .A2(n6771), .Z(\MC_ARK_ARC_1_4/buf_output[103] ) );
  XOR2_X1 U13377 ( .A1(\MC_ARK_ARC_1_4/temp2[103] ), .A2(
        \MC_ARK_ARC_1_4/temp1[103] ), .Z(n6771) );
  NAND3_X1 U13378 ( .A1(\SB1_1_11/i0[9] ), .A2(\SB1_1_11/i0[6] ), .A3(
        \SB1_1_11/i1_5 ), .ZN(\SB1_1_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U13379 ( .A1(\SB4_2/i0[10] ), .A2(\SB4_2/i1[9] ), .A3(\SB4_2/i1_7 ), 
        .ZN(\SB4_2/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U13380 ( .A1(\SB1_4_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_4_27/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_4_27/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_4_27/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_4_27/buf_output[1] ) );
  NAND3_X1 U13381 ( .A1(\SB1_4_27/i0_3 ), .A2(\SB1_4_27/i0[8] ), .A3(
        \SB1_4_27/i1_7 ), .ZN(\SB1_4_27/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U13382 ( .A1(n6772), .A2(n7509), .Z(\MC_ARK_ARC_1_2/temp5[8] ) );
  XOR2_X1 U13383 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), .A2(\RI5[2][2] ), 
        .Z(n6772) );
  NAND4_X2 U13384 ( .A1(\SB4_26/Component_Function_3/NAND4_in[3] ), .A2(n4990), 
        .A3(n1237), .A4(n6773), .ZN(n4790) );
  NAND3_X1 U13385 ( .A1(\SB4_26/i0_3 ), .A2(\SB3_27/buf_output[4] ), .A3(
        \SB3_29/buf_output[2] ), .ZN(n6773) );
  INV_X2 U13386 ( .I(\SB1_1_3/buf_output[2] ), .ZN(\SB2_1_0/i1[9] ) );
  NAND2_X2 U13387 ( .A1(\SB2_2_11/i0_0 ), .A2(\SB2_2_11/i3[0] ), .ZN(n6775) );
  NAND3_X1 U13388 ( .A1(\SB3_29/i0[10] ), .A2(\SB3_29/i1_5 ), .A3(
        \SB3_29/i1[9] ), .ZN(\SB3_29/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U13389 ( .A1(n1534), .A2(n1535), .Z(\MC_ARK_ARC_1_4/buf_output[15] )
         );
  NAND3_X1 U13390 ( .A1(\SB1_3_24/i0_3 ), .A2(\SB1_3_24/i0[10] ), .A3(
        \SB1_3_24/i0_4 ), .ZN(\SB1_3_24/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U13391 ( .A1(\SB2_4_13/Component_Function_2/NAND4_in[0] ), .A2(
        n7541), .A3(\SB2_4_13/Component_Function_2/NAND4_in[2] ), .A4(n6776), 
        .ZN(\SB2_4_13/buf_output[2] ) );
  NAND3_X2 U13392 ( .A1(\SB2_4_13/i0_4 ), .A2(\SB2_4_13/i1_5 ), .A3(
        \SB2_4_13/i0_0 ), .ZN(n6776) );
  NAND4_X2 U13393 ( .A1(n3766), .A2(\SB2_2_7/Component_Function_5/NAND4_in[1] ), .A3(\SB2_2_7/Component_Function_5/NAND4_in[0] ), .A4(n6777), .ZN(
        \SB2_2_7/buf_output[5] ) );
  NAND3_X2 U13394 ( .A1(\SB2_2_7/i0[6] ), .A2(\SB2_2_7/i0[9] ), .A3(
        \SB2_2_7/i0_4 ), .ZN(n6777) );
  NAND3_X1 U13395 ( .A1(\SB3_19/i0_4 ), .A2(\SB3_19/i1_7 ), .A3(\SB3_19/i0[8] ), .ZN(n6779) );
  INV_X1 U13396 ( .I(\SB1_4_14/buf_output[0] ), .ZN(\SB2_4_9/i3[0] ) );
  NAND4_X2 U13397 ( .A1(\SB1_4_14/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_14/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_4_14/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_4_14/buf_output[0] ) );
  XOR2_X1 U13398 ( .A1(\MC_ARK_ARC_1_0/temp4[74] ), .A2(n6780), .Z(n3691) );
  XOR2_X1 U13399 ( .A1(\RI5[0][140] ), .A2(\RI5[0][176] ), .Z(n6780) );
  XOR2_X1 U13400 ( .A1(\MC_ARK_ARC_1_3/temp6[184] ), .A2(n6781), .Z(
        \MC_ARK_ARC_1_3/buf_output[184] ) );
  XOR2_X1 U13401 ( .A1(n6782), .A2(n149), .Z(Ciphertext[86]) );
  NAND4_X2 U13402 ( .A1(\SB4_17/Component_Function_2/NAND4_in[3] ), .A2(n6837), 
        .A3(\SB4_17/Component_Function_2/NAND4_in[1] ), .A4(n7557), .ZN(n6782)
         );
  XOR2_X1 U13403 ( .A1(\RI5[3][56] ), .A2(n61), .Z(n6783) );
  XOR2_X1 U13404 ( .A1(\RI5[3][92] ), .A2(\RI5[3][50] ), .Z(n6784) );
  XOR2_X1 U13405 ( .A1(n6786), .A2(n6785), .Z(\MC_ARK_ARC_1_1/buf_output[104] ) );
  XOR2_X1 U13406 ( .A1(\MC_ARK_ARC_1_1/temp4[104] ), .A2(
        \MC_ARK_ARC_1_1/temp1[104] ), .Z(n6785) );
  NAND3_X2 U13407 ( .A1(\SB1_4_30/i0[9] ), .A2(\SB1_4_30/i0_3 ), .A3(
        \SB1_4_30/i0[8] ), .ZN(n6789) );
  XOR2_X1 U13408 ( .A1(n6790), .A2(\MC_ARK_ARC_1_0/temp5[15] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[15] ) );
  XOR2_X1 U13409 ( .A1(\MC_ARK_ARC_1_0/temp3[15] ), .A2(
        \MC_ARK_ARC_1_0/temp4[15] ), .Z(n6790) );
  NAND4_X2 U13410 ( .A1(n6792), .A2(n6791), .A3(
        \SB2_0_25/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_0_25/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB2_0_25/buf_output[0] ) );
  NAND3_X1 U13411 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB2_0_25/i0[10] ), .A3(
        \SB2_0_25/i0_4 ), .ZN(n6792) );
  XOR2_X1 U13412 ( .A1(\RI5[1][87] ), .A2(\RI5[1][93] ), .Z(n1678) );
  NAND4_X2 U13413 ( .A1(\SB1_2_16/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_16/Component_Function_1/NAND4_in[0] ), .A4(n6793), .ZN(
        \SB1_2_16/buf_output[1] ) );
  NAND3_X1 U13414 ( .A1(\SB1_2_16/i0[8] ), .A2(\SB1_2_16/i0_4 ), .A3(
        \SB1_2_16/i1_7 ), .ZN(n6793) );
  XOR2_X1 U13415 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[24] ), .A2(\RI5[3][30] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[30] ) );
  XOR2_X1 U13416 ( .A1(\MC_ARK_ARC_1_3/temp6[30] ), .A2(
        \MC_ARK_ARC_1_3/temp5[30] ), .Z(\MC_ARK_ARC_1_3/buf_output[30] ) );
  XOR2_X1 U13417 ( .A1(n2525), .A2(\MC_ARK_ARC_1_4/temp5[13] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[13] ) );
  NAND4_X2 U13418 ( .A1(\SB2_3_13/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_13/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_3_13/Component_Function_1/NAND4_in[0] ), .A4(n6794), .ZN(
        \SB2_3_13/buf_output[1] ) );
  XOR2_X1 U13419 ( .A1(\RI5[3][63] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[39] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[93] ) );
  NAND4_X2 U13420 ( .A1(n6927), .A2(\SB1_3_0/Component_Function_0/NAND4_in[1] ), .A3(\SB1_3_0/Component_Function_0/NAND4_in[0] ), .A4(n6796), .ZN(
        \SB1_3_0/buf_output[0] ) );
  NAND3_X2 U13421 ( .A1(\SB1_1_22/i0_3 ), .A2(\SB1_1_22/i0[7] ), .A3(
        \SB1_1_22/i0_0 ), .ZN(n2229) );
  XOR2_X1 U13422 ( .A1(\RI5[0][104] ), .A2(\RI5[0][68] ), .Z(
        \MC_ARK_ARC_1_0/temp3[2] ) );
  AND2_X1 U13423 ( .A1(\SB1_1_3/Component_Function_4/NAND4_in[2] ), .A2(n6798), 
        .Z(n2398) );
  NAND3_X1 U13424 ( .A1(\SB1_1_3/i0_0 ), .A2(\SB1_1_3/i0[8] ), .A3(
        \SB1_1_3/i0[9] ), .ZN(n6798) );
  INV_X2 U13425 ( .I(\SB1_3_29/buf_output[5] ), .ZN(\SB2_3_29/i1_5 ) );
  XOR2_X1 U13426 ( .A1(n6799), .A2(n111), .Z(Ciphertext[60]) );
  NAND4_X2 U13427 ( .A1(n3820), .A2(\SB4_21/Component_Function_0/NAND4_in[2] ), 
        .A3(\SB4_21/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_21/Component_Function_0/NAND4_in[3] ), .ZN(n6799) );
  NAND4_X2 U13428 ( .A1(\SB1_3_0/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_0/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_3_0/Component_Function_1/NAND4_in[3] ), .A4(n6801), .ZN(
        \SB1_3_0/buf_output[1] ) );
  XOR2_X1 U13429 ( .A1(n6802), .A2(n170), .Z(Ciphertext[53]) );
  NAND4_X2 U13430 ( .A1(\SB4_23/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_23/Component_Function_5/NAND4_in[1] ), .A3(n649), .A4(
        \SB4_23/Component_Function_5/NAND4_in[0] ), .ZN(n6802) );
  XOR2_X1 U13431 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[122] ), .A2(\RI5[1][86] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[20] ) );
  NAND3_X2 U13432 ( .A1(\SB2_4_8/i0[10] ), .A2(\SB2_4_8/i0_0 ), .A3(
        \SB2_4_8/i0[6] ), .ZN(n7412) );
  NAND3_X2 U13433 ( .A1(\SB2_2_18/i0[10] ), .A2(\SB2_2_18/i1_5 ), .A3(
        \SB2_2_18/i1[9] ), .ZN(\SB2_2_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U13434 ( .A1(\SB1_2_16/i0[9] ), .A2(\SB1_2_16/i0[6] ), .A3(
        \SB1_2_16/i0_4 ), .ZN(n7212) );
  NAND3_X2 U13435 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0[8] ), .A3(
        \SB2_2_0/i0[9] ), .ZN(\SB2_2_0/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U13436 ( .A1(\SB2_3_31/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_3_31/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_31/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_31/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_3_31/buf_output[2] ) );
  NAND4_X2 U13437 ( .A1(\SB3_23/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_23/Component_Function_3/NAND4_in[1] ), .A3(n5118), .A4(n7071), 
        .ZN(\SB3_23/buf_output[3] ) );
  XOR2_X1 U13438 ( .A1(\RI5[0][59] ), .A2(\RI5[0][5] ), .Z(n6804) );
  XOR2_X1 U13439 ( .A1(n6842), .A2(n1263), .Z(\MC_ARK_ARC_1_1/buf_output[7] )
         );
  XOR2_X1 U13440 ( .A1(n6805), .A2(n54), .Z(Ciphertext[78]) );
  NAND4_X2 U13441 ( .A1(\SB4_18/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_18/Component_Function_0/NAND4_in[3] ), .A4(
        \SB4_18/Component_Function_0/NAND4_in[0] ), .ZN(n6805) );
  NAND4_X2 U13442 ( .A1(\SB1_4_10/Component_Function_2/NAND4_in[0] ), .A2(
        n7146), .A3(\SB1_4_10/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_4_10/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_4_10/buf_output[2] ) );
  NAND4_X2 U13443 ( .A1(n4246), .A2(
        \SB1_4_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_4_10/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_4_10/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_4_10/buf_output[3] ) );
  NAND3_X2 U13444 ( .A1(\SB2_1_29/i0[10] ), .A2(\SB2_1_29/i0_3 ), .A3(
        \SB2_1_29/i0[6] ), .ZN(\SB2_1_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U13445 ( .A1(\SB2_1_20/i0[8] ), .A2(\SB2_1_20/i0_4 ), .A3(
        \SB2_1_20/i1_7 ), .ZN(n4074) );
  NAND4_X2 U13446 ( .A1(\SB2_3_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_21/Component_Function_2/NAND4_in[2] ), .A3(n6853), .A4(n7013), 
        .ZN(\SB2_3_21/buf_output[2] ) );
  XOR2_X1 U13447 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[5] ), .A2(\RI5[3][191] ), 
        .Z(n7339) );
  NAND3_X1 U13448 ( .A1(\SB1_3_30/i0_4 ), .A2(\SB1_3_30/i1[9] ), .A3(
        \SB1_3_30/i1_5 ), .ZN(n6811) );
  INV_X1 U13449 ( .I(\SB3_7/buf_output[3] ), .ZN(\SB4_5/i0[8] ) );
  NAND4_X2 U13450 ( .A1(\SB3_7/Component_Function_3/NAND4_in[1] ), .A2(n2436), 
        .A3(n7577), .A4(\SB3_7/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB3_7/buf_output[3] ) );
  XOR2_X1 U13451 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[20] ), .A2(\RI5[3][56] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[146] ) );
  NAND4_X2 U13452 ( .A1(n4763), .A2(
        \SB1_1_22/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_22/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_1_22/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_1_22/buf_output[4] ) );
  XOR2_X1 U13453 ( .A1(n4743), .A2(n6806), .Z(\MC_ARK_ARC_1_1/buf_output[91] )
         );
  XOR2_X1 U13454 ( .A1(\MC_ARK_ARC_1_1/temp1[91] ), .A2(
        \MC_ARK_ARC_1_1/temp2[91] ), .Z(n6806) );
  XOR2_X1 U13455 ( .A1(\MC_ARK_ARC_1_0/temp1[44] ), .A2(n6807), .Z(n4404) );
  XOR2_X1 U13456 ( .A1(\RI5[0][14] ), .A2(\RI5[0][182] ), .Z(n6807) );
  NAND4_X2 U13457 ( .A1(n3029), .A2(\SB2_4_5/Component_Function_4/NAND4_in[1] ), .A3(\SB2_4_5/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_4_5/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_4_5/buf_output[4] ) );
  NAND4_X2 U13458 ( .A1(\SB3_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_3/NAND4_in[2] ), .A3(
        \SB3_11/Component_Function_3/NAND4_in[3] ), .A4(
        \SB3_11/Component_Function_3/NAND4_in[1] ), .ZN(\SB4_9/i0[10] ) );
  XOR2_X1 U13459 ( .A1(n3049), .A2(n6808), .Z(\MC_ARK_ARC_1_2/buf_output[32] )
         );
  XOR2_X1 U13460 ( .A1(\MC_ARK_ARC_1_3/temp2[25] ), .A2(n6812), .Z(n7031) );
  XOR2_X1 U13461 ( .A1(\RI5[3][25] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[19] ), 
        .Z(n6812) );
  XOR2_X1 U13462 ( .A1(n6814), .A2(n6813), .Z(\MC_ARK_ARC_1_1/temp6[98] ) );
  XOR2_X1 U13463 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[164] ), .A2(n536), .Z(
        n6813) );
  XOR2_X1 U13464 ( .A1(n3168), .A2(\RI5[1][134] ), .Z(n6814) );
  XOR2_X1 U13465 ( .A1(n6815), .A2(\MC_ARK_ARC_1_2/temp2[80] ), .Z(
        \MC_ARK_ARC_1_2/temp5[80] ) );
  XOR2_X1 U13466 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[74] ), .A2(\RI5[2][80] ), 
        .Z(n6815) );
  NAND4_X2 U13467 ( .A1(\SB2_3_7/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_7/Component_Function_1/NAND4_in[1] ), .A3(n5088), .A4(
        \SB2_3_7/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_7/buf_output[1] ) );
  INV_X1 U13468 ( .I(\SB1_3_11/buf_output[1] ), .ZN(\SB2_3_7/i1_7 ) );
  NAND4_X2 U13469 ( .A1(\SB1_3_11/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_3_11/Component_Function_1/NAND4_in[1] ), .A3(n4885), .A4(
        \SB1_3_11/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_11/buf_output[1] ) );
  NAND3_X1 U13470 ( .A1(\SB4_10/i0[6] ), .A2(\SB4_10/i0[7] ), .A3(
        \SB4_10/i0[8] ), .ZN(n6816) );
  INV_X2 U13471 ( .I(\SB1_2_9/buf_output[2] ), .ZN(\SB2_2_6/i1[9] ) );
  NAND4_X2 U13472 ( .A1(\SB1_2_9/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_9/Component_Function_2/NAND4_in[3] ), .A3(n3548), .A4(n4411), 
        .ZN(\SB1_2_9/buf_output[2] ) );
  XOR2_X1 U13473 ( .A1(\MC_ARK_ARC_1_1/temp1[65] ), .A2(n6817), .Z(
        \MC_ARK_ARC_1_1/temp5[65] ) );
  XOR2_X1 U13474 ( .A1(\RI5[1][11] ), .A2(\RI5[1][35] ), .Z(n6817) );
  NAND4_X2 U13475 ( .A1(\SB2_4_23/Component_Function_5/NAND4_in[1] ), .A2(
        n4784), .A3(\SB2_4_23/Component_Function_5/NAND4_in[0] ), .A4(n6818), 
        .ZN(\SB2_4_23/buf_output[5] ) );
  NAND3_X2 U13476 ( .A1(\SB2_4_23/i0[6] ), .A2(\SB2_4_23/i0_4 ), .A3(
        \SB2_4_23/i0[9] ), .ZN(n6818) );
  NAND3_X2 U13477 ( .A1(\SB2_3_5/i0[10] ), .A2(\SB2_3_5/i0_4 ), .A3(
        \SB2_3_5/i0_3 ), .ZN(\SB2_3_5/Component_Function_0/NAND4_in[2] ) );
  INV_X1 U13478 ( .I(\SB1_4_9/buf_output[1] ), .ZN(\SB2_4_5/i1_7 ) );
  NAND4_X2 U13479 ( .A1(\SB1_4_9/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_4_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_4_9/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_4_9/buf_output[1] ) );
  BUF_X2 U13480 ( .I(\SB2_3_20/i0[7] ), .Z(n6819) );
  NAND3_X1 U13481 ( .A1(\SB4_21/i0_3 ), .A2(\SB3_24/buf_output[2] ), .A3(
        \SB4_21/i0[7] ), .ZN(\SB4_21/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U13482 ( .A1(n4393), .A2(\SB3_21/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB3_21/Component_Function_5/NAND4_in[0] ), .A4(n6820), .ZN(
        \SB3_21/buf_output[5] ) );
  NAND3_X1 U13483 ( .A1(\SB2_1_16/i0_3 ), .A2(\SB1_1_17/buf_output[4] ), .A3(
        \SB2_1_16/i1[9] ), .ZN(n3149) );
  NAND4_X2 U13484 ( .A1(\SB2_0_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_0_5/Component_Function_2/NAND4_in[1] ), .A4(n6822), .ZN(
        \SB2_0_5/buf_output[2] ) );
  NAND3_X2 U13485 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0[8] ), .A3(
        \SB2_0_5/i0[9] ), .ZN(n6822) );
  NAND4_X2 U13486 ( .A1(\SB1_2_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_2_28/Component_Function_2/NAND4_in[1] ), .A4(n7352), .ZN(
        \SB1_2_28/buf_output[2] ) );
  NAND4_X2 U13487 ( .A1(\SB3_28/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_28/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_28/Component_Function_4/NAND4_in[3] ), .A4(n6823), .ZN(
        \SB3_28/buf_output[4] ) );
  NAND3_X2 U13488 ( .A1(\SB1_1_13/i0_0 ), .A2(\SB1_1_13/i1_5 ), .A3(
        \SB1_1_13/i0_4 ), .ZN(\SB1_1_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U13489 ( .A1(\SB1_2_8/i0_3 ), .A2(\SB1_2_8/i0_4 ), .A3(
        \SB1_2_8/i1[9] ), .ZN(\SB1_2_8/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U13490 ( .A1(\SB1_0_5/i0_3 ), .A2(\SB1_0_5/i0[9] ), .A3(
        \SB1_0_5/i0[8] ), .ZN(\SB1_0_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U13491 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i0_0 ), .A3(
        \SB2_3_27/i0_4 ), .ZN(\SB2_3_27/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U13492 ( .A1(n2829), .A2(
        \SB1_0_18/Component_Function_2/NAND4_in[2] ), .ZN(n6824) );
  NAND2_X1 U13493 ( .A1(\SB1_0_18/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_18/Component_Function_2/NAND4_in[0] ), .ZN(n6825) );
  XOR2_X1 U13494 ( .A1(n3391), .A2(n7317), .Z(n862) );
  NAND3_X1 U13495 ( .A1(\SB2_0_2/i0_0 ), .A2(\SB2_0_2/i0_3 ), .A3(
        \SB2_0_2/i0[7] ), .ZN(\SB2_0_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U13496 ( .A1(\SB4_19/i0_3 ), .A2(\SB4_19/i1[9] ), .A3(\SB4_19/i0_4 ), .ZN(n7132) );
  NAND3_X1 U13497 ( .A1(\SB4_19/i0_3 ), .A2(\SB4_19/i0[7] ), .A3(\SB4_19/i0_0 ), .ZN(\SB4_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U13498 ( .A1(\SB4_19/i0_3 ), .A2(\SB4_19/i0_0 ), .A3(\SB4_19/i0_4 ), 
        .ZN(\SB4_19/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U13499 ( .A1(\RI5[0][59] ), .A2(\RI5[0][191] ), .Z(n6826) );
  XOR2_X1 U13500 ( .A1(n6827), .A2(\MC_ARK_ARC_1_4/temp6[50] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[50] ) );
  NAND3_X1 U13501 ( .A1(\SB3_20/i0[8] ), .A2(\SB3_20/i1_5 ), .A3(
        \SB3_20/i3[0] ), .ZN(n7240) );
  INV_X2 U13502 ( .I(\RI3[0][171] ), .ZN(\SB2_0_3/i0[8] ) );
  NAND4_X2 U13503 ( .A1(\SB1_0_5/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_5/Component_Function_3/NAND4_in[0] ), .A4(n7475), .ZN(
        \RI3[0][171] ) );
  NAND4_X2 U13504 ( .A1(\SB1_4_14/Component_Function_1/NAND4_in[1] ), .A2(
        n1106), .A3(\SB1_4_14/Component_Function_1/NAND4_in[3] ), .A4(n6829), 
        .ZN(\RI3[4][127] ) );
  NAND3_X2 U13505 ( .A1(\SB2_1_31/i0[6] ), .A2(\SB2_1_31/i0[10] ), .A3(
        \SB2_1_31/i0_3 ), .ZN(\SB2_1_31/Component_Function_2/NAND4_in[1] ) );
  NAND2_X2 U13506 ( .A1(n572), .A2(n959), .ZN(\SB2_3_5/i0_4 ) );
  NAND4_X2 U13507 ( .A1(\SB2_3_20/Component_Function_5/NAND4_in[2] ), .A2(
        n2174), .A3(\SB2_3_20/Component_Function_5/NAND4_in[0] ), .A4(n6830), 
        .ZN(\SB2_3_20/buf_output[5] ) );
  NAND3_X2 U13508 ( .A1(\SB2_3_20/i0[9] ), .A2(\RI3[3][70] ), .A3(
        \SB2_3_20/i0[6] ), .ZN(n6830) );
  XOR2_X1 U13509 ( .A1(n6831), .A2(\MC_ARK_ARC_1_0/temp5[71] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[71] ) );
  NAND3_X2 U13510 ( .A1(\SB1_1_12/i0_3 ), .A2(\SB1_1_12/i1[9] ), .A3(
        \SB1_1_12/i0_4 ), .ZN(\SB1_1_12/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U13511 ( .I(\SB1_4_17/buf_output[2] ), .ZN(\SB2_4_14/i1[9] ) );
  NAND4_X2 U13512 ( .A1(\SB1_4_17/Component_Function_2/NAND4_in[0] ), .A2(
        n7375), .A3(\SB1_4_17/Component_Function_2/NAND4_in[1] ), .A4(n4548), 
        .ZN(\SB1_4_17/buf_output[2] ) );
  XOR2_X1 U13513 ( .A1(n6833), .A2(n6832), .Z(\MC_ARK_ARC_1_4/temp5[69] ) );
  XOR2_X1 U13514 ( .A1(\RI5[4][69] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[15] ), 
        .Z(n6832) );
  XOR2_X1 U13515 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[63] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[39] ), .Z(n6833) );
  XOR2_X1 U13516 ( .A1(n6834), .A2(\MC_ARK_ARC_1_0/temp2[159] ), .Z(n2804) );
  XOR2_X1 U13517 ( .A1(\RI5[0][159] ), .A2(\RI5[0][153] ), .Z(n6834) );
  NAND4_X2 U13518 ( .A1(\SB2_0_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_18/Component_Function_4/NAND4_in[3] ), .A4(n6835), .ZN(
        \SB2_0_18/buf_output[4] ) );
  XOR2_X1 U13519 ( .A1(n6836), .A2(\MC_ARK_ARC_1_0/temp1[142] ), .Z(
        \MC_ARK_ARC_1_0/temp5[142] ) );
  XOR2_X1 U13520 ( .A1(\RI5[0][88] ), .A2(\RI5[0][112] ), .Z(n6836) );
  NAND3_X1 U13521 ( .A1(\SB4_17/i1[9] ), .A2(n3984), .A3(\SB4_17/i0[10] ), 
        .ZN(n6837) );
  XOR2_X1 U13522 ( .A1(n6838), .A2(n95), .Z(Ciphertext[84]) );
  NAND3_X2 U13523 ( .A1(\SB2_2_22/i0_0 ), .A2(\SB2_2_22/i1_7 ), .A3(
        \SB2_2_22/i3[0] ), .ZN(\SB2_2_22/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U13524 ( .A1(\MC_ARK_ARC_1_4/temp5[145] ), .A2(
        \MC_ARK_ARC_1_4/temp6[145] ), .Z(\MC_ARK_ARC_1_4/buf_output[145] ) );
  XOR2_X1 U13525 ( .A1(\MC_ARK_ARC_1_3/temp5[88] ), .A2(
        \MC_ARK_ARC_1_3/temp6[88] ), .Z(\MC_ARK_ARC_1_3/buf_output[88] ) );
  NAND4_X2 U13526 ( .A1(\SB1_0_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_25/Component_Function_3/NAND4_in[1] ), .A3(n4557), .A4(
        \SB1_0_25/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_0_25/buf_output[3] ) );
  NAND4_X2 U13527 ( .A1(\SB1_3_10/Component_Function_3/NAND4_in[1] ), .A2(
        n7040), .A3(n1304), .A4(\SB1_3_10/Component_Function_3/NAND4_in[0] ), 
        .ZN(\SB1_3_10/buf_output[3] ) );
  XOR2_X1 U13528 ( .A1(\RI5[1][116] ), .A2(\RI5[1][140] ), .Z(n6839) );
  NAND3_X1 U13529 ( .A1(\SB4_17/i1[9] ), .A2(\SB4_17/i0[10] ), .A3(
        \SB4_17/i1_7 ), .ZN(\SB4_17/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U13530 ( .A1(\SB4_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB4_18/Component_Function_2/NAND4_in[2] ), .A3(n5130), .A4(
        \SB4_18/Component_Function_2/NAND4_in[3] ), .ZN(n5131) );
  XOR2_X1 U13531 ( .A1(\RI5[4][100] ), .A2(\RI5[4][124] ), .Z(
        \MC_ARK_ARC_1_4/temp2[154] ) );
  XOR2_X1 U13532 ( .A1(\RI5[1][148] ), .A2(\RI5[1][142] ), .Z(n4056) );
  NAND3_X2 U13533 ( .A1(\SB1_3_25/i0_3 ), .A2(\SB1_3_25/i1[9] ), .A3(
        \SB1_3_25/i0_4 ), .ZN(n1075) );
  XOR2_X1 U13534 ( .A1(n6840), .A2(\MC_ARK_ARC_1_2/temp4[162] ), .Z(
        \MC_ARK_ARC_1_2/temp6[162] ) );
  XOR2_X1 U13535 ( .A1(\RI5[2][36] ), .A2(\RI5[2][72] ), .Z(n6840) );
  NAND4_X2 U13536 ( .A1(n4509), .A2(
        \SB2_2_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_30/Component_Function_0/NAND4_in[0] ), .A4(n6841), .ZN(
        \SB2_2_30/buf_output[0] ) );
  NAND3_X1 U13537 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0_0 ), .A3(
        \SB2_2_30/i0[7] ), .ZN(n6841) );
  XOR2_X1 U13538 ( .A1(\MC_ARK_ARC_1_1/temp4[7] ), .A2(
        \MC_ARK_ARC_1_1/temp3[7] ), .Z(n6842) );
  NAND3_X2 U13539 ( .A1(\SB2_3_24/i0[10] ), .A2(\SB2_3_24/i1_5 ), .A3(
        \SB2_3_24/i1[9] ), .ZN(\SB2_3_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U13540 ( .A1(\SB2_2_7/i0_0 ), .A2(\SB2_2_7/i0_4 ), .A3(
        \SB2_2_7/i1_5 ), .ZN(n6843) );
  NAND4_X2 U13541 ( .A1(n1765), .A2(\SB1_4_0/Component_Function_2/NAND4_in[1] ), .A3(\SB1_4_0/Component_Function_2/NAND4_in[0] ), .A4(n6844), .ZN(
        \SB1_4_0/buf_output[2] ) );
  NAND3_X2 U13542 ( .A1(\SB1_4_0/i1_5 ), .A2(\SB1_4_0/i0_4 ), .A3(
        \SB1_4_0/i0_0 ), .ZN(n6844) );
  NAND2_X2 U13543 ( .A1(\SB1_4_16/i1[9] ), .A2(n6846), .ZN(n6845) );
  NAND4_X2 U13544 ( .A1(\SB1_4_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_4_9/Component_Function_2/NAND4_in[2] ), .A3(n2538), .A4(n6847), 
        .ZN(\SB1_4_9/buf_output[2] ) );
  NAND3_X2 U13545 ( .A1(\SB1_4_9/i0_3 ), .A2(\SB1_4_9/i0[10] ), .A3(
        \SB1_4_9/i0[6] ), .ZN(n6847) );
  OR3_X1 U13546 ( .A1(n6737), .A2(\SB1_2_9/buf_output[3] ), .A3(
        \SB1_2_12/buf_output[0] ), .Z(
        \SB2_2_7/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U13547 ( .A1(\MC_ARK_ARC_1_4/temp2[135] ), .A2(n6848), .Z(
        \MC_ARK_ARC_1_4/temp5[135] ) );
  XOR2_X1 U13548 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[135] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[129] ), .Z(n6848) );
  NAND3_X2 U13549 ( .A1(\SB1_4_1/i0[10] ), .A2(\SB1_4_1/i1_7 ), .A3(
        \SB1_4_1/i1[9] ), .ZN(\SB1_4_1/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U13550 ( .A1(n6850), .A2(n6849), .Z(\RI1[5][80] ) );
  XOR2_X1 U13551 ( .A1(\MC_ARK_ARC_1_4/temp2[80] ), .A2(
        \MC_ARK_ARC_1_4/temp1[80] ), .Z(n6850) );
  NAND4_X2 U13552 ( .A1(\SB2_1_24/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_1_24/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_24/Component_Function_3/NAND4_in[3] ), .A4(n6851), .ZN(
        \SB2_1_24/buf_output[3] ) );
  NAND3_X2 U13553 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0_4 ), .A3(
        \SB2_1_24/i0_0 ), .ZN(n6851) );
  XOR2_X1 U13554 ( .A1(\RI5[1][26] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[164] ), 
        .Z(n7121) );
  XOR2_X1 U13555 ( .A1(n6852), .A2(n2667), .Z(\MC_ARK_ARC_1_3/buf_output[143] ) );
  XOR2_X1 U13556 ( .A1(\MC_ARK_ARC_1_3/temp3[143] ), .A2(
        \MC_ARK_ARC_1_3/temp4[143] ), .Z(n6852) );
  NAND3_X2 U13557 ( .A1(\SB1_3_21/i0[9] ), .A2(\SB1_3_21/i0_4 ), .A3(
        \SB1_3_21/i0[6] ), .ZN(n6854) );
  XOR2_X1 U13558 ( .A1(n6856), .A2(n6855), .Z(\MC_ARK_ARC_1_4/buf_output[109] ) );
  XOR2_X1 U13559 ( .A1(\MC_ARK_ARC_1_4/temp3[109] ), .A2(
        \MC_ARK_ARC_1_4/temp2[109] ), .Z(n6855) );
  XOR2_X1 U13560 ( .A1(\MC_ARK_ARC_1_4/temp1[109] ), .A2(
        \MC_ARK_ARC_1_4/temp4[109] ), .Z(n6856) );
  XOR2_X1 U13561 ( .A1(n6857), .A2(\MC_ARK_ARC_1_4/temp4[135] ), .Z(
        \MC_ARK_ARC_1_4/temp6[135] ) );
  XOR2_X1 U13562 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[45] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[9] ), .Z(n6857) );
  NAND3_X2 U13563 ( .A1(\SB2_1_28/i0[10] ), .A2(\SB2_1_28/i1_7 ), .A3(
        \SB2_1_28/i1[9] ), .ZN(n6858) );
  NAND3_X2 U13564 ( .A1(\SB2_1_28/i0[8] ), .A2(\SB2_1_28/i3[0] ), .A3(
        \SB2_1_28/i1_5 ), .ZN(n6859) );
  NAND3_X2 U13565 ( .A1(\SB1_2_1/i0_0 ), .A2(\SB1_2_1/i0_4 ), .A3(
        \SB1_2_1/i1_5 ), .ZN(n6860) );
  NAND4_X2 U13566 ( .A1(\SB1_3_9/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_9/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_3_9/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_3_9/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_9/buf_output[1] ) );
  NAND4_X2 U13567 ( .A1(\SB1_4_3/Component_Function_2/NAND4_in[1] ), .A2(n1571), .A3(\SB1_4_3/Component_Function_2/NAND4_in[3] ), .A4(n6861), .ZN(
        \RI3[4][188] ) );
  NAND3_X2 U13568 ( .A1(\SB1_4_3/i0[10] ), .A2(\SB1_4_3/i1[9] ), .A3(
        \SB1_4_3/i1_5 ), .ZN(n6861) );
  NAND4_X2 U13569 ( .A1(\SB2_2_21/Component_Function_0/NAND4_in[1] ), .A2(
        n4473), .A3(\SB2_2_21/Component_Function_0/NAND4_in[0] ), .A4(n6862), 
        .ZN(\SB2_2_21/buf_output[0] ) );
  XOR2_X1 U13570 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[60] ), .A2(\RI5[2][54] ), 
        .Z(n893) );
  XOR2_X1 U13571 ( .A1(n742), .A2(n741), .Z(n6865) );
  NAND4_X2 U13572 ( .A1(\SB3_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_28/Component_Function_3/NAND4_in[1] ), .A3(n863), .A4(
        \SB3_28/Component_Function_3/NAND4_in[2] ), .ZN(\SB4_26/i0[10] ) );
  NOR2_X2 U13573 ( .A1(n2374), .A2(n6866), .ZN(n1102) );
  NAND3_X2 U13574 ( .A1(\SB2_2_0/i0[6] ), .A2(\SB2_2_0/i0_0 ), .A3(
        \SB2_2_0/i0[10] ), .ZN(n601) );
  NAND3_X2 U13575 ( .A1(\SB2_1_11/i0_3 ), .A2(\SB2_1_11/i0_0 ), .A3(
        \SB2_1_11/i0_4 ), .ZN(\SB2_1_11/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U13576 ( .A1(\RI5[1][75] ), .A2(\RI5[1][39] ), .Z(n3319) );
  XOR2_X1 U13577 ( .A1(\SB2_0_15/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[75] ), .Z(n2206) );
  NAND4_X2 U13578 ( .A1(\SB2_3_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_2/NAND4_in[1] ), .A3(n1034), .A4(n6867), 
        .ZN(\SB2_3_3/buf_output[2] ) );
  NAND3_X2 U13579 ( .A1(\SB2_3_3/i0_0 ), .A2(\SB2_3_3/i0_4 ), .A3(
        \SB2_3_3/i1_5 ), .ZN(n6867) );
  XOR2_X1 U13580 ( .A1(\MC_ARK_ARC_1_3/temp1[189] ), .A2(n6868), .Z(n1131) );
  XOR2_X1 U13581 ( .A1(\RI5[3][135] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[159] ), .Z(n6868) );
  NAND4_X2 U13582 ( .A1(n2593), .A2(\SB1_4_0/Component_Function_0/NAND4_in[1] ), .A3(\SB1_4_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_0/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_4_0/buf_output[0] ) );
  NAND4_X2 U13583 ( .A1(\SB1_3_1/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_1/Component_Function_4/NAND4_in[0] ), .A3(n6869), .A4(
        \SB1_3_1/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_1/buf_output[4] ) );
  NAND3_X2 U13584 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i0[10] ), .A3(
        \SB2_2_27/i0_4 ), .ZN(n1125) );
  NAND4_X2 U13585 ( .A1(n2151), .A2(n7405), .A3(n911), .A4(
        \SB1_2_27/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_27/buf_output[5] ) );
  NAND3_X1 U13586 ( .A1(\SB4_10/i0[6] ), .A2(\SB4_10/i0_3 ), .A3(
        \SB4_10/i0[10] ), .ZN(n5369) );
  XOR2_X1 U13587 ( .A1(\RI5[4][182] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[86] ), 
        .Z(n6870) );
  XOR2_X1 U13588 ( .A1(\RI5[0][123] ), .A2(\RI5[0][147] ), .Z(
        \MC_ARK_ARC_1_0/temp2[177] ) );
  NAND4_X2 U13589 ( .A1(\SB2_4_14/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_4_14/Component_Function_0/NAND4_in[1] ), .A3(n7462), .A4(n6873), 
        .ZN(\SB2_4_14/buf_output[0] ) );
  NAND2_X1 U13590 ( .A1(\SB2_4_14/i0[9] ), .A2(\SB2_4_14/i0[10] ), .ZN(n6873)
         );
  XOR2_X1 U13591 ( .A1(\MC_ARK_ARC_1_4/temp1[186] ), .A2(
        \MC_ARK_ARC_1_4/temp2[186] ), .Z(n6874) );
  XOR2_X1 U13592 ( .A1(n6876), .A2(n6875), .Z(\MC_ARK_ARC_1_0/temp6[32] ) );
  XOR2_X1 U13593 ( .A1(\RI5[0][134] ), .A2(n107), .Z(n6875) );
  XOR2_X1 U13594 ( .A1(\RI5[0][98] ), .A2(\RI5[0][68] ), .Z(n6876) );
  NAND3_X2 U13595 ( .A1(\SB2_2_10/i0_3 ), .A2(\SB2_2_10/i0[9] ), .A3(
        \SB2_2_10/i0[8] ), .ZN(\SB2_2_10/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U13596 ( .A1(\SB1_4_16/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_16/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_4_16/Component_Function_0/NAND4_in[1] ), .A4(n6877), .ZN(
        \SB1_4_16/buf_output[0] ) );
  NAND3_X2 U13597 ( .A1(\SB1_4_16/i0_3 ), .A2(\SB1_4_16/i0[7] ), .A3(
        \SB1_4_16/i0_0 ), .ZN(n6877) );
  XOR2_X1 U13598 ( .A1(n6878), .A2(n176), .Z(Ciphertext[41]) );
  NAND4_X2 U13599 ( .A1(\SB4_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_25/Component_Function_5/NAND4_in[1] ), .A3(n2213), .A4(
        \SB4_25/Component_Function_5/NAND4_in[0] ), .ZN(n6878) );
  NAND3_X1 U13600 ( .A1(\SB2_3_28/i0_0 ), .A2(\SB2_3_28/i0[8] ), .A3(
        \SB2_3_28/i0[9] ), .ZN(\SB2_3_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U13601 ( .A1(\SB4_18/i0[10] ), .A2(\SB4_18/i0_0 ), .A3(
        \SB4_18/i0[6] ), .ZN(\SB4_18/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U13602 ( .A1(\SB2_4_18/i0_0 ), .A2(\SB2_4_18/i0[9] ), .A3(
        \SB2_4_18/i0[8] ), .ZN(\SB2_4_18/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U13603 ( .A1(\SB2_1_0/Component_Function_3/NAND4_in[3] ), .A2(n4516), .A3(n6889), .A4(n4228), .ZN(\SB2_1_0/buf_output[3] ) );
  INV_X2 U13604 ( .I(\SB1_2_15/buf_output[3] ), .ZN(\SB2_2_13/i0[8] ) );
  NAND4_X2 U13605 ( .A1(\SB2_3_23/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_23/Component_Function_1/NAND4_in[2] ), .A4(n6881), .ZN(
        \SB2_3_23/buf_output[1] ) );
  NAND3_X2 U13606 ( .A1(\SB1_3_11/i0[10] ), .A2(\SB1_3_11/i1[9] ), .A3(
        \SB1_3_11/i1_7 ), .ZN(n6897) );
  NAND3_X2 U13607 ( .A1(\SB2_2_15/i0[8] ), .A2(\SB2_2_15/i3[0] ), .A3(
        \SB2_2_15/i1_5 ), .ZN(\SB2_2_15/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U13608 ( .A1(\SB2_3_8/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_3_8/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_3_8/Component_Function_5/NAND4_in[0] ), .A4(n6882), .ZN(
        \SB2_3_8/buf_output[5] ) );
  XOR2_X1 U13609 ( .A1(\MC_ARK_ARC_1_1/temp1[89] ), .A2(n6883), .Z(
        \MC_ARK_ARC_1_1/temp5[89] ) );
  XOR2_X1 U13610 ( .A1(\RI5[1][59] ), .A2(\RI5[1][35] ), .Z(n6883) );
  XOR2_X1 U13611 ( .A1(\MC_ARK_ARC_1_2/temp6[33] ), .A2(n6884), .Z(
        \MC_ARK_ARC_1_2/buf_output[33] ) );
  XOR2_X1 U13612 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[75] ), .A2(\RI5[0][69] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[75] ) );
  XOR2_X1 U13613 ( .A1(n2831), .A2(n6885), .Z(n2846) );
  XOR2_X1 U13614 ( .A1(\RI5[3][41] ), .A2(\RI5[3][65] ), .Z(n6885) );
  NAND4_X2 U13615 ( .A1(\SB1_2_26/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_26/Component_Function_3/NAND4_in[0] ), .A3(n6957), .A4(n1975), 
        .ZN(\SB1_2_26/buf_output[3] ) );
  NAND3_X2 U13616 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i1[9] ), .A3(
        \SB2_2_12/i0[6] ), .ZN(n6886) );
  NAND4_X2 U13617 ( .A1(\SB1_3_16/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_3_16/Component_Function_4/NAND4_in[3] ), .A3(n4813), .A4(
        \SB1_3_16/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_3_16/buf_output[4] ) );
  XOR2_X1 U13618 ( .A1(\RI5[2][189] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[3] ), 
        .Z(n6887) );
  NAND3_X1 U13619 ( .A1(\SB1_0_18/i0_4 ), .A2(n6290), .A3(\SB1_0_18/i1_5 ), 
        .ZN(n2829) );
  INV_X2 U13620 ( .I(n6888), .ZN(\RI1[5][53] ) );
  XNOR2_X1 U13621 ( .A1(\MC_ARK_ARC_1_4/temp5[53] ), .A2(
        \MC_ARK_ARC_1_4/temp6[53] ), .ZN(n6888) );
  NAND3_X1 U13622 ( .A1(\SB1_0_3/i0_4 ), .A2(\SB1_0_3/i0_0 ), .A3(
        \SB1_0_3/i1_5 ), .ZN(\SB1_0_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U13623 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i1_7 ), .A3(
        \SB2_1_0/i1[9] ), .ZN(n6889) );
  NAND4_X2 U13624 ( .A1(\SB1_3_0/Component_Function_2/NAND4_in[0] ), .A2(n5347), .A3(n5114), .A4(n6890), .ZN(\SB1_3_0/buf_output[2] ) );
  NAND3_X2 U13625 ( .A1(\SB1_3_0/i0_0 ), .A2(\SB1_3_0/i0_4 ), .A3(
        \SB1_3_0/i1_5 ), .ZN(n6890) );
  NAND3_X2 U13626 ( .A1(\SB1_4_0/i0[9] ), .A2(\SB1_4_0/i0[8] ), .A3(
        \SB1_4_0/i0_0 ), .ZN(\SB1_4_0/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U13627 ( .A1(\SB2_2_16/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_2_16/Component_Function_2/NAND4_in[2] ), .A3(n3584), .A4(n6891), 
        .ZN(\SB2_2_16/buf_output[2] ) );
  NAND3_X2 U13628 ( .A1(\SB2_2_16/i0[10] ), .A2(\SB2_2_16/i1_5 ), .A3(
        \SB2_2_16/i1[9] ), .ZN(n6891) );
  NAND3_X2 U13629 ( .A1(\SB1_2_29/i0_4 ), .A2(\SB1_2_29/i0[6] ), .A3(
        \SB1_2_29/i0[9] ), .ZN(n6892) );
  NAND3_X2 U13630 ( .A1(\SB1_2_19/i0[10] ), .A2(\SB1_2_19/i1[9] ), .A3(
        \SB1_2_19/i1_5 ), .ZN(n6893) );
  INV_X2 U13631 ( .I(\SB1_1_5/buf_output[2] ), .ZN(\SB2_1_2/i1[9] ) );
  NAND4_X2 U13632 ( .A1(\SB1_1_5/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_5/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_1_5/Component_Function_2/NAND4_in[2] ), .A4(n7474), .ZN(
        \SB1_1_5/buf_output[2] ) );
  NAND3_X2 U13633 ( .A1(\SB1_1_28/i0[9] ), .A2(\SB1_1_28/i0_4 ), .A3(
        \SB1_1_28/i0[6] ), .ZN(n6894) );
  NAND3_X1 U13634 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i0[6] ), .A3(
        \SB1_0_20/i1[9] ), .ZN(n6895) );
  XOR2_X1 U13635 ( .A1(\RI5[0][38] ), .A2(\RI5[0][32] ), .Z(n6896) );
  INV_X2 U13636 ( .I(\RI3[0][1] ), .ZN(\SB2_0_31/i1_7 ) );
  NAND4_X2 U13637 ( .A1(\SB1_0_3/Component_Function_1/NAND4_in[1] ), .A2(n6958), .A3(\SB1_0_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_3/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][1] ) );
  XOR2_X1 U13638 ( .A1(\RI5[3][70] ), .A2(\SB2_3_20/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/temp1[76] ) );
  NAND4_X2 U13639 ( .A1(\SB2_1_23/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_23/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_1_23/Component_Function_4/NAND4_in[0] ), .A4(n6898), .ZN(
        \SB2_1_23/buf_output[4] ) );
  NAND3_X2 U13640 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0[10] ), .A3(
        \SB2_1_23/i0[9] ), .ZN(n6898) );
  XOR2_X1 U13641 ( .A1(\MC_ARK_ARC_1_2/temp6[121] ), .A2(n5161), .Z(
        \MC_ARK_ARC_1_2/buf_output[121] ) );
  XOR2_X1 U13642 ( .A1(n6900), .A2(n6899), .Z(\MC_ARK_ARC_1_3/buf_output[191] ) );
  XOR2_X1 U13643 ( .A1(n7021), .A2(n4437), .Z(n6899) );
  XOR2_X1 U13644 ( .A1(n3073), .A2(n4438), .Z(n6900) );
  XOR2_X1 U13645 ( .A1(n6902), .A2(n6901), .Z(n5105) );
  XOR2_X1 U13646 ( .A1(\RI5[1][57] ), .A2(n456), .Z(n6901) );
  XOR2_X1 U13647 ( .A1(\RI5[1][183] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[21] ), 
        .Z(n6902) );
  NAND3_X2 U13648 ( .A1(\SB1_1_29/i0_0 ), .A2(\SB1_1_29/i1_5 ), .A3(
        \SB1_1_29/i0_4 ), .ZN(\SB1_1_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U13649 ( .A1(\SB2_4_9/i3[0] ), .A2(\SB2_4_9/i1_5 ), .A3(
        \SB2_4_9/i0[8] ), .ZN(n6914) );
  XOR2_X1 U13650 ( .A1(n709), .A2(n6903), .Z(\MC_ARK_ARC_1_1/buf_output[55] )
         );
  XOR2_X1 U13651 ( .A1(\MC_ARK_ARC_1_1/temp1[55] ), .A2(
        \MC_ARK_ARC_1_1/temp4[55] ), .Z(n6903) );
  NAND3_X1 U13652 ( .A1(\SB4_6/i0[9] ), .A2(\SB4_6/i0_3 ), .A3(\SB4_6/i0[10] ), 
        .ZN(\SB4_6/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U13653 ( .A1(\SB1_4_28/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_4_28/Component_Function_5/NAND4_in[1] ), .A3(n1311), .A4(n6906), 
        .ZN(\SB1_4_28/buf_output[5] ) );
  INV_X2 U13654 ( .I(\SB1_2_12/buf_output[3] ), .ZN(\SB2_2_10/i0[8] ) );
  NAND4_X2 U13655 ( .A1(\SB1_2_12/Component_Function_3/NAND4_in[3] ), .A2(
        n4012), .A3(n7025), .A4(\SB1_2_12/Component_Function_3/NAND4_in[1] ), 
        .ZN(\SB1_2_12/buf_output[3] ) );
  XOR2_X1 U13656 ( .A1(\RI5[3][27] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[21] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[27] ) );
  NAND3_X2 U13657 ( .A1(n6908), .A2(
        \SB1_2_10/Component_Function_1/NAND4_in[0] ), .A3(n6907), .ZN(
        \SB1_2_10/buf_output[1] ) );
  XOR2_X1 U13658 ( .A1(n6910), .A2(\MC_ARK_ARC_1_2/temp6[13] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[13] ) );
  NAND3_X2 U13659 ( .A1(\SB2_4_25/i0[10] ), .A2(\SB2_4_25/i0_3 ), .A3(
        \SB2_4_25/i0[6] ), .ZN(n6911) );
  INV_X2 U13660 ( .I(\SB1_3_23/buf_output[2] ), .ZN(\SB2_3_20/i1[9] ) );
  NAND3_X1 U13661 ( .A1(\SB1_1_5/i0[6] ), .A2(\SB1_1_5/i1[9] ), .A3(
        \SB1_1_5/i0_3 ), .ZN(\SB1_1_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U13662 ( .A1(\SB1_1_23/i0_0 ), .A2(\SB1_1_23/i1_5 ), .A3(
        \SB1_1_23/i0_4 ), .ZN(\SB1_1_23/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U13663 ( .A1(\RI5[0][103] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[97] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[103] ) );
  XOR2_X1 U13664 ( .A1(\MC_ARK_ARC_1_2/temp3[109] ), .A2(
        \MC_ARK_ARC_1_2/temp4[109] ), .Z(\MC_ARK_ARC_1_2/temp6[109] ) );
  NAND4_X2 U13665 ( .A1(\SB1_4_1/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_4_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_4_1/Component_Function_0/NAND4_in[0] ), .A4(n6913), .ZN(
        \SB1_4_1/buf_output[0] ) );
  NAND3_X1 U13666 ( .A1(\SB1_4_1/i0_0 ), .A2(\SB1_4_1/i0[7] ), .A3(
        \SB1_4_1/i0_3 ), .ZN(n6913) );
  NAND4_X2 U13667 ( .A1(n4292), .A2(\SB2_4_9/Component_Function_3/NAND4_in[0] ), .A3(n4255), .A4(n6914), .ZN(\SB2_4_9/buf_output[3] ) );
  NAND3_X1 U13668 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0[6] ), .A3(
        \SB1_3_23/i1[9] ), .ZN(\SB1_3_23/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U13669 ( .A1(n6916), .A2(n5057), .Z(\MC_ARK_ARC_1_3/buf_output[183] ) );
  XOR2_X1 U13670 ( .A1(n7458), .A2(n7457), .Z(n6916) );
  NAND4_X2 U13671 ( .A1(\SB2_4_31/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_4_31/Component_Function_4/NAND4_in[0] ), .A3(n3689), .A4(n2469), 
        .ZN(\SB2_4_31/buf_output[4] ) );
  NAND3_X1 U13672 ( .A1(\SB4_20/i0[6] ), .A2(\SB4_20/i0[8] ), .A3(
        \SB4_20/i0[7] ), .ZN(n6917) );
  XOR2_X1 U13673 ( .A1(\RI5[2][155] ), .A2(\RI5[2][119] ), .Z(
        \MC_ARK_ARC_1_2/temp3[53] ) );
  NAND3_X2 U13674 ( .A1(\SB2_1_29/i0[10] ), .A2(\SB2_1_29/i0_0 ), .A3(
        \SB2_1_29/i0[6] ), .ZN(n6919) );
  NAND4_X2 U13675 ( .A1(\SB2_3_21/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_3_21/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_21/Component_Function_3/NAND4_in[0] ), .A4(n6920), .ZN(
        \SB2_3_21/buf_output[3] ) );
  XOR2_X1 U13676 ( .A1(n3089), .A2(n3090), .Z(\MC_ARK_ARC_1_4/buf_output[177] ) );
  NAND3_X2 U13677 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i1[9] ), .A3(
        \SB1_3_5/i0_4 ), .ZN(n6921) );
  XOR2_X1 U13678 ( .A1(n6922), .A2(n10), .Z(Ciphertext[18]) );
  NAND4_X2 U13679 ( .A1(\SB4_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_28/Component_Function_0/NAND4_in[1] ), .A3(n2412), .A4(n3122), 
        .ZN(n6922) );
  NAND3_X2 U13680 ( .A1(\SB2_3_15/i0[6] ), .A2(\SB2_3_15/i0_4 ), .A3(
        \SB2_3_15/i0[9] ), .ZN(n6923) );
  XOR2_X1 U13681 ( .A1(\RI5[0][103] ), .A2(\RI5[0][79] ), .Z(
        \MC_ARK_ARC_1_0/temp2[133] ) );
  NAND3_X1 U13682 ( .A1(\SB1_4_28/i0_4 ), .A2(\SB1_4_28/i1[9] ), .A3(
        \SB1_4_28/i1_5 ), .ZN(n2238) );
  NAND4_X2 U13683 ( .A1(\SB2_3_19/Component_Function_0/NAND4_in[2] ), .A2(
        n2232), .A3(\SB2_3_19/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_3_19/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_19/buf_output[0] ) );
  XOR2_X1 U13684 ( .A1(n4657), .A2(n7275), .Z(\MC_ARK_ARC_1_3/buf_output[20] )
         );
  INV_X2 U13685 ( .I(\SB1_3_9/buf_output[3] ), .ZN(\SB2_3_7/i0[8] ) );
  NAND4_X2 U13686 ( .A1(\SB1_3_9/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_9/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_3_9/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_3_9/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_9/buf_output[3] ) );
  XOR2_X1 U13687 ( .A1(\MC_ARK_ARC_1_2/temp4[134] ), .A2(
        \MC_ARK_ARC_1_2/temp3[134] ), .Z(\MC_ARK_ARC_1_2/temp6[134] ) );
  XOR2_X1 U13688 ( .A1(\MC_ARK_ARC_1_2/temp4[103] ), .A2(n2651), .Z(
        \MC_ARK_ARC_1_2/temp6[103] ) );
  NAND4_X2 U13689 ( .A1(\SB1_2_25/Component_Function_3/NAND4_in[1] ), .A2(
        n7237), .A3(\SB1_2_25/Component_Function_3/NAND4_in[0] ), .A4(n2203), 
        .ZN(\SB1_2_25/buf_output[3] ) );
  INV_X1 U13690 ( .I(\SB3_20/buf_output[1] ), .ZN(\SB4_16/i1_7 ) );
  XOR2_X1 U13691 ( .A1(n6925), .A2(n6924), .Z(\MC_ARK_ARC_1_1/buf_output[27] )
         );
  XOR2_X1 U13692 ( .A1(\MC_ARK_ARC_1_1/temp4[27] ), .A2(n2633), .Z(n6924) );
  XOR2_X1 U13693 ( .A1(\MC_ARK_ARC_1_1/temp3[27] ), .A2(
        \MC_ARK_ARC_1_1/temp1[27] ), .Z(n6925) );
  NAND3_X2 U13694 ( .A1(\SB3_26/i0[9] ), .A2(\SB3_26/i0_3 ), .A3(
        \SB3_26/i0[8] ), .ZN(n6926) );
  NAND3_X1 U13695 ( .A1(\SB2_2_19/i0_0 ), .A2(\SB2_2_19/i1_7 ), .A3(
        \SB2_2_19/i3[0] ), .ZN(\SB2_2_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U13696 ( .A1(\SB1_3_0/i0_3 ), .A2(\SB1_3_0/i0[7] ), .A3(
        \SB1_3_0/i0_0 ), .ZN(n6927) );
  XOR2_X1 U13697 ( .A1(n6928), .A2(n70), .Z(Ciphertext[155]) );
  NAND4_X2 U13698 ( .A1(\SB4_6/Component_Function_5/NAND4_in[3] ), .A2(n2742), 
        .A3(\SB4_6/Component_Function_5/NAND4_in[0] ), .A4(n7149), .ZN(n6928)
         );
  XOR2_X1 U13699 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[79] ), .A2(\RI5[2][103] ), 
        .Z(n6929) );
  NAND3_X1 U13700 ( .A1(\SB1_2_15/i0[10] ), .A2(\SB1_2_15/i0[6] ), .A3(
        \RI1[2][101] ), .ZN(\SB1_2_15/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U13701 ( .A1(\MC_ARK_ARC_1_3/temp6[7] ), .A2(
        \MC_ARK_ARC_1_3/temp5[7] ), .Z(\MC_ARK_ARC_1_3/buf_output[7] ) );
  NAND4_X2 U13702 ( .A1(\SB1_2_12/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_12/Component_Function_1/NAND4_in[1] ), .A3(n598), .A4(n6930), 
        .ZN(\SB1_2_12/buf_output[1] ) );
  NAND3_X2 U13703 ( .A1(\SB1_2_12/i1_5 ), .A2(\SB1_2_12/i0[9] ), .A3(
        \SB1_2_12/i0[6] ), .ZN(n6930) );
  NAND4_X2 U13704 ( .A1(\SB1_4_27/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_4_27/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_4_27/Component_Function_0/NAND4_in[2] ), .A4(n6931), .ZN(
        \SB1_4_27/buf_output[0] ) );
  NAND4_X2 U13705 ( .A1(\SB1_4_13/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_4_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_4_13/Component_Function_4/NAND4_in[0] ), .A4(n6933), .ZN(
        \SB1_4_13/buf_output[4] ) );
  NAND3_X2 U13706 ( .A1(\SB1_4_13/i0[10] ), .A2(\SB1_4_13/i0_3 ), .A3(
        \SB1_4_13/i0[9] ), .ZN(n6933) );
  XOR2_X1 U13707 ( .A1(\MC_ARK_ARC_1_2/temp2[169] ), .A2(n6934), .Z(n597) );
  XOR2_X1 U13708 ( .A1(\RI5[2][163] ), .A2(\RI5[2][169] ), .Z(n6934) );
  NAND3_X1 U13709 ( .A1(n1493), .A2(n3984), .A3(\SB4_17/i3[0] ), .ZN(n6935) );
  XOR2_X1 U13710 ( .A1(n6936), .A2(n76), .Z(Ciphertext[77]) );
  XOR2_X1 U13711 ( .A1(n2669), .A2(\MC_ARK_ARC_1_3/temp6[123] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[123] ) );
  XOR2_X1 U13712 ( .A1(\MC_ARK_ARC_1_3/temp2[123] ), .A2(
        \MC_ARK_ARC_1_3/temp1[123] ), .Z(n2669) );
  XOR2_X1 U13713 ( .A1(n6939), .A2(n201), .Z(Ciphertext[153]) );
  NAND4_X2 U13714 ( .A1(\SB2_3_24/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_24/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_3_24/Component_Function_1/NAND4_in[2] ), .A4(n6940), .ZN(
        \SB2_3_24/buf_output[1] ) );
  NAND4_X2 U13715 ( .A1(\SB2_2_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_2_20/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_2_20/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_20/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_2_20/buf_output[5] ) );
  XOR2_X1 U13716 ( .A1(\RI5[0][116] ), .A2(\RI5[0][110] ), .Z(
        \MC_ARK_ARC_1_0/temp1[116] ) );
  XOR2_X1 U13717 ( .A1(\MC_ARK_ARC_1_4/temp5[111] ), .A2(
        \MC_ARK_ARC_1_4/temp6[111] ), .Z(\MC_ARK_ARC_1_4/buf_output[111] ) );
  XOR2_X1 U13718 ( .A1(n4717), .A2(n6967), .Z(\MC_ARK_ARC_1_4/temp5[111] ) );
  NAND4_X2 U13719 ( .A1(n1623), .A2(\SB2_3_1/Component_Function_5/NAND4_in[0] ), .A3(n2115), .A4(n6942), .ZN(\SB2_3_1/buf_output[5] ) );
  NAND3_X2 U13720 ( .A1(\SB2_3_1/i0[10] ), .A2(\SB2_3_1/i0_0 ), .A3(
        \SB2_3_1/i0[6] ), .ZN(n6942) );
  NAND4_X2 U13721 ( .A1(n2665), .A2(\SB3_15/Component_Function_5/NAND4_in[2] ), 
        .A3(n3476), .A4(n6943), .ZN(\SB3_15/buf_output[5] ) );
  NAND3_X2 U13722 ( .A1(\SB2_1_10/i0[10] ), .A2(\SB2_1_10/i1_7 ), .A3(
        \SB2_1_10/i1[9] ), .ZN(n6944) );
  NAND3_X2 U13723 ( .A1(\SB1_1_12/i0_0 ), .A2(\SB1_1_12/i1_5 ), .A3(
        \SB1_1_12/i0_4 ), .ZN(\SB1_1_12/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U13724 ( .A1(\SB2_3_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_30/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_3_30/Component_Function_1/NAND4_in[0] ), .A4(n6945), .ZN(
        \SB2_3_30/buf_output[1] ) );
  NAND3_X1 U13725 ( .A1(\SB2_3_30/i0[9] ), .A2(\SB2_3_30/i0[6] ), .A3(
        \SB2_3_30/i1_5 ), .ZN(n6945) );
  XOR2_X1 U13726 ( .A1(\MC_ARK_ARC_1_0/temp1[109] ), .A2(n6946), .Z(n3354) );
  XOR2_X1 U13727 ( .A1(\RI5[0][19] ), .A2(\RI5[0][175] ), .Z(n6946) );
  NAND4_X2 U13728 ( .A1(\SB1_3_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_23/Component_Function_3/NAND4_in[1] ), .A3(n1109), .A4(n6947), 
        .ZN(\SB1_3_23/buf_output[3] ) );
  NAND4_X2 U13729 ( .A1(\SB1_4_17/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_4_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_17/Component_Function_1/NAND4_in[0] ), .A4(n6948), .ZN(
        \SB1_4_17/buf_output[1] ) );
  NAND3_X1 U13730 ( .A1(\SB1_4_7/i0[10] ), .A2(\SB1_4_7/i1[9] ), .A3(
        \SB1_4_7/i1_7 ), .ZN(n6949) );
  XOR2_X1 U13731 ( .A1(n6950), .A2(n71), .Z(Ciphertext[54]) );
  NAND4_X2 U13732 ( .A1(\SB4_22/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_22/Component_Function_0/NAND4_in[2] ), .A3(n1746), .A4(
        \SB4_22/Component_Function_0/NAND4_in[0] ), .ZN(n6950) );
  NAND3_X2 U13733 ( .A1(\SB2_1_11/i0_3 ), .A2(\SB2_1_11/i0[9] ), .A3(
        \SB2_1_11/i0[8] ), .ZN(n6951) );
  NAND4_X2 U13734 ( .A1(\SB1_2_13/Component_Function_5/NAND4_in[1] ), .A2(n784), .A3(\SB1_2_13/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_2_13/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_13/buf_output[5] ) );
  NAND3_X2 U13735 ( .A1(\SB1_4_13/i0_3 ), .A2(\SB1_4_13/i0_4 ), .A3(
        \SB1_4_13/i1[9] ), .ZN(n6953) );
  NAND4_X2 U13736 ( .A1(\SB3_13/Component_Function_4/NAND4_in[0] ), .A2(n5229), 
        .A3(\SB3_13/Component_Function_4/NAND4_in[1] ), .A4(n6954), .ZN(
        \SB3_13/buf_output[4] ) );
  XOR2_X1 U13737 ( .A1(n6955), .A2(n146), .Z(Ciphertext[145]) );
  NAND4_X2 U13738 ( .A1(\SB4_7/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_7/Component_Function_1/NAND4_in[3] ), .A3(n2535), .A4(
        \SB4_7/Component_Function_1/NAND4_in[0] ), .ZN(n6955) );
  NAND4_X2 U13739 ( .A1(\SB1_2_4/Component_Function_3/NAND4_in[1] ), .A2(n2564), .A3(\SB1_2_4/Component_Function_3/NAND4_in[0] ), .A4(n6956), .ZN(
        \SB1_2_4/buf_output[3] ) );
  NAND3_X2 U13740 ( .A1(\SB1_2_26/i0[10] ), .A2(\SB1_2_26/i1[9] ), .A3(
        \SB1_2_26/i1_7 ), .ZN(n6957) );
  NAND3_X2 U13741 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0_0 ), .A3(
        \SB1_3_31/i0_4 ), .ZN(\SB1_3_31/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U13742 ( .A1(\MC_ARK_ARC_1_1/temp5[143] ), .A2(
        \MC_ARK_ARC_1_1/temp6[143] ), .Z(\MC_ARK_ARC_1_1/buf_output[143] ) );
  NAND3_X1 U13743 ( .A1(\SB2_0_22/i0[7] ), .A2(\SB2_0_22/i0_3 ), .A3(
        \SB2_0_22/i0_0 ), .ZN(n3535) );
  NAND3_X2 U13744 ( .A1(\SB1_0_3/i0_4 ), .A2(\SB1_0_3/i1_7 ), .A3(
        \SB1_0_3/i0[8] ), .ZN(n6958) );
  XOR2_X1 U13745 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[79] ), .A2(\RI5[2][43] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[169] ) );
  XOR2_X1 U13746 ( .A1(\MC_ARK_ARC_1_3/temp5[26] ), .A2(n7045), .Z(
        \MC_ARK_ARC_1_3/buf_output[26] ) );
  NAND4_X2 U13747 ( .A1(n3652), .A2(
        \SB2_0_22/Component_Function_3/NAND4_in[1] ), .A3(n1617), .A4(
        \SB2_0_22/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_22/buf_output[3] ) );
  XOR2_X1 U13748 ( .A1(\RI5[0][69] ), .A2(\RI5[0][45] ), .Z(n4204) );
  NAND3_X2 U13749 ( .A1(\SB1_2_12/i1[9] ), .A2(\SB1_2_12/i1_7 ), .A3(
        \SB1_2_12/i0[10] ), .ZN(n7025) );
  NAND3_X1 U13750 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i0_0 ), .A3(\SB4_20/i0[7] ), .ZN(n6959) );
  NAND3_X1 U13751 ( .A1(\SB3_20/i0[10] ), .A2(\SB3_20/i1_5 ), .A3(
        \SB3_20/i1[9] ), .ZN(\SB3_20/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U13752 ( .A1(n4226), .A2(n4227), .Z(\MC_ARK_ARC_1_4/buf_output[65] )
         );
  XOR2_X1 U13753 ( .A1(\MC_ARK_ARC_1_4/temp2[65] ), .A2(
        \MC_ARK_ARC_1_4/temp4[65] ), .Z(n4226) );
  NAND2_X1 U13754 ( .A1(\SB1_4_31/Component_Function_4/NAND4_in[1] ), .A2(
        n7047), .ZN(n2347) );
  NAND3_X2 U13755 ( .A1(\SB1_4_30/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_4_30/Component_Function_5/NAND4_in[2] ), .A3(n6960), .ZN(
        \SB1_4_30/buf_output[5] ) );
  AOI21_X2 U13756 ( .A1(\SB1_4_30/i3[0] ), .A2(\SB1_4_30/i0_0 ), .B(n6961), 
        .ZN(n6960) );
  NAND4_X2 U13757 ( .A1(\SB2_1_5/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_5/Component_Function_5/NAND4_in[0] ), .A3(n758), .A4(n6962), 
        .ZN(\SB2_1_5/buf_output[5] ) );
  NAND3_X2 U13758 ( .A1(\SB2_1_5/i0[10] ), .A2(\SB2_1_5/i0_0 ), .A3(
        \SB2_1_5/i0[6] ), .ZN(n6962) );
  NAND3_X2 U13759 ( .A1(\SB1_1_22/i0[9] ), .A2(\SB1_1_22/i0[6] ), .A3(
        \SB1_1_22/i0_4 ), .ZN(n2531) );
  NAND3_X1 U13760 ( .A1(\SB2_4_20/i0_3 ), .A2(\SB2_4_20/i0_0 ), .A3(
        \SB2_4_20/i0_4 ), .ZN(n4900) );
  XOR2_X1 U13761 ( .A1(\MC_ARK_ARC_1_1/temp3[23] ), .A2(n6963), .Z(n3343) );
  XOR2_X1 U13762 ( .A1(\RI5[1][161] ), .A2(\RI5[1][185] ), .Z(n6963) );
  NAND2_X2 U13763 ( .A1(\SB1_4_25/i0_0 ), .A2(\SB1_4_25/i3[0] ), .ZN(
        \SB1_4_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U13764 ( .A1(\SB2_0_22/i0_3 ), .A2(\RI3[0][58] ), .A3(
        \SB2_0_22/i1[9] ), .ZN(\SB2_0_22/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U13765 ( .A1(\MC_ARK_ARC_1_4/temp3[186] ), .A2(
        \MC_ARK_ARC_1_4/temp4[186] ), .Z(n6964) );
  XOR2_X1 U13766 ( .A1(\MC_ARK_ARC_1_4/temp6[5] ), .A2(
        \MC_ARK_ARC_1_4/temp5[5] ), .Z(n3980) );
  XOR2_X1 U13767 ( .A1(n1683), .A2(n4367), .Z(\MC_ARK_ARC_1_4/temp5[5] ) );
  NAND3_X1 U13768 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i1[9] ), .A3(n237), 
        .ZN(n6965) );
  XOR2_X1 U13769 ( .A1(\RI5[0][38] ), .A2(\RI5[0][62] ), .Z(n5283) );
  NAND4_X2 U13770 ( .A1(\SB2_4_17/Component_Function_5/NAND4_in[2] ), .A2(
        n7214), .A3(n1016), .A4(n7109), .ZN(\SB2_4_17/buf_output[5] ) );
  XOR2_X1 U13771 ( .A1(\RI5[4][57] ), .A2(\RI5[4][111] ), .Z(n6967) );
  XOR2_X1 U13772 ( .A1(\RI5[1][57] ), .A2(\RI5[1][123] ), .Z(n6969) );
  NAND4_X2 U13773 ( .A1(\SB1_1_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_7/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_1_7/Component_Function_2/NAND4_in[1] ), .A4(n6971), .ZN(
        \SB1_1_7/buf_output[2] ) );
  NAND3_X2 U13774 ( .A1(\SB1_1_7/i0_0 ), .A2(\SB1_1_7/i1_5 ), .A3(
        \SB1_1_7/i0_4 ), .ZN(n6971) );
  NAND4_X2 U13775 ( .A1(\SB2_0_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_21/Component_Function_5/NAND4_in[3] ), .A3(n7230), .A4(
        \SB2_0_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_21/buf_output[5] ) );
  NAND3_X2 U13776 ( .A1(\SB2_4_17/i0_4 ), .A2(\SB2_4_17/i0_3 ), .A3(
        \SB2_4_17/i1[9] ), .ZN(\SB2_4_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U13777 ( .A1(\RI1[2][107] ), .A2(\SB1_2_14/i0_4 ), .A3(
        \SB1_2_14/i1[9] ), .ZN(n5156) );
  NAND4_X2 U13778 ( .A1(\SB2_1_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_2/NAND4_in[1] ), .A3(n5054), .A4(
        \SB2_1_18/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_1_18/buf_output[2] ) );
  NAND3_X2 U13779 ( .A1(\SB1_4_22/i0[6] ), .A2(\SB1_4_22/i0[10] ), .A3(
        \SB1_4_22/i0_0 ), .ZN(\SB1_4_22/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U13780 ( .A1(\SB1_0_11/i0[10] ), .A2(\SB1_0_11/i1[9] ), .A3(
        \SB1_0_11/i1_5 ), .ZN(n5158) );
  NAND3_X1 U13781 ( .A1(\SB2_3_11/i3[0] ), .A2(\SB2_3_11/i0[8] ), .A3(
        \SB2_3_11/i1_5 ), .ZN(\SB2_3_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U13782 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0[6] ), .A3(
        \SB1_3_23/i0[10] ), .ZN(\SB1_3_23/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U13783 ( .A1(n862), .A2(n6972), .Z(\MC_ARK_ARC_1_3/buf_output[45] )
         );
  XOR2_X1 U13784 ( .A1(\RI5[1][19] ), .A2(\RI5[1][175] ), .Z(n6977) );
  NAND4_X2 U13785 ( .A1(\SB3_0/Component_Function_3/NAND4_in[1] ), .A2(n7176), 
        .A3(n4096), .A4(n1475), .ZN(\SB3_0/buf_output[3] ) );
  NAND3_X2 U13786 ( .A1(\SB2_1_20/i0[7] ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0_0 ), .ZN(n4307) );
  NAND4_X2 U13787 ( .A1(\SB2_0_17/Component_Function_3/NAND4_in[0] ), .A2(
        n7067), .A3(n7247), .A4(\SB2_0_17/Component_Function_3/NAND4_in[3] ), 
        .ZN(\SB2_0_17/buf_output[3] ) );
  NAND4_X2 U13788 ( .A1(n4983), .A2(
        \SB2_1_22/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_22/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_1_22/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_22/buf_output[1] ) );
  XOR2_X1 U13789 ( .A1(\MC_ARK_ARC_1_0/temp6[186] ), .A2(n1653), .Z(
        \MC_ARK_ARC_1_0/buf_output[186] ) );
  NAND4_X2 U13790 ( .A1(\SB2_1_20/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_20/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_20/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_1_20/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_1_20/buf_output[2] ) );
  NAND3_X2 U13791 ( .A1(\SB1_4_24/i0[8] ), .A2(\SB1_4_24/i3[0] ), .A3(
        \SB1_4_24/i1_5 ), .ZN(n6973) );
  XOR2_X1 U13792 ( .A1(\MC_ARK_ARC_1_2/temp5[188] ), .A2(
        \MC_ARK_ARC_1_2/temp6[188] ), .Z(\MC_ARK_ARC_1_2/buf_output[188] ) );
  XOR2_X1 U13793 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[98] ), .A2(\RI5[2][62] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[188] ) );
  NAND4_X2 U13794 ( .A1(\SB1_0_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_2/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_2/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_2/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][179] ) );
  XOR2_X1 U13795 ( .A1(\RI5[1][96] ), .A2(\RI5[1][102] ), .Z(
        \MC_ARK_ARC_1_1/temp1[102] ) );
  XOR2_X1 U13796 ( .A1(\MC_ARK_ARC_1_0/temp3[191] ), .A2(n1399), .Z(n6980) );
  XOR2_X1 U13797 ( .A1(\RI5[1][24] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[0] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[54] ) );
  XOR2_X1 U13798 ( .A1(\RI5[0][180] ), .A2(\RI5[0][186] ), .Z(
        \MC_ARK_ARC_1_0/temp1[186] ) );
  NAND4_X2 U13799 ( .A1(\SB2_0_6/Component_Function_0/NAND4_in[1] ), .A2(n4497), .A3(n4498), .A4(n6974), .ZN(\SB2_0_6/buf_output[0] ) );
  NAND2_X1 U13800 ( .A1(\SB2_0_6/i0[9] ), .A2(\SB2_0_6/i0[10] ), .ZN(n6974) );
  XOR2_X1 U13801 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[60] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[84] ), .Z(\MC_ARK_ARC_1_2/temp2[114] )
         );
  NAND3_X2 U13802 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i0_4 ), .A3(
        \SB1_1_0/i1[9] ), .ZN(n6975) );
  NAND4_X2 U13803 ( .A1(\SB3_17/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_17/Component_Function_2/NAND4_in[2] ), .A3(n7207), .A4(n1787), 
        .ZN(\SB3_17/buf_output[2] ) );
  XOR2_X1 U13804 ( .A1(\MC_ARK_ARC_1_3/temp2[54] ), .A2(
        \MC_ARK_ARC_1_3/temp1[54] ), .Z(n2003) );
  XOR2_X1 U13805 ( .A1(n6977), .A2(\MC_ARK_ARC_1_1/temp4[109] ), .Z(n7563) );
  NAND3_X2 U13806 ( .A1(\SB1_3_14/i0[10] ), .A2(\SB1_3_14/i0_0 ), .A3(
        \SB1_3_14/i0[6] ), .ZN(\SB1_3_14/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U13807 ( .I(\SB1_3_17/buf_output[3] ), .ZN(\SB2_3_15/i0[8] ) );
  XOR2_X1 U13808 ( .A1(n6978), .A2(\MC_ARK_ARC_1_3/temp5[71] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[71] ) );
  XOR2_X1 U13809 ( .A1(\MC_ARK_ARC_1_3/temp4[71] ), .A2(n3546), .Z(n6978) );
  NAND3_X2 U13810 ( .A1(\SB1_0_3/i0_4 ), .A2(\SB1_0_3/i0_0 ), .A3(
        \SB1_0_3/i0_3 ), .ZN(n6981) );
  NAND4_X2 U13811 ( .A1(\SB2_0_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_1/Component_Function_5/NAND4_in[0] ), .A3(n7322), .A4(n6982), 
        .ZN(\SB2_0_1/buf_output[5] ) );
  NAND3_X2 U13812 ( .A1(\SB2_0_1/i0[10] ), .A2(\SB2_0_1/i0_0 ), .A3(
        \SB2_0_1/i0[6] ), .ZN(n6982) );
  NAND3_X2 U13813 ( .A1(\SB2_3_22/i0_0 ), .A2(\SB2_3_22/i0[9] ), .A3(
        \SB2_3_22/i0[8] ), .ZN(\SB2_3_22/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U13814 ( .A1(\SB2_3_23/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_23/Component_Function_0/NAND4_in[0] ), .A3(n4485), .A4(n6983), 
        .ZN(\SB2_3_23/buf_output[0] ) );
  XOR2_X1 U13815 ( .A1(\RI5[4][104] ), .A2(\RI5[4][140] ), .Z(n4869) );
  XOR2_X1 U13816 ( .A1(n6985), .A2(n6984), .Z(n4124) );
  XOR2_X1 U13817 ( .A1(\RI5[2][149] ), .A2(n115), .Z(n6984) );
  XOR2_X1 U13818 ( .A1(\RI5[2][191] ), .A2(\RI5[2][125] ), .Z(n6985) );
  NAND4_X2 U13819 ( .A1(\SB1_1_9/Component_Function_2/NAND4_in[1] ), .A2(n3116), .A3(\SB1_1_9/Component_Function_2/NAND4_in[2] ), .A4(n6986), .ZN(
        \RI3[1][152] ) );
  NAND4_X2 U13820 ( .A1(\SB2_1_24/Component_Function_0/NAND4_in[3] ), .A2(
        n1341), .A3(\SB2_1_24/Component_Function_0/NAND4_in[1] ), .A4(n6987), 
        .ZN(\SB2_1_24/buf_output[0] ) );
  XOR2_X1 U13821 ( .A1(\MC_ARK_ARC_1_0/temp6[135] ), .A2(n6988), .Z(
        \MC_ARK_ARC_1_0/buf_output[135] ) );
  NAND3_X2 U13822 ( .A1(\SB1_1_14/i0[10] ), .A2(\SB1_1_14/i0_3 ), .A3(
        \SB1_1_14/i0[9] ), .ZN(n7564) );
  XOR2_X1 U13823 ( .A1(\MC_ARK_ARC_1_0/temp1[185] ), .A2(n6989), .Z(
        \MC_ARK_ARC_1_0/temp5[185] ) );
  XOR2_X1 U13824 ( .A1(\RI5[0][155] ), .A2(\RI5[0][131] ), .Z(n6989) );
  NAND3_X2 U13825 ( .A1(n590), .A2(\SB2_1_0/i0_0 ), .A3(\SB2_1_0/i1_5 ), .ZN(
        \SB2_1_0/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U13826 ( .A1(\MC_ARK_ARC_1_2/temp5[189] ), .A2(n6991), .Z(
        \MC_ARK_ARC_1_2/buf_output[189] ) );
  XOR2_X1 U13827 ( .A1(\MC_ARK_ARC_1_2/temp3[189] ), .A2(
        \MC_ARK_ARC_1_2/temp4[189] ), .Z(n6991) );
  XOR2_X1 U13828 ( .A1(n4747), .A2(n6992), .Z(\MC_ARK_ARC_1_1/buf_output[43] )
         );
  XOR2_X1 U13829 ( .A1(\MC_ARK_ARC_1_1/temp3[43] ), .A2(
        \MC_ARK_ARC_1_1/temp4[43] ), .Z(n6992) );
  NAND3_X1 U13830 ( .A1(\SB1_2_9/i0_4 ), .A2(\SB1_2_9/i1_5 ), .A3(
        \SB1_2_9/i1[9] ), .ZN(\SB1_2_9/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U13831 ( .A1(\SB3_12/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_12/Component_Function_5/NAND4_in[2] ), .A3(
        \SB3_12/Component_Function_5/NAND4_in[0] ), .A4(n6993), .ZN(
        \SB3_12/buf_output[5] ) );
  NAND3_X2 U13832 ( .A1(\SB3_12/i0[6] ), .A2(\SB3_12/i0[9] ), .A3(
        \SB3_12/i0_4 ), .ZN(n6993) );
  INV_X1 U13833 ( .I(\SB3_22/buf_output[3] ), .ZN(\SB4_20/i0[8] ) );
  NAND4_X2 U13834 ( .A1(\SB3_22/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_22/Component_Function_3/NAND4_in[0] ), .A3(n694), .A4(
        \SB3_22/Component_Function_3/NAND4_in[2] ), .ZN(\SB3_22/buf_output[3] ) );
  NAND4_X2 U13835 ( .A1(\SB1_3_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_28/Component_Function_0/NAND4_in[3] ), .A4(n6994), .ZN(
        \SB1_3_28/buf_output[0] ) );
  XOR2_X1 U13836 ( .A1(n6995), .A2(n4452), .Z(n2623) );
  XOR2_X1 U13837 ( .A1(\RI5[0][101] ), .A2(\RI5[0][155] ), .Z(n6995) );
  XOR2_X1 U13838 ( .A1(\RI5[4][125] ), .A2(\RI5[4][161] ), .Z(
        \MC_ARK_ARC_1_4/temp3[59] ) );
  XOR2_X1 U13839 ( .A1(n6997), .A2(n203), .Z(Ciphertext[69]) );
  XOR2_X1 U13840 ( .A1(\RI5[0][65] ), .A2(\RI5[0][23] ), .Z(n3417) );
  XOR2_X1 U13841 ( .A1(\MC_ARK_ARC_1_2/temp6[174] ), .A2(n6998), .Z(
        \MC_ARK_ARC_1_2/buf_output[174] ) );
  XOR2_X1 U13842 ( .A1(n7584), .A2(\MC_ARK_ARC_1_2/temp1[174] ), .Z(n6998) );
  NAND3_X1 U13843 ( .A1(\SB1_2_9/i0_4 ), .A2(\SB1_2_9/i0[10] ), .A3(
        \SB1_2_9/i0_3 ), .ZN(\SB1_2_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U13844 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0_4 ), .A3(
        \SB1_0_25/i1[9] ), .ZN(\SB1_0_25/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U13845 ( .A1(n4305), .A2(n1061), .A3(n4023), .A4(
        \SB2_1_3/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_3/buf_output[5] ) );
  NAND3_X2 U13846 ( .A1(\SB2_4_15/i0_0 ), .A2(\SB2_4_15/i1_5 ), .A3(
        \SB2_4_15/i0_4 ), .ZN(n4940) );
  XOR2_X1 U13847 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[48] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[72] ), .Z(\MC_ARK_ARC_1_1/temp2[102] )
         );
  NAND4_X2 U13848 ( .A1(\SB2_3_9/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_9/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_3_9/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_3_9/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_9/buf_output[1] ) );
  XOR2_X1 U13849 ( .A1(\MC_ARK_ARC_1_4/temp6[154] ), .A2(
        \MC_ARK_ARC_1_4/temp5[154] ), .Z(\MC_ARK_ARC_1_4/buf_output[154] ) );
  NAND3_X2 U13850 ( .A1(\SB1_2_9/i0[10] ), .A2(\SB1_2_9/i1[9] ), .A3(
        \SB1_2_9/i1_7 ), .ZN(n6999) );
  XOR2_X1 U13851 ( .A1(n7000), .A2(\MC_ARK_ARC_1_1/temp4[15] ), .Z(
        \MC_ARK_ARC_1_1/temp6[15] ) );
  XOR2_X1 U13852 ( .A1(\RI5[1][81] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[117] ), 
        .Z(n7000) );
  NAND3_X2 U13853 ( .A1(\SB2_3_13/i0_3 ), .A2(\SB2_3_13/i0[6] ), .A3(
        \SB2_3_13/i1[9] ), .ZN(n5179) );
  NAND4_X2 U13854 ( .A1(n7141), .A2(
        \SB1_4_27/Component_Function_4/NAND4_in[2] ), .A3(n7093), .A4(n7001), 
        .ZN(\SB1_4_27/buf_output[4] ) );
  XOR2_X1 U13855 ( .A1(\RI5[0][56] ), .A2(\RI5[0][50] ), .Z(n7002) );
  NAND4_X2 U13856 ( .A1(\SB1_3_25/Component_Function_0/NAND4_in[2] ), .A2(n739), .A3(n7188), .A4(\SB1_3_25/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_3_25/buf_output[0] ) );
  INV_X2 U13857 ( .I(\RI3[0][167] ), .ZN(\SB2_0_4/i1_5 ) );
  XOR2_X1 U13858 ( .A1(\RI5[1][65] ), .A2(\RI5[1][101] ), .Z(
        \MC_ARK_ARC_1_1/temp3[191] ) );
  NAND4_X2 U13859 ( .A1(\SB2_2_28/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_2_28/Component_Function_3/NAND4_in[0] ), .A3(n5120), .A4(n922), 
        .ZN(\SB2_2_28/buf_output[3] ) );
  NAND3_X2 U13860 ( .A1(\SB1_4_6/i0[9] ), .A2(\SB1_4_6/i0[10] ), .A3(
        \RI1[4][155] ), .ZN(n7003) );
  XOR2_X1 U13861 ( .A1(\RI5[1][119] ), .A2(\RI5[1][167] ), .Z(n7005) );
  INV_X2 U13862 ( .I(\SB1_2_0/buf_output[2] ), .ZN(\SB2_2_29/i1[9] ) );
  NAND4_X2 U13863 ( .A1(\SB1_2_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_0/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_2_0/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_2_0/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_2_0/buf_output[2] ) );
  NAND3_X1 U13864 ( .A1(\SB4_21/i0[10] ), .A2(\SB3_24/buf_output[2] ), .A3(
        \SB4_21/i0[6] ), .ZN(\SB4_21/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U13865 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i0[9] ), .A3(\SB4_5/i0_3 ), 
        .ZN(n7006) );
  XOR2_X1 U13866 ( .A1(\MC_ARK_ARC_1_4/temp3[174] ), .A2(
        \MC_ARK_ARC_1_4/temp4[174] ), .Z(\MC_ARK_ARC_1_4/temp6[174] ) );
  XOR2_X1 U13867 ( .A1(n7007), .A2(n129), .Z(Ciphertext[159]) );
  NAND4_X2 U13868 ( .A1(n3649), .A2(\SB4_5/Component_Function_3/NAND4_in[3] ), 
        .A3(n1324), .A4(\SB4_5/Component_Function_3/NAND4_in[1] ), .ZN(n7007)
         );
  NAND2_X1 U13869 ( .A1(\SB3_8/i0_0 ), .A2(\SB3_8/i3[0] ), .ZN(n2067) );
  NAND3_X1 U13870 ( .A1(\SB1_2_5/i0[8] ), .A2(\SB1_2_5/i1_5 ), .A3(
        \SB1_2_5/i3[0] ), .ZN(\SB1_2_5/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U13871 ( .A1(\SB3_8/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_2/NAND4_in[0] ), .A4(n7008), .ZN(
        \SB3_8/buf_output[2] ) );
  NAND3_X1 U13872 ( .A1(\SB3_8/i0_0 ), .A2(\SB3_8/i0_4 ), .A3(\SB3_8/i1_5 ), 
        .ZN(n7008) );
  NAND4_X2 U13873 ( .A1(\SB1_4_0/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_4_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_4_0/Component_Function_4/NAND4_in[0] ), .A4(n7009), .ZN(
        \SB1_4_0/buf_output[4] ) );
  NAND3_X2 U13874 ( .A1(\SB1_4_0/i0_4 ), .A2(\SB1_4_0/i1_5 ), .A3(
        \SB1_4_0/i1[9] ), .ZN(n7009) );
  XOR2_X1 U13875 ( .A1(n3484), .A2(n7011), .Z(\MC_ARK_ARC_1_1/buf_output[159] ) );
  XOR2_X1 U13876 ( .A1(\MC_ARK_ARC_1_1/temp4[159] ), .A2(
        \MC_ARK_ARC_1_1/temp1[159] ), .Z(n7011) );
  NAND4_X2 U13877 ( .A1(\SB2_3_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_21/Component_Function_5/NAND4_in[1] ), .A3(n2848), .A4(n7012), 
        .ZN(\SB2_3_21/buf_output[5] ) );
  NAND3_X2 U13878 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0[10] ), .A3(
        \SB2_1_10/i0[9] ), .ZN(n2508) );
  XOR2_X1 U13879 ( .A1(n7015), .A2(n7014), .Z(n4043) );
  XOR2_X1 U13880 ( .A1(\RI5[1][159] ), .A2(n48), .Z(n7014) );
  XOR2_X1 U13881 ( .A1(\RI5[1][9] ), .A2(\RI5[1][165] ), .Z(n7015) );
  INV_X2 U13882 ( .I(\RI3[0][143] ), .ZN(\SB2_0_8/i1_5 ) );
  XOR2_X1 U13883 ( .A1(\RI5[1][183] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[189] ), .Z(\MC_ARK_ARC_1_1/temp1[189] ) );
  NAND3_X2 U13884 ( .A1(\SB2_4_21/i0_4 ), .A2(\SB2_4_21/i0_3 ), .A3(
        \SB2_4_21/i1[9] ), .ZN(\SB2_4_21/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U13885 ( .A1(\SB2_3_23/Component_Function_5/NAND4_in[2] ), .A2(
        n7128), .A3(n7017), .A4(\SB2_3_23/Component_Function_5/NAND4_in[0] ), 
        .ZN(\SB2_3_23/buf_output[5] ) );
  NAND3_X2 U13886 ( .A1(\SB2_3_25/i0_3 ), .A2(n5432), .A3(\SB2_3_25/i0[8] ), 
        .ZN(n7018) );
  NAND4_X2 U13887 ( .A1(\SB2_4_22/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_4_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_4_22/Component_Function_0/NAND4_in[0] ), .A4(n7019), .ZN(
        \SB2_4_22/buf_output[0] ) );
  XOR2_X1 U13888 ( .A1(\MC_ARK_ARC_1_4/temp1[90] ), .A2(
        \MC_ARK_ARC_1_4/temp2[90] ), .Z(\MC_ARK_ARC_1_4/temp5[90] ) );
  NAND3_X2 U13889 ( .A1(\SB2_4_30/i0[10] ), .A2(\SB2_4_30/i0_3 ), .A3(
        \SB2_4_30/i0[6] ), .ZN(n7099) );
  NAND4_X2 U13890 ( .A1(\SB1_2_0/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_2_0/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_0/Component_Function_4/NAND4_in[1] ), .A4(n7020), .ZN(
        \SB1_2_0/buf_output[4] ) );
  NAND3_X2 U13891 ( .A1(\SB2_2_30/i0[10] ), .A2(\SB2_2_30/i1_7 ), .A3(
        \SB2_2_30/i1[9] ), .ZN(n3923) );
  XOR2_X1 U13892 ( .A1(\RI5[3][191] ), .A2(\RI5[3][185] ), .Z(n7021) );
  XOR2_X1 U13893 ( .A1(\SB2_1_29/buf_output[0] ), .A2(\RI5[1][6] ), .Z(
        \MC_ARK_ARC_1_1/temp3[132] ) );
  XOR2_X1 U13894 ( .A1(n7022), .A2(\MC_ARK_ARC_1_2/temp6[51] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[51] ) );
  XOR2_X1 U13895 ( .A1(n7024), .A2(n7023), .Z(n2885) );
  XOR2_X1 U13896 ( .A1(\RI5[1][104] ), .A2(n427), .Z(n7023) );
  INV_X2 U13897 ( .I(\SB1_1_14/buf_output[3] ), .ZN(\SB2_1_12/i0[8] ) );
  NAND3_X1 U13898 ( .A1(\SB1_4_31/i0_3 ), .A2(\SB1_4_31/i1[9] ), .A3(
        \SB1_4_31/i0[6] ), .ZN(\SB1_4_31/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U13899 ( .A1(\MC_ARK_ARC_1_3/temp6[188] ), .A2(
        \MC_ARK_ARC_1_3/temp5[188] ), .Z(n3977) );
  XOR2_X1 U13900 ( .A1(\MC_ARK_ARC_1_3/temp2[103] ), .A2(
        \MC_ARK_ARC_1_3/temp1[103] ), .Z(n5073) );
  XOR2_X1 U13901 ( .A1(\MC_ARK_ARC_1_2/temp1[66] ), .A2(
        \MC_ARK_ARC_1_2/temp2[66] ), .Z(\MC_ARK_ARC_1_2/temp5[66] ) );
  NAND3_X1 U13902 ( .A1(\SB4_1/i0[10] ), .A2(n5442), .A3(\SB4_1/i1[9] ), .ZN(
        \SB4_1/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U13903 ( .I(\RI3[0][133] ), .ZN(\SB2_0_9/i1_7 ) );
  NAND4_X2 U13904 ( .A1(\SB1_0_13/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_13/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_0_13/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_0_13/Component_Function_1/NAND4_in[3] ), .ZN(\RI3[0][133] ) );
  NAND4_X2 U13905 ( .A1(\SB4_3/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_3/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_3/Component_Function_1/NAND4_in[3] ), .ZN(n7395) );
  NAND4_X2 U13906 ( .A1(\SB2_2_26/Component_Function_1/NAND4_in[0] ), .A2(
        n7414), .A3(\SB2_2_26/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_2_26/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_2_26/buf_output[1] ) );
  NAND4_X2 U13907 ( .A1(\SB1_2_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_30/Component_Function_5/NAND4_in[1] ), .A3(n7347), .A4(
        \SB1_2_30/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_30/buf_output[5] ) );
  XOR2_X1 U13908 ( .A1(\MC_ARK_ARC_1_1/temp6[18] ), .A2(n7027), .Z(
        \MC_ARK_ARC_1_1/buf_output[18] ) );
  XOR2_X1 U13909 ( .A1(\MC_ARK_ARC_1_1/temp1[18] ), .A2(
        \MC_ARK_ARC_1_1/temp2[18] ), .Z(n7027) );
  XOR2_X1 U13910 ( .A1(n4219), .A2(n7028), .Z(\MC_ARK_ARC_1_1/buf_output[188] ) );
  NAND3_X1 U13911 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i1_5 ), .A3(\SB4_5/i1[9] ), 
        .ZN(n7029) );
  NAND3_X1 U13912 ( .A1(\SB4_1/i0[9] ), .A2(\SB4_1/i0_3 ), .A3(\SB4_1/i0[8] ), 
        .ZN(n7030) );
  INV_X2 U13913 ( .I(\SB1_2_25/buf_output[3] ), .ZN(\SB2_2_23/i0[8] ) );
  XOR2_X1 U13914 ( .A1(n7031), .A2(\MC_ARK_ARC_1_3/temp6[25] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[25] ) );
  NAND4_X2 U13915 ( .A1(n7048), .A2(\SB2_3_8/Component_Function_0/NAND4_in[3] ), .A3(\SB2_3_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_8/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_8/buf_output[0] ) );
  XOR2_X1 U13916 ( .A1(n7032), .A2(\MC_ARK_ARC_1_2/temp4[48] ), .Z(
        \MC_ARK_ARC_1_2/temp6[48] ) );
  XOR2_X1 U13917 ( .A1(\RI5[2][114] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[150] ), .Z(n7032) );
  XOR2_X1 U13918 ( .A1(\RI5[3][63] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[69] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[69] ) );
  XOR2_X1 U13919 ( .A1(\MC_ARK_ARC_1_2/temp3[173] ), .A2(
        \MC_ARK_ARC_1_2/temp4[173] ), .Z(\MC_ARK_ARC_1_2/temp6[173] ) );
  XOR2_X1 U13920 ( .A1(n4921), .A2(n7033), .Z(\MC_ARK_ARC_1_3/buf_output[87] )
         );
  XOR2_X1 U13921 ( .A1(\MC_ARK_ARC_1_3/temp3[87] ), .A2(
        \MC_ARK_ARC_1_3/temp4[87] ), .Z(n7033) );
  NAND4_X2 U13922 ( .A1(n1012), .A2(
        \SB2_2_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_17/Component_Function_0/NAND4_in[0] ), .A4(n7034), .ZN(
        \SB2_2_17/buf_output[0] ) );
  NAND3_X1 U13923 ( .A1(\SB1_4_24/i0[10] ), .A2(\SB1_4_24/i1[9] ), .A3(
        \SB1_4_24/i1_5 ), .ZN(\SB1_4_24/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U13924 ( .A1(\SB4_21/Component_Function_3/NAND4_in[2] ), .A2(n4239), 
        .A3(\SB4_21/Component_Function_3/NAND4_in[1] ), .A4(n7035), .ZN(n7590)
         );
  NAND3_X1 U13925 ( .A1(\SB4_21/i0[6] ), .A2(\SB4_21/i0_3 ), .A3(n3998), .ZN(
        n7035) );
  INV_X2 U13926 ( .I(\SB1_1_23/buf_output[1] ), .ZN(\SB2_1_19/i1_7 ) );
  NAND4_X2 U13927 ( .A1(\SB1_1_23/Component_Function_1/NAND4_in[1] ), .A2(
        n2261), .A3(\SB1_1_23/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_1_23/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_1_23/buf_output[1] ) );
  NAND3_X1 U13928 ( .A1(\SB3_25/i0[8] ), .A2(\SB3_25/i0_3 ), .A3(\SB3_25/i1_7 ), .ZN(\SB3_25/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U13929 ( .A1(\SB2_3_10/i0[10] ), .A2(\SB2_3_10/i0_0 ), .A3(
        \SB2_3_10/i0[6] ), .ZN(n1291) );
  NAND3_X1 U13930 ( .A1(\SB4_22/i0_4 ), .A2(\SB4_22/i0_0 ), .A3(\SB4_22/i0_3 ), 
        .ZN(n7036) );
  XOR2_X1 U13931 ( .A1(n7039), .A2(n7038), .Z(n4700) );
  XOR2_X1 U13932 ( .A1(\RI5[2][152] ), .A2(\RI5[2][44] ), .Z(n7038) );
  XOR2_X1 U13933 ( .A1(\RI5[2][116] ), .A2(\RI5[2][50] ), .Z(n7039) );
  XOR2_X1 U13934 ( .A1(\RI5[1][89] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[125] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[23] ) );
  NAND3_X1 U13935 ( .A1(\SB1_3_10/i0[10] ), .A2(\SB1_3_10/i1[9] ), .A3(
        \SB1_3_10/i1_7 ), .ZN(n7040) );
  NAND4_X2 U13936 ( .A1(\SB1_3_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_5/NAND4_in[0] ), .A4(n7041), .ZN(
        \SB1_3_13/buf_output[5] ) );
  NAND3_X2 U13937 ( .A1(\SB1_3_13/i0[6] ), .A2(\SB1_3_13/i0_4 ), .A3(
        \SB1_3_13/i0[9] ), .ZN(n7041) );
  XOR2_X1 U13938 ( .A1(n7043), .A2(n7042), .Z(n5057) );
  XOR2_X1 U13939 ( .A1(\SB2_3_24/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_3/buf_keyinput[183] ), .Z(n7042) );
  NAND3_X2 U13940 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0[8] ), .A3(
        \SB2_2_14/i1_7 ), .ZN(\SB2_2_14/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U13941 ( .A1(n1045), .A2(\MC_ARK_ARC_1_3/temp4[26] ), .Z(n7045) );
  XOR2_X1 U13942 ( .A1(n7046), .A2(\MC_ARK_ARC_1_4/temp4[74] ), .Z(n7392) );
  XOR2_X1 U13943 ( .A1(\RI5[4][140] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[176] ), .Z(n7046) );
  NAND3_X1 U13944 ( .A1(\SB1_4_31/i0_0 ), .A2(\SB1_4_31/i0[9] ), .A3(
        \SB1_4_31/i0[8] ), .ZN(n7047) );
  NAND3_X1 U13945 ( .A1(\SB2_3_8/i0[6] ), .A2(\SB2_3_8/i0[7] ), .A3(
        \SB2_3_8/i0[8] ), .ZN(n7048) );
  XOR2_X1 U13946 ( .A1(n7049), .A2(\MC_ARK_ARC_1_1/temp4[152] ), .Z(
        \MC_ARK_ARC_1_1/temp6[152] ) );
  XOR2_X1 U13947 ( .A1(\RI5[1][26] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[62] ), 
        .Z(n7049) );
  XOR2_X1 U13948 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[181] ), .A2(\RI5[2][157] ), .Z(\MC_ARK_ARC_1_2/temp2[19] ) );
  NAND2_X2 U13949 ( .A1(n955), .A2(n954), .ZN(\RI5[2][157] ) );
  XOR2_X1 U13950 ( .A1(n7051), .A2(n159), .Z(Ciphertext[143]) );
  XOR2_X1 U13951 ( .A1(n7053), .A2(n7052), .Z(n1209) );
  XOR2_X1 U13952 ( .A1(\RI5[0][33] ), .A2(\RI5[0][57] ), .Z(n7052) );
  XOR2_X1 U13953 ( .A1(\RI5[0][9] ), .A2(\RI5[0][63] ), .Z(n7053) );
  NAND3_X1 U13954 ( .A1(\SB4_28/i0[6] ), .A2(\SB4_28/i0[7] ), .A3(
        \SB4_28/i0[8] ), .ZN(\SB4_28/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U13955 ( .A1(\SB1_4_10/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_4_10/Component_Function_4/NAND4_in[0] ), .A3(n7425), .A4(n7054), 
        .ZN(\SB1_4_10/buf_output[4] ) );
  NAND3_X2 U13956 ( .A1(\SB1_4_10/i0[10] ), .A2(\RI1[4][131] ), .A3(
        \SB1_4_10/i0[9] ), .ZN(n7054) );
  XOR2_X1 U13957 ( .A1(\RI5[4][157] ), .A2(\RI5[4][1] ), .Z(
        \MC_ARK_ARC_1_4/temp3[91] ) );
  XOR2_X1 U13958 ( .A1(\MC_ARK_ARC_1_0/temp6[35] ), .A2(n7055), .Z(
        \MC_ARK_ARC_1_0/buf_output[35] ) );
  XOR2_X1 U13959 ( .A1(n3445), .A2(n3446), .Z(n7055) );
  NAND4_X2 U13960 ( .A1(\SB2_4_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_4_26/Component_Function_3/NAND4_in[3] ), .A4(n7056), .ZN(
        \SB2_4_26/buf_output[3] ) );
  NAND3_X2 U13961 ( .A1(\SB2_4_26/i1[9] ), .A2(\SB2_4_26/i0[10] ), .A3(
        \SB2_4_26/i1_7 ), .ZN(n7056) );
  NAND4_X2 U13962 ( .A1(\SB1_1_6/Component_Function_2/NAND4_in[1] ), .A2(n4744), .A3(n2100), .A4(n7057), .ZN(\SB1_1_6/buf_output[2] ) );
  NAND3_X2 U13963 ( .A1(\SB1_1_6/i0[9] ), .A2(\SB1_1_6/i0_3 ), .A3(
        \SB1_1_6/i0[8] ), .ZN(n7057) );
  NAND4_X2 U13964 ( .A1(\SB1_1_12/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_12/Component_Function_2/NAND4_in[0] ), .A3(n7210), .A4(
        \SB1_1_12/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_1_12/buf_output[2] ) );
  AND2_X1 U13965 ( .A1(\SB1_4_21/Component_Function_4/NAND4_in[3] ), .A2(n7058), .Z(n5104) );
  NAND3_X1 U13966 ( .A1(\SB1_1_3/i1[9] ), .A2(\SB1_1_3/i0[10] ), .A3(
        \SB1_1_3/i1_5 ), .ZN(\SB1_1_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U13967 ( .A1(\SB3_0/i0[9] ), .A2(\SB3_0/i0[6] ), .A3(\SB3_0/i1_5 ), 
        .ZN(\SB3_0/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U13968 ( .A1(\SB1_4_19/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_4_19/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_4_19/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_4_19/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB1_4_19/buf_output[0] ) );
  NAND4_X2 U13969 ( .A1(\SB1_1_12/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_12/Component_Function_5/NAND4_in[2] ), .A3(n7330), .A4(
        \SB1_1_12/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_12/buf_output[5] ) );
  NAND2_X1 U13970 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i0[9] ), .ZN(
        \SB4_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 U13971 ( .A1(\SB2_0_18/i0[10] ), .A2(\SB2_0_18/i0[6] ), .A3(
        \SB2_0_18/i0_0 ), .ZN(\SB2_0_18/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U13972 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[3] ), .A2(\RI5[2][27] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[57] ) );
  XOR2_X1 U13973 ( .A1(\MC_ARK_ARC_1_0/temp5[153] ), .A2(n4202), .Z(
        \MC_ARK_ARC_1_0/buf_output[153] ) );
  NAND3_X1 U13974 ( .A1(\SB2_4_27/i0[10] ), .A2(\SB2_4_27/i0_3 ), .A3(
        \SB2_4_27/i0[6] ), .ZN(\SB2_4_27/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U13975 ( .A1(n3063), .A2(\MC_ARK_ARC_1_4/temp5[173] ), .Z(
        \RI1[5][173] ) );
  NAND3_X1 U13976 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i1_7 ), .A3(\SB4_16/i0[8] ), .ZN(\SB4_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U13977 ( .A1(\SB1_0_15/i0[9] ), .A2(\SB1_0_15/i0[8] ), .A3(
        \SB1_0_15/i0_0 ), .ZN(\SB1_0_15/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U13978 ( .A1(\MC_ARK_ARC_1_0/temp6[51] ), .A2(n3274), .Z(
        \MC_ARK_ARC_1_0/buf_output[51] ) );
  NAND4_X2 U13979 ( .A1(\SB1_0_2/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_2/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_0_2/Component_Function_4/NAND4_in[2] ), .ZN(\RI3[0][184] ) );
  NAND3_X2 U13980 ( .A1(\SB2_2_15/i0_0 ), .A2(\SB2_2_15/i0[9] ), .A3(
        \SB2_2_15/i0[8] ), .ZN(\SB2_2_15/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U13981 ( .A1(n2588), .A2(n2826), .A3(n798), .A4(
        \SB1_1_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_4/buf_output[5] ) );
  XOR2_X1 U13982 ( .A1(\MC_ARK_ARC_1_4/temp4[44] ), .A2(n7059), .Z(n4263) );
  XOR2_X1 U13983 ( .A1(\RI5[4][110] ), .A2(\RI5[4][146] ), .Z(n7059) );
  NAND4_X2 U13984 ( .A1(\SB1_2_7/Component_Function_5/NAND4_in[1] ), .A2(n3284), .A3(n7112), .A4(\SB1_2_7/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_7/buf_output[5] ) );
  NAND4_X2 U13985 ( .A1(\SB1_3_20/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_20/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_3_20/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_20/buf_output[0] ) );
  NAND4_X2 U13986 ( .A1(\SB1_2_12/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_12/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_12/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_2_12/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_12/buf_output[5] ) );
  XOR2_X1 U13987 ( .A1(\RI5[3][47] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[53] ) );
  XOR2_X1 U13988 ( .A1(n1277), .A2(\MC_ARK_ARC_1_1/temp6[88] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[88] ) );
  XOR2_X1 U13989 ( .A1(\RI5[1][129] ), .A2(\RI5[1][153] ), .Z(n4272) );
  NAND4_X2 U13990 ( .A1(\SB1_0_19/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_19/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_19/Component_Function_1/NAND4_in[3] ), .A4(n3644), .ZN(
        \RI3[0][97] ) );
  NAND3_X1 U13991 ( .A1(\SB4_23/i0_4 ), .A2(\SB4_23/i1_7 ), .A3(n3974), .ZN(
        \SB4_23/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U13992 ( .A1(n3447), .A2(\SB4_10/Component_Function_1/NAND4_in[3] ), 
        .A3(n1087), .A4(\SB4_10/Component_Function_1/NAND4_in[0] ), .ZN(n5370)
         );
  NAND4_X2 U13993 ( .A1(\SB1_2_7/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_2_7/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_7/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_7/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_2_7/buf_output[4] ) );
  NAND4_X2 U13994 ( .A1(\SB2_3_9/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_9/Component_Function_4/NAND4_in[1] ), .A3(n7265), .A4(n7061), 
        .ZN(\SB2_3_9/buf_output[4] ) );
  XOR2_X1 U13995 ( .A1(\RI5[0][21] ), .A2(\RI5[0][189] ), .Z(n7415) );
  XOR2_X1 U13996 ( .A1(\MC_ARK_ARC_1_4/temp4[105] ), .A2(n7062), .Z(n7383) );
  XOR2_X1 U13997 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[15] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[171] ), .Z(n7062) );
  INV_X2 U13998 ( .I(\RI3[0][8] ), .ZN(\SB2_0_30/i1[9] ) );
  NAND4_X2 U13999 ( .A1(n2181), .A2(\SB1_0_1/Component_Function_2/NAND4_in[1] ), .A3(\SB1_0_1/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_0_1/Component_Function_2/NAND4_in[2] ), .ZN(\RI3[0][8] ) );
  NAND3_X1 U14000 ( .A1(\SB4_6/i0_4 ), .A2(\SB4_6/i1_7 ), .A3(\SB4_6/i0[8] ), 
        .ZN(\SB4_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U14001 ( .A1(\SB2_3_30/i0_4 ), .A2(\SB2_3_30/i0_0 ), .A3(
        \SB2_3_30/i0_3 ), .ZN(n7063) );
  NAND3_X1 U14002 ( .A1(\SB1_4_25/i0_3 ), .A2(\SB1_4_25/i0_4 ), .A3(
        \SB1_4_25/i0[10] ), .ZN(\SB1_4_25/Component_Function_0/NAND4_in[2] )
         );
  NAND3_X2 U14003 ( .A1(\SB1_3_7/i0[10] ), .A2(\SB1_3_7/i1_7 ), .A3(
        \SB1_3_7/i1[9] ), .ZN(n2544) );
  NAND3_X1 U14004 ( .A1(\SB3_12/i1_5 ), .A2(\SB3_12/i3[0] ), .A3(
        \SB3_12/i0[8] ), .ZN(\SB3_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U14005 ( .A1(\SB4_19/i0_3 ), .A2(\SB4_19/i0[6] ), .A3(
        \SB4_19/i0[10] ), .ZN(n7065) );
  NAND3_X1 U14006 ( .A1(\SB4_7/i0_4 ), .A2(\SB4_7/i0_0 ), .A3(\SB4_7/i1_5 ), 
        .ZN(n7066) );
  NAND3_X2 U14007 ( .A1(\SB2_0_17/i0[10] ), .A2(\SB2_0_17/i1_7 ), .A3(
        \SB2_0_17/i1[9] ), .ZN(n7067) );
  NAND3_X1 U14008 ( .A1(\SB1_2_14/i3[0] ), .A2(\SB1_2_14/i0[8] ), .A3(
        \SB1_2_14/i1_5 ), .ZN(n7068) );
  NAND3_X1 U14009 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB2_3_19/i0[10] ), .A3(
        \SB1_3_20/buf_output[4] ), .ZN(
        \SB2_3_19/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U14010 ( .A1(\SB2_4_27/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_4_27/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_4_27/Component_Function_0/NAND4_in[0] ), .A4(n7069), .ZN(
        \SB2_4_27/buf_output[0] ) );
  XOR2_X1 U14011 ( .A1(\MC_ARK_ARC_1_0/temp2[29] ), .A2(n7070), .Z(n3942) );
  XOR2_X1 U14012 ( .A1(\RI5[0][95] ), .A2(\RI5[0][131] ), .Z(n7070) );
  NAND3_X1 U14013 ( .A1(\SB2_3_0/i0_0 ), .A2(\SB2_3_0/i0[9] ), .A3(
        \SB2_3_0/i0[8] ), .ZN(n7072) );
  NAND3_X2 U14014 ( .A1(\RI1[2][107] ), .A2(\SB1_2_14/i0[8] ), .A3(
        \SB1_2_14/i0[9] ), .ZN(n7201) );
  XOR2_X1 U14015 ( .A1(n7074), .A2(n7073), .Z(n3113) );
  XOR2_X1 U14016 ( .A1(\SB2_3_21/buf_output[2] ), .A2(n199), .Z(n7073) );
  XOR2_X1 U14017 ( .A1(\RI5[3][44] ), .A2(\RI5[3][14] ), .Z(n7074) );
  NAND4_X2 U14018 ( .A1(\SB2_1_16/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_16/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_1_16/Component_Function_4/NAND4_in[0] ), .A4(n7075), .ZN(
        \SB2_1_16/buf_output[4] ) );
  NAND3_X1 U14019 ( .A1(\SB2_1_16/i0[9] ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i0[10] ), .ZN(n7075) );
  NAND3_X2 U14020 ( .A1(\SB2_3_30/i0_4 ), .A2(\SB2_3_30/i0[9] ), .A3(
        \SB2_3_30/i0[6] ), .ZN(n7076) );
  NAND4_X2 U14021 ( .A1(\SB2_3_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_2/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_2/Component_Function_4/NAND4_in[1] ), .A4(n7077), .ZN(
        \SB2_3_2/buf_output[4] ) );
  NAND4_X2 U14022 ( .A1(\SB1_1_26/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_26/Component_Function_5/NAND4_in[1] ), .A3(n4683), .A4(
        \SB1_1_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_26/buf_output[5] ) );
  XOR2_X1 U14023 ( .A1(\RI5[3][22] ), .A2(n540), .Z(n7078) );
  NAND4_X2 U14024 ( .A1(\SB1_2_7/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_7/Component_Function_1/NAND4_in[0] ), .A4(n7080), .ZN(
        \SB1_2_7/buf_output[1] ) );
  NAND3_X2 U14025 ( .A1(\SB1_2_7/i1_5 ), .A2(\SB1_2_7/i0[6] ), .A3(
        \SB1_2_7/i0[9] ), .ZN(n7080) );
  XOR2_X1 U14026 ( .A1(n5316), .A2(\MC_ARK_ARC_1_4/temp4[111] ), .Z(
        \MC_ARK_ARC_1_4/temp6[111] ) );
  NAND4_X2 U14027 ( .A1(\SB1_4_16/Component_Function_3/NAND4_in[1] ), .A2(
        n4834), .A3(n3236), .A4(n7081), .ZN(\SB1_4_16/buf_output[3] ) );
  NAND3_X2 U14028 ( .A1(\SB2_0_15/i0[6] ), .A2(\SB2_0_15/i0[10] ), .A3(
        \SB1_0_18/buf_output[2] ), .ZN(n7082) );
  NAND3_X2 U14029 ( .A1(\SB2_0_15/i0[9] ), .A2(\SB2_0_15/i0[6] ), .A3(
        \RI3[0][100] ), .ZN(n7083) );
  XOR2_X1 U14030 ( .A1(n7084), .A2(n196), .Z(Ciphertext[62]) );
  NAND4_X2 U14031 ( .A1(\SB4_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB4_21/Component_Function_2/NAND4_in[2] ), .A3(
        \SB4_21/Component_Function_2/NAND4_in[3] ), .A4(
        \SB4_21/Component_Function_2/NAND4_in[1] ), .ZN(n7084) );
  XOR2_X1 U14032 ( .A1(n7085), .A2(n7086), .Z(\MC_ARK_ARC_1_4/buf_output[116] ) );
  XOR2_X1 U14033 ( .A1(n7175), .A2(n7087), .Z(\MC_ARK_ARC_1_4/buf_output[86] )
         );
  XOR2_X1 U14034 ( .A1(\MC_ARK_ARC_1_4/temp3[86] ), .A2(
        \MC_ARK_ARC_1_4/temp1[86] ), .Z(n7087) );
  NAND3_X1 U14035 ( .A1(\SB2_1_22/i0_0 ), .A2(\SB2_1_22/i0_3 ), .A3(
        \SB2_1_22/i0[7] ), .ZN(n1896) );
  NOR2_X2 U14036 ( .A1(n7089), .A2(n7088), .ZN(\SB2_1_22/i0[7] ) );
  NAND2_X2 U14037 ( .A1(\SB1_1_23/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_1_23/Component_Function_4/NAND4_in[2] ), .ZN(n7088) );
  NAND2_X2 U14038 ( .A1(\SB1_1_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_23/Component_Function_4/NAND4_in[1] ), .ZN(n7089) );
  NAND4_X2 U14039 ( .A1(\SB2_4_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_4_29/Component_Function_4/NAND4_in[3] ), .A3(n3726), .A4(n7090), 
        .ZN(\SB2_4_29/buf_output[4] ) );
  NAND3_X1 U14040 ( .A1(\SB2_4_29/i0[10] ), .A2(\SB2_4_29/i0_3 ), .A3(
        \SB2_4_29/i0[9] ), .ZN(n7090) );
  AND2_X1 U14041 ( .A1(n3475), .A2(\SB1_3_8/Component_Function_4/NAND4_in[3] ), 
        .Z(n7091) );
  NAND4_X2 U14042 ( .A1(\SB2_2_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_13/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_2_13/Component_Function_3/NAND4_in[1] ), .A4(n7092), .ZN(
        \SB2_2_13/buf_output[3] ) );
  NAND3_X1 U14043 ( .A1(\SB1_4_27/i0[9] ), .A2(\SB1_4_27/i0[8] ), .A3(
        \RI1[4][26] ), .ZN(n7093) );
  NAND4_X2 U14044 ( .A1(n3730), .A2(n757), .A3(n1928), .A4(
        \SB1_4_12/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_4_12/buf_output[4] ) );
  XOR2_X1 U14045 ( .A1(n4197), .A2(n7361), .Z(n4227) );
  XOR2_X1 U14046 ( .A1(\RI5[4][157] ), .A2(\RI5[4][133] ), .Z(
        \MC_ARK_ARC_1_4/temp2[187] ) );
  NAND4_X2 U14047 ( .A1(\SB1_4_28/Component_Function_0/NAND4_in[2] ), .A2(n655), .A3(\SB1_4_28/Component_Function_0/NAND4_in[0] ), .A4(n7095), .ZN(
        \SB1_4_28/buf_output[0] ) );
  NAND3_X1 U14048 ( .A1(\SB1_4_28/i0[6] ), .A2(\SB1_4_28/i0[8] ), .A3(
        \SB1_4_28/i0[7] ), .ZN(n7095) );
  NAND4_X2 U14049 ( .A1(\SB2_4_3/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_4_3/Component_Function_5/NAND4_in[0] ), .A3(
        \SB2_4_3/Component_Function_5/NAND4_in[1] ), .A4(n7096), .ZN(
        \SB2_4_3/buf_output[5] ) );
  NAND3_X2 U14050 ( .A1(\SB2_4_3/i0_4 ), .A2(\SB2_4_3/i0_3 ), .A3(
        \SB2_4_3/i1[9] ), .ZN(n7096) );
  NAND4_X2 U14051 ( .A1(\SB1_4_30/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_4_30/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_4_30/Component_Function_4/NAND4_in[1] ), .A4(n7097), .ZN(
        \SB1_4_30/buf_output[4] ) );
  NAND3_X1 U14052 ( .A1(\SB1_4_30/i0[9] ), .A2(\SB1_4_30/i0[10] ), .A3(
        \SB1_4_30/i0_3 ), .ZN(n7097) );
  XOR2_X1 U14053 ( .A1(\MC_ARK_ARC_1_3/temp6[150] ), .A2(n7098), .Z(
        \MC_ARK_ARC_1_3/buf_output[150] ) );
  XOR2_X1 U14054 ( .A1(n4371), .A2(\MC_ARK_ARC_1_3/temp2[150] ), .Z(n7098) );
  NAND4_X2 U14055 ( .A1(\SB2_4_30/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_4_30/Component_Function_2/NAND4_in[0] ), .A3(n4321), .A4(n7099), 
        .ZN(\SB2_4_30/buf_output[2] ) );
  NAND4_X2 U14056 ( .A1(\SB2_3_12/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_12/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_12/Component_Function_0/NAND4_in[0] ), .A4(n7100), .ZN(
        \SB2_3_12/buf_output[0] ) );
  NAND3_X2 U14057 ( .A1(\SB2_3_12/i0[6] ), .A2(n7586), .A3(\SB2_3_12/i0[8] ), 
        .ZN(n7100) );
  NAND4_X2 U14058 ( .A1(\SB1_1_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_19/Component_Function_5/NAND4_in[0] ), .A3(n5251), .A4(n7102), 
        .ZN(\SB1_1_19/buf_output[5] ) );
  NAND3_X2 U14059 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i1[9] ), .A3(
        \SB1_1_19/i0_4 ), .ZN(n7102) );
  XOR2_X1 U14060 ( .A1(n7104), .A2(n7103), .Z(\MC_ARK_ARC_1_4/temp5[89] ) );
  XOR2_X1 U14061 ( .A1(\RI5[4][59] ), .A2(\RI5[4][35] ), .Z(n7104) );
  INV_X2 U14062 ( .I(\MC_ARK_ARC_1_3/buf_output[17] ), .ZN(n7105) );
  XOR2_X1 U14063 ( .A1(n7107), .A2(n7106), .Z(\MC_ARK_ARC_1_2/buf_output[105] ) );
  XOR2_X1 U14064 ( .A1(\MC_ARK_ARC_1_2/temp1[105] ), .A2(
        \MC_ARK_ARC_1_2/temp3[105] ), .Z(n7106) );
  XOR2_X1 U14065 ( .A1(\MC_ARK_ARC_1_2/temp4[105] ), .A2(n4998), .Z(n7107) );
  NAND3_X2 U14066 ( .A1(\SB1_2_16/i0[10] ), .A2(\SB1_2_16/i0_0 ), .A3(
        \SB1_2_16/i0[6] ), .ZN(\SB1_2_16/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U14067 ( .A1(\SB3_3/i0_3 ), .A2(\SB3_3/i0[9] ), .A3(\SB3_3/i0[8] ), 
        .ZN(\SB3_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U14068 ( .A1(\SB2_4_0/i0[10] ), .A2(\SB2_4_0/i0_0 ), .A3(
        \SB2_4_0/i0[6] ), .ZN(n7108) );
  NAND2_X2 U14069 ( .A1(\SB2_4_17/i0_0 ), .A2(\SB2_4_17/i3[0] ), .ZN(n7109) );
  NAND3_X2 U14070 ( .A1(\SB1_3_16/i0[10] ), .A2(\SB1_3_16/i1[9] ), .A3(
        \SB1_3_16/i1_5 ), .ZN(n7110) );
  NAND3_X1 U14071 ( .A1(\SB1_4_4/i0[6] ), .A2(\SB1_4_4/i0[9] ), .A3(
        \SB1_4_4/i1_5 ), .ZN(n7111) );
  NAND3_X1 U14072 ( .A1(\SB1_2_26/i0_4 ), .A2(\SB1_2_26/i0_3 ), .A3(
        \SB1_2_26/i0[10] ), .ZN(\SB1_2_26/Component_Function_0/NAND4_in[2] )
         );
  NAND4_X2 U14073 ( .A1(\SB2_4_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_4_18/Component_Function_2/NAND4_in[2] ), .A3(n3201), .A4(n5315), 
        .ZN(\SB2_4_18/buf_output[2] ) );
  XOR2_X1 U14074 ( .A1(\MC_ARK_ARC_1_3/temp4[6] ), .A2(
        \MC_ARK_ARC_1_3/temp3[6] ), .Z(\MC_ARK_ARC_1_3/temp6[6] ) );
  NAND4_X2 U14075 ( .A1(\SB1_1_15/Component_Function_3/NAND4_in[1] ), .A2(
        n4752), .A3(\SB1_1_15/Component_Function_3/NAND4_in[2] ), .A4(n2877), 
        .ZN(\RI3[1][111] ) );
  XOR2_X1 U14076 ( .A1(n7113), .A2(n4155), .Z(\MC_ARK_ARC_1_3/temp6[15] ) );
  NAND4_X2 U14077 ( .A1(\SB2_4_11/Component_Function_3/NAND4_in[0] ), .A2(n904), .A3(\SB2_4_11/Component_Function_3/NAND4_in[3] ), .A4(n7114), .ZN(
        \SB2_4_11/buf_output[3] ) );
  XOR2_X1 U14078 ( .A1(\RI5[0][11] ), .A2(\RI5[0][167] ), .Z(
        \MC_ARK_ARC_1_0/temp3[101] ) );
  NAND4_X2 U14079 ( .A1(\SB2_1_13/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_13/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_13/Component_Function_1/NAND4_in[2] ), .A4(n7115), .ZN(
        \SB2_1_13/buf_output[1] ) );
  NAND3_X2 U14080 ( .A1(\SB2_1_13/i0_3 ), .A2(\SB2_1_13/i0[8] ), .A3(
        \SB2_1_13/i1_7 ), .ZN(n7115) );
  XOR2_X1 U14081 ( .A1(n7118), .A2(n7117), .Z(\MC_ARK_ARC_1_0/buf_output[170] ) );
  XOR2_X1 U14082 ( .A1(\MC_ARK_ARC_1_0/temp1[170] ), .A2(
        \MC_ARK_ARC_1_0/temp4[170] ), .Z(n7117) );
  XOR2_X1 U14083 ( .A1(\MC_ARK_ARC_1_0/temp2[170] ), .A2(
        \MC_ARK_ARC_1_0/temp3[170] ), .Z(n7118) );
  NAND3_X2 U14084 ( .A1(\SB1_4_20/i0_0 ), .A2(\SB1_4_20/i1_5 ), .A3(
        \SB1_4_20/i0_4 ), .ZN(n7119) );
  NAND3_X1 U14085 ( .A1(\SB4_9/i0[6] ), .A2(\SB4_9/i0[10] ), .A3(\SB4_9/i0_0 ), 
        .ZN(\SB4_9/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U14086 ( .I(\SB2_3_7/i0_4 ), .ZN(\SB2_3_7/i0[7] ) );
  XOR2_X1 U14087 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[188] ), .A2(\RI5[1][20] ), 
        .Z(n7122) );
  XOR2_X1 U14088 ( .A1(n3501), .A2(n7123), .Z(\MC_ARK_ARC_1_3/buf_output[135] ) );
  XOR2_X1 U14089 ( .A1(\MC_ARK_ARC_1_3/temp1[135] ), .A2(
        \MC_ARK_ARC_1_3/temp2[135] ), .Z(n7123) );
  NAND4_X2 U14090 ( .A1(\SB1_4_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_4_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_4_7/Component_Function_4/NAND4_in[2] ), .A4(n7124), .ZN(
        \SB1_4_7/buf_output[4] ) );
  NAND3_X1 U14091 ( .A1(\SB1_4_7/i1[9] ), .A2(\SB1_4_7/i1_5 ), .A3(
        \MC_ARK_ARC_1_3/buf_output[148] ), .ZN(n7124) );
  XOR2_X1 U14092 ( .A1(\MC_ARK_ARC_1_3/temp1[174] ), .A2(n7125), .Z(n3195) );
  XOR2_X1 U14093 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[144] ), .A2(\RI5[3][120] ), .Z(n7125) );
  NAND3_X1 U14094 ( .A1(\RI1[2][107] ), .A2(\SB1_2_14/i0[6] ), .A3(
        \SB1_2_14/i1[9] ), .ZN(n7126) );
  NAND4_X2 U14095 ( .A1(\SB1_4_29/Component_Function_4/NAND4_in[0] ), .A2(
        n4533), .A3(n7527), .A4(n7127), .ZN(\SB1_4_29/buf_output[4] ) );
  NAND3_X2 U14096 ( .A1(\SB2_3_17/i0[10] ), .A2(\SB2_3_17/i1_7 ), .A3(
        \SB2_3_17/i1[9] ), .ZN(n7216) );
  NAND3_X2 U14097 ( .A1(\SB2_4_4/i0_3 ), .A2(\SB2_4_4/i0[8] ), .A3(
        \SB2_4_4/i0[9] ), .ZN(\SB2_4_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U14098 ( .A1(\SB1_2_30/i0[10] ), .A2(\SB1_2_30/i1[9] ), .A3(
        \SB1_2_30/i1_7 ), .ZN(n7129) );
  XOR2_X1 U14099 ( .A1(\MC_ARK_ARC_1_3/temp5[33] ), .A2(n7130), .Z(
        \MC_ARK_ARC_1_3/buf_output[33] ) );
  NAND3_X2 U14100 ( .A1(\SB1_3_23/i0_0 ), .A2(\SB1_3_23/i1_5 ), .A3(
        \SB1_3_23/i0_4 ), .ZN(\SB1_3_23/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U14101 ( .A1(\SB4_28/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_28/Component_Function_4/NAND4_in[0] ), .A3(n1199), .A4(n2864), 
        .ZN(n7493) );
  NAND3_X2 U14102 ( .A1(\SB2_4_22/i0[10] ), .A2(\SB2_4_22/i1_7 ), .A3(
        \SB2_4_22/i1[9] ), .ZN(n7131) );
  XOR2_X1 U14103 ( .A1(\RI5[3][28] ), .A2(\RI5[3][52] ), .Z(
        \MC_ARK_ARC_1_3/temp2[82] ) );
  XOR2_X1 U14104 ( .A1(n7133), .A2(n37), .Z(Ciphertext[72]) );
  XOR2_X1 U14105 ( .A1(n2117), .A2(n1557), .Z(n7135) );
  NAND4_X2 U14106 ( .A1(\SB2_3_25/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_25/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_25/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_3_25/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB2_3_25/buf_output[4] ) );
  NAND4_X2 U14107 ( .A1(\SB4_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_19/Component_Function_3/NAND4_in[1] ), .A3(n3746), .A4(
        \SB4_19/Component_Function_3/NAND4_in[3] ), .ZN(n7476) );
  XOR2_X1 U14108 ( .A1(n7136), .A2(n7504), .Z(\MC_ARK_ARC_1_1/buf_output[117] ) );
  XOR2_X1 U14109 ( .A1(\MC_ARK_ARC_1_1/temp1[117] ), .A2(
        \MC_ARK_ARC_1_1/temp2[117] ), .Z(n7136) );
  XOR2_X1 U14110 ( .A1(\MC_ARK_ARC_1_1/temp5[123] ), .A2(n7137), .Z(
        \MC_ARK_ARC_1_1/buf_output[123] ) );
  XOR2_X1 U14111 ( .A1(\MC_ARK_ARC_1_1/temp3[123] ), .A2(
        \MC_ARK_ARC_1_1/temp4[123] ), .Z(n7137) );
  XOR2_X1 U14112 ( .A1(\MC_ARK_ARC_1_2/temp1[122] ), .A2(n7138), .Z(
        \MC_ARK_ARC_1_2/temp5[122] ) );
  XOR2_X1 U14113 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[92] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[68] ), .Z(n7138) );
  NAND2_X1 U14114 ( .A1(\SB1_0_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_15/Component_Function_4/NAND4_in[3] ), .ZN(n2610) );
  NAND3_X1 U14115 ( .A1(\SB2_0_15/i0_3 ), .A2(\SB2_0_15/i0[10] ), .A3(
        \RI3[0][100] ), .ZN(\SB2_0_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U14116 ( .A1(\SB1_1_21/i0[6] ), .A2(\SB1_1_21/i0[10] ), .A3(
        \SB1_1_21/i0_0 ), .ZN(n7139) );
  NAND3_X1 U14117 ( .A1(\SB1_4_27/i1[9] ), .A2(\SB1_4_27/i0_4 ), .A3(
        \SB1_4_27/i1_5 ), .ZN(n7141) );
  NAND3_X2 U14118 ( .A1(\SB2_4_13/i0[10] ), .A2(\SB2_4_13/i1[9] ), .A3(
        \SB2_4_13/i1_7 ), .ZN(n7581) );
  XOR2_X1 U14119 ( .A1(n3185), .A2(n3186), .Z(\MC_ARK_ARC_1_1/temp6[35] ) );
  XOR2_X1 U14120 ( .A1(\MC_ARK_ARC_1_0/temp5[45] ), .A2(
        \MC_ARK_ARC_1_0/temp6[45] ), .Z(\MC_ARK_ARC_1_0/buf_output[45] ) );
  NAND3_X2 U14121 ( .A1(\SB1_3_28/i0[10] ), .A2(\SB1_3_28/i1[9] ), .A3(
        \SB1_3_28/i1_5 ), .ZN(\SB1_3_28/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U14122 ( .A1(\MC_ARK_ARC_1_1/temp5[62] ), .A2(
        \MC_ARK_ARC_1_1/temp6[62] ), .Z(\MC_ARK_ARC_1_1/buf_output[62] ) );
  NAND4_X2 U14123 ( .A1(n980), .A2(\SB2_1_20/Component_Function_5/NAND4_in[1] ), .A3(n1490), .A4(\SB2_1_20/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_20/buf_output[5] ) );
  XOR2_X1 U14124 ( .A1(\RI5[0][111] ), .A2(\RI5[0][147] ), .Z(
        \MC_ARK_ARC_1_0/temp3[45] ) );
  XOR2_X1 U14125 ( .A1(n7142), .A2(n4625), .Z(\MC_ARK_ARC_1_0/buf_output[165] ) );
  XOR2_X1 U14126 ( .A1(\MC_ARK_ARC_1_0/temp2[165] ), .A2(
        \MC_ARK_ARC_1_0/temp3[165] ), .Z(n7142) );
  NAND4_X2 U14127 ( .A1(\SB1_1_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_24/Component_Function_4/NAND4_in[1] ), .A3(n2022), .A4(n7144), 
        .ZN(\SB1_1_24/buf_output[4] ) );
  NAND3_X1 U14128 ( .A1(\SB1_1_24/i0[10] ), .A2(\SB1_1_24/i0[9] ), .A3(
        \RI1[1][47] ), .ZN(n7144) );
  NAND3_X1 U14129 ( .A1(\SB3_11/i0[6] ), .A2(\SB3_11/i0[8] ), .A3(
        \SB3_11/i0[7] ), .ZN(\SB3_11/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U14130 ( .A1(n7147), .A2(n18), .Z(Ciphertext[151]) );
  XOR2_X1 U14131 ( .A1(n3295), .A2(n7148), .Z(\MC_ARK_ARC_1_0/buf_output[17] )
         );
  XOR2_X1 U14132 ( .A1(n7150), .A2(\MC_ARK_ARC_1_0/temp6[127] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[127] ) );
  XOR2_X1 U14133 ( .A1(\MC_ARK_ARC_1_0/temp1[127] ), .A2(
        \MC_ARK_ARC_1_0/temp2[127] ), .Z(n7150) );
  NAND3_X2 U14134 ( .A1(n5188), .A2(n7270), .A3(
        \SB2_0_15/Component_Function_1/NAND4_in[3] ), .ZN(\RI5[0][121] ) );
  XOR2_X1 U14135 ( .A1(n7152), .A2(n7289), .Z(\MC_ARK_ARC_1_3/buf_output[10] )
         );
  INV_X1 U14136 ( .I(\SB1_4_30/buf_output[5] ), .ZN(\SB2_4_30/i1_5 ) );
  NAND3_X2 U14137 ( .A1(\SB1_3_30/i0_4 ), .A2(\SB1_3_30/i0[10] ), .A3(
        \SB1_3_30/i0_3 ), .ZN(n7549) );
  XOR2_X1 U14138 ( .A1(n7153), .A2(\MC_ARK_ARC_1_4/temp6[181] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[181] ) );
  NAND4_X2 U14139 ( .A1(n7378), .A2(
        \SB2_3_12/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_3_12/Component_Function_5/NAND4_in[0] ), .A4(n7154), .ZN(
        \SB2_3_12/buf_output[5] ) );
  NAND3_X2 U14140 ( .A1(\SB2_3_12/i0[6] ), .A2(\SB2_3_12/i0[10] ), .A3(
        \SB2_3_12/i0_0 ), .ZN(n7154) );
  AND2_X1 U14141 ( .A1(\SB2_3_20/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_20/Component_Function_1/NAND4_in[0] ), .Z(n7155) );
  NAND2_X2 U14142 ( .A1(\SB1_3_20/i3[0] ), .A2(\SB1_3_20/i0_0 ), .ZN(
        \SB1_3_20/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 U14143 ( .A1(\SB1_0_15/Component_Function_5/NAND4_in[1] ), .A2(
        n7182), .A3(\SB1_0_15/Component_Function_5/NAND4_in[0] ), .A4(n7156), 
        .ZN(\RI3[0][101] ) );
  XOR2_X1 U14144 ( .A1(\MC_ARK_ARC_1_0/temp6[160] ), .A2(n7157), .Z(
        \MC_ARK_ARC_1_0/buf_output[160] ) );
  INV_X2 U14145 ( .I(\SB1_4_10/buf_output[2] ), .ZN(\SB2_4_7/i1[9] ) );
  XOR2_X1 U14146 ( .A1(\RI5[0][126] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[102] ), .Z(n7158) );
  INV_X2 U14147 ( .I(\RI3[0][176] ), .ZN(\SB2_0_2/i1[9] ) );
  NAND4_X2 U14148 ( .A1(\SB1_0_5/Component_Function_2/NAND4_in[0] ), .A2(n3938), .A3(n4574), .A4(\SB1_0_5/Component_Function_2/NAND4_in[2] ), .ZN(
        \RI3[0][176] ) );
  NAND4_X2 U14149 ( .A1(\SB1_1_7/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_7/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_7/Component_Function_3/NAND4_in[3] ), .A4(n7159), .ZN(
        \SB1_1_7/buf_output[3] ) );
  NAND3_X2 U14150 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i1[9] ), .A3(
        \SB1_1_7/i0[6] ), .ZN(n7159) );
  NAND3_X2 U14151 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i0[6] ), .A3(
        \SB2_1_0/i0_0 ), .ZN(\SB2_1_0/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U14152 ( .I(\SB1_3_16/buf_output[3] ), .ZN(\SB2_3_14/i0[8] ) );
  NOR2_X2 U14153 ( .A1(n2610), .A2(n7160), .ZN(n2822) );
  NAND3_X2 U14154 ( .A1(\SB2_0_11/i0[10] ), .A2(\SB2_0_11/i1_7 ), .A3(
        \SB2_0_11/i1[9] ), .ZN(n3623) );
  NAND4_X2 U14155 ( .A1(\SB2_1_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_29/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_29/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_1_29/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_1_29/buf_output[3] ) );
  INV_X2 U14156 ( .I(\SB1_1_0/buf_output[2] ), .ZN(\SB2_1_29/i1[9] ) );
  NAND3_X1 U14157 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0_0 ), .A3(
        \RI3[0][166] ), .ZN(n1669) );
  XOR2_X1 U14158 ( .A1(\MC_ARK_ARC_1_0/temp6[189] ), .A2(n7162), .Z(
        \MC_ARK_ARC_1_0/buf_output[189] ) );
  NAND4_X2 U14159 ( .A1(\SB1_2_9/Component_Function_1/NAND4_in[1] ), .A2(n3832), .A3(\SB1_2_9/Component_Function_1/NAND4_in[0] ), .A4(n7163), .ZN(
        \SB1_2_9/buf_output[1] ) );
  INV_X2 U14160 ( .I(\SB1_2_9/buf_output[3] ), .ZN(\SB2_2_7/i0[8] ) );
  XOR2_X1 U14161 ( .A1(\RI5[4][33] ), .A2(\RI5[4][189] ), .Z(
        \MC_ARK_ARC_1_4/temp3[123] ) );
  NAND4_X2 U14162 ( .A1(n3743), .A2(\SB2_3_0/Component_Function_5/NAND4_in[3] ), .A3(\SB2_3_0/Component_Function_5/NAND4_in[0] ), .A4(n7165), .ZN(
        \SB2_3_0/buf_output[5] ) );
  NAND3_X2 U14163 ( .A1(\SB2_3_0/i0_0 ), .A2(\SB2_3_0/i0[10] ), .A3(
        \SB2_3_0/i0[6] ), .ZN(n7165) );
  XOR2_X1 U14164 ( .A1(n7166), .A2(\MC_ARK_ARC_1_3/temp5[136] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[136] ) );
  XOR2_X1 U14165 ( .A1(\MC_ARK_ARC_1_3/temp3[136] ), .A2(
        \MC_ARK_ARC_1_3/temp4[136] ), .Z(n7166) );
  NAND3_X1 U14166 ( .A1(\SB1_1_6/i0[10] ), .A2(\SB1_1_6/i1[9] ), .A3(
        \SB1_1_6/i1_7 ), .ZN(\SB1_1_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U14167 ( .A1(\SB1_4_19/i0_4 ), .A2(\SB1_4_19/i1[9] ), .A3(
        \SB1_4_19/i1_5 ), .ZN(\SB1_4_19/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U14168 ( .A1(\SB2_0_0/i0[9] ), .A2(\RI3[0][189] ), .ZN(
        \SB2_0_0/Component_Function_0/NAND4_in[0] ) );
  XOR2_X1 U14169 ( .A1(\MC_ARK_ARC_1_3/temp5[46] ), .A2(
        \MC_ARK_ARC_1_3/temp6[46] ), .Z(\MC_ARK_ARC_1_3/buf_output[46] ) );
  XOR2_X1 U14170 ( .A1(\MC_ARK_ARC_1_0/temp1[4] ), .A2(
        \MC_ARK_ARC_1_0/temp2[4] ), .Z(n4545) );
  NAND3_X1 U14171 ( .A1(\SB1_1_27/i0_0 ), .A2(\SB1_1_27/i1_5 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[28] ), .ZN(n4554) );
  NAND4_X2 U14172 ( .A1(n4604), .A2(
        \SB1_2_23/Component_Function_5/NAND4_in[3] ), .A3(n3256), .A4(
        \SB1_2_23/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_23/buf_output[5] ) );
  XOR2_X1 U14173 ( .A1(\RI5[1][20] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[188] ), 
        .Z(n7168) );
  XOR2_X1 U14174 ( .A1(n7169), .A2(\MC_ARK_ARC_1_2/temp5[53] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[53] ) );
  XOR2_X1 U14175 ( .A1(\MC_ARK_ARC_1_2/temp3[53] ), .A2(
        \MC_ARK_ARC_1_2/temp4[53] ), .Z(n7169) );
  XOR2_X1 U14176 ( .A1(n7235), .A2(\MC_ARK_ARC_1_2/temp1[22] ), .Z(n7170) );
  XOR2_X1 U14177 ( .A1(n3154), .A2(n4654), .Z(\MC_ARK_ARC_1_1/buf_output[127] ) );
  XOR2_X1 U14178 ( .A1(\RI5[1][183] ), .A2(\RI5[1][159] ), .Z(n3664) );
  XOR2_X1 U14179 ( .A1(n7171), .A2(\MC_ARK_ARC_1_3/temp6[52] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[52] ) );
  XOR2_X1 U14180 ( .A1(\MC_ARK_ARC_1_3/temp1[52] ), .A2(
        \MC_ARK_ARC_1_3/temp2[52] ), .Z(n7171) );
  NAND3_X1 U14181 ( .A1(\SB4_1/i0_4 ), .A2(\SB4_1/i0_0 ), .A3(\SB4_1/i0_3 ), 
        .ZN(n7172) );
  NAND3_X1 U14182 ( .A1(\SB4_9/i0_3 ), .A2(n6272), .A3(\SB4_9/i0_0 ), .ZN(
        n7173) );
  NAND3_X1 U14183 ( .A1(\SB1_4_19/i0[6] ), .A2(\SB1_4_19/i0_3 ), .A3(
        \SB1_4_19/i1[9] ), .ZN(\SB1_4_19/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U14184 ( .A1(\MC_ARK_ARC_1_2/temp5[71] ), .A2(n7174), .Z(
        \MC_ARK_ARC_1_2/buf_output[71] ) );
  XOR2_X1 U14185 ( .A1(\MC_ARK_ARC_1_2/temp3[71] ), .A2(
        \MC_ARK_ARC_1_2/temp4[71] ), .Z(n7174) );
  XOR2_X1 U14186 ( .A1(\MC_ARK_ARC_1_4/temp2[86] ), .A2(
        \MC_ARK_ARC_1_4/temp4[86] ), .Z(n7175) );
  NAND4_X2 U14187 ( .A1(n4147), .A2(
        \SB1_4_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_4_25/Component_Function_3/NAND4_in[3] ), .A4(n7177), .ZN(
        \SB1_4_25/buf_output[3] ) );
  INV_X2 U14188 ( .I(\RI3[1][111] ), .ZN(\SB2_1_13/i0[8] ) );
  NAND3_X2 U14189 ( .A1(\SB1_4_7/i0_4 ), .A2(\SB1_4_7/i0_0 ), .A3(
        \SB1_4_7/i0_3 ), .ZN(\SB1_4_7/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U14190 ( .A1(n7178), .A2(\MC_ARK_ARC_1_2/temp2[104] ), .Z(n7363) );
  XOR2_X1 U14191 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[14] ), .A2(\RI5[2][170] ), 
        .Z(n7178) );
  XOR2_X1 U14192 ( .A1(n924), .A2(n7179), .Z(n2667) );
  XOR2_X1 U14193 ( .A1(\RI5[3][137] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[143] ), .Z(n7179) );
  NAND3_X2 U14194 ( .A1(\SB1_0_15/i0[9] ), .A2(\SB1_0_15/i0[6] ), .A3(
        \SB1_0_15/i0_4 ), .ZN(n7182) );
  XOR2_X1 U14195 ( .A1(\MC_ARK_ARC_1_4/temp4[168] ), .A2(n7183), .Z(
        \MC_ARK_ARC_1_4/temp6[168] ) );
  XOR2_X1 U14196 ( .A1(\RI5[4][42] ), .A2(\RI5[4][78] ), .Z(n7183) );
  XOR2_X1 U14197 ( .A1(n7299), .A2(\MC_ARK_ARC_1_2/temp2[160] ), .Z(
        \MC_ARK_ARC_1_2/temp5[160] ) );
  NAND3_X1 U14198 ( .A1(\SB3_3/i0[9] ), .A2(\SB3_3/i1_5 ), .A3(\SB3_3/i0[6] ), 
        .ZN(\SB3_3/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U14199 ( .A1(\SB2_1_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_9/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_1_9/Component_Function_2/NAND4_in[2] ), .A4(n7184), .ZN(
        \SB2_1_9/buf_output[2] ) );
  NAND3_X2 U14200 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0[10] ), .A3(
        \SB2_1_9/i0[6] ), .ZN(n7184) );
  XOR2_X1 U14201 ( .A1(\MC_ARK_ARC_1_4/temp4[98] ), .A2(n7186), .Z(
        \MC_ARK_ARC_1_4/temp6[98] ) );
  XOR2_X1 U14202 ( .A1(\SB2_4_1/buf_output[2] ), .A2(\RI5[4][164] ), .Z(n7186)
         );
  NAND3_X2 U14203 ( .A1(\SB2_0_15/i0[9] ), .A2(\SB2_0_15/i0_3 ), .A3(
        \SB2_0_15/i0[8] ), .ZN(n7187) );
  NAND3_X1 U14204 ( .A1(\SB2_2_13/i0[10] ), .A2(\SB2_2_13/i0_3 ), .A3(
        \SB2_2_13/i0_4 ), .ZN(\SB2_2_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U14205 ( .A1(\SB1_2_29/i0[10] ), .A2(\SB1_2_29/i1_7 ), .A3(
        \SB1_2_29/i1[9] ), .ZN(\SB1_2_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U14206 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i1[9] ), .A3(
        \SB4_24/i0[6] ), .ZN(n7189) );
  NAND4_X2 U14207 ( .A1(\SB2_1_26/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_26/Component_Function_2/NAND4_in[2] ), .A4(n7190), .ZN(
        \SB2_1_26/buf_output[2] ) );
  NAND3_X2 U14208 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0_0 ), .A3(
        \SB1_0_2/i0_4 ), .ZN(\SB1_0_2/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U14209 ( .A1(n7191), .A2(n214), .Z(Ciphertext[67]) );
  NAND4_X2 U14210 ( .A1(\SB4_20/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_20/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_20/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_20/Component_Function_1/NAND4_in[0] ), .ZN(n7191) );
  NAND3_X1 U14211 ( .A1(\SB2_0_1/i0_4 ), .A2(\SB2_0_1/i0[10] ), .A3(
        \SB2_0_1/i0_3 ), .ZN(n7192) );
  NAND3_X2 U14212 ( .A1(\SB1_1_22/i1_5 ), .A2(\SB1_1_22/i0[10] ), .A3(
        \SB1_1_22/i1[9] ), .ZN(n7578) );
  NAND4_X2 U14213 ( .A1(\SB2_2_10/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_10/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_2_10/Component_Function_1/NAND4_in[2] ), .A4(n7194), .ZN(
        \SB2_2_10/buf_output[1] ) );
  NAND3_X2 U14214 ( .A1(\SB2_2_10/i0_4 ), .A2(\SB2_2_10/i1_7 ), .A3(
        \SB2_2_10/i0[8] ), .ZN(n7194) );
  XOR2_X1 U14215 ( .A1(\MC_ARK_ARC_1_0/temp1[57] ), .A2(n7195), .Z(n7413) );
  XOR2_X1 U14216 ( .A1(\SB2_0_1/buf_output[3] ), .A2(\RI5[0][27] ), .Z(n7195)
         );
  XOR2_X1 U14217 ( .A1(n7197), .A2(n7196), .Z(\MC_ARK_ARC_1_1/buf_output[187] ) );
  XOR2_X1 U14218 ( .A1(\MC_ARK_ARC_1_1/temp1[187] ), .A2(
        \MC_ARK_ARC_1_1/temp3[187] ), .Z(n7196) );
  XOR2_X1 U14219 ( .A1(\MC_ARK_ARC_1_1/temp4[187] ), .A2(
        \MC_ARK_ARC_1_1/temp2[187] ), .Z(n7197) );
  NAND3_X1 U14220 ( .A1(\SB2_3_5/i0_4 ), .A2(\SB2_3_5/i1_7 ), .A3(
        \SB2_3_5/i0[8] ), .ZN(\SB2_3_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U14221 ( .A1(\SB2_2_0/i0_0 ), .A2(\SB2_2_0/i3[0] ), .A3(
        \SB2_2_0/i1_7 ), .ZN(\SB2_2_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U14222 ( .A1(\SB1_3_26/i0_4 ), .A2(\SB1_3_26/i1_7 ), .A3(
        \SB1_3_26/i0[8] ), .ZN(\SB1_3_26/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U14223 ( .A1(\SB2_4_28/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_4_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_4_28/Component_Function_4/NAND4_in[2] ), .A4(n7198), .ZN(
        \SB2_4_28/buf_output[4] ) );
  NAND3_X1 U14224 ( .A1(\SB2_3_25/i0_3 ), .A2(\SB2_3_25/i0_0 ), .A3(
        \SB2_3_25/i0_4 ), .ZN(\SB2_3_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U14225 ( .A1(\SB1_2_1/i0[9] ), .A2(\SB1_2_1/i0[8] ), .A3(
        \SB1_2_1/i0_0 ), .ZN(n7199) );
  NAND3_X2 U14226 ( .A1(\SB2_4_30/i0_0 ), .A2(\SB2_4_30/i0_3 ), .A3(
        \SB1_4_31/buf_output[4] ), .ZN(n2683) );
  NAND3_X2 U14227 ( .A1(\SB1_2_14/i0_0 ), .A2(\SB1_2_14/i0_4 ), .A3(
        \SB1_2_14/i1_5 ), .ZN(n7202) );
  XOR2_X1 U14228 ( .A1(\RI5[2][123] ), .A2(\RI5[2][93] ), .Z(n3413) );
  XOR2_X1 U14229 ( .A1(\RI5[3][17] ), .A2(\RI5[3][11] ), .Z(n3361) );
  INV_X2 U14230 ( .I(\SB1_0_19/buf_output[2] ), .ZN(\SB2_0_16/i1[9] ) );
  NAND4_X2 U14231 ( .A1(\SB1_0_19/Component_Function_2/NAND4_in[0] ), .A2(
        n3585), .A3(\SB1_0_19/Component_Function_2/NAND4_in[2] ), .A4(n4146), 
        .ZN(\SB1_0_19/buf_output[2] ) );
  XOR2_X1 U14232 ( .A1(\MC_ARK_ARC_1_1/temp6[99] ), .A2(
        \MC_ARK_ARC_1_1/temp5[99] ), .Z(n1509) );
  XOR2_X1 U14233 ( .A1(\MC_ARK_ARC_1_1/temp1[99] ), .A2(
        \MC_ARK_ARC_1_1/temp2[99] ), .Z(\MC_ARK_ARC_1_1/temp5[99] ) );
  NAND4_X2 U14234 ( .A1(\SB1_2_7/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_2_7/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_7/Component_Function_3/NAND4_in[0] ), .A4(n7284), .ZN(
        \SB1_2_7/buf_output[3] ) );
  XOR2_X1 U14235 ( .A1(\MC_ARK_ARC_1_2/temp5[110] ), .A2(
        \MC_ARK_ARC_1_2/temp6[110] ), .Z(\MC_ARK_ARC_1_2/buf_output[110] ) );
  NAND4_X2 U14236 ( .A1(\SB1_4_8/Component_Function_2/NAND4_in[1] ), .A2(n2393), .A3(\SB1_4_8/Component_Function_2/NAND4_in[3] ), .A4(n7204), .ZN(
        \SB1_4_8/buf_output[2] ) );
  XOR2_X1 U14237 ( .A1(\RI5[3][113] ), .A2(\RI5[3][89] ), .Z(n924) );
  XOR2_X1 U14238 ( .A1(\RI5[0][105] ), .A2(\RI5[0][111] ), .Z(
        \MC_ARK_ARC_1_0/temp1[111] ) );
  XOR2_X1 U14239 ( .A1(n3506), .A2(\MC_ARK_ARC_1_1/temp6[158] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[158] ) );
  XOR2_X1 U14240 ( .A1(\MC_ARK_ARC_1_2/temp6[169] ), .A2(n597), .Z(
        \MC_ARK_ARC_1_2/buf_output[169] ) );
  XOR2_X1 U14241 ( .A1(\RI5[3][59] ), .A2(\RI5[3][89] ), .Z(n5244) );
  XOR2_X1 U14242 ( .A1(n7205), .A2(n130), .Z(Ciphertext[104]) );
  NAND4_X2 U14243 ( .A1(\SB4_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_14/Component_Function_2/NAND4_in[0] ), .A3(n7560), .A4(n4238), 
        .ZN(n7205) );
  XOR2_X1 U14244 ( .A1(\MC_ARK_ARC_1_4/temp6[88] ), .A2(n7206), .Z(
        \MC_ARK_ARC_1_4/buf_output[88] ) );
  XOR2_X1 U14245 ( .A1(\MC_ARK_ARC_1_4/temp2[88] ), .A2(n4424), .Z(n7206) );
  XOR2_X1 U14246 ( .A1(\RI5[3][134] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[158] ), .Z(\MC_ARK_ARC_1_3/temp2[188] ) );
  NAND3_X2 U14247 ( .A1(\SB3_17/i0_4 ), .A2(\SB3_17/i0_0 ), .A3(\SB3_17/i1_5 ), 
        .ZN(n7207) );
  XOR2_X1 U14248 ( .A1(\MC_ARK_ARC_1_3/temp5[187] ), .A2(n7209), .Z(
        \MC_ARK_ARC_1_3/buf_output[187] ) );
  XOR2_X1 U14249 ( .A1(\MC_ARK_ARC_1_3/temp3[187] ), .A2(
        \MC_ARK_ARC_1_3/temp4[187] ), .Z(n7209) );
  NAND3_X2 U14250 ( .A1(\SB1_1_12/i0[10] ), .A2(\SB1_1_12/i0_3 ), .A3(
        \SB1_1_12/i0[6] ), .ZN(n7210) );
  XOR2_X1 U14251 ( .A1(\RI5[1][60] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[36] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[90] ) );
  NAND4_X2 U14252 ( .A1(\SB1_1_17/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_1_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_17/Component_Function_1/NAND4_in[0] ), .A4(n7211), .ZN(
        \SB1_1_17/buf_output[1] ) );
  NAND3_X2 U14253 ( .A1(\SB1_1_17/i0[9] ), .A2(\SB1_1_17/i0[6] ), .A3(
        \SB1_1_17/i1_5 ), .ZN(n7211) );
  NAND4_X2 U14254 ( .A1(\SB1_2_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_16/Component_Function_5/NAND4_in[0] ), .A4(n7212), .ZN(
        \SB1_2_16/buf_output[5] ) );
  NAND4_X2 U14255 ( .A1(\SB2_2_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_8/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_8/Component_Function_5/NAND4_in[0] ), .A4(n7213), .ZN(
        \SB2_2_8/buf_output[5] ) );
  NAND3_X2 U14256 ( .A1(\SB2_2_8/i0[6] ), .A2(\SB2_2_8/i0_4 ), .A3(
        \SB2_2_8/i0[9] ), .ZN(n7213) );
  XOR2_X1 U14257 ( .A1(\RI5[3][67] ), .A2(\RI5[3][91] ), .Z(
        \MC_ARK_ARC_1_3/temp2[121] ) );
  NAND3_X2 U14258 ( .A1(\SB2_4_17/i0[10] ), .A2(\SB2_4_17/i0_0 ), .A3(
        \SB2_4_17/i0[6] ), .ZN(n7214) );
  NAND4_X2 U14259 ( .A1(\SB2_2_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_23/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_2_23/Component_Function_3/NAND4_in[1] ), .A4(n7217), .ZN(
        \SB2_2_23/buf_output[3] ) );
  NAND3_X2 U14260 ( .A1(\SB2_2_23/i0[10] ), .A2(\SB2_2_23/i1_7 ), .A3(
        \SB2_2_23/i1[9] ), .ZN(n7217) );
  XOR2_X1 U14261 ( .A1(n7218), .A2(n219), .Z(Ciphertext[28]) );
  NAND4_X2 U14262 ( .A1(n2217), .A2(n7580), .A3(n1903), .A4(
        \SB4_27/Component_Function_4/NAND4_in[1] ), .ZN(n7218) );
  NAND3_X2 U14263 ( .A1(\SB2_4_22/i0[10] ), .A2(\SB2_4_22/i0_3 ), .A3(
        \SB2_4_22/i0[6] ), .ZN(n7219) );
  INV_X2 U14264 ( .I(\SB1_3_24/buf_output[3] ), .ZN(\SB2_3_22/i0[8] ) );
  NAND4_X2 U14265 ( .A1(\SB1_3_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_3_24/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_3_24/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_24/buf_output[3] ) );
  NAND4_X2 U14266 ( .A1(\SB2_2_21/Component_Function_2/NAND4_in[0] ), .A2(
        n1052), .A3(n7223), .A4(n7220), .ZN(\SB2_2_21/buf_output[2] ) );
  NAND4_X2 U14267 ( .A1(\SB2_4_19/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_4_19/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_4_19/Component_Function_3/NAND4_in[1] ), .A4(n7221), .ZN(
        \SB2_4_19/buf_output[3] ) );
  XOR2_X1 U14268 ( .A1(\MC_ARK_ARC_1_0/temp5[146] ), .A2(n7222), .Z(
        \MC_ARK_ARC_1_0/buf_output[146] ) );
  XOR2_X1 U14269 ( .A1(n7327), .A2(\MC_ARK_ARC_1_0/temp4[146] ), .Z(n7222) );
  BUF_X2 U14270 ( .I(n3104), .Z(n7225) );
  NAND4_X2 U14271 ( .A1(\SB1_1_15/Component_Function_5/NAND4_in[1] ), .A2(
        n2903), .A3(\SB1_1_15/Component_Function_5/NAND4_in[0] ), .A4(n7226), 
        .ZN(\SB1_1_15/buf_output[5] ) );
  NAND3_X2 U14272 ( .A1(\SB1_1_15/i0[6] ), .A2(\SB1_1_15/i0[9] ), .A3(
        \SB1_1_15/i0_4 ), .ZN(n7226) );
  NAND4_X2 U14273 ( .A1(\SB1_2_13/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_13/Component_Function_3/NAND4_in[0] ), .A3(n1573), .A4(
        \SB1_2_13/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_13/buf_output[3] ) );
  NAND3_X1 U14274 ( .A1(\SB2_2_18/i0_3 ), .A2(\SB2_2_18/i0[8] ), .A3(
        \SB2_2_18/i1_7 ), .ZN(\SB2_2_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U14275 ( .A1(\SB2_3_1/i0_4 ), .A2(\SB2_3_1/i1_5 ), .A3(
        \SB2_3_1/i1[9] ), .ZN(n7227) );
  NAND4_X2 U14276 ( .A1(\SB1_1_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_6/Component_Function_3/NAND4_in[2] ), .A3(n1883), .A4(n7228), 
        .ZN(\SB1_1_6/buf_output[3] ) );
  XOR2_X1 U14277 ( .A1(n5090), .A2(n7229), .Z(n1931) );
  XOR2_X1 U14278 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[164] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[170] ), .Z(n7229) );
  NAND3_X2 U14279 ( .A1(\SB2_0_21/i0[6] ), .A2(\SB2_0_21/i0[10] ), .A3(
        \RI3[0][62] ), .ZN(n7230) );
  INV_X2 U14280 ( .I(\SB1_1_12/buf_output[2] ), .ZN(\SB2_1_9/i1[9] ) );
  NAND3_X2 U14281 ( .A1(\SB2_4_5/i0_3 ), .A2(\SB2_4_5/i0_0 ), .A3(
        \SB1_4_6/buf_output[4] ), .ZN(n7384) );
  NAND3_X2 U14282 ( .A1(\SB1_1_23/i0[10] ), .A2(\SB1_1_23/i0_3 ), .A3(
        \SB1_1_23/i0[9] ), .ZN(\SB1_1_23/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U14283 ( .A1(\RI5[2][47] ), .A2(\RI5[2][71] ), .Z(n2388) );
  XOR2_X1 U14284 ( .A1(n7231), .A2(n119), .Z(Ciphertext[48]) );
  NAND4_X2 U14285 ( .A1(\SB4_23/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_23/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_23/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_23/Component_Function_0/NAND4_in[0] ), .ZN(n7231) );
  NAND4_X2 U14286 ( .A1(\SB1_0_25/Component_Function_0/NAND4_in[1] ), .A2(
        n5270), .A3(n5269), .A4(\SB1_0_25/Component_Function_0/NAND4_in[0] ), 
        .ZN(\SB1_0_25/buf_output[0] ) );
  NAND4_X2 U14287 ( .A1(\SB2_3_4/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_3_4/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_3_4/Component_Function_3/NAND4_in[0] ), .A4(n7234), .ZN(
        \SB2_3_4/buf_output[3] ) );
  INV_X2 U14288 ( .I(n6288), .ZN(\SB2_0_22/i1[9] ) );
  XOR2_X1 U14289 ( .A1(\RI5[2][160] ), .A2(\RI5[2][184] ), .Z(n7235) );
  XOR2_X1 U14290 ( .A1(n3762), .A2(n7236), .Z(\MC_ARK_ARC_1_0/temp5[65] ) );
  XOR2_X1 U14291 ( .A1(\RI5[0][11] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[35] ), 
        .Z(n7236) );
  XOR2_X1 U14292 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[50] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[44] ), .Z(\MC_ARK_ARC_1_1/temp1[50] ) );
  NAND3_X2 U14293 ( .A1(\SB1_3_25/i0[9] ), .A2(\SB1_3_25/i1_5 ), .A3(
        \SB1_3_25/i0[6] ), .ZN(\SB1_3_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U14294 ( .A1(\SB1_3_15/i0[10] ), .A2(\SB1_3_15/i1_5 ), .A3(n5431), 
        .ZN(\SB1_3_15/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U14295 ( .A1(\SB1_3_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_26/Component_Function_4/NAND4_in[3] ), .A4(n7238), .ZN(
        \SB1_3_26/buf_output[4] ) );
  NAND4_X2 U14296 ( .A1(\SB2_3_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_25/Component_Function_5/NAND4_in[1] ), .A3(n7367), .A4(
        \SB2_3_25/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_25/buf_output[5] ) );
  NAND3_X1 U14297 ( .A1(\SB4_23/i0_4 ), .A2(\SB4_23/i1[9] ), .A3(\SB4_23/i1_5 ), .ZN(\SB4_23/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U14298 ( .A1(\MC_ARK_ARC_1_2/temp5[35] ), .A2(n5171), .Z(
        \MC_ARK_ARC_1_2/buf_output[35] ) );
  XOR2_X1 U14299 ( .A1(\RI5[2][107] ), .A2(\RI5[2][71] ), .Z(
        \MC_ARK_ARC_1_2/temp3[5] ) );
  XOR2_X1 U14300 ( .A1(\RI5[0][65] ), .A2(\RI5[0][191] ), .Z(n5096) );
  NAND4_X2 U14301 ( .A1(\SB2_2_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_29/Component_Function_5/NAND4_in[0] ), .A4(n7239), .ZN(
        \SB2_2_29/buf_output[5] ) );
  NAND3_X2 U14302 ( .A1(\SB2_2_29/i0[6] ), .A2(\SB2_2_29/i0_4 ), .A3(
        \SB2_2_29/i0[9] ), .ZN(n7239) );
  NAND3_X2 U14303 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0[9] ), .A3(
        \SB1_0_25/i0[8] ), .ZN(n3303) );
  XOR2_X1 U14304 ( .A1(n2623), .A2(\MC_ARK_ARC_1_0/temp6[155] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[155] ) );
  NAND4_X2 U14305 ( .A1(\SB1_0_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_25/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_0_25/Component_Function_1/NAND4_in[3] ), .A4(n7268), .ZN(
        \SB1_0_25/buf_output[1] ) );
  XOR2_X1 U14306 ( .A1(\RI5[0][182] ), .A2(n452), .Z(n7241) );
  XOR2_X1 U14307 ( .A1(\RI5[0][56] ), .A2(\RI5[0][158] ), .Z(n7242) );
  NAND4_X2 U14308 ( .A1(\SB2_1_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_27/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_27/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_1_27/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_1_27/buf_output[2] ) );
  XOR2_X1 U14309 ( .A1(\SB2_4_22/buf_output[4] ), .A2(\RI5[4][88] ), .Z(
        \MC_ARK_ARC_1_4/temp2[118] ) );
  NAND4_X2 U14310 ( .A1(\SB3_10/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_10/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_10/Component_Function_0/NAND4_in[1] ), .A4(
        \SB3_10/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_10/buf_output[0] ) );
  XOR2_X1 U14311 ( .A1(n7243), .A2(n77), .Z(Ciphertext[161]) );
  NAND4_X2 U14312 ( .A1(\SB4_5/Component_Function_5/NAND4_in[2] ), .A2(n3788), 
        .A3(\SB4_5/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_5/Component_Function_5/NAND4_in[0] ), .ZN(n7243) );
  XOR2_X1 U14313 ( .A1(n7244), .A2(\MC_ARK_ARC_1_2/temp5[99] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[99] ) );
  XOR2_X1 U14314 ( .A1(\RI5[1][59] ), .A2(\RI5[1][23] ), .Z(
        \MC_ARK_ARC_1_1/temp3[149] ) );
  XOR2_X1 U14315 ( .A1(\MC_ARK_ARC_1_2/temp6[18] ), .A2(n7245), .Z(
        \MC_ARK_ARC_1_2/buf_output[18] ) );
  XOR2_X1 U14316 ( .A1(\MC_ARK_ARC_1_2/temp1[18] ), .A2(n7470), .Z(n7245) );
  NAND4_X2 U14317 ( .A1(\SB2_4_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_4_27/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_4_27/Component_Function_1/NAND4_in[0] ), .A4(n7246), .ZN(
        \SB2_4_27/buf_output[1] ) );
  NAND3_X1 U14318 ( .A1(\SB2_4_27/i0_4 ), .A2(\SB2_4_27/i1_7 ), .A3(
        \SB2_4_27/i0[8] ), .ZN(n7246) );
  NAND3_X1 U14319 ( .A1(\SB3_29/i0[6] ), .A2(\SB3_29/i1[9] ), .A3(\RI1[5][17] ), .ZN(\SB3_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U14320 ( .A1(\SB4_31/i0_3 ), .A2(\SB4_31/i0[6] ), .A3(
        \SB4_31/i1[9] ), .ZN(n7248) );
  NAND4_X2 U14321 ( .A1(\SB2_0_23/Component_Function_5/NAND4_in[3] ), .A2(
        n4814), .A3(\SB2_0_23/Component_Function_5/NAND4_in[0] ), .A4(n7249), 
        .ZN(\SB2_0_23/buf_output[5] ) );
  NAND3_X2 U14322 ( .A1(\SB2_0_23/i0[10] ), .A2(\RI3[0][49] ), .A3(
        \SB2_0_23/i0_0 ), .ZN(n7249) );
  NAND3_X1 U14323 ( .A1(\SB4_8/i3[0] ), .A2(\SB4_8/i0_0 ), .A3(\SB4_8/i1_7 ), 
        .ZN(\SB4_8/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U14324 ( .A1(\MC_ARK_ARC_1_2/temp2[71] ), .A2(n7251), .Z(
        \MC_ARK_ARC_1_2/temp5[71] ) );
  XOR2_X1 U14325 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[65] ), .A2(\RI5[2][71] ), 
        .Z(n7251) );
  NAND4_X2 U14326 ( .A1(\SB2_1_15/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_15/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_15/Component_Function_4/NAND4_in[3] ), .A4(n7252), .ZN(
        \SB2_1_15/buf_output[4] ) );
  XOR2_X1 U14327 ( .A1(\MC_ARK_ARC_1_3/temp4[27] ), .A2(n7253), .Z(n3840) );
  XOR2_X1 U14328 ( .A1(\RI5[3][165] ), .A2(\RI5[3][189] ), .Z(n7253) );
  NAND3_X2 U14329 ( .A1(\SB3_25/i0[10] ), .A2(\SB3_25/i0[6] ), .A3(
        \SB3_25/i0_3 ), .ZN(n7254) );
  NAND4_X2 U14330 ( .A1(\SB2_3_7/Component_Function_2/NAND4_in[2] ), .A2(n2159), .A3(\SB2_3_7/Component_Function_2/NAND4_in[0] ), .A4(n7255), .ZN(
        \SB2_3_7/buf_output[2] ) );
  NAND3_X1 U14331 ( .A1(\SB2_1_11/i0[6] ), .A2(\SB2_1_11/i0[8] ), .A3(
        \SB2_1_11/i0[7] ), .ZN(\SB2_1_11/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U14332 ( .A1(\SB2_2_11/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_11/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_2_11/Component_Function_0/NAND4_in[0] ), .A4(n7256), .ZN(
        \SB2_2_11/buf_output[0] ) );
  NAND3_X1 U14333 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i0[10] ), .A3(
        \SB2_2_11/i0_3 ), .ZN(n7256) );
  NAND4_X2 U14334 ( .A1(\SB2_4_24/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_4_24/Component_Function_3/NAND4_in[3] ), .A4(n7257), .ZN(
        \SB2_4_24/buf_output[3] ) );
  NAND3_X1 U14335 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i1[9] ), .A3(
        \SB1_0_11/i0_4 ), .ZN(\SB1_0_11/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U14336 ( .A1(\SB3_2/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_2/Component_Function_1/NAND4_in[1] ), .A3(n1176), .A4(n2597), 
        .ZN(\SB3_2/buf_output[1] ) );
  XOR2_X1 U14337 ( .A1(\MC_ARK_ARC_1_2/temp6[167] ), .A2(n7260), .Z(
        \MC_ARK_ARC_1_2/buf_output[167] ) );
  XOR2_X1 U14338 ( .A1(n7408), .A2(\MC_ARK_ARC_1_2/temp1[167] ), .Z(n7260) );
  NAND3_X1 U14339 ( .A1(\SB1_3_21/i0[9] ), .A2(\SB1_3_21/i0_0 ), .A3(
        \SB1_3_21/i0[8] ), .ZN(n7261) );
  XOR2_X1 U14340 ( .A1(n7263), .A2(n7262), .Z(\MC_ARK_ARC_1_2/buf_output[14] )
         );
  XOR2_X1 U14341 ( .A1(n753), .A2(\MC_ARK_ARC_1_2/temp4[14] ), .Z(n7263) );
  XOR2_X1 U14342 ( .A1(\MC_ARK_ARC_1_1/temp5[74] ), .A2(n7264), .Z(
        \MC_ARK_ARC_1_1/buf_output[74] ) );
  XOR2_X1 U14343 ( .A1(\MC_ARK_ARC_1_1/temp3[74] ), .A2(
        \MC_ARK_ARC_1_1/temp4[74] ), .Z(n7264) );
  XOR2_X1 U14344 ( .A1(\RI5[2][19] ), .A2(\RI5[2][13] ), .Z(
        \MC_ARK_ARC_1_2/temp1[19] ) );
  NAND3_X1 U14345 ( .A1(\SB2_4_2/i0[6] ), .A2(\SB2_4_2/i0_0 ), .A3(
        \SB2_4_2/i0[10] ), .ZN(\SB2_4_2/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 U14346 ( .A1(\SB1_1_8/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_8/Component_Function_1/NAND4_in[2] ), .ZN(n2756) );
  XOR2_X1 U14347 ( .A1(\RI5[0][58] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[64] ), 
        .Z(n7266) );
  NAND3_X1 U14348 ( .A1(\SB3_29/i0_0 ), .A2(\SB3_29/i0[7] ), .A3(\RI1[5][17] ), 
        .ZN(\SB3_29/Component_Function_0/NAND4_in[3] ) );
  AND2_X1 U14349 ( .A1(n227), .A2(n265), .Z(n7269) );
  NAND3_X1 U14350 ( .A1(\SB2_0_15/i0[6] ), .A2(\SB2_0_15/i1_5 ), .A3(
        \RI3[0][96] ), .ZN(n7270) );
  XOR2_X1 U14351 ( .A1(\RI5[1][129] ), .A2(\RI5[1][135] ), .Z(n7271) );
  NAND4_X2 U14352 ( .A1(n3162), .A2(n5352), .A3(
        \SB2_3_31/Component_Function_5/NAND4_in[0] ), .A4(n7272), .ZN(
        \SB2_3_31/buf_output[5] ) );
  NAND3_X2 U14353 ( .A1(\SB2_3_31/i0[10] ), .A2(\SB2_3_31/i0_0 ), .A3(
        \SB2_3_31/i0[6] ), .ZN(n7272) );
  NAND3_X1 U14354 ( .A1(\SB1_4_6/i1_5 ), .A2(\SB1_4_6/i0_4 ), .A3(
        \SB1_4_6/i1[9] ), .ZN(\SB1_4_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U14355 ( .A1(\SB1_1_20/i0_0 ), .A2(\SB1_1_20/i1_7 ), .A3(
        \SB1_1_20/i3[0] ), .ZN(n7273) );
  NAND4_X2 U14356 ( .A1(\SB2_3_22/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_3_22/Component_Function_5/NAND4_in[2] ), .A3(n2694), .A4(n7274), 
        .ZN(\SB2_3_22/buf_output[5] ) );
  NAND3_X2 U14357 ( .A1(\SB2_3_22/i0_0 ), .A2(\SB2_3_22/i0[10] ), .A3(
        \SB2_3_22/i0[6] ), .ZN(n7274) );
  XOR2_X1 U14358 ( .A1(\MC_ARK_ARC_1_3/temp2[20] ), .A2(
        \MC_ARK_ARC_1_3/temp4[20] ), .Z(n7275) );
  NAND3_X1 U14359 ( .A1(\SB2_4_17/i0_3 ), .A2(\SB2_4_17/i0[7] ), .A3(
        \SB2_4_17/i0_0 ), .ZN(\SB2_4_17/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U14360 ( .A1(\MC_ARK_ARC_1_3/temp2[134] ), .A2(n4268), .Z(n3495) );
  NAND4_X2 U14361 ( .A1(\SB2_1_29/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_1_29/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_29/Component_Function_4/NAND4_in[1] ), .A4(n7276), .ZN(
        \SB2_1_29/buf_output[4] ) );
  NAND3_X1 U14362 ( .A1(\SB2_1_29/i1[9] ), .A2(\SB2_1_29/i1_5 ), .A3(
        \SB2_1_29/i0_4 ), .ZN(n7276) );
  NAND3_X2 U14363 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i0[10] ), .A3(
        \SB1_3_18/i0[6] ), .ZN(\SB1_3_18/Component_Function_5/NAND4_in[1] ) );
  OR3_X2 U14364 ( .A1(\MC_ARK_ARC_1_0/buf_output[54] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[57] ), .A3(\MC_ARK_ARC_1_0/buf_output[59] ), 
        .Z(n7492) );
  NAND3_X2 U14365 ( .A1(\SB2_0_16/i0[6] ), .A2(n594), .A3(\SB2_0_16/i0[9] ), 
        .ZN(n1283) );
  XOR2_X1 U14366 ( .A1(\RI5[0][74] ), .A2(\RI5[0][110] ), .Z(
        \MC_ARK_ARC_1_0/temp3[8] ) );
  NAND3_X2 U14367 ( .A1(\SB2_2_12/i0[10] ), .A2(\SB2_2_12/i0_0 ), .A3(
        \SB2_2_12/i0[6] ), .ZN(\SB2_2_12/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U14368 ( .A1(\RI5[3][93] ), .A2(\RI5[3][87] ), .Z(n907) );
  NAND4_X2 U14369 ( .A1(\SB1_2_26/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_26/Component_Function_0/NAND4_in[1] ), .A3(n5207), .A4(
        \SB1_2_26/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_26/buf_output[0] ) );
  XOR2_X1 U14370 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[22] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[178] ), .Z(\MC_ARK_ARC_1_1/temp3[112] )
         );
  NAND4_X2 U14371 ( .A1(\SB2_3_22/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_3_22/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_22/Component_Function_2/NAND4_in[2] ), .A4(n7278), .ZN(
        \SB2_3_22/buf_output[2] ) );
  NAND3_X2 U14372 ( .A1(\SB2_3_22/i0_0 ), .A2(\RI3[3][58] ), .A3(
        \SB2_3_22/i1_5 ), .ZN(n7278) );
  NAND4_X2 U14373 ( .A1(n3957), .A2(\SB1_4_6/Component_Function_3/NAND4_in[1] ), .A3(\SB1_4_6/Component_Function_3/NAND4_in[0] ), .A4(n2911), .ZN(
        \SB1_4_6/buf_output[3] ) );
  XOR2_X1 U14374 ( .A1(\RI5[3][180] ), .A2(\RI5[3][150] ), .Z(n7279) );
  XOR2_X1 U14375 ( .A1(n7281), .A2(\MC_ARK_ARC_1_3/temp4[182] ), .Z(n3639) );
  XOR2_X1 U14376 ( .A1(\RI5[3][152] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[128] ), .Z(n7281) );
  XOR2_X1 U14377 ( .A1(n7282), .A2(n7283), .Z(\MC_ARK_ARC_1_2/temp5[172] ) );
  XOR2_X1 U14378 ( .A1(\RI5[2][142] ), .A2(\RI5[2][118] ), .Z(n7282) );
  XOR2_X1 U14379 ( .A1(\RI5[2][166] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[172] ), .Z(n7283) );
  NOR2_X1 U14380 ( .A1(\MC_ARK_ARC_1_1/buf_output[147] ), .A2(
        \MC_ARK_ARC_1_1/buf_output[144] ), .ZN(n7285) );
  NAND3_X2 U14381 ( .A1(\SB1_0_8/i0_0 ), .A2(\SB1_0_8/i0_3 ), .A3(
        \SB1_0_8/i0[7] ), .ZN(n7287) );
  NAND3_X1 U14382 ( .A1(\SB2_3_0/i0_0 ), .A2(\SB2_3_0/i3[0] ), .A3(
        \SB2_3_0/i1_7 ), .ZN(n7288) );
  XOR2_X1 U14383 ( .A1(\MC_ARK_ARC_1_3/temp1[10] ), .A2(
        \MC_ARK_ARC_1_3/temp2[10] ), .Z(n7289) );
  NAND4_X2 U14384 ( .A1(\SB1_4_30/Component_Function_0/NAND4_in[1] ), .A2(
        n4848), .A3(\SB1_4_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_4_30/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_4_30/buf_output[0] ) );
  XOR2_X1 U14385 ( .A1(n7290), .A2(n53), .Z(Ciphertext[24]) );
  NAND4_X2 U14386 ( .A1(n7333), .A2(\SB4_27/Component_Function_0/NAND4_in[2] ), 
        .A3(n898), .A4(\SB4_27/Component_Function_0/NAND4_in[0] ), .ZN(n7290)
         );
  XOR2_X1 U14387 ( .A1(\MC_ARK_ARC_1_0/temp2[40] ), .A2(n7291), .Z(
        \MC_ARK_ARC_1_0/temp5[40] ) );
  XOR2_X1 U14388 ( .A1(\RI5[0][34] ), .A2(\RI5[0][40] ), .Z(n7291) );
  XOR2_X1 U14389 ( .A1(\MC_ARK_ARC_1_0/temp4[41] ), .A2(n7459), .Z(n7292) );
  XOR2_X1 U14390 ( .A1(\RI5[0][24] ), .A2(\RI5[0][0] ), .Z(
        \MC_ARK_ARC_1_0/temp2[54] ) );
  NAND3_X2 U14391 ( .A1(\SB1_3_12/i0_0 ), .A2(\SB1_3_12/i1_5 ), .A3(
        \SB1_3_12/i0_4 ), .ZN(\SB1_3_12/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U14392 ( .A1(\MC_ARK_ARC_1_3/temp3[32] ), .A2(
        \MC_ARK_ARC_1_3/temp4[32] ), .Z(n3956) );
  NAND3_X2 U14393 ( .A1(\SB1_3_22/i0_4 ), .A2(\SB1_3_22/i0_3 ), .A3(
        \SB1_3_22/i1[9] ), .ZN(n7294) );
  XOR2_X1 U14394 ( .A1(\RI5[2][119] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[143] ), .Z(n7295) );
  XOR2_X1 U14395 ( .A1(\MC_ARK_ARC_1_4/temp6[134] ), .A2(n7296), .Z(
        \MC_ARK_ARC_1_4/buf_output[134] ) );
  XOR2_X1 U14396 ( .A1(n7297), .A2(n660), .Z(\MC_ARK_ARC_1_4/temp5[114] ) );
  XOR2_X1 U14397 ( .A1(\RI5[4][114] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[108] ), .Z(n7297) );
  XOR2_X1 U14398 ( .A1(\MC_ARK_ARC_1_1/temp2[177] ), .A2(n7298), .Z(
        \MC_ARK_ARC_1_1/temp5[177] ) );
  XOR2_X1 U14399 ( .A1(\RI5[1][171] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[177] ), .Z(n7298) );
  XOR2_X1 U14400 ( .A1(\RI5[2][160] ), .A2(\RI5[2][154] ), .Z(n7299) );
  AOI21_X1 U14401 ( .A1(n7390), .A2(\SB4_19/i0_0 ), .B(n6273), .ZN(n4679) );
  NAND3_X1 U14402 ( .A1(\SB3_29/i0_0 ), .A2(\SB3_29/i0[9] ), .A3(
        \SB3_29/i0[8] ), .ZN(\SB3_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U14403 ( .A1(\SB1_2_22/i0[6] ), .A2(\SB1_2_22/i0[8] ), .A3(
        \SB1_2_22/i0[7] ), .ZN(\SB1_2_22/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U14404 ( .A1(\SB2_4_9/Component_Function_5/NAND4_in[1] ), .A2(n5140), .A3(n7424), .A4(n7300), .ZN(\SB2_4_9/buf_output[5] ) );
  NAND2_X2 U14405 ( .A1(\SB2_4_9/i0_0 ), .A2(\SB2_4_9/i3[0] ), .ZN(n7300) );
  NAND4_X2 U14406 ( .A1(\SB1_2_30/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_30/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_30/Component_Function_4/NAND4_in[3] ), .A4(n7302), .ZN(
        \SB1_2_30/buf_output[4] ) );
  XOR2_X1 U14407 ( .A1(n7303), .A2(n7389), .Z(\MC_ARK_ARC_1_2/temp5[147] ) );
  XOR2_X1 U14408 ( .A1(\RI5[2][117] ), .A2(\RI5[2][93] ), .Z(n7303) );
  XOR2_X1 U14409 ( .A1(\MC_ARK_ARC_1_0/temp3[173] ), .A2(n7304), .Z(n7422) );
  XOR2_X1 U14410 ( .A1(\RI5[0][143] ), .A2(\RI5[0][119] ), .Z(n7304) );
  XOR2_X1 U14411 ( .A1(n7565), .A2(\MC_ARK_ARC_1_1/temp1[115] ), .Z(n7305) );
  NAND4_X2 U14412 ( .A1(n1146), .A2(n4286), .A3(n5275), .A4(n7306), .ZN(n7569)
         );
  NAND3_X1 U14413 ( .A1(\SB4_10/i1[9] ), .A2(\SB4_10/i0_4 ), .A3(\SB4_10/i1_5 ), .ZN(n7306) );
  XOR2_X1 U14414 ( .A1(n7307), .A2(\MC_ARK_ARC_1_3/temp1[162] ), .Z(
        \MC_ARK_ARC_1_3/temp5[162] ) );
  XOR2_X1 U14415 ( .A1(\RI5[3][132] ), .A2(\RI5[3][108] ), .Z(n7307) );
  XOR2_X1 U14416 ( .A1(\RI5[4][102] ), .A2(\MC_ARK_ARC_1_4/buf_datainput[108] ), .Z(n7308) );
  XOR2_X1 U14417 ( .A1(n7310), .A2(n7309), .Z(\MC_ARK_ARC_1_2/temp6[170] ) );
  XOR2_X1 U14418 ( .A1(\RI5[2][44] ), .A2(n123), .Z(n7309) );
  XOR2_X1 U14419 ( .A1(\RI5[2][87] ), .A2(\RI5[2][81] ), .Z(
        \MC_ARK_ARC_1_2/temp1[87] ) );
  NAND3_X1 U14420 ( .A1(\SB2_4_4/i0_3 ), .A2(\SB2_4_4/i0_0 ), .A3(
        \SB2_4_4/i0[7] ), .ZN(\SB2_4_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U14421 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i0[9] ), .A3(
        \SB1_0_11/i0[10] ), .ZN(\SB1_0_11/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U14422 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i0_0 ), .A3(
        \SB1_0_20/i0_4 ), .ZN(\SB1_0_20/Component_Function_3/NAND4_in[1] ) );
  AND2_X1 U14423 ( .A1(n3668), .A2(\SB1_2_27/Component_Function_4/NAND4_in[3] ), .Z(n7311) );
  XOR2_X1 U14424 ( .A1(n7313), .A2(n7312), .Z(\MC_ARK_ARC_1_0/buf_output[134] ) );
  XOR2_X1 U14425 ( .A1(n4617), .A2(n1993), .Z(n7313) );
  XOR2_X1 U14426 ( .A1(\RI5[4][68] ), .A2(\RI5[4][20] ), .Z(n7314) );
  XOR2_X1 U14427 ( .A1(\RI5[4][44] ), .A2(\RI5[4][74] ), .Z(n7315) );
  NAND4_X2 U14428 ( .A1(\SB2_0_18/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_18/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_0_18/Component_Function_1/NAND4_in[0] ), .A4(n7316), .ZN(
        \SB2_0_18/buf_output[1] ) );
  XOR2_X1 U14429 ( .A1(\RI5[2][129] ), .A2(\RI5[2][93] ), .Z(
        \MC_ARK_ARC_1_2/temp3[27] ) );
  NAND3_X1 U14430 ( .A1(\SB2_0_29/i0[9] ), .A2(\SB2_0_29/i1_5 ), .A3(
        \SB1_0_1/buf_output[1] ), .ZN(
        \SB2_0_29/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U14431 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[39] ), .A2(\RI5[3][45] ), 
        .Z(n7317) );
  NAND3_X1 U14432 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0[10] ), .A3(
        \SB1_0_2/i0_4 ), .ZN(\SB1_0_2/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U14433 ( .A1(\SB1_0_2/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_2/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_0_2/Component_Function_2/NAND4_in[0] ), .A4(n1839), .ZN(
        \SB1_0_2/buf_output[2] ) );
  NAND4_X2 U14434 ( .A1(\SB2_1_11/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_1/NAND4_in[0] ), .A4(n7318), .ZN(
        \SB2_1_11/buf_output[1] ) );
  NAND4_X2 U14435 ( .A1(\SB2_3_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_3/NAND4_in[1] ), .A3(n5332), .A4(
        \SB2_3_3/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_3_3/buf_output[3] ) );
  XOR2_X1 U14436 ( .A1(n6285), .A2(n4652), .Z(\MC_ARK_ARC_1_2/temp5[2] ) );
  XOR2_X1 U14437 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[164] ), .A2(\RI5[2][188] ), .Z(n2961) );
  XOR2_X1 U14438 ( .A1(\RI5[1][25] ), .A2(\RI5[1][19] ), .Z(
        \MC_ARK_ARC_1_1/temp1[25] ) );
  XOR2_X1 U14439 ( .A1(n7319), .A2(n173), .Z(Ciphertext[76]) );
  XOR2_X1 U14440 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[35] ), .A2(\RI5[2][59] ), 
        .Z(n7320) );
  NAND3_X1 U14441 ( .A1(\SB4_21/i0[9] ), .A2(\SB4_21/i0_3 ), .A3(
        \SB4_21/i0[8] ), .ZN(\SB4_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U14442 ( .A1(\SB2_1_31/i0[7] ), .A2(\SB2_1_31/i0_0 ), .A3(
        \SB2_1_31/i0_3 ), .ZN(\SB2_1_31/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U14443 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[169] ), .A2(\RI5[4][1] ), 
        .Z(\MC_ARK_ARC_1_4/temp2[31] ) );
  NAND3_X1 U14444 ( .A1(\SB2_3_29/i1[9] ), .A2(\SB2_3_29/i0_4 ), .A3(
        \SB2_3_29/i1_5 ), .ZN(\SB2_3_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U14445 ( .A1(\SB2_0_1/i0_4 ), .A2(\SB2_0_1/i0[6] ), .A3(
        \SB2_0_1/i0[9] ), .ZN(n7322) );
  NAND4_X2 U14446 ( .A1(\SB2_4_27/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_4_27/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_4_27/Component_Function_2/NAND4_in[2] ), .A4(n4055), .ZN(
        \SB2_4_27/buf_output[2] ) );
  XOR2_X1 U14447 ( .A1(n4542), .A2(\MC_ARK_ARC_1_1/temp4[23] ), .Z(n3344) );
  XOR2_X1 U14448 ( .A1(\RI5[1][28] ), .A2(\RI5[1][52] ), .Z(n7323) );
  XOR2_X1 U14449 ( .A1(\RI5[3][119] ), .A2(\RI5[3][185] ), .Z(n3205) );
  XOR2_X1 U14450 ( .A1(\RI5[2][128] ), .A2(\RI5[2][134] ), .Z(
        \MC_ARK_ARC_1_2/temp1[134] ) );
  XOR2_X1 U14451 ( .A1(\MC_ARK_ARC_1_2/temp5[134] ), .A2(
        \MC_ARK_ARC_1_2/temp6[134] ), .Z(\MC_ARK_ARC_1_2/buf_output[134] ) );
  NAND4_X2 U14452 ( .A1(\SB1_4_18/Component_Function_2/NAND4_in[1] ), .A2(
        n3306), .A3(\SB1_4_18/Component_Function_2/NAND4_in[0] ), .A4(n7427), 
        .ZN(\SB1_4_18/buf_output[2] ) );
  NAND3_X1 U14453 ( .A1(\SB1_2_3/i1[9] ), .A2(\SB1_2_3/i1_5 ), .A3(
        \MC_ARK_ARC_1_1/buf_output[172] ), .ZN(
        \SB1_2_3/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U14454 ( .A1(\MC_ARK_ARC_1_4/temp5[31] ), .A2(n763), .Z(
        \MC_ARK_ARC_1_4/buf_output[31] ) );
  NAND4_X2 U14455 ( .A1(n2337), .A2(\SB3_19/Component_Function_5/NAND4_in[1] ), 
        .A3(n5411), .A4(\SB3_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_19/buf_output[5] ) );
  NAND3_X1 U14456 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i1_7 ), .A3(\SB4_11/i3[0] ), .ZN(n7324) );
  NAND4_X2 U14457 ( .A1(\SB2_1_12/Component_Function_5/NAND4_in[2] ), .A2(
        n3883), .A3(n4405), .A4(n1148), .ZN(\SB2_1_12/buf_output[5] ) );
  XOR2_X1 U14458 ( .A1(\MC_ARK_ARC_1_0/temp6[3] ), .A2(n7326), .Z(
        \MC_ARK_ARC_1_0/buf_output[3] ) );
  XOR2_X1 U14459 ( .A1(\MC_ARK_ARC_1_0/temp1[3] ), .A2(n3648), .Z(n7326) );
  NAND3_X1 U14460 ( .A1(\MC_ARK_ARC_1_2/buf_output[94] ), .A2(\SB1_3_16/i0_0 ), 
        .A3(\SB1_3_16/i1_5 ), .ZN(n3520) );
  XOR2_X1 U14461 ( .A1(\RI5[0][20] ), .A2(\RI5[0][56] ), .Z(n7327) );
  XOR2_X1 U14462 ( .A1(n7328), .A2(n3902), .Z(\MC_ARK_ARC_1_2/buf_output[136] ) );
  XOR2_X1 U14463 ( .A1(\MC_ARK_ARC_1_2/temp3[136] ), .A2(
        \MC_ARK_ARC_1_2/temp1[136] ), .Z(n7328) );
  NAND4_X2 U14464 ( .A1(\SB2_3_4/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_4/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_4/Component_Function_4/NAND4_in[1] ), .A4(n7329), .ZN(
        \SB2_3_4/buf_output[4] ) );
  NAND3_X1 U14465 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i0[10] ), .A3(
        \SB2_3_4/i0[9] ), .ZN(n7329) );
  NAND3_X1 U14466 ( .A1(\SB1_2_27/i0[6] ), .A2(\SB1_2_27/i0[9] ), .A3(
        \SB1_2_27/i1_5 ), .ZN(n7331) );
  XOR2_X1 U14467 ( .A1(n7332), .A2(n7), .Z(Ciphertext[108]) );
  NAND4_X2 U14468 ( .A1(\SB4_13/Component_Function_0/NAND4_in[1] ), .A2(n729), 
        .A3(n2697), .A4(\SB4_13/Component_Function_0/NAND4_in[0] ), .ZN(n7332)
         );
  INV_X2 U14469 ( .I(\SB1_3_15/buf_output[3] ), .ZN(\SB2_3_13/i0[8] ) );
  NAND3_X1 U14470 ( .A1(\SB4_27/i0_3 ), .A2(\SB4_27/i0_0 ), .A3(\SB4_27/i0[7] ), .ZN(n7333) );
  XOR2_X1 U14471 ( .A1(\RI5[2][47] ), .A2(\RI5[2][83] ), .Z(
        \MC_ARK_ARC_1_2/temp3[173] ) );
  XOR2_X1 U14472 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[77] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[53] ), .Z(n7334) );
  NAND3_X1 U14473 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i0[10] ), .A3(
        \SB1_0_11/i0_4 ), .ZN(\SB1_0_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U14474 ( .A1(\SB1_4_18/i0_3 ), .A2(\SB1_4_18/i0[10] ), .A3(
        \SB1_4_18/i0_4 ), .ZN(\SB1_4_18/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U14475 ( .A1(\SB2_2_23/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_23/Component_Function_1/NAND4_in[0] ), .A4(n7336), .ZN(
        \SB2_2_23/buf_output[1] ) );
  NAND3_X1 U14476 ( .A1(\SB2_2_23/i0[6] ), .A2(\SB2_2_23/i1_5 ), .A3(
        \SB2_2_23/i0[9] ), .ZN(n7336) );
  XOR2_X1 U14477 ( .A1(n7337), .A2(n118), .Z(Ciphertext[109]) );
  NAND4_X2 U14478 ( .A1(n2183), .A2(\SB4_13/Component_Function_1/NAND4_in[1] ), 
        .A3(\SB4_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_13/Component_Function_1/NAND4_in[0] ), .ZN(n7337) );
  NAND3_X2 U14479 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i0[9] ), .A3(
        \SB2_3_1/i0[10] ), .ZN(\SB2_3_1/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U14480 ( .A1(\MC_ARK_ARC_1_3/temp2[5] ), .A2(n7339), .Z(
        \MC_ARK_ARC_1_3/temp5[5] ) );
  XOR2_X1 U14481 ( .A1(\MC_ARK_ARC_1_4/temp1[176] ), .A2(n7340), .Z(n7437) );
  XOR2_X1 U14482 ( .A1(\RI5[4][122] ), .A2(\RI5[4][146] ), .Z(n7340) );
  INV_X1 U14483 ( .I(\SB3_2/buf_output[2] ), .ZN(\SB4_31/i1[9] ) );
  NAND4_X2 U14484 ( .A1(n4910), .A2(\SB3_2/Component_Function_2/NAND4_in[1] ), 
        .A3(n7428), .A4(\SB3_2/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB3_2/buf_output[2] ) );
  XOR2_X1 U14485 ( .A1(\MC_ARK_ARC_1_3/temp2[58] ), .A2(
        \MC_ARK_ARC_1_3/temp1[58] ), .Z(\MC_ARK_ARC_1_3/temp5[58] ) );
  NAND3_X1 U14486 ( .A1(\SB1_3_1/i0[6] ), .A2(\SB1_3_1/i0[8] ), .A3(
        \SB1_3_1/i0[7] ), .ZN(\SB1_3_1/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U14487 ( .A1(\SB1_0_11/Component_Function_2/NAND4_in[2] ), .A2(
        n3891), .A3(n5158), .A4(n7342), .ZN(\RI3[0][140] ) );
  NAND3_X2 U14488 ( .A1(\SB1_0_11/i0_0 ), .A2(\SB1_0_11/i0_4 ), .A3(
        \SB1_0_11/i1_5 ), .ZN(n7342) );
  NAND3_X2 U14489 ( .A1(\SB2_2_4/i0_0 ), .A2(\SB2_2_4/i0[10] ), .A3(
        \SB2_2_4/i0[6] ), .ZN(\SB2_2_4/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U14490 ( .A1(\SB4_10/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_10/Component_Function_5/NAND4_in[2] ), .A3(n2925), .A4(n7345), 
        .ZN(n3364) );
  NAND3_X1 U14491 ( .A1(\SB4_10/i0[6] ), .A2(\SB4_10/i0[9] ), .A3(
        \SB4_10/i0_4 ), .ZN(n7345) );
  NAND4_X2 U14492 ( .A1(\SB1_2_5/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_5/Component_Function_0/NAND4_in[0] ), .A4(n7346), .ZN(
        \SB1_2_5/buf_output[0] ) );
  XOR2_X1 U14493 ( .A1(\RI5[2][176] ), .A2(\RI5[2][170] ), .Z(
        \MC_ARK_ARC_1_2/temp1[176] ) );
  NAND3_X2 U14494 ( .A1(\SB2_3_9/i0[10] ), .A2(\SB2_3_9/i1_7 ), .A3(
        \SB2_3_9/i1[9] ), .ZN(n7348) );
  XOR2_X1 U14495 ( .A1(n7350), .A2(n7349), .Z(\MC_ARK_ARC_1_4/buf_output[113] ) );
  XOR2_X1 U14496 ( .A1(n1919), .A2(n4915), .Z(\MC_ARK_ARC_1_2/buf_output[7] )
         );
  XOR2_X1 U14497 ( .A1(n7351), .A2(n4447), .Z(\MC_ARK_ARC_1_4/temp5[185] ) );
  XOR2_X1 U14498 ( .A1(\RI5[4][155] ), .A2(\RI5[4][131] ), .Z(n7351) );
  NAND3_X2 U14499 ( .A1(\SB1_2_28/i0_0 ), .A2(\SB1_2_28/i1_5 ), .A3(
        \SB1_2_28/i0_4 ), .ZN(n7352) );
  NAND4_X2 U14500 ( .A1(n3787), .A2(
        \SB2_0_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_25/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_0_25/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_0_25/buf_output[5] ) );
  NAND4_X2 U14501 ( .A1(\SB1_1_17/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_17/Component_Function_2/NAND4_in[3] ), .A3(n1192), .A4(n7572), 
        .ZN(\SB1_1_17/buf_output[2] ) );
  NAND4_X2 U14502 ( .A1(\SB1_4_13/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_4_13/Component_Function_2/NAND4_in[3] ), .A3(n7353), .A4(n5247), 
        .ZN(\SB1_4_13/buf_output[2] ) );
  NAND3_X1 U14503 ( .A1(\SB2_3_4/i3[0] ), .A2(\SB2_3_4/i0[8] ), .A3(
        \SB2_3_4/i1_5 ), .ZN(\SB2_3_4/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U14504 ( .A1(\MC_ARK_ARC_1_4/temp5[71] ), .A2(n674), .Z(
        \MC_ARK_ARC_1_4/buf_output[71] ) );
  NAND3_X1 U14505 ( .A1(\SB1_4_13/i0[8] ), .A2(\SB1_4_13/i3[0] ), .A3(
        \SB1_4_13/i1_5 ), .ZN(\SB1_4_13/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U14506 ( .A1(\SB1_4_26/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_4_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_4_26/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_4_26/buf_output[1] ) );
  NAND4_X2 U14507 ( .A1(\SB2_0_17/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_17/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_17/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_17/buf_output[5] ) );
  NAND3_X1 U14508 ( .A1(\SB1_2_16/i0[10] ), .A2(\SB1_2_16/i1_5 ), .A3(
        \SB1_2_16/i1[9] ), .ZN(\SB1_2_16/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U14509 ( .A1(n7355), .A2(n7354), .Z(\MC_ARK_ARC_1_2/temp6[92] ) );
  XOR2_X1 U14510 ( .A1(\RI5[2][158] ), .A2(n439), .Z(n7354) );
  XOR2_X1 U14511 ( .A1(\RI5[2][90] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[84] ), 
        .Z(n7356) );
  NAND3_X1 U14512 ( .A1(\SB2_0_14/i1_5 ), .A2(\SB2_0_14/i0[9] ), .A3(
        \SB2_0_14/i0[6] ), .ZN(\SB2_0_14/Component_Function_1/NAND4_in[2] ) );
  NAND2_X2 U14513 ( .A1(n3061), .A2(
        \SB1_0_19/Component_Function_0/NAND4_in[2] ), .ZN(\SB2_0_14/i0[9] ) );
  XOR2_X1 U14514 ( .A1(n3165), .A2(\RI5[4][7] ), .Z(\MC_ARK_ARC_1_4/temp2[37] ) );
  XOR2_X1 U14515 ( .A1(n4963), .A2(n7359), .Z(\MC_ARK_ARC_1_0/buf_output[79] )
         );
  XOR2_X1 U14516 ( .A1(\MC_ARK_ARC_1_0/temp4[79] ), .A2(n1715), .Z(n7359) );
  NAND4_X2 U14517 ( .A1(\SB2_1_16/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_1_16/Component_Function_1/NAND4_in[1] ), .A3(n7360), .A4(
        \SB2_1_16/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_16/buf_output[1] ) );
  NAND3_X1 U14518 ( .A1(\SB2_3_9/i0_0 ), .A2(\SB2_3_9/i3[0] ), .A3(
        \SB2_3_9/i1_7 ), .ZN(\SB2_3_9/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U14519 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[167] ), .A2(\RI5[4][59] ), 
        .Z(n7361) );
  INV_X1 U14520 ( .I(\SB1_3_7/buf_output[1] ), .ZN(\SB2_3_3/i1_7 ) );
  NAND4_X2 U14521 ( .A1(\SB1_3_7/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_7/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_3_7/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_3_7/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_3_7/buf_output[1] ) );
  XOR2_X1 U14522 ( .A1(\MC_ARK_ARC_1_2/temp4[104] ), .A2(
        \MC_ARK_ARC_1_2/temp1[104] ), .Z(n7362) );
  NAND4_X2 U14523 ( .A1(\SB3_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_22/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_5/NAND4_in[0] ), .A4(n7364), .ZN(
        \SB3_22/buf_output[5] ) );
  XOR2_X1 U14524 ( .A1(\RI5[4][52] ), .A2(\RI5[4][16] ), .Z(
        \MC_ARK_ARC_1_4/temp3[142] ) );
  NAND4_X2 U14525 ( .A1(\SB2_1_15/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_15/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_15/Component_Function_0/NAND4_in[0] ), .A4(n7365), .ZN(
        \SB2_1_15/buf_output[0] ) );
  NAND4_X2 U14526 ( .A1(n4806), .A2(n4886), .A3(
        \SB4_22/Component_Function_2/NAND4_in[2] ), .A4(n7366), .ZN(n3215) );
  NAND3_X1 U14527 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i0[10] ), .A3(
        \SB3_26/buf_output[1] ), .ZN(n7366) );
  NAND3_X2 U14528 ( .A1(\SB2_3_25/i0_4 ), .A2(\SB2_3_25/i0[6] ), .A3(n5432), 
        .ZN(n7367) );
  XOR2_X1 U14529 ( .A1(n5206), .A2(n7368), .Z(\MC_ARK_ARC_1_4/buf_output[58] )
         );
  XOR2_X1 U14530 ( .A1(\MC_ARK_ARC_1_4/temp2[58] ), .A2(
        \MC_ARK_ARC_1_4/temp1[58] ), .Z(n7368) );
  XOR2_X1 U14531 ( .A1(\MC_ARK_ARC_1_1/temp1[132] ), .A2(
        \MC_ARK_ARC_1_1/temp2[132] ), .Z(n7369) );
  XOR2_X1 U14532 ( .A1(n7370), .A2(n108), .Z(Ciphertext[149]) );
  NAND4_X2 U14533 ( .A1(\SB4_7/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_7/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_7/Component_Function_5/NAND4_in[2] ), .A4(
        \SB4_7/Component_Function_5/NAND4_in[0] ), .ZN(n7370) );
  XOR2_X1 U14534 ( .A1(n1558), .A2(\MC_ARK_ARC_1_3/temp5[127] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[127] ) );
  NAND4_X2 U14535 ( .A1(\SB1_1_31/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_31/Component_Function_2/NAND4_in[0] ), .A3(n3723), .A4(n7371), 
        .ZN(\SB1_1_31/buf_output[2] ) );
  NAND3_X2 U14536 ( .A1(\SB1_1_31/i0_3 ), .A2(\SB1_1_31/i0[9] ), .A3(
        \SB1_1_31/i0[8] ), .ZN(n7371) );
  INV_X1 U14537 ( .I(\SB3_20/buf_output[2] ), .ZN(\SB4_17/i1[9] ) );
  NAND3_X1 U14538 ( .A1(\SB1_0_6/i0_0 ), .A2(\SB1_0_6/i0[9] ), .A3(
        \SB1_0_6/i0[8] ), .ZN(n7372) );
  XOR2_X1 U14539 ( .A1(\RI5[1][97] ), .A2(\RI5[1][133] ), .Z(n7373) );
  NAND4_X2 U14540 ( .A1(\SB2_2_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_21/Component_Function_5/NAND4_in[1] ), .A3(n7374), .A4(
        \SB2_2_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_21/buf_output[5] ) );
  NAND3_X2 U14541 ( .A1(\SB1_4_18/i0_0 ), .A2(\SB1_4_18/i0_4 ), .A3(
        \SB1_4_18/i1_5 ), .ZN(n7427) );
  NAND3_X2 U14542 ( .A1(\SB1_2_4/i0[6] ), .A2(\SB1_2_4/i0_3 ), .A3(
        \SB1_2_4/i1[9] ), .ZN(\SB1_2_4/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U14543 ( .A1(\RI5[3][42] ), .A2(\RI5[3][36] ), .Z(
        \MC_ARK_ARC_1_3/temp1[42] ) );
  NAND3_X2 U14544 ( .A1(\SB2_2_13/i0[9] ), .A2(\SB2_2_13/i0_4 ), .A3(
        \SB2_2_13/i0[6] ), .ZN(\SB2_2_13/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U14545 ( .A1(n7377), .A2(n7376), .Z(\MC_ARK_ARC_1_0/buf_output[50] )
         );
  XOR2_X1 U14546 ( .A1(n816), .A2(\MC_ARK_ARC_1_0/temp4[50] ), .Z(n7376) );
  NAND3_X2 U14547 ( .A1(\SB2_3_12/i0[9] ), .A2(\SB2_3_12/i0[6] ), .A3(n592), 
        .ZN(n7378) );
  XOR2_X1 U14548 ( .A1(n7380), .A2(\MC_ARK_ARC_1_2/temp6[114] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[114] ) );
  XOR2_X1 U14549 ( .A1(\MC_ARK_ARC_1_2/temp2[114] ), .A2(
        \MC_ARK_ARC_1_2/temp1[114] ), .Z(n7380) );
  INV_X2 U14550 ( .I(\SB1_4_28/buf_output[2] ), .ZN(\SB2_4_25/i1[9] ) );
  NAND3_X2 U14551 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i0[6] ), .A3(
        \SB2_1_20/i0_0 ), .ZN(\SB2_1_20/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U14552 ( .A1(\MC_ARK_ARC_1_0/temp1[21] ), .A2(n2434), .Z(n5134) );
  NAND4_X2 U14553 ( .A1(\SB3_23/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_23/Component_Function_0/NAND4_in[3] ), .A3(
        \SB3_23/Component_Function_0/NAND4_in[0] ), .A4(n7381), .ZN(
        \SB3_23/buf_output[0] ) );
  NAND3_X1 U14554 ( .A1(\SB3_23/i0[6] ), .A2(\SB3_23/i0[8] ), .A3(
        \SB3_23/i0[7] ), .ZN(n7381) );
  NAND3_X1 U14555 ( .A1(\SB1_2_18/i0[6] ), .A2(\MC_ARK_ARC_1_1/buf_output[78] ), .A3(\MC_ARK_ARC_1_1/buf_output[82] ), .ZN(n4149) );
  XOR2_X1 U14556 ( .A1(\RI5[0][28] ), .A2(\RI5[0][34] ), .Z(n3948) );
  XOR2_X1 U14557 ( .A1(\MC_ARK_ARC_1_0/temp5[59] ), .A2(n5004), .Z(
        \MC_ARK_ARC_1_0/buf_output[59] ) );
  XOR2_X1 U14558 ( .A1(\MC_ARK_ARC_1_1/temp2[79] ), .A2(n7382), .Z(
        \MC_ARK_ARC_1_1/temp5[79] ) );
  XOR2_X1 U14559 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[73] ), .A2(\RI5[1][79] ), 
        .Z(n7382) );
  NAND3_X1 U14560 ( .A1(\SB1_4_2/i0_3 ), .A2(\SB1_4_2/i0[8] ), .A3(
        \SB1_4_2/i1_7 ), .ZN(\SB1_4_2/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U14561 ( .A1(\SB2_1_16/Component_Function_5/NAND4_in[0] ), .A2(
        n3149), .A3(n7409), .A4(n1137), .ZN(\SB2_1_16/buf_output[5] ) );
  NAND4_X2 U14562 ( .A1(n917), .A2(\SB2_1_0/Component_Function_0/NAND4_in[2] ), 
        .A3(\SB2_1_0/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_1_0/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_1_0/buf_output[0] ) );
  XOR2_X1 U14563 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[71] ), .A2(\RI5[0][65] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[71] ) );
  XOR2_X1 U14564 ( .A1(n3777), .A2(n3776), .Z(\MC_ARK_ARC_1_3/buf_output[167] ) );
  XOR2_X1 U14565 ( .A1(n3085), .A2(n1391), .Z(\MC_ARK_ARC_1_3/buf_output[177] ) );
  NAND3_X1 U14566 ( .A1(\SB1_2_7/i1_5 ), .A2(\SB1_2_7/i1[9] ), .A3(
        \SB1_2_7/i0_4 ), .ZN(\SB1_2_7/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U14567 ( .A1(\MC_ARK_ARC_1_4/temp5[105] ), .A2(n7383), .Z(
        \MC_ARK_ARC_1_4/buf_output[105] ) );
  NAND4_X2 U14568 ( .A1(\SB3_6/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_6/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_6/Component_Function_4/NAND4_in[1] ), .A4(n7385), .ZN(
        \SB3_6/buf_output[4] ) );
  NAND4_X2 U14569 ( .A1(\SB1_4_5/Component_Function_5/NAND4_in[1] ), .A2(n5238), .A3(\SB1_4_5/Component_Function_5/NAND4_in[0] ), .A4(n7386), .ZN(
        \SB1_4_5/buf_output[5] ) );
  NAND3_X2 U14570 ( .A1(\SB1_4_5/i0_4 ), .A2(\SB1_4_5/i1[9] ), .A3(
        \SB1_4_5/i0_3 ), .ZN(n7386) );
  NAND3_X1 U14571 ( .A1(\SB4_5/i0_4 ), .A2(\SB4_5/i1[9] ), .A3(\SB4_5/i1_5 ), 
        .ZN(n7387) );
  NAND3_X1 U14572 ( .A1(\SB1_4_12/i0[8] ), .A2(\RI1[4][119] ), .A3(
        \SB1_4_12/i1_7 ), .ZN(\SB1_4_12/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U14573 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[141] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[147] ), .Z(n7389) );
  NAND2_X1 U14574 ( .A1(\SB4_19/i1_7 ), .A2(\SB4_19/i0[8] ), .ZN(n7390) );
  NAND4_X2 U14575 ( .A1(\SB2_2_8/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_8/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_2_8/Component_Function_1/NAND4_in[2] ), .A4(n7391), .ZN(
        \SB2_2_8/buf_output[1] ) );
  NAND3_X1 U14576 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i0[9] ), .A3(
        \SB3_26/buf_output[3] ), .ZN(n5026) );
  XOR2_X1 U14577 ( .A1(n1818), .A2(n7393), .Z(\MC_ARK_ARC_1_1/buf_output[82] )
         );
  XOR2_X1 U14578 ( .A1(\MC_ARK_ARC_1_1/temp3[82] ), .A2(
        \MC_ARK_ARC_1_1/temp4[82] ), .Z(n7393) );
  XOR2_X1 U14579 ( .A1(\RI5[2][138] ), .A2(\RI5[2][132] ), .Z(n7394) );
  XOR2_X1 U14580 ( .A1(n7395), .A2(n105), .Z(Ciphertext[169]) );
  XOR2_X1 U14581 ( .A1(n7589), .A2(\MC_ARK_ARC_1_4/temp6[165] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[165] ) );
  NAND3_X1 U14582 ( .A1(\SB3_31/i0[6] ), .A2(\SB3_31/i0[7] ), .A3(
        \SB3_31/i0[8] ), .ZN(\SB3_31/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U14583 ( .A1(\SB1_1_14/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_14/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_14/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_1_14/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_14/buf_output[0] ) );
  NAND4_X2 U14584 ( .A1(\SB2_3_1/Component_Function_2/NAND4_in[2] ), .A2(n7518), .A3(\SB2_3_1/Component_Function_2/NAND4_in[0] ), .A4(n7396), .ZN(
        \SB2_3_1/buf_output[2] ) );
  NAND3_X2 U14585 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i0[10] ), .A3(
        \SB2_3_1/i0[6] ), .ZN(n7396) );
  NAND4_X2 U14586 ( .A1(\SB2_2_5/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_5/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_5/Component_Function_2/NAND4_in[3] ), .A4(n7397), .ZN(
        \SB2_2_5/buf_output[2] ) );
  NAND3_X2 U14587 ( .A1(\SB2_2_5/i0[10] ), .A2(\SB2_2_5/i1_5 ), .A3(
        \SB2_2_5/i1[9] ), .ZN(n7397) );
  XOR2_X1 U14588 ( .A1(n7398), .A2(n199), .Z(Ciphertext[34]) );
  NAND4_X2 U14589 ( .A1(n2882), .A2(n2938), .A3(
        \SB4_26/Component_Function_4/NAND4_in[0] ), .A4(
        \SB4_26/Component_Function_4/NAND4_in[1] ), .ZN(n7398) );
  XOR2_X1 U14590 ( .A1(n2292), .A2(n7399), .Z(\MC_ARK_ARC_1_3/buf_output[55] )
         );
  XOR2_X1 U14591 ( .A1(\MC_ARK_ARC_1_3/temp4[55] ), .A2(
        \MC_ARK_ARC_1_3/temp3[55] ), .Z(n7399) );
  INV_X2 U14592 ( .I(\RI3[0][140] ), .ZN(\SB2_0_8/i1[9] ) );
  XOR2_X1 U14593 ( .A1(\MC_ARK_ARC_1_1/temp6[11] ), .A2(n4943), .Z(
        \MC_ARK_ARC_1_1/buf_output[11] ) );
  NAND4_X2 U14594 ( .A1(\SB1_2_30/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_30/Component_Function_0/NAND4_in[0] ), .A4(n7400), .ZN(
        \SB1_2_30/buf_output[0] ) );
  NAND3_X1 U14595 ( .A1(\SB1_4_9/i1[9] ), .A2(\SB1_4_9/i0[10] ), .A3(
        \SB1_4_9/i1_7 ), .ZN(\SB1_4_9/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U14596 ( .A1(\MC_ARK_ARC_1_4/temp3[96] ), .A2(
        \MC_ARK_ARC_1_4/temp4[96] ), .Z(\MC_ARK_ARC_1_4/temp6[96] ) );
  NAND3_X1 U14597 ( .A1(\SB2_0_8/i0_0 ), .A2(\SB2_0_8/i0[8] ), .A3(
        \SB2_0_8/i0[9] ), .ZN(n7401) );
  NAND4_X2 U14598 ( .A1(\SB1_1_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_5/NAND4_in[0] ), .A4(n7402), .ZN(
        \SB1_1_13/buf_output[5] ) );
  NAND3_X2 U14599 ( .A1(\SB1_1_13/i0_4 ), .A2(\SB1_1_13/i0[6] ), .A3(
        \SB1_1_13/i0[9] ), .ZN(n7402) );
  NAND3_X2 U14600 ( .A1(\SB1_2_16/i0[8] ), .A2(\SB1_2_16/i3[0] ), .A3(
        \SB1_2_16/i1_5 ), .ZN(n3812) );
  XOR2_X1 U14601 ( .A1(\MC_ARK_ARC_1_1/temp4[99] ), .A2(n7403), .Z(
        \MC_ARK_ARC_1_1/temp6[99] ) );
  XOR2_X1 U14602 ( .A1(\RI5[1][9] ), .A2(\RI5[1][165] ), .Z(n7403) );
  NAND3_X1 U14603 ( .A1(\SB4_31/i0_3 ), .A2(\SB4_31/i0_0 ), .A3(\SB4_31/i0[7] ), .ZN(n7404) );
  NAND3_X2 U14604 ( .A1(\SB1_2_27/i0_0 ), .A2(\SB1_2_27/i0[6] ), .A3(
        \SB1_2_27/i0[10] ), .ZN(n7405) );
  NAND3_X1 U14605 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i0_3 ), .A3(\SB4_13/i0_4 ), 
        .ZN(n4284) );
  XOR2_X1 U14606 ( .A1(\MC_ARK_ARC_1_0/temp5[103] ), .A2(n7406), .Z(
        \MC_ARK_ARC_1_0/buf_output[103] ) );
  XOR2_X1 U14607 ( .A1(\MC_ARK_ARC_1_0/temp3[103] ), .A2(
        \MC_ARK_ARC_1_0/temp4[103] ), .Z(n7406) );
  INV_X2 U14608 ( .I(\SB1_2_26/buf_output[5] ), .ZN(\SB2_2_26/i1_5 ) );
  XOR2_X1 U14609 ( .A1(\MC_ARK_ARC_1_0/temp1[143] ), .A2(n7407), .Z(n861) );
  XOR2_X1 U14610 ( .A1(\RI5[0][89] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[113] ), 
        .Z(n7407) );
  XOR2_X1 U14611 ( .A1(\RI5[2][113] ), .A2(\RI5[2][137] ), .Z(n7408) );
  NAND3_X2 U14612 ( .A1(\SB2_1_16/i0[9] ), .A2(\SB2_1_16/i0_4 ), .A3(
        \SB2_1_16/i0[6] ), .ZN(n7409) );
  XOR2_X1 U14613 ( .A1(n7410), .A2(n133), .Z(Ciphertext[129]) );
  XOR2_X1 U14614 ( .A1(\RI5[3][134] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[140] ), .Z(\MC_ARK_ARC_1_3/temp1[140] ) );
  NAND4_X2 U14615 ( .A1(\SB2_0_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_22/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_0_22/Component_Function_4/NAND4_in[1] ), .A4(n7411), .ZN(
        \SB2_0_22/buf_output[4] ) );
  NAND3_X2 U14616 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0[9] ), .A3(
        \SB2_0_22/i0[10] ), .ZN(n7411) );
  NAND3_X2 U14617 ( .A1(\SB1_3_7/i0_0 ), .A2(\SB1_3_7/i0[10] ), .A3(
        \SB1_3_7/i0[6] ), .ZN(\SB1_3_7/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U14618 ( .A1(n7413), .A2(n3103), .Z(\MC_ARK_ARC_1_0/buf_output[57] )
         );
  XOR2_X1 U14619 ( .A1(n1882), .A2(\MC_ARK_ARC_1_2/temp6[70] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[70] ) );
  NAND3_X1 U14620 ( .A1(\SB4_18/i0[9] ), .A2(\SB4_18/i0_0 ), .A3(
        \SB4_18/i0[8] ), .ZN(n7416) );
  NAND4_X2 U14621 ( .A1(\SB2_4_9/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_4_9/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_4_9/Component_Function_4/NAND4_in[2] ), .A4(n7417), .ZN(
        \SB2_4_9/buf_output[4] ) );
  NAND3_X1 U14622 ( .A1(\SB2_4_9/i0_4 ), .A2(\SB2_4_9/i1[9] ), .A3(
        \SB2_4_9/i1_5 ), .ZN(n7417) );
  NAND3_X1 U14623 ( .A1(\SB4_21/i0[10] ), .A2(\SB4_21/i0_3 ), .A3(
        \SB4_21/i0_4 ), .ZN(\SB4_21/Component_Function_0/NAND4_in[2] ) );
  INV_X1 U14624 ( .I(\SB3_29/buf_output[3] ), .ZN(\SB4_27/i0[8] ) );
  XOR2_X1 U14625 ( .A1(\RI5[4][107] ), .A2(\RI5[4][101] ), .Z(n7419) );
  INV_X1 U14626 ( .I(\SB1_1_19/buf_output[1] ), .ZN(\SB2_1_15/i1_7 ) );
  NAND4_X2 U14627 ( .A1(\SB1_1_19/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_1_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_1_19/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_1_19/buf_output[1] ) );
  NAND4_X2 U14628 ( .A1(\SB1_0_1/Component_Function_5/NAND4_in[1] ), .A2(n4575), .A3(\SB1_0_1/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_1/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_0_1/buf_output[5] ) );
  XOR2_X1 U14629 ( .A1(\MC_ARK_ARC_1_3/temp1[42] ), .A2(n7420), .Z(n7490) );
  XOR2_X1 U14630 ( .A1(\RI5[3][180] ), .A2(\RI5[3][12] ), .Z(n7420) );
  NAND3_X1 U14631 ( .A1(\SB2_4_3/i0[6] ), .A2(\SB2_4_3/i0[9] ), .A3(
        \SB1_4_4/buf_output[4] ), .ZN(
        \SB2_4_3/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U14632 ( .A1(n7422), .A2(n7421), .Z(\MC_ARK_ARC_1_0/buf_output[173] ) );
  NAND3_X2 U14633 ( .A1(\SB2_4_9/i0[9] ), .A2(\SB2_4_9/i0_4 ), .A3(
        \SB2_4_9/i0[6] ), .ZN(n7424) );
  NAND3_X1 U14634 ( .A1(\SB1_4_10/i0_0 ), .A2(\SB1_4_10/i1_7 ), .A3(
        \SB1_4_10/i3[0] ), .ZN(n7425) );
  NAND4_X2 U14635 ( .A1(\SB2_4_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_4_1/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_4_1/Component_Function_3/NAND4_in[1] ), .A4(n7426), .ZN(
        \SB2_4_1/buf_output[3] ) );
  NAND3_X2 U14636 ( .A1(\SB3_25/i0[6] ), .A2(\SB3_25/i0_4 ), .A3(
        \SB3_25/i0[9] ), .ZN(n7429) );
  XOR2_X1 U14637 ( .A1(\MC_ARK_ARC_1_1/temp5[144] ), .A2(n7430), .Z(
        \MC_ARK_ARC_1_1/buf_output[144] ) );
  XOR2_X1 U14638 ( .A1(\MC_ARK_ARC_1_1/temp4[144] ), .A2(n4712), .Z(n7430) );
  NAND4_X2 U14639 ( .A1(\SB1_4_18/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_4_18/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_4_18/Component_Function_4/NAND4_in[3] ), .A4(n7431), .ZN(
        \SB1_4_18/buf_output[4] ) );
  XOR2_X1 U14640 ( .A1(n1853), .A2(n7432), .Z(\MC_ARK_ARC_1_1/buf_output[41] )
         );
  XOR2_X1 U14641 ( .A1(n3486), .A2(\MC_ARK_ARC_1_1/temp2[41] ), .Z(n7432) );
  NAND4_X2 U14642 ( .A1(\SB2_0_21/Component_Function_2/NAND4_in[0] ), .A2(
        n7433), .A3(\SB2_0_21/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_21/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_0_21/buf_output[2] ) );
  NAND4_X2 U14643 ( .A1(\SB2_1_30/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_30/Component_Function_0/NAND4_in[0] ), .A4(n7434), .ZN(
        \SB2_1_30/buf_output[0] ) );
  NAND3_X2 U14644 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i0_0 ), .A3(
        \SB2_1_30/i0[7] ), .ZN(n7434) );
  NAND3_X2 U14645 ( .A1(\SB2_0_21/i0_0 ), .A2(\SB2_0_21/i0_4 ), .A3(
        \SB2_0_21/i0_3 ), .ZN(\SB2_0_21/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U14646 ( .A1(\RI5[2][95] ), .A2(\RI5[2][71] ), .Z(n7435) );
  NAND3_X1 U14647 ( .A1(\SB2_4_9/i0_0 ), .A2(\SB2_4_9/i0_4 ), .A3(
        \SB2_4_9/i1_5 ), .ZN(n1799) );
  XOR2_X1 U14648 ( .A1(\RI5[1][89] ), .A2(\RI5[1][113] ), .Z(
        \MC_ARK_ARC_1_1/temp2[143] ) );
  XOR2_X1 U14649 ( .A1(\MC_ARK_ARC_1_1/temp6[139] ), .A2(
        \MC_ARK_ARC_1_1/temp5[139] ), .Z(\MC_ARK_ARC_1_1/buf_output[139] ) );
  XOR2_X1 U14650 ( .A1(\RI5[4][85] ), .A2(\RI5[4][91] ), .Z(n7436) );
  XOR2_X1 U14651 ( .A1(\MC_ARK_ARC_1_4/temp4[179] ), .A2(n4037), .Z(n3145) );
  NAND4_X2 U14652 ( .A1(\SB4_12/Component_Function_1/NAND4_in[1] ), .A2(n1287), 
        .A3(\SB4_12/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_12/Component_Function_1/NAND4_in[2] ), .ZN(n7449) );
  XOR2_X1 U14653 ( .A1(\MC_ARK_ARC_1_0/temp1[122] ), .A2(
        \MC_ARK_ARC_1_0/temp2[122] ), .Z(\MC_ARK_ARC_1_0/temp5[122] ) );
  XOR2_X1 U14654 ( .A1(\MC_ARK_ARC_1_0/temp5[23] ), .A2(n2422), .Z(
        \RI1[1][23] ) );
  XOR2_X1 U14655 ( .A1(\MC_ARK_ARC_1_1/temp5[163] ), .A2(
        \MC_ARK_ARC_1_1/temp6[163] ), .Z(\MC_ARK_ARC_1_1/buf_output[163] ) );
  XOR2_X1 U14656 ( .A1(\MC_ARK_ARC_1_1/temp6[99] ), .A2(
        \MC_ARK_ARC_1_1/temp5[99] ), .Z(\MC_ARK_ARC_1_1/buf_output[99] ) );
  XOR2_X1 U14657 ( .A1(\MC_ARK_ARC_1_2/temp5[172] ), .A2(
        \MC_ARK_ARC_1_2/temp6[172] ), .Z(\MC_ARK_ARC_1_2/buf_output[172] ) );
  NAND4_X2 U14658 ( .A1(\SB2_1_31/Component_Function_3/NAND4_in[3] ), .A2(
        n7443), .A3(\SB2_1_31/Component_Function_3/NAND4_in[2] ), .A4(n2266), 
        .ZN(\SB2_1_31/buf_output[3] ) );
  XOR2_X1 U14659 ( .A1(\MC_ARK_ARC_1_4/temp6[176] ), .A2(n7437), .Z(
        \MC_ARK_ARC_1_4/buf_output[176] ) );
  NAND4_X2 U14660 ( .A1(\SB2_1_29/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_29/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_1_29/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_29/buf_output[1] ) );
  NAND4_X2 U14661 ( .A1(\SB2_3_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_14/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_3_14/Component_Function_3/NAND4_in[1] ), .A4(n7438), .ZN(
        \SB2_3_14/buf_output[3] ) );
  NAND3_X2 U14662 ( .A1(\SB2_3_14/i0[10] ), .A2(\SB2_3_14/i1[9] ), .A3(
        \SB2_3_14/i1_7 ), .ZN(n7438) );
  NAND3_X1 U14663 ( .A1(\SB3_29/i0_0 ), .A2(\SB3_29/i0[10] ), .A3(
        \SB3_29/i0[6] ), .ZN(\SB3_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U14664 ( .A1(\SB4_29/i0_3 ), .A2(\SB4_29/i0[6] ), .A3(
        \SB4_29/i1[9] ), .ZN(n1029) );
  XOR2_X1 U14665 ( .A1(\RI5[0][83] ), .A2(\RI5[0][89] ), .Z(
        \MC_ARK_ARC_1_0/temp1[89] ) );
  XOR2_X1 U14666 ( .A1(\MC_ARK_ARC_1_0/temp5[53] ), .A2(n7439), .Z(
        \MC_ARK_ARC_1_0/buf_output[53] ) );
  XOR2_X1 U14667 ( .A1(\MC_ARK_ARC_1_0/temp4[53] ), .A2(
        \MC_ARK_ARC_1_0/temp3[53] ), .Z(n7439) );
  XOR2_X1 U14668 ( .A1(n5231), .A2(n7440), .Z(\MC_ARK_ARC_1_1/buf_output[71] )
         );
  XOR2_X1 U14669 ( .A1(n2263), .A2(\MC_ARK_ARC_1_1/temp4[71] ), .Z(n7440) );
  XOR2_X1 U14670 ( .A1(n7441), .A2(n3532), .Z(\MC_ARK_ARC_1_3/buf_output[77] )
         );
  XOR2_X1 U14671 ( .A1(\MC_ARK_ARC_1_3/temp4[77] ), .A2(n2741), .Z(n7441) );
  INV_X2 U14672 ( .I(\SB1_4_19/buf_output[2] ), .ZN(\SB2_4_16/i1[9] ) );
  NAND3_X2 U14673 ( .A1(\SB2_0_15/i3[0] ), .A2(\SB2_0_15/i1_5 ), .A3(
        \SB2_0_15/i0[8] ), .ZN(\SB2_0_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U14674 ( .A1(\SB2_1_31/i0[6] ), .A2(\SB2_1_31/i1[9] ), .A3(
        \SB2_1_31/i0_3 ), .ZN(n7443) );
  NAND3_X2 U14675 ( .A1(\SB2_3_4/i0_0 ), .A2(\SB2_3_4/i0[10] ), .A3(
        \SB2_3_4/i0[6] ), .ZN(n7444) );
  XOR2_X1 U14676 ( .A1(n7445), .A2(n60), .Z(Ciphertext[37]) );
  NAND4_X2 U14677 ( .A1(\SB4_25/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_25/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_25/Component_Function_1/NAND4_in[1] ), .A4(n946), .ZN(n7445) );
  NAND4_X2 U14678 ( .A1(\SB2_4_25/Component_Function_0/NAND4_in[1] ), .A2(
        n2606), .A3(\SB2_4_25/Component_Function_0/NAND4_in[0] ), .A4(n7446), 
        .ZN(\SB2_4_25/buf_output[0] ) );
  NAND3_X2 U14679 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i0[6] ), .A3(
        \SB1_0_2/i1[9] ), .ZN(\SB1_0_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U14680 ( .A1(\SB1_0_3/i0[10] ), .A2(\SB1_0_3/i0_3 ), .A3(
        \SB1_0_3/i0[6] ), .ZN(n7447) );
  NAND3_X2 U14681 ( .A1(n851), .A2(\SB2_3_10/i1[9] ), .A3(\SB2_3_10/i0_3 ), 
        .ZN(\SB2_3_10/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U14682 ( .A1(\MC_ARK_ARC_1_3/temp5[29] ), .A2(n7448), .Z(
        \MC_ARK_ARC_1_3/buf_output[29] ) );
  XOR2_X1 U14683 ( .A1(\MC_ARK_ARC_1_3/temp3[29] ), .A2(
        \MC_ARK_ARC_1_3/temp4[29] ), .Z(n7448) );
  XOR2_X1 U14684 ( .A1(n7449), .A2(n192), .Z(Ciphertext[115]) );
  NAND4_X2 U14685 ( .A1(n1609), .A2(n4901), .A3(
        \SB2_2_20/Component_Function_2/NAND4_in[2] ), .A4(n7450), .ZN(
        \SB2_2_20/buf_output[2] ) );
  NAND3_X2 U14686 ( .A1(\SB2_2_20/i0[10] ), .A2(\SB2_2_20/i1_5 ), .A3(
        \SB2_2_20/i1[9] ), .ZN(n7450) );
  XOR2_X1 U14687 ( .A1(\RI5[2][104] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[68] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[2] ) );
  NAND3_X1 U14688 ( .A1(\SB1_4_4/i0_3 ), .A2(\SB1_4_4/i1[9] ), .A3(
        \SB1_4_4/i0[6] ), .ZN(\SB1_4_4/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U14689 ( .A1(\SB3_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_27/Component_Function_2/NAND4_in[1] ), .A3(n7512), .A4(n7452), 
        .ZN(\SB3_27/buf_output[2] ) );
  XOR2_X1 U14690 ( .A1(\MC_ARK_ARC_1_2/temp2[78] ), .A2(
        \MC_ARK_ARC_1_2/temp1[78] ), .Z(n1967) );
  NAND3_X2 U14691 ( .A1(\SB2_2_3/i0_4 ), .A2(n3994), .A3(\SB2_2_3/i0_0 ), .ZN(
        n687) );
  NAND4_X2 U14692 ( .A1(\SB2_0_16/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_0_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_16/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_16/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_0_16/buf_output[1] ) );
  XOR2_X1 U14693 ( .A1(n4113), .A2(n4112), .Z(\MC_ARK_ARC_1_4/buf_output[191] ) );
  XOR2_X1 U14694 ( .A1(\MC_ARK_ARC_1_0/temp2[125] ), .A2(
        \MC_ARK_ARC_1_0/temp1[125] ), .Z(n1957) );
  XOR2_X1 U14695 ( .A1(n1856), .A2(\MC_ARK_ARC_1_1/temp4[29] ), .Z(n1935) );
  NAND4_X2 U14696 ( .A1(\SB2_2_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_24/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_24/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_2_24/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_24/buf_output[2] ) );
  NAND4_X2 U14697 ( .A1(\SB1_0_21/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_21/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_21/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_0_21/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_0_21/buf_output[3] ) );
  NAND4_X2 U14698 ( .A1(\SB1_3_4/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_4/Component_Function_2/NAND4_in[0] ), .A3(n7545), .A4(n4414), 
        .ZN(\SB1_3_4/buf_output[2] ) );
  XOR2_X1 U14699 ( .A1(\RI5[1][63] ), .A2(\RI5[1][39] ), .Z(
        \MC_ARK_ARC_1_1/temp2[93] ) );
  NAND3_X2 U14700 ( .A1(\SB2_3_1/i0[10] ), .A2(\SB2_3_1/i1[9] ), .A3(
        \SB2_3_1/i1_5 ), .ZN(\SB2_3_1/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U14701 ( .A1(\SB1_1_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_1_5/Component_Function_3/NAND4_in[1] ), .A4(n7453), .ZN(
        \SB1_1_5/buf_output[3] ) );
  XOR2_X1 U14702 ( .A1(\MC_ARK_ARC_1_2/temp5[47] ), .A2(n1355), .Z(
        \MC_ARK_ARC_1_2/buf_output[47] ) );
  NAND4_X2 U14703 ( .A1(\SB3_23/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_23/Component_Function_5/NAND4_in[2] ), .A3(
        \SB3_23/Component_Function_5/NAND4_in[3] ), .A4(
        \SB3_23/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_23/buf_output[5] ) );
  NAND3_X2 U14704 ( .A1(\SB2_2_1/i0[10] ), .A2(\SB2_2_1/i1_5 ), .A3(
        \SB2_2_1/i1[9] ), .ZN(\SB2_2_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U14705 ( .A1(\SB1_1_10/i0_0 ), .A2(\SB1_1_10/i0_4 ), .A3(
        \SB1_1_10/i1_5 ), .ZN(n7454) );
  OAI21_X2 U14706 ( .A1(n5435), .A2(n5436), .B(\SB1_0_10/i0[10] ), .ZN(n7489)
         );
  NAND3_X2 U14707 ( .A1(\SB1_1_17/i0[10] ), .A2(\SB1_1_17/i1[9] ), .A3(
        \SB1_1_17/i1_5 ), .ZN(n7572) );
  NAND3_X1 U14708 ( .A1(\SB3_15/i0[9] ), .A2(\SB3_15/i0[8] ), .A3(
        \SB3_15/i0_0 ), .ZN(\SB3_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U14709 ( .A1(\SB3_15/i0[9] ), .A2(\SB3_15/i0[6] ), .A3(
        \SB3_15/i0_4 ), .ZN(n2665) );
  XOR2_X1 U14710 ( .A1(\RI5[2][127] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[151] ), .Z(\MC_ARK_ARC_1_2/temp2[181] ) );
  XOR2_X1 U14711 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[129] ), .A2(\RI5[3][153] ), .Z(n7457) );
  XOR2_X1 U14712 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[177] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[183] ), .Z(n7458) );
  NAND3_X2 U14713 ( .A1(\SB1_1_2/i1[9] ), .A2(\SB1_1_2/i0_3 ), .A3(
        \SB1_1_2/i0[6] ), .ZN(\SB1_1_2/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U14714 ( .A1(\RI5[0][11] ), .A2(\RI5[0][179] ), .Z(n7459) );
  NAND3_X2 U14715 ( .A1(\SB2_1_11/i0[10] ), .A2(\SB2_1_11/i1[9] ), .A3(
        \SB2_1_11/i1_7 ), .ZN(\SB2_1_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U14716 ( .A1(\SB1_2_7/i0[10] ), .A2(\RI1[2][149] ), .A3(
        \SB1_2_7/i0[6] ), .ZN(\SB1_2_7/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U14717 ( .A1(n1861), .A2(\SB2_1_1/Component_Function_3/NAND4_in[0] ), .A3(\SB2_1_1/Component_Function_3/NAND4_in[3] ), .A4(n4597), .ZN(
        \SB2_1_1/buf_output[3] ) );
  NAND4_X2 U14718 ( .A1(\SB1_0_12/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_12/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_12/Component_Function_3/NAND4_in[0] ), .A4(n4748), .ZN(
        \RI3[0][129] ) );
  XOR2_X1 U14719 ( .A1(n7461), .A2(n7460), .Z(n2858) );
  XOR2_X1 U14720 ( .A1(\RI5[0][40] ), .A2(n204), .Z(n7460) );
  XOR2_X1 U14721 ( .A1(\RI5[0][10] ), .A2(\RI5[0][76] ), .Z(n7461) );
  XOR2_X1 U14722 ( .A1(n3921), .A2(\MC_ARK_ARC_1_1/temp1[179] ), .Z(n7463) );
  NAND4_X2 U14723 ( .A1(\SB2_2_14/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_14/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_2_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_14/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_14/buf_output[0] ) );
  NAND3_X1 U14724 ( .A1(\SB1_3_9/i0_0 ), .A2(n3979), .A3(\SB1_3_9/i0[8] ), 
        .ZN(\SB1_3_9/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U14725 ( .A1(\MC_ARK_ARC_1_2/temp5[132] ), .A2(
        \MC_ARK_ARC_1_2/temp6[132] ), .Z(n3979) );
  XOR2_X1 U14726 ( .A1(\MC_ARK_ARC_1_3/temp4[180] ), .A2(
        \MC_ARK_ARC_1_3/temp1[180] ), .Z(n7465) );
  XOR2_X1 U14727 ( .A1(n7466), .A2(n35), .Z(Ciphertext[179]) );
  NAND4_X2 U14728 ( .A1(\SB1_2_0/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_2_0/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_2_0/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_2_0/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB1_2_0/buf_output[3] ) );
  XOR2_X1 U14729 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[83] ), .A2(\RI5[1][107] ), 
        .Z(n4385) );
  NAND3_X1 U14730 ( .A1(\SB1_2_17/i0_4 ), .A2(\SB1_2_17/i0[10] ), .A3(
        \SB1_2_17/i0_3 ), .ZN(n7467) );
  NAND3_X1 U14731 ( .A1(\SB3_15/buf_output[2] ), .A2(\SB4_12/i1_7 ), .A3(
        \SB4_12/i3[0] ), .ZN(\SB4_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U14732 ( .A1(\SB2_1_11/i0[6] ), .A2(\SB2_1_11/i0[9] ), .A3(
        \SB2_1_11/i0_4 ), .ZN(n7469) );
  INV_X1 U14733 ( .I(\RI3[5][149] ), .ZN(\SB4_7/i1_5 ) );
  NAND4_X2 U14734 ( .A1(\SB3_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_7/Component_Function_5/NAND4_in[3] ), .A3(n1594), .A4(
        \SB3_7/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[5][149] ) );
  NAND3_X2 U14735 ( .A1(\SB2_2_1/i0[10] ), .A2(\SB2_2_1/i0_3 ), .A3(
        \SB1_2_2/buf_output[4] ), .ZN(
        \SB2_2_1/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U14736 ( .A1(\RI5[2][156] ), .A2(\RI5[2][180] ), .Z(n7470) );
  NAND3_X1 U14737 ( .A1(\SB2_2_13/i0_3 ), .A2(\SB2_2_13/i0[6] ), .A3(
        \SB2_2_13/i1[9] ), .ZN(\SB2_2_13/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U14738 ( .A1(\MC_ARK_ARC_1_1/temp2[185] ), .A2(n7471), .Z(n3198) );
  XOR2_X1 U14739 ( .A1(\RI5[1][179] ), .A2(\RI5[1][185] ), .Z(n7471) );
  XOR2_X1 U14740 ( .A1(\MC_ARK_ARC_1_4/buf_datainput[94] ), .A2(
        \MC_ARK_ARC_1_4/buf_datainput[118] ), .Z(\MC_ARK_ARC_1_4/temp2[148] )
         );
  XOR2_X1 U14741 ( .A1(n7472), .A2(n3064), .Z(\MC_ARK_ARC_1_2/buf_output[87] )
         );
  XOR2_X1 U14742 ( .A1(\RI5[2][138] ), .A2(\RI5[2][114] ), .Z(
        \MC_ARK_ARC_1_2/temp2[168] ) );
  NAND3_X2 U14743 ( .A1(\SB2_2_10/i0_0 ), .A2(\SB2_2_10/i0[7] ), .A3(
        \SB2_2_10/i0_3 ), .ZN(\SB2_2_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U14744 ( .A1(\SB1_1_5/i0[10] ), .A2(\SB1_1_5/i1_5 ), .A3(
        \SB1_1_5/i1[9] ), .ZN(n7474) );
  NAND4_X2 U14745 ( .A1(\SB2_4_1/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_4_1/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_4_1/Component_Function_2/NAND4_in[0] ), .A4(n7473), .ZN(
        \SB2_4_1/buf_output[2] ) );
  NAND3_X2 U14746 ( .A1(\SB2_4_1/i0[10] ), .A2(\SB2_4_1/i0_3 ), .A3(
        \SB2_4_1/i0[6] ), .ZN(n7473) );
  NAND3_X2 U14747 ( .A1(\SB1_0_5/i0[10] ), .A2(\SB1_0_5/i1[9] ), .A3(
        \SB1_0_5/i1_7 ), .ZN(n7475) );
  XOR2_X1 U14748 ( .A1(\MC_ARK_ARC_1_3/temp3[79] ), .A2(
        \MC_ARK_ARC_1_3/temp4[79] ), .Z(\MC_ARK_ARC_1_3/temp6[79] ) );
  XOR2_X1 U14749 ( .A1(n7476), .A2(n117), .Z(Ciphertext[75]) );
  XOR2_X1 U14750 ( .A1(\MC_ARK_ARC_1_3/temp1[43] ), .A2(
        \MC_ARK_ARC_1_3/temp2[43] ), .Z(n7477) );
  NAND3_X1 U14751 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB2_3_7/i0[8] ), .A3(
        \SB2_3_7/i1_7 ), .ZN(\SB2_3_7/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U14752 ( .A1(\MC_ARK_ARC_1_4/temp4[15] ), .A2(n1128), .Z(n1534) );
  XOR2_X1 U14753 ( .A1(n3302), .A2(n3301), .Z(\MC_ARK_ARC_1_0/buf_output[110] ) );
  XOR2_X1 U14754 ( .A1(\RI5[2][69] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[63] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[69] ) );
  XOR2_X1 U14755 ( .A1(\RI5[0][80] ), .A2(\RI5[0][56] ), .Z(
        \MC_ARK_ARC_1_0/temp2[110] ) );
  XOR2_X1 U14756 ( .A1(n1720), .A2(n7479), .Z(\MC_ARK_ARC_1_4/buf_output[95] )
         );
  XOR2_X1 U14757 ( .A1(n7519), .A2(\MC_ARK_ARC_1_4/temp4[95] ), .Z(n7479) );
  NAND4_X2 U14758 ( .A1(n4483), .A2(\SB1_4_3/Component_Function_1/NAND4_in[1] ), .A3(\SB1_4_3/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_4_3/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_4_3/buf_output[1] ) );
  XOR2_X1 U14759 ( .A1(\MC_ARK_ARC_1_0/temp2[52] ), .A2(n7480), .Z(n4882) );
  XOR2_X1 U14760 ( .A1(\RI5[0][46] ), .A2(\RI5[0][52] ), .Z(n7480) );
  AND2_X1 U14761 ( .A1(n2011), .A2(\SB3_25/Component_Function_3/NAND4_in[2] ), 
        .Z(n3385) );
  NAND3_X1 U14762 ( .A1(\SB3_18/i1[9] ), .A2(\SB3_18/i0[10] ), .A3(
        \SB3_18/i1_5 ), .ZN(\SB3_18/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U14763 ( .A1(n3485), .A2(n7482), .Z(\RI1[5][41] ) );
  XOR2_X1 U14764 ( .A1(\MC_ARK_ARC_1_4/temp4[41] ), .A2(
        \MC_ARK_ARC_1_4/temp3[41] ), .Z(n7482) );
  XOR2_X1 U14765 ( .A1(\MC_ARK_ARC_1_3/temp5[98] ), .A2(n7483), .Z(
        \MC_ARK_ARC_1_3/buf_output[98] ) );
  XOR2_X1 U14766 ( .A1(\MC_ARK_ARC_1_3/temp4[98] ), .A2(n5067), .Z(n7483) );
  XOR2_X1 U14767 ( .A1(\MC_ARK_ARC_1_0/temp2[45] ), .A2(
        \MC_ARK_ARC_1_0/temp1[45] ), .Z(\MC_ARK_ARC_1_0/temp5[45] ) );
  NAND3_X1 U14768 ( .A1(\SB4_27/i0_3 ), .A2(\SB4_27/i0[8] ), .A3(\SB4_27/i1_7 ), .ZN(\SB4_27/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U14769 ( .A1(n5060), .A2(\MC_ARK_ARC_1_1/temp2[33] ), .Z(n7484) );
  XOR2_X1 U14770 ( .A1(\MC_ARK_ARC_1_3/temp6[128] ), .A2(
        \MC_ARK_ARC_1_3/temp5[128] ), .Z(\MC_ARK_ARC_1_3/buf_output[128] ) );
  NAND3_X2 U14771 ( .A1(\SB1_0_18/i0[10] ), .A2(\SB1_0_18/i1[9] ), .A3(
        \SB1_0_18/i1_7 ), .ZN(n7485) );
  NAND3_X2 U14772 ( .A1(\SB1_4_5/i0[10] ), .A2(\SB1_4_5/i1_7 ), .A3(
        \SB1_4_5/i1[9] ), .ZN(n2350) );
  NAND4_X2 U14773 ( .A1(n5364), .A2(
        \SB2_4_14/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_4_14/Component_Function_4/NAND4_in[1] ), .A4(n7486), .ZN(
        \SB2_4_14/buf_output[4] ) );
  NAND4_X2 U14774 ( .A1(\SB1_1_26/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_26/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_1_26/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_1_26/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_26/buf_output[4] ) );
  NAND3_X2 U14775 ( .A1(\SB2_4_10/i0[10] ), .A2(\SB2_4_10/i0_0 ), .A3(
        \SB2_4_10/i0[6] ), .ZN(n7487) );
  XOR2_X1 U14776 ( .A1(\MC_ARK_ARC_1_0/temp2[141] ), .A2(n3822), .Z(n1351) );
  XOR2_X1 U14777 ( .A1(\MC_ARK_ARC_1_2/temp5[86] ), .A2(n7488), .Z(
        \MC_ARK_ARC_1_2/buf_output[86] ) );
  XOR2_X1 U14778 ( .A1(\MC_ARK_ARC_1_2/temp3[86] ), .A2(
        \MC_ARK_ARC_1_2/temp4[86] ), .Z(n7488) );
  NAND4_X2 U14779 ( .A1(\SB2_0_22/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_22/Component_Function_1/NAND4_in[3] ), .A3(n3352), .A4(
        \SB2_0_22/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_22/buf_output[1] ) );
  NAND4_X2 U14780 ( .A1(n3322), .A2(
        \SB2_3_27/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_27/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_3_27/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_27/buf_output[0] ) );
  NAND4_X2 U14781 ( .A1(n3500), .A2(\SB2_3_7/Component_Function_4/NAND4_in[0] ), .A3(\SB2_3_7/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_7/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_3_7/buf_output[4] ) );
  NAND4_X2 U14782 ( .A1(\SB1_0_30/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_30/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_30/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_0_30/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_0_30/buf_output[1] ) );
  NAND2_X2 U14783 ( .A1(n1364), .A2(n7489), .ZN(\SB1_0_10/buf_output[2] ) );
  NAND4_X2 U14784 ( .A1(\SB1_0_8/Component_Function_5/NAND4_in[1] ), .A2(n2816), .A3(\SB1_0_8/Component_Function_5/NAND4_in[0] ), .A4(n2672), .ZN(
        \RI3[0][143] ) );
  XOR2_X1 U14785 ( .A1(n2340), .A2(n7490), .Z(\MC_ARK_ARC_1_3/buf_output[42] )
         );
  XOR2_X1 U14786 ( .A1(n7493), .A2(n181), .Z(Ciphertext[22]) );
  XOR2_X1 U14787 ( .A1(n7494), .A2(\MC_ARK_ARC_1_3/temp6[163] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[163] ) );
  XOR2_X1 U14788 ( .A1(n7495), .A2(\MC_ARK_ARC_1_4/temp6[1] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[1] ) );
  XOR2_X1 U14789 ( .A1(\MC_ARK_ARC_1_4/temp1[1] ), .A2(n3573), .Z(n7495) );
  NAND4_X2 U14790 ( .A1(n4960), .A2(
        \SB2_2_31/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_2_31/Component_Function_3/NAND4_in[1] ), .A4(n7496), .ZN(
        \SB2_2_31/buf_output[3] ) );
  NAND3_X2 U14791 ( .A1(\SB2_2_31/i0[6] ), .A2(\SB2_2_31/i0_3 ), .A3(
        \SB2_2_31/i1[9] ), .ZN(n7496) );
  NAND4_X2 U14792 ( .A1(n5237), .A2(n5303), .A3(
        \SB4_28/Component_Function_3/NAND4_in[2] ), .A4(n7497), .ZN(n4879) );
  NAND4_X2 U14793 ( .A1(\SB1_1_4/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_1_4/Component_Function_4/NAND4_in[1] ), .A3(n2660), .A4(n7498), 
        .ZN(\SB1_1_4/buf_output[4] ) );
  NAND3_X1 U14794 ( .A1(\MC_ARK_ARC_1_0/buf_output[166] ), .A2(\SB1_1_4/i1[9] ), .A3(\SB1_1_4/i1_5 ), .ZN(n7498) );
  NAND3_X1 U14795 ( .A1(\SB4_23/i0_3 ), .A2(n3974), .A3(\SB4_23/i1_7 ), .ZN(
        \SB4_23/Component_Function_1/NAND4_in[1] ) );
  NOR2_X2 U14796 ( .A1(n7500), .A2(n7499), .ZN(n3974) );
  NAND2_X2 U14797 ( .A1(\SB3_25/Component_Function_3/NAND4_in[2] ), .A2(n2011), 
        .ZN(n7499) );
  NAND3_X1 U14798 ( .A1(\SB1_2_3/i0_4 ), .A2(\SB1_2_3/i1_7 ), .A3(
        \SB1_2_3/i0[8] ), .ZN(\SB1_2_3/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U14799 ( .A1(n7501), .A2(\MC_ARK_ARC_1_3/temp6[108] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[108] ) );
  XOR2_X1 U14800 ( .A1(\MC_ARK_ARC_1_3/temp2[108] ), .A2(
        \MC_ARK_ARC_1_3/temp1[108] ), .Z(n7501) );
  NAND4_X2 U14801 ( .A1(n1242), .A2(\SB3_23/Component_Function_4/NAND4_in[1] ), 
        .A3(\SB3_23/Component_Function_4/NAND4_in[3] ), .A4(n7502), .ZN(
        \SB3_23/buf_output[4] ) );
  NAND3_X1 U14802 ( .A1(\SB3_23/i0[9] ), .A2(\SB3_23/i0_0 ), .A3(
        \SB3_23/i0[8] ), .ZN(n7502) );
  XOR2_X1 U14803 ( .A1(n7503), .A2(\MC_ARK_ARC_1_4/temp6[48] ), .Z(
        \MC_ARK_ARC_1_4/buf_output[48] ) );
  NAND3_X1 U14804 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i0_0 ), .A3(
        \SB1_2_13/i0_4 ), .ZN(\SB1_2_13/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U14805 ( .A1(\MC_ARK_ARC_1_1/temp3[117] ), .A2(
        \MC_ARK_ARC_1_1/temp4[117] ), .Z(n7504) );
  NAND3_X2 U14806 ( .A1(\SB2_1_8/i0_3 ), .A2(\SB2_1_8/i1[9] ), .A3(
        \SB2_1_8/i0[6] ), .ZN(\SB2_1_8/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U14807 ( .A1(\MC_ARK_ARC_1_3/temp5[23] ), .A2(
        \MC_ARK_ARC_1_3/temp6[23] ), .Z(\MC_ARK_ARC_1_3/buf_output[23] ) );
  XOR2_X1 U14808 ( .A1(n7505), .A2(n131), .Z(Ciphertext[65]) );
  NAND4_X2 U14809 ( .A1(\SB4_21/Component_Function_5/NAND4_in[1] ), .A2(n2860), 
        .A3(\SB4_21/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_21/Component_Function_5/NAND4_in[0] ), .ZN(n7505) );
  NAND3_X2 U14810 ( .A1(n5403), .A2(n5402), .A3(n7506), .ZN(
        \SB2_4_12/buf_output[5] ) );
  NAND3_X2 U14811 ( .A1(\SB2_4_12/i0_4 ), .A2(\SB2_4_12/i0_3 ), .A3(
        \SB2_4_12/i1[9] ), .ZN(n7506) );
  INV_X2 U14812 ( .I(\SB1_2_1/buf_output[5] ), .ZN(\SB2_2_1/i1_5 ) );
  XOR2_X1 U14813 ( .A1(n7507), .A2(n195), .Z(Ciphertext[64]) );
  NAND4_X2 U14814 ( .A1(\SB2_0_30/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_0_30/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_0_30/Component_Function_2/NAND4_in[1] ), .A4(n7508), .ZN(
        \SB2_0_30/buf_output[2] ) );
  XOR2_X1 U14815 ( .A1(\RI5[2][8] ), .A2(\RI5[2][170] ), .Z(n7509) );
  XOR2_X1 U14816 ( .A1(n2055), .A2(n2054), .Z(n5017) );
  XOR2_X1 U14817 ( .A1(\MC_ARK_ARC_1_0/temp3[147] ), .A2(
        \MC_ARK_ARC_1_0/temp4[147] ), .Z(\MC_ARK_ARC_1_0/temp6[147] ) );
  XOR2_X1 U14818 ( .A1(n7510), .A2(n212), .Z(Ciphertext[29]) );
  NAND4_X2 U14819 ( .A1(\SB4_27/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_27/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_27/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_27/Component_Function_5/NAND4_in[0] ), .ZN(n7510) );
  NAND3_X1 U14820 ( .A1(\SB3_16/i0[8] ), .A2(\SB3_16/i0_4 ), .A3(\SB3_16/i1_7 ), .ZN(\SB3_16/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U14821 ( .A1(\MC_ARK_ARC_1_2/temp6[11] ), .A2(n7511), .Z(
        \MC_ARK_ARC_1_2/buf_output[11] ) );
  XOR2_X1 U14822 ( .A1(\MC_ARK_ARC_1_2/temp2[11] ), .A2(n710), .Z(n7511) );
  NAND3_X2 U14823 ( .A1(\SB2_0_19/i0[8] ), .A2(\SB2_0_19/i0[9] ), .A3(
        \SB2_0_19/i0_0 ), .ZN(\SB2_0_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U14824 ( .A1(\SB1_1_20/i0[9] ), .A2(\SB1_1_20/i0_4 ), .A3(
        \SB1_1_20/i0[6] ), .ZN(n7513) );
  NAND3_X1 U14825 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i1[9] ), .A3(\SB4_2/i0[6] ), 
        .ZN(n7514) );
  NAND3_X1 U14826 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i0_0 ), .A3(
        \SB2_3_27/i0[7] ), .ZN(n3322) );
  NAND4_X2 U14827 ( .A1(n2620), .A2(n2286), .A3(
        \SB2_2_10/Component_Function_4/NAND4_in[1] ), .A4(n7516), .ZN(
        \SB2_2_10/buf_output[4] ) );
  NAND3_X2 U14828 ( .A1(\SB2_2_10/i0_0 ), .A2(\SB2_2_10/i0[9] ), .A3(
        \SB2_2_10/i0[8] ), .ZN(n7516) );
  XOR2_X1 U14829 ( .A1(\SB2_0_2/buf_output[0] ), .A2(\RI5[0][36] ), .Z(
        \MC_ARK_ARC_1_0/temp2[66] ) );
  NAND4_X2 U14830 ( .A1(\SB1_4_20/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_4_20/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_4_20/Component_Function_1/NAND4_in[0] ), .A4(n7517), .ZN(
        \SB1_4_20/buf_output[1] ) );
  NAND3_X1 U14831 ( .A1(\SB1_0_30/i0_4 ), .A2(\SB1_0_30/i0[10] ), .A3(
        \SB1_0_30/i0_3 ), .ZN(\SB1_0_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U14832 ( .A1(\SB2_3_1/i0_0 ), .A2(\SB2_3_1/i0_4 ), .A3(
        \SB2_3_1/i1_5 ), .ZN(n7518) );
  NAND3_X2 U14833 ( .A1(\SB1_4_25/i0[6] ), .A2(\SB1_4_25/i0[9] ), .A3(
        \SB1_4_25/i1_5 ), .ZN(n3698) );
  XOR2_X1 U14834 ( .A1(n7521), .A2(n7520), .Z(\MC_ARK_ARC_1_2/buf_output[116] ) );
  XOR2_X1 U14835 ( .A1(\MC_ARK_ARC_1_2/temp2[116] ), .A2(
        \MC_ARK_ARC_1_2/temp4[116] ), .Z(n7520) );
  XOR2_X1 U14836 ( .A1(\MC_ARK_ARC_1_2/temp1[116] ), .A2(
        \MC_ARK_ARC_1_2/temp3[116] ), .Z(n7521) );
  NAND3_X1 U14837 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0_0 ), .A3(n2748), .ZN(
        \SB2_2_1/Component_Function_0/NAND4_in[3] ) );
  NAND2_X2 U14838 ( .A1(n5255), .A2(n7523), .ZN(\SB2_3_10/i0_4 ) );
  XOR2_X1 U14839 ( .A1(\MC_ARK_ARC_1_0/temp5[65] ), .A2(n7524), .Z(
        \MC_ARK_ARC_1_0/buf_output[65] ) );
  XOR2_X1 U14840 ( .A1(n7525), .A2(\MC_ARK_ARC_1_0/temp2[176] ), .Z(
        \MC_ARK_ARC_1_0/temp5[176] ) );
  XOR2_X1 U14841 ( .A1(\RI5[0][176] ), .A2(\RI5[0][170] ), .Z(n7525) );
  NAND3_X1 U14842 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i0[6] ), .A3(
        \SB4_16/i1[9] ), .ZN(\SB4_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U14843 ( .A1(\SB2_1_7/i0_4 ), .A2(\SB2_1_7/i0[6] ), .A3(
        \SB2_1_7/i0[9] ), .ZN(n7585) );
  INV_X2 U14844 ( .I(\RI3[0][158] ), .ZN(\SB2_0_5/i1[9] ) );
  NAND4_X2 U14845 ( .A1(n1294), .A2(\SB1_0_8/Component_Function_2/NAND4_in[1] ), .A3(n5214), .A4(\SB1_0_8/Component_Function_2/NAND4_in[2] ), .ZN(
        \RI3[0][158] ) );
  NAND3_X1 U14846 ( .A1(\SB1_1_2/i1[9] ), .A2(\SB1_1_2/i0[10] ), .A3(
        \SB1_1_2/i1_7 ), .ZN(n2291) );
  NAND2_X2 U14847 ( .A1(n3169), .A2(n7528), .ZN(\SB2_2_23/i0_4 ) );
  AND2_X1 U14848 ( .A1(\SB1_2_24/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_24/Component_Function_4/NAND4_in[3] ), .Z(n7528) );
  NAND4_X2 U14849 ( .A1(\SB2_2_1/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_1/Component_Function_4/NAND4_in[1] ), .A3(n3672), .A4(n7529), 
        .ZN(\SB2_2_1/buf_output[4] ) );
  NAND3_X2 U14850 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0[10] ), .A3(
        \SB2_2_1/i0[9] ), .ZN(n7529) );
  XOR2_X1 U14851 ( .A1(\MC_ARK_ARC_1_2/temp1[69] ), .A2(n7530), .Z(
        \MC_ARK_ARC_1_2/temp5[69] ) );
  XOR2_X1 U14852 ( .A1(\RI5[2][39] ), .A2(\RI5[2][15] ), .Z(n7530) );
  NAND4_X2 U14853 ( .A1(\SB4_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_24/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_24/Component_Function_0/NAND4_in[0] ), .A4(n7531), .ZN(n2872) );
  NAND4_X2 U14854 ( .A1(\SB2_2_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_14/Component_Function_3/NAND4_in[1] ), .A3(n882), .A4(
        \SB2_2_14/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_14/buf_output[3] ) );
  XOR2_X1 U14855 ( .A1(\MC_ARK_ARC_1_3/temp5[69] ), .A2(n7532), .Z(
        \MC_ARK_ARC_1_3/buf_output[69] ) );
  NAND4_X2 U14856 ( .A1(\SB2_1_19/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_19/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_19/Component_Function_1/NAND4_in[0] ), .A4(n7533), .ZN(
        \SB2_1_19/buf_output[1] ) );
  XOR2_X1 U14857 ( .A1(n7534), .A2(n83), .Z(Ciphertext[90]) );
  NAND4_X2 U14858 ( .A1(\SB4_16/Component_Function_0/NAND4_in[2] ), .A2(n4957), 
        .A3(\SB4_16/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_16/Component_Function_0/NAND4_in[0] ), .ZN(n7534) );
  NAND3_X1 U14859 ( .A1(\SB3_29/i0[9] ), .A2(\RI1[5][17] ), .A3(\SB3_29/i0[8] ), .ZN(\SB3_29/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U14860 ( .A1(\MC_ARK_ARC_1_2/temp5[34] ), .A2(
        \MC_ARK_ARC_1_2/temp6[34] ), .Z(\MC_ARK_ARC_1_2/buf_output[34] ) );
  XOR2_X1 U14861 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[28] ), .A2(\RI5[2][34] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[34] ) );
  NAND3_X1 U14862 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i0[9] ), .A3(
        \SB4_14/i0[8] ), .ZN(n7536) );
  XOR2_X1 U14863 ( .A1(\MC_ARK_ARC_1_1/temp6[106] ), .A2(n7538), .Z(
        \MC_ARK_ARC_1_1/buf_output[106] ) );
  XOR2_X1 U14864 ( .A1(\MC_ARK_ARC_1_1/temp1[106] ), .A2(
        \MC_ARK_ARC_1_1/temp2[106] ), .Z(n7538) );
  XOR2_X1 U14865 ( .A1(\RI5[2][64] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[28] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[154] ) );
  NAND3_X1 U14866 ( .A1(\SB1_1_8/i0_3 ), .A2(\SB1_1_8/i0_0 ), .A3(
        \SB1_1_8/i0_4 ), .ZN(\SB1_1_8/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U14867 ( .A1(\MC_ARK_ARC_1_3/temp5[145] ), .A2(
        \MC_ARK_ARC_1_3/temp6[145] ), .Z(\MC_ARK_ARC_1_3/buf_output[145] ) );
  NAND4_X2 U14868 ( .A1(\SB2_4_5/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_4_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_4_5/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_4_5/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_4_5/buf_output[1] ) );
  NAND4_X2 U14869 ( .A1(\SB1_4_21/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_4_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_4_21/Component_Function_1/NAND4_in[0] ), .A4(n7540), .ZN(
        \SB1_4_21/buf_output[1] ) );
  XOR2_X1 U14870 ( .A1(\MC_ARK_ARC_1_3/temp5[181] ), .A2(n7542), .Z(
        \MC_ARK_ARC_1_3/buf_output[181] ) );
  XOR2_X1 U14871 ( .A1(\MC_ARK_ARC_1_3/temp3[181] ), .A2(
        \MC_ARK_ARC_1_3/temp4[181] ), .Z(n7542) );
  XOR2_X1 U14872 ( .A1(n7543), .A2(n2806), .Z(\MC_ARK_ARC_1_3/buf_output[109] ) );
  XOR2_X1 U14873 ( .A1(\MC_ARK_ARC_1_3/temp2[109] ), .A2(
        \MC_ARK_ARC_1_3/temp1[109] ), .Z(n7543) );
  XOR2_X1 U14874 ( .A1(n4581), .A2(\MC_ARK_ARC_1_4/temp1[102] ), .Z(
        \MC_ARK_ARC_1_4/temp5[102] ) );
  NAND4_X2 U14875 ( .A1(\SB3_31/Component_Function_4/NAND4_in[3] ), .A2(
        \SB3_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_4/NAND4_in[0] ), .A4(n7544), .ZN(
        \SB3_31/buf_output[4] ) );
  NAND3_X2 U14876 ( .A1(\SB3_31/i0[9] ), .A2(\SB3_31/i0_3 ), .A3(
        \SB3_31/i0[10] ), .ZN(n7544) );
  NAND3_X2 U14877 ( .A1(\SB1_3_4/i1_5 ), .A2(\SB1_3_4/i0_0 ), .A3(
        \SB1_3_4/i0_4 ), .ZN(n7545) );
  NAND3_X1 U14878 ( .A1(\SB1_4_10/i0[10] ), .A2(\SB1_4_10/i1_5 ), .A3(
        \SB1_4_10/i1[9] ), .ZN(\SB1_4_10/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U14879 ( .A1(\RI5[3][17] ), .A2(\RI5[3][185] ), .Z(n804) );
  NAND3_X2 U14880 ( .A1(\SB1_3_29/i0[9] ), .A2(\SB1_3_29/i0[6] ), .A3(
        \SB1_3_29/i0_4 ), .ZN(n7546) );
  XOR2_X1 U14881 ( .A1(n7547), .A2(n1910), .Z(\MC_ARK_ARC_1_1/buf_output[51] )
         );
  XOR2_X1 U14882 ( .A1(\MC_ARK_ARC_1_1/temp4[51] ), .A2(n5224), .Z(n7547) );
  NAND3_X1 U14883 ( .A1(\SB1_2_28/i0[10] ), .A2(\SB1_2_28/i1[9] ), .A3(
        \SB1_2_28/i1_7 ), .ZN(n7548) );
  INV_X2 U14884 ( .I(\SB1_0_6/buf_output[3] ), .ZN(\SB2_0_4/i0[8] ) );
  NAND4_X2 U14885 ( .A1(\SB1_0_6/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_0_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_6/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_0_6/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB1_0_6/buf_output[3] ) );
  NAND3_X1 U14886 ( .A1(\SB1_1_24/i0_4 ), .A2(\SB1_1_24/i0[10] ), .A3(
        \RI1[1][47] ), .ZN(\SB1_1_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U14887 ( .A1(\SB2_1_1/i0_4 ), .A2(\SB2_1_1/i0[9] ), .A3(
        \SB2_1_1/i0[6] ), .ZN(n4543) );
  NAND3_X1 U14888 ( .A1(\SB4_31/i1_5 ), .A2(\SB4_31/i3[0] ), .A3(
        \SB4_31/i0[8] ), .ZN(n7550) );
  XOR2_X1 U14889 ( .A1(\RI5[4][95] ), .A2(\RI5[4][47] ), .Z(n7551) );
  XOR2_X1 U14890 ( .A1(\RI5[0][47] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[41] ), 
        .Z(n7552) );
  XOR2_X1 U14891 ( .A1(n7553), .A2(\MC_ARK_ARC_1_1/temp5[24] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[24] ) );
  XOR2_X1 U14892 ( .A1(\MC_ARK_ARC_1_1/temp3[24] ), .A2(
        \MC_ARK_ARC_1_1/temp4[24] ), .Z(n7553) );
  NAND3_X2 U14893 ( .A1(\SB2_1_30/i0_4 ), .A2(\SB2_1_30/i0_0 ), .A3(
        \SB2_1_30/i1_5 ), .ZN(n7554) );
  NAND4_X2 U14894 ( .A1(\SB1_1_31/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_1_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_31/Component_Function_4/NAND4_in[0] ), .A4(n7555), .ZN(
        \SB1_1_31/buf_output[4] ) );
  XOR2_X1 U14895 ( .A1(\MC_ARK_ARC_1_0/temp5[168] ), .A2(n7556), .Z(
        \MC_ARK_ARC_1_0/buf_output[168] ) );
  XOR2_X1 U14896 ( .A1(\MC_ARK_ARC_1_0/temp3[168] ), .A2(
        \MC_ARK_ARC_1_0/temp4[168] ), .Z(n7556) );
  NAND3_X1 U14897 ( .A1(\SB3_16/i0[8] ), .A2(\SB3_16/i3[0] ), .A3(
        \SB3_16/i1_5 ), .ZN(n4773) );
  INV_X1 U14898 ( .I(\SB1_1_26/buf_output[1] ), .ZN(\SB2_1_22/i1_7 ) );
  NAND4_X2 U14899 ( .A1(\SB1_1_26/Component_Function_1/NAND4_in[1] ), .A2(
        n3642), .A3(\SB1_1_26/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_1_26/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_1_26/buf_output[1] ) );
  NAND4_X2 U14900 ( .A1(n4796), .A2(
        \SB1_4_24/Component_Function_4/NAND4_in[2] ), .A3(n5149), .A4(n7559), 
        .ZN(\SB1_4_24/buf_output[4] ) );
  NAND3_X1 U14901 ( .A1(\SB4_14/i0_0 ), .A2(n1495), .A3(\SB4_14/i0_4 ), .ZN(
        n7560) );
  NAND4_X2 U14902 ( .A1(\SB1_0_20/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_20/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_20/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_0_20/Component_Function_2/NAND4_in[0] ), .ZN(\RI3[0][86] ) );
  XOR2_X1 U14903 ( .A1(n4479), .A2(n4480), .Z(\MC_ARK_ARC_1_0/buf_output[38] )
         );
  XOR2_X1 U14904 ( .A1(n7561), .A2(n7562), .Z(\MC_ARK_ARC_1_1/buf_output[120] ) );
  XOR2_X1 U14905 ( .A1(n971), .A2(n806), .Z(n7561) );
  XOR2_X1 U14906 ( .A1(n4513), .A2(\MC_ARK_ARC_1_1/temp4[120] ), .Z(n7562) );
  XOR2_X1 U14907 ( .A1(n7563), .A2(n1197), .Z(\MC_ARK_ARC_1_1/buf_output[109] ) );
  NAND4_X2 U14908 ( .A1(\SB1_1_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_14/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_1_14/Component_Function_4/NAND4_in[1] ), .A4(n7564), .ZN(
        \SB1_1_14/buf_output[4] ) );
  XOR2_X1 U14909 ( .A1(\MC_ARK_ARC_1_1/temp5[118] ), .A2(
        \MC_ARK_ARC_1_1/temp6[118] ), .Z(\MC_ARK_ARC_1_1/buf_output[118] ) );
  NAND4_X2 U14910 ( .A1(\SB1_1_15/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_15/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_1_15/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_1_15/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_1_15/buf_output[1] ) );
  XOR2_X1 U14911 ( .A1(\RI5[4][149] ), .A2(\RI5[4][185] ), .Z(
        \MC_ARK_ARC_1_4/temp3[83] ) );
  INV_X2 U14912 ( .I(\SB1_4_12/buf_output[2] ), .ZN(\SB2_4_9/i1[9] ) );
  NAND3_X2 U14913 ( .A1(n600), .A2(\SB2_2_23/i1[9] ), .A3(\SB2_2_23/i1_5 ), 
        .ZN(n7573) );
  NAND3_X1 U14914 ( .A1(\SB2_4_20/i0[7] ), .A2(\SB2_4_20/i0_0 ), .A3(
        \SB2_4_20/i0_3 ), .ZN(\SB2_4_20/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U14915 ( .A1(\RI5[2][188] ), .A2(\RI5[2][32] ), .Z(
        \MC_ARK_ARC_1_2/temp3[122] ) );
  XOR2_X1 U14916 ( .A1(\MC_ARK_ARC_1_2/temp5[17] ), .A2(n2372), .Z(n3125) );
  NAND3_X1 U14917 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0[10] ), .A3(
        \SB2_2_30/i0[9] ), .ZN(n7567) );
  XOR2_X1 U14918 ( .A1(\MC_ARK_ARC_1_3/temp5[152] ), .A2(n7568), .Z(
        \MC_ARK_ARC_1_3/buf_output[152] ) );
  XOR2_X1 U14919 ( .A1(n2013), .A2(\MC_ARK_ARC_1_3/temp4[152] ), .Z(n7568) );
  XOR2_X1 U14920 ( .A1(n7569), .A2(n211), .Z(Ciphertext[130]) );
  XOR2_X1 U14921 ( .A1(\MC_ARK_ARC_1_0/temp1[86] ), .A2(
        \MC_ARK_ARC_1_0/temp4[86] ), .Z(n7571) );
  NAND4_X2 U14922 ( .A1(\SB2_2_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_23/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_2_23/Component_Function_4/NAND4_in[1] ), .A4(n7573), .ZN(
        \SB2_2_23/buf_output[4] ) );
  XOR2_X1 U14923 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[32] ), .A2(\RI5[1][68] ), 
        .Z(n5219) );
  NAND3_X2 U14924 ( .A1(\SB2_1_3/i0_4 ), .A2(\SB2_1_3/i0_3 ), .A3(
        \SB2_1_3/i0_0 ), .ZN(n7574) );
  NAND3_X2 U14925 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0[10] ), .A3(
        \RI3[0][58] ), .ZN(\SB2_0_22/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U14926 ( .A1(\SB2_1_3/Component_Function_3/NAND4_in[2] ), .A2(n2999), .A3(n3472), .A4(n7574), .ZN(\SB2_1_3/buf_output[3] ) );
  NAND3_X2 U14927 ( .A1(\SB1_1_3/i0_4 ), .A2(\SB1_1_3/i0[6] ), .A3(
        \SB1_1_3/i0[9] ), .ZN(n7575) );
  NAND4_X2 U14928 ( .A1(\SB2_3_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_7/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_3_7/Component_Function_3/NAND4_in[3] ), .A4(n7576), .ZN(
        \SB2_3_7/buf_output[3] ) );
  NAND3_X2 U14929 ( .A1(\SB3_7/i0_3 ), .A2(\SB3_7/i1[9] ), .A3(\SB3_7/i0[6] ), 
        .ZN(n7577) );
  NAND3_X2 U14930 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i0_4 ), .A3(\SB3_0/i1[9] ), 
        .ZN(n3309) );
  NAND3_X1 U14931 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i0_3 ), .A3(\SB4_5/i0[6] ), 
        .ZN(n3541) );
  XOR2_X1 U14932 ( .A1(\MC_ARK_ARC_1_2/temp3[115] ), .A2(
        \MC_ARK_ARC_1_2/temp2[115] ), .Z(n7579) );
  XOR2_X1 U14933 ( .A1(\RI5[4][71] ), .A2(\RI5[4][35] ), .Z(
        \MC_ARK_ARC_1_4/temp3[161] ) );
  NAND3_X1 U14934 ( .A1(\SB4_27/i0[9] ), .A2(\SB4_27/i0_3 ), .A3(
        \SB4_27/i0[10] ), .ZN(n7580) );
  NAND4_X2 U14935 ( .A1(\SB2_4_13/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_4_13/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_4_13/Component_Function_3/NAND4_in[3] ), .A4(n7581), .ZN(
        \SB2_4_13/buf_output[3] ) );
  NAND4_X2 U14936 ( .A1(\SB2_2_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_31/Component_Function_2/NAND4_in[1] ), .A3(n4443), .A4(n7582), 
        .ZN(\SB2_2_31/buf_output[2] ) );
  NAND3_X2 U14937 ( .A1(\SB2_2_31/i0[9] ), .A2(\SB2_2_31/i0_3 ), .A3(
        \SB2_2_31/i0[8] ), .ZN(n7582) );
  NAND3_X1 U14938 ( .A1(\SB1_1_15/i0[8] ), .A2(\SB1_1_15/i0_4 ), .A3(
        \SB1_1_15/i1_7 ), .ZN(\SB1_1_15/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U14939 ( .A1(\SB2_4_4/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_4_4/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_4_4/Component_Function_4/NAND4_in[3] ), .A4(n7583), .ZN(
        \SB2_4_4/buf_output[4] ) );
  NAND3_X2 U14940 ( .A1(\SB2_4_4/i0_3 ), .A2(\SB2_4_4/i0[10] ), .A3(
        \SB2_4_4/i0[9] ), .ZN(n7583) );
  XOR2_X1 U14941 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[120] ), .A2(\RI5[2][144] ), .Z(n7584) );
  NAND4_X2 U14942 ( .A1(\SB1_2_25/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_2_25/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_25/Component_Function_4/NAND4_in[1] ), .A4(n7588), .ZN(
        \SB1_2_25/buf_output[4] ) );
  XOR2_X1 U14943 ( .A1(\MC_ARK_ARC_1_4/temp1[165] ), .A2(
        \MC_ARK_ARC_1_4/temp2[165] ), .Z(n7589) );
  XOR2_X1 U14944 ( .A1(n7590), .A2(n210), .Z(Ciphertext[63]) );
  NAND4_X2 U14945 ( .A1(n2406), .A2(\SB3_15/Component_Function_3/NAND4_in[1] ), 
        .A3(\SB3_15/Component_Function_3/NAND4_in[0] ), .A4(
        \SB3_15/Component_Function_3/NAND4_in[3] ), .ZN(\SB3_15/buf_output[3] ) );
endmodule


module SPEEDY_Top ( clk, Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  input clk;

  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFFSNQ_X1 \reg_in_reg[191]  ( .D(Plaintext[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[191]) );
  DFFSNQ_X1 \reg_in_reg[190]  ( .D(Plaintext[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[190]) );
  DFFSNQ_X1 \reg_in_reg[189]  ( .D(Plaintext[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[189]) );
  DFFSNQ_X1 \reg_in_reg[188]  ( .D(Plaintext[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[188]) );
  DFFSNQ_X1 \reg_in_reg[187]  ( .D(Plaintext[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[187]) );
  DFFSNQ_X1 \reg_in_reg[186]  ( .D(Plaintext[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[186]) );
  DFFSNQ_X1 \reg_in_reg[185]  ( .D(Plaintext[185]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[185]) );
  DFFSNQ_X1 \reg_in_reg[184]  ( .D(Plaintext[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[184]) );
  DFFSNQ_X1 \reg_in_reg[183]  ( .D(Plaintext[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[183]) );
  DFFSNQ_X1 \reg_in_reg[182]  ( .D(Plaintext[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[182]) );
  DFFSNQ_X1 \reg_in_reg[181]  ( .D(Plaintext[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[181]) );
  DFFSNQ_X1 \reg_in_reg[180]  ( .D(Plaintext[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[180]) );
  DFFSNQ_X1 \reg_in_reg[179]  ( .D(Plaintext[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[179]) );
  DFFSNQ_X1 \reg_in_reg[178]  ( .D(Plaintext[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[178]) );
  DFFSNQ_X1 \reg_in_reg[177]  ( .D(Plaintext[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[177]) );
  DFFSNQ_X1 \reg_in_reg[176]  ( .D(Plaintext[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[176]) );
  DFFSNQ_X1 \reg_in_reg[175]  ( .D(Plaintext[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[175]) );
  DFFSNQ_X1 \reg_in_reg[174]  ( .D(Plaintext[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[174]) );
  DFFSNQ_X1 \reg_in_reg[173]  ( .D(Plaintext[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[173]) );
  DFFSNQ_X1 \reg_in_reg[172]  ( .D(Plaintext[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[172]) );
  DFFSNQ_X1 \reg_in_reg[171]  ( .D(Plaintext[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[171]) );
  DFFSNQ_X1 \reg_in_reg[170]  ( .D(Plaintext[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[170]) );
  DFFSNQ_X1 \reg_in_reg[169]  ( .D(Plaintext[169]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[169]) );
  DFFSNQ_X1 \reg_in_reg[168]  ( .D(Plaintext[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[168]) );
  DFFSNQ_X1 \reg_in_reg[167]  ( .D(Plaintext[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[167]) );
  DFFSNQ_X1 \reg_in_reg[166]  ( .D(Plaintext[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[166]) );
  DFFSNQ_X1 \reg_in_reg[165]  ( .D(Plaintext[165]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[165]) );
  DFFSNQ_X1 \reg_in_reg[164]  ( .D(Plaintext[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[164]) );
  DFFSNQ_X1 \reg_in_reg[163]  ( .D(Plaintext[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[163]) );
  DFFSNQ_X1 \reg_in_reg[162]  ( .D(Plaintext[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[162]) );
  DFFSNQ_X1 \reg_in_reg[161]  ( .D(Plaintext[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[161]) );
  DFFSNQ_X1 \reg_in_reg[160]  ( .D(Plaintext[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[160]) );
  DFFSNQ_X1 \reg_in_reg[159]  ( .D(Plaintext[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[159]) );
  DFFSNQ_X1 \reg_in_reg[158]  ( .D(Plaintext[158]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[158]) );
  DFFSNQ_X1 \reg_in_reg[157]  ( .D(Plaintext[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[157]) );
  DFFSNQ_X1 \reg_in_reg[156]  ( .D(Plaintext[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[156]) );
  DFFSNQ_X1 \reg_in_reg[155]  ( .D(Plaintext[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[155]) );
  DFFSNQ_X1 \reg_in_reg[154]  ( .D(Plaintext[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[154]) );
  DFFSNQ_X1 \reg_in_reg[153]  ( .D(Plaintext[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[153]) );
  DFFSNQ_X1 \reg_in_reg[152]  ( .D(Plaintext[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[152]) );
  DFFSNQ_X1 \reg_in_reg[151]  ( .D(Plaintext[151]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[151]) );
  DFFSNQ_X1 \reg_in_reg[150]  ( .D(Plaintext[150]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[150]) );
  DFFSNQ_X1 \reg_in_reg[149]  ( .D(Plaintext[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[149]) );
  DFFSNQ_X1 \reg_in_reg[148]  ( .D(Plaintext[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[148]) );
  DFFSNQ_X1 \reg_in_reg[147]  ( .D(Plaintext[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[147]) );
  DFFSNQ_X1 \reg_in_reg[146]  ( .D(Plaintext[146]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[146]) );
  DFFSNQ_X1 \reg_in_reg[145]  ( .D(Plaintext[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[145]) );
  DFFSNQ_X1 \reg_in_reg[144]  ( .D(Plaintext[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[144]) );
  DFFSNQ_X1 \reg_in_reg[143]  ( .D(Plaintext[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[143]) );
  DFFSNQ_X1 \reg_in_reg[142]  ( .D(Plaintext[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[142]) );
  DFFSNQ_X1 \reg_in_reg[141]  ( .D(Plaintext[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[141]) );
  DFFSNQ_X1 \reg_in_reg[140]  ( .D(Plaintext[140]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[140]) );
  DFFSNQ_X1 \reg_in_reg[139]  ( .D(Plaintext[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[139]) );
  DFFSNQ_X1 \reg_in_reg[138]  ( .D(Plaintext[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[138]) );
  DFFSNQ_X1 \reg_in_reg[137]  ( .D(Plaintext[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[137]) );
  DFFSNQ_X1 \reg_in_reg[136]  ( .D(Plaintext[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[136]) );
  DFFSNQ_X1 \reg_in_reg[135]  ( .D(Plaintext[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[135]) );
  DFFSNQ_X1 \reg_in_reg[134]  ( .D(Plaintext[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[134]) );
  DFFSNQ_X1 \reg_in_reg[133]  ( .D(Plaintext[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[133]) );
  DFFSNQ_X1 \reg_in_reg[132]  ( .D(Plaintext[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[132]) );
  DFFSNQ_X1 \reg_in_reg[131]  ( .D(Plaintext[131]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[131]) );
  DFFSNQ_X1 \reg_in_reg[130]  ( .D(Plaintext[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[130]) );
  DFFSNQ_X1 \reg_in_reg[129]  ( .D(Plaintext[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[129]) );
  DFFSNQ_X1 \reg_in_reg[128]  ( .D(Plaintext[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[128]) );
  DFFSNQ_X1 \reg_in_reg[127]  ( .D(Plaintext[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[127]) );
  DFFSNQ_X1 \reg_in_reg[126]  ( .D(Plaintext[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[126]) );
  DFFSNQ_X1 \reg_in_reg[125]  ( .D(Plaintext[125]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[125]) );
  DFFSNQ_X1 \reg_in_reg[124]  ( .D(Plaintext[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[124]) );
  DFFSNQ_X1 \reg_in_reg[123]  ( .D(Plaintext[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[123]) );
  DFFSNQ_X1 \reg_in_reg[122]  ( .D(Plaintext[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[122]) );
  DFFSNQ_X1 \reg_in_reg[121]  ( .D(Plaintext[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[121]) );
  DFFSNQ_X1 \reg_in_reg[120]  ( .D(Plaintext[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[120]) );
  DFFSNQ_X1 \reg_in_reg[119]  ( .D(Plaintext[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[119]) );
  DFFSNQ_X1 \reg_in_reg[118]  ( .D(Plaintext[118]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[118]) );
  DFFSNQ_X1 \reg_in_reg[117]  ( .D(Plaintext[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[117]) );
  DFFSNQ_X1 \reg_in_reg[116]  ( .D(Plaintext[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[116]) );
  DFFSNQ_X1 \reg_in_reg[115]  ( .D(Plaintext[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[115]) );
  DFFSNQ_X1 \reg_in_reg[114]  ( .D(Plaintext[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[114]) );
  DFFSNQ_X1 \reg_in_reg[113]  ( .D(Plaintext[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[113]) );
  DFFSNQ_X1 \reg_in_reg[112]  ( .D(Plaintext[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[112]) );
  DFFSNQ_X1 \reg_in_reg[111]  ( .D(Plaintext[111]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[111]) );
  DFFSNQ_X1 \reg_in_reg[110]  ( .D(Plaintext[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[110]) );
  DFFSNQ_X1 \reg_in_reg[109]  ( .D(Plaintext[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[109]) );
  DFFSNQ_X1 \reg_in_reg[108]  ( .D(Plaintext[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[108]) );
  DFFSNQ_X1 \reg_in_reg[107]  ( .D(Plaintext[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[107]) );
  DFFSNQ_X1 \reg_in_reg[106]  ( .D(Plaintext[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[106]) );
  DFFSNQ_X1 \reg_in_reg[105]  ( .D(Plaintext[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[105]) );
  DFFSNQ_X1 \reg_in_reg[104]  ( .D(Plaintext[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[104]) );
  DFFSNQ_X1 \reg_in_reg[103]  ( .D(Plaintext[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[103]) );
  DFFSNQ_X1 \reg_in_reg[102]  ( .D(Plaintext[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[102]) );
  DFFSNQ_X1 \reg_in_reg[101]  ( .D(Plaintext[101]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[101]) );
  DFFSNQ_X1 \reg_in_reg[100]  ( .D(Plaintext[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[100]) );
  DFFSNQ_X1 \reg_in_reg[99]  ( .D(Plaintext[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[99]) );
  DFFSNQ_X1 \reg_in_reg[98]  ( .D(Plaintext[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[98]) );
  DFFSNQ_X1 \reg_in_reg[97]  ( .D(Plaintext[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[97]) );
  DFFSNQ_X1 \reg_in_reg[96]  ( .D(Plaintext[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[96]) );
  DFFSNQ_X1 \reg_in_reg[95]  ( .D(Plaintext[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[95]) );
  DFFSNQ_X1 \reg_in_reg[94]  ( .D(Plaintext[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[94]) );
  DFFSNQ_X1 \reg_in_reg[93]  ( .D(Plaintext[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[93]) );
  DFFSNQ_X1 \reg_in_reg[92]  ( .D(Plaintext[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[92]) );
  DFFSNQ_X1 \reg_in_reg[91]  ( .D(Plaintext[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[91]) );
  DFFSNQ_X1 \reg_in_reg[90]  ( .D(Plaintext[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[90]) );
  DFFSNQ_X1 \reg_in_reg[89]  ( .D(Plaintext[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[89]) );
  DFFSNQ_X1 \reg_in_reg[88]  ( .D(Plaintext[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[88]) );
  DFFSNQ_X1 \reg_in_reg[87]  ( .D(Plaintext[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[87]) );
  DFFSNQ_X1 \reg_in_reg[86]  ( .D(Plaintext[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[86]) );
  DFFSNQ_X1 \reg_in_reg[85]  ( .D(Plaintext[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[85]) );
  DFFSNQ_X1 \reg_in_reg[84]  ( .D(Plaintext[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[84]) );
  DFFSNQ_X1 \reg_in_reg[83]  ( .D(Plaintext[83]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[83]) );
  DFFSNQ_X1 \reg_in_reg[82]  ( .D(Plaintext[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[82]) );
  DFFSNQ_X1 \reg_in_reg[81]  ( .D(Plaintext[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[81]) );
  DFFSNQ_X1 \reg_in_reg[80]  ( .D(Plaintext[80]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[80]) );
  DFFSNQ_X1 \reg_in_reg[79]  ( .D(Plaintext[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[79]) );
  DFFSNQ_X1 \reg_in_reg[78]  ( .D(Plaintext[78]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[78]) );
  DFFSNQ_X1 \reg_in_reg[77]  ( .D(Plaintext[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[77]) );
  DFFSNQ_X1 \reg_in_reg[76]  ( .D(Plaintext[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[76]) );
  DFFSNQ_X1 \reg_in_reg[75]  ( .D(Plaintext[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[75]) );
  DFFSNQ_X1 \reg_in_reg[74]  ( .D(Plaintext[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[74]) );
  DFFSNQ_X1 \reg_in_reg[73]  ( .D(Plaintext[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[73]) );
  DFFSNQ_X1 \reg_in_reg[72]  ( .D(Plaintext[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[72]) );
  DFFSNQ_X1 \reg_in_reg[71]  ( .D(Plaintext[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[71]) );
  DFFSNQ_X1 \reg_in_reg[70]  ( .D(Plaintext[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[70]) );
  DFFSNQ_X1 \reg_in_reg[69]  ( .D(Plaintext[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[69]) );
  DFFSNQ_X1 \reg_in_reg[68]  ( .D(Plaintext[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[68]) );
  DFFSNQ_X1 \reg_in_reg[67]  ( .D(Plaintext[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[67]) );
  DFFSNQ_X1 \reg_in_reg[66]  ( .D(Plaintext[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[66]) );
  DFFSNQ_X1 \reg_in_reg[65]  ( .D(Plaintext[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[65]) );
  DFFSNQ_X1 \reg_in_reg[64]  ( .D(Plaintext[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[64]) );
  DFFSNQ_X1 \reg_in_reg[63]  ( .D(Plaintext[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[63]) );
  DFFSNQ_X1 \reg_in_reg[62]  ( .D(Plaintext[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[62]) );
  DFFSNQ_X1 \reg_in_reg[61]  ( .D(Plaintext[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[61]) );
  DFFSNQ_X1 \reg_in_reg[60]  ( .D(Plaintext[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[60]) );
  DFFSNQ_X1 \reg_in_reg[59]  ( .D(Plaintext[59]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[59]) );
  DFFSNQ_X1 \reg_in_reg[58]  ( .D(Plaintext[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[58]) );
  DFFSNQ_X1 \reg_in_reg[57]  ( .D(Plaintext[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[57]) );
  DFFSNQ_X1 \reg_in_reg[56]  ( .D(Plaintext[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[56]) );
  DFFSNQ_X1 \reg_in_reg[55]  ( .D(Plaintext[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[55]) );
  DFFSNQ_X1 \reg_in_reg[54]  ( .D(Plaintext[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[54]) );
  DFFSNQ_X1 \reg_in_reg[53]  ( .D(Plaintext[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[53]) );
  DFFSNQ_X1 \reg_in_reg[52]  ( .D(Plaintext[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[52]) );
  DFFSNQ_X1 \reg_in_reg[51]  ( .D(Plaintext[51]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[51]) );
  DFFSNQ_X1 \reg_in_reg[50]  ( .D(Plaintext[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[50]) );
  DFFSNQ_X1 \reg_in_reg[49]  ( .D(Plaintext[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[49]) );
  DFFSNQ_X1 \reg_in_reg[48]  ( .D(Plaintext[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[48]) );
  DFFSNQ_X1 \reg_in_reg[47]  ( .D(Plaintext[47]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[47]) );
  DFFSNQ_X1 \reg_in_reg[46]  ( .D(Plaintext[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[46]) );
  DFFSNQ_X1 \reg_in_reg[45]  ( .D(Plaintext[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[45]) );
  DFFSNQ_X1 \reg_in_reg[44]  ( .D(Plaintext[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[44]) );
  DFFSNQ_X1 \reg_in_reg[43]  ( .D(Plaintext[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[43]) );
  DFFSNQ_X1 \reg_in_reg[42]  ( .D(Plaintext[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[42]) );
  DFFSNQ_X1 \reg_in_reg[41]  ( .D(Plaintext[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[41]) );
  DFFSNQ_X1 \reg_in_reg[40]  ( .D(Plaintext[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[40]) );
  DFFSNQ_X1 \reg_in_reg[39]  ( .D(Plaintext[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[39]) );
  DFFSNQ_X1 \reg_in_reg[38]  ( .D(Plaintext[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[38]) );
  DFFSNQ_X1 \reg_in_reg[37]  ( .D(Plaintext[37]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[37]) );
  DFFSNQ_X1 \reg_in_reg[36]  ( .D(Plaintext[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[36]) );
  DFFSNQ_X1 \reg_in_reg[35]  ( .D(Plaintext[35]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[35]) );
  DFFSNQ_X1 \reg_in_reg[34]  ( .D(Plaintext[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[34]) );
  DFFSNQ_X1 \reg_in_reg[33]  ( .D(Plaintext[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[33]) );
  DFFSNQ_X1 \reg_in_reg[32]  ( .D(Plaintext[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[32]) );
  DFFSNQ_X1 \reg_in_reg[31]  ( .D(Plaintext[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[31]) );
  DFFSNQ_X1 \reg_in_reg[30]  ( .D(Plaintext[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[30]) );
  DFFSNQ_X1 \reg_in_reg[29]  ( .D(Plaintext[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[29]) );
  DFFSNQ_X1 \reg_in_reg[28]  ( .D(Plaintext[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[28]) );
  DFFSNQ_X1 \reg_in_reg[27]  ( .D(Plaintext[27]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[27]) );
  DFFSNQ_X1 \reg_in_reg[26]  ( .D(Plaintext[26]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[26]) );
  DFFSNQ_X1 \reg_in_reg[25]  ( .D(Plaintext[25]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[25]) );
  DFFSNQ_X1 \reg_in_reg[24]  ( .D(Plaintext[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[24]) );
  DFFSNQ_X1 \reg_in_reg[23]  ( .D(Plaintext[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[23]) );
  DFFSNQ_X1 \reg_in_reg[22]  ( .D(Plaintext[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[22]) );
  DFFSNQ_X1 \reg_in_reg[21]  ( .D(Plaintext[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[21]) );
  DFFSNQ_X1 \reg_in_reg[20]  ( .D(Plaintext[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[20]) );
  DFFSNQ_X1 \reg_in_reg[19]  ( .D(Plaintext[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[19]) );
  DFFSNQ_X1 \reg_in_reg[18]  ( .D(Plaintext[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[18]) );
  DFFSNQ_X1 \reg_in_reg[17]  ( .D(Plaintext[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[17]) );
  DFFSNQ_X1 \reg_in_reg[16]  ( .D(Plaintext[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[16]) );
  DFFSNQ_X1 \reg_in_reg[15]  ( .D(Plaintext[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[15]) );
  DFFSNQ_X1 \reg_in_reg[14]  ( .D(Plaintext[14]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[14]) );
  DFFSNQ_X1 \reg_in_reg[13]  ( .D(Plaintext[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[13]) );
  DFFSNQ_X1 \reg_in_reg[12]  ( .D(Plaintext[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[12]) );
  DFFSNQ_X1 \reg_in_reg[11]  ( .D(Plaintext[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[11]) );
  DFFSNQ_X1 \reg_in_reg[10]  ( .D(Plaintext[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[10]) );
  DFFSNQ_X1 \reg_in_reg[9]  ( .D(Plaintext[9]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[9]) );
  DFFSNQ_X1 \reg_in_reg[8]  ( .D(Plaintext[8]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[8]) );
  DFFSNQ_X1 \reg_in_reg[7]  ( .D(Plaintext[7]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[7]) );
  DFFSNQ_X1 \reg_in_reg[6]  ( .D(Plaintext[6]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[6]) );
  DFFSNQ_X1 \reg_in_reg[5]  ( .D(Plaintext[5]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[5]) );
  DFFSNQ_X1 \reg_in_reg[4]  ( .D(Plaintext[4]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[4]) );
  DFFSNQ_X1 \reg_in_reg[3]  ( .D(Plaintext[3]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[3]) );
  DFFSNQ_X1 \reg_in_reg[2]  ( .D(Plaintext[2]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[2]) );
  DFFSNQ_X1 \reg_in_reg[1]  ( .D(Plaintext[1]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[1]) );
  DFFSNQ_X1 \reg_in_reg[0]  ( .D(Plaintext[0]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[0]) );
  DFFSNQ_X1 \reg_key_reg[191]  ( .D(Key[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[191]) );
  DFFSNQ_X1 \reg_key_reg[190]  ( .D(Key[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[190]) );
  DFFSNQ_X1 \reg_key_reg[189]  ( .D(Key[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[189]) );
  DFFSNQ_X1 \reg_key_reg[188]  ( .D(Key[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[188]) );
  DFFSNQ_X1 \reg_key_reg[187]  ( .D(Key[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[187]) );
  DFFSNQ_X1 \reg_key_reg[186]  ( .D(Key[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[186]) );
  DFFSNQ_X1 \reg_key_reg[185]  ( .D(Key[185]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[185]) );
  DFFSNQ_X1 \reg_key_reg[184]  ( .D(Key[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[184]) );
  DFFSNQ_X1 \reg_key_reg[183]  ( .D(Key[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[183]) );
  DFFSNQ_X1 \reg_key_reg[182]  ( .D(Key[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[182]) );
  DFFSNQ_X1 \reg_key_reg[181]  ( .D(Key[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[181]) );
  DFFSNQ_X1 \reg_key_reg[180]  ( .D(Key[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[180]) );
  DFFSNQ_X1 \reg_key_reg[179]  ( .D(Key[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[179]) );
  DFFSNQ_X1 \reg_key_reg[178]  ( .D(Key[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[178]) );
  DFFSNQ_X1 \reg_key_reg[177]  ( .D(Key[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[177]) );
  DFFSNQ_X1 \reg_key_reg[176]  ( .D(Key[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[176]) );
  DFFSNQ_X1 \reg_key_reg[175]  ( .D(Key[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[175]) );
  DFFSNQ_X1 \reg_key_reg[174]  ( .D(Key[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[174]) );
  DFFSNQ_X1 \reg_key_reg[173]  ( .D(Key[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[173]) );
  DFFSNQ_X1 \reg_key_reg[172]  ( .D(Key[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[172]) );
  DFFSNQ_X1 \reg_key_reg[171]  ( .D(Key[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[171]) );
  DFFSNQ_X1 \reg_key_reg[170]  ( .D(Key[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[170]) );
  DFFSNQ_X1 \reg_key_reg[169]  ( .D(Key[169]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[169]) );
  DFFSNQ_X1 \reg_key_reg[168]  ( .D(Key[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[168]) );
  DFFSNQ_X1 \reg_key_reg[167]  ( .D(Key[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[167]) );
  DFFSNQ_X1 \reg_key_reg[166]  ( .D(Key[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[166]) );
  DFFSNQ_X1 \reg_key_reg[165]  ( .D(Key[165]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[165]) );
  DFFSNQ_X1 \reg_key_reg[164]  ( .D(Key[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[164]) );
  DFFSNQ_X1 \reg_key_reg[163]  ( .D(Key[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[163]) );
  DFFSNQ_X1 \reg_key_reg[162]  ( .D(Key[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[162]) );
  DFFSNQ_X1 \reg_key_reg[161]  ( .D(Key[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[161]) );
  DFFSNQ_X1 \reg_key_reg[160]  ( .D(Key[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[160]) );
  DFFSNQ_X1 \reg_key_reg[159]  ( .D(Key[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[159]) );
  DFFSNQ_X1 \reg_key_reg[158]  ( .D(Key[158]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[158]) );
  DFFSNQ_X1 \reg_key_reg[157]  ( .D(Key[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[157]) );
  DFFSNQ_X1 \reg_key_reg[156]  ( .D(Key[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[156]) );
  DFFSNQ_X1 \reg_key_reg[155]  ( .D(Key[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[155]) );
  DFFSNQ_X1 \reg_key_reg[154]  ( .D(Key[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[154]) );
  DFFSNQ_X1 \reg_key_reg[153]  ( .D(Key[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[153]) );
  DFFSNQ_X1 \reg_key_reg[152]  ( .D(Key[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[152]) );
  DFFSNQ_X1 \reg_key_reg[151]  ( .D(Key[151]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[151]) );
  DFFSNQ_X1 \reg_key_reg[150]  ( .D(Key[150]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[150]) );
  DFFSNQ_X1 \reg_key_reg[149]  ( .D(Key[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[149]) );
  DFFSNQ_X1 \reg_key_reg[148]  ( .D(Key[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[148]) );
  DFFSNQ_X1 \reg_key_reg[147]  ( .D(Key[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[147]) );
  DFFSNQ_X1 \reg_key_reg[146]  ( .D(Key[146]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[146]) );
  DFFSNQ_X1 \reg_key_reg[145]  ( .D(Key[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[145]) );
  DFFSNQ_X1 \reg_key_reg[144]  ( .D(Key[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[144]) );
  DFFSNQ_X1 \reg_key_reg[143]  ( .D(Key[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[143]) );
  DFFSNQ_X1 \reg_key_reg[142]  ( .D(Key[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[142]) );
  DFFSNQ_X1 \reg_key_reg[141]  ( .D(Key[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[141]) );
  DFFSNQ_X1 \reg_key_reg[140]  ( .D(Key[140]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[140]) );
  DFFSNQ_X1 \reg_key_reg[139]  ( .D(Key[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[139]) );
  DFFSNQ_X1 \reg_key_reg[138]  ( .D(Key[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[138]) );
  DFFSNQ_X1 \reg_key_reg[137]  ( .D(Key[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[137]) );
  DFFSNQ_X1 \reg_key_reg[136]  ( .D(Key[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[136]) );
  DFFSNQ_X1 \reg_key_reg[135]  ( .D(Key[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[135]) );
  DFFSNQ_X1 \reg_key_reg[134]  ( .D(Key[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[134]) );
  DFFSNQ_X1 \reg_key_reg[133]  ( .D(Key[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[133]) );
  DFFSNQ_X1 \reg_key_reg[132]  ( .D(Key[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[132]) );
  DFFSNQ_X1 \reg_key_reg[131]  ( .D(Key[131]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[131]) );
  DFFSNQ_X1 \reg_key_reg[130]  ( .D(Key[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[130]) );
  DFFSNQ_X1 \reg_key_reg[129]  ( .D(Key[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[129]) );
  DFFSNQ_X1 \reg_key_reg[128]  ( .D(Key[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[128]) );
  DFFSNQ_X1 \reg_key_reg[127]  ( .D(Key[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[127]) );
  DFFSNQ_X1 \reg_key_reg[126]  ( .D(Key[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[126]) );
  DFFSNQ_X1 \reg_key_reg[125]  ( .D(Key[125]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[125]) );
  DFFSNQ_X1 \reg_key_reg[124]  ( .D(Key[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[124]) );
  DFFSNQ_X1 \reg_key_reg[123]  ( .D(Key[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[123]) );
  DFFSNQ_X1 \reg_key_reg[122]  ( .D(Key[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[122]) );
  DFFSNQ_X1 \reg_key_reg[121]  ( .D(Key[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[121]) );
  DFFSNQ_X1 \reg_key_reg[120]  ( .D(Key[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[120]) );
  DFFSNQ_X1 \reg_key_reg[119]  ( .D(Key[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[119]) );
  DFFSNQ_X1 \reg_key_reg[118]  ( .D(Key[118]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[118]) );
  DFFSNQ_X1 \reg_key_reg[117]  ( .D(Key[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[117]) );
  DFFSNQ_X1 \reg_key_reg[116]  ( .D(Key[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[116]) );
  DFFSNQ_X1 \reg_key_reg[115]  ( .D(Key[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[115]) );
  DFFSNQ_X1 \reg_key_reg[114]  ( .D(Key[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[114]) );
  DFFSNQ_X1 \reg_key_reg[113]  ( .D(Key[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[113]) );
  DFFSNQ_X1 \reg_key_reg[112]  ( .D(Key[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[112]) );
  DFFSNQ_X1 \reg_key_reg[111]  ( .D(Key[111]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[111]) );
  DFFSNQ_X1 \reg_key_reg[110]  ( .D(Key[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[110]) );
  DFFSNQ_X1 \reg_key_reg[109]  ( .D(Key[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[109]) );
  DFFSNQ_X1 \reg_key_reg[108]  ( .D(Key[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[108]) );
  DFFSNQ_X1 \reg_key_reg[107]  ( .D(Key[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[107]) );
  DFFSNQ_X1 \reg_key_reg[106]  ( .D(Key[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[106]) );
  DFFSNQ_X1 \reg_key_reg[105]  ( .D(Key[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[105]) );
  DFFSNQ_X1 \reg_key_reg[104]  ( .D(Key[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[104]) );
  DFFSNQ_X1 \reg_key_reg[103]  ( .D(Key[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[103]) );
  DFFSNQ_X1 \reg_key_reg[102]  ( .D(Key[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[102]) );
  DFFSNQ_X1 \reg_key_reg[101]  ( .D(Key[101]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[101]) );
  DFFSNQ_X1 \reg_key_reg[100]  ( .D(Key[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[100]) );
  DFFSNQ_X1 \reg_key_reg[99]  ( .D(Key[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[99]) );
  DFFSNQ_X1 \reg_key_reg[98]  ( .D(Key[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[98]) );
  DFFSNQ_X1 \reg_key_reg[97]  ( .D(Key[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[97]) );
  DFFSNQ_X1 \reg_key_reg[96]  ( .D(Key[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[96]) );
  DFFSNQ_X1 \reg_key_reg[95]  ( .D(Key[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[95]) );
  DFFSNQ_X1 \reg_key_reg[94]  ( .D(Key[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[94]) );
  DFFSNQ_X1 \reg_key_reg[93]  ( .D(Key[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[93]) );
  DFFSNQ_X1 \reg_key_reg[92]  ( .D(Key[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[92]) );
  DFFSNQ_X1 \reg_key_reg[91]  ( .D(Key[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[91]) );
  DFFSNQ_X1 \reg_key_reg[90]  ( .D(Key[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[90]) );
  DFFSNQ_X1 \reg_key_reg[89]  ( .D(Key[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[89]) );
  DFFSNQ_X1 \reg_key_reg[88]  ( .D(Key[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[88]) );
  DFFSNQ_X1 \reg_key_reg[87]  ( .D(Key[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[87]) );
  DFFSNQ_X1 \reg_key_reg[86]  ( .D(Key[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[86]) );
  DFFSNQ_X1 \reg_key_reg[85]  ( .D(Key[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[85]) );
  DFFSNQ_X1 \reg_key_reg[84]  ( .D(Key[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[84]) );
  DFFSNQ_X1 \reg_key_reg[83]  ( .D(Key[83]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[83]) );
  DFFSNQ_X1 \reg_key_reg[82]  ( .D(Key[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[82]) );
  DFFSNQ_X1 \reg_key_reg[81]  ( .D(Key[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[81]) );
  DFFSNQ_X1 \reg_key_reg[80]  ( .D(Key[80]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[80]) );
  DFFSNQ_X1 \reg_key_reg[79]  ( .D(Key[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[79]) );
  DFFSNQ_X1 \reg_key_reg[78]  ( .D(Key[78]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[78]) );
  DFFSNQ_X1 \reg_key_reg[77]  ( .D(Key[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[77]) );
  DFFSNQ_X1 \reg_key_reg[76]  ( .D(Key[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[76]) );
  DFFSNQ_X1 \reg_key_reg[75]  ( .D(Key[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[75]) );
  DFFSNQ_X1 \reg_key_reg[74]  ( .D(Key[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[74]) );
  DFFSNQ_X1 \reg_key_reg[73]  ( .D(Key[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[73]) );
  DFFSNQ_X1 \reg_key_reg[72]  ( .D(Key[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[72]) );
  DFFSNQ_X1 \reg_key_reg[71]  ( .D(Key[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[71]) );
  DFFSNQ_X1 \reg_key_reg[70]  ( .D(Key[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[70]) );
  DFFSNQ_X1 \reg_key_reg[69]  ( .D(Key[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[69]) );
  DFFSNQ_X1 \reg_key_reg[68]  ( .D(Key[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[68]) );
  DFFSNQ_X1 \reg_key_reg[67]  ( .D(Key[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[67]) );
  DFFSNQ_X1 \reg_key_reg[66]  ( .D(Key[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[66]) );
  DFFSNQ_X1 \reg_key_reg[65]  ( .D(Key[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[65]) );
  DFFSNQ_X1 \reg_key_reg[64]  ( .D(Key[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[64]) );
  DFFSNQ_X1 \reg_key_reg[63]  ( .D(Key[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[63]) );
  DFFSNQ_X1 \reg_key_reg[62]  ( .D(Key[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[62]) );
  DFFSNQ_X1 \reg_key_reg[61]  ( .D(Key[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[61]) );
  DFFSNQ_X1 \reg_key_reg[60]  ( .D(Key[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[60]) );
  DFFSNQ_X1 \reg_key_reg[59]  ( .D(Key[59]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[59]) );
  DFFSNQ_X1 \reg_key_reg[58]  ( .D(Key[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[58]) );
  DFFSNQ_X1 \reg_key_reg[57]  ( .D(Key[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[57]) );
  DFFSNQ_X1 \reg_key_reg[56]  ( .D(Key[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[56]) );
  DFFSNQ_X1 \reg_key_reg[55]  ( .D(Key[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[55]) );
  DFFSNQ_X1 \reg_key_reg[54]  ( .D(Key[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[54]) );
  DFFSNQ_X1 \reg_key_reg[53]  ( .D(Key[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[53]) );
  DFFSNQ_X1 \reg_key_reg[52]  ( .D(Key[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[52]) );
  DFFSNQ_X1 \reg_key_reg[51]  ( .D(Key[51]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[51]) );
  DFFSNQ_X1 \reg_key_reg[50]  ( .D(Key[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[50]) );
  DFFSNQ_X1 \reg_key_reg[49]  ( .D(Key[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[49]) );
  DFFSNQ_X1 \reg_key_reg[48]  ( .D(Key[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[48]) );
  DFFSNQ_X1 \reg_key_reg[47]  ( .D(Key[47]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[47]) );
  DFFSNQ_X1 \reg_key_reg[46]  ( .D(Key[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[46]) );
  DFFSNQ_X1 \reg_key_reg[45]  ( .D(Key[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[45]) );
  DFFSNQ_X1 \reg_key_reg[44]  ( .D(Key[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[44]) );
  DFFSNQ_X1 \reg_key_reg[43]  ( .D(Key[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[43]) );
  DFFSNQ_X1 \reg_key_reg[42]  ( .D(Key[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[42]) );
  DFFSNQ_X1 \reg_key_reg[41]  ( .D(Key[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[41]) );
  DFFSNQ_X1 \reg_key_reg[40]  ( .D(Key[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[40]) );
  DFFSNQ_X1 \reg_key_reg[39]  ( .D(Key[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[39]) );
  DFFSNQ_X1 \reg_key_reg[38]  ( .D(Key[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[38]) );
  DFFSNQ_X1 \reg_key_reg[37]  ( .D(Key[37]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[37]) );
  DFFSNQ_X1 \reg_key_reg[36]  ( .D(Key[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[36]) );
  DFFSNQ_X1 \reg_key_reg[35]  ( .D(Key[35]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[35]) );
  DFFSNQ_X1 \reg_key_reg[34]  ( .D(Key[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[34]) );
  DFFSNQ_X1 \reg_key_reg[33]  ( .D(Key[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[33]) );
  DFFSNQ_X1 \reg_key_reg[32]  ( .D(Key[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[32]) );
  DFFSNQ_X1 \reg_key_reg[31]  ( .D(Key[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[31]) );
  DFFSNQ_X1 \reg_key_reg[30]  ( .D(Key[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[30]) );
  DFFSNQ_X1 \reg_key_reg[29]  ( .D(Key[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[29]) );
  DFFSNQ_X1 \reg_key_reg[28]  ( .D(Key[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[28]) );
  DFFSNQ_X1 \reg_key_reg[27]  ( .D(Key[27]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[27]) );
  DFFSNQ_X1 \reg_key_reg[26]  ( .D(Key[26]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[26]) );
  DFFSNQ_X1 \reg_key_reg[25]  ( .D(Key[25]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[25]) );
  DFFSNQ_X1 \reg_key_reg[24]  ( .D(Key[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[24]) );
  DFFSNQ_X1 \reg_key_reg[23]  ( .D(Key[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[23]) );
  DFFSNQ_X1 \reg_key_reg[22]  ( .D(Key[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[22]) );
  DFFSNQ_X1 \reg_key_reg[21]  ( .D(Key[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[21]) );
  DFFSNQ_X1 \reg_key_reg[20]  ( .D(Key[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[20]) );
  DFFSNQ_X1 \reg_key_reg[19]  ( .D(Key[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[19]) );
  DFFSNQ_X1 \reg_key_reg[18]  ( .D(Key[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[18]) );
  DFFSNQ_X1 \reg_key_reg[17]  ( .D(Key[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[17]) );
  DFFSNQ_X1 \reg_key_reg[16]  ( .D(Key[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[16]) );
  DFFSNQ_X1 \reg_key_reg[15]  ( .D(Key[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[15]) );
  DFFSNQ_X1 \reg_key_reg[14]  ( .D(Key[14]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[14]) );
  DFFSNQ_X1 \reg_key_reg[13]  ( .D(Key[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[13]) );
  DFFSNQ_X1 \reg_key_reg[12]  ( .D(Key[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[12]) );
  DFFSNQ_X1 \reg_key_reg[11]  ( .D(Key[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[11]) );
  DFFSNQ_X1 \reg_key_reg[10]  ( .D(Key[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[10]) );
  DFFSNQ_X1 \reg_key_reg[9]  ( .D(Key[9]), .CLK(clk), .SN(1'b1), .Q(reg_key[9]) );
  DFFSNQ_X1 \reg_key_reg[8]  ( .D(Key[8]), .CLK(clk), .SN(1'b1), .Q(reg_key[8]) );
  DFFSNQ_X1 \reg_key_reg[7]  ( .D(Key[7]), .CLK(clk), .SN(1'b1), .Q(reg_key[7]) );
  DFFSNQ_X1 \reg_key_reg[6]  ( .D(Key[6]), .CLK(clk), .SN(1'b1), .Q(reg_key[6]) );
  DFFSNQ_X1 \reg_key_reg[5]  ( .D(Key[5]), .CLK(clk), .SN(1'b1), .Q(reg_key[5]) );
  DFFSNQ_X1 \reg_key_reg[4]  ( .D(Key[4]), .CLK(clk), .SN(1'b1), .Q(reg_key[4]) );
  DFFSNQ_X1 \reg_key_reg[3]  ( .D(Key[3]), .CLK(clk), .SN(1'b1), .Q(reg_key[3]) );
  DFFSNQ_X1 \reg_key_reg[2]  ( .D(Key[2]), .CLK(clk), .SN(1'b1), .Q(reg_key[2]) );
  DFFSNQ_X1 \reg_key_reg[1]  ( .D(Key[1]), .CLK(clk), .SN(1'b1), .Q(reg_key[1]) );
  DFFSNQ_X1 \reg_key_reg[0]  ( .D(Key[0]), .CLK(clk), .SN(1'b1), .Q(reg_key[0]) );
  DFFRNQ_X1 \Ciphertext_reg[181]  ( .D(reg_out[181]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[181]) );
  DFFRNQ_X1 \Ciphertext_reg[79]  ( .D(reg_out[79]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[79]) );
  DFFRNQ_X1 \Ciphertext_reg[165]  ( .D(reg_out[165]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[165]) );
  DFFRNQ_X1 \Ciphertext_reg[153]  ( .D(reg_out[153]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[153]) );
  DFFRNQ_X1 \Ciphertext_reg[80]  ( .D(reg_out[80]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[80]) );
  DFFRNQ_X1 \Ciphertext_reg[85]  ( .D(reg_out[85]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[85]) );
  DFFRNQ_X1 \Ciphertext_reg[152]  ( .D(reg_out[152]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[152]) );
  DFFRNQ_X1 \Ciphertext_reg[105]  ( .D(reg_out[105]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[105]) );
  DFFRNQ_X1 \Ciphertext_reg[185]  ( .D(reg_out[185]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[185]) );
  DFFRNQ_X1 \Ciphertext_reg[93]  ( .D(reg_out[93]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[93]) );
  DFFRNQ_X1 \Ciphertext_reg[146]  ( .D(reg_out[146]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[146]) );
  DFFRNQ_X1 \Ciphertext_reg[139]  ( .D(reg_out[139]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[139]) );
  DFFRNQ_X1 \Ciphertext_reg[69]  ( .D(reg_out[69]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[69]) );
  DFFRNQ_X1 \Ciphertext_reg[179]  ( .D(reg_out[179]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[179]) );
  DFFRNQ_X1 \Ciphertext_reg[50]  ( .D(reg_out[50]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[50]) );
  DFFRNQ_X1 \Ciphertext_reg[72]  ( .D(reg_out[72]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[72]) );
  DFFRNQ_X1 \Ciphertext_reg[39]  ( .D(reg_out[39]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[39]) );
  DFFRNQ_X1 \Ciphertext_reg[67]  ( .D(reg_out[67]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[67]) );
  DFFRNQ_X1 \Ciphertext_reg[54]  ( .D(reg_out[54]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[54]) );
  DFFRNQ_X1 \Ciphertext_reg[44]  ( .D(reg_out[44]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[44]) );
  DFFRNQ_X1 \Ciphertext_reg[184]  ( .D(reg_out[184]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[184]) );
  DFFRNQ_X1 \Ciphertext_reg[174]  ( .D(reg_out[174]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[174]) );
  DFFRNQ_X1 \Ciphertext_reg[134]  ( .D(reg_out[134]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[134]) );
  DFFRNQ_X1 \Ciphertext_reg[151]  ( .D(reg_out[151]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[151]) );
  DFFRNQ_X1 \Ciphertext_reg[35]  ( .D(reg_out[35]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[35]) );
  DFFRNQ_X1 \Ciphertext_reg[31]  ( .D(reg_out[31]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[31]) );
  DFFRNQ_X1 \Ciphertext_reg[109]  ( .D(reg_out[109]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[109]) );
  DFFRNQ_X1 \Ciphertext_reg[3]  ( .D(reg_out[3]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[3]) );
  DFFRNQ_X1 \Ciphertext_reg[84]  ( .D(reg_out[84]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[84]) );
  DFFRNQ_X1 \Ciphertext_reg[58]  ( .D(reg_out[58]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[58]) );
  DFFRNQ_X1 \Ciphertext_reg[145]  ( .D(reg_out[145]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[145]) );
  DFFRNQ_X1 \Ciphertext_reg[46]  ( .D(reg_out[46]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[46]) );
  DFFRNQ_X1 \Ciphertext_reg[71]  ( .D(reg_out[71]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[71]) );
  DFFRNQ_X1 \Ciphertext_reg[33]  ( .D(reg_out[33]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[33]) );
  DFFRNQ_X1 \Ciphertext_reg[183]  ( .D(reg_out[183]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[183]) );
  DFFRNQ_X1 \Ciphertext_reg[43]  ( .D(reg_out[43]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[43]) );
  DFFRNQ_X1 \Ciphertext_reg[182]  ( .D(reg_out[182]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[182]) );
  DFFRNQ_X1 \Ciphertext_reg[154]  ( .D(reg_out[154]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[154]) );
  DFFRNQ_X1 \Ciphertext_reg[22]  ( .D(reg_out[22]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[22]) );
  DFFRNQ_X1 \Ciphertext_reg[66]  ( .D(reg_out[66]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[66]) );
  DFFRNQ_X1 \Ciphertext_reg[86]  ( .D(reg_out[86]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[86]) );
  DFFRNQ_X1 \Ciphertext_reg[82]  ( .D(reg_out[82]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[82]) );
  DFFRNQ_X1 \Ciphertext_reg[68]  ( .D(reg_out[68]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[68]) );
  DFFRNQ_X1 \Ciphertext_reg[64]  ( .D(reg_out[64]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[64]) );
  DFFRNQ_X1 \Ciphertext_reg[6]  ( .D(reg_out[6]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[6]) );
  DFFRNQ_X1 \Ciphertext_reg[178]  ( .D(reg_out[178]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[178]) );
  DFFRNQ_X1 \Ciphertext_reg[148]  ( .D(reg_out[148]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[148]) );
  DFFRNQ_X1 \Ciphertext_reg[10]  ( .D(reg_out[10]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[10]) );
  DFFRNQ_X1 \Ciphertext_reg[171]  ( .D(reg_out[171]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[171]) );
  DFFRNQ_X1 \Ciphertext_reg[156]  ( .D(reg_out[156]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[156]) );
  DFFRNQ_X1 \Ciphertext_reg[30]  ( .D(reg_out[30]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[30]) );
  DFFRNQ_X1 \Ciphertext_reg[102]  ( .D(reg_out[102]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[102]) );
  DFFRNQ_X1 \Ciphertext_reg[155]  ( .D(reg_out[155]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[155]) );
  DFFRNQ_X1 \Ciphertext_reg[7]  ( .D(reg_out[7]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[7]) );
  DFFRNQ_X1 \Ciphertext_reg[76]  ( .D(reg_out[76]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[76]) );
  DFFRNQ_X1 \Ciphertext_reg[175]  ( .D(reg_out[175]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[175]) );
  DFFRNQ_X1 \Ciphertext_reg[57]  ( .D(reg_out[57]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[57]) );
  DFFRNQ_X1 \Ciphertext_reg[166]  ( .D(reg_out[166]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[166]) );
  DFFRNQ_X1 \Ciphertext_reg[63]  ( .D(reg_out[63]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[63]) );
  DFFRNQ_X1 \Ciphertext_reg[90]  ( .D(reg_out[90]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[90]) );
  DFFRNQ_X1 \Ciphertext_reg[163]  ( .D(reg_out[163]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[163]) );
  DFFRNQ_X1 \Ciphertext_reg[162]  ( .D(reg_out[162]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[162]) );
  DFFRNQ_X1 \Ciphertext_reg[113]  ( .D(reg_out[113]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[113]) );
  DFFRNQ_X1 \Ciphertext_reg[77]  ( .D(reg_out[77]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[77]) );
  DFFRNQ_X1 \Ciphertext_reg[150]  ( .D(reg_out[150]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[150]) );
  DFFRNQ_X1 \Ciphertext_reg[83]  ( .D(reg_out[83]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[83]) );
  DFFRNQ_X1 \Ciphertext_reg[176]  ( .D(reg_out[176]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[176]) );
  DFFRNQ_X1 \Ciphertext_reg[149]  ( .D(reg_out[149]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[149]) );
  DFFRNQ_X1 \Ciphertext_reg[60]  ( .D(reg_out[60]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[60]) );
  DFFRNQ_X1 \Ciphertext_reg[118]  ( .D(reg_out[118]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[118]) );
  DFFRNQ_X1 \Ciphertext_reg[94]  ( .D(reg_out[94]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[94]) );
  DFFRNQ_X1 \Ciphertext_reg[73]  ( .D(reg_out[73]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[73]) );
  DFFRNQ_X1 \Ciphertext_reg[74]  ( .D(reg_out[74]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[74]) );
  DFFRNQ_X1 \Ciphertext_reg[47]  ( .D(reg_out[47]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[47]) );
  DFFRNQ_X1 \Ciphertext_reg[144]  ( .D(reg_out[144]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[144]) );
  DFFRNQ_X1 \Ciphertext_reg[13]  ( .D(reg_out[13]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[13]) );
  DFFRNQ_X1 \Ciphertext_reg[42]  ( .D(reg_out[42]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[42]) );
  DFFRNQ_X1 \Ciphertext_reg[37]  ( .D(reg_out[37]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[37]) );
  DFFRNQ_X1 \Ciphertext_reg[132]  ( .D(reg_out[132]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[132]) );
  DFFRNQ_X1 \Ciphertext_reg[78]  ( .D(reg_out[78]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[78]) );
  DFFRNQ_X1 \Ciphertext_reg[133]  ( .D(reg_out[133]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[133]) );
  DFFRNQ_X1 \Ciphertext_reg[103]  ( .D(reg_out[103]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[103]) );
  DFFRNQ_X1 \Ciphertext_reg[164]  ( .D(reg_out[164]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[164]) );
  DFFRNQ_X1 \Ciphertext_reg[38]  ( .D(reg_out[38]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[38]) );
  DFFRNQ_X1 \Ciphertext_reg[115]  ( .D(reg_out[115]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[115]) );
  DFFRNQ_X1 \Ciphertext_reg[27]  ( .D(reg_out[27]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[27]) );
  DFFRNQ_X1 \Ciphertext_reg[70]  ( .D(reg_out[70]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[70]) );
  DFFRNQ_X1 \Ciphertext_reg[36]  ( .D(reg_out[36]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[36]) );
  DFFRNQ_X1 \Ciphertext_reg[180]  ( .D(reg_out[180]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[180]) );
  DFFRNQ_X1 \Ciphertext_reg[41]  ( .D(reg_out[41]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[41]) );
  DFFRNQ_X1 \Ciphertext_reg[23]  ( .D(reg_out[23]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[23]) );
  DFFRNQ_X1 \Ciphertext_reg[173]  ( .D(reg_out[173]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[173]) );
  DFFRNQ_X1 \Ciphertext_reg[123]  ( .D(reg_out[123]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[123]) );
  DFFRNQ_X1 \Ciphertext_reg[4]  ( .D(reg_out[4]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[4]) );
  DFFRNQ_X1 \Ciphertext_reg[119]  ( .D(reg_out[119]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[119]) );
  DFFRNQ_X1 \Ciphertext_reg[8]  ( .D(reg_out[8]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[8]) );
  DFFRNQ_X1 \Ciphertext_reg[161]  ( .D(reg_out[161]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[161]) );
  DFFRNQ_X1 \Ciphertext_reg[14]  ( .D(reg_out[14]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[14]) );
  DFFRNQ_X1 \Ciphertext_reg[136]  ( .D(reg_out[136]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[136]) );
  DFFRNQ_X1 \Ciphertext_reg[108]  ( .D(reg_out[108]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[108]) );
  DFFRNQ_X1 \Ciphertext_reg[29]  ( .D(reg_out[29]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[29]) );
  DFFRNQ_X1 \Ciphertext_reg[28]  ( .D(reg_out[28]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[28]) );
  DFFRNQ_X1 \Ciphertext_reg[40]  ( .D(reg_out[40]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[40]) );
  DFFRNQ_X1 \Ciphertext_reg[49]  ( .D(reg_out[49]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[49]) );
  DFFRNQ_X1 \Ciphertext_reg[117]  ( .D(reg_out[117]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[117]) );
  DFFRNQ_X1 \Ciphertext_reg[158]  ( .D(reg_out[158]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[158]) );
  DFFRNQ_X1 \Ciphertext_reg[137]  ( .D(reg_out[137]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[137]) );
  DFFRNQ_X1 \Ciphertext_reg[0]  ( .D(reg_out[0]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[0]) );
  DFFRNQ_X1 \Ciphertext_reg[11]  ( .D(reg_out[11]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[11]) );
  DFFRNQ_X1 \Ciphertext_reg[75]  ( .D(reg_out[75]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[75]) );
  DFFRNQ_X1 \Ciphertext_reg[159]  ( .D(reg_out[159]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[159]) );
  DFFRNQ_X1 \Ciphertext_reg[65]  ( .D(reg_out[65]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[65]) );
  DFFRNQ_X1 \Ciphertext_reg[56]  ( .D(reg_out[56]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[56]) );
  DFFRNQ_X1 \Ciphertext_reg[168]  ( .D(reg_out[168]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[168]) );
  DFFRNQ_X1 \Ciphertext_reg[5]  ( .D(reg_out[5]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[5]) );
  DFFRNQ_X1 \Ciphertext_reg[157]  ( .D(reg_out[157]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[157]) );
  DFFRNQ_X1 \Ciphertext_reg[140]  ( .D(reg_out[140]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[140]) );
  DFFRNQ_X1 \Ciphertext_reg[52]  ( .D(reg_out[52]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[52]) );
  DFFRNQ_X1 \Ciphertext_reg[53]  ( .D(reg_out[53]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[53]) );
  DFFRNQ_X1 \Ciphertext_reg[55]  ( .D(reg_out[55]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[55]) );
  DFFRNQ_X1 \Ciphertext_reg[34]  ( .D(reg_out[34]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[34]) );
  DFFRNQ_X1 \Ciphertext_reg[160]  ( .D(reg_out[160]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[160]) );
  DFFRNQ_X1 \Ciphertext_reg[104]  ( .D(reg_out[104]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[104]) );
  DFFRNQ_X1 \Ciphertext_reg[135]  ( .D(reg_out[135]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[135]) );
  DFFRNQ_X1 \Ciphertext_reg[120]  ( .D(reg_out[120]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[120]) );
  DFFRNQ_X1 \Ciphertext_reg[188]  ( .D(reg_out[188]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[188]) );
  DFFRNQ_X1 \Ciphertext_reg[12]  ( .D(reg_out[12]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[12]) );
  DFFRNQ_X1 \Ciphertext_reg[20]  ( .D(reg_out[20]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[20]) );
  DFFRNQ_X1 \Ciphertext_reg[62]  ( .D(reg_out[62]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[62]) );
  DFFRNQ_X1 \Ciphertext_reg[19]  ( .D(reg_out[19]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[19]) );
  DFFRNQ_X1 \Ciphertext_reg[167]  ( .D(reg_out[167]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[167]) );
  DFFRNQ_X1 \Ciphertext_reg[143]  ( .D(reg_out[143]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[143]) );
  DFFRNQ_X1 \Ciphertext_reg[48]  ( .D(reg_out[48]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[48]) );
  DFFRNQ_X1 \Ciphertext_reg[45]  ( .D(reg_out[45]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[45]) );
  DFFRNQ_X1 \Ciphertext_reg[59]  ( .D(reg_out[59]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[59]) );
  DFFRNQ_X1 \Ciphertext_reg[172]  ( .D(reg_out[172]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[172]) );
  DFFRNQ_X1 \Ciphertext_reg[89]  ( .D(reg_out[89]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[89]) );
  DFFRNQ_X1 \Ciphertext_reg[16]  ( .D(reg_out[16]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[16]) );
  DFFRNQ_X1 \Ciphertext_reg[18]  ( .D(reg_out[18]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[18]) );
  DFFRNQ_X1 \Ciphertext_reg[51]  ( .D(reg_out[51]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[51]) );
  DFFRNQ_X1 \Ciphertext_reg[141]  ( .D(reg_out[141]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[141]) );
  DFFRNQ_X1 \Ciphertext_reg[32]  ( .D(reg_out[32]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[32]) );
  DFFRNQ_X1 \Ciphertext_reg[87]  ( .D(reg_out[87]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[87]) );
  DFFRNQ_X1 \Ciphertext_reg[15]  ( .D(reg_out[15]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[15]) );
  DFFRNQ_X1 \Ciphertext_reg[61]  ( .D(reg_out[61]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[61]) );
  DFFRNQ_X1 \Ciphertext_reg[170]  ( .D(reg_out[170]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[170]) );
  DFFRNQ_X1 \Ciphertext_reg[21]  ( .D(reg_out[21]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[21]) );
  DFFRNQ_X1 \Ciphertext_reg[142]  ( .D(reg_out[142]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[142]) );
  DFFRNQ_X1 \Ciphertext_reg[169]  ( .D(reg_out[169]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[169]) );
  DFFRNQ_X1 \Ciphertext_reg[92]  ( .D(reg_out[92]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[92]) );
  DFFRNQ_X1 \Ciphertext_reg[17]  ( .D(reg_out[17]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[17]) );
  DFFRNQ_X1 \Ciphertext_reg[177]  ( .D(reg_out[177]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[177]) );
  DFFRNQ_X1 \Ciphertext_reg[138]  ( .D(reg_out[138]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[138]) );
  DFFRNQ_X1 \Ciphertext_reg[187]  ( .D(reg_out[187]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[187]) );
  DFFRNQ_X1 \Ciphertext_reg[81]  ( .D(reg_out[81]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[81]) );
  DFFRNQ_X1 \Ciphertext_reg[111]  ( .D(reg_out[111]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[111]) );
  DFFRNQ_X1 \Ciphertext_reg[110]  ( .D(reg_out[110]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[110]) );
  DFFRNQ_X1 \Ciphertext_reg[25]  ( .D(reg_out[25]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[25]) );
  DFFRNQ_X1 \Ciphertext_reg[189]  ( .D(reg_out[189]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[189]) );
  DFFRNQ_X1 \Ciphertext_reg[124]  ( .D(reg_out[124]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[124]) );
  DFFRNQ_X1 \Ciphertext_reg[106]  ( .D(reg_out[106]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[106]) );
  DFFRNQ_X1 \Ciphertext_reg[88]  ( .D(reg_out[88]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[88]) );
  DFFRNQ_X1 \Ciphertext_reg[95]  ( .D(reg_out[95]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[95]) );
  DFFRNQ_X1 \Ciphertext_reg[107]  ( .D(reg_out[107]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[107]) );
  DFFRNQ_X1 \Ciphertext_reg[1]  ( .D(reg_out[1]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[1]) );
  DFFRNQ_X1 \Ciphertext_reg[91]  ( .D(reg_out[91]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[91]) );
  DFFRNQ_X1 \Ciphertext_reg[26]  ( .D(reg_out[26]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[26]) );
  DFFRNQ_X1 \Ciphertext_reg[2]  ( .D(reg_out[2]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[2]) );
  DFFRNQ_X1 \Ciphertext_reg[112]  ( .D(reg_out[112]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[112]) );
  DFFRNQ_X1 \Ciphertext_reg[24]  ( .D(reg_out[24]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[24]) );
  DFFRNQ_X1 \Ciphertext_reg[9]  ( .D(reg_out[9]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[9]) );
  DFFRNQ_X1 \Ciphertext_reg[129]  ( .D(reg_out[129]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[129]) );
  DFFRNQ_X1 \Ciphertext_reg[114]  ( .D(reg_out[114]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[114]) );
  DFFRNQ_X1 \Ciphertext_reg[122]  ( .D(reg_out[122]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[122]) );
  DFFRNQ_X1 \Ciphertext_reg[130]  ( .D(reg_out[130]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[130]) );
  DFFRNQ_X1 \Ciphertext_reg[126]  ( .D(reg_out[126]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[126]) );
  DFFRNQ_X1 \Ciphertext_reg[186]  ( .D(reg_out[186]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[186]) );
  DFFRNQ_X1 \Ciphertext_reg[97]  ( .D(reg_out[97]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[97]) );
  DFFRNQ_X1 \Ciphertext_reg[191]  ( .D(reg_out[191]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[191]) );
  DFFRNQ_X1 \Ciphertext_reg[121]  ( .D(reg_out[121]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[121]) );
  DFFRNQ_X1 \Ciphertext_reg[190]  ( .D(reg_out[190]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[190]) );
  DFFRNQ_X1 \Ciphertext_reg[131]  ( .D(reg_out[131]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[131]) );
  DFFRNQ_X1 \Ciphertext_reg[125]  ( .D(reg_out[125]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[125]) );
  DFFRNQ_X1 \Ciphertext_reg[116]  ( .D(reg_out[116]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[116]) );
  DFFRNQ_X1 \Ciphertext_reg[128]  ( .D(reg_out[128]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[128]) );
  DFFRNQ_X1 \Ciphertext_reg[127]  ( .D(reg_out[127]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[127]) );
  DFFRNQ_X1 \Ciphertext_reg[98]  ( .D(reg_out[98]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[98]) );
  DFFRNQ_X1 \Ciphertext_reg[100]  ( .D(reg_out[100]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[100]) );
  DFFRNQ_X1 \Ciphertext_reg[96]  ( .D(reg_out[96]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[96]) );
  DFFRNQ_X1 \Ciphertext_reg[99]  ( .D(reg_out[99]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[99]) );
  DFFRNQ_X1 \Ciphertext_reg[101]  ( .D(reg_out[101]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[101]) );
  DFFRNQ_X1 \Ciphertext_reg[147]  ( .D(reg_out[147]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[147]) );
  SPEEDY_Rounds6_0 SPEEDY_instance ( .Plaintext(reg_in), .Key(reg_key), 
        .Ciphertext(reg_out) );
endmodule

