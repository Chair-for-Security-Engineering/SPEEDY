library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SB is
    Port ( input : in STD_LOGIC_VECTOR (5 downto 0);
           output : out STD_LOGIC_VECTOR (5 downto 0));
end SB;

architecture Behavioral of SB is

begin

    with input select
    output <= "001000" when "000000",
              "000000" when "000001",
              "001001" when "000010",
              "000011" when "000011",
              "111000" when "000100",
              "010000" when "000101",
              "101001" when "000110",
              "010011" when "000111",
              "001100" when "001000",
              "001101" when "001001",
              "000100" when "001010",
              "000111" when "001011",
              "110000" when "001100",
              "000001" when "001101",
              "100000" when "001110",
              "100011" when "001111",
              "011010" when "010000",
              "010010" when "010001",
              "011000" when "010010",
              "110010" when "010011",
              "111110" when "010100",
              "010110" when "010101",
              "101100" when "010110",
              "110110" when "010111",
              "011100" when "011000",
              "011101" when "011001",
              "010100" when "011010",
              "110111" when "011011",
              "110100" when "011100",
              "000101" when "011101",
              "100100" when "011110",
              "100111" when "011111",
              "000010" when "100000",
              "000110" when "100001",
              "001011" when "100010",
              "001111" when "100011",
              "110011" when "100100",
              "010111" when "100101",
              "100001" when "100110",
              "010101" when "100111",
              "001010" when "101000",
              "011011" when "101001",
              "001110" when "101010",
              "011111" when "101011",
              "110001" when "101100",
              "010001" when "101101",
              "100101" when "101110",
              "110101" when "101111",
              "100010" when "110000",
              "100110" when "110001",
              "101010" when "110010",
              "101110" when "110011",
              "111010" when "110100",
              "011110" when "110101",
              "101000" when "110110",
              "111100" when "110111",
              "101011" when "111000",
              "111011" when "111001",
              "101111" when "111010",
              "111111" when "111011",
              "111001" when "111100",
              "011001" when "111101",
              "101101" when "111110",
              "111101" when others;

end Behavioral;