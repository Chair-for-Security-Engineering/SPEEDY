
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_SPEEDY_Top is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_SPEEDY_Top;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Rounds5_0 is

   port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : out
         std_logic_vector (191 downto 0));

end SPEEDY_Rounds5_0;

architecture SYN_Behavioral of SPEEDY_Rounds5_0 is

   component OAI21_X2
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( I0, I1, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X12
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X4
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X8
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X8
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5, n8, n11, n13, n14, n19, n20, n23, n25, n30, n33, n34, n35, 
      n36, n41, n45, n47, n50, n51, n53, n56, n57, n58, n60, n61, n62, n63, n65
      , n67, n68, n72, n73, n74, n75, n76, n78, n79, n82, n84, n87, n89, n92, 
      n94, n95, n97, n100, n102, n103, n110, n111, n113, n114, n116, n120, n121
      , n123, n124, n125, n126, n128, n132, n133, n135, n136, n137, n139, n142,
      n143, n145, n147, n148, n149, n150, n153, n155, n159, n161, n162, n166, 
      n167, n170, n171, n172, n173, n174, n175, n180, n182, n183, n184, n188, 
      n190, n193, n194, n195, n198, n199, n201, n203, n204, n205, n206, n209, 
      n210, n211, n212, n213, n215, n216, n217, n218, n220, n224, n229, n231, 
      n233, n235, n237, n238, n242, n243, n247, n248, n249, n250, n251, n252, 
      n253, n254, n256, n257, n260, n263, n265, n266, n270, n272, n273, n274, 
      n275, n277, n278, n280, n281, n283, n287, n288, n293, n294, n295, n299, 
      n300, n301, n302, n303, n304, n305, n308, n309, n311, n315, n316, n319, 
      n322, n323, n327, n329, n333, n334, n336, n337, n338, n341, n347, n348, 
      n350, n356, n357, n359, n360, n361, n369, n370, n372, n375, n376, n379, 
      n383, n385, n386, n390, n391, n401, n402, n404, n406, n407, n413, n415, 
      n421, n422, n427, n431, n434, n437, n438, n442, n443, n444, n446, n447, 
      n448, n450, n451, n452, n454, n456, n457, n458, n460, n461, n463, n464, 
      n465, n467, n469, n473, n476, n477, n479, n480, n481, n482, n484, n488, 
      n489, n491, n492, n500, n502, n503, n505, n506, n507, n508, n510, n511, 
      n514, n516, n517, n521, n523, n524, n527, n529, n531, n532, n534, n535, 
      n536, n537, n538, n539, n540, n542, n543, n544, n545, n546, n548, n549, 
      n550, n552, n553, n554, n556, n558, n559, n560, n561, n562, n563, n564, 
      n566, n567, n569, n571, n573, n574, n575, n576, n577, n578, n580, n584, 
      n587, n589, n590, n592, n594, n595, n596, n597, n598, n599, n600, n602, 
      n603, n604, n605, n606, n608, n609, n610, n611, n612, n613, n615, n616, 
      n617, n619, n620, n622, n624, n625, n626, n627, n628, n630, n631, n632, 
      n633, n634, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, 
      n647, n649, n650, n652, n653, n655, n656, n657, n658, n659, n663, n664, 
      n665, n666, n668, n669, n670, n671, n672, n674, n675, n677, n679, n680, 
      n682, n683, n684, n686, n687, n689, n690, n692, n693, n694, n696, n698, 
      n699, n703, n704, n705, n708, n709, n713, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n727, n728, n729, n730, n731, n732, n733, 
      n734, n735, n736, n737, n738, n739, n740, n741, n742, n744, n745, n748, 
      n749, n751, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n769, n770, n772, n773, n774, n775, n777, n778, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n802, n803, n806, 
      n807, n808, n809, n810, n811, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n838, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n855, n856, n857, n858, n859, 
      n860, n863, n864, n865, n866, n867, n868, n869, n873, n874, n875, n877, 
      n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n890, n891, 
      n892, n894, n896, n897, n898, n899, n900, n901, n902, n904, n905, n906, 
      n907, n908, n910, n912, n913, n914, n915, n918, n919, n920, n921, n922, 
      n923, n924, n925, n927, n928, n929, n932, n933, n934, n935, n936, n937, 
      n939, n940, n943, n944, n945, n946, n948, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n964, n965, n966, n967, n968, 
      n969, n971, n972, n974, n975, n976, n977, n978, n979, n980, n981, n982, 
      n984, n985, n986, n987, n988, n989, n990, n992, n993, n994, n996, n997, 
      n998, n999, n1000, n1001, n1003, n1004, n1005, n1006, n1009, n1010, n1011
      , n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, 
      n1022, n1023, n1024, n1025, n1026, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1045, 
      n1046, n1047, n1048, n1049, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1058, n1059, n1061, n1062, n1064, n1065, n1067, n1068, n1070, n1071, 
      n1072, n1073, n1074, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1087, n1090, n1091, n1092, n1094, n1096, n1097, 
      n1098, n1099, n1101, n1102, n1103, n1104, n1105, n1106, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1125, n1127, n1128, n1129, n1130, n1131, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1140, n1142, n1149, n1150, n1152, 
      n1153, n1154, n1156, n1158, n1159, n1163, n1164, n1165, n1166, n1167, 
      n1168, n1169, n1172, n1174, n1175, n1177, n1179, n1180, n1184, n1185, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1197, n1198, 
      n1199, n1200, n1202, n1203, n1207, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1219, n1222, n1223, n1224, n1227, n1228, 
      n1229, n1231, n1232, n1233, n1234, n1235, n1237, n1241, n1242, n1243, 
      n1246, n1247, n1251, n1252, n1253, n1255, n1256, n1257, n1258, n1259, 
      n1260, n1261, n1262, n1263, n1264, n1266, n1267, n1268, n1269, n1270, 
      n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, 
      n1281, n1283, n1284, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1313, 
      n1314, n1316, n1317, n1318, n1319, n1320, n1321, n1325, n1326, n1328, 
      n1329, n1330, n1331, n1334, n1335, n1338, n1339, n1342, n1348, n1349, 
      n1350, n1353, n1354, n1355, n1357, n1358, n1359, n1362, n1363, n1364, 
      n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, 
      n1376, n1377, n1378, n1380, n1381, n1383, n1385, n1387, n1389, n1392, 
      n1396, n1397, n1398, n1400, n1401, n1402, n1403, n1406, n1407, n1408, 
      n1410, n1411, n1412, n1413, n1415, n1416, n1418, n1419, n1420, n1421, 
      n1422, n1424, n1425, n1428, n1429, n1431, n1435, n1436, n1437, n1438, 
      n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1451, n1454, 
      n1455, n1457, n1458, n1459, n1460, n1464, n1465, n1468, n1470, n1472, 
      n1473, n1475, n1478, n1480, n1481, n1483, n1485, n1489, n1491, n1493, 
      n1494, n1495, n1496, n1497, n1499, n1500, n1502, n1503, n1504, n1506, 
      n1512, n1513, n1515, n1516, n1517, n1518, n1519, n1520, n1525, n1526, 
      n1527, n1530, n1534, n1535, n1536, n1539, n1540, n1541, n1543, n1544, 
      n1545, n1546, n1547, n1548, n1550, n1551, n1557, n1558, n1562, n1563, 
      n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1572, n1573, n1577, 
      n1579, n1580, n1581, n1582, n1583, n1585, n1587, n1588, n1589, n1591, 
      n1593, n1595, n1596, n1597, n1598, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1613, n1616, n1617, n1618, 
      n1622, n1624, n1626, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1637, n1638, n1639, n1640, n1642, n1643, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1655, n1658, n1659, n1661, n1664, 
      n1665, n1667, n1671, n1676, n1679, n1680, n1681, n1683, n1684, n1685, 
      n1687, n1689, n1690, n1692, n1693, n1696, n1697, n1699, n1701, n1703, 
      n1704, n1706, n1709, n1710, n1711, n1712, n1713, n1715, n1716, n1717, 
      n1718, n1720, n1721, n1722, n1725, n1726, n1727, n1728, n1729, n1731, 
      n1732, n1733, n1734, n1737, n1738, n1739, n1741, n1742, n1743, n1746, 
      n1748, n1749, n1750, n1755, n1756, n1757, n1758, n1759, n1760, n1761, 
      n1763, n1764, n1765, n1767, n1768, n1769, n1771, n1772, n1776, n1777, 
      n1780, n1783, n1784, n1785, n1786, n1789, n1790, n1791, n1792, n1793, 
      n1794, n1795, n1797, n1798, n1799, n1800, n1801, n1802, n1804, n1806, 
      n1807, n1809, n1811, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1824, n1825, n1831, n1832, n1833, n1834, n1835, n1839, n1840, n1841, 
      n1842, n1843, n1845, n1846, n1848, n1851, n1853, n1854, n1856, n1858, 
      n1859, n1863, n1864, n1865, n1866, n1869, n1870, n1872, n1874, n1875, 
      n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1886, n1887, 
      n1888, n1890, n1891, n1892, n1893, n1895, n1896, n1897, n1898, n1902, 
      n1905, n1906, n1908, n1911, n1912, n1914, n1916, n1918, n1919, n1920, 
      n1922, n1923, n1924, n1925, n1926, n1927, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1937, n1938, n1940, n1943, n1944, n1946, n1947, n1948, 
      n1949, n1950, n1951, n1952, n1954, n1955, n1956, n1959, n1960, n1961, 
      n1964, n1965, n1966, n1968, n1970, n1974, n1975, n1976, n1977, n1980, 
      n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1990, n1991, 
      n1992, n1994, n1995, n1996, n1997, n1998, n2004, n2007, n2012, n2013, 
      n2015, n2016, n2018, n2019, n2020, n2021, n2023, n2025, n2026, n2029, 
      n2031, n2034, n2035, n2036, n2037, n2038, n2039, n2041, n2044, n2045, 
      n2047, n2049, n2051, n2052, n2057, n2060, n2061, n2062, n2064, n2065, 
      n2068, n2070, n2071, n2072, n2074, n2076, n2079, n2081, n2082, n2083, 
      n2084, n2085, n2086, n2087, n2091, n2093, n2094, n2095, n2097, n2098, 
      n2099, n2100, n2101, n2102, n2105, n2108, n2109, n2110, n2111, n2114, 
      n2115, n2116, n2118, n2120, n2121, n2123, n2124, n2126, n2127, n2128, 
      n2129, n2131, n2132, n2133, n2135, n2136, n2137, n2138, n2139, n2140, 
      n2145, n2147, n2148, n2149, n2150, n2154, n2155, n2156, n2157, n2158, 
      n2159, n2160, n2161, n2163, n2164, n2167, n2168, n2170, n2171, n2173, 
      n2174, n2176, n2177, n2178, n2179, n2181, n2183, n2184, n2185, n2188, 
      n2189, n2190, n2191, n2192, n2193, n2195, n2198, n2199, n2201, n2202, 
      n2203, n2206, n2208, n2209, n2210, n2212, n2213, n2214, n2215, n2218, 
      n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2228, n2230, n2231, 
      n2232, n2233, n2234, n2235, n2236, n2238, n2245, n2247, n2248, n2249, 
      n2251, n2252, n2253, n2254, n2256, n2257, n2258, n2261, n2262, n2264, 
      n2265, n2266, n2268, n2271, n2273, n2274, n2276, n2277, n2278, n2279, 
      n2281, n2282, n2283, n2284, n2285, n2287, n2290, n2292, n2293, n2294, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2306, n2307, 
      n2308, n2309, n2311, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
      n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2328, n2329, n2331, 
      n2337, n2339, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, 
      n2350, n2351, n2352, n2353, n2356, n2357, n2358, n2359, n2361, n2362, 
      n2363, n2365, n2366, n2367, n2369, n2370, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2385, n2388, n2389, n2390, 
      n2391, n2394, n2395, n2396, n2398, n2399, n2401, n2403, n2404, n2405, 
      n2406, n2407, n2409, n2410, n2413, n2415, n2418, n2420, n2422, n2423, 
      n2425, n2427, n2430, n2432, n2433, n2434, n2435, n2436, n2437, n2439, 
      n2440, n2441, n2444, n2445, n2447, n2448, n2449, n2450, n2452, n2453, 
      n2454, n2455, n2457, n2458, n2459, n2460, n2462, n2463, n2465, n2466, 
      n2467, n2469, n2470, n2471, n2472, n2474, n2476, n2477, n2478, n2481, 
      n2482, n2483, n2484, n2487, n2488, n2490, n2491, n2492, n2495, n2496, 
      n2497, n2499, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, 
      n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, 
      n2520, n2522, n2523, n2524, n2525, n2527, n2528, n2529, n2530, n2533, 
      n2536, n2537, n2538, n2540, n2541, n2542, n2543, n2544, n2545, n2549, 
      n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2560, n2561, 
      n2562, n2563, n2564, n2565, n2566, n2567, n2569, n2570, n2571, n2572, 
      n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2581, n2582, n2585, 
      n2586, n2587, n2588, n2590, n2591, n2592, n2594, n2595, n2596, n2597, 
      n2599, n2602, n2603, n2604, n2605, n2607, n2609, n2610, n2611, n2614, 
      n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
      n2626, n2627, n2629, n2631, n2632, n2633, n2635, n2636, n2639, n2641, 
      n2642, n2647, n2648, n2649, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2658, n2659, n2660, n2661, n2664, n2665, n2666, n2667, n2668, n2670, 
      n2671, n2673, n2675, n2676, n2679, n2680, n2681, n2686, n2687, n2689, 
      n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
      n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2708, n2709, n2710, 
      n2711, n2712, n2713, n2716, n2717, n2718, n2719, n2722, n2723, n2725, 
      n2726, n2727, n2728, n2729, n2730, n2733, n2735, n2736, n2739, n2740, 
      n2742, n2743, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, 
      n2753, n2754, n2755, n2756, n2757, n2759, n2760, n2761, n2762, n2765, 
      n2766, n2767, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2798, n2799, 
      n2800, n2802, n2804, n2805, n2808, n2809, n2811, n2812, n2813, n2814, 
      n2815, n2816, n2817, n2818, n2820, n2823, n2824, n2825, n2826, n2827, 
      n2828, n2829, n2831, n2832, n2833, n2834, n2835, n2837, n2838, n2840, 
      n2841, n2842, n2844, n2848, n2850, n2852, n2853, n2855, n2857, n2858, 
      n2862, n2863, n2864, n2865, n2868, n2869, n2871, n2872, n2873, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2884, n2885, n2886, n2887, 
      n2888, n2889, n2890, n2891, n2894, n2895, n2897, n2898, n2900, n2901, 
      n2902, n2903, n2904, n2906, n2908, n2910, n2911, n2912, n2914, n2915, 
      n2916, n2919, n2920, n2921, n2922, n2925, n2927, n2928, n2934, n2936, 
      n2937, n2938, n2939, n2941, n2944, n2945, n2946, n2947, n2948, n2949, 
      n2950, n2952, n2953, n2955, n2956, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2964, n2965, n2966, n2967, n2971, n2973, n2974, n2975, n2976, 
      n2978, n2979, n2980, n2981, n2982, n2985, n2986, n2989, n2990, n2991, 
      n2993, n2994, n2995, n2997, n2998, n2999, n3000, n3001, n3003, n3005, 
      n3006, n3007, n3009, n3010, n3012, n3013, n3014, n3015, n3016, n3017, 
      n3018, n3019, n3020, n3022, n3029, n3030, n3031, n3032, n3033, n3034, 
      n3036, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3053, n3054, n3057, n3059, n3060, n3062, n3063, n3067, n3070, 
      n3071, n3072, n3073, n3074, n3076, n3077, n3078, n3080, n3081, n3082, 
      n3083, n3084, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3099, n3100, n3101, n3102, n3105, n3106, n3107, 
      n3109, n3110, n3112, n3113, n3115, n3118, n3119, n3121, n3122, n3123, 
      n3124, n3125, n3128, n3132, n3133, n3134, n3138, n3141, n3144, n3146, 
      n3147, n3150, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, 
      n3160, n3163, n3164, n3165, n3166, n3170, n3171, n3172, n3173, n3175, 
      n3176, n3178, n3179, n3181, n3182, n3186, n3190, n3193, n3195, n3196, 
      n3198, n3199, n3202, n3203, n3204, n3205, n3207, n3211, n3212, n3215, 
      n3216, n3217, n3218, n3219, n3220, n3221, n3223, n3224, n3225, n3226, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3238, n3239, 
      n3243, n3249, n3251, n3255, n3259, n3260, n3261, n3262, n3267, n3268, 
      n3269, n3271, n3272, n3273, n3275, n3276, n3277, n3278, n3279, n3283, 
      n3286, n3288, n3289, n3290, n3291, n3292, n3293, n3296, n3297, n3298, 
      n3299, n3300, n3302, n3303, n3304, n3310, n3312, n3313, n3315, n3316, 
      n3317, n3319, n3323, n3325, n3326, n3329, n3330, n3331, n3335, n3336, 
      n3338, n3342, n3343, n3344, n3346, n3347, n3348, n3350, n3351, n3353, 
      n3355, n3356, n3358, n3360, n3361, n3362, n3363, n3364, n3368, n3369, 
      n3370, n3372, n3373, n3376, n3380, n3382, n3383, n3386, n3387, n3388, 
      n3389, n3390, n3391, n3392, n3394, n3398, n3399, n3401, n3404, n3405, 
      n3406, n3410, n3411, n3414, n3415, n3416, n3417, n3418, n3419, n3422, 
      n3423, n3424, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, 
      n3435, n3437, n3438, n3439, n3440, n3442, n3443, n3448, n3451, n3452, 
      n3454, n3456, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3467, n3469, n3470, n3473, n3474, n3477, n3479, n3480, n3481, n3484, 
      n3486, n3487, n3489, n3490, n3491, n3493, n3494, n3495, n3496, n3497, 
      n3499, n3501, n3502, n3504, n3505, n3506, n3508, n3509, n3510, n3511, 
      n3514, n3515, n3516, n3517, n3518, n3521, n3524, n3525, n3527, n3529, 
      n3530, n3531, n3533, n3534, n3535, n3537, n3538, n3539, n3540, n3541, 
      n3544, n3545, n3547, n3549, n3550, n3551, n3552, n3553, n3554, n3556, 
      n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
      n3567, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3578, 
      n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3590, 
      n3592, n3593, n3594, n3595, n3597, n3598, n3600, n3601, n3602, n3603, 
      n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, 
      n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3627, n3629, n3631, 
      n3633, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, 
      n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3654, n3655, n3657, 
      n3658, n3660, n3661, n3662, n3663, n3664, n3665, n3667, n3668, n3670, 
      n3671, n3674, n3675, n3676, n3678, n3682, n3684, n3685, n3686, n3688, 
      n3691, n3693, n3694, n3695, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3710, n3711, n3716, n3717, n3723, 
      n3724, n3725, n3726, n3727, n3728, n3729, n3731, n3732, n3733, n3734, 
      n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3744, n3745, 
      n3746, n3748, n3751, n3752, n3753, n3754, n3755, n3756, n3759, n3760, 
      n3762, n3763, n3764, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3775, n3777, n3778, n3779, n3780, n3783, n3786, n3787, n3788, 
      n3789, n3790, n3792, n3793, n3794, n3797, n3798, n3799, n3801, n3802, 
      n3803, n3806, n3807, n3808, n3809, n3810, n3812, n3814, n3815, n3816, 
      n3818, n3820, n3821, n3822, n3824, n3825, n3826, n3828, n3830, n3832, 
      n3833, n3834, n3835, n3836, n3838, n3839, n3840, n3843, n3845, n3846, 
      n3847, n3848, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3861, n3862, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3872, 
      n3873, n3874, n3875, n3877, n3878, n3879, n3880, n3882, n3883, n3885, 
      n3886, n3887, n3889, n3891, n3893, n3895, n3897, n3898, n3899, n3900, 
      n3902, n3903, n3905, n3906, n3908, n3910, n3913, n3914, n3916, n3918, 
      n3920, n3921, n3923, n3925, n3927, n3928, n3929, n3932, n3933, n3934, 
      n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3943, n3945, n3946, 
      n3948, n3949, n3953, n3954, n3956, n3958, n3959, n3960, n3961, n3963, 
      n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3974, 
      n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, 
      n3986, n3988, n3989, n3990, n3991, n3992, n3994, n3995, n3996, n3997, 
      n4001, n4002, n4005, n4006, n4010, n4013, n4014, n4015, n4016, n4018, 
      n4019, n4020, n4021, n4022, n4025, n4026, n4028, n4029, n4030, n4031, 
      n4032, n4034, n4035, n4038, n4040, n4043, n4044, n4045, n4048, n4049, 
      n4050, n4051, n4053, n4054, n4055, n4057, n4058, n4059, n4060, n4062, 
      n4063, n4064, n4067, n4068, n4069, n4070, n4071, n4072, n4074, n4075, 
      n4076, n4077, n4079, n4080, n4081, n4082, n4084, n4085, n4086, n4087, 
      n4088, n4089, n4090, n4091, n4093, n4094, n4095, n4096, n4097, n4098, 
      n4100, n4101, n4103, n4104, n4106, n4107, n4108, n4109, n4110, n4111, 
      n4112, n4113, n4114, n4115, n4116, n4118, n4119, n4120, n4121, n4122, 
      n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4131, n4132, n4133, 
      n4136, n4137, n4138, n4140, n4143, n4147, n4150, n4151, n4155, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4168, 
      n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4178, n4179, n4180, 
      n4181, n4182, n4183, n4184, n4185, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4197, n4198, n4199, n4200, n4201, n4203, n4204, n4206, 
      n4208, n4209, n4211, n4212, n4215, n4217, n4222, n4223, n4224, n4225, 
      n4226, n4227, n4228, n4231, n4234, n4236, n4237, n4238, n4239, n4241, 
      n4244, n4245, n4246, n4247, n4250, n4252, n4253, n4254, n4255, n4256, 
      n4258, n4259, n4260, n4262, n4263, n4264, n4265, n4267, n4268, n4269, 
      n4271, n4272, n4273, n4274, n4277, n4279, n4280, n4281, n4282, n4285, 
      n4286, n4287, n4288, n4290, n4291, n4292, n4293, n4294, n4295, n4296, 
      n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, 
      n4310, n4311, n4314, n4315, n4317, n4318, n4319, n4320, n4321, n4324, 
      n4326, n4327, n4328, n4329, n4331, n4332, n4333, n4334, n4337, n4339, 
      n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4348, n4351, n4353, 
      n4354, n4355, n4356, n4357, n4358, n4360, n4361, n4362, n4364, n4366, 
      n4370, n4371, n4372, n4373, n4375, n4376, n4377, n4378, n4379, n4380, 
      n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, 
      n4391, n4392, n4393, n4394, n4395, n4397, n4398, n4399, n4401, n4402, 
      n4403, n4404, n4405, n4409, n4410, n4411, n4412, n4413, n4414, n4415, 
      n4416, n4417, n4420, n4422, n4423, n4424, n4425, n4426, n4427, n4428, 
      n4430, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, 
      n4441, n4442, n4443, n4445, n4446, n4447, n4448, n4449, n4450, n4452, 
      n4453, n4455, n4456, n4457, n4458, n4459, n4461, n4462, n4463, n4465, 
      n4469, n4470, n4471, n4472, n4474, n4475, n4478, n4479, n4480, n4481, 
      n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4490, n4491, n4493, 
      n4495, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, 
      n4507, n4508, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, 
      n4520, n4521, n4522, n4524, n4525, n4530, n4531, n4532, n4533, n4534, 
      n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, 
      n4546, n4548, n4549, n4552, n4553, n4554, n4555, n4556, n4557, n4558, 
      n4559, n4560, n4561, n4563, n4564, n4565, n4566, n4568, n4574, n4575, 
      n4577, n4580, n4581, n4582, n4585, n4587, n4589, n4590, n4591, n4592, 
      n4593, n4595, n4596, n4597, n4601, n4604, n4605, n4606, n4607, n4608, 
      n4609, n4610, n4611, n4613, n4615, n4618, n4619, n4620, n4621, n4622, 
      n4623, n4624, n4625, n4626, n4627, n4628, n4630, n4631, n4632, n4633, 
      n4634, n4635, n4636, n4637, n4638, n4639, n4642, n4644, n4645, n4647, 
      n4648, n4649, n4650, n4653, n4654, n4655, n4656, n4657, n4658, n4659, 
      n4660, n4661, n4662, n4664, n4665, n4667, n4668, n4669, n4673, n4674, 
      n4675, n4679, n4680, n4681, n4683, n4684, n4685, n4686, n4687, n4688, 
      n4689, n4690, n4696, n4697, n4698, n4701, n4702, n4703, n4704, n4705, 
      n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4715, n4716, n4719, 
      n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4728, n4729, n4730, 
      n4731, n4734, n4735, n4736, n4737, n4738, n4739, n4742, n4743, n4744, 
      n4747, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4759, 
      n4760, n4761, n4762, n4763, n4764, n4766, n4767, n4768, n4770, n4771, 
      n4774, n4775, n4776, n4777, n4779, n4780, n4781, n4782, n4783, n4784, 
      n4786, n4787, n4788, n4789, n4790, n4791, n4793, n4794, n4795, n4797, 
      n4798, n4799, n4800, n4801, n4802, n4803, n4805, n4807, n4808, n4809, 
      n4810, n4811, n4812, n4813, n4814, n4816, n4819, n4820, n4821, n4822, 
      n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4832, n4833, n4834, 
      n4836, n4837, n4838, n4839, n4840, n4841, n4843, n4844, n4846, n4847, 
      n4848, n4849, n4850, n4851, n4852, n4857, n4858, n4859, n4860, n4861, 
      n4864, n4865, n4866, n4867, n4869, n4870, n4871, n4873, n4875, n4876, 
      n4877, n4878, n4879, n4880, n4881, n4883, n4885, n4887, n4888, n4889, 
      n4890, n4891, n4892, n4893, n4895, n4896, n4897, n4898, n4899, n4901, 
      n4903, n4904, n4905, n4907, n4908, n4910, n4911, n4912, n4914, n4915, 
      n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4925, n4926, n4928, 
      n4929, n4931, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, 
      n4942, n4943, n4945, n4947, n4949, n4950, n4952, n4953, n4954, n4956, 
      n4957, n4958, n4959, n4960, n4961, n4964, n4965, n4966, n4967, n4969, 
      n4970, n4972, n4973, n4974, n4976, n4981, n4983, n4984, n4985, n4986, 
      n4987, n4988, n4990, n4992, n4993, n4994, n4995, n4996, n4998, n4999, 
      n5000, n5001, n5002, n5004, n5005, n5007, n5008, n5009, n5010, n5011, 
      n5012, n5013, n5014, n5015, n5016, n5020, n5021, n5022, n5024, n5025, 
      n5026, n5028, n5029, n5030, n5031, n5034, n5036, n5037, n5038, n5040, 
      n5042, n5043, n5044, n5045, n5047, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5055, n5057, n5059, n5060, n5061, n5062, n5063, n5064, n5065, 
      n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, 
      n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5089, 
      n5090, n5092, n5093, n5095, n5096, n5097, n5098, n5099, n5100, n5102, 
      n5103, n5105, n5108, n5109, n5110, n5112, n5113, n5114, n5115, n5116, 
      n5117, n5118, n5120, n5121, n5122, n5124, n5125, n5126, n5127, n5129, 
      n5130, n5131, n5133, n5134, n5138, n5139, n5140, n5141, n5142, n5143, 
      n5144, n5145, n5146, n5147, n5149, n5150, n5152, n5153, n5159, n5161, 
      n5163, n5164, n5165, n5166, n5168, n5169, n5171, n5172, n5173, n5174, 
      n5176, n5178, n5179, n5182, n5186, n5187, n5188, n5189, n5192, n5194, 
      n5195, n5196, n5197, n5198, n5202, n5203, n5204, n5205, n5206, n5209, 
      n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5218, n5221, n5222, 
      n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5234, n5235, 
      n5236, n5238, n5240, n5243, n5244, n5245, n5246, n5247, n5248, n5249, 
      n5250, n5251, n5252, n5253, n5254, n5257, n5258, n5261, n5263, n5264, 
      n5265, n5266, n5268, n5271, n5272, n5274, n5275, n5277, n5280, n5281, 
      n5282, n5283, n5285, n5287, n5288, n5289, n5291, n5292, n5294, n5295, 
      n5296, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, 
      n5307, n5308, n5310, n5311, n5312, n5314, n5315, n5316, n5317, n5320, 
      n5324, n5325, n5326, n5327, n5328, n5331, n5332, n5333, n5334, n5335, 
      n5338, n5341, n5342, n5344, n5345, n5346, n5349, n5350, n5351, n5353, 
      n5354, n5355, n5357, n5359, n5360, n5361, n5362, n5363, n5367, n5368, 
      n5369, n5370, n5371, n5373, n5375, n5376, n5378, n5379, n5381, n5382, 
      n5388, n5391, n5393, n5394, n5395, n5396, n5398, n5400, n5401, n5402, 
      n5403, n5406, n5407, n5408, n5409, n5412, n5413, n5415, n5416, n5417, 
      n5420, n5421, n5424, n5425, n5429, n5432, n5433, n5434, n5435, n5438, 
      n5439, n5441, n5442, n5445, n5446, n5447, n5448, n5449, n5450, n5452, 
      n5454, n5455, n5456, n5457, n5458, n5459, n5461, n5462, n5463, n5464, 
      n5467, n5468, n5471, n5473, n5474, n5475, n5478, n5479, n5480, n5481, 
      n5482, n5483, n5486, n5488, n5489, n5490, n5491, n5492, n5494, n5497, 
      n5499, n5500, n5502, n5503, n5505, n5506, n5509, n5510, n5511, n5512, 
      n5513, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, 
      n5525, n5529, n5530, n5531, n5532, n5535, n5537, n5539, n5540, n5541, 
      n5542, n5543, n5545, n5547, n5550, n5554, n5556, n5557, n5558, n5559, 
      n5560, n5561, n5562, n5563, n5566, n5568, n5569, n5570, n5571, n5573, 
      n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5582, n5583, n5584, 
      n5585, n5586, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, 
      n5596, n5597, n5599, n5600, n5601, n5602, n5603, n5605, n5606, n5609, 
      n5610, n5612, n5613, n5614, n5615, n5616, n5617, n5619, n5621, n5623, 
      n5624, n5625, n5626, n5627, n5630, n5631, n5632, n5634, n5637, n5639, 
      n5642, n5645, n5646, n5647, n5648, n5649, n5652, n5653, n5655, n5656, 
      n5658, n5659, n5660, n5662, n5663, n5664, n5666, n5667, n5668, n5669, 
      n5670, n5673, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, 
      n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5693, 
      n5696, n5697, n5698, n5700, n5701, n5702, n5704, n5705, n5706, n5707, 
      n5708, n5709, n5710, n5711, n5712, n5713, n5715, n5716, n5718, n5721, 
      n5722, n5724, n5725, n5726, n5727, n5729, n5730, n5731, n5732, n5734, 
      n5736, n5738, n5739, n5740, n5741, n5742, n5744, n5746, n5748, n5749, 
      n5750, n5751, n5752, n5753, n5755, n5756, n5757, n5759, n5760, n5761, 
      n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5771, n5772, n5773, 
      n5775, n5776, n5777, n5779, n5780, n5781, n5782, n5783, n5784, n5785, 
      n5786, n5788, n5789, n5790, n5792, n5793, n5796, n5797, n5798, n5799, 
      n5801, n5804, n5805, n5806, n5807, n5808, n5809, n5811, n5812, n5813, 
      n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5823, n5825, n5826, 
      n5827, n5828, n5830, n5833, n5834, n5835, n5836, n5837, n5838, n5839, 
      n5840, n5841, n5844, n5845, n5847, n5849, n5850, n5852, n5853, n5854, 
      n5856, n5858, n5859, n5860, n5861, n5862, n5865, n5866, n5867, n5868, 
      n5870, n5871, n5872, n5874, n5875, n5876, n5877, n5879, n5880, n5881, 
      n5883, n5884, n5885, n5887, n5889, n5890, n5892, n5894, n5895, n5896, 
      n5897, n5900, n5903, n5904, n5905, n5906, n5908, n5909, n5910, n5911, 
      n5912, n5913, n5914, n5915, n5917, n5919, n5920, n5921, n5922, n5923, 
      n5926, n5927, n5928, n5929, n5930, n5931, n5934, n5936, n5937, n5938, 
      n5939, n5940, n5941, n5942, n5943, n5944, n5946, n5949, n5950, n5951, 
      n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5961, n5962, 
      n5963, n5964, n5965, n5967, n5969, n5971, n5972, n5973, n5974, n5977, 
      n5978, n5981, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
      n5993, n5994, n5995, n5997, n5999, n6001, n6004, n6005, n6006, n6007, 
      n6013, n6014, n6015, n6018, n6019, n6021, n6022, n6024, n6025, n6026, 
      n6029, n6030, n6031, n6034, n6035, n6037, n6038, n6040, n6041, n6042, 
      n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, 
      n6056, n6057, n6058, n6059, n6060, n6062, n6063, n6064, n6065, n6066, 
      n6068, n6070, n6071, n6073, n6074, n6075, n6076, n6077, n6080, n6081, 
      n6082, n6085, n6087, n6089, n6090, n6091, n6092, n6095, n6096, n6097, 
      n6098, n6101, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6112, 
      n6113, n6115, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6126, 
      n6129, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6140, 
      n6141, n6142, n6143, n6144, n6145, n6147, n6148, n6149, n6150, n6152, 
      n6154, n6155, n6157, n6158, n6159, n6160, n6162, n6164, n6166, n6168, 
      n6169, n6170, n6171, n6173, n6174, n6175, n6176, n6177, n6179, n6180, 
      n6181, n6182, n6183, n6185, n6186, n6188, n6189, n6190, n6191, n6192, 
      n6193, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6205, 
      n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, 
      n6216, n6217, n6218, n6219, n6220, n6223, n6226, n6229, n6231, n6232, 
      n6233, n6234, n6235, n6236, n6237, n6239, n6240, n6241, n6242, n6243, 
      n6245, n6246, n6247, n6248, n6249, n6251, n6253, n6254, n6255, n6256, 
      n6257, n6258, n6259, n6260, n6262, n6263, n6264, n6265, n6268, n6269, 
      n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, 
      n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6291, 
      n6293, n6294, n6295, n6296, n6297, n6298, n6301, n6303, n6304, n6306, 
      n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, 
      n6317, n6318, n6319, n6320, n6321, n6323, n6327, n6330, n6332, n6334, 
      n6336, n6338, n6339, n6342, n6344, n6345, n6346, n6347, n6348, n6349, 
      n6351, n6353, n6354, n6355, n6359, n6362, n6364, n6365, n6367, n6368, 
      n6369, n6370, n6371, n6372, n6373, n6375, n6376, n6377, n6378, n6379, 
      n6380, n6381, n6382, n6384, n6385, n6386, n6387, n6388, n6389, n6391, 
      n6392, n6393, n6394, n6395, n6396, n6397, n6399, n6400, n6402, n6403, 
      n6405, n6406, n6407, n6408, n6410, n6413, n6415, n6416, n6417, n6418, 
      n6419, n6420, n6421, n6422, n6423, n6425, n6426, n6427, n6428, n6429, 
      n6430, n6432, n6433, n6434, n6435, n6438, n6439, n6440, n6442, n6443, 
      n6444, n6445, n6447, n6449, n6451, n6452, n6453, n6455, n6456, n6457, 
      n6459, n6460, n6462, n6463, n6465, n6466, n6469, n6470, n6471, n6472, 
      n6473, n6475, n6476, n6477, n6479, n6480, n6481, n6482, n6483, n6484, 
      n6485, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, 
      n6496, n6498, n6500, n6501, n6502, n6503, n6504, n6507, n6508, n6509, 
      n6511, n6512, n6513, n6515, n6516, n6517, n6518, n6520, n6522, n6523, 
      n6525, n6528, n6529, n6530, n6533, n6534, n6535, n6536, n6538, n6539, 
      n6540, n6541, n6542, n6543, n6545, n6547, n6548, n6549, n6550, n6551, 
      n6552, n6554, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, 
      n6567, n6568, n6570, n6571, n6572, n6573, n6574, n6575, n6581, n6582, 
      n6584, n6585, n6586, n6588, n6589, n6590, n6591, n6592, n6593, n6594, 
      n6595, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, 
      n6606, n6608, n6611, n6612, n6614, n6615, n6616, n6617, n6618, n6619, 
      n6620, n6621, n6622, n6624, n6625, n6627, n6628, n6629, n6630, n6631, 
      n6633, n6634, n6635, n6637, n6638, n6640, n6642, n6643, n6644, n6646, 
      n6647, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, 
      n6658, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6668, n6670, 
      n6672, n6673, n6675, n6676, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6695, 
      n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, 
      n6708, n6709, n6712, n6713, n6716, n6718, n6719, n6722, n6725, n6727, 
      n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, 
      n6739, n6740, n6743, n6744, n6745, n6746, n6748, n6749, n6751, n6752, 
      n6753, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6770, n6773, n6774, n6775, n6776, 
      n6777, n6778, n6779, n6780, n6782, n6783, n6784, n6786, n6788, n6789, 
      n6790, n6791, n6792, n6794, n6795, n6798, n6799, n6800, n6801, n6802, 
      n6803, n6804, n6805, n6806, n6808, n6809, n6811, n6812, n6813, n6814, 
      n6815, n6819, n6820, n6821, n6822, n6823, n6825, n6826, n6827, n6830, 
      n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
      n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, 
      n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, 
      n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6874, n6875, 
      n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6885, n6886, n6887, 
      n6889, n6891, n6892, n6893, n6894, n6895, n6897, n6898, n6902, n6903, 
      n6904, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6916, 
      n6917, n6921, n6923, n6924, n6925, n6926, n6927, n6928, n6930, n6931, 
      n6932, n6933, n6934, n6935, n6936, n6937, n6939, n6941, n6943, n6944, 
      n6945, n6946, n6951, n6952, n6954, n6955, n6957, n6958, n6959, n6960, 
      n6962, n6964, n6965, n6966, n6967, n6968, n6969, n6972, n6975, n6976, 
      n6977, n6978, n6979, n6981, n6982, n6983, n6984, n6985, n6986, n6987, 
      n6991, n6996, n6997, n6998, n6999, n7000, n7002, n7003, n7004, n7007, 
      n7008, n7009, n7010, n7011, n7012, n7014, n7015, n7016, n7017, n7018, 
      n7022, n7023, n7025, n7027, n7029, n7030, n7031, n7032, n7033, n7036, 
      n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7046, n7047, 
      n7048, n7050, n7052, n7053, n7054, n7055, n7057, n7059, n7060, n7061, 
      n7062, n7063, n7064, n7065, n7067, n7068, n7069, n7071, n7072, n7073, 
      n7074, n7076, n7077, n7078, n7079, n7080, n7082, n7084, n7085, n7086, 
      n7087, n7088, n7090, n7091, n7092, n7094, n7095, n7096, n7097, n7099, 
      n7100, n7102, n7103, n7105, n7106, n7107, n7108, n7110, n7112, n7113, 
      n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7122, n7123, n7124, 
      n7125, n7126, n7129, n7130, n7131, n7132, n7134, n7138, n7140, n7142, 
      n7143, n7144, n7145, n7147, n7148, n7150, n7151, n7152, n7153, n7154, 
      n7155, n7156, n7158, n7162, n7165, n7167, n7168, n7169, n7170, n7171, 
      n7174, n7175, n7176, n7178, n7180, n7181, n7182, n7183, n7184, n7185, 
      n7186, n7187, n7189, n7190, n7192, n7193, n7194, n7196, n7199, n7200, 
      n7201, n7203, n7204, n7209, n7211, n7212, n7213, n7215, n7218, n7219, 
      n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7231, 
      n7232, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7244, 
      n7245, n7247, n7248, n7250, n7251, n7252, n7253, n7254, n7255, n7256, 
      n7257, n7258, n7260, n7261, n7263, n7264, n7265, n7266, n7267, n7268, 
      n7269, n7270, n7271, n7274, n7275, n7276, n7277, n7279, n7280, n7281, 
      n7282, n7284, n7285, n7288, n7289, n7291, n7293, n7294, n7296, n7298, 
      n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7307, n7308, n7309, 
      n7311, n7312, n7313, n7314, n7315, n7317, n7319, n7320, n7321, n7322, 
      n7323, n7324, n7325, n7326, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7336, n7338, n7339, n7340, n7341, n7342, n7345, n7346, n7347, n7348, 
      n7349, n7350, n7351, n7354, n7355, n7356, n7357, n7358, n7359, n7361, 
      n7362, n7363, n7364, n7365, n7368, n7370, n7371, n7372, n7374, n7375, 
      n7376, n7377, n7378, n7379, n7381, n7382, n7383, n7384, n7385, n7386, 
      n7387, n7388, n7390, n7391, n7395, n7396, n7397, n7398, n7399, n7403, 
      n7405, n7406, n7407, n7408, n7409, n7411, n7412, n7413, n7416, n7418, 
      n7420, n7421, n7422, n7423, n7424, n7425, n7427, n7428, n7429, n7430, 
      n7431, n7432, n7433, n7435, n7437, n7440, n7441, n7442, n7443, n7445, 
      n7446, n7447, n7449, n7450, n7451, n7452, n7453, n7454, n7456, n7457, 
      n7458, n7460, n7463, n7464, n7466, n7467, n7468, n7471, n7472, n7474, 
      n7475, n7476, n7478, n7480, n7481, n7482, n7483, n7484, n7485, n7486, 
      n7487, n7492, n7495, n7496, n7497, n7498, n7499, n7500, n7502, n7503, 
      n7506, n7507, n7509, n7510, n7513, n7514, n7515, n7516, n7517, n7518, 
      n7520, n7522, n7523, n7524, n7525, n7526, n7527, n7529, n7530, n7531, 
      n7533, n7535, n7536, n7537, n7539, n7540, n7541, n7542, n7543, n7545, 
      n7546, n7547, n7548, n7551, n7552, n7553, n7554, n7555, n7556, n7557, 
      n7559, n7560, n7561, n7562, n7563, n7565, n7566, n7567, n7568, n7569, 
      n7570, n7571, n7577, n7578, n7581, n7582, n7583, n7584, n7585, n7586, 
      n7587, n7588, n7589, n7590, n7591, n7592, n7594, n7595, n7596, n7597, 
      n7598, n7599, n7601, n7602, n7603, n7604, n7605, n7607, n7608, n7609, 
      n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, 
      n7621, n7622, n7625, n7628, n7629, n7630, n7631, n7634, n7635, n7636, 
      n7638, n7639, n7640, n7644, n7645, n7647, n7648, n7649, n7650, n7651, 
      n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, 
      n7662, n7663, n7664, n7665, n7667, n7668, n7671, n7672, n7673, n7675, 
      n7676, n7677, n7678, n7679, n7681, n7682, n7684, n7687, n7688, n7689, 
      n7690, n7691, n7693, n7694, n7695, n7696, n7697, n7698, n7700, n7701, 
      n7702, n7703, n7704, n7705, n7706, n7707, n7709, n7710, n7711, n7712, 
      n7713, n7714, n7715, n7716, n7717, n7720, n7721, n7722, n7723, n7725, 
      n7726, n7727, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7737, 
      n7738, n7739, n7740, n7741, n7742, n7744, n7745, n7748, n7749, n7750, 
      n7751, n7752, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7762, 
      n7763, n7764, n7767, n7769, n7770, n7771, n7772, n7774, n7776, n7778, 
      n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, 
      n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, 
      n7801, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7811, n7812, 
      n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, 
      n7823, n7824, n7825, n7826, n7827, n7830, n7831, n7832, n7833, n7834, 
      n7835, n7836, n7837, n7839, n7840, n7841, n7843, n7844, n7845, n7846, 
      n7848, n7849, n7850, n7852, n7854, n7855, n7856, n7857, n7858, n7859, 
      n7861, n7862, n7864, n7865, n7867, n7868, n7869, n7870, n7873, n7874, 
      n7875, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, 
      n7886, n7887, n7888, n7890, n7893, n7894, n7895, n7896, n7897, n7898, 
      n7899, n7900, n7901, n7902, n7903, n7904, n7906, n7907, n7908, n7910, 
      n7911, n7912, n7913, n7914, n7916, n7917, n7918, n7919, n7921, n7922, 
      n7923, n7925, n7927, n7930, n7931, n7932, n7933, n7934, n7935, n7937, 
      n7938, n7939, n7940, n7941, n7942, n7944, n7945, n7946, n7947, n7948, 
      n7949, n7950, n7951, n7952, n7954, n7955, n7956, n7957, n7960, n7961, 
      n7963, n7964, n7965, n7966, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7975, n7976, n7977, n7978, n7980, n7981, n7982, n7983, n7984, n7985, 
      n7986, n7987, n7988, n7990, n7991, n7994, n7995, n7996, n7998, n7999, 
      n8000, n8001, n8002, n8003, n8004, n8006, n8007, n8009, n8010, n8011, 
      n8012, n8013, n8016, n8017, n8018, n8019, n8021, n8022, n8024, n8025, 
      n8026, n8027, n8029, n8030, n8031, n8032, n8033, n8035, n8037, n8039, 
      n8040, n8041, n8042, n8043, n8044, n8045, n8048, n8049, n8050, n8051, 
      n8052, n8054, n8057, n8059, n8060, n8063, n8064, n8069, n8070, n8071, 
      n8072, n8073, n8075, n8077, n8079, n8080, n8082, n8083, n8084, n8085, 
      n8086, n8087, n8088, n8089, n8090, n8091, n8093, n8094, n8095, n8097, 
      n8098, n8099, n8100, n8102, n8106, n8107, n8108, n8109, n8111, n8112, 
      n8113, n8114, n8115, n8117, n8118, n8119, n8120, n8121, n8122, n8123, 
      n8125, n8126, n8127, n8128, n8130, n8131, n8132, n8133, n8134, n8135, 
      n8137, n8138, n8139, n8140, n8143, n8144, n8145, n8146, n8147, n8148, 
      n8149, n8150, n8151, n8152, n8154, n8155, n8156, n8157, n8160, n8161, 
      n8162, n8163, n8165, n8166, n8167, n8169, n8171, n8172, n8173, n8174, 
      n8175, n8177, n8178, n8180, n8181, n8182, n8183, n8184, n8185, n8186, 
      n8187, n8190, n8191, n8192, n8193, n8194, n8195, n8197, n8198, n8199, 
      n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8211, 
      n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, 
      n8222, n8223, n8224, n8225, n8226, n8227, n8230, n8232, n8233, n8234, 
      n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8244, n8245, 
      n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, 
      n8256, n8257, n8259, n8260, n8262, n8263, n8264, n8265, n8267, n8268, 
      n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, 
      n8280, n8281, n8283, n8286, n8287, n8290, n8293, n8295, n8299, n8300, 
      n8301, n8303, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8318, n8319, n8320, n8321, n8322, n8323, n8325, 
      n8326, n8327, n8329, n8330, n8331, n8332, n8333, n8335, n8337, n8338, 
      n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, 
      n8351, n8354, n8357, n8358, n8359, n8361, n8363, n8365, n8366, n8367, 
      n8370, n8371, n8372, n8373, n8374, n8377, n8378, n8379, n8380, n8381, 
      n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8393, 
      n8396, n8398, n8399, n8401, n8405, n8406, n8407, n8408, n8409, n8410, 
      n8411, n8412, n8413, n8416, n8417, n8418, n8419, n8422, n8423, n8424, 
      n8425, n8428, n8429, n8430, n8431, n8432, n8433, n8435, n8436, n8438, 
      n8439, n8440, n8441, n8442, n8444, n8446, n8447, n8448, n8449, n8450, 
      n8451, n8452, n8453, n8459, n8461, n8462, n8463, n8464, n8467, n8468, 
      n8469, n8470, n8471, n8472, n8473, n8477, n8478, n8479, n8480, n8481, 
      n8482, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, 
      n8493, n8495, n8498, n8500, n8501, n8502, n8503, n8504, n8505, n8506, 
      n8507, n8508, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, 
      n8518, n8519, n8521, n8524, n8525, n8527, n8528, n8529, n8530, n8532, 
      n8533, n8534, n8535, n8536, n8538, n8541, n8542, n8543, n8544, n8545, 
      n8546, n8547, n8548, n8549, n8551, n8552, n8553, n8554, n8555, n8557, 
      n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8568, n8569, n8570, 
      n8573, n8574, n8575, n8576, n8579, n8580, n8581, n8582, n8584, n8585, 
      n8586, n8588, n8593, n8594, n8595, n8596, n8597, n8598, n8600, n8601, 
      n8602, n8603, n8604, n8605, n8608, n8609, n8610, n8611, n8612, n8613, 
      n8614, n8616, n8617, n8618, n8619, n8620, n8621, n8623, n8624, n8625, 
      n8626, n8627, n8628, n8629, n8630, n8632, n8635, n8636, n8637, n8638, 
      n8639, n8640, n8641, n8642, n8645, n8646, n8647, n8648, n8649, n8650, 
      n8651, n8652, n8654, n8655, n8656, n8657, n8658, n8660, n8661, n8663, 
      n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, 
      n8675, n8677, n8678, n8681, n8682, n8683, n8684, n8685, n8686, n8687, 
      n8688, n8689, n8690, n8691, n8692, n8694, n8695, n8696, n8697, n8698, 
      n8699, n8700, n8702, n8703, n8704, n8705, n8707, n8708, n8710, n8711, 
      n8714, n8716, n8717, n8721, n8722, n8723, n8724, n8726, n8727, n8728, 
      n8729, n8730, n8731, n8733, n8735, n8736, n8738, n8740, n8741, n8742, 
      n8745, n8746, n8748, n8749, n8750, n8751, n8753, n8754, n8755, n8756, 
      n8757, n8758, n8759, n8760, n8762, n8763, n8764, n8765, n8766, n8767, 
      n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8781, 
      n8782, n8784, n8786, n8788, n8789, n8790, n8792, n8793, n8794, n8795, 
      n8796, n8797, n8798, n8799, n8800, n8802, n8804, n8805, n8807, n8808, 
      n8810, n8811, n8812, n8814, n8815, n8816, n8817, n8819, n8820, n8821, 
      n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8831, n8832, 
      n8834, n8835, n8836, n8837, n8838, n8843, n8844, n8845, n8846, n8848, 
      n8849, n8851, n8852, n8853, n8854, n8855, n8857, n8858, n8860, n8861, 
      n8863, n8864, n8867, n8868, n8872, n8873, n8875, n8876, n8877, n8879, 
      n8880, n8881, n8882, n8883, n8884, n8885, n8887, n8888, n8889, n8890, 
      n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8900, n8901, n8902, 
      n8903, n8904, n8905, n8906, n8907, n8908, n8910, n8911, n8912, n8913, 
      n8914, n8915, n8916, n8917, n8921, n8922, n8923, n8925, n8926, n8927, 
      n8928, n8929, n8931, n8932, n8934, n8935, n8937, n8938, n8939, n8940, 
      n8943, n8944, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, 
      n8954, n8955, n8957, n8959, n8963, n8964, n8965, n8968, n8970, n8972, 
      n8974, n8976, n8978, n8980, n8982, n8983, n8984, n8985, n8986, n8988, 
      n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, 
      n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, 
      n9010, n9012, n9013, n9016, n9017, n9018, n9019, n9020, n9021, n9022, 
      n9023, n9024, n9025, n9026, n9027, n9029, n9030, n9031, n9032, n9034, 
      n9035, n9036, n9037, n9038, n9040, n9041, n9042, n9044, n9047, n9049, 
      n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, 
      n9060, n9062, n9063, n9065, n9070, n9071, n9072, n9073, n9074, n9076, 
      n9077, n9078, n9079, n9080, n9081, n9083, n9084, n9085, n9087, n9088, 
      n9089, n9092, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9102, 
      n9103, n9104, n9105, n9107, n9108, n9109, n9110, n9111, n9115, n9116, 
      n9117, n9119, n9121, n9123, n9124, n9125, n9129, n9130, n9131, n9132, 
      n9133, n9134, n9135, n9137, n9138, n9139, n9140, n9141, n9142, n9143, 
      n9144, n9145, n9147, n9148, n9149, n9150, n9152, n9154, n9156, n9157, 
      n9158, n9159, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, 
      n9173, n9174, n9175, n9176, n9178, n9179, n9180, n9181, n9186, n9188, 
      n9189, n9190, n9191, n9192, n9193, n9197, n9198, n9201, n9202, n9203, 
      n9204, n9205, n9210, n9211, n9214, n9215, n9216, n9217, n9218, n9219, 
      n9220, n9222, n9223, n9224, n9226, n9228, n9229, n9230, n9232, n9233, 
      n9234, n9236, n9237, n9241, n9242, n9244, n9248, n9249, n9250, n9252, 
      n9254, n9255, n9256, n9257, n9258, n9259, n9261, n9262, n9263, n9264, 
      n9265, n9266, n9267, n9268, n9269, n9270, n9272, n9273, n9274, n9275, 
      n9276, n9279, n9280, n9281, n9283, n9284, n9285, n9286, n9287, n9288, 
      n9289, n9292, n9294, n9295, n9296, n9298, n9301, n9302, n9304, n9305, 
      n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9314, n9315, n9316, 
      n9317, n9318, n9319, n9320, n9322, n9323, n9324, n9325, n9326, n9327, 
      n9328, n9329, n9330, n9331, n9332, n9333, n9335, n9337, n9338, n9339, 
      n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9348, n9349, n9350, 
      n9351, n9353, n9354, n9356, n9357, n9358, n9359, n9360, n9361, n9362, 
      n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, 
      n9373, n9374, n9376, n9377, n9378, n9379, n9381, n9382, n9383, n9384, 
      n9386, n9390, n9391, n9392, n9393, n9394, n9396, n9397, n9399, n9400, 
      n9401, n9402, n9405, n9407, n9408, n9409, n9410, n9411, n9414, n9417, 
      n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9429, 
      n9430, n9431, n9432, n9433, n9434, n9437, n9438, n9439, n9440, n9441, 
      n9443, n9445, n9446, n9447, n9449, n9450, n9451, n9452, n9453, n9454, 
      n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, 
      n9466, n9468, n9469, n9470, n9472, n9473, n9474, n9477, n9480, n9481, 
      n9482, n9483, n9484, n9485, n9489, n9490, n9493, n9494, n9495, n9497, 
      n9498, n9499, n9500, n9502, n9503, n9504, n9505, n9507, n9508, n9509, 
      n9510, n9511, n9512, n9513, n9514, n9517, n9518, n9519, n9520, n9521, 
      n9522, n9523, n9524, n9525, n9526, n9527, n9529, n9530, n9531, n9532, 
      n9533, n9534, n9535, n9536, n9538, n9539, n9541, n9542, n9543, n9544, 
      n9545, n9546, n9548, n9549, n9550, n9552, n9553, n9554, n9555, n9556, 
      n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9567, 
      n9568, n9569, n9570, n9571, n9573, n9574, n9575, n9576, n9577, n9578, 
      n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9588, n9590, n9593, 
      n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9602, n9603, n9604, 
      n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, 
      n9615, n9616, n9617, n9618, n9619, n9620, n9627, n9628, n9629, n9630, 
      n9631, n9632, n9634, n9635, n9636, n9637, n9638, n9640, n9641, n9642, 
      n9644, n9645, n9646, n9648, n9650, n9651, n9652, n9653, n9654, n9655, 
      n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9667, n9668, 
      n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, 
      n9680, n9682, n9683, n9684, n9686, n9687, n9689, n9690, n9691, n9692, 
      n9694, n9696, n9697, n9698, n9699, n9701, n9702, n9704, n9705, n9706, 
      n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9718, 
      n9719, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9730, n9731, 
      n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, 
      n9742, n9743, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9753, 
      n9754, n9756, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9766, 
      n9767, n9768, n9769, n9771, n9772, n9773, n9774, n9775, n9776, n9778, 
      n9779, n9780, n9784, n9785, n9786, n9787, n9789, n9790, n9791, n9792, 
      n9793, n9794, n9797, n9799, n9800, n9801, n9802, n9803, n9804, n9805, 
      n9807, n9809, n9811, n9812, n9813, n9814, n9819, n9820, n9822, n9823, 
      n9825, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9836, n9840, 
      n9841, n9842, n9845, n9846, n9847, n9848, n9850, n9851, n9854, n9855, 
      n9856, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, 
      n9867, n9868, n9869, n9870, n9871, n9873, n9875, n9876, n9877, n9878, 
      n9879, n9880, n9881, n9887, n9888, n9889, n9891, n9892, n9893, n9894, 
      n9896, n9898, n9899, n9900, n9902, n9903, n9904, n9905, n9906, n9907, 
      n9910, n9911, n9912, n9914, n9916, n9917, n9918, n9919, n9920, n9921, 
      n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9932, 
      n9933, n9934, n9939, n9943, n9945, n9946, n9948, n9949, n9950, n9952, 
      n9955, n9956, n9957, n9960, n9961, n9964, n9965, n9966, n9967, n9969, 
      n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, 
      n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9989, n9990, 
      n9991, n9992, n9993, n9994, n9995, n9996, n9998, n9999, n10000, n10001, 
      n10002, n10004, n10007, n10008, n10009, n10011, n10012, n10013, n10014, 
      n10015, n10016, n10018, n10019, n10023, n10024, n10025, n10026, n10027, 
      n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, 
      n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10045, n10046, 
      n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10055, n10056, 
      n10057, n10058, n10059, n10061, n10062, n10063, n10064, n10066, n10067, 
      n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, 
      n10078, n10080, n10081, n10082, n10083, n10084, n10086, n10087, n10088, 
      n10090, n10091, n10093, n10094, n10095, n10096, n10097, n10100, n10101, 
      n10103, n10104, n10105, n10107, n10111, n10112, n10114, n10116, n10117, 
      n10118, n10119, n10121, n10122, n10123, n10124, n10125, n10126, n10128, 
      n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10139, n10140, 
      n10141, n10142, n10144, n10145, n10146, n10147, n10149, n10150, n10151, 
      n10152, n10153, n10154, n10155, n10156, n10159, n10160, n10161, n10163, 
      n10164, n10165, n10167, n10168, n10169, n10170, n10171, n10173, n10174, 
      n10175, n10176, n10177, n10178, n10179, n10181, n10182, n10183, n10186, 
      n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, 
      n10196, n10197, n10201, n10202, n10203, n10204, n10205, n10206, n10207, 
      n10208, n10209, n10210, n10211, n10213, n10214, n10215, n10216, n10217, 
      n10220, n10221, n10222, n10224, n10225, n10226, n10227, n10228, n10229, 
      n10230, n10231, n10232, n10234, n10236, n10237, n10238, n10239, n10240, 
      n10241, n10242, n10243, n10246, n10248, n10249, n10250, n10251, n10252, 
      n10253, n10254, n10255, n10257, n10258, n10259, n10260, n10261, n10263, 
      n10264, n10265, n10267, n10268, n10269, n10270, n10271, n10272, n10273, 
      n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10284, 
      n10285, n10287, n10288, n10289, n10291, n10293, n10294, n10295, n10296, 
      n10297, n10298, n10299, n10300, n10301, n10303, n10304, n10305, n10310, 
      n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, 
      n10320, n10321, n10322, n10323, n10327, n10328, n10329, n10331, n10332, 
      n10333, n10335, n10337, n10338, n10339, n10341, n10344, n10345, n10346, 
      n10347, n10348, n10350, n10351, n10352, n10355, n10356, n10357, n10358, 
      n10359, n10360, n10362, n10363, n10364, n10365, n10366, n10367, n10369, 
      n10370, n10371, n10372, n10373, n10374, n10376, n10378, n10379, n10382, 
      n10383, n10385, n10387, n10388, n10389, n10390, n10391, n10392, n10393, 
      n10394, n10395, n10396, n10397, n10399, n10400, n10401, n10405, n10409, 
      n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10422, n10423, 
      n10425, n10427, n10428, n10430, n10431, n10432, n10433, n10435, n10436, 
      n10437, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10447, 
      n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, 
      n10458, n10460, n10461, n10462, n10464, n10465, n10466, n10467, n10469, 
      n10470, n10474, n10475, n10477, n10478, n10479, n10480, n10481, n10482, 
      n10483, n10484, n10486, n10487, n10488, n10490, n10491, n10492, n10493, 
      n10494, n10495, n10497, n10498, n10499, n10500, n10501, n10502, n10503, 
      n10504, n10505, n10507, n10508, n10509, n10510, n10512, n10513, n10514, 
      n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10524, 
      n10525, n10526, n10527, n10529, n10530, n10531, n10532, n10533, n10534, 
      n10535, n10536, n10537, n10538, n10539, n10541, n10542, n10543, n10544, 
      n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10554, 
      n10555, n10556, n10557, n10558, n10559, n10561, n10562, n10563, n10564, 
      n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10573, n10574, 
      n10575, n10576, n10577, n10578, n10579, n10580, n10582, n10583, n10584, 
      n10585, n10586, n10587, n10588, n10591, n10593, n10594, n10595, n10596, 
      n10597, n10598, n10599, n10601, n10602, n10603, n10604, n10605, n10608, 
      n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, 
      n10618, n10620, n10621, n10622, n10623, n10627, n10629, n10630, n10631, 
      n10632, n10634, n10635, n10636, n10638, n10639, n10640, n10641, n10642, 
      n10643, n10646, n10647, n10648, n10649, n10650, n10652, n10654, n10655, 
      n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, 
      n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, 
      n10677, n10678, n10680, n10681, n10683, n10684, n10685, n10686, n10687, 
      n10688, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, 
      n10698, n10700, n10701, n10702, n10704, n10705, n10707, n10708, n10709, 
      n10710, n10711, n10713, n10714, n10715, n10716, n10717, n10720, n10721, 
      n10724, n10725, n10727, n10728, n10729, n10730, n10732, n10733, n10734, 
      n10735, n10736, n10737, n10739, n10740, n10741, n10742, n10743, n10745, 
      n10746, n10747, n10748, n10749, n10751, n10752, n10754, n10755, n10756, 
      n10759, n10761, n10763, n10764, n10766, n10767, n10768, n10770, n10771, 
      n10772, n10773, n10774, n10775, n10777, n10779, n10780, n10783, n10784, 
      n10785, n10786, n10787, n10789, n10790, n10791, n10792, n10793, n10794, 
      n10795, n10797, n10798, n10800, n10801, n10804, n10807, n10808, n10809, 
      n10810, n10811, n10812, n10813, n10815, n10816, n10817, n10818, n10819, 
      n10820, n10821, n10823, n10826, n10827, n10828, n10829, n10830, n10832, 
      n10833, n10834, n10838, n10839, n10840, n10841, n10842, n10843, n10844, 
      n10845, n10847, n10849, n10850, n10851, n10852, n10853, n10854, n10855, 
      n10856, n10858, n10862, n10863, n10864, n10865, n10866, n10868, n10869, 
      n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10878, n10880, 
      n10881, n10882, n10883, n10884, n10885, n10887, n10889, n10890, n10891, 
      n10893, n10894, n10895, n10897, n10898, n10901, n10903, n10904, n10905, 
      n10906, n10907, n10908, n10911, n10912, n10913, n10914, n10917, n10918, 
      n10919, n10920, n10921, n10922, n10923, n10924, n10926, n10927, n10928, 
      n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, 
      n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, 
      n10947, n10948, n10950, n10951, n10952, n10953, n10954, n10956, n10957, 
      n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, 
      n10967, n10968, n10970, n10971, n10972, n10974, n10975, n10976, n10977, 
      n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, 
      n10988, n10989, n10990, n10992, n10993, n10995, n10996, n10997, n10998, 
      n10999, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11010, 
      n11011, n11012, n11013, n11014, n11015, n11017, n11018, n11021, n11022, 
      n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, 
      n11032, n11033, n11034, n11035, n11037, n11038, n11039, n11040, n11041, 
      n11042, n11044, n11046, n11047, n11048, n11049, n11051, n11052, n11053, 
      n11054, n11058, n11059, n11061, n11062, n11063, n11067, n11068, n11069, 
      n11070, n11071, n11072, n11073, n11074, n11076, n11077, n11078, n11079, 
      n11080, n11081, n11082, n11084, n11085, n11087, n11088, n11089, n11090, 
      n11092, n11093, n11094, n11095, n11097, n11098, n11100, n11102, n11103, 
      n11105, n11107, n11108, n11110, n11111, n11112, n11113, n11114, n11117, 
      n11118, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11129, 
      n11130, n11132, n11134, n11136, n11137, n11138, n11140, n11141, n11142, 
      n11143, n11144, n11147, n11148, n11150, n11151, n11152, n11153, n11154, 
      n11155, n11156, n11157, n11160, n11161, n11163, n11164, n11165, n11166, 
      n11167, n11168, n11170, n11171, n11174, n11175, n11176, n11177, n11178, 
      n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, 
      n11189, n11190, n11191, n11193, n11194, n11195, n11196, n11197, n11198, 
      n11200, n11201, n11203, n11204, n11205, n11206, n11207, n11209, n11210, 
      n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11219, n11220, 
      n11222, n11223, n11224, n11225, n11226, n11228, n11229, n11230, n11231, 
      n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, 
      n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, 
      n11251, n11253, n11255, n11256, n11257, n11259, n11261, n11262, n11263, 
      n11264, n11267, n11270, n11275, n11276, n11277, n11278, n11279, n11280, 
      n11281, n11282, n11283, n11284, n11286, n11287, n11288, n11289, n11290, 
      n11291, n11292, n11293, n11294, n11295, n11296, n11299, n11300, n11303, 
      n11306, n11307, n11309, n11312, n11313, n11314, n11315, n11316, n11317, 
      n11318, n11319, n11320, n11321, n11322, n11323, n11325, n11326, n11327, 
      n11328, n11329, n11330, n11331, n11334, n11336, n11337, n11339, n11341, 
      n11342, n11343, n11344, n11345, n11353, n11354, n11355, n11356, n11359, 
      n11360, n11361, n11363, n11364, n11366, n11369, n11370, n11371, n11372, 
      n11373, n11374, n11376, n11377, n11378, n11379, n11380, n11382, n11383, 
      n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11395, 
      n11396, n11397, n11398, n11400, n11401, n11402, n11403, n11404, n11405, 
      n11407, n11408, n11409, n11410, n11411, n11413, n11414, n11415, n11416, 
      n11417, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, 
      n11427, n11429, n11430, n11431, n11432, n11434, n11435, n11436, n11438, 
      n11439, n11440, n11442, n11443, n11444, n11445, n11447, n11450, n11452, 
      n11453, n11454, n11456, n11457, n11458, n11459, n11460, n11461, n11462, 
      n11463, n11464, n11465, n11466, n11467, n11468, n11470, n11471, n11472, 
      n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, 
      n11483, n11485, n11486, n11487, n11488, n11490, n11491, n11492, n11493, 
      n11494, n11495, n11497, n11498, n11499, n11501, n11502, n11503, n11504, 
      n11505, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, 
      n11519, n11521, n11522, n11524, n11525, n11528, n11532, n11533, n11535, 
      n11539, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, 
      n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, 
      n11558, n11559, n11560, n11562, n11564, n11565, n11566, n11567, n11568, 
      n11569, n11571, n11572, n11574, n11575, n11576, n11577, n11578, n11579, 
      n11580, n11581, n11583, n11587, n11589, n11590, n11591, n11592, n11593, 
      n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, 
      n11605, n11606, n11607, n11609, n11610, n11611, n11612, n11613, n11614, 
      n11616, n11617, n11618, n11619, n11622, n11623, n11624, n11626, n11627, 
      n11628, n11629, n11630, n11631, n11632, n11633, n11636, n11637, n11640, 
      n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11651, 
      n11652, n11653, n11655, n11656, n11658, n11660, n11661, n11663, n11664, 
      n11667, n11668, n11670, n11671, n11672, n11674, n11675, n11676, n11677, 
      n11678, n11679, n11680, n11681, n11682, n11684, n11685, n11687, n11689, 
      n11691, n11692, n11693, n11694, n11696, n11698, n11699, n11701, n11702, 
      n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11711, n11712, 
      n11714, n11715, n11716, n11718, n11719, n11721, n11722, n11723, n11726, 
      n11728, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, 
      n11739, n11741, n11743, n11744, n11746, n11747, n11748, n11750, n11751, 
      n11752, n11753, n11755, n11756, n11757, n11759, n11760, n11761, n11762, 
      n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, 
      n11773, n11775, n11776, n11777, n11778, n11780, n11781, n11782, n11783, 
      n11785, n11786, n11787, n11789, n11792, n11793, n11794, n11795, n11796, 
      n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11805, n11806, 
      n11808, n11809, n11811, n11812, n11813, n11815, n11816, n11817, n11818, 
      n11819, n11820, n11821, n11822, n11824, n11826, n11828, n11829, n11830, 
      n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, 
      n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11852, 
      n11854, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11865, 
      n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, 
      n11875, n11876, n11877, n11878, n11880, n11885, n11886, n11887, n11890, 
      n11891, n11892, n11893, n11894, n11896, n11897, n11898, n11899, n11900, 
      n11901, n11902, n11904, n11905, n11906, n11907, n11908, n11909, n11910, 
      n11911, n11912, n11913, n11917, n11918, n11919, n11920, n11923, n11924, 
      n11925, n11926, n11927, n11932, n11933, n11934, n11935, n11936, n11937, 
      n11938, n11939, n11940, n11943, n11944, n11945, n11946, n11947, n11950, 
      n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, 
      n11961, n11962, n11964, n11965, n11966, n11967, n11968, n11969, n11970, 
      n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11980, n11981, 
      n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, 
      n11991, n11992, n11994, n11995, n11996, n11997, n11999, n12001, n12002, 
      n12003, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, 
      n12014, n12015, n12016, n12018, n12019, n12020, n12021, n12022, n12023, 
      n12024, n12025, n12026, n12027, n12030, n12031, n12033, n12034, n12035, 
      n12036, n12037, n12039, n12040, n12041, n12042, n12044, n12045, n12046, 
      n12047, n12048, n12049, n12050, n12053, n12054, n12055, n12056, n12057, 
      n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12066, n12067, 
      n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12077, n12078, 
      n12079, n12080, n12081, n12082, n12083, n12085, n12086, n12087, n12089, 
      n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, 
      n12099, n12100, n12102, n12104, n12105, n12106, n12107, n12108, n12109, 
      n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12120, 
      n12122, n12124, n12125, n12126, n12128, n12129, n12130, n12131, n12132, 
      n12135, n12136, n12138, n12139, n12140, n12142, n12143, n12144, n12145, 
      n12146, n12147, n12149, n12151, n12152, n12153, n12154, n12156, n12157, 
      n12159, n12160, n12162, n12164, n12166, n12169, n12170, n12171, n12172, 
      n12175, n12176, n12177, n12179, n12180, n12181, n12182, n12184, n12185, 
      n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, 
      n12195, n12196, n12197, n12200, n12202, n12203, n12204, n12205, n12206, 
      n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12217, n12218, 
      n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, 
      n12228, n12230, n12233, n12234, n12235, n12236, n12239, n12241, n12242, 
      n12244, n12245, n12246, n12247, n12249, n12250, n12251, n12252, n12253, 
      n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12263, 
      n12264, n12265, n12266, n12267, n12270, n12271, n12272, n12274, n12275, 
      n12276, n12277, n12278, n12279, n12281, n12282, n12283, n12285, n12286, 
      n12287, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, 
      n12300, n12302, n12304, n12305, n12306, n12307, n12308, n12309, n12310, 
      n12311, n12312, n12314, n12315, n12316, n12317, n12318, n12320, n12321, 
      n12322, n12323, n12324, n12325, n12327, n12328, n12329, n12331, n12334, 
      n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, 
      n12344, n12346, n12348, n12351, n12352, n12353, n12354, n12355, n12357, 
      n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, 
      n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, 
      n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12389, n12391, 
      n12393, n12394, n12395, n12396, n12397, n12399, n12401, n12402, n12403, 
      n12405, n12406, n12407, n12410, n12411, n12413, n12414, n12416, n12417, 
      n12419, n12421, n12423, n12424, n12425, n12426, n12428, n12429, n12430, 
      n12431, n12432, n12433, n12434, n12437, n12438, n12439, n12440, n12441, 
      n12443, n12444, n12445, n12446, n12449, n12450, n12451, n12452, n12453, 
      n12454, n12455, n12457, n12458, n12459, n12463, n12464, n12465, n12466, 
      n12467, n12468, n12470, n12472, n12473, n12474, n12475, n12476, n12477, 
      n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, 
      n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, 
      n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12506, n12507, 
      n12508, n12509, n12510, n12512, n12515, n12516, n12517, n12518, n12519, 
      n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, 
      n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12540, 
      n12542, n12545, n12546, n12548, n12549, n12551, n12553, n12554, n12555, 
      n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12569, 
      n12570, n12571, n12572, n12573, n12574, n12576, n12577, n12579, n12580, 
      n12581, n12583, n12584, n12585, n12586, n12588, n12589, n12590, n12593, 
      n12594, n12595, n12596, n12598, n12599, n12600, n12601, n12602, n12603, 
      n12604, n12605, n12607, n12608, n12610, n12611, n12612, n12613, n12614, 
      n12615, n12617, n12618, n12619, n12620, n12621, n12623, n12625, n12626, 
      n12627, n12628, n12629, n12631, n12632, n12633, n12634, n12635, n12637, 
      n12638, n12639, n12641, n12643, n12644, n12645, n12646, n12647, n12648, 
      n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12658, 
      n12659, n12661, n12664, n12665, n12666, n12667, n12668, n12669, n12670, 
      n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, 
      n12681, n12682, n12684, n12686, n12689, n12690, n12691, n12692, n12693, 
      n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, 
      n12703, n12704, n12706, n12707, n12708, n12709, n12711, n12712, n12713, 
      n12714, n12715, n12717, n12718, n12719, n12720, n12721, n12722, n12723, 
      n12724, n12725, n12726, n12728, n12729, n12731, n12732, n12733, n12734, 
      n12735, n12736, n12738, n12739, n12742, n12746, n12748, n12749, n12750, 
      n12751, n12752, n12754, n12755, n12757, n12759, n12760, n12761, n12763, 
      n12765, n12766, n12767, n12769, n12771, n12772, n12773, n12775, n12776, 
      n12777, n12778, n12779, n12781, n12783, n12784, n12785, n12786, n12788, 
      n12789, n12790, n12791, n12795, n12797, n12800, n12801, n12802, n12803, 
      n12806, n12807, n12809, n12810, n12812, n12813, n12815, n12816, n12817, 
      n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, 
      n12829, n12830, n12831, n12832, n12834, n12836, n12837, n12839, n12840, 
      n12843, n12845, n12846, n12847, n12849, n12850, n12851, n12852, n12853, 
      n12854, n12855, n12857, n12860, n12862, n12863, n12866, n12870, n12871, 
      n12872, n12874, n12875, n12876, n12879, n12881, n12882, n12884, n12885, 
      n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, 
      n12895, n12896, n12897, n12899, n12900, n12902, n12903, n12904, n12906, 
      n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12915, n12916, 
      n12918, n12919, n12922, n12925, n12926, n12928, n12930, n12931, n12932, 
      n12933, n12934, n12935, n12937, n12938, n12939, n12941, n12942, n12943, 
      n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, 
      n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, 
      n12962, n12964, n12967, n12969, n12973, n12974, n12976, n12977, n12978, 
      n12979, n12980, n12981, n12982, n12983, n12986, n12989, n12991, n12992, 
      n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13005, 
      n13007, n13008, n13009, n13011, n13012, n13013, n13015, n13018, n13019, 
      n13020, n13021, n13022, n13023, n13025, n13028, n13030, n13031, n13032, 
      n13033, n13034, n13035, n13036, n13037, n13039, n13040, n13042, n13043, 
      n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, 
      n13054, n13055, n13056, n13057, n13059, n13061, n13062, n13063, n13064, 
      n13066, n13067, n13069, n13070, n13071, n13072, n13073, n13074, n13075, 
      n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13084, n13085, 
      n13086, n13088, n13089, n13090, n13091, n13092, n13093, n13095, n13096, 
      n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, 
      n13106, n13107, n13109, n13110, n13112, n13113, n13114, n13115, n13116, 
      n13117, n13118, n13119, n13121, n13122, n13123, n13125, n13126, n13127, 
      n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13136, n13137, 
      n13138, n13140, n13142, n13145, n13146, n13147, n13148, n13150, n13151, 
      n13152, n13153, n13154, n13155, n13156, n13157, n13159, n13160, n13161, 
      n13164, n13165, n13167, n13169, n13170, n13171, n13172, n13174, n13178, 
      n13179, n13180, n13181, n13183, n13184, n13185, n13186, n13187, n13188, 
      n13189, n13190, n13191, n13192, n13194, n13195, n13196, n13197, n13198, 
      n13200, n13201, n13202, n13203, n13205, n13207, n13208, n13209, n13210, 
      n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, 
      n13220, n13223, n13224, n13225, n13226, n13228, n13229, n13230, n13232, 
      n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13242, n13244, 
      n13245, n13246, n13247, n13248, n13250, n13252, n13253, n13255, n13256, 
      n13259, n13261, n13263, n13264, n13265, n13267, n13268, n13269, n13270, 
      n13271, n13272, n13274, n13275, n13276, n13278, n13280, n13281, n13282, 
      n13283, n13284, n13285, n13287, n13288, n13289, n13291, n13293, n13294, 
      n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13303, n13305, 
      n13306, n13307, n13308, n13309, n13310, n13311, n13314, n13315, n13319, 
      n13320, n13321, n13325, n13326, n13327, n13329, n13330, n13332, n13333, 
      n13334, n13335, n13337, n13338, n13339, n13340, n13341, n13342, n13343, 
      n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, 
      n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, 
      n13362, n13363, n13364, n13365, n13369, n13370, n13371, n13372, n13373, 
      n13374, n13375, n13376, n13378, n13379, n13380, n13382, n13383, n13385, 
      n13386, n13387, n13388, n13389, n13390, n13391, n13395, n13396, n13398, 
      n13399, n13400, n13401, n13402, n13403, n13404, n13406, n13407, n13410, 
      n13411, n13412, n13415, n13416, n13417, n13418, n13420, n13421, n13422, 
      n13423, n13424, n13425, n13426, n13428, n13429, n13430, n13431, n13432, 
      n13433, n13434, n13435, n13436, n13437, n13438, n13440, n13443, n13444, 
      n13445, n13446, n13447, n13448, n13449, n13450, n13453, n13454, n13455, 
      n13457, n13458, n13459, n13460, n13461, n13463, n13464, n13466, n13467, 
      n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, 
      n13477, n13478, n13480, n13481, n13482, n13483, n13485, n13486, n13488, 
      n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, 
      n13498, n13499, n13502, n13503, n13504, n13505, n13506, n13507, n13508, 
      n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13517, n13518, 
      n13519, n13522, n13524, n13525, n13526, n13528, n13530, n13532, n13533, 
      n13534, n13535, n13536, n13537, n13538, n13539, n13541, n13545, n13546, 
      n13547, n13548, n13549, n13550, n13551, n13553, n13554, n13557, n13560, 
      n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13570, 
      n13571, n13572, n13573, n13574, n13577, n13578, n13579, n13580, n13581, 
      n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, 
      n13592, n13593, n13594, n13595, n13596, n13597, n13599, n13600, n13601, 
      n13602, n13604, n13605, n13606, n13607, n13608, n13610, n13612, n13613, 
      n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, 
      n13623, n13624, n13625, n13628, n13629, n13631, n13632, n13633, n13636, 
      n13637, n13638, n13642, n13643, n13644, n13645, n13646, n13647, n13648, 
      n13649, n13650, n13651, n13652, n13655, n13656, n13657, n13658, n13659, 
      n13660, n13661, n13662, n13663, n13665, n13666, n13669, n13671, n13673, 
      n13674, n13676, n13677, n13678, n13679, n13680, n13682, n13684, n13685, 
      n13686, n13687, n13688, n13690, n13693, n13694, n13695, n13697, n13698, 
      n13699, n13700, n13701, n13702, n13704, n13705, n13709, n13710, n13711, 
      n13712, n13714, n13715, n13716, n13717, n13718, n13719, n13721, n13722, 
      n13723, n13726, n13727, n13729, n13730, n13731, n13732, n13734, n13735, 
      n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13746, 
      n13747, n13748, n13749, n13750, n13751, n13752, n13754, n13755, n13756, 
      n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, 
      n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, 
      n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, 
      n13784, n13785, n13786, n13787, n13788, n13790, n13791, n13793, n13794, 
      n13796, n13797, n13798, n13799, n13802, n13803, n13805, n13806, n13807, 
      n13808, n13809, n13810, n13811, n13812, n13813, n13815, n13816, n13818, 
      n13819, n13821, n13822, n13824, n13825, n13826, n13829, n13830, n13831, 
      n13832, n13833, n13834, n13835, n13837, n13838, n13840, n13841, n13842, 
      n13843, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, 
      n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, 
      n13862, n13863, n13864, n13865, n13866, n13868, n13869, n13870, n13872, 
      n13873, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, 
      n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13894, 
      n13895, n13896, n13897, n13900, n13902, n13903, n13904, n13905, n13906, 
      n13908, n13909, n13911, n13912, n13914, n13915, n13916, n13917, n13918, 
      n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, 
      n13928, n13929, n13930, n13932, n13933, n13934, n13936, n13937, n13938, 
      n13939, n13940, n13942, n13943, n13944, n13945, n13946, n13948, n13949, 
      n13950, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, 
      n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, 
      n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, 
      n13981, n13982, n13983, n13984, n13986, n13987, n13988, n13989, n13990, 
      n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, 
      n14001, n14002, n14006, n14007, n14008, n14009, n14010, n14011, n14012, 
      n14014, n14015, n14016, n14017, n14019, n14020, n14021, n14022, n14023, 
      n14024, n14025, n14026, n14027, n14028, n14032, n14033, n14034, n14035, 
      n14036, n14037, n14038, n14039, n14041, n14042, n14043, n14044, n14046, 
      n14047, n14048, n14052, n14053, n14054, n14055, n14056, n14058, n14059, 
      n14060, n14061, n14062, n14063, n14065, n14066, n14067, n14068, n14069, 
      n14070, n14071, n14073, n14075, n14077, n14078, n14079, n14080, n14082, 
      n14085, n14088, n14089, n14090, n14091, n14093, n14094, n14095, n14096, 
      n14097, n14098, n14099, n14100, n14102, n14103, n14104, n14105, n14106, 
      n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14116, 
      n14117, n14119, n14120, n14121, n14122, n14123, n14126, n14127, n14128, 
      n14129, n14132, n14134, n14136, n14137, n14138, n14139, n14140, n14141, 
      n14142, n14143, n14144, n14145, n14146, n14148, n14150, n14151, n14152, 
      n14153, n14154, n14156, n14157, n14162, n14163, n14165, n14166, n14167, 
      n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14176, n14177, 
      n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14187, 
      n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, 
      n14197, n14198, n14201, n14202, n14203, n14204, n14206, n14207, n14208, 
      n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, 
      n14219, n14220, n14221, n14222, n14224, n14225, n14227, n14228, n14229, 
      n14230, n14234, n14235, n14237, n14238, n14239, n14240, n14241, n14242, 
      n14243, n14244, n14245, n14246, n14248, n14250, n14252, n14253, n14254, 
      n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, 
      n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, 
      n14273, n14274, n14275, n14277, n14278, n14279, n14281, n14282, n14283, 
      n14284, n14285, n14287, n14288, n14289, n14291, n14292, n14293, n14294, 
      n14300, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, 
      n14310, n14311, n14312, n14313, n14314, n14317, n14318, n14319, n14320, 
      n14321, n14322, n14324, n14325, n14326, n14328, n14332, n14334, n14335, 
      n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, 
      n14345, n14346, n14347, n14348, n14350, n14351, n14352, n14353, n14354, 
      n14356, n14357, n14358, n14360, n14361, n14362, n14364, n14367, n14368, 
      n14369, n14370, n14371, n14372, n14375, n14376, n14377, n14378, n14382, 
      n14383, n14384, n14385, n14386, n14390, n14391, n14392, n14393, n14395, 
      n14396, n14397, n14398, n14399, n14401, n14402, n14403, n14404, n14405, 
      n14406, n14407, n14408, n14409, n14410, n14411, n14414, n14415, n14416, 
      n14417, n14418, n14419, n14420, n14421, n14423, n14424, n14425, n14426, 
      n14427, n14428, n14429, n14430, n14432, n14433, n14434, n14435, n14436, 
      n14437, n14438, n14440, n14441, n14442, n14443, n14445, n14446, n14447, 
      n14448, n14450, n14451, n14452, n14453, n14455, n14456, n14457, n14458, 
      n14459, n14460, n14461, n14463, n14465, n14466, n14467, n14468, n14469, 
      n14472, n14473, n14474, n14478, n14479, n14480, n14481, n14483, n14484, 
      n14485, n14487, n14488, n14489, n14491, n14492, n14494, n14495, n14496, 
      n14497, n14498, n14500, n14501, n14502, n14503, n14504, n14505, n14506, 
      n14507, n14508, n14509, n14510, n14512, n14513, n14514, n14515, n14516, 
      n14518, n14519, n14520, n14521, n14522, n14525, n14526, n14528, n14529, 
      n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, 
      n14539, n14540, n14542, n14543, n14544, n14545, n14546, n14548, n14549, 
      n14550, n14551, n14552, n14554, n14555, n14556, n14557, n14558, n14559, 
      n14560, n14561, n14562, n14564, n14565, n14566, n14567, n14568, n14569, 
      n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14578, n14579, 
      n14580, n14581, n14582, n14583, n14584, n14586, n14587, n14588, n14589, 
      n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, 
      n14599, n14600, n14601, n14602, n14604, n14605, n14606, n14607, n14608, 
      n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, 
      n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14626, n14627, 
      n14628, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, 
      n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, 
      n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, 
      n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, 
      n14665, n14666, n14668, n14669, n14670, n14671, n14672, n14673, n14675, 
      n14676, n14677, n14678, n14679, n14681, n14682, n14683, n14684, n14685, 
      n14686, n14687, n14688, n14689, n14690, n14693, n14694, n14695, n14697, 
      n14698, n14699, n14700, n14701, n14702, n14704, n14705, n14706, n14707, 
      n14708, n14709, n14710, n14712, n14715, n14716, n14717, n14718, n14719, 
      n14720, n14721, n14723, n14724, n14726, n14728, n14732, n14733, n14734, 
      n14735, n14737, n14739, n14740, n14741, n14743, n14744, n14745, n14746, 
      n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14757, 
      n14758, n14759, n14761, n14762, n14763, n14764, n14765, n14766, n14767, 
      n14771, n14772, n14775, n14776, n14777, n14778, n14779, n14780, n14781, 
      n14782, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, 
      n14792, n14793, n14795, n14796, n14797, n14800, n14801, n14802, n14803, 
      n14804, n14806, n14808, n14810, n14811, n14813, n14814, n14815, n14816, 
      n14819, n14820, n14821, n14823, n14826, n14828, n14829, n14830, n14831, 
      n14832, n14833, n14835, n14836, n14837, n14838, n14840, n14841, n14842, 
      n14843, n14844, n14845, n14848, n14850, n14851, n14852, n14853, n14854, 
      n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, 
      n14864, n14865, n14866, n14868, n14870, n14872, n14873, n14876, n14878, 
      n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, 
      n14888, n14889, n14891, n14892, n14893, n14894, n14895, n14896, n14900, 
      n14901, n14902, n14903, n14904, n14906, n14907, n14908, n14909, n14910, 
      n14911, n14912, n14914, n14915, n14916, n14917, n14920, n14921, n14922, 
      n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14931, n14932, 
      n14933, n14934, n14939, n14940, n14941, n14942, n14943, n14944, n14945, 
      n14947, n14948, n14950, n14951, n14952, n14954, n14955, n14956, n14957, 
      n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, 
      n14968, n14969, n14971, n14972, n14973, n14974, n14975, n14976, n14977, 
      n14978, n14979, n14980, n14981, n14982, n14984, n14986, n14989, n14990, 
      n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, 
      n15000, n15001, n15002, n15003, n15004, n15005, n15007, n15008, n15009, 
      n15010, n15012, n15013, n15015, n15016, n15017, n15018, n15019, n15021, 
      n15022, n15023, n15025, n15026, n15027, n15028, n15029, n15030, n15031, 
      n15034, n15036, n15037, n15038, n15039, n15040, n15041, n15043, n15044, 
      n15046, n15048, n15049, n15052, n15053, n15054, n15055, n15056, n15057, 
      n15058, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, 
      n15069, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, 
      n15081, n15084, n15085, n15088, n15089, n15090, n15091, n15093, n15094, 
      n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, 
      n15105, n15106, n15107, n15108, n15109, n15111, n15112, n15113, n15114, 
      n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15124, 
      n15125, n15126, n15128, n15129, n15130, n15131, n15132, n15133, n15134, 
      n15135, n15136, n15137, n15138, n15142, n15143, n15144, n15145, n15146, 
      n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15155, n15156, 
      n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15167, n15168, 
      n15169, n15172, n15173, n15174, n15175, n15177, n15178, n15179, n15180, 
      n15181, n15182, n15183, n15186, n15187, n15188, n15189, n15190, n15192, 
      n15193, n15194, n15195, n15197, n15198, n15199, n15201, n15202, n15203, 
      n15205, n15207, n15208, n15209, n15210, n15211, n15213, n15214, n15215, 
      n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, 
      n15226, n15227, n15228, n15230, n15231, n15234, n15235, n15236, n15237, 
      n15239, n15241, n15242, n15243, n15244, n15246, n15249, n15250, n15253, 
      n15255, n15256, n15258, n15260, n15261, n15262, n15265, n15266, n15268, 
      n15269, n15270, n15271, n15272, n15273, n15276, n15277, n15278, n15279, 
      n15280, n15281, n15282, n15284, n15285, n15286, n15287, n15288, n15290, 
      n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, 
      n15300, n15301, n15302, n15303, n15305, n15307, n15308, n15309, n15310, 
      n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, 
      n15320, n15321, n15322, n15324, n15325, n15326, n15329, n15330, n15331, 
      n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, 
      n15341, n15342, n15343, n15344, n15345, n15347, n15348, n15349, n15351, 
      n15352, n15353, n15354, n15356, n15358, n15359, n15360, n15361, n15362, 
      n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15372, n15373, 
      n15374, n15375, n15376, n15378, n15379, n15380, n15381, n15382, n15383, 
      n15384, n15385, n15386, n15387, n15390, n15391, n15392, n15393, n15394, 
      n15395, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15405, 
      n15406, n15407, n15408, n15411, n15412, n15413, n15414, n15415, n15416, 
      n15418, n15419, n15420, n15421, n15423, n15424, n15425, n15426, n15427, 
      n15428, n15429, n15430, n15431, n15432, n15434, n15435, n15436, n15437, 
      n15438, n15439, n15440, n15441, n15442, n15443, n15447, n15448, n15449, 
      n15450, n15451, n15453, n15454, n15455, n15456, n15457, n15458, n15459, 
      n15460, n15461, n15462, n15463, n15466, n15468, n15469, n15470, n15471, 
      n15472, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, 
      n15482, n15483, n15485, n15486, n15487, n15488, n15489, n15490, n15491, 
      n15492, n15493, n15494, n15496, n15497, n15498, n15499, n15500, n15501, 
      n15502, n15503, n15504, n15506, n15507, n15509, n15510, n15511, n15512, 
      n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, 
      n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, 
      n15532, n15533, n15534, n15536, n15537, n15538, n15539, n15540, n15542, 
      n15544, n15545, n15546, n15547, n15548, n15550, n15551, n15552, n15553, 
      n15554, n15556, n15557, n15558, n15559, n15560, n15562, n15563, n15564, 
      n15565, n15568, n15570, n15571, n15573, n15575, n15576, n15577, n15578, 
      n15579, n15580, n15582, n15583, n15584, n15586, n15589, n15592, n15593, 
      n15594, n15596, n15597, n15598, n15599, n15600, n15603, n15604, n15606, 
      n15607, n15609, n15610, n15611, n15613, n15614, n15615, n15616, n15618, 
      n15619, n15620, n15621, n15622, n15623, n15624, n15627, n15631, n15632, 
      n15633, n15634, n15636, n15637, n15638, n15639, n15640, n15641, n15642, 
      n15643, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, 
      n15653, n15655, n15656, n15657, n15658, n15660, n15661, n15662, n15663, 
      n15664, n15667, n15669, n15670, n15673, n15674, n15675, n15676, n15677, 
      n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, 
      n15688, n15689, n15690, n15691, n15693, n15694, n15696, n15697, n15698, 
      n15699, n15701, n15702, n15703, n15704, n15705, n15706, n15708, n15709, 
      n15710, n15711, n15712, n15713, n15714, n15717, n15718, n15719, n15720, 
      n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, 
      n15730, n15731, n15732, n15733, n15734, n15735, n15737, n15738, n15739, 
      n15740, n15742, n15743, n15744, n15748, n15751, n15752, n15754, n15756, 
      n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, 
      n15766, n15767, n15768, n15769, n15770, n15772, n15773, n15774, n15775, 
      n15776, n15777, n15778, n15779, n15781, n15782, n15783, n15784, n15786, 
      n15787, n15788, n15790, n15793, n15794, n15795, n15796, n15797, n15798, 
      n15799, n15800, n15801, n15803, n15804, n15805, n15806, n15807, n15808, 
      n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, 
      n15819, n15820, n15821, n15822, n15824, n15825, n15826, n15827, n15828, 
      n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, 
      n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15847, 
      n15848, n15850, n15851, n15852, n15853, n15855, n15856, n15857, n15858, 
      n15859, n15860, n15861, n15862, n15864, n15865, n15866, n15867, n15868, 
      n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15877, n15878, 
      n15879, n15880, n15881, n15882, n15884, n15885, n15886, n15887, n15888, 
      n15889, n15890, n15891, n15892, n15894, n15895, n15897, n15898, n15900, 
      n15901, n15903, n15904, n15905, n15906, n15908, n15909, n15912, n15913, 
      n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, 
      n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, 
      n15932, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, 
      n15942, n15943, n15945, n15946, n15947, n15949, n15950, n15951, n15952, 
      n15953, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, 
      n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, 
      n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, 
      n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, 
      n15991, n15992, n15994, n15995, n15996, n15997, n15998, n15999, n16001, 
      n16002, n16003, n16005, n16006, n16007, n16008, n16009, n16010, n16011, 
      n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, 
      n16021, n16022, n16023, n16025, n16026, n16027, n16028, n16029, n16030, 
      n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16041, 
      n16042, n16043, n16044, n16046, n16047, n16048, n16049, n16050, n16051, 
      n16055, n16056, n16057, n16058, n16059, n16062, n16063, n16064, n16065, 
      n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, 
      n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, 
      n16085, n16086, n16088, n16089, n16090, n16091, n16092, n16093, n16094, 
      n16095, n16096, n16097, n16098, n16100, n16102, n16103, n16104, n16105, 
      n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, 
      n16115, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, 
      n16125, n16126, n16127, n16128, n16130, n16131, n16132, n16133, n16134, 
      n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, 
      n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, 
      n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, 
      n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, 
      n16171, n16172, n16175, n16176, n16177, n16178, n16179, n16181, n16182, 
      n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, 
      n16193, n16194, n16195, n16196, n16197, n16198, n16200, n16201, n16202, 
      n16203, n16204, n16206, n16207, n16209, n16212, n16213, n16214, n16215, 
      n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, 
      n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, 
      n16234, n16235, n16236, n16237, n16239, n16240, n16241, n16242, n16244, 
      n16245, n16246, n16247, n16249, n16250, n16251, n16252, n16253, n16254, 
      n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, 
      n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, 
      n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16282, 
      n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, 
      n16292, n16293, n16295, n16298, n16299, n16300, n16301, n16302, n16303, 
      n16304, n16305, n16306, n16307, n16308, n16309, n16311, n16312, n16313, 
      n16314, n16315, n16316, n16317, n16318, n16320, n16321, n16323, n16324, 
      n16325, n16326, n16329, n16330, n16331, n16332, n16333, n16334, n16335, 
      n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, 
      n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, 
      n16354, n16355, n16356, n16358, n16359, n16360, n16361, n16362, n16363, 
      n16366, n16367, n16368, n16370, n16371, n16372, n16374, n16375, n16376, 
      n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, 
      n16386, n16387, n16389, n16391, n16392, n16393, n16394, n16397, n16398, 
      n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, 
      n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, 
      n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16426, 
      n16428, n16429, n16430, n16432, n16433, n16434, n16435, n16437, n16438, 
      n16439, n16440, n16441, n16443, n16444, n16445, n16446, n16447, n16448, 
      n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, 
      n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16466, n16467, 
      n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, 
      n16478, n16481, n16483, n16484, n16485, n16486, n16488, n16490, n16491, 
      n16493, n16494, n16496, n16497, n16498, n16500, n16501, n16502, n16503, 
      n16505, n16507, n16508, n16510, n16511, n16512, n16513, n16514, n16515, 
      n16516, n16517, n16518, n16519, n16520, n16521, n16523, n16524, n16525, 
      n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, 
      n16535, n16537, n16538, n16540, n16542, n16544, n16545, n16546, n16547, 
      n16548, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, 
      n16558, n16559, n16561, n16562, n16563, n16564, n16565, n16566, n16567, 
      n16568, n16569, n16571, n16572, n16573, n16574, n16575, n16576, n16577, 
      n16578, n16579, n16580, n16583, n16584, n16585, n16587, n16588, n16589, 
      n16590, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, 
      n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, 
      n16611, n16612, n16614, n16615, n16616, n16617, n16618, n16619, n16620, 
      n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16629, n16630, 
      n16632, n16633, n16634, n16635, n16636, n16638, n16639, n16640, n16642, 
      n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16651, n16652, 
      n16653, n16654, n16656, n16657, n16658, n16660, n16661, n16662, n16663, 
      n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, 
      n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16684, n16685, 
      n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, 
      n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16704, 
      n16705, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, 
      n16715, n16716, n16718, n16719, n16720, n16722, n16723, n16724, n16725, 
      n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, 
      n16735, n16736, n16737, n16739, n16740, n16741, n16742, n16743, n16744, 
      n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, 
      n16754, n16755, n16756, n16757, n16759, n16760, n16762, n16763, n16764, 
      n16765, n16767, n16768, n16769, n16770, n16771, n16773, n16774, n16778, 
      n16779, n16780, n16781, n16783, n16784, n16785, n16786, n16787, n16788, 
      n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, 
      n16798, n16799, n16800, n16801, n16803, n16804, n16805, n16806, n16807, 
      n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, 
      n16817, n16818, n16819, n16820, n16822, n16823, n16825, n16826, n16828, 
      n16829, n16830, n16832, n16834, n16835, n16836, n16838, n16839, n16840, 
      n16841, n16842, n16845, n16846, n16847, n16848, n16849, n16850, n16851, 
      n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, 
      n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, 
      n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, 
      n16879, n16880, n16881, n16883, n16884, n16885, n16886, n16887, n16889, 
      n16890, n16893, n16894, n16895, n16897, n16898, n16899, n16900, n16901, 
      n16902, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, 
      n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, 
      n16922, n16924, n16928, n16929, n16930, n16931, n16932, n16933, n16934, 
      n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, 
      n16944, n16945, n16946, n16947, n16948, n16950, n16951, n16955, n16957, 
      n16958, n16959, n16960, n16961, n16962, n16964, n16965, n16966, n16967, 
      n16968, n16969, n16970, n16971, n16972, n16973, n16975, n16976, n16977, 
      n16980, n16981, n16982, n16985, n16987, n16988, n16989, n16990, n16991, 
      n16992, n16993, n16994, n16995, n16996, n16998, n16999, n17000, n17001, 
      n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, 
      n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17021, 
      n17022, n17023, n17024, n17025, n17026, n17028, n17029, n17030, n17031, 
      n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, 
      n17041, n17042, n17044, n17045, n17046, n17047, n17049, n17051, n17053, 
      n17054, n17055, n17056, n17057, n17058, n17059, n17061, n17062, n17063, 
      n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, 
      n17073, n17074, n17075, n17076, n17077, n17078, n17080, n17081, n17082, 
      n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, 
      n17092, n17094, n17095, n17096, n17097, n17098, n17100, n17101, n17102, 
      n17103, n17104, n17105, n17106, n17108, n17109, n17110, n17112, n17113, 
      n17114, n17115, n17116, n17117, n17119, n17120, n17121, n17122, n17123, 
      n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, 
      n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, 
      n17142, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, 
      n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, 
      n17164, n17166, n17168, n17169, n17172, n17173, n17174, n17175, n17176, 
      n17177, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17187, 
      n17188, n17191, n17192, n17193, n17195, n17196, n17197, n17198, n17199, 
      n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17208, n17209, 
      n17210, n17211, n17213, n17214, n17216, n17217, n17218, n17219, n17220, 
      n17221, n17222, n17223, n17224, n17226, n17227, n17228, n17229, n17230, 
      n17231, n17232, n17234, n17235, n17236, n17238, n17240, n17241, n17242, 
      n17243, n17244, n17246, n17247, n17248, n17249, n17250, n17251, n17252, 
      n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17261, n17262, 
      n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, 
      n17277, n17278, n17279, n17280, n17281, n17286, n17287, n17288, n17290, 
      n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17300, 
      n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, 
      n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, 
      n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17328, 
      n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, 
      n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, 
      n17350, n17351, n17352, n17353, n17354, n17355, n17357, n17358, n17359, 
      n17360, n17362, n17363, n17364, n17365, n17366, n17367, n17369, n17370, 
      n17372, n17374, n17376, n17379, n17380, n17381, n17383, n17384, n17385, 
      n17386, n17388, n17390, n17391, n17393, n17396, n17397, n17398, n17399, 
      n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, 
      n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, 
      n17418, n17419, n17421, n17422, n17424, n17426, n17427, n17429, n17431, 
      n17432, n17433, n17435, n17436, n17437, n17440, n17441, n17442, n17443, 
      n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, 
      n17454, n17457, n17458, n17460, n17461, n17462, n17463, n17464, n17465, 
      n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, 
      n17475, n17476, n17477, n17478, n17479, n17480, n17482, n17483, n17485, 
      n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, 
      n17495, n17496, n17497, n17498, n17499, n17501, n17502, n17503, n17504, 
      n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17513, n17514, 
      n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, 
      n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, 
      n17533, n17534, n17538, n17539, n17540, n17541, n17542, n17543, n17545, 
      n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17554, n17555, 
      n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, 
      n17565, n17566, n17567, n17568, n17569, n17570, n17573, n17574, n17575, 
      n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, 
      n17586, n17587, n17588, n17591, n17594, n17595, n17596, n17597, n17598, 
      n17599, n17600, n17601, n17602, n17603, n17605, n17606, n17607, n17608, 
      n17609, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, 
      n17619, n17620, n17621, n17623, n17625, n17627, n17628, n17629, n17630, 
      n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17640, n17641, 
      n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17651, 
      n17653, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, 
      n17664, n17665, n17666, n17669, n17670, n17671, n17672, n17674, n17675, 
      n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, 
      n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17694, n17695, 
      n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17707, 
      n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17718, 
      n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, 
      n17729, n17731, n17732, n17733, n17734, n17735, n17737, n17738, n17739, 
      n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, 
      n17750, n17751, n17752, n17753, n17754, n17755, n17757, n17758, n17759, 
      n17760, n17761, n17762, n17764, n17765, n17766, n17767, n17768, n17769, 
      n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, 
      n17779, n17780, n17782, n17783, n17784, n17785, n17787, n17788, n17789, 
      n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, 
      n17800, n17801, n17802, n17803, n17805, n17806, n17807, n17809, n17810, 
      n17811, n17812, n17813, n17815, n17816, n17817, n17818, n17819, n17820, 
      n17822, n17823, n17824, n17826, n17827, n17828, n17830, n17831, n17833, 
      n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17842, n17843, 
      n17844, n17845, n17847, n17848, n17850, n17852, n17854, n17855, n17856, 
      n17858, n17859, n17860, n17861, n17862, n17864, n17865, n17866, n17867, 
      n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17876, n17878, 
      n17880, n17881, n17884, n17885, n17887, n17888, n17889, n17891, n17892, 
      n17893, n17894, n17895, n17897, n17898, n17900, n17902, n17903, n17904, 
      n17905, n17906, n17909, n17910, n17912, n17914, n17915, n17917, n17918, 
      n17919, n17920, n17921, n17922, n17924, n17925, n17926, n17927, n17928, 
      n17929, n17931, n17933, n17934, n17935, n17937, n17938, n17939, n17940, 
      n17941, n17942, n17943, n17945, n17947, n17948, n17950, n17952, n17953, 
      n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, 
      n17963, n17964, n17966, n17967, n17968, n17969, n17970, n17971, n17972, 
      n17974, n17975, n17976, n17977, n17979, n17980, n17981, n17983, n17984, 
      n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, 
      n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18002, n18003, 
      n18004, n18005, n18006, n18008, n18009, n18010, n18011, n18012, n18013, 
      n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, 
      n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, 
      n18033, n18034, n18035, n18036, n18038, n18039, n18040, n18041, n18043, 
      n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18052, n18053, 
      n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, 
      n18063, n18064, n18065, n18066, n18068, n18069, n18070, n18071, n18072, 
      n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, 
      n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, 
      n18091, n18092, n18095, n18097, n18099, n18100, n18101, n18102, n18103, 
      n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, 
      n18113, n18114, n18115, n18116, n18118, n18119, n18120, n18121, n18122, 
      n18123, n18124, n18125, n18128, n18129, n18130, n18131, n18132, n18133, 
      n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18142, n18144, 
      n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, 
      n18154, n18155, n18157, n18158, n18159, n18160, n18161, n18162, n18163, 
      n18164, n18166, n18167, n18168, n18169, n18171, n18172, n18173, n18174, 
      n18175, n18176, n18177, n18179, n18180, n18181, n18182, n18183, n18184, 
      n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18193, n18194, 
      n18196, n18197, n18198, n18199, n18201, n18202, n18203, n18204, n18205, 
      n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18214, n18215, 
      n18216, n18217, n18218, n18219, n18221, n18222, n18223, n18224, n18225, 
      n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, 
      n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, 
      n18244, n18245, n18246, n18249, n18250, n18251, n18253, n18254, n18256, 
      n18257, n18258, n18260, n18261, n18262, n18263, n18264, n18265, n18266, 
      n18267, n18269, n18270, n18272, n18273, n18274, n18275, n18276, n18278, 
      n18279, n18280, n18282, n18283, n18284, n18286, n18287, n18288, n18289, 
      n18290, n18291, n18292, n18293, n18294, n18297, n18299, n18300, n18301, 
      n18302, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, 
      n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18321, n18322, 
      n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, 
      n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, 
      n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18350, n18351, 
      n18352, n18353, n18355, n18356, n18357, n18359, n18360, n18361, n18362, 
      n18363, n18365, n18366, n18368, n18369, n18370, n18371, n18372, n18375, 
      n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18385, 
      n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, 
      n18396, n18398, n18399, n18401, n18402, n18404, n18405, n18406, n18407, 
      n18409, n18410, n18412, n18413, n18414, n18415, n18416, n18417, n18418, 
      n18419, n18420, n18421, n18422, n18424, n18425, n18426, n18427, n18428, 
      n18429, n18432, n18434, n18435, n18436, n18437, n18438, n18439, n18442, 
      n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, 
      n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18460, n18461, 
      n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18472, 
      n18473, n18474, n18475, n18476, n18478, n18479, n18480, n18481, n18482, 
      n18483, n18484, n18487, n18488, n18489, n18490, n18491, n18493, n18494, 
      n18495, n18496, n18497, n18498, n18499, n18501, n18504, n18505, n18506, 
      n18507, n18509, n18510, n18511, n18512, n18515, n18516, n18518, n18519, 
      n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, 
      n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18537, n18538, 
      n18539, n18540, n18541, n18543, n18544, n18545, n18546, n18547, n18548, 
      n18549, n18551, n18552, n18554, n18555, n18556, n18557, n18561, n18563, 
      n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, 
      n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, 
      n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, 
      n18592, n18595, n18597, n18599, n18600, n18601, n18602, n18603, n18604, 
      n18605, n18606, n18608, n18609, n18610, n18611, n18612, n18613, n18615, 
      n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, 
      n18625, n18626, n18627, n18628, n18629, n18630, n18633, n18634, n18635, 
      n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18645, n18646, 
      n18648, n18649, n18651, n18653, n18654, n18655, n18656, n18657, n18658, 
      n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, 
      n18669, n18670, n18672, n18673, n18674, n18675, n18676, n18677, n18682, 
      n18683, n18684, n18685, n18686, n18687, n18688, n18690, n18691, n18692, 
      n18693, n18694, n18696, n18697, n18698, n18699, n18700, n18702, n18703, 
      n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, 
      n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, 
      n18723, n18724, n18725, n18726, n18727, n18728, n18730, n18731, n18732, 
      n18733, n18736, n18737, n18739, n18740, n18741, n18742, n18743, n18744, 
      n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, 
      n18755, n18756, n18757, n18759, n18760, n18761, n18763, n18764, n18765, 
      n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18776, 
      n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, 
      n18786, n18787, n18789, n18790, n18791, n18793, n18794, n18795, n18796, 
      n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18806, 
      n18807, n18808, n18810, n18811, n18812, n18813, n18814, n18815, n18816, 
      n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, 
      n18826, n18827, n18828, n18829, n18830, n18831, n18833, n18836, n18837, 
      n18838, n18839, n18840, n18841, n18845, n18847, n18851, n18852, n18854, 
      n18855, n18856, n18857, n18858, n18860, n18861, n18862, n18863, n18864, 
      n18866, n18869, n18871, n18872, n18873, n18875, n18876, n18877, n18879, 
      n18882, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, 
      n18897, n18898, n18899, n18900, n18903, n18904, n18905, n18906, n18907, 
      n18908, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, 
      n18918, n18919, n18920, n18921, n18923, n18924, n18925, n18926, n18927, 
      n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, 
      n18937, n18938, n18939, n18940, n18942, n18943, n18944, n18945, n18946, 
      n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18956, n18958, 
      n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18968, 
      n18970, n18971, n18972, n18974, n18975, n18976, n18977, n18980, n18982, 
      n18983, n18984, n18985, n18990, n18991, n18992, n18993, n18994, n18995, 
      n18996, n18997, n18999, n19000, n19001, n19002, n19003, n19004, n19005, 
      n19006, n19007, n19008, n19009, n19010, n19011, n19013, n19014, n19015, 
      n19016, n19017, n19018, n19019, n19021, n19022, n19023, n19024, n19025, 
      n19026, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, 
      n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, 
      n19045, n19046, n19048, n19052, n19053, n19054, n19055, n19056, n19057, 
      n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, 
      n19067, n19068, n19071, n19072, n19073, n19074, n19075, n19077, n19078, 
      n19079, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, 
      n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, 
      n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, 
      n19108, n19109, n19110, n19112, n19113, n19114, n19115, n19116, n19117, 
      n19120, n19121, n19122, n19123, n19124, n19126, n19128, n19129, n19131, 
      n19132, n19133, n19134, n19135, n19136, n19138, n19140, n19141, n19142, 
      n19143, n19144, n19145, n19146, n19147, n19148, n19150, n19151, n19152, 
      n19153, n19154, n19155, n19156, n19157, n19159, n19160, n19161, n19163, 
      n19164, n19165, n19166, n19167, n19168, n19169, n19171, n19172, n19173, 
      n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19182, n19183, 
      n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, 
      n19193, n19194, n19195, n19196, n19198, n19199, n19200, n19201, n19202, 
      n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, 
      n19212, n19213, n19214, n19216, n19218, n19219, n19220, n19222, n19223, 
      n19224, n19225, n19226, n19227, n19228, n19231, n19233, n19234, n19235, 
      n19236, n19237, n19238, n19239, n19240, n19242, n19243, n19244, n19246, 
      n19247, n19248, n19250, n19251, n19252, n19253, n19254, n19255, n19256, 
      n19257, n19258, n19260, n19261, n19262, n19264, n19265, n19266, n19267, 
      n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19276, n19277, 
      n19278, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, 
      n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, 
      n19298, n19299, n19300, n19302, n19303, n19304, n19305, n19306, n19307, 
      n19308, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, 
      n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, 
      n19328, n19329, n19330, n19331, n19333, n19334, n19335, n19336, n19338, 
      n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, 
      n19348, n19349, n19350, n19351, n19352, n19353, n19355, n19356, n19357, 
      n19358, n19359, n19360, n19361, n19362, n19363, n19365, n19366, n19367, 
      n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, 
      n19377, n19378, n19379, n19382, n19383, n19384, n19385, n19386, n19387, 
      n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19397, 
      n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, 
      n19408, n19409, n19410, n19411, n19412, n19414, n19415, n19416, n19418, 
      n19419, n19420, n19421, n19423, n19424, n19425, n19426, n19427, n19428, 
      n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, 
      n19440, n19441, n19443, n19444, n19445, n19446, n19447, n19448, n19449, 
      n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19460, n19461, 
      n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19472, 
      n19473, n19474, n19477, n19478, n19479, n19480, n19481, n19482, n19483, 
      n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19492, n19493, 
      n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, 
      n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, 
      n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, 
      n19521, n19522, n19523, n19524, n19526, n19527, n19528, n19529, n19530, 
      n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, 
      n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, 
      n19550, n19551, n19552, n19554, n19555, n19556, n19557, n19558, n19559, 
      n19560, n19562, n19563, n19564, n19565, n19568, n19570, n19571, n19572, 
      n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19582, 
      n19584, n19585, n19586, n19587, n19590, n19592, n19593, n19595, n19596, 
      n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, 
      n19606, n19607, n19608, n19610, n19611, n19612, n19614, n19615, n19616, 
      n19617, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, 
      n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, 
      n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, 
      n19647, n19649, n19650, n19651, n19652, n19656, n19658, n19659, n19660, 
      n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, 
      n19670, n19671, n19672, n19673, n19675, n19676, n19677, n19678, n19679, 
      n19681, n19682, n19683, n19684, n19685, n19688, n19689, n19690, n19691, 
      n19692, n19693, n19694, n19695, n19696, n19697, n19699, n19700, n19701, 
      n19702, n19705, n19706, n19707, n19709, n19711, n19712, n19713, n19714, 
      n19715, n19716, n19717, n19718, n19720, n19721, n19722, n19723, n19724, 
      n19725, n19726, n19727, n19728, n19730, n19731, n19733, n19734, n19735, 
      n19736, n19737, n19738, n19739, n19741, n19742, n19743, n19744, n19745, 
      n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, 
      n19755, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, 
      n19765, n19766, n19767, n19768, n19770, n19771, n19774, n19775, n19776, 
      n19778, n19779, n19781, n19782, n19783, n19784, n19785, n19786, n19788, 
      n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, 
      n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19808, 
      n19809, n19810, n19812, n19813, n19814, n19815, n19816, n19817, n19818, 
      n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, 
      n19828, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, 
      n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, 
      n19847, n19848, n19849, n19850, n19853, n19854, n19855, n19857, n19858, 
      n19859, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, 
      n19869, n19870, n19871, n19872, n19873, n19875, n19876, n19877, n19878, 
      n19880, n19882, n19883, n19884, n19885, n19886, n19888, n19889, n19890, 
      n19891, n19892, n19893, n19895, n19898, n19899, n19901, n19903, n19905, 
      n19906, n19907, n19908, n19911, n19912, n19913, n19914, n19915, n19916, 
      n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19925, n19926, 
      n19928, n19930, n19931, n19932, n19934, n19935, n19936, n19937, n19938, 
      n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, 
      n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, 
      n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, 
      n19968, n19969, n19971, n19972, n19973, n19974, n19975, n19976, n19978, 
      n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, 
      n19988, n19989, n19991, n19992, n19996, n19998, n19999, n20000, n20001, 
      n20003, n20005, n20006, n20007, n20008, n20011, n20012, n20016, n20018, 
      n20019, n20021, n20022, n20023, n20024, n20025, n20029, n20030, n20031, 
      n20032, n20033, n20034, n20036, n20037, n20038, n20039, n20040, n20041, 
      n20043, n20044, n20045, n20047, n20049, n20050, n20051, n20052, n20053, 
      n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, 
      n20063, n20064, n20065, n20066, n20068, n20070, n20071, n20072, n20073, 
      n20074, n20075, n20076, n20078, n20080, n20082, n20083, n20084, n20085, 
      n20087, n20088, n20089, n20090, n20091, n20092, n20094, n20096, n20097, 
      n20098, n20099, n20100, n20101, n20102, n20105, n20106, n20107, n20108, 
      n20110, n20111, n20112, n20113, n20114, n20116, n20118, n20119, n20121, 
      n20122, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, 
      n20132, n20133, n20135, n20136, n20137, n20138, n20139, n20141, n20142, 
      n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, 
      n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20161, n20162, 
      n20163, n20164, n20165, n20166, n20168, n20171, n20173, n20174, n20176, 
      n20177, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, 
      n20188, n20189, n20190, n20192, n20193, n20194, n20195, n20196, n20197, 
      n20198, n20199, n20200, n20201, n20203, n20205, n20206, n20207, n20208, 
      n20209, n20210, n20213, n20214, n20215, n20216, n20217, n20219, n20220, 
      n20221, n20222, n20223, n20224, n20225, n20226, n20231, n20232, n20233, 
      n20234, n20235, n20237, n20238, n20239, n20240, n20241, n20244, n20245, 
      n20246, n20247, n20248, n20249, n20250, n20252, n20253, n20254, n20255, 
      n20256, n20259, n20260, n20261, n20262, n20263, n20267, n20268, n20269, 
      n20270, n20271, n20272, n20273, n20276, n20277, n20278, n20279, n20280, 
      n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, 
      n20290, n20291, n20292, n20294, n20295, n20298, n20300, n20301, n20302, 
      n20303, n20304, n20307, n20308, n20309, n20310, n20311, n20312, n20313, 
      n20314, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, 
      n20324, n20326, n20328, n20329, n20330, n20332, n20334, n20335, n20336, 
      n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, 
      n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, 
      n20356, n20357, n20358, n20359, n20361, n20362, n20363, n20364, n20365, 
      n20366, n20367, n20368, n20369, n20370, n20371, n20373, n20374, n20375, 
      n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, 
      n20385, n20387, n20388, n20389, n20392, n20393, n20394, n20395, n20396, 
      n20398, n20399, n20401, n20402, n20403, n20404, n20405, n20406, n20408, 
      n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, 
      n20418, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, 
      n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, 
      n20437, n20438, n20440, n20442, n20443, n20445, n20446, n20447, n20448, 
      n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, 
      n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, 
      n20467, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, 
      n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, 
      n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, 
      n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20504, 
      n20505, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, 
      n20515, n20516, n20517, n20518, n20519, n20521, n20522, n20523, n20524, 
      n20525, n20526, n20527, n20529, n20530, n20531, n20532, n20533, n20534, 
      n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20543, n20544, 
      n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, 
      n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, 
      n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, 
      n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, 
      n20583, n20584, n20585, n20586, n20587, n20588, n20590, n20591, n20592, 
      n20593, n20595, n20596, n20598, n20599, n20600, n20601, n20602, n20603, 
      n20604, n20605, n20607, n20608, n20609, n20610, n20611, n20612, n20613, 
      n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20623, 
      n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20633, 
      n20634, n20635, n20636, n20637, n20638, n20639, n20642, n20643, n20644, 
      n20645, n20647, n20648, n20649, n20650, n20652, n20653, n20654, n20655, 
      n20656, n20657, n20658, n20659, n20660, n20662, n20663, n20664, n20665, 
      n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, 
      n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20687, 
      n20688, n20689, n20691, n20692, n20693, n20694, n20695, n20696, n20697, 
      n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20707, n20709, 
      n20710, n20711, n20713, n20714, n20716, n20718, n20719, n20720, n20721, 
      n20722, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, 
      n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, 
      n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, 
      n20750, n20751, n20752, n20753, n20754, n20755, n20757, n20758, n20760, 
      n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, 
      n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20779, 
      n20780, n20781, n20783, n20784, n20785, n20786, n20787, n20788, n20789, 
      n20791, n20792, n20793, n20795, n20796, n20797, n20798, n20799, n20800, 
      n20801, n20802, n20803, n20804, n20807, n20809, n20810, n20811, n20812, 
      n20813, n20815, n20816, n20817, n20818, n20819, n20821, n20822, n20823, 
      n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20833, n20835, 
      n20836, n20837, n20838, n20840, n20842, n20843, n20844, n20845, n20846, 
      n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, 
      n20856, n20857, n20858, n20860, n20861, n20862, n20863, n20864, n20865, 
      n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, 
      n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, 
      n20884, n20885, n20887, n20888, n20889, n20890, n20891, n20892, n20893, 
      n20894, n20895, n20897, n20898, n20899, n20900, n20901, n20902, n20903, 
      n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, 
      n20913, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, 
      n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, 
      n20932, n20933, n20935, n20936, n20938, n20939, n20940, n20941, n20943, 
      n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, 
      n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, 
      n20965, n20966, n20967, n20968, n20969, n20971, n20972, n20973, n20974, 
      n20975, n20976, n20977, n20979, n20980, n20981, n20982, n20984, n20986, 
      n20987, n20988, n20989, n20990, n20992, n20993, n20994, n20995, n20997, 
      n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, 
      n21007, n21008, n21009, n21010, n21012, n21013, n21014, n21015, n21016, 
      n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, 
      n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, 
      n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21047, n21048, 
      n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, 
      n21059, n21061, n21062, n21063, n21064, n21066, n21068, n21069, n21070, 
      n21071, n21072, n21073, n21074, n21075, n21077, n21078, n21079, n21080, 
      n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21090, 
      n21091, n21092, n21094, n21095, n21096, n21097, n21098, n21099, n21100, 
      n21101, n21102, n21104, n21105, n21106, n21107, n21109, n21110, n21111, 
      n21112, n21113, n21114, n21116, n21118, n21120, n21121, n21122, n21123, 
      n21124, n21125, n21126, n21127, n21128, n21129, n21131, n21133, n21134, 
      n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, 
      n21144, n21145, n21147, n21148, n21149, n21150, n21151, n21152, n21153, 
      n21154, n21155, n21156, n21157, n21158, n21160, n21161, n21162, n21163, 
      n21164, n21165, n21166, n21168, n21169, n21170, n21172, n21173, n21174, 
      n21175, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, 
      n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, 
      n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, 
      n21205, n21208, n21210, n21211, n21212, n21213, n21214, n21215, n21216, 
      n21217, n21218, n21219, n21220, n21221, n21222, n21225, n21226, n21227, 
      n21228, n21230, n21232, n21233, n21234, n21235, n21237, n21238, n21239, 
      n21240, n21241, n21243, n21244, n21245, n21247, n21249, n21250, n21251, 
      n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, 
      n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21270, 
      n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, 
      n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21288, n21289, 
      n21290, n21291, n21292, n21293, n21294, n21295, n21297, n21298, n21299, 
      n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, 
      n21309, n21311, n21313, n21314, n21315, n21316, n21317, n21318, n21320, 
      n21322, n21323, n21324, n21325, n21327, n21328, n21330, n21331, n21332, 
      n21335, n21336, n21338, n21339, n21340, n21341, n21342, n21343, n21344, 
      n21345, n21347, n21348, n21349, n21352, n21353, n21354, n21355, n21356, 
      n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, 
      n21366, n21367, n21368, n21369, n21370, n21371, n21373, n21374, n21375, 
      n21376, n21377, n21378, n21379, n21380, n21381, n21383, n21384, n21385, 
      n21386, n21387, n21388, n21389, n21392, n21393, n21394, n21395, n21396, 
      n21397, n21398, n21399, n21401, n21402, n21403, n21404, n21405, n21406, 
      n21407, n21408, n21409, n21411, n21412, n21413, n21414, n21415, n21416, 
      n21418, n21419, n21420, n21421, n21422, n21424, n21426, n21427, n21428, 
      n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21438, 
      n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21449, 
      n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, 
      n21459, n21460, n21462, n21463, n21464, n21465, n21467, n21468, n21469, 
      n21470, n21471, n21473, n21474, n21475, n21476, n21477, n21478, n21479, 
      n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, 
      n21490, n21491, n21495, n21496, n21498, n21499, n21500, n21501, n21502, 
      n21504, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, 
      n21514, n21515, n21516, n21517, n21519, n21520, n21521, n21522, n21523, 
      n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, 
      n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21542, 
      n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, 
      n21552, n21553, n21554, n21555, n21556, n21557, n21561, n21563, n21564, 
      n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21574, 
      n21576, n21578, n21579, n21580, n21581, n21584, n21586, n21587, n21588, 
      n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, 
      n21599, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, 
      n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21618, 
      n21619, n21620, n21621, n21622, n21623, n21624, n21626, n21627, n21628, 
      n21629, n21630, n21631, n21632, n21634, n21635, n21636, n21637, n21638, 
      n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, 
      n21648, n21649, n21650, n21651, n21653, n21655, n21656, n21658, n21659, 
      n21660, n21663, n21664, n21666, n21667, n21668, n21669, n21670, n21671, 
      n21673, n21674, n21675, n21676, n21678, n21679, n21680, n21681, n21682, 
      n21683, n21684, n21685, n21686, n21689, n21690, n21691, n21692, n21693, 
      n21695, n21696, n21697, n21698, n21699, n21700, n21702, n21703, n21704, 
      n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, 
      n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, 
      n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21732, 
      n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, 
      n21742, n21753, n21754, n21756, n21757, n21758, n21759, n21760, n21761, 
      n21764, n21765, n21767, n21768, n21769, n21772, n21773, n21774, n21775, 
      n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, 
      n21785, n21786, n21787, n21788, n21790, n21791, n21792, n21793, n21795, 
      n21798, n21799, n21800, n21801, n21804, n21807, n21808, n21809, n21812, 
      n21813, n21814, n21816, n21818, n21819, n21820, n21821, n21822, n21824, 
      n21825, n21826, n21827, n21829, n21830, n21831, n21832, n21833, n21834, 
      n21837, n21838, n21839, n21841, n21842, n21843, n21845, n21846, n21848, 
      n21850, n21852, n21854, n21855, n21856, n21857, n21859, n21860, n21861, 
      n21863, n21865, n21866, n21867, n21868, n21869, n21871, n21872, n21873, 
      n21874, n21875, n21876, n21877, n21879, n21880, n21881, n21882, n21885, 
      n21886, n21888, n21890, n21891, n21892, n21893, n21894, n21895, n21896, 
      n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, 
      n21906, n21907, n21908, n21909, n21911, n21912, n21914, n21915, n21916, 
      n21917, n21918, n21919, n21920, n21922, n21923, n21924, n21926, n21927, 
      n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21936, n21937, 
      n21938, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21948, 
      n21949, n21952, n21957, n21958, n21959, n21961, n21962, n21963, n21964, 
      n21965, n21969, n21970, n21974, n21979, n21980, n21983, n21984, n21985, 
      n21986, n21987, n21988, n21989, n21992, n21993, n21994, n21995, n21998, 
      n21999, n22000, n22001, n22005, n22008, n22010, n22011, n22012, n22015, 
      n22016, n22017, n22018, n22019, n22022, n22025, n22027, n22031, n22033, 
      n22035, n22036, n22040, n22041, n22043, n22044, n22045, n22046, n22047, 
      n22050, n22051, n22052, n22054, n22055, n22056, n22057, n22060, n22061, 
      n22066, n22069, n22071, n22073, n22075, n22077, n22080, n22081, n22082, 
      n22085, n22086, n22087, n22091, n22092, n22093, n22096, n22097, n22099, 
      n22102, n22104, n22105, n22106, n22108, n22109, n22110, n22111, n22112, 
      n22113, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, 
      n22123, n22126, n22127, n22128, n22129, n22130, n22135, n22139, n22140, 
      n22142, n22143, n22144, n22146, n22148, n22150, n22153, n22154, n22155, 
      n22157, n22158, n22159, n22162, n22163, n22164, n22165, n22169, n22170, 
      n22171, n22172, n22174, n22175, n22176, n22178, n22183, n22184, n22185, 
      n22190, n22191, n22192, n22194, n22195, n22196, n22197, n22198, n22199, 
      n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, 
      n22212, n22213, n22214, n22216, n22217, n22218, n22221, n22224, n22226, 
      n22227, n22234, n22237, n22238, n22239, n22240, n22241, n22242, n22244, 
      n22247, n22252, n22253, n22254, n22256, n22257, n22259, n22260, n22263, 
      n22264, n22265, n22266, n22267, n22269, n22272, n22273, n22274, n22275, 
      n22277, n22279, n22280, n22281, n22282, n22285, n22287, n22288, n22289, 
      n22290, n22291, n22295, n22296, n22299, n22302, n22303, n22305, n22306, 
      n22307, n22309, n22311, n22312, n22313, n22314, n22315, n22319, n22322, 
      n22325, n22326, n22329, n22330, n22331, n22333, n22335, n22337, n22338, 
      n22339, n22340, n22341, n22342, n22343, n22345, n22346, n22347, n22349, 
      n22353, n22354, n22357, n22358, n22363, n22364, n22365, n22370, n22371, 
      n22373, n22374, n22376, n22377, n22378, n22380, n22381, n22383, n22385, 
      n22386, n22387, n22388, n22391, n22392, n22393, n22396, n22398, n22399, 
      n22401, n22402, n22404, n22405, n22407, n22409, n22411, n22415, n22417, 
      n22418, n22420, n22421, n22422, n22423, n22424, n22425, n22427, n22429, 
      n22430, n22432, n22436, n22437, n22438, n22439, n22440, n22444, n22445, 
      n22446, n22449, n22450, n22451, n22453, n22454, n22457, n22458, n22459, 
      n22460, n22463, n22466, n22470, n22471, n22472, n22475, n22478, n22482, 
      n22483, n22484, n22485, n22487, n22489, n22490, n22492, n22493, n22494, 
      n22496, n22498, n22500, n22501, n22504, n22505, n22506, n22508, n22510, 
      n22511, n22512, n22514, n22515, n22516, n22517, n22518, n22519, n22522, 
      n22523, n22524, n22525, n22526, n22528, n22529, n22531, n22533, n22536, 
      n22537, n22538, n22540, n22541, n22542, n22544, n22546, n22547, n22548, 
      n22551, n22552, n22554, n22555, n22556, n22557, n22558, n22559, n22560, 
      n22561, n22563, n22566, n22567, n22568, n22569, n22570, n22571, n22572, 
      n22574, n22575, n22576, n22577, n22578, n22579, n22581, n22584, n22585, 
      n22587, n22589, n22590, n22591, n22592, n22594, n22596, n22597, n22598, 
      n22599, n22600, n22602, n22603, n22604, n22605, n22607, n22609, n22612, 
      n22613, n22614, n22616, n22617, n22619, n22620, n22621, n22622, n22623, 
      n22624, n22625, n22626, n22628, n22629, n22630, n22631, n22632, n22633, 
      n22634, n22635, n22637, n22640, n22641, n22642, n22643, n22645, n22646, 
      n22647, n22648, n22649, n22650, n22652, n22653, n22654, n22655, n22657, 
      n22658, n22659, n22660, n22666, n22668, n22671, n22672, n22673, n22674, 
      n22676, n22678, n22679, n22680, n22681, n22684, n22686, n22687, n22688, 
      n22689, n22691, n22692, n22693, n22694, n22695, n22696, n22698, n22699, 
      n22700, n22701, n22703, n22704, n22705, n22707, n22709, n22710, n22711, 
      n22712, n22715, n22716, n22718, n22719, n22724, n22725, n22726, n22727, 
      n22728, n22729, n22730, n22731, n22732, n22734, n22735, n22736, n22737, 
      n22738, n22739, n22740, n22741, n22743, n22744, n22745, n22746, n22747, 
      n22748, n22749, n22750, n22751, n22753, n22755, n22756, n22757, n22758, 
      n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, 
      n22768, n22770, n22771, n22773, n22774, n22775, n22776, n22777, n22778, 
      n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22788, 
      n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, 
      n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22806, n22807, 
      n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22817, n22818, 
      n22819, n22820, n22821, n22823, n22824, n22825, n22826, n22828, n22829, 
      n22830, n22831, n22832, n22834, n22835, n22836, n22837, n22838, n22839, 
      n22840, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, 
      n22851, n22855, n22856, n22860, n22862, n22863, n22864, n22865, n22866, 
      n22868, n22869, n22871, n22873, n22875, n22876, n22877, n22879, n22880, 
      n22881, n22882, n22883, n22886, n22887, n22888, n22889, n22890, n22891, 
      n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22900, n22901, 
      n22902, n22903, n22905, n22906, n22907, n22908, n22910, n22912, n22913, 
      n22914, n22916, n22918, n22919, n22920, n22921, n22924, n22925, n22926, 
      n22927, n22929, n22931, n22932, n22935, n22936, n22937, n22938, n22939, 
      n22940, n22942, n22943, n22944, n22946, n22949, n22950, n22954, n22955, 
      n22956, n22958, n22959, n22960, n22961, n22962, n22965, n22967, n22969, 
      n22973, n22974, n22975, n22977, n22978, n22979, n22981, n22983, n22984, 
      n22986, n22987, n22988, n22990, n22991, n22993, n22994, n22995, n22996, 
      n22997, n22998, n23000, n23001, n23002, n23004, n23005, n23006, n23007, 
      n23010, n23011, n23012, n23013, n23014, n23017, n23018, n23019, n23020, 
      n23021, n23022, n23023, n23025, n23026, n23029, n23030, n23031, n23032, 
      n23034, n23035, n23036, n23037, n23040, n23041, n23042, n23043, n23044, 
      n23046, n23047, n23048, n23053, n23054, n23055, n23056, n23057, n23059, 
      n23060, n23062, n23063, n23064, n23065, n23066, n23067, n23069, n23070, 
      n23071, n23072, n23073, n23074, n23075, n23079, n23081, n23083, n23086, 
      n23087, n23088, n23092, n23093, n23094, n23096, n23097, n23098, n23102, 
      n23103, n23104, n23105, n23107, n23109, n23110, n23111, n23113, n23115, 
      n23116, n23117, n23118, n23119, n23120, n23124, n23125, n23126, n23127, 
      n23128, n23129, n23130, n23134, n23135, n23137, n23138, n23139, n23141, 
      n23142, n23143, n23145, n23146, n23147, n23150, n23151, n23154, n23156, 
      n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23165, n23166, 
      n23167, n23168, n23169, n23170, n23171, n23173, n23175, n23178, n23180, 
      n23181, n23183, n23184, n23185, n23186, n23187, n23188, n23191, n23196, 
      n23197, n23198, n23199, n23201, n23202, n23203, n23204, n23205, n23209, 
      n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23219, n23220, 
      n23221, n23222, n23223, n23225, n23226, n23227, n23228, n23229, n23231, 
      n23232, n23233, n23236, n23238, n23239, n23243, n23244, n23245, n23247, 
      n23248, n23251, n23253, n23255, n23256, n23258, n23259, n23260, n23261, 
      n23264, n23267, n23268, n23269, n23270, n23274, n23275, n23276, n23277, 
      n23278, n23279, n23283, n23284, n23285, n23287, n23288, n23291, n23294, 
      n23295, n23296, n23301, n23302, n23304, n23305, n23306, n23307, n23309, 
      n23311, n23312, n23313, n23314, n23315, n23318, n23319, n23322, n23323, 
      n23325, n23327, n23329, n23331, n23332, n23333, n23334, n23335, n23336, 
      n23337, n23338, n23339, n23341, n23343, n23344, n23345, n23346, n23347, 
      n23349, n23352, n23354, n23355, n23356, n23357, n23359, n23361, n23362, 
      n23363, n23365, n23367, n23368, n23369, n23371, n23373, n23374, n23375, 
      n23379, n23380, n23383, n23386, n23390, n23391, n23392, n23393, n23395, 
      n23399, n23401, n23405, n23407, n23408, n23409, n23411, n23413, n23414, 
      n23415, n23416, n23418, n23419, n23420, n23421, n23422, n23423, n23424, 
      n23426, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, 
      n23436, n23437, n23438, n23439, n23440, n23441, n23443, n23444, n23445, 
      n23448, n23449, n23450, n23453, n23454, n23455, n23456, n23457, n23462, 
      n23463, n23466, n23467, n23469, n23471, n23474, n23475, n23477, n23478, 
      n23479, n23480, n23481, n23482, n23484, n23485, n23486, n23488, n23492, 
      n23494, n23497, n23499, n23500, n23501, n23502, n23504, n23505, n23507, 
      n23508, n23510, n23512, n23514, n23515, n23518, n23525, n23528, n23529, 
      n23530, n23531, n23533, n23534, n23535, n23536, n23537, n23538, n23539, 
      n23540, n23542, n23544, n23546, n23547, n23548, n23552, n23553, n23554, 
      n23556, n23557, n23558, n23559, n23561, n23563, n23564, n23565, n23567, 
      n23568, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, 
      n23579, n23581, n23582, n23583, n23585, n23589, n23591, n23592, n23593, 
      n23594, n23597, n23599, n23600, n23601, n23602, n23604, n23607, n23608, 
      n23609, n23610, n23613, n23614, n23616, n23617, n23618, n23620, n23621, 
      n23622, n23623, n23624, n23626, n23628, n23630, n23633, n23634, n23635, 
      n23636, n23637, n23638, n23641, n23642, n23643, n23644, n23645, n23646, 
      n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23656, n23657, 
      n23659, n23662, n23663, n23665, n23666, n23667, n23668, n23669, n23671, 
      n23672, n23674, n23676, n23677, n23678, n23679, n23680, n23681, n23682, 
      n23683, n23684, n23686, n23687, n23689, n23691, n23692, n23694, n23696, 
      n23697, n23698, n23700, n23703, n23704, n23706, n23709, n23713, n23716, 
      n23717, n23718, n23719, n23720, n23722, n23723, n23724, n23725, n23726, 
      n23727, n23728, n23730, n23731, n23732, n23735, n23736, n23737, n23739, 
      n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23748, n23749, 
      n23750, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23760, 
      n23761, n23764, n23765, n23770, n23771, n23772, n23774, n23776, n23777, 
      n23778, n23779, n23780, n23781, n23782, n23784, n23786, n23787, n23788, 
      n23791, n23793, n23794, n23797, n23798, n23799, n23800, n23802, n23804, 
      n23805, n23806, n23808, n23809, n23810, n23811, n23812, n23815, n23816, 
      n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, 
      n23827, n23828, n23829, n23830, n23831, n23833, n23834, n23835, n23836, 
      n23837, n23839, n23840, n23841, n23842, n23844, n23845, n23846, n23849, 
      n23852, n23853, n23856, n23857, n23858, n23859, n23860, n23861, n23863, 
      n23864, n23865, n23867, n23868, n23869, n23870, n23871, n23872, n23873, 
      n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23883, 
      n23884, n23886, n23887, n23888, n23889, n23891, n23892, n23893, n23895, 
      n23896, n23897, n23898, n23899, n23903, n23904, n23905, n23906, n23907, 
      n23908, n23910, n23912, n23913, n23914, n23915, n23916, n23917, n23918, 
      n23919, n23920, n23922, n23923, n23926, n23927, n23928, n23929, n23931, 
      n23934, n23935, n23936, n23937, n23938, n23940, n23945, n23946, n23948, 
      n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, 
      n23960, n23963, n23966, n23967, n23968, n23969, n23970, n23971, n23973, 
      n23974, n23976, n23977, n23978, n23979, n23980, n23984, n23986, n23987, 
      n23990, n23991, n23992, n23993, n23996, n23998, n23999, n24000, n24003, 
      n24004, n24006, n24007, n24008, n24009, n24010, n24012, n24013, n24017, 
      n24018, n24019, n24022, n24025, n24026, n24027, n24028, n24029, n24032, 
      n24033, n24034, n24035, n24036, n24037, n24038, n24040, n24044, n24045, 
      n24047, n24048, n24049, n24050, n24051, n24052, n24054, n24055, n24056, 
      n24059, n24060, n24061, n24062, n24064, n24065, n24066, n24067, n24069, 
      n24070, n24071, n24072, n24075, n24076, n24077, n24078, n24079, n24080, 
      n24081, n24083, n24085, n24087, n24088, n24089, n24090, n24091, n24092, 
      n24093, n24094, n24095, n24096, n24097, n24098, n24102, n24103, n24104, 
      n24105, n24107, n24108, n24109, n24111, n24112, n24114, n24115, n24116, 
      n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24126, 
      n24127, n24130, n24132, n24133, n24134, n24135, n24136, n24138, n24141, 
      n24142, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, 
      n24152, n24153, n24154, n24155, n24156, n24157, n24159, n24160, n24162, 
      n24163, n24166, n24167, n24168, n24170, n24172, n24173, n24175, n24176, 
      n24177, n24178, n24179, n24181, n24182, n24183, n24184, n24185, n24186, 
      n24187, n24188, n24189, n24190, n24193, n24194, n24195, n24196, n24197, 
      n24198, n24199, n24200, n24201, n24202, n24205, n24206, n24207, n24208, 
      n24209, n24210, n24212, n24213, n24214, n24215, n24216, n24219, n24220, 
      n24221, n24223, n24224, n24225, n24227, n24228, n24230, n24231, n24232, 
      n24234, n24235, n24236, n24239, n24241, n24242, n24243, n24244, n24245, 
      n24247, n24248, n24249, n24251, n24253, n24254, n24255, n24258, n24259, 
      n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, 
      n24270, n24271, n24273, n24275, n24276, n24277, n24278, n24279, n24280, 
      n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24289, n24292, 
      n24293, n24294, n24295, n24297, n24299, n24302, n24304, n24306, n24307, 
      n24308, n24309, n24311, n24312, n24315, n24316, n24317, n24318, n24320, 
      n24321, n24322, n24323, n24324, n24325, n24327, n24328, n24329, n24330, 
      n24331, n24332, n24334, n24335, n24336, n24337, n24339, n24340, n24341, 
      n24343, n24344, n24345, n24347, n24349, n24350, n24351, n24356, n24357, 
      n24358, n24361, n24363, n24364, n24365, n24368, n24371, n24373, n24374, 
      n24376, n24377, n24379, n24380, n24381, n24382, n24383, n24384, n24386, 
      n24387, n24388, n24390, n24391, n24392, n24394, n24397, n24399, n24400, 
      n24403, n24405, n24406, n24407, n24408, n24413, n24414, n24415, n24416, 
      n24418, n24419, n24421, n24422, n24423, n24424, n24425, n24426, n24427, 
      n24429, n24430, n24431, n24432, n24433, n24437, n24438, n24439, n24440, 
      n24442, n24443, n24444, n24445, n24447, n24449, n24450, n24451, n24453, 
      n24454, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24466, 
      n24468, n24469, n24470, n24472, n24473, n24474, n24476, n24477, n24478, 
      n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24487, n24489, 
      n24491, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, 
      n24501, n24502, n24506, n24507, n24509, n24513, n24514, n24517, n24518, 
      n24520, n24522, n24523, n24524, n24525, n24528, n24529, n24530, n24531, 
      n24532, n24533, n24534, n24536, n24538, n24539, n24540, n24541, n24542, 
      n24545, n24547, n24548, n24549, n24550, n24552, n24553, n24554, n24558, 
      n24560, n24562, n24563, n24564, n24566, n24567, n24568, n24570, n24572, 
      n24573, n24574, n24575, n24576, n24577, n24579, n24580, n24581, n24582, 
      n24583, n24584, n24585, n24586, n24588, n24589, n24590, n24591, n24592, 
      n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, 
      n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24610, n24611, 
      n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620, 
      n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24630, 
      n24632, n24633, n24634, n24635, n24638, n24639, n24640, n24641, n24642, 
      n24643, n24644, n24645, n24646, n24648, n24649, n24650, n24651, n24652, 
      n24653, n24654, n24657, n24658, n24659, n24661, n24662, n24663, n24664, 
      n24665, n24666, n24667, n24668, n24669, n24670, n24672, n24673, n24674, 
      n24676, n24677, n24679, n24680, n24681, n24682, n24684, n24685, n24686, 
      n24687, n24688, n24691, n24693, n24695, n24696, n24697, n24699, n24700, 
      n24701, n24702, n24703, n24705, n24706, n24707, n24709, n24710, n24711, 
      n24712, n24714, n24715, n24718, n24719, n24720, n24723, n24725, n24727, 
      n24728, n24729, n24730, n24732, n24734, n24735, n24738, n24739, n24740, 
      n24741, n24742, n24743, n24744, n24745, n24747, n24749, n24750, n24752, 
      n24754, n24756, n24761, n24763, n24764, n24765, n24766, n24770, n24771, 
      n24772, n24773, n24774, n24775, n24779, n24781, n24783, n24785, n24786, 
      n24787, n24788, n24790, n24791, n24792, n24793, n24794, n24795, n24796, 
      n24797, n24798, n24800, n24801, n24802, n24804, n24805, n24806, n24807, 
      n24808, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, 
      n24818, n24820, n24821, n24825, n24829, n24830, n24831, n24832, n24833, 
      n24834, n24835, n24839, n24840, n24841, n24842, n24843, n24844, n24845, 
      n24846, n24847, n24848, n24849, n24851, n24852, n24853, n24854, n24855, 
      n24856, n24858, n24859, n24861, n24862, n24863, n24864, n24865, n24866, 
      n24867, n24868, n24870, n24872, n24874, n24875, n24877, n24878, n24879, 
      n24880, n24881, n24882, n24883, n24885, n24886, n24887, n24894, n24895, 
      n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, 
      n24906, n24910, n24912, n24914, n24916, n24917, n24919, n24921, n24922, 
      n24924, n24925, n24926, n24927, n24929, n24930, n24932, n24933, n24934, 
      n24935, n24936, n24937, n24938, n24941, n24944, n24946, n24950, n24951, 
      n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24960, n24961, 
      n24962, n24963, n24964, n24966, n24967, n24968, n24969, n24970, n24971, 
      n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24980, n24981, 
      n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, 
      n24995, n24996, n24997, n24998, n25000, n25002, n25003, n25004, n25005, 
      n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, 
      n25015, n25016, n25017, n25018, n25023, n25024, n25028, n25029, n25030, 
      n25034, n25035, n25036, n25037, n25038, n25039, n25042, n25043, n25045, 
      n25048, n25049, n25051, n25052, n25054, n25056, n25057, n25059, n25061, 
      n25063, n25064, n25066, n25067, n25068, n25069, n25070, n25071, n25072, 
      n25074, n25075, n25076, n25077, n25078, n25080, n25081, n25082, n25084, 
      n25086, n25087, n25090, n25092, n25093, n25094, n25095, n25096, n25097, 
      n25098, n25099, n25102, n25103, n25104, n25105, n25106, n25107, n25109, 
      n25110, n25111, n25113, n25114, n25115, n25116, n25118, n25119, n25120, 
      n25123, n25125, n25126, n25128, n25129, n25130, n25133, n25134, n25135, 
      n25136, n25137, n25138, n25140, n25141, n25143, n25144, n25145, n25147, 
      n25149, n25150, n25151, n25152, n25154, n25155, n25156, n25158, n25159, 
      n25161, n25162, n25163, n25165, n25166, n25167, n25168, n25170, n25171, 
      n25173, n25174, n25175, n25176, n25178, n25179, n25180, n25181, n25183, 
      n25184, n25185, n25186, n25188, n25191, n25192, n25195, n25196, n25197, 
      n25198, n25199, n25200, n25201, n25202, n25203, n25206, n25208, n25209, 
      n25212, n25214, n25215, n25216, n25217, n25218, n25222, n25224, n25225, 
      n25227, n25230, n25233, n25234, n25235, n25236, n25237, n25238, n25239, 
      n25240, n25241, n25242, n25243, n25245, n25246, n25247, n25249, n25252, 
      n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25261, n25262, 
      n25263, n25264, n25265, n25266, n25267, n25270, n25271, n25275, n25276, 
      n25277, n25278, n25279, n25280, n25282, n25283, n25284, n25287, n25288, 
      n25289, n25290, n25292, n25293, n25294, n25296, n25297, n25298, n25300, 
      n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, 
      n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25321, 
      n25322, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, 
      n25332, n25333, n25334, n25336, n25337, n25338, n25339, n25340, n25342, 
      n25343, n25345, n25346, n25347, n25348, n25349, n25351, n25352, n25353, 
      n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, 
      n25363, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, 
      n25373, n25374, n25375, n25376, n25377, n25378, n25380, n25381, n25382, 
      n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, 
      n25392, n25393, n25394, n25395, n25396, n25397, n25399, n25400, n25401, 
      n25403, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, 
      n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, 
      n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, 
      n25432, n25436, n25439, n25440, n25441, n25442, n25444, n25445, n25448, 
      n25449, n25450, n25451, n25453, n25455, n25457, n25458, n25459, n25460, 
      n25461, n25462, n25464, n25465, n25466, n25468, n25469, n25470, n25471, 
      n25474, n25476, n25477, n25478, n25479, n25481, n25482, n25484, n25485, 
      n25487, n25488, n25489, n25491, n25492, n25493, n25494, n25496, n25497, 
      n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25506, n25507, 
      n25508, n25509, n25511, n25514, n25515, n25517, n25518, n25520, n25521, 
      n25523, n25524, n25525, n25526, n25527, n25528, n25530, n25531, n25532, 
      n25533, n25534, n25535, n25536, n25538, n25540, n25541, n25542, n25543, 
      n25544, n25545, n25547, n25548, n25549, n25550, n25551, n25552, n25553, 
      n25554, n25557, n25559, n25560, n25561, n25562, n25563, n25564, n25566, 
      n25567, n25568, n25570, n25571, n25572, n25573, n25575, n25576, n25577, 
      n25578, n25579, n25582, n25583, n25584, n25585, n25586, n25590, n25591, 
      n25592, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, 
      n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, 
      n25614, n25616, n25617, n25618, n25619, n25621, n25622, n25624, n25626, 
      n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, 
      n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25644, n25645, 
      n25646, n25647, n25648, n25650, n25651, n25652, n25653, n25654, n25655, 
      n25657, n25658, n25659, n25660, n25662, n25664, n25665, n25666, n25668, 
      n25670, n25671, n25672, n25674, n25675, n25676, n25677, n25679, n25680, 
      n25681, n25683, n25684, n25685, n25687, n25688, n25689, n25692, n25693, 
      n25694, n25695, n25696, n25697, n25698, n25699, n25701, n25704, n25705, 
      n25707, n25708, n25709, n25710, n25712, n25713, n25714, n25717, n25718, 
      n25719, n25720, n25721, n25722, n25723, n25724, n25726, n25727, n25728, 
      n25729, n25730, n25731, n25732, n25733, n25734, n25736, n25738, n25739, 
      n25740, n25741, n25744, n25745, n25747, n25748, n25750, n25751, n25752, 
      n25753, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, 
      n25763, n25764, n25766, n25767, n25768, n25769, n25770, n25772, n25773, 
      n25774, n25778, n25779, n25780, n25781, n25784, n25785, n25786, n25787, 
      n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, 
      n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25806, n25807, 
      n25808, n25809, n25811, n25812, n25813, n25816, n25818, n25819, n25821, 
      n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, 
      n25831, n25833, n25834, n25835, n25837, n25838, n25840, n25841, n25843, 
      n25845, n25846, n25847, n25850, n25852, n25853, n25854, n25855, n25856, 
      n25857, n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, 
      n25867, n25868, n25869, n25870, n25871, n25873, n25874, n25875, n25877, 
      n25879, n25881, n25882, n25883, n25884, n25885, n25889, n25891, n25892, 
      n25894, n25896, n25898, n25899, n25900, n25901, n25902, n25903, n25904, 
      n25906, n25907, n25908, n25910, n25911, n25912, n25914, n25917, n25922, 
      n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25933, 
      n25934, n25935, n25936, n25938, n25939, n25940, n25941, n25942, n25943, 
      n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, 
      n25953, n25955, n25956, n25959, n25960, n25961, n25963, n25965, n25966, 
      n25968, n25969, n25970, n25971, n25973, n25975, n25977, n25979, n25980, 
      n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25991, n25993, 
      n25994, n25995, n25998, n25999, n26001, n26003, n26004, n26005, n26006, 
      n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, 
      n26017, n26018, n26020, n26021, n26022, n26023, n26024, n26027, n26028, 
      n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, 
      n26038, n26039, n26041, n26042, n26043, n26044, n26046, n26048, n26049, 
      n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, 
      n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, 
      n26068, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26078, 
      n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26087, n26088, 
      n26089, n26091, n26092, n26093, n26096, n26097, n26098, n26099, n26100, 
      n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110, 
      n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119, 
      n26120, n26121, n26122, n26123, n26124, n26126, n26128, n26129, n26130, 
      n26132, n26133, n26134, n26135, n26136, n26137, n26140, n26141, n26142, 
      n26143, n26144, n26145, n26146, n26147, n26149, n26150, n26152, n26153, 
      n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162, 
      n26163, n26165, n26166, n26167, n26168, n26169, n26170, n26172, n26173, 
      n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182, 
      n26183, n26186, n26187, n26189, n26191, n26192, n26193, n26194, n26195, 
      n26196, n26197, n26198, n26201, n26202, n26205, n26206, n26207, n26208, 
      n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, 
      n26218, n26219, n26220, n26221, n26222, n26223, n26226, n26227, n26228, 
      n26229, n26231, n26233, n26234, n26235, n26237, n26238, n26240, n26241, 
      n26243, n26244, n26246, n26248, n26252, n26254, n26255, n26256, n26257, 
      n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26266, n26267, 
      n26268, n26270, n26271, n26272, n26273, n26274, n26276, n26277, n26278, 
      n26279, n26280, n26281, n26282, n26283, n26284, n26286, n26287, n26288, 
      n26289, n26290, n26292, n26293, n26294, n26295, n26296, n26297, n26298, 
      n26299, n26300, n26301, n26302, n26303, n26305, n26306, n26307, n26308, 
      n26309, n26310, n26311, n26312, n26314, n26315, n26316, n26317, n26318, 
      n26319, n26321, n26323, n26324, n26325, n26326, n26327, n26329, n26330, 
      n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26342, 
      n26343, n26344, n26345, n26347, n26348, n26349, n26350, n26351, n26353, 
      n26354, n26355, n26356, n26357, n26358, n26361, n26362, n26363, n26364, 
      n26365, n26367, n26368, n26371, n26372, n26373, n26374, n26375, n26377, 
      n26378, n26380, n26381, n26382, n26384, n26386, n26387, n26388, n26389, 
      n26391, n26392, n26395, n26396, n26398, n26399, n26400, n26401, n26402, 
      n26403, n26405, n26406, n26408, n26409, n26410, n26412, n26413, n26414, 
      n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, 
      n26425, n26426, n26427, n26429, n26430, n26431, n26432, n26434, n26435, 
      n26436, n26437, n26438, n26439, n26440, n26443, n26445, n26446, n26447, 
      n26448, n26449, n26451, n26453, n26455, n26456, n26457, n26459, n26461, 
      n26462, n26463, n26464, n26465, n26469, n26471, n26472, n26473, n26476, 
      n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26485, n26486, 
      n26488, n26489, n26491, n26492, n26493, n26494, n26495, n26496, n26497, 
      n26498, n26499, n26500, n26501, n26503, n26504, n26505, n26507, n26510, 
      n26512, n26513, n26514, n26515, n26517, n26518, n26519, n26520, n26521, 
      n26522, n26523, n26527, n26528, n26531, n26532, n26533, n26535, n26536, 
      n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, 
      n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, 
      n26555, n26556, n26557, n26559, n26560, n26561, n26562, n26566, n26568, 
      n26569, n26570, n26574, n26575, n26576, n26577, n26578, n26579, n26580, 
      n26583, n26584, n26585, n26586, n26589, n26590, n26592, n26593, n26594, 
      n26598, n26599, n26600, n26601, n26603, n26604, n26606, n26607, n26608, 
      n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26620, 
      n26621, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, 
      n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, 
      n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26649, 
      n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, 
      n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, 
      n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, 
      n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, 
      n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, 
      n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, 
      n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, 
      n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, 
      n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, 
      n26731, n26732, n26733, n26734, n26737, n26738, n26739, n26740, n26741, 
      n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, 
      n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, 
      n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, 
      n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, 
      n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, 
      n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, 
      n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, 
      n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, 
      n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, 
      n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, 
      n26832, n26833, n26834, n26835, n26836, n26837, n26839, n26840, n26841, 
      n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, 
      n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, 
      n26860, n26861, n26862, n26863, n26864, n26866, n26867, n26868, n26869, 
      n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, 
      n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, 
      n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, 
      n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, 
      n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, 
      n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, 
      n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, 
      n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, 
      n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, 
      n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, 
      n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, 
      n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, 
      n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, 
      n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, 
      n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, 
      n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, 
      n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, 
      n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, 
      n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27041, 
      n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, 
      n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, 
      n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, 
      n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077, 
      n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086, 
      n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095, 
      n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, 
      n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113, 
      n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, 
      n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131, 
      n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, 
      n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, 
      n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158, 
      n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167, 
      n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176, 
      n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185, 
      n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194, 
      n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, 
      n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, 
      n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, 
      n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, 
      n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, 
      n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, 
      n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, 
      n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, 
      n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, 
      n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, 
      n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, 
      n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, 
      n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, 
      n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, 
      n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, 
      n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, 
      n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, 
      n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, 
      n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, 
      n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, 
      n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383, 
      n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392, 
      n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401, 
      n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410, 
      n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419, 
      n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428, 
      n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437, 
      n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446, 
      n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, 
      n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, 
      n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473, 
      n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482, 
      n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491, 
      n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500, 
      n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509, 
      n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, 
      n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, 
      n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, 
      n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, 
      n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, 
      n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, 
      n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, 
      n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, 
      n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, 
      n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, 
      n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, 
      n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, 
      n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, 
      n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, 
      n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, 
      n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, 
      n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, 
      n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, 
      n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, 
      n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, 
      n27691, n27692, n27694, n27695, n27696, n27697, n27698, n27699, n27700, 
      n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, 
      n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, 
      n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, 
      n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, 
      n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, 
      n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, 
      n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, 
      n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, 
      n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, 
      n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, 
      n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, 
      n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, 
      n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, 
      n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, 
      n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, 
      n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, 
      n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, 
      n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, 
      n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, 
      n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, 
      n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, 
      n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, 
      n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, 
      n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, 
      n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, 
      n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, 
      n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, 
      n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, 
      n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, 
      n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, 
      n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, 
      n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, 
      n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, 
      n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, 
      n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015, 
      n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, 
      n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, 
      n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, 
      n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, 
      n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, 
      n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, 
      n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, 
      n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087, 
      n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, 
      n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, 
      n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114, 
      n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123, 
      n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132, 
      n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141, 
      n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150, 
      n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159, 
      n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168, 
      n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, 
      n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186, 
      n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195, 
      n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204, 
      n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, 
      n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, 
      n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, 
      n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240, 
      n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249, 
      n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, 
      n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267, 
      n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276, 
      n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, 
      n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294, 
      n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, 
      n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312, 
      n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321, 
      n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330, 
      n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339, 
      n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, 
      n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, 
      n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366, 
      n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375, 
      n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384, 
      n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393, 
      n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402, 
      n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411, 
      n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420, 
      n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, 
      n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438, 
      n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447, 
      n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, 
      n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, 
      n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, 
      n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, 
      n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, 
      n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, 
      n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, 
      n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, 
      n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, 
      n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, 
      n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, 
      n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554 : 
      std_logic;

begin
   
   U15 : NOR2_X1 port map( A1 => n7009, A2 => n696, ZN => n3273);
   U67 : NAND2_X1 port map( A1 => n21574, A2 => n4623, ZN => n203);
   U72 : NOR2_X1 port map( A1 => n20736, A2 => n20739, ZN => n15714);
   U77 : INV_X1 port map( I => n21499, ZN => n21464);
   U82 : INV_X1 port map( I => n79, ZN => n78);
   U107 : INV_X2 port map( I => n13424, ZN => n15378);
   U150 : INV_X1 port map( I => n21141, ZN => n402);
   U184 : NAND2_X1 port map( A1 => n10602, A2 => n11052, ZN => n19982);
   U189 : NAND3_X1 port map( A1 => n8300, A2 => n26738, A3 => n21772, ZN => 
                           n19996);
   U234 : OR2_X1 port map( A1 => n9644, A2 => n7767, Z => n10742);
   U251 : NAND2_X1 port map( A1 => n19608, A2 => n211, ZN => n210);
   U291 : NAND2_X1 port map( A1 => n10881, A2 => n814, ZN => n9840);
   U351 : INV_X1 port map( I => n25376, ZN => n1142);
   U353 : INV_X1 port map( I => n21453, ZN => n1286);
   U369 : INV_X1 port map( I => n20381, ZN => n20603);
   U378 : NAND3_X1 port map( A1 => n10159, A2 => n14378, A3 => n23835, ZN => 
                           n4447);
   U386 : INV_X1 port map( I => n7568, ZN => n14837);
   U392 : NAND2_X1 port map( A1 => n11981, A2 => n21776, ZN => n15516);
   U423 : NOR2_X1 port map( A1 => n9050, A2 => n11485, ZN => n13347);
   U472 : INV_X1 port map( I => n5881, ZN => n266);
   U479 : NOR2_X1 port map( A1 => n24523, A2 => n41, ZN => n10649);
   U535 : NOR2_X1 port map( A1 => n1001, A2 => n26639, ZN => n18768);
   U560 : NOR2_X1 port map( A1 => n2192, A2 => n18612, ZN => n2191);
   U569 : INV_X1 port map( I => n20694, ZN => n918);
   U574 : INV_X2 port map( I => n24363, ZN => n1192);
   U575 : INV_X2 port map( I => n13851, ZN => n13686);
   U585 : INV_X1 port map( I => n14203, ZN => n7150);
   U606 : OAI21_X1 port map( A1 => n506, A2 => n3621, B => n505, ZN => n17836);
   U621 : NOR2_X1 port map( A1 => n890, A2 => n4486, ZN => n506);
   U690 : OAI21_X1 port map( A1 => n7912, A2 => n12225, B => n900, ZN => n4843)
                           ;
   U699 : NOR2_X1 port map( A1 => n17564, A2 => n10539, ZN => n17338);
   U719 : INV_X1 port map( I => n17183, ZN => n17564);
   U730 : OR2_X1 port map( A1 => n17493, A2 => n8125, Z => n8750);
   U805 : OAI21_X1 port map( A1 => n10153, A2 => n10154, B => n10027, ZN => 
                           n9542);
   U821 : AND2_X1 port map( A1 => n162, A2 => n12224, Z => n4761);
   U827 : NAND2_X1 port map( A1 => n15490, A2 => n22061, ZN => n10145);
   U829 : NAND2_X1 port map( A1 => n15029, A2 => n12224, ZN => n9072);
   U840 : INV_X1 port map( I => n16378, ZN => n2300);
   U878 : NOR2_X1 port map( A1 => n3479, A2 => n16466, ZN => n12384);
   U896 : NAND2_X1 port map( A1 => n9828, A2 => n23842, ZN => n9617);
   U913 : NAND2_X1 port map( A1 => n14370, A2 => n15932, ZN => n13334);
   U921 : INV_X1 port map( I => n15943, ZN => n16168);
   U925 : NAND2_X1 port map( A1 => n9986, A2 => n10001, ZN => n15797);
   U931 : INV_X1 port map( I => n333, ZN => n10905);
   U958 : INV_X1 port map( I => n16128, ZN => n14370);
   U978 : AOI22_X2 port map( A1 => n7429, A2 => n7759, B1 => n16503, B2 => 
                           n26835, ZN => n5326);
   U1009 : AOI21_X2 port map( A1 => n17476, A2 => n1035, B => n14275, ZN => 
                           n14274);
   U1014 : AOI21_X2 port map( A1 => n10565, A2 => n987, B => n10348, ZN => 
                           n15101);
   U1068 : INV_X2 port map( I => n14137, ZN => n16632);
   U1080 : BUF_X2 port map( I => n17293, Z => n14367);
   U1086 : NAND2_X2 port map( A1 => n1011, A2 => n1440, ZN => n2564);
   U1091 : INV_X4 port map( I => n4928, ZN => n20430);
   U1109 : NAND2_X1 port map( A1 => n11571, A2 => n11763, ZN => n217);
   U1111 : NOR2_X2 port map( A1 => n9831, A2 => n14267, ZN => n9828);
   U1112 : NAND2_X1 port map( A1 => n4721, A2 => n4754, ZN => n4720);
   U1116 : NOR2_X2 port map( A1 => n4787, A2 => n4786, ZN => n4702);
   U1121 : OAI21_X2 port map( A1 => n14777, A2 => n17826, B => n8502, ZN => 
                           n8501);
   U1134 : AND2_X1 port map( A1 => n4639, A2 => n5434, Z => n8881);
   U1141 : NAND2_X2 port map( A1 => n1362, A2 => n2111, ZN => n3768);
   U1179 : NAND3_X2 port map( A1 => n17720, A2 => n11411, A3 => n28495, ZN => 
                           n6982);
   U1210 : NAND2_X2 port map( A1 => n26730, A2 => n10028, ZN => n10435);
   U1214 : OR2_X1 port map( A1 => n11597, A2 => n11598, Z => n10194);
   U1216 : INV_X2 port map( I => n11775, ZN => n14766);
   U1241 : NOR2_X2 port map( A1 => n11776, A2 => n22201, ZN => n11598);
   U1275 : OAI21_X2 port map( A1 => n4788, A2 => n16484, B => n14264, ZN => 
                           n7855);
   U1278 : INV_X1 port map( I => n13344, ZN => n5327);
   U1282 : NOR2_X1 port map( A1 => n24563, A2 => n17580, ZN => n5478);
   U1287 : INV_X1 port map( I => n13628, ZN => n850);
   U1290 : INV_X1 port map( I => n11395, ZN => n13435);
   U1320 : OAI21_X1 port map( A1 => n28136, A2 => n14664, B => n24062, ZN => 
                           n4409);
   U1323 : NAND2_X1 port map( A1 => n5726, A2 => n20881, ZN => n8030);
   U1325 : OAI22_X2 port map( A1 => n7730, A2 => n6856, B1 => n18470, B2 => 
                           n15693, ZN => n12047);
   U1339 : INV_X1 port map( I => n21638, ZN => n932);
   U1355 : INV_X1 port map( I => n18578, ZN => n1326);
   U1359 : OAI21_X1 port map( A1 => n2939, A2 => n20697, B => n25329, ZN => 
                           n2938);
   U1361 : NOR2_X1 port map( A1 => n22763, A2 => n20608, ZN => n8536);
   U1371 : OAI21_X1 port map( A1 => n25298, A2 => n28314, B => n944, ZN => 
                           n1851);
   U1380 : INV_X1 port map( I => n7184, ZN => n305);
   U1387 : NAND2_X1 port map( A1 => n25214, A2 => n21768, ZN => n15509);
   U1416 : INV_X1 port map( I => n26058, ZN => n14);
   U1421 : NAND2_X1 port map( A1 => n3621, A2 => n17349, ZN => n505);
   U1436 : OAI21_X2 port map( A1 => n6254, A2 => n6253, B => n26652, ZN => 
                           n4155);
   U1437 : INV_X1 port map( I => n21394, ZN => n21405);
   U1444 : NOR2_X1 port map( A1 => n2097, A2 => n305, ZN => n692);
   U1494 : NAND2_X1 port map( A1 => n10217, A2 => n9494, ZN => n8892);
   U1525 : NAND3_X1 port map( A1 => n12290, A2 => n21723, A3 => n21724, ZN => 
                           n6336);
   U1526 : INV_X1 port map( I => n16165, ZN => n11291);
   U1534 : NOR2_X1 port map( A1 => n13538, A2 => n24523, ZN => n532);
   U1535 : NAND2_X1 port map( A1 => n10289, A2 => n13538, ZN => n41);
   U1560 : NAND2_X1 port map( A1 => n7162, A2 => n12510, ZN => n15855);
   U1571 : INV_X1 port map( I => n5420, ZN => n1136);
   U1579 : NAND2_X1 port map( A1 => n21880, A2 => n20963, ZN => n4082);
   U1580 : NOR2_X1 port map( A1 => n20964, A2 => n20963, ZN => n20944);
   U1589 : NAND2_X1 port map( A1 => n14319, A2 => n4246, ZN => n4120);
   U1591 : OAI21_X1 port map( A1 => n19831, A2 => n14319, B => n19830, ZN => 
                           n14472);
   U1592 : NAND2_X1 port map( A1 => n20732, A2 => n27416, ZN => n79);
   U1604 : NAND2_X2 port map( A1 => n1794, A2 => n1795, ZN => n16610);
   U1616 : INV_X2 port map( I => n5680, ZN => n1058);
   U1623 : NOR2_X1 port map( A1 => n26652, A2 => n5577, ZN => n5);
   U1652 : XNOR2_X1 port map( A1 => n17140, A2 => n4807, ZN => n61);
   U1661 : XOR2_X1 port map( A1 => Plaintext(8), A2 => Key(8), Z => n333);
   U1670 : NAND2_X2 port map( A1 => n8102, A2 => n7531, ZN => n16246);
   U1696 : BUF_X4 port map( I => n1869, Z => n1780);
   U1718 : XOR2_X1 port map( A1 => n12222, A2 => n4837, Z => n12220);
   U1728 : AOI21_X1 port map( A1 => n10666, A2 => n20598, B => n21714, ZN => 
                           n3992);
   U1732 : NAND2_X2 port map( A1 => n3991, A2 => n3994, ZN => n7319);
   U1743 : BUF_X2 port map( I => n19603, Z => n45);
   U1768 : NAND2_X2 port map( A1 => n5165, A2 => n5164, ZN => n391);
   U1773 : INV_X2 port map( I => n2025, ZN => n16744);
   U1775 : BUF_X2 port map( I => n13613, Z => n51);
   U1785 : XOR2_X1 port map( A1 => n18132, A2 => n18081, Z => n12783);
   U1789 : XOR2_X1 port map( A1 => n5406, A2 => n10648, Z => n10519);
   U1790 : OAI21_X2 port map( A1 => n53, A2 => n15496, B => n9889, ZN => n9888)
                           ;
   U1793 : AOI21_X2 port map( A1 => n4079, A2 => n25770, B => n4077, ZN => 
                           n3617);
   U1794 : XOR2_X1 port map( A1 => n56, A2 => n20650, Z => Ciphertext(12));
   U1796 : XOR2_X1 port map( A1 => n57, A2 => n25387, Z => n16889);
   U1808 : BUF_X2 port map( I => n10704, Z => n5421);
   U1814 : AOI21_X2 port map( A1 => n17471, A2 => n17534, B => n15394, ZN => 
                           n15393);
   U1815 : OAI21_X1 port map( A1 => n11379, A2 => n22740, B => n21647, ZN => 
                           n11378);
   U1827 : XOR2_X1 port map( A1 => n4809, A2 => n61, Z => n542);
   U1829 : NAND3_X1 port map( A1 => n14858, A2 => n25873, A3 => n15930, ZN => 
                           n9085);
   U1830 : XOR2_X1 port map( A1 => Plaintext(40), A2 => Key(40), Z => n16141);
   U1836 : NOR2_X2 port map( A1 => n3347, A2 => n17728, ZN => n17594);
   U1852 : NAND2_X1 port map( A1 => n68, A2 => n20263, ZN => n67);
   U1861 : INV_X4 port map( I => n13372, ZN => n882);
   U1882 : NAND2_X1 port map( A1 => n10346, A2 => n19803, ZN => n72);
   U1902 : XOR2_X1 port map( A1 => n10999, A2 => n22818, Z => n8115);
   U1906 : INV_X2 port map( I => n658, ZN => n979);
   U1914 : XOR2_X1 port map( A1 => n17399, A2 => n17398, Z => n18753);
   U1918 : NOR2_X2 port map( A1 => n1485, A2 => n4160, ZN => n1483);
   U1925 : BUF_X4 port map( I => n19901, Z => n815);
   U1930 : OR2_X1 port map( A1 => n421, A2 => n1964, Z => n11070);
   U1937 : XOR2_X1 port map( A1 => n89, A2 => n20707, Z => Ciphertext(28));
   U1941 : XOR2_X1 port map( A1 => n8042, A2 => n8041, Z => n8040);
   U1953 : XOR2_X1 port map( A1 => n19482, A2 => n14652, Z => n19483);
   U1960 : NAND2_X2 port map( A1 => n13782, A2 => n5205, ZN => n16251);
   U1985 : NAND2_X2 port map( A1 => n3415, A2 => n4998, ZN => n16485);
   U1987 : AOI22_X2 port map( A1 => n2635, A2 => n11044, B1 => n2057, B2 => 
                           n2633, ZN => n9417);
   U2013 : XOR2_X1 port map( A1 => n19353, A2 => n19228, Z => n2020);
   U2035 : OAI21_X2 port map( A1 => n5230, A2 => n5860, B => n6031, ZN => n5859
                           );
   U2045 : NAND2_X2 port map( A1 => n1112, A2 => n5931, ZN => n6646);
   U2068 : NOR2_X1 port map( A1 => n3223, A2 => n20279, ZN => n8197);
   U2069 : XOR2_X1 port map( A1 => n2477, A2 => n12156, Z => n2476);
   U2077 : NAND2_X2 port map( A1 => n13421, A2 => n17898, ZN => n17768);
   U2120 : OAI21_X1 port map( A1 => n10124, A2 => n8753, B => n26682, ZN => 
                           n1635);
   U2147 : XOR2_X1 port map( A1 => n19300, A2 => n5105, Z => n2611);
   U2149 : OAI21_X2 port map( A1 => n4282, A2 => n4280, B => n28231, ZN => 
                           n4279);
   U2150 : XOR2_X1 port map( A1 => n17074, A2 => n16756, Z => n4031);
   U2158 : INV_X2 port map( I => n18427, ZN => n738);
   U2164 : XOR2_X1 port map( A1 => n10671, A2 => n7304, Z => n137);
   U2174 : AOI21_X1 port map( A1 => n20940, A2 => n23088, B => n139, ZN => 
                           n20943);
   U2180 : INV_X2 port map( I => n7308, ZN => n14676);
   U2181 : OAI21_X1 port map( A1 => n10936, A2 => n10217, B => n21213, ZN => 
                           n5350);
   U2182 : OAI21_X1 port map( A1 => n15345, A2 => n23578, B => n12784, ZN => 
                           n11767);
   U2183 : NAND2_X1 port map( A1 => n25352, A2 => n10635, ZN => n12075);
   U2190 : AND2_X1 port map( A1 => n19826, A2 => n27606, Z => n278);
   U2197 : XOR2_X1 port map( A1 => n3086, A2 => n24529, Z => n3084);
   U2208 : AOI21_X2 port map( A1 => n11061, A2 => n143, B => n11062, ZN => 
                           n20195);
   U2219 : NAND2_X2 port map( A1 => n1617, A2 => n11112, ZN => n5632);
   U2224 : NOR2_X1 port map( A1 => n150, A2 => n10272, ZN => n149);
   U2230 : INV_X2 port map( I => n6603, ZN => n16289);
   U2239 : XOR2_X1 port map( A1 => n2885, A2 => n153, Z => n2882);
   U2240 : XOR2_X1 port map( A1 => n2884, A2 => n21760, Z => n153);
   U2246 : NAND2_X2 port map( A1 => n13815, A2 => n4462, ZN => n16647);
   U2249 : XOR2_X1 port map( A1 => n16876, A2 => n16877, Z => n155);
   U2268 : NAND2_X2 port map( A1 => n2516, A2 => n25412, ZN => n19022);
   U2271 : XOR2_X1 port map( A1 => n3567, A2 => n7824, Z => n3566);
   U2281 : BUF_X4 port map( I => n18232, Z => n18685);
   U2284 : INV_X2 port map( I => n4762, ZN => n14326);
   U2292 : AOI21_X2 port map( A1 => n12445, A2 => n791, B => n15735, ZN => 
                           n8626);
   U2295 : NAND2_X2 port map( A1 => n11600, A2 => n11599, ZN => n17032);
   U2299 : AOI21_X1 port map( A1 => n11755, A2 => n14787, B => n14786, ZN => 
                           n14785);
   U2324 : INV_X2 port map( I => n167, ZN => n631);
   U2333 : XOR2_X1 port map( A1 => n13808, A2 => n25383, Z => n15016);
   U2335 : XOR2_X1 port map( A1 => n170, A2 => n24255, Z => n1481);
   U2336 : XOR2_X1 port map( A1 => n22207, A2 => n21607, Z => n170);
   U2340 : INV_X4 port map( I => n341, ZN => n11579);
   U2343 : INV_X2 port map( I => n18739, ZN => n18653);
   U2345 : OAI21_X2 port map( A1 => n24648, A2 => n3399, B => n13881, ZN => 
                           n3278);
   U2349 : AOI21_X1 port map( A1 => n175, A2 => n15803, B => n16072, ZN => 
                           n15804);
   U2366 : XOR2_X1 port map( A1 => n9904, A2 => n18174, Z => n7831);
   U2368 : NAND2_X2 port map( A1 => n15855, A2 => n182, ZN => n16813);
   U2369 : AOI22_X2 port map( A1 => n15853, A2 => n16279, B1 => n15852, B2 => 
                           n11291, ZN => n182);
   U2401 : XOR2_X1 port map( A1 => n3598, A2 => n11190, Z => n3597);
   U2405 : AND2_X1 port map( A1 => n6425, A2 => n24368, Z => n198);
   U2409 : INV_X2 port map( I => n205, ZN => n7767);
   U2410 : XOR2_X1 port map( A1 => n14129, A2 => n19223, Z => n205);
   U2417 : XOR2_X1 port map( A1 => n6806, A2 => n502, Z => n20345);
   U2419 : XOR2_X1 port map( A1 => n11025, A2 => n15183, Z => n206);
   U2425 : XOR2_X1 port map( A1 => n10107, A2 => n18209, Z => n18056);
   U2433 : BUF_X2 port map( I => n19160, Z => n209);
   U2434 : NAND2_X1 port map( A1 => n212, A2 => n210, ZN => n19611);
   U2436 : OAI21_X1 port map( A1 => n21837, A2 => n213, B => n10549, ZN => n212
                           );
   U2437 : NOR2_X1 port map( A1 => n19720, A2 => n19898, ZN => n213);
   U2444 : XOR2_X1 port map( A1 => n215, A2 => n11450, Z => n20405);
   U2448 : XOR2_X1 port map( A1 => n2264, A2 => n16583, Z => n10049);
   U2453 : XOR2_X1 port map( A1 => n218, A2 => n16781, Z => n8549);
   U2454 : XOR2_X1 port map( A1 => n8547, A2 => n9614, Z => n218);
   U2467 : XOR2_X1 port map( A1 => n19434, A2 => n19195, Z => n220);
   U2469 : BUF_X2 port map( I => n10401, Z => n8594);
   U2483 : OR2_X1 port map( A1 => n15886, A2 => n15989, Z => n10866);
   U2492 : INV_X4 port map( I => n14815, ZN => n16280);
   U2504 : NAND2_X1 port map( A1 => n16471, A2 => n15029, ZN => n10710);
   U2521 : NAND2_X1 port map( A1 => n2190, A2 => n9249, ZN => n233);
   U2524 : XOR2_X1 port map( A1 => n6582, A2 => n16794, Z => n16796);
   U2554 : NAND2_X2 port map( A1 => n11803, A2 => n7341, ZN => n15524);
   U2556 : BUF_X2 port map( I => n5169, Z => n242);
   U2563 : NAND2_X1 port map( A1 => n576, A2 => n5139, ZN => n9969);
   U2566 : INV_X1 port map( I => n21641, ZN => n803);
   U2572 : XOR2_X1 port map( A1 => n248, A2 => n13643, Z => n13642);
   U2576 : NAND2_X1 port map( A1 => n9996, A2 => n249, ZN => n9999);
   U2577 : OR3_X1 port map( A1 => n14314, A2 => n11152, A3 => n14313, Z => n249
                           );
   U2579 : NAND2_X2 port map( A1 => n17674, A2 => n17675, ZN => n11502);
   U2597 : AOI21_X2 port map( A1 => n9178, A2 => n19948, B => n9176, ZN => 
                           n9175);
   U2616 : XOR2_X1 port map( A1 => n1353, A2 => n2529, Z => n20502);
   U2618 : NAND2_X2 port map( A1 => n7525, A2 => n8620, ZN => n16139);
   U2619 : XOR2_X1 port map( A1 => n256, A2 => n9292, Z => n5226);
   U2620 : XOR2_X1 port map( A1 => n26719, A2 => n257, Z => n256);
   U2623 : AOI22_X2 port map( A1 => n18480, A2 => n18481, B1 => n18723, B2 => 
                           n9163, ZN => n19164);
   U2631 : INV_X2 port map( I => n615, ZN => n831);
   U2650 : NAND2_X2 port map( A1 => n22614, A2 => n15159, ZN => n1802);
   U2655 : NAND2_X2 port map( A1 => n3875, A2 => n7175, ZN => n14862);
   U2664 : NOR2_X1 port map( A1 => n6246, A2 => n6248, ZN => n272);
   U2665 : INV_X4 port map( I => n15886, ZN => n1271);
   U2666 : OAI21_X2 port map( A1 => n7737, A2 => n23889, B => n273, ZN => 
                           n11485);
   U2667 : XOR2_X1 port map( A1 => n274, A2 => n10373, Z => n4025);
   U2671 : XOR2_X1 port map( A1 => n23641, A2 => n14479, Z => n14058);
   U2681 : NAND3_X2 port map( A1 => n8251, A2 => n8253, A3 => n8252, ZN => 
                           n12600);
   U2690 : BUF_X4 port map( I => n11819, Z => n913);
   U2695 : NOR2_X2 port map( A1 => n13275, A2 => n17831, ZN => n18236);
   U2696 : NOR2_X1 port map( A1 => n18776, A2 => n1005, ZN => n281);
   U2700 : INV_X2 port map( I => n14193, ZN => n19805);
   U2705 : NOR2_X1 port map( A1 => n9422, A2 => n21035, ZN => n21036);
   U2712 : AOI21_X1 port map( A1 => n21168, A2 => n27368, B => n936, ZN => 
                           n15657);
   U2726 : NAND3_X1 port map( A1 => n7944, A2 => n13987, A3 => n12784, ZN => 
                           n6466);
   U2728 : NOR2_X2 port map( A1 => n1026, A2 => n14548, ZN => n6415);
   U2747 : NAND2_X1 port map( A1 => n18705, A2 => n25709, ZN => n293);
   U2748 : INV_X1 port map( I => n15405, ZN => n294);
   U2752 : XOR2_X1 port map( A1 => n295, A2 => n4568, Z => n8995);
   U2757 : INV_X2 port map( I => n7183, ZN => n13578);
   U2759 : NAND2_X2 port map( A1 => n22614, A2 => n5861, ZN => n16689);
   U2769 : NAND2_X1 port map( A1 => n7555, A2 => n7554, ZN => n299);
   U2772 : NAND2_X2 port map( A1 => n23540, A2 => n15137, ZN => n18145);
   U2777 : NAND2_X1 port map( A1 => n16049, A2 => n23880, ZN => n301);
   U2783 : XOR2_X1 port map( A1 => n17153, A2 => n303, Z => n302);
   U2792 : XOR2_X1 port map( A1 => n17072, A2 => n11769, Z => n1789);
   U2793 : NAND2_X2 port map( A1 => n1791, A2 => n1790, ZN => n17072);
   U2795 : INV_X4 port map( I => n22614, ZN => n5557);
   U2796 : XOR2_X1 port map( A1 => n4305, A2 => n4304, Z => n4303);
   U2800 : XOR2_X1 port map( A1 => n16779, A2 => n8080, Z => n8079);
   U2806 : OR2_X1 port map( A1 => n17591, A2 => n26610, Z => n2809);
   U2814 : BUF_X2 port map( I => n13727, Z => n309);
   U2815 : NAND2_X2 port map( A1 => n12581, A2 => n10675, ZN => n10992);
   U2817 : NOR2_X2 port map( A1 => n13964, A2 => n13927, ZN => n16399);
   U2818 : XOR2_X1 port map( A1 => n18347, A2 => n311, Z => n18160);
   U2819 : XOR2_X1 port map( A1 => n1193, A2 => n18329, Z => n311);
   U2822 : NOR2_X1 port map( A1 => n10268, A2 => n6756, ZN => n21225);
   U2832 : OR2_X1 port map( A1 => n21446, A2 => n14017, Z => n21178);
   U2841 : XOR2_X1 port map( A1 => n23359, A2 => n567, Z => n316);
   U2843 : NAND2_X2 port map( A1 => n10135, A2 => n10137, ZN => n12439);
   U2862 : XOR2_X1 port map( A1 => n12289, A2 => n21906, Z => n319);
   U2867 : INV_X1 port map( I => n18353, ZN => n13314);
   U2868 : NAND3_X2 port map( A1 => n8219, A2 => n8222, A3 => n8218, ZN => 
                           n18353);
   U2875 : INV_X2 port map( I => n12694, ZN => n729);
   U2878 : NAND2_X2 port map( A1 => n4720, A2 => n16847, ZN => n4719);
   U2880 : NAND2_X2 port map( A1 => n9714, A2 => n10928, ZN => n9494);
   U2890 : OAI21_X2 port map( A1 => n1038, A2 => n14126, B => n892, ZN => n7785
                           );
   U2898 : AND2_X1 port map( A1 => n2478, A2 => n18685, Z => n12385);
   U2912 : NAND2_X1 port map( A1 => n21490, A2 => n21491, ZN => n5186);
   U2933 : XOR2_X1 port map( A1 => Plaintext(26), A2 => Key(26), Z => n338);
   U2935 : INV_X2 port map( I => n12498, ZN => n17502);
   U2939 : NOR2_X2 port map( A1 => n18804, A2 => n18803, ZN => n19324);
   U2947 : XOR2_X1 port map( A1 => n20761, A2 => n13092, Z => n20353);
   U2952 : INV_X2 port map( I => n28551, ZN => n4308);
   U2972 : XOR2_X1 port map( A1 => n10248, A2 => n21239, Z => n4965);
   U2980 : AOI21_X2 port map( A1 => n19844, A2 => n19876, B => n19842, ZN => 
                           n19737);
   U3027 : XOR2_X1 port map( A1 => n5420, A2 => n14360, Z => n6025);
   U3037 : OAI21_X2 port map( A1 => n17499, A2 => n9018, B => n17497, ZN => 
                           n8609);
   U3040 : OR2_X1 port map( A1 => n10045, A2 => n10937, Z => n359);
   U3046 : XOR2_X1 port map( A1 => n15851, A2 => Key(114), Z => n1321);
   U3049 : NAND2_X1 port map( A1 => n4821, A2 => n14146, ZN => n8586);
   U3054 : XOR2_X1 port map( A1 => n4133, A2 => n24520, Z => n1550);
   U3055 : NAND2_X2 port map( A1 => n9250, A2 => n8432, ZN => n1587);
   U3071 : AOI21_X2 port map( A1 => n1491, A2 => n8621, B => n3928, ZN => 
                           n12267);
   U3073 : INV_X2 port map( I => n10251, ZN => n10545);
   U3086 : OAI21_X2 port map( A1 => n13335, A2 => n14370, B => n13334, ZN => 
                           n16698);
   U3090 : XOR2_X1 port map( A1 => n12411, A2 => n6809, Z => n21301);
   U3096 : XOR2_X1 port map( A1 => n19331, A2 => n369, Z => n599);
   U3097 : XOR2_X1 port map( A1 => n370, A2 => n19330, Z => n369);
   U3103 : NAND2_X1 port map( A1 => n25324, A2 => n28176, ZN => n12519);
   U3126 : XOR2_X1 port map( A1 => n383, A2 => n8194, Z => n6229);
   U3141 : XOR2_X1 port map( A1 => n13537, A2 => n19414, Z => n5930);
   U3149 : INV_X4 port map( I => n18645, ZN => n10872);
   U3173 : NAND2_X2 port map( A1 => n5959, A2 => n5958, ZN => n5955);
   U3178 : AOI21_X2 port map( A1 => n14452, A2 => n21787, B => n10740, ZN => 
                           n7144);
   U3182 : AOI22_X2 port map( A1 => n15953, A2 => n840, B1 => n2719, B2 => 
                           n1261, ZN => n2590);
   U3187 : NAND2_X2 port map( A1 => n13964, A2 => n16530, ZN => n16400);
   U3188 : INV_X2 port map( I => n13888, ZN => n847);
   U3195 : XOR2_X1 port map( A1 => n8726, A2 => n402, Z => n6059);
   U3202 : INV_X4 port map( I => n14671, ZN => n19758);
   U3205 : XOR2_X1 port map( A1 => n406, A2 => n21281, Z => Ciphertext(115));
   U3206 : AOI22_X1 port map( A1 => n21293, A2 => n11891, B1 => n21284, B2 => 
                           n21280, ZN => n406);
   U3209 : AOI21_X1 port map( A1 => n21477, A2 => n22844, B => n407, ZN => 
                           n10834);
   U3212 : XOR2_X1 port map( A1 => n2994, A2 => n10294, Z => n17063);
   U3225 : NAND2_X2 port map( A1 => n11423, A2 => n8620, ZN => n16138);
   U3245 : NOR2_X2 port map( A1 => n8513, A2 => n3423, ZN => n1879);
   U3246 : AND2_X1 port map( A1 => n8536, A2 => n25315, Z => n693);
   U3255 : NAND2_X1 port map( A1 => n7571, A2 => n21774, ZN => n17241);
   U3259 : XOR2_X1 port map( A1 => n20513, A2 => n21196, Z => n14678);
   U3260 : XOR2_X1 port map( A1 => n20538, A2 => n11885, Z => n21196);
   U3263 : XOR2_X1 port map( A1 => n6932, A2 => n2290, Z => n1946);
   U3285 : NAND2_X2 port map( A1 => n16137, A2 => n10457, ZN => n16728);
   U3286 : NAND2_X2 port map( A1 => n20930, A2 => n20929, ZN => n20963);
   U3288 : NAND2_X1 port map( A1 => n13086, A2 => n20623, ZN => n13085);
   U3293 : NAND2_X1 port map( A1 => n7700, A2 => n26198, ZN => n7003);
   U3296 : OAI21_X2 port map( A1 => n26693, A2 => n422, B => n14651, ZN => 
                           n3100);
   U3306 : INV_X2 port map( I => n13101, ZN => n15038);
   U3308 : NAND2_X2 port map( A1 => n9797, A2 => n9800, ZN => n13101);
   U3320 : AOI21_X2 port map( A1 => n24634, A2 => n18509, B => n6712, ZN => 
                           n7478);
   U3323 : NAND2_X2 port map( A1 => n9772, A2 => n4455, ZN => n7986);
   U3332 : NOR2_X1 port map( A1 => n7472, A2 => n16234, ZN => n10696);
   U3338 : XOR2_X1 port map( A1 => n437, A2 => n21411, Z => Ciphertext(130));
   U3343 : OAI21_X2 port map( A1 => n5939, A2 => n10583, B => n5938, ZN => 
                           n17914);
   U3347 : NOR2_X2 port map( A1 => n15744, A2 => n13396, ZN => n7086);
   U3351 : NAND3_X1 port map( A1 => n22775, A2 => n27443, A3 => n12617, ZN => 
                           n19699);
   U3367 : XOR2_X1 port map( A1 => n442, A2 => n26082, Z => n1859);
   U3387 : INV_X2 port map( I => n14321, ZN => n12711);
   U3389 : NAND2_X2 port map( A1 => n2976, A2 => n3479, ZN => n4166);
   U3399 : AOI22_X2 port map( A1 => n6655, A2 => n19619, B1 => n12425, B2 => 
                           n7849, ZN => n5415);
   U3431 : XOR2_X1 port map( A1 => n8366, A2 => n21570, Z => n6960);
   U3433 : AOI22_X1 port map( A1 => n456, A2 => n12270, B1 => n12904, B2 => 
                           n28308, ZN => n12903);
   U3434 : NAND2_X1 port map( A1 => n21567, A2 => n22789, ZN => n456);
   U3438 : INV_X2 port map( I => n19559, ZN => n19387);
   U3439 : NAND3_X2 port map( A1 => n3012, A2 => n3010, A3 => n3015, ZN => 
                           n19559);
   U3462 : BUF_X2 port map( I => n13538, Z => n467);
   U3468 : NAND2_X2 port map( A1 => n21623, A2 => n11198, ZN => n21546);
   U3473 : NOR3_X2 port map( A1 => n16555, A2 => n4630, A3 => n23505, ZN => 
                           n16368);
   U3476 : BUF_X4 port map( I => n10134, Z => n9675);
   U3480 : OAI21_X2 port map( A1 => n28461, A2 => n12875, B => n8867, ZN => 
                           n8826);
   U3484 : XOR2_X1 port map( A1 => n1622, A2 => n10736, Z => n473);
   U3490 : XOR2_X1 port map( A1 => n6864, A2 => n20148, Z => n1534);
   U3505 : XOR2_X1 port map( A1 => n8259, A2 => n14238, Z => n21430);
   U3509 : INV_X2 port map( I => n28551, ZN => n21444);
   U3529 : NAND2_X2 port map( A1 => n6975, A2 => n15098, ZN => n17688);
   U3531 : NOR2_X2 port map( A1 => n16698, A2 => n16697, ZN => n10144);
   U3532 : INV_X2 port map( I => n16103, ZN => n14385);
   U3536 : BUF_X2 port map( I => n15997, Z => n14584);
   U3539 : NAND2_X2 port map( A1 => n5562, A2 => n5566, ZN => n17607);
   U3542 : INV_X2 port map( I => n21729, ZN => n1076);
   U3544 : NAND2_X2 port map( A1 => n17688, A2 => n12815, ZN => n2329);
   U3549 : INV_X4 port map( I => n17487, ZN => n15077);
   U3559 : INV_X2 port map( I => n7281, ZN => n14887);
   U3570 : XOR2_X1 port map( A1 => n6507, A2 => n9505, Z => n7252);
   U3581 : XOR2_X1 port map( A1 => n18327, A2 => n10996, Z => n10995);
   U3583 : XOR2_X1 port map( A1 => n13136, A2 => n9803, Z => n502);
   U3599 : NAND3_X2 port map( A1 => n17341, A2 => n17339, A3 => n17340, ZN => 
                           n2636);
   U3607 : INV_X4 port map( I => n10539, ZN => n17565);
   U3608 : INV_X2 port map( I => n16677, ZN => n6937);
   U3620 : XOR2_X1 port map( A1 => n4889, A2 => n15230, Z => n511);
   U3628 : XOR2_X1 port map( A1 => n517, A2 => n22771, Z => n5490);
   U3632 : INV_X4 port map( I => n13049, ZN => n1084);
   U3637 : OAI21_X2 port map( A1 => n16607, A2 => n16608, B => n16606, ZN => 
                           n2290);
   U3643 : XOR2_X1 port map( A1 => n16863, A2 => n2290, Z => n17086);
   U3663 : NOR3_X1 port map( A1 => n4802, A2 => n12257, A3 => n17950, ZN => 
                           n3124);
   U3677 : NAND2_X1 port map( A1 => n529, A2 => n527, ZN => n13335);
   U3678 : NAND2_X1 port map( A1 => n14512, A2 => n12116, ZN => n529);
   U3681 : NOR2_X2 port map( A1 => n16113, A2 => n3262, ZN => n1908);
   U3683 : INV_X2 port map( I => n11407, ZN => n3773);
   U3684 : XOR2_X1 port map( A1 => n531, A2 => n18209, Z => n13364);
   U3686 : AOI22_X2 port map( A1 => n11359, A2 => n17759, B1 => n26681, B2 => 
                           n17954, ZN => n18209);
   U3719 : NAND2_X1 port map( A1 => n2394, A2 => n2177, ZN => n2396);
   U3729 : NOR2_X1 port map( A1 => n8824, A2 => n19861, ZN => n19575);
   U3741 : AND2_X1 port map( A1 => n21699, A2 => n21724, Z => n689);
   U3747 : INV_X1 port map( I => n21199, ZN => n1305);
   U3748 : INV_X1 port map( I => n14576, ZN => n1303);
   U3750 : XNOR2_X1 port map( A1 => n10773, A2 => n21476, ZN => n535);
   U3751 : XNOR2_X1 port map( A1 => n16960, A2 => n16962, ZN => n536);
   U3754 : XNOR2_X1 port map( A1 => n21895, A2 => n14016, ZN => n539);
   U3757 : XNOR2_X1 port map( A1 => n14143, A2 => n584, ZN => n543);
   U3758 : XNOR2_X1 port map( A1 => n8819, A2 => n14558, ZN => n544);
   U3759 : XNOR2_X1 port map( A1 => n2850, A2 => n1279, ZN => n545);
   U3760 : XNOR2_X1 port map( A1 => n11684, A2 => n21077, ZN => n546);
   U3763 : XNOR2_X1 port map( A1 => n19478, A2 => n20872, ZN => n549);
   U3764 : XNOR2_X1 port map( A1 => n27448, A2 => n21523, ZN => n550);
   U3767 : XNOR2_X1 port map( A1 => n17754, A2 => n10544, ZN => n553);
   U3768 : XOR2_X1 port map( A1 => n16937, A2 => n14418, Z => n554);
   U3770 : XNOR2_X1 port map( A1 => n20449, A2 => n21732, ZN => n556);
   U3772 : XNOR2_X1 port map( A1 => n19330, A2 => n14404, ZN => n558);
   U3773 : XNOR2_X1 port map( A1 => n9534, A2 => n14560, ZN => n559);
   U3774 : XNOR2_X1 port map( A1 => n13469, A2 => n14488, ZN => n560);
   U3775 : XOR2_X1 port map( A1 => Key(89), A2 => Plaintext(89), Z => n561);
   U3777 : XOR2_X1 port map( A1 => Plaintext(168), A2 => Key(168), Z => n563);
   U3779 : XOR2_X1 port map( A1 => n1801, A2 => Plaintext(19), Z => n564);
   U3781 : XNOR2_X1 port map( A1 => n15708, A2 => n13678, ZN => n566);
   U3782 : XNOR2_X1 port map( A1 => n18161, A2 => n20877, ZN => n567);
   U3786 : INV_X2 port map( I => n13757, ZN => n19015);
   U3790 : XOR2_X1 port map( A1 => Plaintext(102), A2 => Key(102), Z => n573);
   U3796 : XNOR2_X1 port map( A1 => n16502, A2 => n16501, ZN => n578);
   U3798 : XNOR2_X1 port map( A1 => n18130, A2 => n1278, ZN => n580);
   U3801 : XNOR2_X1 port map( A1 => n12204, A2 => n20208, ZN => n584);
   U3804 : XNOR2_X1 port map( A1 => n8657, A2 => n19500, ZN => n587);
   U3808 : XNOR2_X1 port map( A1 => n18161, A2 => n18360, ZN => n590);
   U3810 : XNOR2_X1 port map( A1 => n14187, A2 => n1305, ZN => n592);
   U3812 : XNOR2_X1 port map( A1 => n24318, A2 => n26793, ZN => n594);
   U3813 : XNOR2_X1 port map( A1 => n19527, A2 => n10544, ZN => n595);
   U3814 : XNOR2_X1 port map( A1 => n19445, A2 => n14503, ZN => n596);
   U3815 : XNOR2_X1 port map( A1 => n19445, A2 => n19391, ZN => n597);
   U3819 : XNOR2_X1 port map( A1 => n22135, A2 => n14623, ZN => n602);
   U3820 : XNOR2_X1 port map( A1 => n5351, A2 => n21419, ZN => n603);
   U3821 : XNOR2_X1 port map( A1 => n6562, A2 => n14550, ZN => n604);
   U3823 : XNOR2_X1 port map( A1 => n19334, A2 => n21044, ZN => n605);
   U3825 : XNOR2_X1 port map( A1 => n19306, A2 => n14540, ZN => n608);
   U3826 : XNOR2_X1 port map( A1 => n11389, A2 => n21190, ZN => n609);
   U3828 : XNOR2_X1 port map( A1 => n19487, A2 => n14591, ZN => n610);
   U3829 : XNOR2_X1 port map( A1 => n19532, A2 => n20683, ZN => n611);
   U3839 : INV_X2 port map( I => n10431, ZN => n9593);
   U3844 : XOR2_X1 port map( A1 => n1548, A2 => n1890, Z => n619);
   U3850 : XOR2_X1 port map( A1 => n9006, A2 => n9007, Z => n624);
   U3851 : AND2_X1 port map( A1 => n23863, A2 => n28389, Z => n625);
   U3853 : XNOR2_X1 port map( A1 => n6705, A2 => n6704, ZN => n626);
   U3856 : AND2_X1 port map( A1 => n9675, A2 => n10816, Z => n628);
   U3857 : INV_X2 port map( I => n14426, ZN => n2963);
   U3866 : XNOR2_X1 port map( A1 => n27137, A2 => n14480, ZN => n634);
   U3872 : XNOR2_X1 port map( A1 => n18168, A2 => n10853, ZN => n637);
   U3875 : XOR2_X1 port map( A1 => n22165, A2 => n21281, Z => n639);
   U3876 : XNOR2_X1 port map( A1 => n1019, A2 => n1454, ZN => n641);
   U3877 : XNOR2_X1 port map( A1 => n18162, A2 => n10734, ZN => n642);
   U3879 : XNOR2_X1 port map( A1 => n4580, A2 => n18021, ZN => n644);
   U3892 : INV_X2 port map( I => n27797, ZN => n18475);
   U3896 : INV_X2 port map( I => n15674, ZN => n15693);
   U3897 : NOR2_X2 port map( A1 => n12579, A2 => n15133, ZN => n18794);
   U3904 : XNOR2_X1 port map( A1 => n4777, A2 => n27451, ZN => n653);
   U3915 : XNOR2_X1 port map( A1 => n14570, A2 => n9545, ZN => n655);
   U3917 : XNOR2_X1 port map( A1 => n22810, A2 => n11995, ZN => n657);
   U3918 : XOR2_X1 port map( A1 => n19496, A2 => n19495, Z => n659);
   U3925 : INV_X2 port map( I => n7240, ZN => n8330);
   U3926 : XOR2_X1 port map( A1 => n8337, A2 => n8338, Z => n666);
   U3929 : XNOR2_X1 port map( A1 => n11245, A2 => n11244, ZN => n668);
   U3930 : INV_X2 port map( I => n7854, ZN => n11369);
   U3935 : XNOR2_X1 port map( A1 => n11551, A2 => n6200, ZN => n672);
   U3954 : XOR2_X1 port map( A1 => n14144, A2 => n20034, Z => n682);
   U3955 : XNOR2_X1 port map( A1 => n9859, A2 => n9858, ZN => n684);
   U3957 : XNOR2_X1 port map( A1 => n20450, A2 => n14600, ZN => n686);
   U3965 : INV_X2 port map( I => n14795, ZN => n21161);
   U3974 : NOR2_X2 port map( A1 => n15986, A2 => n15983, ZN => n16016);
   U3978 : INV_X2 port map( I => n19661, ZN => n19782);
   U3995 : NOR2_X2 port map( A1 => n8931, A2 => n8929, ZN => n8928);
   U4011 : NOR3_X2 port map( A1 => n7722, A2 => n7721, A3 => n16339, ZN => 
                           n7720);
   U4019 : NAND2_X1 port map( A1 => n19140, A2 => n2398, ZN => n1848);
   U4026 : INV_X2 port map( I => n14385, ZN => n7266);
   U4048 : AOI21_X2 port map( A1 => n19824, A2 => n14752, B => n13911, ZN => 
                           n14751);
   U4052 : AND2_X2 port map( A1 => n15545, A2 => n21054, Z => n21098);
   U4058 : NAND2_X2 port map( A1 => n14887, A2 => n13721, ZN => n14894);
   U4059 : NAND2_X2 port map( A1 => n25415, A2 => n16336, ZN => n16660);
   U4075 : OAI21_X2 port map( A1 => n16497, A2 => n14483, B => n14894, ZN => 
                           n15301);
   U4088 : NAND2_X2 port map( A1 => n9273, A2 => n9270, ZN => n18891);
   U4095 : AOI22_X2 port map( A1 => n683, A2 => n9103, B1 => n1102, B2 => 
                           n24394, ZN => n9955);
   U4098 : INV_X2 port map( I => n9618, ZN => n10555);
   U4127 : INV_X1 port map( I => n16306, ZN => n11407);
   U4134 : NOR2_X2 port map( A1 => n8573, A2 => n12379, ZN => n14162);
   U4170 : INV_X4 port map( I => n8939, ZN => n17941);
   U4176 : NAND2_X1 port map( A1 => n21405, A2 => n13741, ZN => n4984);
   U4177 : NOR2_X1 port map( A1 => n21409, A2 => n22794, ZN => n5004);
   U4193 : NAND2_X1 port map( A1 => n1074, A2 => n21500, ZN => n4514);
   U4207 : INV_X1 port map( I => n13188, ZN => n20635);
   U4216 : INV_X2 port map( I => n14567, ZN => n21629);
   U4217 : INV_X1 port map( I => n3353, ZN => n20921);
   U4223 : INV_X1 port map( I => n13684, ZN => n1098);
   U4233 : INV_X1 port map( I => n23253, ZN => n709);
   U4253 : INV_X2 port map( I => n7186, ZN => n9583);
   U4275 : INV_X1 port map( I => n14138, ZN => n785);
   U4281 : NOR2_X2 port map( A1 => n8613, A2 => n8612, ZN => n18221);
   U4284 : NAND3_X1 port map( A1 => n6910, A2 => n17676, A3 => n9330, ZN => 
                           n4458);
   U4286 : INV_X1 port map( I => n27947, ZN => n6109);
   U4293 : NAND3_X2 port map( A1 => n3625, A2 => n3623, A3 => n3622, ZN => 
                           n13043);
   U4298 : NAND3_X1 port map( A1 => n17036, A2 => n17415, A3 => n14250, ZN => 
                           n10903);
   U4300 : INV_X1 port map( I => n11610, ZN => n8094);
   U4310 : NAND2_X1 port map( A1 => n16512, A2 => n16657, ZN => n10988);
   U4326 : NOR2_X1 port map( A1 => n16220, A2 => n16255, ZN => n7229);
   U4327 : OAI21_X1 port map( A1 => n16256, A2 => n16253, B => n16220, ZN => 
                           n16446);
   U4328 : INV_X1 port map( I => n15188, ZN => n1056);
   U4336 : INV_X2 port map( I => n14425, ZN => n16111);
   U4352 : NAND3_X1 port map( A1 => n4057, A2 => n4428, A3 => n21116, ZN => 
                           n4430);
   U4376 : INV_X2 port map( I => n15374, ZN => n722);
   U4381 : INV_X1 port map( I => n14601, ZN => n1092);
   U4394 : INV_X1 port map( I => n7289, ZN => n15320);
   U4416 : NAND2_X1 port map( A1 => n867, A2 => n204, ZN => n19096);
   U4440 : INV_X1 port map( I => n24525, ZN => n18781);
   U4465 : OAI21_X2 port map( A1 => n12194, A2 => n12193, B => n8379, ZN => 
                           n9772);
   U4469 : OAI21_X2 port map( A1 => n17568, A2 => n17567, B => n17566, ZN => 
                           n17578);
   U4472 : NAND2_X2 port map( A1 => n16880, A2 => n16879, ZN => n17989);
   U4499 : OAI21_X2 port map( A1 => n7631, A2 => n16313, B => n16312, ZN => 
                           n7596);
   U4500 : NAND3_X1 port map( A1 => n26879, A2 => n1419, A3 => n1056, ZN => 
                           n2281);
   U4511 : BUF_X1 port map( I => Key(78), Z => n21742);
   U4518 : INV_X1 port map( I => n2588, ZN => n15742);
   U4527 : INV_X1 port map( I => n20755, ZN => n8232);
   U4536 : INV_X1 port map( I => n21671, ZN => n4879);
   U4547 : NAND2_X1 port map( A1 => n20493, A2 => n1731, ZN => n14054);
   U4559 : OAI21_X1 port map( A1 => n21788, A2 => n7182, B => n8562, ZN => 
                           n5295);
   U4573 : INV_X2 port map( I => n7025, ZN => n11175);
   U4577 : INV_X1 port map( I => n19593, ZN => n1128);
   U4578 : INV_X2 port map( I => n6166, ZN => n735);
   U4579 : INV_X1 port map( I => n8704, ZN => n11708);
   U4597 : INV_X1 port map( I => n7770, ZN => n14245);
   U4603 : INV_X4 port map( I => n11426, ZN => n737);
   U4604 : INV_X1 port map( I => n11809, ZN => n14138);
   U4608 : AOI21_X1 port map( A1 => n17952, A2 => n28495, B => n786, ZN => 
                           n5765);
   U4623 : INV_X1 port map( I => n17247, ZN => n8108);
   U4639 : BUF_X2 port map( I => n17469, Z => n748);
   U4641 : NAND3_X1 port map( A1 => n9072, A2 => n16553, A3 => n162, ZN => 
                           n6495);
   U4653 : INV_X1 port map( I => n16343, ZN => n9526);
   U4657 : BUF_X2 port map( I => n16343, Z => n14644);
   U4660 : BUF_X1 port map( I => Key(140), Z => n19218);
   U4663 : NAND2_X1 port map( A1 => n21644, A2 => n21636, ZN => n21646);
   U4664 : INV_X1 port map( I => n21608, ZN => n21604);
   U4676 : NAND2_X1 port map( A1 => n11198, A2 => n21626, ZN => n11251);
   U4684 : NAND2_X1 port map( A1 => n8246, A2 => n10610, ZN => n20755);
   U4705 : NAND2_X1 port map( A1 => n4393, A2 => n14256, ZN => n7060);
   U4723 : NAND3_X1 port map( A1 => n6394, A2 => n24579, A3 => n1120, ZN => 
                           n19943);
   U4728 : NAND2_X1 port map( A1 => n28377, A2 => n19823, ZN => n3190);
   U4729 : AND2_X1 port map( A1 => n19642, A2 => n19918, Z => n2652);
   U4747 : NOR2_X1 port map( A1 => n24454, A2 => n23488, ZN => n4453);
   U4751 : NOR2_X1 port map( A1 => n114, A2 => n18891, ZN => n18984);
   U4754 : INV_X1 port map( I => n24190, ZN => n18925);
   U4759 : INV_X1 port map( I => n18768, ZN => n5582);
   U4762 : NAND2_X1 port map( A1 => n22873, A2 => n18366, ZN => n10672);
   U4770 : OR2_X1 port map( A1 => n18785, A2 => n2072, Z => n3202);
   U4771 : AND2_X1 port map( A1 => n8576, A2 => n26639, Z => n11416);
   U4772 : INV_X1 port map( I => n18609, ZN => n18698);
   U4783 : AOI21_X1 port map( A1 => n11410, A2 => n788, B => n3124, ZN => 
                           n11409);
   U4809 : NAND2_X2 port map( A1 => n7405, A2 => n9990, ZN => n6770);
   U4823 : NOR2_X1 port map( A1 => n26298, A2 => n6937, ZN => n6933);
   U4825 : NAND3_X1 port map( A1 => n742, A2 => n23096, A3 => n741, ZN => n9110
                           );
   U4848 : INV_X1 port map( I => n16342, ZN => n16115);
   U4849 : INV_X1 port map( I => n16190, ZN => n7022);
   U4875 : INV_X4 port map( I => n7587, ZN => n20932);
   U4890 : NAND2_X1 port map( A1 => n14179, A2 => n9446, ZN => n20162);
   U4895 : NAND3_X1 port map( A1 => n9994, A2 => n13771, A3 => n964, ZN => 
                           n6665);
   U4897 : NOR2_X1 port map( A1 => n20339, A2 => n7618, ZN => n9961);
   U4918 : NAND2_X1 port map( A1 => n13665, A2 => n19744, ZN => n19765);
   U4922 : INV_X2 port map( I => n14757, ZN => n756);
   U4930 : NOR2_X1 port map( A1 => n10474, A2 => n19140, ZN => n10265);
   U4937 : OR2_X1 port map( A1 => n11576, A2 => n10362, Z => n4001);
   U4953 : NAND2_X1 port map( A1 => n18566, A2 => n14498, ZN => n18567);
   U4959 : INV_X2 port map( I => n2013, ZN => n758);
   U4970 : INV_X1 port map( I => n18725, ZN => n18667);
   U4979 : INV_X2 port map( I => n12094, ZN => n761);
   U5002 : NAND3_X1 port map( A1 => n10566, A2 => n10920, A3 => n17843, ZN => 
                           n17752);
   U5005 : NAND2_X1 port map( A1 => n622, A2 => n28367, ZN => n16847);
   U5020 : AOI21_X1 port map( A1 => n6462, A2 => n28539, B => n748, ZN => n6460
                           );
   U5024 : INV_X1 port map( I => n12450, ZN => n6112);
   U5037 : INV_X2 port map( I => n10190, ZN => n767);
   U5045 : NAND2_X1 port map( A1 => n16514, A2 => n27353, ZN => n16760);
   U5048 : AND2_X1 port map( A1 => n5310, A2 => n23935, Z => n1992);
   U5058 : NOR3_X1 port map( A1 => n14198, A2 => n14197, A3 => n16195, ZN => 
                           n8762);
   U5068 : NAND2_X1 port map( A1 => n16351, A2 => n16086, ZN => n6844);
   U5076 : NAND2_X1 port map( A1 => n21876, A2 => n16342, ZN => n16341);
   U5077 : NOR2_X1 port map( A1 => n7608, A2 => n10303, ZN => n16353);
   U5079 : BUF_X2 port map( I => n16165, Z => n16278);
   U5082 : INV_X1 port map( I => n9437, ZN => n8925);
   U5092 : AND2_X1 port map( A1 => n25329, A2 => n8388, Z => n2115);
   U5117 : INV_X2 port map( I => n15642, ZN => n773);
   U5118 : BUF_X2 port map( I => n5914, Z => n5904);
   U5125 : NOR2_X1 port map( A1 => n7978, A2 => n20253, ZN => n7062);
   U5129 : CLKBUF_X2 port map( I => n20339, Z => n11920);
   U5130 : INV_X1 port map( I => n20336, ZN => n960);
   U5139 : NAND2_X1 port map( A1 => n19760, A2 => n1122, ZN => n19964);
   U5151 : NAND2_X1 port map( A1 => n19935, A2 => n814, ZN => n12738);
   U5170 : INV_X4 port map( I => n14459, ZN => n867);
   U5176 : INV_X2 port map( I => n14423, ZN => n777);
   U5194 : INV_X1 port map( I => n12667, ZN => n19010);
   U5199 : NAND2_X1 port map( A1 => n19147, A2 => n736, ZN => n14378);
   U5207 : NAND2_X1 port map( A1 => n18343, A2 => n18342, ZN => n15133);
   U5210 : AOI21_X1 port map( A1 => n18589, A2 => n8254, B => n1016, ZN => 
                           n8257);
   U5225 : OAI21_X1 port map( A1 => n10702, A2 => n9618, B => n14424, ZN => 
                           n5134);
   U5246 : OAI21_X1 port map( A1 => n13944, A2 => n13943, B => n21703, ZN => 
                           n2261);
   U5253 : NAND2_X1 port map( A1 => n6910, A2 => n15539, ZN => n17975);
   U5257 : NAND2_X1 port map( A1 => n17990, A2 => n17991, ZN => n17995);
   U5262 : AOI21_X1 port map( A1 => n17663, A2 => n1024, B => n1209, ZN => 
                           n6413);
   U5274 : NAND2_X1 port map( A1 => n5317, A2 => n5368, ZN => n17663);
   U5280 : INV_X2 port map( I => n17952, ZN => n788);
   U5284 : NOR2_X1 port map( A1 => n23105, A2 => n17520, ZN => n9778);
   U5302 : INV_X1 port map( I => n13727, ZN => n17498);
   U5311 : INV_X2 port map( I => n6624, ZN => n17401);
   U5321 : INV_X2 port map( I => n4334, ZN => n8424);
   U5327 : NAND3_X1 port map( A1 => n10597, A2 => n10502, A3 => n16652, ZN => 
                           n10295);
   U5336 : INV_X1 port map( I => n12224, ZN => n15203);
   U5340 : INV_X1 port map( I => n1241, ZN => n15107);
   U5342 : AOI21_X1 port map( A1 => n15951, A2 => n16224, B => n4644, ZN => 
                           n6661);
   U5345 : INV_X1 port map( I => n6687, ZN => n16715);
   U5355 : INV_X1 port map( I => n22296, ZN => n7758);
   U5357 : AND2_X1 port map( A1 => n26578, A2 => n12434, Z => n12669);
   U5359 : OR2_X1 port map( A1 => n12482, A2 => n11908, Z => n11005);
   U5372 : NAND2_X1 port map( A1 => n16219, A2 => n16076, ZN => n11081);
   U5375 : OAI21_X1 port map( A1 => n16083, A2 => n15497, B => n12035, ZN => 
                           n11006);
   U5378 : INV_X1 port map( I => n16316, ZN => n14942);
   U5379 : NOR2_X1 port map( A1 => n16329, A2 => n720, ZN => n5615);
   U5381 : NOR2_X1 port map( A1 => n7022, A2 => n13430, ZN => n7064);
   U5383 : INV_X1 port map( I => n15982, ZN => n16017);
   U5399 : CLKBUF_X2 port map( I => n16190, Z => n11568);
   U5404 : INV_X1 port map( I => n15892, ZN => n13306);
   U5407 : CLKBUF_X2 port map( I => Key(191), Z => n21642);
   U5411 : AOI22_X1 port map( A1 => n5004, A2 => n25369, B1 => n5360, B2 => 
                           n21413, ZN => n5002);
   U5413 : OAI22_X1 port map( A1 => n8446, A2 => n25325, B1 => n3650, B2 => 
                           n6051, ZN => n7119);
   U5420 : INV_X2 port map( I => n14437, ZN => n933);
   U5427 : NOR2_X1 port map( A1 => n21588, A2 => n21589, ZN => n8272);
   U5431 : OAI22_X1 port map( A1 => n5752, A2 => n20921, B1 => n15021, B2 => 
                           n5797, ZN => n4244);
   U5437 : INV_X1 port map( I => n1083, ZN => n4847);
   U5439 : OAI21_X1 port map( A1 => n21020, A2 => n1090, B => n2865, ZN => 
                           n3303);
   U5445 : INV_X1 port map( I => n21443, ZN => n21593);
   U5451 : INV_X1 port map( I => n21619, ZN => n21616);
   U5452 : INV_X1 port map( I => n13855, ZN => n21149);
   U5454 : OAI21_X1 port map( A1 => n956, A2 => n260, B => n25418, ZN => n8508)
                           ;
   U5490 : NOR2_X1 port map( A1 => n8326, A2 => n19689, ZN => n19826);
   U5498 : NAND2_X1 port map( A1 => n19889, A2 => n15067, ZN => n3988);
   U5500 : AOI21_X1 port map( A1 => n12738, A2 => n10881, B => n10601, ZN => 
                           n3102);
   U5504 : NOR2_X1 port map( A1 => n10957, A2 => n1129, ZN => n10863);
   U5513 : NOR2_X1 port map( A1 => n971, A2 => n14319, ZN => n1609);
   U5516 : INV_X2 port map( I => n19899, ZN => n19836);
   U5517 : NOR2_X1 port map( A1 => n19889, A2 => n19888, ZN => n3920);
   U5528 : NAND2_X1 port map( A1 => n24135, A2 => n968, ZN => n11063);
   U5543 : OAI21_X1 port map( A1 => n11445, A2 => n9873, B => n3830, ZN => 
                           n6749);
   U5544 : INV_X1 port map( I => n11445, ZN => n1135);
   U5549 : NAND2_X1 port map( A1 => n13229, A2 => n778, ZN => n1895);
   U5555 : NAND2_X1 port map( A1 => n19143, A2 => n25514, ZN => n18861);
   U5565 : AOI22_X1 port map( A1 => n14119, A2 => n15502, B1 => n19159, B2 => 
                           n22345, ZN => n2818);
   U5590 : NOR2_X1 port map( A1 => n760, A2 => n9041, ZN => n9272);
   U5592 : NOR2_X1 port map( A1 => n11035, A2 => n8624, ZN => n8623);
   U5601 : NAND2_X1 port map( A1 => n18666, A2 => n2081, ZN => n7578);
   U5602 : NOR2_X1 port map( A1 => n22973, A2 => n10556, ZN => n8944);
   U5626 : INV_X1 port map( I => n18414, ZN => n18413);
   U5634 : INV_X2 port map( I => n15349, ZN => n18344);
   U5654 : NAND2_X1 port map( A1 => n6098, A2 => n7981, ZN => n7984);
   U5679 : INV_X1 port map( I => n17458, ZN => n7656);
   U5687 : NOR2_X1 port map( A1 => n17498, A2 => n17497, ZN => n3936);
   U5689 : INV_X2 port map( I => n1038, ZN => n896);
   U5696 : AND2_X1 port map( A1 => n898, A2 => n15514, Z => n7016);
   U5706 : INV_X1 port map( I => n619, ZN => n17413);
   U5712 : INV_X1 port map( I => n17221, ZN => n17557);
   U5729 : NAND2_X1 port map( A1 => n8722, A2 => n26262, ZN => n5731);
   U5736 : OR2_X1 port map( A1 => n16693, A2 => n912, Z => n5849);
   U5740 : AND3_X1 port map( A1 => n9683, A2 => n16610, A3 => n4683, Z => 
                           n15912);
   U5744 : NAND2_X1 port map( A1 => n13039, A2 => n7132, ZN => n16578);
   U5749 : NOR2_X1 port map( A1 => n23107, A2 => n16678, ZN => n6403);
   U5755 : NOR2_X1 port map( A1 => n25940, A2 => n5324, ZN => n16684);
   U5758 : INV_X1 port map( I => n5310, ZN => n16688);
   U5761 : NAND2_X1 port map( A1 => n16618, A2 => n11908, ZN => n16634);
   U5771 : OAI21_X1 port map( A1 => n14150, A2 => n16135, B => n15878, ZN => 
                           n14793);
   U5776 : NOR2_X1 port map( A1 => n13343, A2 => n22623, ZN => n11518);
   U5777 : NAND2_X1 port map( A1 => n16089, A2 => n16226, ZN => n3405);
   U5778 : OAI21_X1 port map( A1 => n13103, A2 => n16254, B => n5050, ZN => 
                           n11007);
   U5781 : AND2_X1 port map( A1 => n11291, A2 => n14218, Z => n16051);
   U5783 : NAND2_X1 port map( A1 => n16278, A2 => n16279, ZN => n8972);
   U5785 : NOR2_X1 port map( A1 => n13430, A2 => n16300, ZN => n12760);
   U5791 : NAND2_X1 port map( A1 => n8684, A2 => n1059, ZN => n15920);
   U5797 : NOR2_X1 port map( A1 => n3193, A2 => n16115, ZN => n13955);
   U5799 : INV_X1 port map( I => n21876, ZN => n15615);
   U5804 : NOR3_X1 port map( A1 => n16334, A2 => n15282, A3 => n7266, ZN => 
                           n12919);
   U5807 : NAND2_X1 port map( A1 => n16343, A2 => n16342, ZN => n16344);
   U5809 : INV_X2 port map( I => n563, ZN => n16069);
   U5814 : INV_X1 port map( I => n16253, ZN => n13103);
   U5817 : INV_X1 port map( I => n14463, ZN => n1279);
   U5818 : BUF_X2 port map( I => n14433, Z => n5680);
   U5820 : INV_X1 port map( I => n20605, ZN => n920);
   U5825 : INV_X1 port map( I => n7397, ZN => n1301);
   U5827 : INV_X1 port map( I => n15834, ZN => n921);
   U5829 : INV_X1 port map( I => n21143, ZN => n924);
   U5830 : INV_X1 port map( I => n20952, ZN => n922);
   U5831 : INV_X1 port map( I => n14518, ZN => n923);
   U5832 : INV_X1 port map( I => n21742, ZN => n925);
   U5833 : INV_X1 port map( I => n14473, ZN => n919);
   U5836 : BUF_X1 port map( I => Key(75), Z => n21341);
   U5838 : CLKBUF_X2 port map( I => Key(97), Z => n21703);
   U5839 : INV_X2 port map( I => n9218, ZN => n841);
   U5840 : CLKBUF_X2 port map( I => Key(67), Z => n14550);
   U5842 : CLKBUF_X2 port map( I => Key(91), Z => n21143);
   U5844 : CLKBUF_X2 port map( I => Key(172), Z => n14633);
   U5850 : NOR2_X1 port map( A1 => n21040, A2 => n10635, ZN => n5659);
   U5857 : NAND3_X1 port map( A1 => n7827, A2 => n24562, A3 => n7826, ZN => 
                           n9302);
   U5860 : NOR2_X1 port map( A1 => n22764, A2 => n4315, ZN => n6248);
   U5861 : NAND3_X1 port map( A1 => n24562, A2 => n20878, A3 => n802, ZN => 
                           n4849);
   U5864 : OAI21_X1 port map( A1 => n8447, A2 => n25325, B => n20752, ZN => 
                           n20743);
   U5867 : NOR2_X1 port map( A1 => n22794, A2 => n25370, ZN => n11466);
   U5871 : NOR2_X1 port map( A1 => n12061, A2 => n2777, ZN => n1659);
   U5875 : NAND2_X1 port map( A1 => n20691, A2 => n934, ZN => n3756);
   U5880 : NAND3_X1 port map( A1 => n21290, A2 => n21286, A3 => n749, ZN => 
                           n6092);
   U5883 : NAND2_X1 port map( A1 => n802, A2 => n20875, ZN => n7826);
   U5884 : NAND2_X1 port map( A1 => n8389, A2 => n934, ZN => n2916);
   U5892 : NAND3_X1 port map( A1 => n15742, A2 => n20910, A3 => n26006, ZN => 
                           n2840);
   U5894 : OR2_X1 port map( A1 => n12846, A2 => n11385, Z => n11384);
   U5896 : NAND2_X1 port map( A1 => n21212, A2 => n9494, ZN => n21220);
   U5898 : NOR2_X1 port map( A1 => n20878, A2 => n3971, ZN => n4170);
   U5903 : OAI21_X1 port map( A1 => n14583, A2 => n21008, B => n937, ZN => 
                           n3740);
   U5906 : NAND2_X1 port map( A1 => n20875, A2 => n20879, ZN => n8163);
   U5907 : INV_X1 port map( I => n20748, ZN => n5812);
   U5908 : AND2_X1 port map( A1 => n15287, A2 => n4822, Z => n4821);
   U5910 : AOI22_X1 port map( A1 => n25329, A2 => n20704, B1 => n9563, B2 => 
                           n27429, ZN => n2114);
   U5912 : NOR2_X1 port map( A1 => n12251, A2 => n13888, ZN => n21284);
   U5919 : INV_X2 port map( I => n10992, ZN => n845);
   U5923 : OAI21_X1 port map( A1 => n21094, A2 => n14341, B => n25173, ZN => 
                           n3788);
   U5932 : AOI21_X1 port map( A1 => n2184, A2 => n20860, B => n20857, ZN => 
                           n2183);
   U5941 : NAND2_X1 port map( A1 => n20882, A2 => n20932, ZN => n20883);
   U5942 : AND2_X1 port map( A1 => n12140, A2 => n20755, Z => n6407);
   U5945 : OR2_X1 port map( A1 => n772, A2 => n24209, Z => n10675);
   U5949 : AND2_X1 port map( A1 => n21387, A2 => n21275, Z => n5252);
   U5959 : INV_X1 port map( I => n21162, ZN => n13052);
   U5973 : NAND2_X1 port map( A1 => n21667, A2 => n21629, ZN => n21574);
   U5974 : NOR2_X1 port map( A1 => n20730, A2 => n9728, ZN => n8492);
   U5983 : OAI21_X1 port map( A1 => n15689, A2 => n20739, B => n20633, ZN => 
                           n20507);
   U5984 : INV_X1 port map( I => n20975, ZN => n21070);
   U5985 : NOR2_X1 port map( A1 => n20781, A2 => n20739, ZN => n5540);
   U5990 : INV_X1 port map( I => n20899, ZN => n7880);
   U5993 : NOR2_X1 port map( A1 => n10031, A2 => n23036, ZN => n6788);
   U5996 : NAND3_X1 port map( A1 => n20633, A2 => n20786, A3 => n20781, ZN => 
                           n6735);
   U6004 : NOR2_X1 port map( A1 => n5550, A2 => n20736, ZN => n5806);
   U6007 : INV_X1 port map( I => n20901, ZN => n20857);
   U6015 : NAND3_X1 port map( A1 => n3060, A2 => n15703, A3 => n21759, ZN => 
                           n5649);
   U6018 : NOR2_X1 port map( A1 => n2718, A2 => n9960, ZN => n2717);
   U6036 : AND2_X1 port map( A1 => n20237, A2 => n28519, Z => n10616);
   U6039 : OAI21_X1 port map( A1 => n20323, A2 => n12712, B => n1756, ZN => 
                           n1755);
   U6040 : INV_X1 port map( I => n8910, ZN => n9219);
   U6048 : NOR2_X1 port map( A1 => n8905, A2 => n2185, ZN => n8908);
   U6054 : NAND2_X1 port map( A1 => n1640, A2 => n20255, ZN => n1639);
   U6057 : INV_X1 port map( I => n20174, ZN => n20270);
   U6066 : OAI21_X1 port map( A1 => n6264, A2 => n23771, B => n26252, ZN => 
                           n5378);
   U6076 : OAI21_X1 port map( A1 => n20190, A2 => n13104, B => n26710, ZN => 
                           n2718);
   U6112 : NOR2_X1 port map( A1 => n19520, A2 => n974, ZN => n8911);
   U6128 : NAND2_X1 port map( A1 => n24196, A2 => n4246, ZN => n19520);
   U6135 : NOR2_X1 port map( A1 => n814, A2 => n10601, ZN => n10095);
   U6156 : NOR3_X1 port map( A1 => n10881, A2 => n814, A3 => n19819, ZN => 
                           n9627);
   U6163 : AOI22_X1 port map( A1 => n15383, A2 => n14319, B1 => n19948, B2 => 
                           n19830, ZN => n1610);
   U6169 : NOR2_X1 port map( A1 => n19883, A2 => n9887, ZN => n6570);
   U6183 : NOR2_X1 port map( A1 => n19951, A2 => n19714, ZN => n6552);
   U6184 : INV_X1 port map( I => n7340, ZN => n19941);
   U6197 : AND2_X1 port map( A1 => n3563, A2 => n14929, Z => n8417);
   U6234 : NAND2_X1 port map( A1 => n1658, A2 => n3619, ZN => n7570);
   U6249 : AOI21_X1 port map( A1 => n18924, A2 => n14382, B => n14925, ZN => 
                           n13636);
   U6259 : NOR3_X1 port map( A1 => n7533, A2 => n19140, A3 => n4224, ZN => 
                           n1331);
   U6266 : NAND2_X1 port map( A1 => n996, A2 => n9538, ZN => n2395);
   U6278 : NAND3_X1 port map( A1 => n23060, A2 => n11476, A3 => n11475, ZN => 
                           n11477);
   U6282 : INV_X1 port map( I => n12338, ZN => n18948);
   U6283 : INV_X2 port map( I => n1716, ZN => n869);
   U6292 : OR2_X2 port map( A1 => n18365, A2 => n18368, Z => n18396);
   U6299 : AOI22_X1 port map( A1 => n9272, A2 => n647, B1 => n18494, B2 => 
                           n9041, ZN => n9270);
   U6310 : NAND2_X1 port map( A1 => n8257, A2 => n2564, ZN => n2563);
   U6319 : NAND2_X1 port map( A1 => n18653, A2 => n9041, ZN => n7099);
   U6324 : AND2_X1 port map( A1 => n9041, A2 => n18741, Z => n18495);
   U6330 : AOI21_X1 port map( A1 => n1009, A2 => n25828, B => n18752, ZN => 
                           n5621);
   U6333 : AOI21_X1 port map( A1 => n9464, A2 => n18773, B => n22814, ZN => 
                           n3310);
   U6338 : OAI22_X1 port map( A1 => n11161, A2 => n1004, B1 => n15449, B2 => 
                           n14207, ZN => n2946);
   U6345 : AOI21_X1 port map( A1 => n18682, A2 => n24054, B => n11911, ZN => 
                           n8616);
   U6350 : NAND3_X1 port map( A1 => n3202, A2 => n24243, A3 => n7095, ZN => 
                           n14500);
   U6351 : NOR2_X1 port map( A1 => n18715, A2 => n1014, ZN => n2154);
   U6352 : NAND3_X1 port map( A1 => n5434, A2 => n18583, A3 => n4639, ZN => 
                           n7742);
   U6359 : OAI22_X1 port map( A1 => n1180, A2 => n7960, B1 => n18776, B2 => 
                           n1017, ZN => n11142);
   U6370 : NAND2_X1 port map( A1 => n14308, A2 => n24047, ZN => n15172);
   U6403 : INV_X2 port map( I => n10542, ZN => n879);
   U6413 : INV_X1 port map( I => n18155, ZN => n1193);
   U6415 : INV_X1 port map( I => n13840, ZN => n12102);
   U6449 : NOR2_X1 port map( A1 => n15539, A2 => n5153, ZN => n5152);
   U6464 : NAND2_X1 port map( A1 => n7599, A2 => n17935, ZN => n8614);
   U6493 : NAND2_X1 port map( A1 => n1349, A2 => n17935, ZN => n8521);
   U6510 : INV_X2 port map( I => n2636, ZN => n890);
   U6528 : NAND2_X1 port map( A1 => n17427, A2 => n26532, ZN => n11029);
   U6531 : NOR3_X1 port map( A1 => n27648, A2 => n24070, A3 => n461, ZN => 
                           n5563);
   U6541 : NAND2_X1 port map( A1 => n25504, A2 => n9827, ZN => n5187);
   U6544 : NOR2_X1 port map( A1 => n15699, A2 => n9132, ZN => n10911);
   U6545 : NOR2_X1 port map( A1 => n2963, A2 => n17175, ZN => n9287);
   U6556 : NAND2_X1 port map( A1 => n9570, A2 => n9569, ZN => n9568);
   U6572 : INV_X1 port map( I => n17485, ZN => n11436);
   U6576 : NOR2_X1 port map( A1 => n1231, A2 => n17522, ZN => n4687);
   U6577 : NOR2_X1 port map( A1 => n636, A2 => n17519, ZN => n9984);
   U6591 : OR2_X1 port map( A1 => n5473, A2 => n13048, Z => n17576);
   U6598 : NOR2_X1 port map( A1 => n17317, A2 => n17318, ZN => n5258);
   U6600 : NAND2_X1 port map( A1 => n10150, A2 => n10577, ZN => n11435);
   U6605 : AND2_X1 port map( A1 => n613, A2 => n14997, Z => n8661);
   U6622 : INV_X1 port map( I => n5169, ZN => n17346);
   U6625 : INV_X1 port map( I => n28025, ZN => n1222);
   U6627 : INV_X2 port map( I => n8193, ZN => n17522);
   U6632 : INV_X1 port map( I => n17185, ZN => n2537);
   U6641 : INV_X2 port map( I => n11966, ZN => n899);
   U6642 : INV_X2 port map( I => n8795, ZN => n900);
   U6651 : NAND2_X1 port map( A1 => n16400, A2 => n8901, ZN => n9392);
   U6657 : NAND2_X1 port map( A1 => n14632, A2 => n10282, ZN => n10281);
   U6664 : OAI21_X1 port map( A1 => n1992, A2 => n15351, B => n13025, ZN => 
                           n6565);
   U6665 : OAI22_X1 port map( A1 => n16713, A2 => n3297, B1 => n1053, B2 => 
                           n6373, ZN => n6880);
   U6667 : INV_X1 port map( I => n15912, ZN => n8845);
   U6669 : AND2_X1 port map( A1 => n22061, A2 => n26262, Z => n8511);
   U6672 : AOI21_X1 port map( A1 => n16413, A2 => n1053, B => n16713, ZN => 
                           n14698);
   U6676 : NAND2_X1 port map( A1 => n14137, A2 => n24646, ZN => n16621);
   U6678 : NOR3_X1 port map( A1 => n16688, A2 => n1048, A3 => n2149, ZN => 
                           n2301);
   U6679 : NAND2_X1 port map( A1 => n16715, A2 => n6688, ZN => n16414);
   U6683 : NAND2_X1 port map( A1 => n16605, A2 => n2131, ZN => n16606);
   U6685 : NOR2_X1 port map( A1 => n8901, A2 => n13690, ZN => n9391);
   U6690 : INV_X1 port map( I => n16587, ZN => n1242);
   U6694 : INV_X1 port map( I => n6110, ZN => n11383);
   U6696 : OAI21_X1 port map( A1 => n24552, A2 => n16518, B => n434, ZN => 
                           n7542);
   U6702 : NAND2_X1 port map( A1 => n16711, A2 => n23128, ZN => n12368);
   U6707 : NAND4_X1 port map( A1 => n15777, A2 => n15794, A3 => n15778, A4 => 
                           n13402, ZN => n16577);
   U6711 : INV_X1 port map( I => n3443, ZN => n16702);
   U6712 : NAND2_X1 port map( A1 => n7132, A2 => n11122, ZN => n16437);
   U6718 : AND2_X1 port map( A1 => n16630, A2 => n23744, Z => n11721);
   U6727 : NAND2_X1 port map( A1 => n6683, A2 => n16571, ZN => n1646);
   U6730 : INV_X1 port map( I => n3479, ZN => n9500);
   U6737 : NOR2_X1 port map( A1 => n11565, A2 => n11564, ZN => n11567);
   U6747 : NOR2_X1 port map( A1 => n1881, A2 => n3370, ZN => n3369);
   U6750 : NOR2_X1 port map( A1 => n16202, A2 => n8684, ZN => n8241);
   U6751 : NAND2_X1 port map( A1 => n1843, A2 => n2148, ZN => n1841);
   U6754 : NAND2_X1 port map( A1 => n14644, A2 => n16115, ZN => n3370);
   U6757 : NOR2_X1 port map( A1 => n13776, A2 => n15930, ZN => n8087);
   U6762 : NOR2_X1 port map( A1 => n16242, A2 => n9768, ZN => n7649);
   U6766 : NAND2_X1 port map( A1 => n6122, A2 => n16321, ZN => n6118);
   U6768 : AOI22_X1 port map( A1 => n12760, A2 => n16188, B1 => n16189, B2 => 
                           n16300, ZN => n12763);
   U6769 : AOI22_X1 port map( A1 => n5455, A2 => n1058, B1 => n16353, B2 => 
                           n23270, ZN => n6635);
   U6772 : NOR2_X1 port map( A1 => n16069, A2 => n16088, ZN => n7869);
   U6780 : NOR2_X1 port map( A1 => n16188, A2 => n24271, ZN => n11564);
   U6781 : NOR2_X1 port map( A1 => n14293, A2 => n1062, ZN => n1866);
   U6784 : NAND2_X1 port map( A1 => n1260, A2 => n16287, ZN => n5789);
   U6793 : NAND2_X1 port map( A1 => n13307, A2 => n7053, ZN => n2556);
   U6794 : AOI21_X1 port map( A1 => n836, A2 => n16062, B => n16063, ZN => 
                           n2555);
   U6796 : NOR2_X1 port map( A1 => n28166, A2 => n14293, ZN => n11647);
   U6797 : OAI21_X1 port map( A1 => n12010, A2 => n5362, B => n121, ZN => n3956
                           );
   U6799 : NAND2_X1 port map( A1 => n5681, A2 => n6886, ZN => n1843);
   U6801 : AND3_X1 port map( A1 => n16069, A2 => n14142, A3 => n13562, Z => 
                           n11875);
   U6802 : NAND2_X1 port map( A1 => n5580, A2 => n15924, ZN => n10452);
   U6805 : AOI21_X1 port map( A1 => n16344, A2 => n25570, B => n28166, ZN => 
                           n16345);
   U6808 : NOR2_X1 port map( A1 => n16320, A2 => n16317, ZN => n6120);
   U6809 : AOI21_X1 port map( A1 => n28152, A2 => n16335, B => n7053, ZN => 
                           n1718);
   U6811 : NOR2_X1 port map( A1 => n16320, A2 => n7311, ZN => n4784);
   U6814 : NAND2_X1 port map( A1 => n16321, A2 => n16317, ZN => n15947);
   U6821 : NOR2_X1 port map( A1 => n14385, A2 => n798, ZN => n13602);
   U6826 : NOR2_X1 port map( A1 => n16193, A2 => n14989, ZN => n12154);
   U6835 : INV_X1 port map( I => n16354, ZN => n1266);
   U6837 : INV_X1 port map( I => n4346, ZN => n16277);
   U6838 : AND2_X1 port map( A1 => n7608, A2 => n6886, Z => n5455);
   U6839 : INV_X1 port map( I => n10573, ZN => n13857);
   U6850 : INV_X1 port map( I => n14433, ZN => n5681);
   U6851 : INV_X1 port map( I => n21044, ZN => n1064);
   U6852 : INV_X1 port map( I => n19218, ZN => n1061);
   U6853 : INV_X2 port map( I => n15354, ZN => n16321);
   U6854 : INV_X1 port map( I => n11628, ZN => n16225);
   U6860 : CLKBUF_X2 port map( I => Key(35), Z => n14623);
   U6866 : CLKBUF_X2 port map( I => Key(96), Z => n20467);
   U6868 : CLKBUF_X2 port map( I => Key(175), Z => n14631);
   U6875 : CLKBUF_X2 port map( I => Key(72), Z => n20880);
   U6876 : CLKBUF_X2 port map( I => Key(109), Z => n21313);
   U6877 : CLKBUF_X2 port map( I => Key(169), Z => n21210);
   U6878 : OAI21_X1 port map( A1 => n5660, A2 => n5659, B => n25352, ZN => 
                           n5658);
   U6880 : OAI21_X1 port map( A1 => n9425, A2 => n21040, B => n21030, ZN => 
                           n5662);
   U6881 : NAND2_X1 port map( A1 => n6037, A2 => n20878, ZN => n9301);
   U6882 : AOI21_X1 port map( A1 => n21290, A2 => n14024, B => n847, ZN => 
                           n6055);
   U6885 : NAND2_X1 port map( A1 => n2778, A2 => n1659, ZN => n6034);
   U6892 : NAND3_X1 port map( A1 => n5813, A2 => n20750, A3 => n5812, ZN => 
                           n5811);
   U6893 : NAND2_X1 port map( A1 => n842, A2 => n8935, ZN => n10430);
   U6894 : NAND2_X1 port map( A1 => n20697, A2 => n480, ZN => n20698);
   U6895 : AOI21_X1 port map( A1 => n13553, A2 => n20879, B => n24562, ZN => 
                           n8160);
   U6897 : AOI21_X1 port map( A1 => n8163, A2 => n8162, B => n1070, ZN => n8161
                           );
   U6901 : OAI21_X1 port map( A1 => n13743, A2 => n5360, B => n25370, ZN => 
                           n11459);
   U6902 : INV_X1 port map( I => n20696, ZN => n3755);
   U6904 : NAND2_X1 port map( A1 => n9460, A2 => n845, ZN => n21704);
   U6913 : AOI21_X1 port map( A1 => n22797, A2 => n10635, B => n21052, ZN => 
                           n21047);
   U6916 : NOR3_X1 port map( A1 => n4170, A2 => n27468, A3 => n20875, ZN => 
                           n5736);
   U6918 : NOR2_X1 port map( A1 => n21355, A2 => n21342, ZN => n7291);
   U6920 : NAND3_X1 port map( A1 => n4766, A2 => n848, A3 => n844, ZN => n4935)
                           ;
   U6921 : OAI21_X1 port map( A1 => n21291, A2 => n21290, B => n749, ZN => 
                           n5847);
   U6923 : AOI21_X1 port map( A1 => n25377, A2 => n3642, B => n21173, ZN => 
                           n3641);
   U6930 : NAND2_X1 port map( A1 => n22824, A2 => n13888, ZN => n6095);
   U6933 : INV_X1 port map( I => n21111, ZN => n21113);
   U6939 : NAND2_X1 port map( A1 => n15742, A2 => n20917, ZN => n4729);
   U6945 : NAND2_X1 port map( A1 => n847, A2 => n12251, ZN => n6056);
   U6946 : OR2_X1 port map( A1 => n13021, A2 => n7454, Z => n7453);
   U6953 : INV_X2 port map( I => n7085, ZN => n21564);
   U6955 : INV_X4 port map( I => n22730, ZN => n934);
   U6959 : NAND2_X1 port map( A1 => n7663, A2 => n3992, ZN => n3991);
   U6969 : NOR2_X1 port map( A1 => n20643, A2 => n10588, ZN => n3995);
   U6971 : AND2_X1 port map( A1 => n5726, A2 => n20931, Z => n20780);
   U6972 : AOI21_X1 port map( A1 => n15365, A2 => n15364, B => n25326, ZN => 
                           n13400);
   U6979 : NOR2_X1 port map( A1 => n20938, A2 => n10483, ZN => n10482);
   U6980 : NOR2_X1 port map( A1 => n8594, A2 => n20732, ZN => n20731);
   U6993 : OR2_X1 port map( A1 => n20710, A2 => n10610, Z => n20747);
   U7004 : AND2_X1 port map( A1 => n852, A2 => n22823, Z => n21359);
   U7006 : NAND2_X1 port map( A1 => n21727, A2 => n1091, ZN => n10394);
   U7009 : OAI21_X1 port map( A1 => n13432, A2 => n773, B => n5781, ZN => 
                           n12586);
   U7010 : NAND2_X1 port map( A1 => n26505, A2 => n21457, ZN => n11164);
   U7012 : OAI21_X1 port map( A1 => n24576, A2 => n28305, B => n15103, ZN => 
                           n21726);
   U7014 : NAND2_X1 port map( A1 => n21586, A2 => n13979, ZN => n21588);
   U7016 : OR2_X1 port map( A1 => n26650, A2 => n21324, Z => n10254);
   U7025 : AND2_X1 port map( A1 => n21099, A2 => n26512, Z => n9676);
   U7030 : NAND2_X1 port map( A1 => n20507, A2 => n20635, ZN => n2623);
   U7037 : AND2_X1 port map( A1 => n21058, A2 => n20972, Z => n20973);
   U7042 : NOR2_X1 port map( A1 => n21161, A2 => n13049, ZN => n21162);
   U7048 : AND2_X1 port map( A1 => n21714, A2 => n20642, Z => n9672);
   U7058 : INV_X1 port map( I => n1090, ZN => n21069);
   U7060 : NAND2_X1 port map( A1 => n9378, A2 => n3559, ZN => n3561);
   U7067 : BUF_X2 port map( I => n12585, Z => n8668);
   U7069 : INV_X1 port map( I => n21728, ZN => n20591);
   U7072 : INV_X2 port map( I => n15353, ZN => n952);
   U7080 : OR2_X2 port map( A1 => n9083, A2 => n10026, Z => n7011);
   U7085 : NAND2_X1 port map( A1 => n3967, A2 => n27398, ZN => n3966);
   U7087 : NAND2_X1 port map( A1 => n4782, A2 => n22758, ZN => n4781);
   U7088 : NAND2_X1 port map( A1 => n20239, A2 => n20238, ZN => n2470);
   U7090 : NAND2_X1 port map( A1 => n20256, A2 => n1106, ZN => n2074);
   U7091 : NAND2_X1 port map( A1 => n1639, A2 => n1106, ZN => n1642);
   U7099 : NOR2_X1 port map( A1 => n8932, A2 => n5378, ZN => n8931);
   U7100 : NAND2_X1 port map( A1 => n1108, A2 => n6670, ZN => n14398);
   U7107 : AOI21_X1 port map( A1 => n8642, A2 => n20021, B => n5575, ZN => 
                           n9341);
   U7110 : AOI21_X1 port map( A1 => n20316, A2 => n14513, B => n22815, ZN => 
                           n13716);
   U7137 : INV_X1 port map( I => n20073, ZN => n20144);
   U7138 : NAND2_X1 port map( A1 => n9579, A2 => n6511, ZN => n1640);
   U7146 : NOR2_X1 port map( A1 => n24533, A2 => n27091, ZN => n20272);
   U7148 : INV_X4 port map( I => n27349, ZN => n956);
   U7153 : INV_X1 port map( I => n27091, ZN => n8507);
   U7158 : INV_X1 port map( I => n20183, ZN => n13995);
   U7168 : NAND2_X1 port map( A1 => n20273, A2 => n25389, ZN => n19664);
   U7170 : INV_X1 port map( I => n10007, ZN => n20313);
   U7179 : NAND2_X1 port map( A1 => n12401, A2 => n19625, ZN => n13655);
   U7180 : OAI21_X1 port map( A1 => n15027, A2 => n19782, B => n3954, ZN => 
                           n19641);
   U7189 : NOR2_X1 port map( A1 => n10498, A2 => n863, ZN => n1655);
   U7190 : OAI21_X1 port map( A1 => n10096, A2 => n10095, B => n10881, ZN => 
                           n10094);
   U7203 : NOR2_X1 port map( A1 => n14170, A2 => n811, ZN => n2209);
   U7208 : NAND2_X1 port map( A1 => n4432, A2 => n14279, ZN => n4435);
   U7215 : NAND2_X1 port map( A1 => n19696, A2 => n11353, ZN => n3424);
   U7224 : INV_X1 port map( I => n19099, ZN => n1348);
   U7225 : OR3_X1 port map( A1 => n25236, A2 => n34, A3 => n12863, Z => n19576)
                           ;
   U7230 : OAI21_X1 port map( A1 => n4432, A2 => n19759, B => n26522, ZN => 
                           n6560);
   U7232 : AOI21_X1 port map( A1 => n4132, A2 => n19743, B => n24235, ZN => 
                           n2739);
   U7238 : AND3_X1 port map( A1 => n19915, A2 => n14459, A3 => n204, Z => n7293
                           );
   U7239 : NOR2_X1 port map( A1 => n11078, A2 => n10978, ZN => n8172);
   U7246 : AND2_X1 port map( A1 => n1122, A2 => n19758, Z => n4437);
   U7247 : NAND2_X1 port map( A1 => n13278, A2 => n19913, ZN => n7068);
   U7249 : NAND2_X1 port map( A1 => n19859, A2 => n1119, ZN => n11987);
   U7259 : NAND2_X1 port map( A1 => n3835, A2 => n19752, ZN => n6191);
   U7264 : NAND2_X1 port map( A1 => n1129, A2 => n8326, ZN => n10207);
   U7266 : NOR2_X1 port map( A1 => n1122, A2 => n19758, ZN => n6189);
   U7272 : AOI21_X1 port map( A1 => n19955, A2 => n19468, B => n19949, ZN => 
                           n13383);
   U7276 : NAND2_X1 port map( A1 => n28285, A2 => n10121, ZN => n9646);
   U7285 : NAND2_X1 port map( A1 => n3584, A2 => n14307, ZN => n5331);
   U7287 : INV_X1 port map( I => n3954, ZN => n19783);
   U7290 : INV_X1 port map( I => n11287, ZN => n15310);
   U7292 : NAND2_X1 port map( A1 => n19828, A2 => n19714, ZN => n19716);
   U7294 : OR2_X1 port map( A1 => n19843, A2 => n15457, Z => n19841);
   U7304 : INV_X2 port map( I => n5209, ZN => n14929);
   U7305 : INV_X2 port map( I => n8838, ZN => n10613);
   U7308 : BUF_X2 port map( I => n12286, Z => n11213);
   U7309 : BUF_X2 port map( I => n19666, Z => n12431);
   U7326 : NOR2_X1 port map( A1 => n18966, A2 => n14272, ZN => n5109);
   U7352 : INV_X1 port map( I => n13636, ZN => n2168);
   U7357 : AOI21_X1 port map( A1 => n10164, A2 => n19043, B => n26097, ZN => 
                           n6784);
   U7361 : INV_X1 port map( I => n21767, ZN => n13659);
   U7365 : NAND2_X1 port map( A1 => n21915, A2 => n8729, ZN => n8728);
   U7373 : NAND2_X1 port map( A1 => n11477, A2 => n13563, ZN => n7032);
   U7377 : NAND2_X1 port map( A1 => n18931, A2 => n13887, ZN => n12750);
   U7385 : NAND2_X1 port map( A1 => n13946, A2 => n13371, ZN => n13671);
   U7386 : INV_X1 port map( I => n18917, ZN => n1415);
   U7390 : AOI21_X1 port map( A1 => n27175, A2 => n24061, B => n5114, ZN => 
                           n8914);
   U7391 : NAND2_X1 port map( A1 => n3383, A2 => n15058, ZN => n5441);
   U7393 : NAND2_X1 port map( A1 => n10171, A2 => n26764, ZN => n10170);
   U7401 : NOR2_X1 port map( A1 => n19033, A2 => n447, ZN => n19031);
   U7407 : NAND2_X1 port map( A1 => n28136, A2 => n6145, ZN => n9226);
   U7414 : NAND2_X1 port map( A1 => n12047, A2 => n11386, ZN => n15480);
   U7416 : NOR2_X1 port map( A1 => n13563, A2 => n12338, ZN => n4118);
   U7423 : NOR2_X1 port map( A1 => n15502, A2 => n22345, ZN => n19034);
   U7431 : OAI21_X1 port map( A1 => n12721, A2 => n14922, B => n19150, ZN => 
                           n8802);
   U7433 : INV_X1 port map( I => n4199, ZN => n18829);
   U7436 : NAND2_X1 port map( A1 => n19110, A2 => n28547, ZN => n8312);
   U7439 : NAND2_X1 port map( A1 => n13812, A2 => n4703, ZN => n5942);
   U7440 : OAI21_X1 port map( A1 => n18912, A2 => n26645, B => n18944, ZN => 
                           n9346);
   U7442 : NAND2_X1 port map( A1 => n4199, A2 => n25176, ZN => n4381);
   U7448 : NAND2_X1 port map( A1 => n25176, A2 => n11376, ZN => n15058);
   U7449 : NOR2_X1 port map( A1 => n8049, A2 => n27965, ZN => n18907);
   U7459 : INV_X2 port map( I => n14210, ZN => n11696);
   U7466 : OR2_X1 port map( A1 => n875, A2 => n26234, Z => n10271);
   U7471 : NAND4_X1 port map( A1 => n15725, A2 => n18376, A3 => n18382, A4 => 
                           n18375, ZN => n18913);
   U7472 : NOR2_X1 port map( A1 => n13483, A2 => n6277, ZN => n13482);
   U7489 : INV_X1 port map( I => n14037, ZN => n19128);
   U7493 : AOI21_X1 port map( A1 => n18424, A2 => n18755, B => n18674, ZN => 
                           n9600);
   U7495 : OAI21_X1 port map( A1 => n18719, A2 => n1189, B => n13372, ZN => 
                           n4331);
   U7507 : OR2_X1 port map( A1 => n18490, A2 => n27281, Z => n4387);
   U7513 : AND3_X1 port map( A1 => n27281, A2 => n10594, A3 => n18424, Z => 
                           n18006);
   U7514 : AOI21_X1 port map( A1 => n18715, A2 => n26317, B => n8746, ZN => 
                           n8745);
   U7521 : INV_X1 port map( I => n8333, ZN => n14121);
   U7526 : NOR2_X1 port map( A1 => n18783, A2 => n6031, ZN => n5880);
   U7533 : AOI21_X1 port map( A1 => n7591, A2 => n26036, B => n18728, ZN => 
                           n2135);
   U7535 : NOR2_X1 port map( A1 => n4639, A2 => n18377, ZN => n4642);
   U7543 : NAND2_X1 port map( A1 => n18706, A2 => n27895, ZN => n18707);
   U7553 : NOR2_X1 port map( A1 => n14138, A2 => n18629, ZN => n18404);
   U7557 : AND2_X1 port map( A1 => n2982, A2 => n24207, Z => n4089);
   U7558 : NAND2_X1 port map( A1 => n18727, A2 => n14594, ZN => n10216);
   U7564 : NOR2_X1 port map( A1 => n24207, A2 => n738, ZN => n12424);
   U7567 : INV_X2 port map( I => n5919, ZN => n18715);
   U7572 : NOR2_X1 port map( A1 => n10962, A2 => n1179, ZN => n10961);
   U7574 : NOR2_X1 port map( A1 => n881, A2 => n18124, ZN => n4542);
   U7575 : NAND2_X1 port map( A1 => n18344, A2 => n14369, ZN => n18461);
   U7578 : OAI21_X1 port map( A1 => n18448, A2 => n27241, B => n3554, ZN => 
                           n5827);
   U7581 : NAND2_X1 port map( A1 => n18753, A2 => n24522, ZN => n6312);
   U7601 : NOR2_X1 port map( A1 => n7383, A2 => n15137, ZN => n7739);
   U7604 : INV_X1 port map( I => n18457, ZN => n18474);
   U7606 : OAI21_X1 port map( A1 => n26051, A2 => n23361, B => n10958, ZN => 
                           n6205);
   U7615 : INV_X2 port map( I => n15423, ZN => n15660);
   U7627 : NAND2_X1 port map( A1 => n7314, A2 => n11514, ZN => n8306);
   U7633 : OAI21_X1 port map( A1 => n5953, A2 => n4237, B => n6287, ZN => n4236
                           );
   U7636 : INV_X1 port map( I => n18038, ZN => n18022);
   U7641 : OAI21_X1 port map( A1 => n4357, A2 => n4356, B => n4355, ZN => n4354
                           );
   U7642 : NAND3_X1 port map( A1 => n15682, A2 => n15681, A3 => n21712, ZN => 
                           n7800);
   U7653 : NAND2_X1 port map( A1 => n1569, A2 => n2524, ZN => n1567);
   U7655 : INV_X1 port map( I => n7002, ZN => n2435);
   U7657 : AND2_X1 port map( A1 => n1215, A2 => n6018, Z => n17641);
   U7661 : AND2_X1 port map( A1 => n21779, A2 => n17817, Z => n17820);
   U7664 : NOR2_X1 port map( A1 => n13237, A2 => n13236, ZN => n9164);
   U7673 : AND2_X1 port map( A1 => n2238, A2 => n25966, Z => n8323);
   U7674 : NOR2_X1 port map( A1 => n17798, A2 => n8070, ZN => n8183);
   U7677 : NOR2_X1 port map( A1 => n1512, A2 => n17678, ZN => n14599);
   U7683 : NAND2_X1 port map( A1 => n17635, A2 => n12964, ZN => n1864);
   U7684 : NAND2_X1 port map( A1 => n17963, A2 => n27947, ZN => n4503);
   U7693 : NAND2_X1 port map( A1 => n8521, A2 => n8009, ZN => n13236);
   U7711 : NOR2_X1 port map( A1 => n22812, A2 => n26643, ZN => n11632);
   U7733 : NOR2_X1 port map( A1 => n8849, A2 => n17349, ZN => n7991);
   U7736 : NAND3_X1 port map( A1 => n8889, A2 => n8888, A3 => n7834, ZN => 
                           n3716);
   U7749 : NAND2_X1 port map( A1 => n17683, A2 => n22851, ZN => n17684);
   U7750 : NOR2_X1 port map( A1 => n21791, A2 => n17605, ZN => n8784);
   U7751 : NOR2_X1 port map( A1 => n1893, A2 => n10779, ZN => n14053);
   U7754 : NAND2_X1 port map( A1 => n25106, A2 => n7108, ZN => n4245);
   U7755 : OAI21_X1 port map( A1 => n7961, A2 => n890, B => n23633, ZN => n4593
                           );
   U7764 : NOR2_X1 port map( A1 => n25926, A2 => n17969, ZN => n2222);
   U7793 : OAI21_X1 port map( A1 => n9984, A2 => n2756, B => n1701, ZN => n2755
                           );
   U7794 : NAND3_X1 port map( A1 => n1232, A2 => n831, A3 => n14354, ZN => 
                           n14353);
   U7799 : OR2_X1 port map( A1 => n17545, A2 => n14697, Z => n7082);
   U7807 : INV_X1 port map( I => n8609, ZN => n3118);
   U7815 : NAND2_X1 port map( A1 => n17440, A2 => n765, ZN => n15112);
   U7818 : OAI21_X1 port map( A1 => n9776, A2 => n23105, B => n14917, ZN => 
                           n9775);
   U7825 : NAND2_X1 port map( A1 => n24419, A2 => n12882, ZN => n4770);
   U7846 : NAND2_X1 port map( A1 => n17503, A2 => n1233, ZN => n1350);
   U7854 : NOR2_X1 port map( A1 => n26213, A2 => n27959, ZN => n5093);
   U7863 : NOR2_X1 port map( A1 => n17565, A2 => n13230, ZN => n9766);
   U7869 : NAND2_X1 port map( A1 => n10559, A2 => n14509, ZN => n10160);
   U7875 : OR2_X1 port map( A1 => n17342, A2 => n24214, Z => n7716);
   U7878 : AND3_X1 port map( A1 => n17335, A2 => n10539, A3 => n7361, Z => 
                           n13480);
   U7882 : NAND2_X1 port map( A1 => n6370, A2 => n24566, ZN => n6369);
   U7885 : OR2_X1 port map( A1 => n5500, A2 => n17315, Z => n17316);
   U7887 : AND2_X1 port map( A1 => n17337, A2 => n17335, Z => n7621);
   U7893 : OAI21_X1 port map( A1 => n13230, A2 => n10539, B => n17335, ZN => 
                           n17182);
   U7894 : NAND3_X1 port map( A1 => n26161, A2 => n3875, A3 => n17569, ZN => 
                           n3018);
   U7896 : NAND2_X1 port map( A1 => n17569, A2 => n615, ZN => n4172);
   U7901 : NOR2_X1 port map( A1 => n4415, A2 => n17558, ZN => n4417);
   U7906 : AND2_X1 port map( A1 => n17230, A2 => n17495, Z => n3147);
   U7913 : INV_X1 port map( I => n17250, ZN => n1223);
   U7914 : NOR2_X1 port map( A1 => n17036, A2 => n17204, ZN => n1951);
   U7921 : INV_X1 port map( I => n17336, ZN => n13230);
   U7926 : BUF_X2 port map( I => n16972, Z => n17181);
   U7930 : NOR2_X1 port map( A1 => n6624, A2 => n5516, ZN => n6762);
   U7932 : INV_X2 port map( I => n6625, ZN => n17318);
   U7938 : INV_X1 port map( I => n17293, ZN => n14762);
   U7941 : INV_X1 port map( I => n17003, ZN => n17454);
   U7948 : INV_X1 port map( I => n16862, ZN => n16861);
   U7951 : NAND2_X1 port map( A1 => n7046, A2 => n1242, ZN => n3144);
   U7955 : INV_X1 port map( I => n23641, ZN => n4958);
   U7956 : NAND2_X1 port map( A1 => n7092, A2 => n7091, ZN => n13140);
   U7959 : NOR2_X1 port map( A1 => n16532, A2 => n8901, ZN => n13953);
   U7962 : AOI21_X1 port map( A1 => n16736, A2 => n10281, B => n14968, ZN => 
                           n10280);
   U7967 : INV_X1 port map( I => n2576, ZN => n2573);
   U7968 : INV_X1 port map( I => n11597, ZN => n10192);
   U7969 : NAND2_X1 port map( A1 => n2576, A2 => n14620, ZN => n2575);
   U7975 : NAND2_X1 port map( A1 => n22572, A2 => n7542, ZN => n7541);
   U7978 : NAND2_X1 port map( A1 => n1042, A2 => n793, ZN => n16532);
   U7979 : NAND2_X1 port map( A1 => n7432, A2 => n7429, ZN => n7428);
   U7984 : NAND3_X1 port map( A1 => n11383, A2 => n16336, A3 => n7688, ZN => 
                           n6978);
   U7988 : AND3_X1 port map( A1 => n16559, A2 => n8199, A3 => n16558, Z => 
                           n10599);
   U7990 : NOR2_X1 port map( A1 => n16689, A2 => n7180, ZN => n6396);
   U7993 : NOR2_X1 port map( A1 => n16575, A2 => n16572, ZN => n1759);
   U7996 : OAI22_X1 port map( A1 => n16415, A2 => n6373, B1 => n10304, B2 => 
                           n16414, ZN => n16416);
   U8007 : NOR2_X1 port map( A1 => n16658, A2 => n28400, ZN => n9754);
   U8011 : AOI21_X1 port map( A1 => n3914, A2 => n12647, B => n16604, ZN => 
                           n15437);
   U8013 : NAND2_X1 port map( A1 => n16813, A2 => n12224, ZN => n12881);
   U8014 : NAND2_X1 port map( A1 => n16469, A2 => n16702, ZN => n15420);
   U8017 : NAND2_X1 port map( A1 => n14165, A2 => n23744, ZN => n2754);
   U8020 : OR2_X1 port map( A1 => n15061, A2 => n11137, Z => n16359);
   U8021 : NOR2_X1 port map( A1 => n7113, A2 => n23758, ZN => n7047);
   U8028 : NAND2_X1 port map( A1 => n905, A2 => n8223, ZN => n2578);
   U8038 : NAND2_X1 port map( A1 => n7395, A2 => n16525, ZN => n4840);
   U8041 : NAND2_X1 port map( A1 => n1251, A2 => n11224, ZN => n7091);
   U8042 : NAND3_X1 port map( A1 => n11005, A2 => n16632, A3 => n5062, ZN => 
                           n16372);
   U8047 : AND2_X1 port map( A1 => n6815, A2 => n4940, Z => n4939);
   U8053 : NAND2_X1 port map( A1 => n16498, A2 => n7668, ZN => n16500);
   U8054 : INV_X1 port map( I => n16578, ZN => n7647);
   U8057 : NAND2_X1 port map( A1 => n5777, A2 => n5776, ZN => n5775);
   U8059 : INV_X1 port map( I => n8223, ZN => n7805);
   U8060 : NOR2_X1 port map( A1 => n16702, A2 => n4295, ZN => n4575);
   U8061 : NOR2_X1 port map( A1 => n25415, A2 => n1251, ZN => n7691);
   U8062 : AOI21_X1 port map( A1 => n16645, A2 => n16644, B => n1681, ZN => 
                           n6049);
   U8064 : NAND2_X1 port map( A1 => n11504, A2 => n16433, ZN => n10156);
   U8072 : NAND2_X1 port map( A1 => n4737, A2 => n16810, ZN => n1597);
   U8086 : NOR2_X1 port map( A1 => n26814, A2 => n5861, ZN => n15571);
   U8088 : OR3_X1 port map( A1 => n25487, A2 => n22510, A3 => n16469, Z => 
                           n14028);
   U8089 : NAND2_X1 port map( A1 => n5324, A2 => n479, ZN => n5265);
   U8090 : NAND2_X1 port map( A1 => n5310, A2 => n28113, ZN => n15951);
   U8095 : NAND2_X1 port map( A1 => n16535, A2 => n9484, ZN => n5777);
   U8098 : AND2_X1 port map( A1 => n10868, A2 => n16468, Z => n3629);
   U8099 : NOR2_X1 port map( A1 => n22529, A2 => n913, ZN => n11342);
   U8102 : NAND2_X1 port map( A1 => n26760, A2 => n3537, ZN => n8250);
   U8110 : NAND2_X1 port map( A1 => n12726, A2 => n16707, ZN => n4867);
   U8117 : NAND2_X1 port map( A1 => n16639, A2 => n16640, ZN => n4596);
   U8118 : INV_X1 port map( I => n24552, ZN => n16444);
   U8119 : INV_X2 port map( I => n13039, ZN => n1253);
   U8121 : INV_X1 port map( I => n15239, ZN => n15536);
   U8130 : NAND2_X1 port map( A1 => n16105, A2 => n1263, ZN => n7227);
   U8132 : INV_X2 port map( I => n11819, ZN => n10422);
   U8133 : AOI21_X1 port map( A1 => n6122, A2 => n6120, B => n16112, ZN => 
                           n6119);
   U8140 : NOR2_X1 port map( A1 => n11223, A2 => n16335, ZN => n9706);
   U8143 : OAI21_X1 port map( A1 => n7300, A2 => n3773, B => n3770, ZN => n3769
                           );
   U8144 : INV_X2 port map( I => n16426, ZN => n16557);
   U8145 : NAND2_X1 port map( A1 => n16313, A2 => n9768, ZN => n13186);
   U8153 : OAI22_X1 port map( A1 => n16157, A2 => n25135, B1 => n16156, B2 => 
                           n6122, ZN => n16162);
   U8154 : NAND2_X1 port map( A1 => n12560, A2 => n1931, ZN => n1930);
   U8158 : NAND2_X1 port map( A1 => n16275, A2 => n13562, ZN => n7427);
   U8164 : OAI21_X1 port map( A1 => n12628, A2 => n6605, B => n5050, ZN => 
                           n2661);
   U8166 : NAND2_X1 port map( A1 => n13776, A2 => n796, ZN => n9084);
   U8177 : AND2_X1 port map( A1 => n15994, A2 => n14512, Z => n16001);
   U8178 : NAND2_X1 port map( A1 => n7869, A2 => n11628, ZN => n7407);
   U8185 : NOR2_X1 port map( A1 => n2654, A2 => n15904, ZN => n12628);
   U8189 : OAI21_X1 port map( A1 => n16069, A2 => n24702, B => n14142, ZN => 
                           n7630);
   U8193 : NAND2_X1 port map( A1 => n16186, A2 => n13533, ZN => n7162);
   U8194 : NOR2_X1 port map( A1 => n12507, A2 => n16280, ZN => n15852);
   U8196 : AOI21_X1 port map( A1 => n16270, A2 => n16271, B => n16269, ZN => 
                           n3260);
   U8199 : AOI21_X1 port map( A1 => n13577, A2 => n14763, B => n14142, ZN => 
                           n14277);
   U8200 : NOR2_X1 port map( A1 => n16112, A2 => n16321, ZN => n13582);
   U8202 : AND2_X1 port map( A1 => n15797, A2 => n21786, Z => n11909);
   U8204 : NAND2_X1 port map( A1 => n16269, A2 => n5853, ZN => n8212);
   U8206 : AOI21_X1 port map( A1 => n16269, A2 => n23104, B => n21786, ZN => 
                           n10367);
   U8209 : OAI21_X1 port map( A1 => n5569, A2 => n15756, B => n24485, ZN => 
                           n1840);
   U8211 : NOR2_X1 port map( A1 => n16353, A2 => n3735, ZN => n5668);
   U8212 : NOR2_X1 port map( A1 => n1267, A2 => n7374, ZN => n9205);
   U8213 : NOR2_X1 port map( A1 => n15946, A2 => n836, ZN => n15262);
   U8215 : NOR2_X1 port map( A1 => n8925, A2 => n16120, ZN => n9259);
   U8216 : NAND2_X1 port map( A1 => n9095, A2 => n27162, ZN => n6121);
   U8220 : NOR2_X1 port map( A1 => n7270, A2 => n5095, ZN => n15768);
   U8222 : AND2_X1 port map( A1 => n1261, A2 => n1268, Z => n2626);
   U8228 : AOI21_X1 port map( A1 => n9526, A2 => n28166, B => n15615, ZN => 
                           n9439);
   U8233 : NAND2_X1 port map( A1 => n16163, A2 => n1260, ZN => n8580);
   U8237 : NAND2_X1 port map( A1 => n1262, A2 => n16140, ZN => n9263);
   U8239 : NAND2_X1 port map( A1 => n16320, A2 => n16317, ZN => n9100);
   U8242 : INV_X1 port map( I => n21873, ZN => n9204);
   U8243 : NOR2_X1 port map( A1 => n7536, A2 => n16226, ZN => n7071);
   U8245 : NAND2_X1 port map( A1 => n15822, A2 => n14306, ZN => n4379);
   U8247 : INV_X1 port map( I => n16280, ZN => n16282);
   U8249 : AND2_X1 port map( A1 => n21787, A2 => n16283, Z => n14346);
   U8250 : NAND2_X1 port map( A1 => n24485, A2 => n10303, ZN => n1472);
   U8253 : INV_X1 port map( I => n16321, ZN => n2558);
   U8261 : NOR2_X1 port map( A1 => n16130, A2 => n4485, ZN => n15840);
   U8262 : NAND2_X1 port map( A1 => n16189, A2 => n3298, ZN => n6359);
   U8276 : NOR2_X1 port map( A1 => n7608, A2 => n6886, ZN => n10177);
   U8278 : NOR2_X1 port map( A1 => n12528, A2 => n14306, ZN => n4115);
   U8283 : INV_X1 port map( I => n20369, ZN => n1297);
   U8284 : BUF_X2 port map( I => n15905, Z => n11080);
   U8286 : INV_X1 port map( I => n21732, ZN => n1289);
   U8287 : INV_X1 port map( I => n20683, ZN => n1275);
   U8289 : INV_X1 port map( I => n14591, ZN => n1306);
   U8290 : INV_X1 port map( I => n20607, ZN => n1295);
   U8292 : INV_X1 port map( I => n21733, ZN => n1302);
   U8293 : INV_X1 port map( I => n20766, ZN => n1318);
   U8296 : INV_X1 port map( I => n15980, ZN => n15925);
   U8298 : INV_X1 port map( I => n20871, ZN => n1293);
   U8300 : INV_X1 port map( I => n20906, ZN => n1317);
   U8301 : INV_X1 port map( I => n21164, ZN => n1310);
   U8302 : INV_X1 port map( I => n20877, ZN => n1288);
   U8305 : INV_X1 port map( I => n2799, ZN => n16354);
   U8306 : BUF_X2 port map( I => n14607, Z => n7460);
   U8308 : INV_X1 port map( I => n14607, ZN => n14415);
   U8309 : INV_X2 port map( I => n5333, ZN => n7608);
   U8313 : INV_X1 port map( I => n14621, ZN => n1300);
   U8314 : INV_X1 port map( I => n21288, ZN => n1291);
   U8316 : INV_X1 port map( I => n20467, ZN => n1319);
   U8317 : INV_X1 port map( I => n14555, ZN => n1311);
   U8318 : INV_X1 port map( I => n14405, ZN => n1290);
   U8320 : INV_X1 port map( I => n21523, ZN => n1278);
   U8321 : INV_X1 port map( I => n21341, ZN => n1296);
   U8322 : CLKBUF_X2 port map( I => Key(56), Z => n14621);
   U8324 : CLKBUF_X2 port map( I => Key(23), Z => n21482);
   U8326 : CLKBUF_X2 port map( I => Key(165), Z => n21039);
   U8327 : CLKBUF_X2 port map( I => Key(77), Z => n14609);
   U8329 : CLKBUF_X2 port map( I => Key(156), Z => n20967);
   U8330 : CLKBUF_X2 port map( I => Key(22), Z => n14604);
   U8332 : CLKBUF_X2 port map( I => Key(44), Z => n20872);
   U8334 : CLKBUF_X2 port map( I => Key(32), Z => n21597);
   U8335 : CLKBUF_X2 port map( I => Key(170), Z => n20989);
   U8336 : CLKBUF_X2 port map( I => Key(121), Z => n21594);
   U8339 : CLKBUF_X2 port map( I => Key(95), Z => n21199);
   U8340 : CLKBUF_X2 port map( I => Key(46), Z => n7362);
   U8341 : CLKBUF_X2 port map( I => Key(92), Z => n20381);
   U8342 : CLKBUF_X2 port map( I => Key(86), Z => n20906);
   U8343 : INV_X2 port map( I => n3493, ZN => n1062);
   U8344 : CLKBUF_X2 port map( I => Key(36), Z => n21712);
   U8347 : CLKBUF_X2 port map( I => Key(5), Z => n21227);
   U8348 : CLKBUF_X2 port map( I => Key(159), Z => n21449);
   U8350 : CLKBUF_X2 port map( I => Key(158), Z => n21679);
   U8351 : CLKBUF_X2 port map( I => Key(38), Z => n21164);
   U8352 : CLKBUF_X2 port map( I => Key(15), Z => n21077);
   U8357 : CLKBUF_X2 port map( I => Key(21), Z => n20766);
   U8358 : CLKBUF_X2 port map( I => Key(14), Z => n14643);
   U8361 : CLKBUF_X2 port map( I => Key(50), Z => n21732);
   U8363 : CLKBUF_X2 port map( I => Key(79), Z => n21553);
   U8364 : CLKBUF_X2 port map( I => Key(185), Z => n20707);
   U8367 : CLKBUF_X2 port map( I => Key(70), Z => n21453);
   U8368 : CLKBUF_X2 port map( I => Key(47), Z => n21288);
   U8371 : CLKBUF_X2 port map( I => Key(171), Z => n20694);
   U8373 : CLKBUF_X2 port map( I => Key(58), Z => n14518);
   U8378 : CLKBUF_X2 port map( I => Key(94), Z => n14505);
   U8381 : CLKBUF_X2 port map( I => Key(146), Z => n21106);
   U8382 : CLKBUF_X2 port map( I => Key(10), Z => n14463);
   U8383 : CLKBUF_X2 port map( I => Key(80), Z => n21216);
   U8387 : CLKBUF_X2 port map( I => Key(176), Z => n20652);
   U8390 : CLKBUF_X2 port map( I => Key(139), Z => n14576);
   U8393 : CLKBUF_X2 port map( I => Key(183), Z => n21218);
   U8396 : CLKBUF_X2 port map( I => Key(153), Z => n21733);
   U8397 : CLKBUF_X2 port map( I => Key(125), Z => n21709);
   U8400 : NAND2_X1 port map( A1 => n7527, A2 => n7526, ZN => n5303);
   U8402 : OAI21_X1 port map( A1 => n5663, A2 => n5662, B => n5658, ZN => n9229
                           );
   U8414 : AOI21_X1 port map( A1 => n21648, A2 => n11380, B => n15658, ZN => 
                           n11377);
   U8417 : AOI21_X1 port map( A1 => n4728, A2 => n4729, B => n4725, ZN => n7223
                           );
   U8428 : AOI21_X1 port map( A1 => n11147, A2 => n27375, B => n20797, ZN => 
                           n8947);
   U8430 : NAND2_X1 port map( A1 => n21040, A2 => n21041, ZN => n9423);
   U8435 : OAI21_X1 port map( A1 => n4937, A2 => n4936, B => n4935, ZN => n7336
                           );
   U8439 : INV_X1 port map( I => n21042, ZN => n5660);
   U8440 : NAND2_X1 port map( A1 => n21477, A2 => n11865, ZN => n21478);
   U8446 : NOR2_X1 port map( A1 => n13297, A2 => n21335, ZN => n14225);
   U8449 : NOR2_X1 port map( A1 => n13127, A2 => n13126, ZN => n13125);
   U8452 : AOI21_X1 port map( A1 => n937, A2 => n21005, B => n21006, ZN => 
                           n2308);
   U8456 : AND2_X1 port map( A1 => n9166, A2 => n6247, Z => n6926);
   U8459 : NOR2_X1 port map( A1 => n20795, A2 => n10477, ZN => n8946);
   U8462 : NAND2_X1 port map( A1 => n27248, A2 => n2749, ZN => n1692);
   U8464 : NOR2_X1 port map( A1 => n6433, A2 => n927, ZN => n3442);
   U8465 : NAND2_X1 port map( A1 => n22844, A2 => n21488, ZN => n7349);
   U8468 : NAND2_X1 port map( A1 => n13638, A2 => n4057, ZN => n7313);
   U8471 : AND2_X1 port map( A1 => n696, A2 => n27390, Z => n7008);
   U8472 : AND2_X1 port map( A1 => n2766, A2 => n6181, Z => n6180);
   U8476 : OAI21_X1 port map( A1 => n20846, A2 => n12407, B => n25378, ZN => 
                           n14606);
   U8477 : OAI21_X1 port map( A1 => n22789, A2 => n24574, B => n21567, ZN => 
                           n9220);
   U8479 : NAND2_X1 port map( A1 => n12728, A2 => n4851, ZN => n4850);
   U8480 : INV_X1 port map( I => n7291, ZN => n21339);
   U8481 : NAND2_X1 port map( A1 => n7443, A2 => n15026, ZN => n7442);
   U8482 : NAND3_X1 port map( A1 => n20611, A2 => n14146, A3 => n20624, ZN => 
                           n20613);
   U8483 : OAI21_X1 port map( A1 => n4892, A2 => n4891, B => n20879, ZN => 
                           n4852);
   U8486 : NAND2_X1 port map( A1 => n27407, A2 => n21739, ZN => n6897);
   U8488 : NAND2_X1 port map( A1 => n1547, A2 => n20662, ZN => n8482);
   U8491 : NAND2_X1 port map( A1 => n25307, A2 => n9493, ZN => n21215);
   U8492 : OR2_X1 port map( A1 => n20684, A2 => n7698, Z => n10410);
   U8493 : NAND2_X1 port map( A1 => n2587, A2 => n2838, ZN => n2837);
   U8495 : NOR2_X1 port map( A1 => n4345, A2 => n20917, ZN => n7441);
   U8498 : INV_X1 port map( I => n20750, ZN => n5815);
   U8499 : INV_X1 port map( I => n21114, ZN => n11587);
   U8500 : NOR2_X1 port map( A1 => n21050, A2 => n25352, ZN => n15720);
   U8501 : NAND3_X1 port map( A1 => n20618, A2 => n24597, A3 => n22766, ZN => 
                           n8585);
   U8502 : NAND2_X1 port map( A1 => n4829, A2 => n21347, ZN => n2454);
   U8509 : NAND2_X1 port map( A1 => n933, A2 => n2359, ZN => n1585);
   U8513 : INV_X1 port map( I => n9141, ZN => n5713);
   U8517 : NAND2_X1 port map( A1 => n20992, A2 => n12046, ZN => n8758);
   U8519 : AND2_X1 port map( A1 => n21409, A2 => n21413, Z => n10372);
   U8521 : AND2_X1 port map( A1 => n20963, A2 => n705, Z => n4607);
   U8522 : NOR4_X1 port map( A1 => n21166, A2 => n21163, A3 => n12191, A4 => 
                           n21162, ZN => n15655);
   U8524 : NAND2_X1 port map( A1 => n28308, A2 => n21564, ZN => n10103);
   U8529 : AND2_X1 port map( A1 => n23976, A2 => n13472, Z => n10724);
   U8535 : CLKBUF_X2 port map( I => n20626, Z => n14146);
   U8537 : NAND2_X1 port map( A1 => n10675, A2 => n12581, ZN => n5768);
   U8538 : AND2_X1 port map( A1 => n9851, A2 => n21071, Z => n9866);
   U8539 : OAI21_X1 port map( A1 => n11263, A2 => n772, B => n12172, ZN => 
                           n12171);
   U8541 : INV_X1 port map( I => n13400, ZN => n9031);
   U8543 : NAND2_X1 port map( A1 => n20746, A2 => n10610, ZN => n6408);
   U8551 : NAND2_X1 port map( A1 => n12063, A2 => n15169, ZN => n12062);
   U8555 : INV_X1 port map( I => n21028, ZN => n12060);
   U8560 : OAI21_X1 port map( A1 => n20864, A2 => n20863, B => n14183, ZN => 
                           n20870);
   U8568 : OAI21_X1 port map( A1 => n26627, A2 => n14341, B => n3790, ZN => 
                           n3789);
   U8572 : NAND2_X1 port map( A1 => n11165, A2 => n11164, ZN => n11163);
   U8582 : NOR2_X1 port map( A1 => n21137, A2 => n12287, ZN => n3362);
   U8585 : OR3_X1 port map( A1 => n13772, A2 => n27455, A3 => n21444, Z => 
                           n10551);
   U8594 : OAI21_X1 port map( A1 => n13912, A2 => n21671, B => n25829, ZN => 
                           n13310);
   U8596 : NOR2_X1 port map( A1 => n11802, A2 => n13050, ZN => n11801);
   U8602 : NOR2_X1 port map( A1 => n12129, A2 => n14806, ZN => n12128);
   U8605 : INV_X1 port map( I => n10795, ZN => n6516);
   U8609 : INV_X1 port map( I => n21726, ZN => n10405);
   U8615 : NOR2_X1 port map( A1 => n21442, A2 => n21591, ZN => n8817);
   U8617 : INV_X1 port map( I => n4513, ZN => n4512);
   U8619 : NAND2_X1 port map( A1 => n20738, A2 => n20737, ZN => n10086);
   U8621 : AND2_X1 port map( A1 => n22942, A2 => n13447, Z => n15180);
   U8626 : NAND2_X1 port map( A1 => n20889, A2 => n25841, ZN => n3044);
   U8628 : NOR2_X1 port map( A1 => n21690, A2 => n952, ZN => n5311);
   U8631 : OR3_X1 port map( A1 => n21622, A2 => n13426, A3 => n21627, Z => 
                           n21581);
   U8633 : OAI21_X1 port map( A1 => n10829, A2 => n21208, B => n21325, ZN => 
                           n3691);
   U8639 : NAND2_X1 port map( A1 => n21697, A2 => n21721, ZN => n9119);
   U8643 : NAND2_X1 port map( A1 => n3561, A2 => n3560, ZN => n1853);
   U8647 : AND2_X1 port map( A1 => n10730, A2 => n10558, Z => n21056);
   U8657 : NAND2_X1 port map( A1 => n612, A2 => n20881, ZN => n15364);
   U8658 : INV_X1 port map( I => n5367, ZN => n20862);
   U8663 : NOR2_X1 port map( A1 => n21160, A2 => n13049, ZN => n2137);
   U8668 : INV_X2 port map( I => n7706, ZN => n5367);
   U8676 : AND2_X1 port map( A1 => n7228, A2 => n12598, Z => n21021);
   U8679 : AND2_X1 port map( A1 => n20395, A2 => n20502, Z => n3820);
   U8687 : CLKBUF_X2 port map( I => n9756, Z => n9005);
   U8688 : AND2_X1 port map( A1 => n21161, A2 => n21160, Z => n10608);
   U8692 : BUF_X2 port map( I => n21728, Z => n5042);
   U8709 : INV_X1 port map( I => n20555, ZN => n5043);
   U8713 : INV_X1 port map( I => n20773, ZN => n4865);
   U8717 : INV_X1 port map( I => n21157, ZN => n4895);
   U8718 : OAI21_X1 port map( A1 => n8852, A2 => n8854, B => n21039, ZN => 
                           n8851);
   U8720 : NOR2_X1 port map( A1 => n11859, A2 => n11860, ZN => n3082);
   U8722 : INV_X1 port map( I => n20470, ZN => n1536);
   U8725 : INV_X1 port map( I => n8448, ZN => n20402);
   U8726 : NAND2_X1 port map( A1 => n4908, A2 => n4907, ZN => n4910);
   U8730 : INV_X1 port map( I => n21304, ZN => n8140);
   U8748 : OAI22_X1 port map( A1 => n3799, A2 => n20101, B1 => n28525, B2 => 
                           n3798, ZN => n19855);
   U8758 : NAND2_X1 port map( A1 => n12014, A2 => n12713, ZN => n8853);
   U8761 : OAI21_X1 port map( A1 => n956, A2 => n20271, B => n5905, ZN => n5908
                           );
   U8764 : INV_X1 port map( I => n20448, ZN => n5335);
   U8773 : NAND2_X1 port map( A1 => n11203, A2 => n26652, ZN => n7359);
   U8774 : NAND2_X1 port map( A1 => n20041, A2 => n745, ZN => n8927);
   U8780 : NAND2_X1 port map( A1 => n20413, A2 => n15320, ZN => n14185);
   U8792 : NAND2_X1 port map( A1 => n3302, A2 => n20166, ZN => n9307);
   U8797 : AOI21_X1 port map( A1 => n3060, A2 => n20245, B => n957, ZN => 
                           n15165);
   U8805 : NOR2_X1 port map( A1 => n20147, A2 => n5271, ZN => n19810);
   U8809 : NAND2_X1 port map( A1 => n12723, A2 => n1835, ZN => n12722);
   U8811 : INV_X1 port map( I => n9341, ZN => n9340);
   U8814 : NAND2_X1 port map( A1 => n1451, A2 => n9875, ZN => n1447);
   U8823 : INV_X1 port map( I => n1605, ZN => n11230);
   U8826 : NOR2_X1 port map( A1 => n25959, A2 => n27235, ZN => n4650);
   U8830 : NAND2_X1 port map( A1 => n2877, A2 => n23558, ZN => n2876);
   U8835 : NAND2_X1 port map( A1 => n13460, A2 => n20215, ZN => n9083);
   U8848 : NAND2_X1 port map( A1 => n12131, A2 => n12130, ZN => n19959);
   U8851 : OAI21_X1 port map( A1 => n2890, A2 => n20084, B => n20085, ZN => 
                           n14089);
   U8858 : INV_X1 port map( I => n20192, ZN => n19986);
   U8866 : NOR2_X1 port map( A1 => n13252, A2 => n733, ZN => n10733);
   U8869 : NOR2_X1 port map( A1 => n13429, A2 => n22815, ZN => n8477);
   U8875 : NAND2_X1 port map( A1 => n1605, A2 => n9579, ZN => n3509);
   U8877 : NAND2_X1 port map( A1 => n4858, A2 => n25045, ZN => n4857);
   U8880 : INV_X1 port map( I => n20054, ZN => n11925);
   U8885 : INV_X1 port map( I => n13269, ZN => n20271);
   U8890 : AND2_X1 port map( A1 => n9087, A2 => n260, Z => n14646);
   U8894 : AND2_X1 port map( A1 => n25795, A2 => n4311, Z => n6525);
   U8901 : NOR2_X1 port map( A1 => n22000, A2 => n20087, ZN => n12339);
   U8902 : NAND2_X1 port map( A1 => n20158, A2 => n2878, ZN => n2877);
   U8904 : NAND2_X1 port map( A1 => n20235, A2 => n1835, ZN => n6286);
   U8908 : INV_X1 port map( I => n3883, ZN => n3882);
   U8912 : NOR2_X1 port map( A1 => n8907, A2 => n8906, ZN => n8905);
   U8914 : INV_X2 port map( I => n20087, ZN => n20209);
   U8918 : AND2_X1 port map( A1 => n20190, A2 => n15732, Z => n10717);
   U8920 : AND2_X1 port map( A1 => n28091, A2 => n10221, Z => n14399);
   U8922 : NAND2_X1 port map( A1 => n20190, A2 => n15733, ZN => n2716);
   U8924 : NAND3_X1 port map( A1 => n7667, A2 => n11033, A3 => n10979, ZN => 
                           n8907);
   U8930 : NOR2_X1 port map( A1 => n7618, A2 => n7704, ZN => n7703);
   U8933 : NAND2_X1 port map( A1 => n8032, A2 => n14221, ZN => n8733);
   U8934 : NOR2_X1 port map( A1 => n13145, A2 => n22000, ZN => n12006);
   U8944 : NOR2_X1 port map( A1 => n12364, A2 => n22374, ZN => n5299);
   U8955 : NAND2_X1 port map( A1 => n4434, A2 => n14672, ZN => n4433);
   U8957 : AND2_X1 port map( A1 => n19095, A2 => n19096, Z => n8769);
   U8966 : NAND2_X1 port map( A1 => n19884, A2 => n12219, ZN => n9294);
   U8982 : NAND2_X1 port map( A1 => n8325, A2 => n977, ZN => n5503);
   U8987 : AOI21_X1 port map( A1 => n6758, A2 => n6757, B => n22422, ZN => 
                           n4563);
   U8989 : INV_X1 port map( I => n11950, ZN => n7148);
   U8995 : NAND2_X1 port map( A1 => n19770, A2 => n28134, ZN => n11237);
   U8996 : NAND2_X1 port map( A1 => n6758, A2 => n6757, ZN => n4566);
   U8998 : NAND2_X1 port map( A1 => n19577, A2 => n19919, ZN => n5291);
   U9003 : INV_X1 port map( I => n4439, ZN => n19760);
   U9006 : OAI21_X1 port map( A1 => n19758, A2 => n24997, B => n4435, ZN => 
                           n4434);
   U9010 : OR2_X1 port map( A1 => n19832, A2 => n26654, Z => n10727);
   U9012 : NAND2_X1 port map( A1 => n19694, A2 => n12512, ZN => n5785);
   U9025 : NAND2_X1 port map( A1 => n28402, A2 => n2087, ZN => n2086);
   U9032 : INV_X1 port map( I => n19635, ZN => n5315);
   U9033 : NOR2_X1 port map( A1 => n24558, A2 => n724, ZN => n8307);
   U9037 : NOR2_X1 port map( A1 => n21813, A2 => n19623, ZN => n5316);
   U9038 : AND3_X1 port map( A1 => n19843, A2 => n19842, A3 => n3584, Z => 
                           n19739);
   U9060 : INV_X1 port map( I => n11044, ZN => n10522);
   U9062 : NOR2_X1 port map( A1 => n11329, A2 => n28068, ZN => n7820);
   U9066 : NAND2_X1 port map( A1 => n11167, A2 => n4136, ZN => n2444);
   U9069 : INV_X1 port map( I => n9296, ZN => n9295);
   U9073 : INV_X1 port map( I => n2102, ZN => n2173);
   U9074 : INV_X1 port map( I => n3452, ZN => n4182);
   U9076 : NAND2_X1 port map( A1 => n24545, A2 => n22174, ZN => n5057);
   U9079 : NAND2_X1 port map( A1 => n24558, A2 => n735, ZN => n7069);
   U9086 : INV_X1 port map( I => n19711, ZN => n10096);
   U9088 : NOR2_X1 port map( A1 => n19762, A2 => n11213, ZN => n4227);
   U9089 : AND2_X1 port map( A1 => n19742, A2 => n26129, Z => n9162);
   U9091 : INV_X1 port map( I => n19820, ZN => n8119);
   U9096 : OAI21_X1 port map( A1 => n3584, A2 => n2941, B => n5331, ZN => 
                           n19738);
   U9097 : NAND2_X1 port map( A1 => n14726, A2 => n19730, ZN => n6391);
   U9099 : NAND2_X1 port map( A1 => n27588, A2 => n724, ZN => n2087);
   U9106 : NAND2_X1 port map( A1 => n19666, A2 => n2320, ZN => n19667);
   U9108 : OR2_X1 port map( A1 => n19623, A2 => n866, Z => n10745);
   U9110 : OR2_X1 port map( A1 => n19499, A2 => n10978, Z => n11132);
   U9112 : INV_X1 port map( I => n19727, ZN => n11167);
   U9113 : AOI21_X1 port map( A1 => n15618, A2 => n19895, B => n28377, ZN => 
                           n3452);
   U9116 : AND2_X1 port map( A1 => n6976, A2 => n12666, Z => n12665);
   U9118 : OR2_X1 port map( A1 => n19937, A2 => n24336, Z => n12928);
   U9126 : AND2_X1 port map( A1 => n9887, A2 => n19883, Z => n19283);
   U9127 : OR2_X1 port map( A1 => n19947, A2 => n19948, Z => n14947);
   U9135 : INV_X2 port map( I => n3940, ZN => n19899);
   U9144 : NAND2_X1 port map( A1 => n19843, A2 => n15457, ZN => n2794);
   U9146 : AND2_X1 port map( A1 => n14423, A2 => n25650, Z => n8276);
   U9153 : AND2_X1 port map( A1 => n19930, A2 => n11354, Z => n19751);
   U9156 : INV_X1 port map( I => n19757, ZN => n8255);
   U9162 : NOR2_X1 port map( A1 => n25650, A2 => n12256, ZN => n8277);
   U9165 : INV_X1 port map( I => n12286, ZN => n5889);
   U9180 : INV_X1 port map( I => n19394, ZN => n8339);
   U9184 : INV_X1 port map( I => n19469, ZN => n9594);
   U9185 : INV_X1 port map( I => n13382, ZN => n19513);
   U9189 : NAND2_X1 port map( A1 => n19213, A2 => n19212, ZN => n11549);
   U9191 : INV_X1 port map( I => n9345, ZN => n13715);
   U9192 : INV_X1 port map( I => n19315, ZN => n7304);
   U9195 : INV_X1 port map( I => n19313, ZN => n19391);
   U9202 : NOR2_X1 port map( A1 => n3054, A2 => n14181, ZN => n3053);
   U9206 : OR2_X1 port map( A1 => n14920, A2 => n14921, Z => n3469);
   U9220 : INV_X2 port map( I => n6699, ZN => n1137);
   U9228 : OR2_X1 port map( A1 => n986, A2 => n19060, Z => n10756);
   U9232 : NAND2_X1 port map( A1 => n11706, A2 => n11705, ZN => n18892);
   U9239 : OAI21_X1 port map( A1 => n13563, A2 => n23268, B => n7032, ZN => 
                           n5467);
   U9240 : NAND2_X1 port map( A1 => n9354, A2 => n18996, ZN => n12806);
   U9243 : OAI21_X1 port map( A1 => n8120, A2 => n8121, B => n14457, ZN => 
                           n7594);
   U9248 : BUF_X2 port map( I => n11552, Z => n5147);
   U9254 : NOR2_X1 port map( A1 => n11840, A2 => n9354, ZN => n9353);
   U9256 : AND2_X1 port map( A1 => n9658, A2 => n18963, Z => n6581);
   U9257 : INV_X1 port map( I => n13059, ZN => n6444);
   U9258 : NAND2_X1 port map( A1 => n18828, A2 => n2928, ZN => n2927);
   U9262 : NAND2_X1 port map( A1 => n18990, A2 => n8095, ZN => n9396);
   U9263 : NAND2_X1 port map( A1 => n5441, A2 => n11874, ZN => n3316);
   U9266 : OR2_X1 port map( A1 => n13671, A2 => n24937, Z => n8147);
   U9270 : NOR2_X1 port map( A1 => n10229, A2 => n13482, ZN => n8128);
   U9274 : INV_X1 port map( I => n8063, ZN => n19192);
   U9278 : INV_X1 port map( I => n9873, ZN => n11444);
   U9279 : NAND2_X1 port map( A1 => n18907, A2 => n19190, ZN => n11646);
   U9300 : NAND2_X1 port map( A1 => n18730, A2 => n990, ZN => n5539);
   U9301 : INV_X1 port map( I => n18984, ZN => n11706);
   U9305 : NAND2_X1 port map( A1 => n2298, A2 => n2297, ZN => n5701);
   U9312 : NAND2_X1 port map( A1 => n19089, A2 => n6906, ZN => n13764);
   U9315 : INV_X1 port map( I => n19025, ZN => n6378);
   U9331 : NAND2_X1 port map( A1 => n11486, A2 => n6999, ZN => n1441);
   U9334 : NAND2_X1 port map( A1 => n1445, A2 => n4953, ZN => n1444);
   U9336 : INV_X1 port map( I => n8802, ZN => n1817);
   U9341 : NAND2_X1 port map( A1 => n14036, A2 => n19128, ZN => n13645);
   U9344 : NOR2_X1 port map( A1 => n18829, A2 => n28491, ZN => n2928);
   U9355 : NAND2_X1 port map( A1 => n8516, A2 => n18866, ZN => n8515);
   U9356 : NAND2_X1 port map( A1 => n26631, A2 => n28303, ZN => n15620);
   U9364 : NOR2_X1 port map( A1 => n18968, A2 => n13946, ZN => n1603);
   U9369 : NAND2_X1 port map( A1 => n18576, A2 => n19124, ZN => n3238);
   U9373 : INV_X1 port map( I => n5458, ZN => n19032);
   U9382 : NOR2_X1 port map( A1 => n12667, A2 => n19045, ZN => n6217);
   U9388 : AND2_X1 port map( A1 => n992, A2 => n19057, Z => n1926);
   U9389 : NAND2_X1 port map( A1 => n2516, A2 => n12111, ZN => n12890);
   U9390 : NAND2_X1 port map( A1 => n18946, A2 => n11485, ZN => n8083);
   U9393 : NAND2_X1 port map( A1 => n11626, A2 => n19089, ZN => n9349);
   U9398 : INV_X1 port map( I => n13482, ZN => n10171);
   U9401 : NAND2_X1 port map( A1 => n12781, A2 => n18793, ZN => n18876);
   U9404 : NAND2_X1 port map( A1 => n18913, A2 => n26645, ZN => n15294);
   U9406 : INV_X2 port map( I => n13967, ZN => n1150);
   U9407 : NAND2_X1 port map( A1 => n18946, A2 => n9050, ZN => n3166);
   U9409 : NOR2_X1 port map( A1 => n26631, A2 => n18925, ZN => n18962);
   U9415 : NOR2_X1 port map( A1 => n994, A2 => n27965, ZN => n14960);
   U9417 : NOR2_X1 port map( A1 => n11388, A2 => n11387, ZN => n11386);
   U9425 : AND4_X1 port map( A1 => n18818, A2 => n18817, A3 => n18816, A4 => 
                           n18815, Z => n18819);
   U9426 : AND2_X1 port map( A1 => n7468, A2 => n18921, Z => n2256);
   U9430 : NAND2_X1 port map( A1 => n19128, A2 => n13573, ZN => n14038);
   U9436 : OAI21_X1 port map( A1 => n14300, A2 => n18546, B => n10014, ZN => 
                           n10013);
   U9440 : AOI21_X1 port map( A1 => n18769, A2 => n18768, B => n10493, ZN => 
                           n10492);
   U9442 : NAND2_X1 port map( A1 => n8745, A2 => n1014, ZN => n2745);
   U9446 : OAI21_X1 port map( A1 => n18424, A2 => n14569, B => n9600, ZN => 
                           n9599);
   U9452 : NAND2_X1 port map( A1 => n9590, A2 => n9588, ZN => n18450);
   U9462 : OAI21_X1 port map( A1 => n26031, A2 => n17732, B => n10455, ZN => 
                           n10454);
   U9463 : NOR2_X1 port map( A1 => n12424, A2 => n4391, ZN => n5585);
   U9465 : NAND2_X1 port map( A1 => n11187, A2 => n1326, ZN => n1325);
   U9467 : INV_X1 port map( I => n12682, ZN => n4038);
   U9479 : NOR2_X1 port map( A1 => n7960, A2 => n28160, ZN => n4864);
   U9486 : OR2_X1 port map( A1 => n5885, A2 => n10594, Z => n18677);
   U9498 : NAND2_X1 port map( A1 => n8944, A2 => n14649, ZN => n5881);
   U9499 : NAND2_X1 port map( A1 => n18711, A2 => n13968, ZN => n18712);
   U9500 : NAND3_X1 port map( A1 => n18721, A2 => n15660, A3 => n26292, ZN => 
                           n12773);
   U9504 : NAND2_X1 port map( A1 => n8618, A2 => n18256, ZN => n8617);
   U9514 : INV_X1 port map( I => n14808, ZN => n6650);
   U9518 : INV_X1 port map( I => n5561, ZN => n18604);
   U9520 : OAI21_X1 port map( A1 => n11919, A2 => n11382, B => n2191, ZN => 
                           n2190);
   U9521 : INV_X1 port map( I => n8619, ZN => n8618);
   U9522 : NAND2_X1 port map( A1 => n12954, A2 => n15137, ZN => n12953);
   U9525 : NAND3_X1 port map( A1 => n18454, A2 => n877, A3 => n1015, ZN => 
                           n7937);
   U9526 : NOR2_X1 port map( A1 => n1015, A2 => n18455, ZN => n6712);
   U9529 : NAND2_X1 port map( A1 => n10961, A2 => n10960, ZN => n10959);
   U9530 : NAND2_X1 port map( A1 => n1001, A2 => n18402, ZN => n10655);
   U9538 : NAND2_X1 port map( A1 => n18565, A2 => n760, ZN => n1652);
   U9548 : NAND2_X1 port map( A1 => n13369, A2 => n10930, ZN => n8281);
   U9549 : NOR2_X1 port map( A1 => n28543, A2 => n18445, ZN => n8640);
   U9552 : NAND2_X1 port map( A1 => n18510, A2 => n18532, ZN => n9590);
   U9561 : NAND2_X1 port map( A1 => n18507, A2 => n7739, ZN => n7738);
   U9562 : NOR2_X1 port map( A1 => n18461, A2 => n13564, ZN => n4960);
   U9564 : AOI21_X1 port map( A1 => n17747, A2 => n8025, B => n18667, ZN => 
                           n17748);
   U9566 : NAND2_X1 port map( A1 => n482, A2 => n12671, ZN => n6733);
   U9567 : INV_X4 port map( I => n11842, ZN => n18546);
   U9571 : NOR2_X1 port map( A1 => n8113, A2 => n6800, ZN => n11047);
   U9572 : INV_X1 port map( I => n2325, ZN => n8943);
   U9583 : AOI21_X1 port map( A1 => n7212, A2 => n27867, B => n17815, ZN => 
                           n3494);
   U9585 : NOR2_X1 port map( A1 => n3554, A2 => n25500, ZN => n7276);
   U9587 : NAND2_X1 port map( A1 => n18201, A2 => n11919, ZN => n12991);
   U9599 : NOR2_X1 port map( A1 => n457, A2 => n26639, ZN => n5098);
   U9601 : INV_X1 port map( I => n10152, ZN => n18551);
   U9605 : AOI21_X1 port map( A1 => n13210, A2 => n10297, B => n14649, ZN => 
                           n14808);
   U9613 : OR2_X1 port map( A1 => n7168, A2 => n24846, Z => n2203);
   U9619 : AND2_X1 port map( A1 => n26051, A2 => n10958, Z => n10746);
   U9623 : AND2_X1 port map( A1 => n11919, A2 => n26880, Z => n6856);
   U9625 : OR2_X1 port map( A1 => n14427, A2 => n2081, Z => n17732);
   U9626 : NOR2_X1 port map( A1 => n2081, A2 => n11262, ZN => n18481);
   U9628 : INV_X2 port map( I => n10363, ZN => n15137);
   U9629 : OR2_X1 port map( A1 => n1018, A2 => n11262, Z => n18724);
   U9630 : NAND2_X1 port map( A1 => n7960, A2 => n18445, ZN => n5656);
   U9634 : INV_X2 port map( I => n18466, ZN => n18684);
   U9641 : INV_X1 port map( I => n6144, ZN => n18743);
   U9645 : NOR2_X1 port map( A1 => n10971, A2 => n1406, ZN => n1407);
   U9648 : NAND2_X1 port map( A1 => n15423, A2 => n22832, ZN => n4091);
   U9657 : INV_X2 port map( I => n18456, ZN => n5704);
   U9663 : INV_X2 port map( I => n11261, ZN => n1190);
   U9664 : OAI21_X1 port map( A1 => n2435, A2 => n2434, B => n2436, ZN => n2433
                           );
   U9668 : INV_X2 port map( I => n18597, ZN => n1191);
   U9675 : INV_X1 port map( I => n4681, ZN => n12902);
   U9679 : INV_X1 port map( I => n1397, ZN => n18060);
   U9684 : INV_X1 port map( I => n18072, ZN => n3775);
   U9685 : INV_X1 port map( I => n18270, ZN => n14693);
   U9688 : INV_X1 port map( I => n8383, ZN => n7763);
   U9693 : INV_X1 port map( I => n27816, ZN => n18078);
   U9695 : NAND2_X1 port map( A1 => n12421, A2 => n13586, ZN => n7705);
   U9704 : INV_X1 port map( I => n17788, ZN => n4072);
   U9706 : NAND2_X1 port map( A1 => n11910, A2 => n11715, ZN => n7314);
   U9708 : INV_X1 port map( I => n5895, ZN => n5894);
   U9711 : INV_X1 port map( I => n18077, ZN => n5871);
   U9714 : INV_X1 port map( I => n13891, ZN => n18312);
   U9717 : INV_X1 port map( I => n12935, ZN => n7492);
   U9723 : AOI21_X1 port map( A1 => n12086, A2 => n21778, B => n17817, ZN => 
                           n12085);
   U9730 : INV_X1 port map( I => n17977, ZN => n4474);
   U9733 : INV_X1 port map( I => n4100, ZN => n4356);
   U9734 : NAND2_X1 port map( A1 => n10025, A2 => n12078, ZN => n3186);
   U9735 : OR2_X1 port map( A1 => n5957, A2 => n4306, Z => n4016);
   U9738 : AOI21_X1 port map( A1 => n8169, A2 => n17638, B => n885, ZN => n5895
                           );
   U9740 : NOR2_X1 port map( A1 => n25493, A2 => n25214, ZN => n10659);
   U9741 : AND2_X1 port map( A1 => n17256, A2 => n17928, Z => n4074);
   U9749 : NAND2_X1 port map( A1 => n5865, A2 => n7140, ZN => n3172);
   U9757 : OR2_X1 port map( A1 => n17681, A2 => n9480, Z => n9138);
   U9760 : NAND2_X1 port map( A1 => n17333, A2 => n17332, ZN => n6213);
   U9764 : OAI21_X1 port map( A1 => n14114, A2 => n8186, B => n25576, ZN => 
                           n8185);
   U9767 : INV_X1 port map( I => n5296, ZN => n2605);
   U9769 : OAI21_X1 port map( A1 => n1617, A2 => n2222, B => n2221, ZN => n2339
                           );
   U9771 : NOR2_X1 port map( A1 => n7017, A2 => n11579, ZN => n16971);
   U9772 : INV_X1 port map( I => n17740, ZN => n4010);
   U9788 : INV_X1 port map( I => n17774, ZN => n17775);
   U9793 : NAND2_X1 port map( A1 => n25607, A2 => n17787, ZN => n4343);
   U9795 : NAND2_X1 port map( A1 => n12334, A2 => n17929, ZN => n5394);
   U9796 : NAND3_X1 port map( A1 => n6209, A2 => n22337, A3 => n763, ZN => 
                           n6208);
   U9800 : AND3_X1 port map( A1 => n17645, A2 => n17646, A3 => n7140, Z => 
                           n6657);
   U9805 : NOR3_X1 port map( A1 => n17683, A2 => n25966, A3 => n25903, ZN => 
                           n17619);
   U9809 : NOR2_X1 port map( A1 => n17350, A2 => n17594, ZN => n12449);
   U9816 : NAND2_X1 port map( A1 => n3041, A2 => n2212, ZN => n17625);
   U9820 : AND2_X1 port map( A1 => n9691, A2 => n23110, Z => n9690);
   U9822 : NAND2_X1 port map( A1 => n11777, A2 => n5368, ZN => n3717);
   U9824 : NOR2_X1 port map( A1 => n17663, A2 => n14548, ZN => n13849);
   U9825 : OAI21_X1 port map( A1 => n11834, A2 => n18005, B => n11579, ZN => 
                           n5828);
   U9826 : NAND2_X1 port map( A1 => n9636, A2 => n11391, ZN => n17940);
   U9830 : NAND2_X1 port map( A1 => n12372, A2 => n8009, ZN => n12371);
   U9833 : NOR2_X1 port map( A1 => n443, A2 => n13389, ZN => n3289);
   U9838 : NOR2_X1 port map( A1 => n25214, A2 => n17898, ZN => n17279);
   U9839 : NOR3_X1 port map( A1 => n7781, A2 => n3146, A3 => n7784, ZN => n7823
                           );
   U9843 : AND2_X1 port map( A1 => n828, A2 => n22253, Z => n17700);
   U9855 : AOI21_X1 port map( A1 => n10800, A2 => n12022, B => n14548, ZN => 
                           n6171);
   U9857 : AND2_X1 port map( A1 => n11937, A2 => n27146, Z => n11793);
   U9862 : INV_X1 port map( I => n17761, ZN => n4504);
   U9865 : INV_X1 port map( I => n17752, ZN => n14052);
   U9868 : INV_X1 port map( I => n8888, ZN => n11777);
   U9873 : NAND2_X1 port map( A1 => n17810, A2 => n21792, ZN => n10449);
   U9875 : NAND2_X1 port map( A1 => n27068, A2 => n17752, ZN => n6169);
   U9877 : NOR2_X1 port map( A1 => n4531, A2 => n17941, ZN => n17807);
   U9887 : OR2_X1 port map( A1 => n3621, A2 => n22724, Z => n3611);
   U9893 : NAND2_X1 port map( A1 => n17959, A2 => n27074, ZN => n6965);
   U9918 : NAND2_X1 port map( A1 => n13687, A2 => n7785, ZN => n7782);
   U9920 : AND2_X1 port map( A1 => n13687, A2 => n372, Z => n3146);
   U9922 : NAND2_X1 port map( A1 => n6112, A2 => n347, ZN => n6979);
   U9933 : INV_X1 port map( I => n12455, ZN => n17441);
   U9946 : NAND2_X1 port map( A1 => n16969, A2 => n16970, ZN => n5568);
   U9960 : NAND3_X1 port map( A1 => n17533, A2 => n17531, A3 => n1035, ZN => 
                           n14772);
   U9966 : AND2_X1 port map( A1 => n9651, A2 => n896, Z => n9217);
   U9970 : NAND2_X1 port map( A1 => n7757, A2 => n6826, ZN => n4321);
   U9971 : NAND2_X1 port map( A1 => n17223, A2 => n17495, ZN => n8517);
   U9975 : AOI21_X1 port map( A1 => n14324, A2 => n10015, B => n17421, ZN => 
                           n9991);
   U9978 : INV_X1 port map( I => n4446, ZN => n15515);
   U9981 : OR2_X1 port map( A1 => n9018, A2 => n17498, Z => n17158);
   U9985 : NOR2_X1 port map( A1 => n17380, A2 => n17547, ZN => n13374);
   U9986 : NAND2_X1 port map( A1 => n13063, A2 => n1036, ZN => n5939);
   U9993 : NAND2_X1 port map( A1 => n17508, A2 => n4755, ZN => n4754);
   U9998 : NAND2_X1 port map( A1 => n17216, A2 => n11857, ZN => n2082);
   U10007 : NOR2_X1 port map( A1 => n17268, A2 => n15031, ZN => n17199);
   U10008 : INV_X1 port map( I => n2966, ZN => n17298);
   U10010 : NAND2_X1 port map( A1 => n17296, A2 => n11992, ZN => n17297);
   U10017 : AND2_X1 port map( A1 => n10082, A2 => n17454, Z => n17006);
   U10024 : AND2_X1 port map( A1 => n740, A2 => n24299, Z => n17494);
   U10029 : NOR2_X1 port map( A1 => n5978, A2 => n14578, ZN => n6198);
   U10032 : INV_X1 port map( I => n10182, ZN => n9635);
   U10041 : NOR2_X1 port map( A1 => n9975, A2 => n17403, ZN => n5346);
   U10045 : AND2_X1 port map( A1 => n17528, A2 => n17196, Z => n10771);
   U10054 : NAND3_X1 port map( A1 => n17036, A2 => n9865, A3 => n9132, ZN => 
                           n9133);
   U10055 : AND2_X1 port map( A1 => n10577, A2 => n11284, Z => n17249);
   U10057 : NAND2_X1 port map( A1 => n17485, A2 => n10559, ZN => n4819);
   U10060 : AOI21_X1 port map( A1 => n17421, A2 => n23571, B => n7370, ZN => 
                           n17271);
   U10061 : INV_X2 port map( I => n17526, ZN => n9989);
   U10067 : AND2_X1 port map( A1 => n17501, A2 => n12498, Z => n17344);
   U10069 : AND2_X1 port map( A1 => n24335, A2 => n17381, Z => n10583);
   U10071 : AND3_X1 port map( A1 => n1036, A2 => n24373, A3 => n17381, Z => 
                           n17383);
   U10077 : NAND2_X1 port map( A1 => n896, A2 => n9546, ZN => n16908);
   U10081 : OR2_X1 port map( A1 => n26363, A2 => n17447, Z => n17448);
   U10084 : INV_X1 port map( I => n17226, ZN => n16743);
   U10086 : AND2_X1 port map( A1 => n6021, A2 => n8093, Z => n9555);
   U10087 : INV_X1 port map( I => n13358, ZN => n8593);
   U10092 : NOR2_X1 port map( A1 => n898, A2 => n8094, ZN => n9546);
   U10094 : NOR2_X1 port map( A1 => n12871, A2 => n17557, ZN => n7901);
   U10095 : OR2_X1 port map( A1 => n17532, A2 => n17474, Z => n17477);
   U10098 : OR2_X1 port map( A1 => n17577, A2 => n23787, Z => n5164);
   U10101 : NOR2_X1 port map( A1 => n17556, A2 => n17557, ZN => n17222);
   U10103 : NOR2_X1 port map( A1 => n17557, A2 => n17495, ZN => n9181);
   U10115 : INV_X1 port map( I => n17454, ZN => n3376);
   U10116 : CLKBUF_X2 port map( I => n10923, Z => n7175);
   U10124 : INV_X1 port map( I => n16975, ZN => n16529);
   U10125 : INV_X1 port map( I => n17055, ZN => n15062);
   U10127 : INV_X1 port map( I => n27393, ZN => n9530);
   U10133 : NAND2_X1 port map( A1 => n2574, A2 => n2571, ZN => n16374);
   U10135 : INV_X1 port map( I => n9614, ZN => n8904);
   U10147 : INV_X1 port map( I => n12523, ZN => n6456);
   U10152 : INV_X1 port map( I => n10280, ZN => n1563);
   U10155 : INV_X1 port map( I => n16957, ZN => n8707);
   U10156 : INV_X1 port map( I => n16938, ZN => n16580);
   U10160 : INV_X1 port map( I => n27599, ZN => n10188);
   U10166 : AND2_X1 port map( A1 => n14964, A2 => n14966, Z => n7917);
   U10170 : OAI21_X1 port map( A1 => n14314, A2 => n14313, B => n11152, ZN => 
                           n9996);
   U10171 : OAI21_X1 port map( A1 => n2573, A2 => n2577, B => n2572, ZN => 
                           n2571);
   U10173 : OR2_X1 port map( A1 => n2575, A2 => n2577, Z => n2574);
   U10174 : NAND2_X1 port map( A1 => n27599, A2 => n11143, ZN => n5716);
   U10175 : AOI21_X1 port map( A1 => n8916, A2 => n8915, B => n15912, ZN => 
                           n15044);
   U10179 : AND2_X1 port map( A1 => n16635, A2 => n16636, Z => n14168);
   U10181 : NAND2_X1 port map( A1 => n4630, A2 => n4761, ZN => n16814);
   U10184 : INV_X1 port map( I => n10156, ZN => n10154);
   U10185 : INV_X1 port map( I => n8820, ZN => n10153);
   U10188 : AOI21_X1 port map( A1 => n16633, A2 => n16617, B => n14127, ZN => 
                           n14536);
   U10190 : NOR2_X1 port map( A1 => n16737, A2 => n25766, ZN => n1564);
   U10191 : OAI21_X1 port map( A1 => n7691, A2 => n7688, B => n7689, ZN => 
                           n12608);
   U10193 : INV_X1 port map( I => n10906, ZN => n4808);
   U10201 : AOI21_X1 port map( A1 => n12891, A2 => n16391, B => n24845, ZN => 
                           n2642);
   U10205 : NAND2_X1 port map( A1 => n16622, A2 => n14337, ZN => n14102);
   U10206 : INV_X1 port map( I => n11341, ZN => n9503);
   U10207 : NAND2_X1 port map( A1 => n2303, A2 => n7180, ZN => n2302);
   U10216 : AOI21_X1 port map( A1 => n7964, A2 => n7850, B => n24845, ZN => 
                           n9473);
   U10217 : INV_X1 port map( I => n7855, ZN => n2695);
   U10218 : AND2_X1 port map( A1 => n6859, A2 => n16644, Z => n9019);
   U10219 : NAND2_X1 port map( A1 => n7690, A2 => n7688, ZN => n7689);
   U10224 : OR2_X1 port map( A1 => n16443, A2 => n10597, Z => n10743);
   U10227 : OAI21_X1 port map( A1 => n16719, A2 => n16718, B => n23163, ZN => 
                           n12822);
   U10228 : INV_X1 port map( I => n8518, ZN => n10748);
   U10233 : AND2_X1 port map( A1 => n10145, A2 => n24845, Z => n2641);
   U10237 : NAND2_X1 port map( A1 => n834, A2 => n4575, ZN => n8001);
   U10243 : INV_X1 port map( I => n15437, ZN => n15436);
   U10247 : NAND2_X1 port map( A1 => n16639, A2 => n16405, ZN => n4215);
   U10248 : INV_X1 port map( I => n16621, ZN => n16622);
   U10250 : NAND2_X1 port map( A1 => n7487, A2 => n16619, ZN => n16620);
   U10251 : INV_X1 port map( I => n11343, ZN => n9502);
   U10253 : NAND2_X1 port map( A1 => n16402, A2 => n16645, ZN => n6494);
   U10258 : AND2_X1 port map( A1 => n15203, A2 => n12223, Z => n10768);
   U10264 : NAND2_X1 port map( A1 => n6859, A2 => n14632, ZN => n6955);
   U10265 : NAND2_X1 port map( A1 => n794, A2 => n9801, ZN => n9800);
   U10277 : INV_X1 port map( I => n1645, ZN => n1644);
   U10286 : NAND2_X1 port map( A1 => n913, A2 => n906, ZN => n9605);
   U10288 : OR2_X1 port map( A1 => n16813, A2 => n16810, Z => n5235);
   U10289 : INV_X1 port map( I => n4166, ZN => n16460);
   U10296 : NAND2_X1 port map( A1 => n16437, A2 => n4867, ZN => n4871);
   U10302 : NOR2_X1 port map( A1 => n10502, A2 => n1052, ZN => n9429);
   U10303 : NAND2_X1 port map( A1 => n16564, A2 => n22570, ZN => n5732);
   U10308 : NAND2_X1 port map( A1 => n24028, A2 => n6766, ZN => n6619);
   U10313 : NOR2_X1 port map( A1 => n16401, A2 => n6058, ZN => n6492);
   U10319 : AND2_X1 port map( A1 => n16461, A2 => n4162, Z => n12383);
   U10322 : NAND2_X1 port map( A1 => n16619, A2 => n16617, ZN => n12211);
   U10324 : NOR2_X1 port map( A1 => n16444, A2 => n10597, ZN => n5382);
   U10332 : NAND2_X1 port map( A1 => n11505, A2 => n11819, ZN => n12369);
   U10334 : INV_X1 port map( I => n16393, ZN => n8799);
   U10335 : INV_X1 port map( I => n16634, ZN => n14127);
   U10337 : OAI21_X1 port map( A1 => n9785, A2 => n16455, B => n16393, ZN => 
                           n10893);
   U10338 : AND2_X1 port map( A1 => n1519, A2 => n26396, Z => n14093);
   U10341 : AND2_X1 port map( A1 => n15536, A2 => n13815, Z => n4282);
   U10342 : AND2_X1 port map( A1 => n22529, A2 => n11505, Z => n11504);
   U10344 : INV_X2 port map( I => n10282, ZN => n1241);
   U10352 : INV_X1 port map( I => n16651, ZN => n9785);
   U10357 : NOR2_X1 port map( A1 => n16698, A2 => n16697, ZN => n8097);
   U10361 : INV_X2 port map( I => n11908, ZN => n16617);
   U10369 : NAND3_X1 port map( A1 => n16651, A2 => n16250, A3 => n16251, ZN => 
                           n8798);
   U10375 : NAND2_X1 port map( A1 => n8410, A2 => n11223, ZN => n2483);
   U10378 : NAND2_X1 port map( A1 => n16037, A2 => n25135, ZN => n5225);
   U10382 : INV_X1 port map( I => n15104, ZN => n14977);
   U10391 : NOR2_X1 port map( A1 => n15783, A2 => n15089, ZN => n15784);
   U10399 : NAND2_X1 port map( A1 => n10161, A2 => n1472, ZN => n3590);
   U10401 : INV_X1 port map( I => n14785, ZN => n16091);
   U10402 : INV_X1 port map( I => n10791, ZN => n3857);
   U10403 : INV_X1 port map( I => n10790, ZN => n3856);
   U10405 : AOI21_X1 port map( A1 => n719, A2 => n14107, B => n16330, ZN => 
                           n2824);
   U10408 : NAND2_X1 port map( A1 => n16229, A2 => n7124, ZN => n7123);
   U10410 : NAND2_X1 port map( A1 => n9439, A2 => n9438, ZN => n1839);
   U10414 : NAND2_X1 port map( A1 => n14884, A2 => n14108, ZN => n4557);
   U10416 : AND2_X1 port map( A1 => n10296, A2 => n16242, Z => n8686);
   U10421 : NAND2_X1 port map( A1 => n14942, A2 => n16312, ZN => n9763);
   U10423 : AOI21_X1 port map( A1 => n16142, A2 => n9263, B => n25873, ZN => 
                           n9262);
   U10424 : INV_X1 port map( I => n16242, ZN => n15089);
   U10426 : NAND2_X1 port map( A1 => n1718, A2 => n13123, ZN => n1717);
   U10428 : NAND2_X1 port map( A1 => n11396, A2 => n16350, ZN => n6845);
   U10429 : NAND2_X1 port map( A1 => n13582, A2 => n13583, ZN => n7254);
   U10432 : OAI21_X1 port map( A1 => n12509, A2 => n16320, B => n9100, ZN => 
                           n9099);
   U10433 : INV_X1 port map( I => n16157, ZN => n16037);
   U10434 : NAND2_X1 port map( A1 => n15967, A2 => n11080, ZN => n2659);
   U10440 : NAND2_X1 port map( A1 => n11289, A2 => n16282, ZN => n5000);
   U10442 : OAI21_X1 port map( A1 => n15074, A2 => n15075, B => n16316, ZN => 
                           n9562);
   U10448 : NAND2_X1 port map( A1 => n3261, A2 => n3260, ZN => n3259);
   U10452 : OAI21_X1 port map( A1 => n16259, A2 => n16262, B => n21904, ZN => 
                           n16071);
   U10454 : OAI22_X1 port map( A1 => n16074, A2 => n21904, B1 => n16262, B2 => 
                           n16073, ZN => n14657);
   U10456 : NAND2_X1 port map( A1 => n7071, A2 => n8811, ZN => n1795);
   U10461 : NAND2_X1 port map( A1 => n10176, A2 => n16206, ZN => n5178);
   U10463 : NAND2_X1 port map( A1 => n16059, A2 => n22801, ZN => n7118);
   U10464 : NAND2_X1 port map( A1 => n15814, A2 => n4346, ZN => n7628);
   U10468 : NOR2_X1 port map( A1 => n13588, A2 => n11518, ZN => n10305);
   U10469 : NAND2_X1 port map( A1 => n11755, A2 => n7630, ZN => n7629);
   U10470 : NAND2_X1 port map( A1 => n14941, A2 => n16240, ZN => n10503);
   U10471 : NAND2_X1 port map( A1 => n9595, A2 => n16167, ZN => n15939);
   U10475 : INV_X1 port map( I => n14884, ZN => n16195);
   U10478 : INV_X1 port map( I => n15611, ZN => n16028);
   U10479 : AOI21_X1 port map( A1 => n11291, A2 => n16283, B => n11290, ZN => 
                           n11289);
   U10480 : NAND2_X1 port map( A1 => n15839, A2 => n13857, ZN => n15440);
   U10481 : INV_X1 port map( I => n21216, ZN => n4698);
   U10487 : NOR2_X1 port map( A1 => n2558, A2 => n25135, ZN => n2557);
   U10488 : INV_X1 port map( I => n15975, ZN => n8603);
   U10491 : NOR2_X1 port map( A1 => n15887, A2 => n7460, ZN => n7540);
   U10492 : AND2_X1 port map( A1 => n3193, A2 => n16341, Z => n1911);
   U10493 : NOR2_X1 port map( A1 => n16257, A2 => n15497, ZN => n6857);
   U10497 : NOR2_X1 port map( A1 => n16265, A2 => n16263, ZN => n5371);
   U10500 : NAND2_X1 port map( A1 => n16332, A2 => n13417, ZN => n16039);
   U10504 : NAND2_X1 port map( A1 => n16112, A2 => n14224, ZN => n7253);
   U10507 : NAND2_X1 port map( A1 => n4114, A2 => n10813, ZN => n10793);
   U10508 : NOR2_X1 port map( A1 => n16062, A2 => n5928, ZN => n15261);
   U10511 : AOI21_X1 port map( A1 => n8926, A2 => n15960, B => n13677, ZN => 
                           n8922);
   U10514 : NAND2_X1 port map( A1 => n10001, A2 => n21786, ZN => n3261);
   U10516 : OR2_X1 port map( A1 => n16123, A2 => n12116, Z => n16124);
   U10518 : NAND3_X1 port map( A1 => n16241, A2 => n16312, A3 => n16240, ZN => 
                           n10296);
   U10519 : INV_X1 port map( I => n8812, ZN => n8811);
   U10520 : INV_X1 port map( I => n16355, ZN => n1878);
   U10521 : NOR2_X1 port map( A1 => n14442, A2 => n16244, ZN => n9432);
   U10524 : INV_X1 port map( I => n9769, ZN => n15105);
   U10526 : NAND3_X1 port map( A1 => n10269, A2 => n798, A3 => n14385, ZN => 
                           n12937);
   U10528 : NOR2_X1 port map( A1 => n15908, A2 => n9986, ZN => n10091);
   U10531 : OAI21_X1 port map( A1 => n16083, A2 => n16254, B => n16255, ZN => 
                           n5977);
   U10532 : NAND2_X1 port map( A1 => n10002, A2 => n10001, ZN => n7125);
   U10534 : NAND2_X1 port map( A1 => n10177, A2 => n5680, ZN => n5179);
   U10535 : OR2_X1 port map( A1 => n16081, A2 => n5744, Z => n5725);
   U10536 : NOR2_X1 port map( A1 => n16270, A2 => n7351, ZN => n10002);
   U10537 : CLKBUF_X2 port map( I => n16166, Z => n14218);
   U10540 : CLKBUF_X2 port map( I => n14311, Z => n14303);
   U10543 : OR2_X1 port map( A1 => n7460, A2 => n4532, Z => n4589);
   U10552 : AOI21_X1 port map( A1 => n3735, A2 => n5680, B => n16207, ZN => 
                           n3451);
   U10553 : AND2_X1 port map( A1 => n6315, A2 => n5139, Z => n3232);
   U10557 : AND2_X1 port map( A1 => n16270, A2 => n7351, Z => n14435);
   U10560 : CLKBUF_X2 port map( I => n16126, Z => n14512);
   U10567 : INV_X1 port map( I => n7368, ZN => n21635);
   U10568 : INV_X1 port map( I => n16133, ZN => n6278);
   U10572 : INV_X1 port map( I => n21649, ZN => n2158);
   U10575 : NAND2_X1 port map( A1 => n16354, A2 => n24643, ZN => n2044);
   U10576 : AND2_X1 port map( A1 => n14695, A2 => n16335, Z => n9704);
   U10577 : AND2_X1 port map( A1 => n15909, A2 => n27877, Z => n16094);
   U10578 : CLKBUF_X2 port map( I => n15957, Z => n15960);
   U10579 : CLKBUF_X2 port map( I => n15922, Z => n3262);
   U10580 : INV_X1 port map( I => n15922, ZN => n16340);
   U10581 : INV_X1 port map( I => n20621, ZN => n5601);
   U10582 : INV_X1 port map( I => n21357, ZN => n21358);
   U10583 : INV_X1 port map( I => n20433, ZN => n2517);
   U10584 : INV_X1 port map( I => n14445, ZN => n11226);
   U10590 : INV_X1 port map( I => n21642, ZN => n21643);
   U10591 : INV_X1 port map( I => n20769, ZN => n9159);
   U10592 : INV_X1 port map( I => n14638, ZN => n5596);
   U10593 : INV_X1 port map( I => n14614, ZN => n7225);
   U10596 : INV_X1 port map( I => n20908, ZN => n20909);
   U10598 : INV_X1 port map( I => n14620, ZN => n2572);
   U10599 : INV_X1 port map( I => n14610, ZN => n15503);
   U10602 : INV_X1 port map( I => n14640, ZN => n5592);
   U10604 : INV_X1 port map( I => n20872, ZN => n5734);
   U10609 : INV_X1 port map( I => n21449, ZN => n21450);
   U10610 : INV_X1 port map( I => n8648, ZN => n8684);
   U10612 : INV_X1 port map( I => n21037, ZN => n6186);
   U10613 : INV_X1 port map( I => n14526, ZN => n9512);
   U10614 : INV_X1 port map( I => n21597, ZN => n14480);
   U10616 : INV_X1 port map( I => n21210, ZN => n21211);
   U10617 : INV_X1 port map( I => n20650, ZN => n9663);
   U10621 : INV_X2 port map( I => n14814, ZN => n16283);
   U10623 : INV_X1 port map( I => n20989, ZN => n20990);
   U10626 : INV_X1 port map( I => n21218, ZN => n14782);
   U10628 : INV_X1 port map( I => n16228, ZN => n15685);
   U10629 : INV_X1 port map( I => n21422, ZN => n6289);
   U10630 : INV_X1 port map( I => n21454, ZN => n12190);
   U10631 : INV_X1 port map( I => n14404, ZN => n2423);
   U10632 : INV_X1 port map( I => n20702, ZN => n13669);
   U10634 : INV_X1 port map( I => n14622, ZN => n6381);
   U10635 : INV_X1 port map( I => n14624, ZN => n9499);
   U10636 : INV_X1 port map( I => n21077, ZN => n8091);
   U10637 : OR2_X1 port map( A1 => n16006, A2 => n11024, Z => n15882);
   U10640 : CLKBUF_X2 port map( I => Key(9), Z => n14587);
   U10641 : CLKBUF_X2 port map( I => Key(87), Z => n7365);
   U10642 : INV_X1 port map( I => n21367, ZN => n1272);
   U10645 : INV_X1 port map( I => n20617, ZN => n1274);
   U10646 : CLKBUF_X2 port map( I => Key(33), Z => n7387);
   U10647 : CLKBUF_X2 port map( I => Key(26), Z => n20671);
   U10648 : INV_X1 port map( I => n21482, ZN => n1276);
   U10650 : CLKBUF_X2 port map( I => Key(155), Z => n21170);
   U10651 : INV_X1 port map( I => Key(0), ZN => n9861);
   U10652 : CLKBUF_X2 port map( I => Key(12), Z => n14581);
   U10654 : CLKBUF_X2 port map( I => Key(2), Z => n14488);
   U10655 : INV_X1 port map( I => n21227, ZN => n1280);
   U10657 : INV_X1 port map( I => n14505, ZN => n1281);
   U10662 : INV_X1 port map( I => n14418, ZN => n1284);
   U10663 : CLKBUF_X2 port map( I => Key(110), Z => n20741);
   U10664 : INV_X1 port map( I => n21553, ZN => n1287);
   U10670 : CLKBUF_X2 port map( I => Key(17), Z => n20727);
   U10671 : CLKBUF_X2 port map( I => Key(41), Z => n14645);
   U10672 : INV_X1 port map( I => n14560, ZN => n1294);
   U10673 : CLKBUF_X2 port map( I => Key(62), Z => n21037);
   U10674 : CLKBUF_X2 port map( I => Key(147), Z => n20873);
   U10675 : CLKBUF_X2 port map( I => Key(90), Z => n14572);
   U10678 : CLKBUF_X2 port map( I => Key(83), Z => n21683);
   U10684 : INV_X1 port map( I => n21313, ZN => n1299);
   U10686 : CLKBUF_X2 port map( I => Key(152), Z => n7409);
   U10687 : INV_X1 port map( I => n21709, ZN => n1304);
   U10688 : CLKBUF_X2 port map( I => Key(64), Z => n14637);
   U10689 : CLKBUF_X2 port map( I => Key(138), Z => n14540);
   U10690 : INV_X1 port map( I => n14623, ZN => n1307);
   U10691 : CLKBUF_X2 port map( I => Key(145), Z => n7399);
   U10693 : INV_X1 port map( I => n21594, ZN => n1308);
   U10694 : CLKBUF_X2 port map( I => Key(135), Z => n21602);
   U10695 : INV_X1 port map( I => n14643, ZN => n1309);
   U10696 : CLKBUF_X2 port map( I => Key(6), Z => n14556);
   U10699 : CLKBUF_X2 port map( I => Key(167), Z => n14489);
   U10700 : INV_X1 port map( I => n21679, ZN => n1313);
   U10701 : CLKBUF_X2 port map( I => Key(8), Z => n21705);
   U10703 : INV_X1 port map( I => n14604, ZN => n1314);
   U10704 : CLKBUF_X2 port map( I => Key(168), Z => n7408);
   U10705 : CLKBUF_X2 port map( I => Key(18), Z => n14596);
   U10706 : CLKBUF_X2 port map( I => Key(20), Z => n14503);
   U10709 : CLKBUF_X2 port map( I => Key(182), Z => n21554);
   U10710 : INV_X1 port map( I => n21033, ZN => n1316);
   U10712 : CLKBUF_X2 port map( I => Key(144), Z => n14457);
   U10713 : INV_X1 port map( I => n20967, ZN => n1320);
   U10715 : INV_X2 port map( I => n1321, ZN => n12507);
   U10724 : INV_X2 port map( I => n1335, ZN => n19141);
   U10726 : OR2_X1 port map( A1 => n1335, A2 => n15187, Z => n1334);
   U10739 : NAND3_X2 port map( A1 => n6420, A2 => n10939, A3 => n10940, ZN => 
                           n12320);
   U10752 : NOR2_X2 port map( A1 => n13545, A2 => n14456, ZN => n1362);
   U10755 : XOR2_X1 port map( A1 => n19219, A2 => n19416, Z => n1363);
   U10756 : XOR2_X1 port map( A1 => n13949, A2 => n23480, Z => n19416);
   U10758 : XOR2_X1 port map( A1 => n6559, A2 => n6748, Z => n1364);
   U10764 : XOR2_X1 port map( A1 => n1370, A2 => n1367, Z => n1406);
   U10765 : XOR2_X1 port map( A1 => n1368, A2 => n1369, Z => n1367);
   U10766 : XOR2_X1 port map( A1 => n10056, A2 => n20949, Z => n1368);
   U10768 : XOR2_X1 port map( A1 => n9250, A2 => n18355, Z => n1369);
   U10772 : NAND2_X2 port map( A1 => n3814, A2 => n12370, ZN => n11787);
   U10777 : XOR2_X1 port map( A1 => n16778, A2 => n767, Z => n1372);
   U10784 : XOR2_X1 port map( A1 => n12142, A2 => n6652, Z => n20375);
   U10791 : XOR2_X1 port map( A1 => n16929, A2 => n17078, Z => n16753);
   U10799 : XOR2_X1 port map( A1 => n1397, A2 => n18171, Z => n18011);
   U10801 : XNOR2_X1 port map( A1 => Plaintext(141), A2 => Key(141), ZN => 
                           n1398);
   U10808 : INV_X2 port map( I => n1406, ZN => n13538);
   U10809 : XOR2_X1 port map( A1 => n17132, A2 => n17134, Z => n2595);
   U10815 : XOR2_X1 port map( A1 => Plaintext(92), A2 => Key(92), Z => n15916);
   U10820 : INV_X1 port map( I => n1412, ZN => n2542);
   U10821 : NAND2_X1 port map( A1 => n17576, A2 => n1228, ZN => n5166);
   U10822 : OAI21_X1 port map( A1 => n13053, A2 => n13054, B => n1228, ZN => 
                           n2592);
   U10823 : NAND2_X1 port map( A1 => n1413, A2 => n2131, ZN => n15439);
   U10825 : XOR2_X1 port map( A1 => n1420, A2 => n2999, Z => n9671);
   U10837 : XOR2_X1 port map( A1 => n1888, A2 => n3985, Z => n9699);
   U10849 : NAND2_X1 port map( A1 => n716, A2 => n22307, ZN => n2212);
   U10858 : OAI21_X1 port map( A1 => n3547, A2 => n8770, B => n1435, ZN => 
                           n14106);
   U10860 : XOR2_X1 port map( A1 => n1436, A2 => n19435, Z => n19437);
   U10861 : XOR2_X1 port map( A1 => n26496, A2 => n27362, Z => n10318);
   U10870 : INV_X1 port map( I => n11485, ZN => n1445);
   U10876 : XOR2_X1 port map( A1 => n26443, A2 => n13738, Z => n13737);
   U10880 : XOR2_X1 port map( A1 => n15443, A2 => n18062, Z => n1454);
   U10886 : NAND3_X2 port map( A1 => n9615, A2 => n16552, A3 => n1465, ZN => 
                           n11408);
   U10889 : AOI21_X1 port map( A1 => n8546, A2 => n28490, B => n14990, ZN => 
                           n1468);
   U10894 : INV_X2 port map( I => n1473, ZN => n9661);
   U10906 : XOR2_X1 port map( A1 => n25651, A2 => n14479, Z => n1489);
   U10907 : NOR2_X1 port map( A1 => n28402, A2 => n724, ZN => n10739);
   U10918 : XOR2_X1 port map( A1 => n1099, A2 => n21153, Z => n1506);
   U10920 : INV_X2 port map( I => n20059, ZN => n20225);
   U10926 : XOR2_X1 port map( A1 => n1518, A2 => n1516, Z => n13308);
   U10927 : XOR2_X1 port map( A1 => n14694, A2 => n1517, Z => n1516);
   U10928 : XOR2_X1 port map( A1 => n27437, A2 => n14621, Z => n1517);
   U10932 : AOI21_X1 port map( A1 => n16557, A2 => n1519, B => n12637, ZN => 
                           n14478);
   U10941 : XOR2_X1 port map( A1 => n13242, A2 => n1275, Z => n1525);
   U10951 : OAI22_X2 port map( A1 => n1955, A2 => n20205, B1 => n9949, B2 => 
                           n5049, ZN => n1912);
   U10953 : XOR2_X1 port map( A1 => n21386, A2 => n8885, Z => n20470);
   U10965 : NAND2_X1 port map( A1 => n4933, A2 => n1547, ZN => n4936);
   U10966 : NAND2_X2 port map( A1 => n4767, A2 => n4934, ZN => n1547);
   U10972 : INV_X2 port map( I => n1550, ZN => n4131);
   U10975 : XOR2_X1 port map( A1 => n18226, A2 => n18106, Z => n1557);
   U10982 : NOR2_X1 port map( A1 => n21863, A2 => n5573, ZN => n9343);
   U10983 : NAND3_X1 port map( A1 => n20255, A2 => n21863, A3 => n9579, ZN => 
                           n20094);
   U10984 : NOR2_X1 port map( A1 => n5577, A2 => n21863, ZN => n6253);
   U10986 : NOR2_X1 port map( A1 => n20021, A2 => n21863, ZN => n11203);
   U10990 : OAI21_X2 port map( A1 => n1568, A2 => n1570, B => n1567, ZN => 
                           n13840);
   U11004 : XOR2_X1 port map( A1 => n1582, A2 => n1313, Z => Ciphertext(175));
   U11005 : AOI21_X1 port map( A1 => n21678, A2 => n1585, B => n1583, ZN => 
                           n1582);
   U11008 : NAND2_X1 port map( A1 => n22734, A2 => n26491, ZN => n11715);
   U11014 : XOR2_X1 port map( A1 => n491, A2 => n13093, Z => n1589);
   U11015 : XOR2_X1 port map( A1 => n20776, A2 => n20060, Z => n1591);
   U11016 : XOR2_X1 port map( A1 => n21299, A2 => n22771, Z => n20060);
   U11032 : INV_X2 port map( I => n6859, ZN => n14968);
   U11033 : NAND2_X2 port map( A1 => n1616, A2 => n9020, ZN => n6859);
   U11046 : NAND2_X2 port map( A1 => n14964, A2 => n14966, ZN => n16941);
   U11052 : AOI21_X2 port map( A1 => n27580, A2 => n1632, B => n1630, ZN => 
                           n14548);
   U11053 : MUX2_X1 port map( I0 => n2960, I1 => n7055, S => n2963, Z => n1632)
                           ;
   U11059 : XOR2_X1 port map( A1 => Plaintext(35), A2 => Key(35), Z => n3493);
   U11069 : INV_X2 port map( I => n1650, ZN => n9677);
   U11071 : NAND2_X2 port map( A1 => n7904, A2 => n21020, ZN => n1650);
   U11074 : XOR2_X1 port map( A1 => n1651, A2 => n16941, Z => n16877);
   U11090 : NAND2_X2 port map( A1 => n4426, A2 => n1664, ZN => n9902);
   U11097 : XOR2_X1 port map( A1 => n21432, A2 => n1308, Z => n1667);
   U11113 : NAND2_X1 port map( A1 => n1681, A2 => n27372, ZN => n12786);
   U11119 : XOR2_X1 port map( A1 => n13661, A2 => n17014, Z => n1689);
   U11120 : XOR2_X1 port map( A1 => n12480, A2 => n19146, Z => n1876);
   U11121 : XNOR2_X1 port map( A1 => n19365, A2 => n27369, ZN => n19146);
   U11125 : XOR2_X1 port map( A1 => n1690, A2 => n1314, Z => Ciphertext(183));
   U11127 : INV_X2 port map( I => n1696, ZN => n7464);
   U11128 : NAND2_X1 port map( A1 => n20312, A2 => n2525, ZN => n11557);
   U11137 : INV_X2 port map( I => n14844, ZN => n8263);
   U11140 : NOR2_X1 port map( A1 => n999, A2 => n28019, ZN => n18416);
   U11141 : NAND2_X1 port map( A1 => n24454, A2 => n28019, ZN => n19063);
   U11142 : INV_X1 port map( I => n1703, ZN => n11980);
   U11143 : NAND2_X2 port map( A1 => n21457, A2 => n13791, ZN => n1703);
   U11152 : XOR2_X1 port map( A1 => n7279, A2 => n9096, Z => n1713);
   U11154 : AOI21_X1 port map( A1 => n14928, A2 => n21347, B => n27439, ZN => 
                           n13297);
   U11156 : XOR2_X1 port map( A1 => n491, A2 => n1280, Z => n8310);
   U11159 : NAND2_X1 port map( A1 => n782, A2 => n869, ZN => n18852);
   U11162 : INV_X2 port map( I => n16104, ZN => n7053);
   U11163 : NOR2_X1 port map( A1 => n16104, A2 => n16062, ZN => n1721);
   U11168 : XOR2_X1 port map( A1 => n1725, A2 => n11535, Z => n3688);
   U11173 : XOR2_X1 port map( A1 => n1734, A2 => n1732, Z => n14094);
   U11174 : XOR2_X1 port map( A1 => n20445, A2 => n1733, Z => n1732);
   U11175 : XOR2_X1 port map( A1 => n20912, A2 => n9161, Z => n1733);
   U11177 : XOR2_X1 port map( A1 => n12320, A2 => n11815, Z => n20445);
   U11186 : XOR2_X1 port map( A1 => n24501, A2 => n7355, Z => n1742);
   U11188 : XOR2_X1 port map( A1 => n11097, A2 => n19375, Z => n19530);
   U11193 : OAI21_X2 port map( A1 => n1758, A2 => n1757, B => n1755, ZN => 
                           n20767);
   U11202 : OAI21_X1 port map( A1 => n24397, A2 => n7599, B => n17824, ZN => 
                           n12372);
   U11209 : XOR2_X1 port map( A1 => n25000, A2 => n14540, Z => n1776);
   U11216 : NOR2_X1 port map( A1 => n9150, A2 => n1784, ZN => n1783);
   U11217 : NOR2_X1 port map( A1 => n1010, A2 => n18537, ZN => n1784);
   U11235 : OAI22_X1 port map( A1 => n15198, A2 => n26682, B1 => n14032, B2 => 
                           n15199, ZN => n15197);
   U11236 : OAI22_X1 port map( A1 => n6180, A2 => n27412, B1 => n21660, B2 => 
                           n26682, ZN => n10146);
   U11238 : INV_X1 port map( I => n21693, ZN => n8980);
   U11246 : XOR2_X1 port map( A1 => n15073, A2 => n1832, Z => n1831);
   U11247 : XOR2_X1 port map( A1 => n19312, A2 => n1304, Z => n1832);
   U11251 : XOR2_X1 port map( A1 => n19377, A2 => n9414, Z => n19184);
   U11254 : OAI21_X2 port map( A1 => n1842, A2 => n1841, B => n1840, ZN => 
                           n16629);
   U11256 : NAND2_X2 port map( A1 => n1846, A2 => n1845, ZN => n2467);
   U11262 : XOR2_X1 port map( A1 => n17032, A2 => n17090, Z => n6382);
   U11263 : XOR2_X1 port map( A1 => n17090, A2 => n20433, Z => n17010);
   U11264 : XOR2_X1 port map( A1 => n3477, A2 => n17090, Z => n17091);
   U11268 : XOR2_X1 port map( A1 => n8378, A2 => n16897, Z => n16931);
   U11275 : NOR2_X1 port map( A1 => n21087, A2 => n22796, ZN => n21072);
   U11281 : XOR2_X1 port map( A1 => n22879, A2 => n6123, Z => n18346);
   U11287 : XOR2_X1 port map( A1 => n19351, A2 => n600, Z => n1875);
   U11299 : NOR2_X1 port map( A1 => n13843, A2 => n1891, ZN => n13842);
   U11301 : NAND2_X1 port map( A1 => n1892, A2 => n17497, ZN => n17359);
   U11302 : OAI21_X1 port map( A1 => n17497, A2 => n1892, B => n3961, ZN => 
                           n17220);
   U11307 : XOR2_X1 port map( A1 => n18270, A2 => n6108, Z => n3153);
   U11309 : OR2_X1 port map( A1 => n6501, A2 => n22786, Z => n9521);
   U11320 : XOR2_X1 port map( A1 => n16932, A2 => n16389, Z => n1918);
   U11324 : OAI21_X2 port map( A1 => n1926, A2 => n1925, B => n1922, ZN => 
                           n7346);
   U11325 : OAI21_X1 port map( A1 => n180, A2 => n19057, B => n23305, ZN => 
                           n1925);
   U11338 : XOR2_X1 port map( A1 => n16988, A2 => n20584, Z => n1947);
   U11339 : NAND2_X2 port map( A1 => n1949, A2 => n17316, ZN => n4110);
   U11344 : INV_X1 port map( I => n11839, ZN => n1960);
   U11345 : XOR2_X1 port map( A1 => Plaintext(143), A2 => Key(143), Z => n16103
                           );
   U11350 : NAND2_X2 port map( A1 => n10953, A2 => n1965, ZN => n2895);
   U11353 : NOR2_X1 port map( A1 => n13563, A2 => n23060, ZN => n13549);
   U11354 : XOR2_X1 port map( A1 => n28315, A2 => n10456, Z => n9490);
   U11355 : XOR2_X1 port map( A1 => n28315, A2 => n14215, Z => n8650);
   U11366 : OAI21_X1 port map( A1 => n1982, A2 => n1048, B => n1981, ZN => 
                           n1980);
   U11370 : NAND2_X1 port map( A1 => n4750, A2 => n1987, ZN => n15790);
   U11374 : INV_X2 port map( I => n16325, ZN => n1987);
   U11376 : MUX2_X1 port map( I0 => n19748, I1 => n19153, S => n24187, Z => 
                           n1988);
   U11381 : NOR2_X1 port map( A1 => n2149, A2 => n4644, ZN => n1994);
   U11386 : INV_X2 port map( I => n1998, ZN => n17520);
   U11389 : XOR2_X1 port map( A1 => n4957, A2 => n16912, Z => n17017);
   U11396 : NAND2_X2 port map( A1 => n6695, A2 => n23700, ZN => n5213);
   U11400 : OAI21_X1 port map( A1 => n13961, A2 => n21005, B => n2007, ZN => 
                           n2425);
   U11411 : XOR2_X1 port map( A1 => n19479, A2 => n15661, Z => n2015);
   U11415 : XOR2_X1 port map( A1 => n8777, A2 => n1298, Z => n2018);
   U11424 : INV_X1 port map( I => n23575, ZN => n19121);
   U11428 : INV_X1 port map( I => n2026, ZN => n17024);
   U11429 : NAND2_X1 port map( A1 => n16550, A2 => n24028, ZN => n10518);
   U11437 : NAND2_X2 port map( A1 => n14468, A2 => n14467, ZN => n18106);
   U11441 : XOR2_X1 port map( A1 => n18227, A2 => n16961, Z => n2031);
   U11448 : NOR2_X1 port map( A1 => n907, A2 => n25336, ZN => n16625);
   U11450 : NOR2_X1 port map( A1 => n25336, A2 => n6612, ZN => n2039);
   U11452 : XOR2_X1 port map( A1 => n4994, A2 => n1235, Z => n4993);
   U11458 : INV_X2 port map( I => n2049, ZN => n5008);
   U11488 : OAI21_X1 port map( A1 => n17977, A2 => n10030, B => n2068, ZN => 
                           n12370);
   U11498 : NAND2_X2 port map( A1 => n2466, A2 => n2465, ZN => n6308);
   U11502 : AND2_X1 port map( A1 => n14583, A2 => n1068, Z => n3738);
   U11503 : XOR2_X1 port map( A1 => n28370, A2 => n1276, Z => n3777);
   U11506 : XOR2_X1 port map( A1 => n5090, A2 => n2098, Z => n5089);
   U11508 : XOR2_X1 port map( A1 => n3179, A2 => n10078, Z => n10387);
   U11512 : XOR2_X1 port map( A1 => n9650, A2 => n925, Z => n2105);
   U11518 : NOR2_X2 port map( A1 => n18890, A2 => n3053, ZN => n19447);
   U11521 : NAND2_X2 port map( A1 => n2110, A2 => n2109, ZN => n2617);
   U11523 : NAND2_X2 port map( A1 => n13956, A2 => n17023, ZN => n14826);
   U11529 : INV_X2 port map( I => n22643, ZN => n15435);
   U11533 : XOR2_X1 port map( A1 => n3810, A2 => n10018, Z => n2123);
   U11539 : XOR2_X1 port map( A1 => n2128, A2 => n2127, Z => n2126);
   U11540 : XOR2_X1 port map( A1 => n18027, A2 => n20707, Z => n2127);
   U11541 : XOR2_X1 port map( A1 => n7764, A2 => n18135, Z => n2128);
   U11542 : XOR2_X1 port map( A1 => n5420, A2 => n1299, Z => n19293);
   U11545 : NOR3_X1 port map( A1 => n1031, A2 => n24560, A3 => n17492, ZN => 
                           n2138);
   U11548 : XOR2_X1 port map( A1 => n2515, A2 => n13242, Z => n16899);
   U11549 : NAND2_X2 port map( A1 => n2299, A2 => n6348, ZN => n2515);
   U11550 : NAND3_X2 port map( A1 => n2302, A2 => n6346, A3 => n11360, ZN => 
                           n13242);
   U11555 : XOR2_X1 port map( A1 => n26922, A2 => n20912, Z => n2145);
   U11557 : NOR2_X1 port map( A1 => n2148, A2 => n23270, ZN => n10176);
   U11559 : AOI22_X1 port map( A1 => n9906, A2 => n1058, B1 => n23270, B2 => 
                           n2148, ZN => n15956);
   U11562 : XOR2_X1 port map( A1 => n2159, A2 => n2156, Z => n5919);
   U11566 : XOR2_X1 port map( A1 => n13891, A2 => n2158, Z => n2157);
   U11573 : INV_X2 port map( I => n2164, ZN => n14570);
   U11597 : XOR2_X1 port map( A1 => n17081, A2 => n2189, Z => n2188);
   U11598 : XOR2_X1 port map( A1 => n17117, A2 => n17077, Z => n2189);
   U11604 : NOR2_X1 port map( A1 => n242, A2 => n1233, ZN => n13053);
   U11605 : OAI22_X2 port map( A1 => n2195, A2 => n25015, B1 => n16194, B2 => 
                           n14989, ZN => n16286);
   U11606 : NAND2_X1 port map( A1 => n4557, A2 => n2195, ZN => n7898);
   U11607 : INV_X1 port map( I => n25003, ZN => n21009);
   U11618 : XOR2_X1 port map( A1 => n11550, A2 => n2210, Z => n5359);
   U11619 : XOR2_X1 port map( A1 => n14570, A2 => n14576, Z => n2210);
   U11622 : INV_X2 port map( I => n16538, ZN => n16611);
   U11627 : XOR2_X1 port map( A1 => n16510, A2 => n16417, Z => n2219);
   U11628 : XOR2_X1 port map( A1 => n16411, A2 => n16871, Z => n2220);
   U11629 : NAND2_X2 port map( A1 => n17310, A2 => n17309, ZN => n17722);
   U11633 : XOR2_X1 port map( A1 => n27854, A2 => n2225, Z => n9497);
   U11640 : NOR2_X1 port map( A1 => n4829, A2 => n2232, ZN => n14080);
   U11641 : XOR2_X1 port map( A1 => n2236, A2 => n2233, Z => n7972);
   U11642 : XOR2_X1 port map( A1 => n2235, A2 => n2234, Z => n2233);
   U11643 : XOR2_X1 port map( A1 => n7200, A2 => n14576, Z => n2234);
   U11649 : OAI21_X2 port map( A1 => n15816, A2 => n10643, B => n13203, ZN => 
                           n3477);
   U11650 : NOR2_X2 port map( A1 => n12942, A2 => n12537, ZN => n16950);
   U11652 : NAND2_X1 port map( A1 => n1022, A2 => n2238, ZN => n17621);
   U11659 : XOR2_X1 port map( A1 => n3574, A2 => n15547, Z => n5593);
   U11665 : NAND2_X1 port map( A1 => n14408, A2 => n2253, ZN => n18815);
   U11667 : NAND2_X1 port map( A1 => n4934, A2 => n2254, ZN => n11439);
   U11676 : XOR2_X1 port map( A1 => n8486, A2 => n2262, Z => n8490);
   U11677 : XOR2_X1 port map( A1 => n12468, A2 => n20602, Z => n2262);
   U11683 : XOR2_X1 port map( A1 => n7431, A2 => n21482, Z => n2268);
   U11690 : XOR2_X1 port map( A1 => n2273, A2 => n2729, Z => n21055);
   U11703 : NAND2_X2 port map( A1 => n15260, A2 => n15945, ZN => n13025);
   U11704 : XOR2_X1 port map( A1 => n2279, A2 => n2278, Z => n18660);
   U11705 : XOR2_X1 port map( A1 => n17811, A2 => n2985, Z => n2278);
   U11715 : XOR2_X1 port map( A1 => n17142, A2 => n2290, Z => n2351);
   U11716 : XOR2_X1 port map( A1 => n17141, A2 => n2290, Z => n4129);
   U11717 : XOR2_X1 port map( A1 => n17088, A2 => n2290, Z => n16800);
   U11720 : AOI21_X1 port map( A1 => n15679, A2 => n9115, B => n923, ZN => 
                           n2293);
   U11721 : XOR2_X1 port map( A1 => n22780, A2 => n20527, Z => n2294);
   U11724 : NAND2_X1 port map( A1 => n9376, A2 => n2820, ZN => n2297);
   U11725 : OAI21_X1 port map( A1 => n14583, A2 => n937, B => n24764, ZN => 
                           n21003);
   U11726 : XOR2_X1 port map( A1 => n2140, A2 => n14560, Z => n7833);
   U11728 : XOR2_X1 port map( A1 => n6535, A2 => n14421, Z => n8983);
   U11733 : XOR2_X1 port map( A1 => n2515, A2 => n16746, Z => n14800);
   U11734 : NOR2_X2 port map( A1 => n16222, A2 => n16223, ZN => n16746);
   U11735 : NOR2_X1 port map( A1 => n5874, A2 => n23935, ZN => n2313);
   U11739 : XOR2_X1 port map( A1 => n20714, A2 => n2319, Z => n2922);
   U11741 : XOR2_X1 port map( A1 => n2673, A2 => n663, Z => n19791);
   U11743 : OR2_X1 port map( A1 => n2939, A2 => n2322, Z => n20699);
   U11745 : AOI21_X1 port map( A1 => n27429, A2 => n20704, B => n8388, ZN => 
                           n2323);
   U11748 : NAND3_X2 port map( A1 => n7530, A2 => n2326, A3 => n3304, ZN => 
                           n18008);
   U11749 : XOR2_X1 port map( A1 => n11780, A2 => n24740, Z => n10237);
   U11751 : INV_X2 port map( I => n7382, ZN => n7910);
   U11752 : XOR2_X1 port map( A1 => Plaintext(98), A2 => Key(98), Z => n7382);
   U11753 : AND2_X1 port map( A1 => n15513, A2 => n15512, Z => n10984);
   U11760 : XOR2_X1 port map( A1 => n18180, A2 => n26486, Z => n17397);
   U11766 : XOR2_X1 port map( A1 => n10705, A2 => n2349, Z => n2348);
   U11767 : XOR2_X1 port map( A1 => n26761, A2 => n20807, Z => n2349);
   U11770 : NAND2_X2 port map( A1 => n14536, A2 => n16372, ZN => n16937);
   U11771 : XOR2_X1 port map( A1 => n8673, A2 => n2351, Z => n2350);
   U11774 : INV_X1 port map( I => n2352, ZN => n14238);
   U11775 : XOR2_X1 port map( A1 => n9123, A2 => n2352, Z => n2366);
   U11777 : XOR2_X1 port map( A1 => n20713, A2 => n2352, Z => n11964);
   U11781 : NOR2_X1 port map( A1 => n4351, A2 => n4864, ZN => n2357);
   U11783 : NAND2_X1 port map( A1 => n2359, A2 => n2800, ZN => n2812);
   U11784 : NAND3_X1 port map( A1 => n2359, A2 => n21681, A3 => n12061, ZN => 
                           n21673);
   U11787 : XOR2_X1 port map( A1 => n8309, A2 => n2361, Z => n2565);
   U11788 : XOR2_X1 port map( A1 => n23750, A2 => n20919, Z => n2361);
   U11789 : NAND2_X2 port map( A1 => n2362, A2 => n2488, ZN => n8309);
   U11790 : XOR2_X1 port map( A1 => n2363, A2 => n16762, Z => n3809);
   U11793 : NOR2_X1 port map( A1 => n945, A2 => n21719, ZN => n21698);
   U11798 : XOR2_X1 port map( A1 => n15226, A2 => n14637, Z => n2365);
   U11800 : OAI21_X2 port map( A1 => n11880, A2 => n10435, B => n3071, ZN => 
                           n10445);
   U11803 : INV_X2 port map( I => n2369, ZN => n20852);
   U11815 : NAND2_X2 port map( A1 => n5076, A2 => n9533, ZN => n17124);
   U11816 : INV_X2 port map( I => n10571, ZN => n10533);
   U11818 : XOR2_X1 port map( A1 => n18327, A2 => n2379, Z => n2378);
   U11819 : XOR2_X1 port map( A1 => n15284, A2 => n22839, Z => n2379);
   U11820 : OAI21_X2 port map( A1 => n2382, A2 => n2381, B => n2380, ZN => 
                           n19133);
   U11821 : NAND3_X1 port map( A1 => n18752, A2 => n25828, A3 => n24429, ZN => 
                           n2380);
   U11822 : AOI21_X1 port map( A1 => n18750, A2 => n1003, B => n18751, ZN => 
                           n2381);
   U11825 : NAND2_X2 port map( A1 => n7622, A2 => n7619, ZN => n15462);
   U11827 : NAND2_X1 port map( A1 => n10289, A2 => n1010, ZN => n9149);
   U11831 : OAI21_X2 port map( A1 => n11084, A2 => n11082, B => n11081, ZN => 
                           n16562);
   U11834 : OAI22_X2 port map( A1 => n3649, A2 => n3921, B1 => n3648, B2 => 
                           n17223, ZN => n10779);
   U11837 : NAND2_X1 port map( A1 => n18003, A2 => n17843, ZN => n2401);
   U11840 : XOR2_X1 port map( A1 => Plaintext(24), A2 => Key(24), Z => n2799);
   U11844 : XOR2_X1 port map( A1 => n699, A2 => n21453, Z => n2409);
   U11850 : XOR2_X1 port map( A1 => n23686, A2 => n13092, Z => n11649);
   U11852 : XOR2_X1 port map( A1 => n23686, A2 => n14573, Z => n12343);
   U11854 : NOR2_X1 port map( A1 => n102, A2 => n21111, ZN => n8544);
   U11872 : XOR2_X1 port map( A1 => n2432, A2 => n11275, Z => n2430);
   U11877 : XOR2_X1 port map( A1 => n7697, A2 => n18313, Z => n2440);
   U11885 : XOR2_X1 port map( A1 => n16887, A2 => n16830, Z => n16832);
   U11886 : XOR2_X1 port map( A1 => n27463, A2 => n2455, Z => n16887);
   U11890 : XOR2_X1 port map( A1 => n23111, A2 => n2459, Z => n2457);
   U11892 : XOR2_X1 port map( A1 => n15361, A2 => n9137, Z => n2463);
   U11903 : XOR2_X1 port map( A1 => n20537, A2 => n28502, Z => n2474);
   U11907 : INV_X2 port map( I => n2478, ZN => n18682);
   U11920 : AND2_X1 port map( A1 => n11070, A2 => n18784, Z => n2487);
   U11922 : NAND2_X2 port map( A1 => n2490, A2 => n2576, ZN => n4776);
   U11923 : AOI22_X1 port map( A1 => n9295, A2 => n2491, B1 => n9296, B2 => 
                           n19885, ZN => n8099);
   U11938 : XOR2_X1 port map( A1 => n2504, A2 => n2503, Z => n7639);
   U11939 : XOR2_X1 port map( A1 => n19405, A2 => n14645, Z => n2503);
   U11943 : XOR2_X1 port map( A1 => n2509, A2 => n8844, Z => n8838);
   U11953 : NAND2_X1 port map( A1 => n19133, A2 => n2516, ZN => n18760);
   U11955 : AOI22_X1 port map( A1 => n18970, A2 => n2516, B1 => n18971, B2 => 
                           n13573, ZN => n11267);
   U11958 : XOR2_X1 port map( A1 => n2140, A2 => n2517, Z => n8037);
   U11959 : XOR2_X1 port map( A1 => n2750, A2 => n2520, Z => n2522);
   U11962 : NOR2_X1 port map( A1 => n2524, A2 => n5368, ZN => n13848);
   U11971 : XOR2_X1 port map( A1 => n5698, A2 => n63, Z => n2528);
   U11973 : XOR2_X1 port map( A1 => n20398, A2 => n12457, Z => n2529);
   U11979 : NAND2_X2 port map( A1 => n4592, A2 => n2538, ZN => n17754);
   U11986 : NOR2_X1 port map( A1 => n9734, A2 => n2549, ZN => n5149);
   U11987 : NOR2_X1 port map( A1 => n17629, A2 => n2549, ZN => n7603);
   U11991 : XOR2_X1 port map( A1 => n2552, A2 => n2551, Z => n2689);
   U11993 : XOR2_X1 port map( A1 => n19537, A2 => n19538, Z => n2552);
   U11997 : NAND2_X2 port map( A1 => n6132, A2 => n13616, ZN => n19453);
   U11998 : NAND2_X2 port map( A1 => n5875, A2 => n6133, ZN => n9002);
   U12003 : XOR2_X1 port map( A1 => n12633, A2 => n18075, Z => n3489);
   U12005 : XOR2_X1 port map( A1 => n5525, A2 => n2565, Z => n9224);
   U12006 : NAND2_X1 port map( A1 => n17259, A2 => n10985, ZN => n2567);
   U12012 : INV_X2 port map( I => n7749, ZN => n7927);
   U12013 : NAND3_X1 port map( A1 => n23416, A2 => n23368, A3 => n20280, ZN => 
                           n13581);
   U12014 : NOR2_X1 port map( A1 => n20278, A2 => n7749, ZN => n9520);
   U12017 : INV_X1 port map( I => n16577, ZN => n2579);
   U12021 : XOR2_X1 port map( A1 => n19478, A2 => n2581, Z => n19187);
   U12026 : OAI21_X1 port map( A1 => n20911, A2 => n20910, B => n2587, ZN => 
                           n8151);
   U12032 : NOR2_X1 port map( A1 => n10251, A2 => n1001, ZN => n2594);
   U12048 : XOR2_X1 port map( A1 => n2615, A2 => n21411, Z => n4457);
   U12049 : XOR2_X1 port map( A1 => n18106, A2 => n2615, Z => n18107);
   U12050 : XOR2_X1 port map( A1 => n27145, A2 => n2615, Z => n2915);
   U12051 : XOR2_X1 port map( A1 => n18361, A2 => n2615, Z => n18363);
   U12056 : XOR2_X1 port map( A1 => n2620, A2 => n2619, Z => n2618);
   U12057 : XOR2_X1 port map( A1 => n12995, A2 => n22673, Z => n2619);
   U12060 : XOR2_X1 port map( A1 => n2621, A2 => n11974, Z => n6633);
   U12061 : XOR2_X1 port map( A1 => n2621, A2 => n5988, Z => n5987);
   U12073 : INV_X2 port map( I => n8598, ZN => n14595);
   U12074 : NAND2_X1 port map( A1 => n17349, A2 => n22724, ZN => n7110);
   U12082 : NAND2_X1 port map( A1 => n22997, A2 => n26097, ZN => n2746);
   U12087 : NAND3_X2 port map( A1 => n2950, A2 => n2947, A3 => n18551, ZN => 
                           n2647);
   U12088 : XOR2_X1 port map( A1 => n2648, A2 => n2651, Z => n4309);
   U12090 : XOR2_X1 port map( A1 => n5529, A2 => n1273, Z => n2649);
   U12092 : XOR2_X1 port map( A1 => n17967, A2 => n18163, Z => n2651);
   U12101 : XOR2_X1 port map( A1 => n2655, A2 => n12344, Z => n9724);
   U12102 : NAND2_X1 port map( A1 => n28468, A2 => n2890, ZN => n12203);
   U12110 : XOR2_X1 port map( A1 => n16875, A2 => n1302, Z => n2664);
   U12113 : XOR2_X1 port map( A1 => n9455, A2 => n8274, Z => n2667);
   U12115 : XOR2_X1 port map( A1 => n16930, A2 => n8378, Z => n2668);
   U12121 : NOR2_X1 port map( A1 => n15584, A2 => n2670, ZN => n15583);
   U12122 : OAI22_X1 port map( A1 => n27013, A2 => n2670, B1 => n4739, B2 => 
                           n11052, ZN => n20414);
   U12126 : XOR2_X1 port map( A1 => n18279, A2 => n2680, Z => n2679);
   U12127 : XOR2_X1 port map( A1 => n28148, A2 => n14564, Z => n2680);
   U12130 : XOR2_X1 port map( A1 => n18085, A2 => n18086, Z => n2681);
   U12142 : NAND2_X2 port map( A1 => n2808, A2 => n2809, ZN => n5529);
   U12144 : XOR2_X1 port map( A1 => n5718, A2 => n922, Z => n2691);
   U12148 : OAI21_X2 port map( A1 => n27463, A2 => n16818, B => n2694, ZN => 
                           n10191);
   U12150 : XOR2_X1 port map( A1 => n2700, A2 => n2697, Z => n12834);
   U12151 : XOR2_X1 port map( A1 => n2699, A2 => n2698, Z => n2697);
   U12152 : XOR2_X1 port map( A1 => n16858, A2 => n923, Z => n2698);
   U12161 : NAND2_X1 port map( A1 => n15018, A2 => n2703, ZN => n15072);
   U12169 : XOR2_X1 port map( A1 => n25383, A2 => n20614, Z => n5103);
   U12171 : XOR2_X1 port map( A1 => n15391, A2 => n25383, Z => n4878);
   U12176 : INV_X2 port map( I => n2711, ZN => n2901);
   U12177 : INV_X2 port map( I => n2712, ZN => n7269);
   U12181 : NOR2_X1 port map( A1 => n24216, A2 => n27456, ZN => n2719);
   U12188 : XOR2_X1 port map( A1 => n4197, A2 => n2904, Z => n2729);
   U12195 : NAND2_X1 port map( A1 => n4343, A2 => n47, ZN => n17788);
   U12199 : XOR2_X1 port map( A1 => n984, A2 => n24528, Z => n2743);
   U12202 : XOR2_X1 port map( A1 => n2978, A2 => n2748, Z => n2747);
   U12206 : NAND2_X2 port map( A1 => n2757, A2 => n2755, ZN => n18005);
   U12210 : INV_X1 port map( I => n2766, ZN => n3205);
   U12214 : XOR2_X1 port map( A1 => n2771, A2 => n2770, Z => n2769);
   U12216 : XNOR2_X1 port map( A1 => n5597, A2 => n18217, ZN => n18076);
   U12218 : XOR2_X1 port map( A1 => n2776, A2 => n2773, Z => n15353);
   U12219 : XOR2_X1 port map( A1 => n2775, A2 => n2774, Z => n2773);
   U12220 : XOR2_X1 port map( A1 => n9161, A2 => n1275, Z => n2774);
   U12221 : XOR2_X1 port map( A1 => n4501, A2 => n22806, Z => n2775);
   U12228 : XOR2_X1 port map( A1 => n17970, A2 => n22315, Z => n7875);
   U12236 : NAND3_X1 port map( A1 => n19843, A2 => n23748, A3 => n19878, ZN => 
                           n2791);
   U12240 : XOR2_X1 port map( A1 => n26495, A2 => n24384, Z => n2795);
   U12247 : NOR2_X1 port map( A1 => n2813, A2 => n1079, ZN => n2805);
   U12256 : NAND2_X1 port map( A1 => n2812, A2 => n933, ZN => n2811);
   U12262 : XOR2_X1 port map( A1 => n2829, A2 => n2826, Z => n20901);
   U12263 : XOR2_X1 port map( A1 => n2828, A2 => n2827, Z => n2826);
   U12264 : XOR2_X1 port map( A1 => n20488, A2 => n14564, Z => n2827);
   U12265 : XOR2_X1 port map( A1 => n21258, A2 => n20538, Z => n2828);
   U12266 : XOR2_X1 port map( A1 => n20443, A2 => n20442, Z => n2829);
   U12268 : NAND2_X1 port map( A1 => n7298, A2 => n12600, ZN => n10800);
   U12269 : NAND2_X1 port map( A1 => n12022, A2 => n7298, ZN => n8888);
   U12277 : XOR2_X1 port map( A1 => n2881, A2 => n2879, Z => n2848);
   U12278 : INV_X2 port map( I => n2848, ZN => n19400);
   U12286 : XOR2_X1 port map( A1 => n17081, A2 => n16799, Z => n2858);
   U12289 : NAND2_X1 port map( A1 => n19728, A2 => n679, ZN => n19727);
   U12290 : INV_X2 port map( I => n2864, ZN => n7228);
   U12291 : NOR2_X1 port map( A1 => n7904, A2 => n7228, ZN => n2865);
   U12295 : XOR2_X1 port map( A1 => n2871, A2 => n2872, Z => n18232);
   U12296 : XOR2_X1 port map( A1 => n18231, A2 => n14704, Z => n2872);
   U12299 : XOR2_X1 port map( A1 => n6912, A2 => n2880, Z => n2879);
   U12300 : XOR2_X1 port map( A1 => n19166, A2 => n14621, Z => n2880);
   U12306 : XOR2_X1 port map( A1 => n1098, A2 => n21435, Z => n2884);
   U12307 : XOR2_X1 port map( A1 => n21196, A2 => n2886, Z => n2885);
   U12308 : XOR2_X1 port map( A1 => n7284, A2 => n5904, Z => n2886);
   U12309 : XOR2_X1 port map( A1 => n12816, A2 => n10341, Z => n2887);
   U12317 : XOR2_X1 port map( A1 => n16780, A2 => n559, Z => n2902);
   U12319 : XOR2_X1 port map( A1 => n16988, A2 => n16862, Z => n16803);
   U12320 : XOR2_X1 port map( A1 => n12411, A2 => n10352, Z => n2904);
   U12321 : NAND2_X1 port map( A1 => n19627, A2 => n24674, ZN => n19186);
   U12333 : INV_X2 port map( I => n2919, ZN => n14997);
   U12334 : XOR2_X1 port map( A1 => n7712, A2 => n7710, Z => n2919);
   U12335 : XOR2_X1 port map( A1 => n2922, A2 => n2920, Z => n20587);
   U12336 : XOR2_X1 port map( A1 => n13071, A2 => n2921, Z => n2920);
   U12337 : XOR2_X1 port map( A1 => n21237, A2 => n21044, Z => n2921);
   U12345 : NAND2_X1 port map( A1 => n6683, A2 => n6373, ZN => n16716);
   U12348 : NAND3_X1 port map( A1 => n20693, A2 => n20695, A3 => n9563, ZN => 
                           n2936);
   U12351 : XOR2_X1 port map( A1 => n13834, A2 => n27417, Z => n20544);
   U12352 : XOR2_X1 port map( A1 => n20480, A2 => n27417, Z => n3939);
   U12353 : XOR2_X1 port map( A1 => n27418, A2 => n1272, Z => n5143);
   U12354 : XOR2_X1 port map( A1 => n11815, A2 => n27418, Z => n4258);
   U12355 : XOR2_X1 port map( A1 => n27370, A2 => n27417, Z => n11025);
   U12363 : INV_X1 port map( I => Plaintext(51), ZN => n2959);
   U12364 : XNOR2_X1 port map( A1 => n2962, A2 => n2961, ZN => n2960);
   U12365 : XOR2_X1 port map( A1 => n17024, A2 => n16745, Z => n2961);
   U12368 : XOR2_X1 port map( A1 => n17062, A2 => n9154, Z => n2965);
   U12371 : OAI22_X2 port map( A1 => n10034, A2 => n2976, B1 => n2975, B2 => 
                           n28257, ZN => n16868);
   U12373 : XOR2_X1 port map( A1 => n3862, A2 => n13118, Z => n2979);
   U12374 : OAI21_X2 port map( A1 => n16822, A2 => n13852, B => n2980, ZN => 
                           n9505);
   U12383 : XOR2_X1 port map( A1 => n10149, A2 => n1303, Z => n2985);
   U12384 : XOR2_X1 port map( A1 => n2873, A2 => n11022, Z => n2986);
   U12387 : NAND2_X2 port map( A1 => n9211, A2 => n9210, ZN => n15604);
   U12393 : XNOR2_X1 port map( A1 => n7480, A2 => n2990, ZN => n2989);
   U12394 : XOR2_X1 port map( A1 => n7280, A2 => n2991, Z => n2990);
   U12395 : XOR2_X1 port map( A1 => n18134, A2 => n9748, Z => n2991);
   U12396 : XOR2_X1 port map( A1 => n8777, A2 => n13001, Z => n4919);
   U12397 : XOR2_X1 port map( A1 => n8777, A2 => n19563, Z => n12283);
   U12398 : XOR2_X1 port map( A1 => n8777, A2 => n19451, Z => n19386);
   U12401 : XOR2_X1 port map( A1 => n2994, A2 => n14600, Z => n10018);
   U12402 : XOR2_X1 port map( A1 => n2994, A2 => n24033, Z => n7729);
   U12405 : XOR2_X1 port map( A1 => n9655, A2 => n2997, Z => n2999);
   U12406 : XOR2_X1 port map( A1 => n3868, A2 => n3001, Z => n2997);
   U12407 : INV_X1 port map( I => n1283, ZN => n3001);
   U12420 : NAND2_X1 port map( A1 => n10221, A2 => n3016, ZN => n13460);
   U12423 : INV_X2 port map( I => n3019, ZN => n7182);
   U12432 : XOR2_X1 port map( A1 => n16951, A2 => n924, Z => n3036);
   U12439 : INV_X2 port map( I => n18401, ZN => n8576);
   U12440 : NAND2_X1 port map( A1 => n27433, A2 => n18633, ZN => n7952);
   U12441 : XOR2_X1 port map( A1 => n9332, A2 => n644, Z => n18401);
   U12442 : NAND2_X1 port map( A1 => n4345, A2 => n3043, ZN => n7907);
   U12443 : NAND2_X1 port map( A1 => n12486, A2 => n22803, ZN => n3043);
   U12444 : NAND2_X2 port map( A1 => n3045, A2 => n3044, ZN => n20911);
   U12447 : NAND2_X2 port map( A1 => n9417, A2 => n10167, ZN => n5934);
   U12450 : NAND2_X1 port map( A1 => n15703, A2 => n3060, ZN => n20246);
   U12455 : NOR2_X1 port map( A1 => n6889, A2 => n6487, ZN => n6040);
   U12460 : NAND2_X2 port map( A1 => n3073, A2 => n19054, ZN => n19302);
   U12463 : XOR2_X1 port map( A1 => n12816, A2 => n14575, Z => n3078);
   U12465 : INV_X2 port map( I => n3083, ZN => n19714);
   U12466 : INV_X2 port map( I => n3084, ZN => n19468);
   U12467 : INV_X1 port map( I => n19714, ZN => n19954);
   U12476 : INV_X2 port map( I => n3105, ZN => n10904);
   U12482 : NAND2_X1 port map( A1 => n6814, A2 => n3009, ZN => n3112);
   U12483 : XOR2_X1 port map( A1 => n12279, A2 => n3115, Z => n6806);
   U12484 : XOR2_X1 port map( A1 => n5224, A2 => n8726, Z => n3115);
   U12491 : NAND2_X2 port map( A1 => n9879, A2 => n23956, ZN => n13673);
   U12494 : AND2_X1 port map( A1 => n27424, A2 => n17586, Z => n3269);
   U12499 : XOR2_X1 port map( A1 => n3665, A2 => n609, Z => n20389);
   U12509 : XOR2_X1 port map( A1 => n9914, A2 => n3128, Z => n14285);
   U12510 : XOR2_X1 port map( A1 => n9076, A2 => n10907, Z => n3128);
   U12520 : XOR2_X1 port map( A1 => n6808, A2 => n19039, Z => n3134);
   U12532 : NAND2_X2 port map( A1 => n4124, A2 => n9189, ZN => n8910);
   U12538 : XOR2_X1 port map( A1 => n18026, A2 => n18025, Z => n18649);
   U12546 : XOR2_X1 port map( A1 => n12094, A2 => n18013, Z => n18272);
   U12570 : XOR2_X1 port map( A1 => n9088, A2 => n3154, Z => n15619);
   U12571 : XOR2_X1 port map( A1 => n19415, A2 => n19416, Z => n3154);
   U12577 : OR2_X1 port map( A1 => n24552, A2 => n1052, Z => n5729);
   U12581 : INV_X2 port map( I => n3157, ZN => n3953);
   U12583 : NAND2_X2 port map( A1 => n3158, A2 => n12105, ZN => n16530);
   U12586 : NOR2_X1 port map( A1 => n16726, A2 => n16725, ZN => n3159);
   U12587 : NAND2_X1 port map( A1 => n24297, A2 => n18665, ZN => n3160);
   U12588 : XOR2_X1 port map( A1 => n17149, A2 => n17148, Z => n15360);
   U12593 : XOR2_X1 port map( A1 => n3163, A2 => n17015, Z => n12107);
   U12594 : XOR2_X1 port map( A1 => n11780, A2 => n21651, Z => n3163);
   U12598 : NAND2_X1 port map( A1 => n4990, A2 => n22623, ZN => n15965);
   U12606 : XNOR2_X1 port map( A1 => n16537, A2 => n13729, ZN => n5530);
   U12618 : NOR2_X1 port map( A1 => n10209, A2 => n17317, ZN => n3175);
   U12621 : XOR2_X1 port map( A1 => n16757, A2 => n16859, Z => n3176);
   U12626 : AND2_X1 port map( A1 => n8805, A2 => n21719, Z => n3822);
   U12627 : NAND3_X2 port map( A1 => n12132, A2 => n3182, A3 => n3181, ZN => 
                           n12612);
   U12629 : NAND2_X1 port map( A1 => n4185, A2 => n15040, ZN => n3182);
   U12634 : INV_X4 port map( I => n9450, ZN => n8265);
   U12636 : XOR2_X1 port map( A1 => Plaintext(100), A2 => Key(100), Z => n14893
                           );
   U12642 : AND2_X1 port map( A1 => n13505, A2 => n20730, Z => n3826);
   U12655 : XOR2_X1 port map( A1 => n18306, A2 => n18308, Z => n4075);
   U12656 : XOR2_X1 port map( A1 => n280, A2 => n11555, Z => n18306);
   U12659 : NOR2_X1 port map( A1 => n7251, A2 => n7041, ZN => n7040);
   U12661 : NAND2_X1 port map( A1 => n9368, A2 => n12665, ZN => n3198);
   U12662 : NAND2_X1 port map( A1 => n3516, A2 => n21290, ZN => n3515);
   U12663 : NOR2_X1 port map( A1 => n3514, A2 => n3518, ZN => n21285);
   U12665 : XOR2_X1 port map( A1 => n6559, A2 => n597, Z => n8652);
   U12670 : XOR2_X1 port map( A1 => n18938, A2 => n18937, Z => n8844);
   U12673 : OR2_X1 port map( A1 => n7030, A2 => n19191, Z => n12589);
   U12675 : NOR2_X1 port map( A1 => n10173, A2 => n6182, ZN => n3204);
   U12676 : XOR2_X1 port map( A1 => n1138, A2 => n19402, Z => n14971);
   U12686 : INV_X2 port map( I => n3216, ZN => n15454);
   U12699 : XNOR2_X1 port map( A1 => n5740, A2 => n5741, ZN => n8331);
   U12704 : INV_X1 port map( I => n4793, ZN => n11969);
   U12722 : XOR2_X1 port map( A1 => n3230, A2 => n21106, Z => Ciphertext(91));
   U12723 : NAND3_X1 port map( A1 => n15124, A2 => n21114, A3 => n21105, ZN => 
                           n3230);
   U12724 : AND2_X1 port map( A1 => n6438, A2 => n12699, Z => n3434);
   U12725 : XOR2_X1 port map( A1 => n3231, A2 => n1273, Z => Ciphertext(102));
   U12729 : XOR2_X1 port map( A1 => n3236, A2 => n3550, Z => n3410);
   U12732 : INV_X2 port map( I => n15557, ZN => n21667);
   U12733 : XOR2_X1 port map( A1 => n18016, A2 => n18202, Z => n8789);
   U12739 : NAND2_X1 port map( A1 => n13492, A2 => n27132, ZN => n9468);
   U12745 : INV_X1 port map( I => n17197, ZN => n7981);
   U12746 : NAND2_X1 port map( A1 => n15640, A2 => n12667, ZN => n6814);
   U12765 : XOR2_X1 port map( A1 => n12574, A2 => n5328, Z => n3251);
   U12772 : OAI21_X2 port map( A1 => n11909, A2 => n10367, B => n3259, ZN => 
                           n16618);
   U12787 : XOR2_X1 port map( A1 => n14800, A2 => n3268, Z => n6951);
   U12796 : XOR2_X1 port map( A1 => n11900, A2 => n15392, Z => n11899);
   U12814 : OR2_X1 port map( A1 => n23274, A2 => n21107, Z => n3293);
   U12817 : XNOR2_X1 port map( A1 => n12411, A2 => n14432, ZN => n11276);
   U12819 : NAND2_X2 port map( A1 => n4340, A2 => n4341, ZN => n20537);
   U12825 : NAND3_X1 port map( A1 => n17240, A2 => n17355, A3 => n17241, ZN => 
                           n17242);
   U12829 : XNOR2_X1 port map( A1 => n16867, A2 => n16866, ZN => n3300);
   U12841 : OR2_X1 port map( A1 => n17185, A2 => n12498, Z => n12999);
   U12862 : OAI21_X1 port map( A1 => n173, A2 => n12482, B => n5060, ZN => 
                           n5059);
   U12865 : AND2_X1 port map( A1 => n16677, A2 => n23107, Z => n6812);
   U12871 : NOR2_X1 port map( A1 => n3772, A2 => n16307, ZN => n3770);
   U12877 : OR2_X1 port map( A1 => n20917, A2 => n15026, Z => n20904);
   U12885 : XOR2_X1 port map( A1 => n14294, A2 => n22818, Z => n16788);
   U12891 : INV_X1 port map( I => n21095, ZN => n3790);
   U12895 : XNOR2_X1 port map( A1 => n19334, A2 => n14436, ZN => n4498);
   U12898 : OAI21_X1 port map( A1 => n3517, A2 => n21284, B => n3515, ZN => 
                           n3514);
   U12900 : XOR2_X1 port map( A1 => n10169, A2 => n3323, Z => n7852);
   U12908 : NAND2_X2 port map( A1 => n11148, A2 => n11150, ZN => n9899);
   U12911 : XOR2_X1 port map( A1 => n9244, A2 => n4949, Z => n4947);
   U12916 : XNOR2_X1 port map( A1 => n19282, A2 => n7529, ZN => n4018);
   U12917 : XOR2_X1 port map( A1 => n13680, A2 => n9680, Z => n9679);
   U12919 : XOR2_X1 port map( A1 => n27816, A2 => n24255, Z => n17659);
   U12941 : XOR2_X1 port map( A1 => n6500, A2 => n3338, Z => n4344);
   U12945 : XNOR2_X1 port map( A1 => n22741, A2 => n20949, ZN => n6986);
   U12956 : NAND2_X2 port map( A1 => n19973, A2 => n12897, ZN => n20773);
   U12963 : XOR2_X1 port map( A1 => n21245, A2 => n21244, Z => n3348);
   U12966 : XNOR2_X1 port map( A1 => n18203, A2 => n639, ZN => n3474);
   U12977 : XOR2_X1 port map( A1 => n8669, A2 => n8670, Z => n3355);
   U12984 : NOR2_X1 port map( A1 => n8263, A2 => n17520, ZN => n9776);
   U12996 : INV_X2 port map( I => n3363, ZN => n12340);
   U12998 : AOI21_X1 port map( A1 => n9864, A2 => n21081, B => n3364, ZN => 
                           n9862);
   U12999 : AOI21_X1 port map( A1 => n9863, A2 => n13476, B => n11923, ZN => 
                           n3364);
   U13007 : NAND2_X1 port map( A1 => n16051, A2 => n12866, ZN => n13870);
   U13010 : NAND2_X1 port map( A1 => n4609, A2 => n4608, ZN => n4613);
   U13020 : INV_X2 port map( I => n3382, ZN => n9125);
   U13023 : NAND2_X1 port map( A1 => n27235, A2 => n23916, ZN => n4654);
   U13030 : OR2_X1 port map( A1 => n21027, A2 => n7421, Z => n8010);
   U13039 : NOR2_X2 port map( A1 => n13428, A2 => n14195, ZN => n18027);
   U13040 : XOR2_X1 port map( A1 => n3707, A2 => n3392, Z => n12278);
   U13042 : NAND2_X1 port map( A1 => n8386, A2 => n7228, ZN => n20888);
   U13047 : XOR2_X1 port map( A1 => n5103, A2 => n12779, Z => n3394);
   U13063 : XOR2_X1 port map( A1 => n4193, A2 => n4194, Z => n3404);
   U13064 : XOR2_X1 port map( A1 => n16790, A2 => n16789, Z => n16972);
   U13074 : OAI22_X1 port map( A1 => n10141, A2 => n17352, B1 => n17479, B2 => 
                           n17353, ZN => n11432);
   U13075 : NOR2_X1 port map( A1 => n7102, A2 => n9635, ZN => n9634);
   U13080 : OR2_X1 port map( A1 => n21787, A2 => n16280, Z => n12866);
   U13082 : XOR2_X1 port map( A1 => n4794, A2 => n4795, Z => n18597);
   U13085 : NAND2_X1 port map( A1 => n6315, A2 => n28088, ZN => n15900);
   U13086 : INV_X2 port map( I => n3410, ZN => n21016);
   U13087 : OR2_X1 port map( A1 => n23706, A2 => n4610, Z => n4609);
   U13097 : NAND2_X2 port map( A1 => n15950, A2 => n15949, ZN => n5310);
   U13098 : OAI21_X1 port map( A1 => n15375, A2 => n6066, B => n6065, ZN => 
                           n21283);
   U13100 : INV_X2 port map( I => n3417, ZN => n11842);
   U13104 : XOR2_X1 port map( A1 => n3418, A2 => n9159, Z => Ciphertext(5));
   U13109 : XOR2_X1 port map( A1 => n3422, A2 => n20364, Z => n13325);
   U13118 : AOI21_X1 port map( A1 => n11384, A2 => n3427, B => n23919, ZN => 
                           n15205);
   U13119 : NAND2_X1 port map( A1 => n21173, A2 => n11385, ZN => n3427);
   U13120 : NAND2_X1 port map( A1 => n27469, A2 => n5680, ZN => n5637);
   U13121 : NOR2_X2 port map( A1 => n3429, A2 => n3428, ZN => n16975);
   U13125 : XOR2_X1 port map( A1 => n15109, A2 => n3432, Z => n18574);
   U13126 : XOR2_X1 port map( A1 => n15108, A2 => n17934, Z => n3432);
   U13133 : NAND2_X1 port map( A1 => n8240, A2 => n16198, ZN => n3440);
   U13137 : NAND2_X1 port map( A1 => n13545, A2 => n1270, ZN => n8240);
   U13148 : OAI21_X1 port map( A1 => n564, A2 => n3735, B => n3451, ZN => 
                           n14561);
   U13155 : NAND2_X2 port map( A1 => n10980, A2 => n10979, ZN => n20023);
   U13167 : XOR2_X1 port map( A1 => n12480, A2 => n3464, Z => n9324);
   U13188 : NOR2_X1 port map( A1 => n3851, A2 => n19110, ZN => n4077);
   U13189 : XOR2_X1 port map( A1 => n12100, A2 => n1320, Z => n4305);
   U13196 : INV_X4 port map( I => n13693, ZN => n3980);
   U13206 : INV_X2 port map( I => n3484, ZN => n3850);
   U13207 : XOR2_X1 port map( A1 => Plaintext(87), A2 => Key(87), Z => n3484);
   U13209 : NAND2_X2 port map( A1 => n3486, A2 => n10869, ZN => n10868);
   U13211 : XOR2_X1 port map( A1 => n3487, A2 => n11714, Z => n20366);
   U13215 : INV_X2 port map( I => n26638, ZN => n7612);
   U13217 : NAND2_X2 port map( A1 => n13503, A2 => n16908, ZN => n7017);
   U13218 : XOR2_X1 port map( A1 => n3491, A2 => n27589, Z => Ciphertext(114));
   U13221 : NAND2_X1 port map( A1 => n15991, A2 => n16013, ZN => n3893);
   U13225 : XOR2_X1 port map( A1 => n3501, A2 => n3499, Z => n3502);
   U13226 : XOR2_X1 port map( A1 => n24542, A2 => n9613, Z => n3499);
   U13234 : XOR2_X1 port map( A1 => n19276, A2 => n3511, Z => n3510);
   U13235 : XOR2_X1 port map( A1 => n27863, A2 => n21164, Z => n3511);
   U13239 : OAI21_X1 port map( A1 => n21286, A2 => n21279, B => n6066, ZN => 
                           n3517);
   U13244 : INV_X2 port map( I => n3527, ZN => n17546);
   U13246 : INV_X1 port map( I => n16936, ZN => n3529);
   U13251 : NAND2_X2 port map( A1 => n7325, A2 => n8387, ZN => n6821);
   U13252 : INV_X1 port map( I => n4485, ZN => n15828);
   U13253 : NAND2_X2 port map( A1 => n3570, A2 => n8580, ZN => n3537);
   U13255 : XOR2_X1 port map( A1 => n15073, A2 => n3539, Z => n3538);
   U13256 : XOR2_X1 port map( A1 => n2508, A2 => n21683, Z => n3539);
   U13257 : XOR2_X1 port map( A1 => n6308, A2 => n3541, Z => n3540);
   U13258 : XOR2_X1 port map( A1 => n19236, A2 => n2507, Z => n3541);
   U13262 : XOR2_X1 port map( A1 => n14840, A2 => n19725, Z => n3550);
   U13264 : XOR2_X1 port map( A1 => Plaintext(61), A2 => Key(61), Z => n3633);
   U13267 : XOR2_X1 port map( A1 => n25445, A2 => n27245, Z => n3556);
   U13268 : AOI21_X2 port map( A1 => n18243, A2 => n6562, B => n3557, ZN => 
                           n18128);
   U13269 : XOR2_X1 port map( A1 => n18129, A2 => n10688, Z => n3558);
   U13270 : INV_X2 port map( I => n5403, ZN => n3593);
   U13272 : INV_X2 port map( I => n3562, ZN => n8326);
   U13277 : XOR2_X1 port map( A1 => n28373, A2 => n12190, Z => n3567);
   U13279 : XOR2_X1 port map( A1 => n17037, A2 => n16869, Z => n3569);
   U13280 : XOR2_X1 port map( A1 => n7431, A2 => n16868, Z => n16869);
   U13283 : NAND2_X2 port map( A1 => n15290, A2 => n15291, ZN => n15287);
   U13284 : XOR2_X1 port map( A1 => n3575, A2 => n15730, Z => n15727);
   U13285 : XOR2_X1 port map( A1 => n23198, A2 => n22784, Z => n3575);
   U13289 : NOR2_X2 port map( A1 => n11239, A2 => n19023, ZN => n19260);
   U13290 : INV_X2 port map( I => n3579, ZN => n18639);
   U13293 : XOR2_X1 port map( A1 => n3581, A2 => n3582, Z => n3631);
   U13301 : XOR2_X1 port map( A1 => n3880, A2 => n15683, Z => n3585);
   U13303 : XOR2_X1 port map( A1 => n19549, A2 => n19262, Z => n3587);
   U13306 : INV_X2 port map( I => n3592, ZN => n20180);
   U13308 : XOR2_X1 port map( A1 => n20456, A2 => n11592, Z => n3595);
   U13315 : XOR2_X1 port map( A1 => n4288, A2 => n18206, Z => n18158);
   U13317 : AOI21_X2 port map( A1 => n17258, A2 => n17257, B => n4074, ZN => 
                           n4288);
   U13320 : XOR2_X1 port map( A1 => n7065, A2 => n14609, Z => n3602);
   U13331 : XOR2_X1 port map( A1 => n4688, A2 => n19175, Z => n3616);
   U13337 : NAND3_X1 port map( A1 => n1232, A2 => n5096, A3 => n17188, ZN => 
                           n3622);
   U13341 : INV_X2 port map( I => n3631, ZN => n7168);
   U13343 : INV_X2 port map( I => n3633, ZN => n4485);
   U13344 : XOR2_X1 port map( A1 => n26216, A2 => n4656, Z => n11102);
   U13347 : XOR2_X1 port map( A1 => n3638, A2 => n3637, Z => n3636);
   U13348 : XOR2_X1 port map( A1 => n16886, A2 => n14505, Z => n3637);
   U13349 : XOR2_X1 port map( A1 => n699, A2 => n9902, Z => n3638);
   U13361 : AOI22_X1 port map( A1 => n20754, A2 => n3650, B1 => n14242, B2 => 
                           n20740, ZN => n20742);
   U13362 : NAND2_X1 port map( A1 => n21272, A2 => n3593, ZN => n3660);
   U13363 : XOR2_X1 port map( A1 => n3663, A2 => n4943, Z => n3662);
   U13364 : XOR2_X1 port map( A1 => n25330, A2 => n20716, Z => n3664);
   U13367 : XOR2_X1 port map( A1 => n3668, A2 => n8707, Z => n3667);
   U13369 : OAI21_X1 port map( A1 => n5407, A2 => n1180, B => n4410, ZN => 
                           n4351);
   U13373 : NAND2_X2 port map( A1 => n3676, A2 => n3675, ZN => n17996);
   U13379 : XOR2_X1 port map( A1 => n7244, A2 => n22774, Z => n18152);
   U13381 : XOR2_X1 port map( A1 => n3686, A2 => n3685, Z => n3684);
   U13382 : XOR2_X1 port map( A1 => n16991, A2 => n17125, Z => n3685);
   U13389 : XOR2_X1 port map( A1 => n3701, A2 => n14535, Z => n12302);
   U13393 : XOR2_X1 port map( A1 => n3704, A2 => n3703, Z => n3702);
   U13394 : XOR2_X1 port map( A1 => n25328, A2 => n14473, Z => n3703);
   U13395 : XOR2_X1 port map( A1 => n20761, A2 => n3707, Z => n3704);
   U13401 : XNOR2_X1 port map( A1 => n12209, A2 => n2508, ZN => n19494);
   U13413 : XOR2_X1 port map( A1 => n20530, A2 => n8139, Z => n8138);
   U13414 : XNOR2_X1 port map( A1 => n20448, A2 => n20511, ZN => n20530);
   U13416 : AOI22_X2 port map( A1 => n11926, A2 => n11925, B1 => n20223, B2 => 
                           n13694, ZN => n20448);
   U13419 : MUX2_X1 port map( I0 => n16026, I1 => n16025, S => n3729, Z => 
                           n16033);
   U13420 : XOR2_X1 port map( A1 => n3734, A2 => n3731, Z => n12952);
   U13421 : XOR2_X1 port map( A1 => n3733, A2 => n3732, Z => n3731);
   U13422 : XOR2_X1 port map( A1 => n22837, A2 => n21288, Z => n3732);
   U13428 : NAND2_X1 port map( A1 => n6373, A2 => n16712, ZN => n3736);
   U13430 : INV_X2 port map( I => n3746, ZN => n20972);
   U13440 : XOR2_X1 port map( A1 => n19465, A2 => n4223, Z => n3754);
   U13443 : NOR2_X2 port map( A1 => n15313, A2 => n15312, ZN => n20704);
   U13446 : XOR2_X1 port map( A1 => n18164, A2 => n15558, Z => n3760);
   U13449 : NOR2_X1 port map( A1 => n25500, A2 => n877, ZN => n3766);
   U13454 : OAI21_X2 port map( A1 => n9222, A2 => n6917, B => n18090, ZN => 
                           n18135);
   U13460 : XOR2_X1 port map( A1 => n10029, A2 => n15669, Z => n21188);
   U13461 : XOR2_X1 port map( A1 => n10029, A2 => n14421, Z => n15403);
   U13462 : XOR2_X1 port map( A1 => n9055, A2 => n10029, Z => n6761);
   U13463 : XOR2_X1 port map( A1 => n25313, A2 => n10029, Z => n12958);
   U13470 : NAND2_X1 port map( A1 => n15717, A2 => n20288, ZN => n3798);
   U13479 : XOR2_X1 port map( A1 => n8366, A2 => n20537, Z => n20481);
   U13481 : XOR2_X1 port map( A1 => n3808, A2 => n3810, Z => n3807);
   U13482 : XOR2_X1 port map( A1 => n1593, A2 => n13859, Z => n3808);
   U13484 : XOR2_X1 port map( A1 => n20510, A2 => n20387, Z => n7808);
   U13488 : XOR2_X1 port map( A1 => n11643, A2 => n20470, Z => n3816);
   U13491 : XOR2_X1 port map( A1 => n1638, A2 => n26273, Z => n3818);
   U13496 : NAND2_X1 port map( A1 => n19759, A2 => n3835, ZN => n5571);
   U13499 : NAND2_X1 port map( A1 => n6189, A2 => n22748, ZN => n6188);
   U13503 : XOR2_X1 port map( A1 => n3840, A2 => n9080, Z => n18718);
   U13504 : OAI21_X2 port map( A1 => n5922, A2 => n17772, B => n17771, ZN => 
                           n5921);
   U13509 : XOR2_X1 port map( A1 => n337, A2 => n16862, Z => n14016);
   U13514 : XOR2_X1 port map( A1 => n4137, A2 => n20208, Z => n11071);
   U13520 : NAND2_X1 port map( A1 => n19836, A2 => n3861, ZN => n6757);
   U13524 : XNOR2_X1 port map( A1 => n19236, A2 => n19298, ZN => n3864);
   U13528 : INV_X2 port map( I => n16203, ZN => n3874);
   U13532 : INV_X2 port map( I => n3879, ZN => n15886);
   U13533 : XNOR2_X1 port map( A1 => Plaintext(75), A2 => Key(75), ZN => n3879)
                           ;
   U13544 : INV_X2 port map( I => n3895, ZN => n21020);
   U13547 : XOR2_X1 port map( A1 => n16545, A2 => n13749, Z => n3899);
   U13549 : XOR2_X1 port map( A1 => n16941, A2 => n21597, Z => n3897);
   U13550 : XOR2_X1 port map( A1 => n1593, A2 => n12481, Z => n3898);
   U13552 : XOR2_X1 port map( A1 => n8225, A2 => n18033, Z => n3900);
   U13554 : NOR2_X1 port map( A1 => n18003, A2 => n22153, ZN => n11483);
   U13556 : OAI21_X2 port map( A1 => n14227, A2 => n4501, B => n3908, ZN => 
                           n6616);
   U13571 : NOR3_X1 port map( A1 => n22842, A2 => n19913, A3 => n735, ZN => 
                           n3928);
   U13575 : XOR2_X1 port map( A1 => n15088, A2 => n3939, Z => n6201);
   U13580 : XOR2_X1 port map( A1 => n27661, A2 => n27573, Z => n16502);
   U13581 : XOR2_X1 port map( A1 => n27573, A2 => n14537, Z => n11844);
   U13582 : XOR2_X1 port map( A1 => n17133, A2 => n27462, Z => n3945);
   U13590 : INV_X4 port map( I => n3953, ZN => n3954);
   U13591 : XOR2_X1 port map( A1 => Plaintext(79), A2 => Key(79), Z => n10813);
   U13593 : NOR2_X1 port map( A1 => n14658, A2 => n24774, ZN => n3964);
   U13594 : INV_X2 port map( I => n14392, ZN => n14658);
   U13596 : XOR2_X1 port map( A1 => n20533, A2 => n3969, Z => n3968);
   U13597 : XOR2_X1 port map( A1 => n20535, A2 => n14619, Z => n3969);
   U13605 : XOR2_X1 port map( A1 => n27393, A2 => n1273, Z => n7857);
   U13607 : XOR2_X1 port map( A1 => n20399, A2 => n3978, Z => n3977);
   U13608 : XOR2_X1 port map( A1 => n28278, A2 => n20508, Z => n3978);
   U13614 : XOR2_X1 port map( A1 => n18362, A2 => n18363, Z => n3985);
   U13616 : OR2_X1 port map( A1 => n19889, A2 => n12393, Z => n3989);
   U13619 : XOR2_X1 port map( A1 => n3996, A2 => n3997, Z => n21695);
   U13622 : XOR2_X1 port map( A1 => n20497, A2 => n20500, Z => n3997);
   U13626 : XOR2_X1 port map( A1 => n5624, A2 => n21894, Z => n10943);
   U13631 : NOR2_X1 port map( A1 => n4404, A2 => n16055, ZN => n4005);
   U13636 : XOR2_X1 port map( A1 => n4019, A2 => n4018, Z => n19614);
   U13643 : XOR2_X1 port map( A1 => n16918, A2 => n20614, Z => n4030);
   U13650 : XOR2_X1 port map( A1 => n4045, A2 => n4044, Z => n4043);
   U13651 : XOR2_X1 port map( A1 => n27415, A2 => n14643, Z => n4044);
   U13656 : XOR2_X1 port map( A1 => n4051, A2 => n4050, Z => n4049);
   U13657 : XOR2_X1 port map( A1 => n27462, A2 => n14491, Z => n4050);
   U13663 : XOR2_X1 port map( A1 => n10641, A2 => n4054, Z => n4053);
   U13664 : XOR2_X1 port map( A1 => n18106, A2 => n21454, Z => n4054);
   U13671 : NAND2_X1 port map( A1 => n961, A2 => n11487, ZN => n19976);
   U13694 : INV_X2 port map( I => n4123, ZN => n15103);
   U13695 : NAND2_X1 port map( A1 => n13628, A2 => n4123, ZN => n4085);
   U13696 : NOR2_X1 port map( A1 => n5042, A2 => n4122, ZN => n4087);
   U13697 : INV_X1 port map( I => n4088, ZN => n5634);
   U13701 : XOR2_X1 port map( A1 => n7200, A2 => n1293, Z => n4093);
   U13707 : XOR2_X1 port map( A1 => n4098, A2 => n4097, Z => n4096);
   U13708 : XOR2_X1 port map( A1 => n6275, A2 => n11275, Z => n4097);
   U13709 : XOR2_X1 port map( A1 => n13904, A2 => n10358, Z => n4098);
   U13711 : XOR2_X1 port map( A1 => n4106, A2 => n15477, Z => n15476);
   U13716 : NAND2_X1 port map( A1 => n4112, A2 => n10980, ZN => n8906);
   U13729 : XOR2_X1 port map( A1 => n16990, A2 => n4129, Z => n4128);
   U13739 : INV_X1 port map( I => n12362, ZN => n4138);
   U13749 : XOR2_X1 port map( A1 => n4147, A2 => n19480, Z => n18897);
   U13755 : XOR2_X1 port map( A1 => n4157, A2 => n4952, Z => n5463);
   U13759 : XOR2_X1 port map( A1 => n6774, A2 => n605, Z => n11821);
   U13764 : NAND2_X1 port map( A1 => n5655, A2 => n4161, ZN => n6469);
   U13766 : NAND2_X1 port map( A1 => n16466, A2 => n9261, ZN => n4165);
   U13769 : XOR2_X1 port map( A1 => n16991, A2 => n7878, Z => n4173);
   U13772 : XOR2_X1 port map( A1 => n14421, A2 => n21650, Z => n4174);
   U13776 : XOR2_X1 port map( A1 => n24528, A2 => n4175, Z => n11460);
   U13778 : XOR2_X1 port map( A1 => n19427, A2 => n19429, Z => n4178);
   U13782 : XOR2_X1 port map( A1 => n4179, A2 => n14503, Z => n9833);
   U13788 : XOR2_X1 port map( A1 => n26717, A2 => n18009, Z => n4183);
   U13789 : XOR2_X1 port map( A1 => n4310, A2 => n13686, Z => n4184);
   U13790 : NOR2_X1 port map( A1 => n25559, A2 => n22643, ZN => n4185);
   U13793 : XOR2_X1 port map( A1 => n4189, A2 => n18333, Z => n4188);
   U13798 : NAND2_X1 port map( A1 => n4191, A2 => n25254, ZN => n11954);
   U13804 : XOR2_X1 port map( A1 => n6554, A2 => n23816, Z => n4193);
   U13806 : XOR2_X1 port map( A1 => n12276, A2 => n18137, Z => n4194);
   U13810 : XOR2_X1 port map( A1 => n25317, A2 => n20952, Z => n4197);
   U13815 : XOR2_X1 port map( A1 => n4203, A2 => n4200, Z => n8529);
   U13816 : XOR2_X1 port map( A1 => n19255, A2 => n4201, Z => n4200);
   U13817 : XOR2_X1 port map( A1 => n19377, A2 => n1292, Z => n4201);
   U13821 : XOR2_X1 port map( A1 => n4204, A2 => n9250, Z => n4838);
   U13822 : XOR2_X1 port map( A1 => n4204, A2 => n18355, Z => n17910);
   U13823 : NOR2_X1 port map( A1 => n23060, A2 => n25339, ZN => n4206);
   U13824 : XOR2_X1 port map( A1 => n4716, A2 => n10974, Z => n4208);
   U13825 : INV_X2 port map( I => n4209, ZN => n7421);
   U13826 : XOR2_X1 port map( A1 => n13680, A2 => n20578, Z => n4211);
   U13838 : XOR2_X1 port map( A1 => n7403, A2 => n21170, Z => n4223);
   U13845 : NAND2_X1 port map( A1 => n5145, A2 => n5952, ZN => n4237);
   U13847 : XOR2_X1 port map( A1 => n16917, A2 => n9505, Z => n4239);
   U13856 : XOR2_X1 port map( A1 => n4260, A2 => n21298, Z => n4259);
   U13861 : INV_X2 port map( I => n4263, ZN => n19913);
   U13863 : AOI21_X1 port map( A1 => n18920, A2 => n26641, B => n9354, ZN => 
                           n14156);
   U13865 : NOR3_X1 port map( A1 => n1164, A2 => n6906, A3 => n26641, ZN => 
                           n13866);
   U13866 : INV_X2 port map( I => n4268, ZN => n18719);
   U13870 : XOR2_X1 port map( A1 => n17073, A2 => n9574, Z => n4273);
   U13874 : NOR3_X1 port map( A1 => n11522, A2 => n4277, A3 => n13021, ZN => 
                           n8541);
   U13879 : XOR2_X1 port map( A1 => n15537, A2 => n20377, Z => n4285);
   U13880 : XOR2_X1 port map( A1 => n12992, A2 => n12316, Z => n4286);
   U13883 : XOR2_X1 port map( A1 => n22756, A2 => n4294, Z => n4293);
   U13884 : NAND2_X2 port map( A1 => n7086, A2 => n9371, ZN => n20377);
   U13885 : XOR2_X1 port map( A1 => n9161, A2 => n21422, Z => n4294);
   U13888 : XOR2_X1 port map( A1 => n16825, A2 => n6765, Z => n4301);
   U13889 : XOR2_X1 port map( A1 => n16875, A2 => n17015, Z => n16825);
   U13895 : NAND2_X1 port map( A1 => n1105, A2 => n4311, ZN => n6498);
   U13898 : NAND2_X1 port map( A1 => n4315, A2 => n6543, ZN => n10366);
   U13904 : AOI21_X2 port map( A1 => n4321, A2 => n17530, B => n4320, ZN => 
                           n8314);
   U13911 : XOR2_X1 port map( A1 => n23041, A2 => n18142, Z => n10365);
   U13912 : XOR2_X1 port map( A1 => n5212, A2 => n4333, Z => n4332);
   U13913 : XOR2_X1 port map( A1 => n4811, A2 => n1280, Z => n4333);
   U13918 : MUX2_X1 port map( I0 => n20074, I1 => n20075, S => n20071, Z => 
                           n4340);
   U13922 : NAND2_X1 port map( A1 => n1013, A2 => n15137, ZN => n12955);
   U13928 : XOR2_X1 port map( A1 => n18174, A2 => n18148, Z => n4360);
   U13929 : XOR2_X1 port map( A1 => n18008, A2 => n12718, Z => n18174);
   U13932 : XOR2_X1 port map( A1 => n19343, A2 => n4373, Z => n4372);
   U13933 : XOR2_X1 port map( A1 => n13752, A2 => n1274, Z => n4373);
   U13934 : XOR2_X1 port map( A1 => n8438, A2 => n19260, Z => n19343);
   U13935 : XOR2_X1 port map( A1 => n4377, A2 => n4376, Z => n4375);
   U13936 : XOR2_X1 port map( A1 => n6878, A2 => n1311, Z => n4376);
   U13937 : XOR2_X1 port map( A1 => n16950, A2 => n23137, Z => n4377);
   U13938 : XOR2_X1 port map( A1 => n15487, A2 => n4382, Z => n4411);
   U13939 : XOR2_X1 port map( A1 => n18112, A2 => n21039, Z => n4382);
   U13940 : XOR2_X1 port map( A1 => n4383, A2 => n20527, Z => n9513);
   U13942 : INV_X2 port map( I => n4384, ZN => n21544);
   U13945 : INV_X2 port map( I => n4386, ZN => n13387);
   U13947 : NAND2_X2 port map( A1 => n4388, A2 => n4387, ZN => n8611);
   U13948 : NOR2_X1 port map( A1 => n14420, A2 => n18428, ZN => n4391);
   U13950 : XOR2_X1 port map( A1 => n5599, A2 => n4399, Z => n7307);
   U13951 : XOR2_X1 port map( A1 => n4398, A2 => n14746, Z => n4399);
   U13956 : NAND2_X1 port map( A1 => n3913, A2 => n26105, ZN => n4404);
   U13957 : NOR2_X1 port map( A1 => n13545, A2 => n1270, ZN => n4405);
   U13964 : XOR2_X1 port map( A1 => n18204, A2 => n604, Z => n4412);
   U13965 : MUX2_X1 port map( I0 => n4413, I1 => n20963, S => n20964, Z => 
                           n20948);
   U13967 : NOR2_X1 port map( A1 => n27468, A2 => n24562, ZN => n4891);
   U13973 : XOR2_X1 port map( A1 => n18244, A2 => n14360, Z => n4422);
   U13976 : XOR2_X1 port map( A1 => n19486, A2 => n4424, Z => n4423);
   U13977 : XOR2_X1 port map( A1 => n24528, A2 => n21341, Z => n4424);
   U13979 : XOR2_X1 port map( A1 => n19231, A2 => n7776, Z => n19042);
   U13984 : XOR2_X1 port map( A1 => n3663, A2 => n20025, Z => n4427);
   U13988 : NAND2_X2 port map( A1 => n4436, A2 => n4433, ZN => n20030);
   U13989 : NAND3_X1 port map( A1 => n18732, A2 => n18733, A3 => n11552, ZN => 
                           n4442);
   U13995 : XNOR2_X1 port map( A1 => n13101, A2 => n14006, ZN => n13131);
   U13996 : AOI22_X2 port map( A1 => n5059, A2 => n14337, B1 => n5061, B2 => 
                           n16472, ZN => n14006);
   U13997 : NAND2_X1 port map( A1 => n4455, A2 => n3292, ZN => n17800);
   U14007 : XOR2_X1 port map( A1 => n26216, A2 => n21679, Z => n6984);
   U14015 : AOI22_X2 port map( A1 => n11211, A2 => n20205, B1 => n11212, B2 => 
                           n5163, ZN => n9397);
   U14016 : XOR2_X1 port map( A1 => n4482, A2 => n4481, Z => n19781);
   U14017 : XOR2_X1 port map( A1 => n19358, A2 => n19410, Z => n4481);
   U14018 : XOR2_X1 port map( A1 => n19388, A2 => n27374, Z => n19410);
   U14019 : XOR2_X1 port map( A1 => n19359, A2 => n4483, Z => n4482);
   U14021 : XOR2_X1 port map( A1 => n25332, A2 => n26566, Z => n4483);
   U14022 : XOR2_X1 port map( A1 => n4484, A2 => Plaintext(122), Z => n15861);
   U14023 : INV_X1 port map( I => Key(122), ZN => n4484);
   U14024 : OAI22_X1 port map( A1 => n15775, A2 => n26371, B1 => n15839, B2 => 
                           n14386, ZN => n8156);
   U14025 : NAND2_X1 port map( A1 => n4486, A2 => n23391, ZN => n13216);
   U14027 : NAND2_X1 port map( A1 => n7961, A2 => n4486, ZN => n17833);
   U14033 : XOR2_X1 port map( A1 => n19268, A2 => n4498, Z => n4497);
   U14035 : XOR2_X1 port map( A1 => n28186, A2 => n14597, Z => n4500);
   U14037 : OAI21_X1 port map( A1 => n7116, A2 => n21499, B => n4516, ZN => 
                           n4515);
   U14039 : XOR2_X1 port map( A1 => n4558, A2 => n4517, Z => n6737);
   U14045 : NAND2_X2 port map( A1 => n4519, A2 => n20196, ZN => n11059);
   U14047 : NAND2_X1 port map( A1 => n20194, A2 => n20195, ZN => n4521);
   U14051 : XOR2_X1 port map( A1 => n24659, A2 => n12633, Z => n13978);
   U14055 : XOR2_X1 port map( A1 => n19236, A2 => n4530, Z => n19465);
   U14064 : XOR2_X1 port map( A1 => n10387, A2 => n4534, Z => n4533);
   U14065 : XOR2_X1 port map( A1 => n12523, A2 => n14543, Z => n4534);
   U14071 : AOI21_X1 port map( A1 => n13822, A2 => n11385, B => n4539, ZN => 
                           n4538);
   U14073 : OAI22_X1 port map( A1 => n4541, A2 => n13822, B1 => n21169, B2 => 
                           n27368, ZN => n4540);
   U14075 : XOR2_X1 port map( A1 => n11644, A2 => n14693, Z => n6545);
   U14079 : NOR2_X1 port map( A1 => n4549, A2 => n7468, ZN => n8555);
   U14080 : NAND2_X1 port map( A1 => n7770, A2 => n24286, ZN => n8214);
   U14081 : NAND2_X2 port map( A1 => n16286, A2 => n14893, ZN => n7897);
   U14083 : XOR2_X1 port map( A1 => n26486, A2 => n21732, Z => n4560);
   U14085 : AOI21_X2 port map( A1 => n4566, A2 => n4565, B => n4564, ZN => 
                           n15703);
   U14087 : XOR2_X1 port map( A1 => n17130, A2 => n17128, Z => n4568);
   U14092 : OR2_X1 port map( A1 => n18633, A2 => n457, Z => n4574);
   U14095 : XOR2_X1 port map( A1 => n18144, A2 => n11364, Z => n4580);
   U14096 : AOI21_X1 port map( A1 => n21021, A2 => n22737, B => n4581, ZN => 
                           n9426);
   U14101 : XOR2_X1 port map( A1 => n4585, A2 => n4587, Z => n10458);
   U14102 : XOR2_X1 port map( A1 => n27438, A2 => n25980, Z => n4587);
   U14104 : XOR2_X1 port map( A1 => n4601, A2 => n11933, Z => n16942);
   U14106 : AND2_X1 port map( A1 => n11932, A2 => n15029, Z => n11095);
   U14107 : INV_X1 port map( I => n20963, ZN => n20951);
   U14110 : OAI21_X1 port map( A1 => n20950, A2 => n4607, B => n23088, ZN => 
                           n4606);
   U14116 : XOR2_X1 port map( A1 => n4619, A2 => n4621, Z => n9022);
   U14117 : XOR2_X1 port map( A1 => n17080, A2 => n4620, Z => n4619);
   U14118 : XOR2_X1 port map( A1 => n17055, A2 => n1278, Z => n4620);
   U14120 : XOR2_X1 port map( A1 => n9399, A2 => n4622, Z => n4621);
   U14121 : XOR2_X1 port map( A1 => n16975, A2 => n26141, Z => n4622);
   U14122 : AOI21_X2 port map( A1 => n12615, A2 => n4623, B => n15570, ZN => 
                           n15499);
   U14129 : XOR2_X1 port map( A1 => n19323, A2 => n4628, Z => n4627);
   U14130 : XOR2_X1 port map( A1 => n27397, A2 => n20912, Z => n4628);
   U14135 : XOR2_X1 port map( A1 => n20459, A2 => n8885, Z => n20522);
   U14136 : OAI21_X2 port map( A1 => n28121, A2 => n19799, B => n4632, ZN => 
                           n20294);
   U14139 : XOR2_X1 port map( A1 => n21376, A2 => n20949, Z => n4635);
   U14140 : XOR2_X1 port map( A1 => n26029, A2 => n24887, Z => n4636);
   U14142 : XOR2_X1 port map( A1 => n20551, A2 => n4638, Z => n4637);
   U14143 : XOR2_X1 port map( A1 => n21185, A2 => n20552, Z => n4638);
   U14145 : XOR2_X1 port map( A1 => n20424, A2 => n20447, Z => n20551);
   U14148 : OAI21_X2 port map( A1 => n20276, A2 => n4660, B => n4648, ZN => 
                           n21258);
   U14149 : AOI22_X1 port map( A1 => n751, A2 => n4650, B1 => n10931, B2 => 
                           n4649, ZN => n4648);
   U14150 : XOR2_X1 port map( A1 => n8636, A2 => n24384, Z => n19341);
   U14151 : NOR2_X2 port map( A1 => n19662, A2 => n19663, ZN => n20273);
   U14162 : XOR2_X1 port map( A1 => n7476, A2 => n7474, Z => n13181);
   U14168 : XOR2_X1 port map( A1 => n17026, A2 => n919, Z => n4673);
   U14173 : XOR2_X1 port map( A1 => n18229, A2 => n4681, Z => n4680);
   U14181 : XOR2_X1 port map( A1 => n20547, A2 => n4685, Z => n4684);
   U14182 : XOR2_X1 port map( A1 => n136, A2 => n20617, Z => n4685);
   U14186 : XOR2_X1 port map( A1 => n5097, A2 => n20548, Z => n4686);
   U14187 : XOR2_X1 port map( A1 => n21374, A2 => n20449, Z => n20548);
   U14198 : XOR2_X1 port map( A1 => n3830, A2 => n4698, Z => n4697);
   U14199 : XOR2_X1 port map( A1 => n4707, A2 => n16966, Z => n16967);
   U14200 : XOR2_X1 port map( A1 => n4708, A2 => n19367, Z => n12351);
   U14201 : XOR2_X1 port map( A1 => n4708, A2 => n13938, Z => n13937);
   U14203 : NAND2_X2 port map( A1 => n4711, A2 => n15748, ZN => n14641);
   U14209 : XOR2_X1 port map( A1 => n4722, A2 => n4724, Z => n5689);
   U14210 : XOR2_X1 port map( A1 => n21893, A2 => n4723, Z => n4722);
   U14215 : XOR2_X1 port map( A1 => n26719, A2 => n9498, Z => n4724);
   U14219 : AND2_X1 port map( A1 => n2844, A2 => n1071, Z => n4728);
   U14222 : INV_X2 port map( I => n15414, ZN => n10764);
   U14226 : XOR2_X1 port map( A1 => n4744, A2 => n4743, Z => n10497);
   U14231 : XOR2_X1 port map( A1 => n27936, A2 => n1289, Z => n4747);
   U14232 : XOR2_X1 port map( A1 => Plaintext(128), A2 => Key(128), Z => n4762)
                           ;
   U14234 : NAND2_X1 port map( A1 => n24513, A2 => n17509, ZN => n4755);
   U14235 : XOR2_X1 port map( A1 => n4966, A2 => n27438, Z => n20524);
   U14236 : MUX2_X1 port map( I0 => n18841, I1 => n7468, S => n26570, Z => 
                           n4759);
   U14237 : NAND2_X1 port map( A1 => n4760, A2 => n13709, ZN => n11388);
   U14244 : NOR2_X1 port map( A1 => n20662, A2 => n4767, ZN => n4937);
   U14246 : NAND2_X2 port map( A1 => n12047, A2 => n18453, ZN => n7468);
   U14247 : NAND3_X1 port map( A1 => n27905, A2 => n972, A3 => n19748, ZN => 
                           n4771);
   U14248 : XOR2_X1 port map( A1 => n4776, A2 => n20769, Z => n16864);
   U14249 : XOR2_X1 port map( A1 => n4776, A2 => n4808, Z => n4807);
   U14250 : INV_X1 port map( I => Plaintext(136), ZN => n9023);
   U14257 : NAND2_X1 port map( A1 => n4783, A2 => n20030, ZN => n15412);
   U14258 : NOR2_X1 port map( A1 => n4790, A2 => n4783, ZN => n11747);
   U14260 : XOR2_X1 port map( A1 => n27369, A2 => n4789, Z => n11004);
   U14261 : XOR2_X1 port map( A1 => n4789, A2 => n7408, Z => n19196);
   U14262 : XOR2_X1 port map( A1 => n1140, A2 => n4789, Z => n19339);
   U14267 : XOR2_X1 port map( A1 => n2462, A2 => n7403, Z => n12228);
   U14268 : XOR2_X1 port map( A1 => n9736, A2 => n22836, Z => n4794);
   U14269 : XOR2_X1 port map( A1 => n18116, A2 => n5079, Z => n4795);
   U14271 : XOR2_X1 port map( A1 => n8673, A2 => n16808, Z => n4809);
   U14273 : XOR2_X1 port map( A1 => n4811, A2 => n21085, Z => n8959);
   U14274 : XOR2_X1 port map( A1 => n10123, A2 => n4811, Z => n16735);
   U14277 : NAND2_X1 port map( A1 => n20618, A2 => n4822, ZN => n20611);
   U14278 : NOR2_X1 port map( A1 => n20618, A2 => n4822, ZN => n20616);
   U14284 : XOR2_X1 port map( A1 => n27370, A2 => n20377, Z => n6941);
   U14285 : OAI21_X1 port map( A1 => n9575, A2 => n21524, B => n4827, ZN => 
                           n9578);
   U14293 : XOR2_X1 port map( A1 => n21199, A2 => n28186, Z => n4836);
   U14295 : XOR2_X1 port map( A1 => n10887, A2 => n4838, Z => n4837);
   U14298 : XOR2_X1 port map( A1 => n4848, A2 => n20877, Z => Ciphertext(52));
   U14300 : NAND2_X1 port map( A1 => n4859, A2 => n12265, ZN => n12263);
   U14302 : NAND2_X1 port map( A1 => n4860, A2 => n20703, ZN => n8389);
   U14307 : INV_X2 port map( I => n4873, ZN => n9887);
   U14310 : XOR2_X1 port map( A1 => n15647, A2 => n4878, Z => n7559);
   U14315 : OAI22_X2 port map( A1 => n10981, A2 => n16366, B1 => n16368, B2 => 
                           n16367, ZN => n16863);
   U14316 : INV_X1 port map( I => n27468, ZN => n12729);
   U14317 : AND2_X1 port map( A1 => n11869, A2 => n3971, Z => n4892);
   U14322 : XOR2_X1 port map( A1 => n20776, A2 => n20775, Z => n4897);
   U14325 : XOR2_X1 port map( A1 => n4901, A2 => n5940, Z => n4952);
   U14329 : NOR2_X1 port map( A1 => n7733, A2 => n23817, ZN => n7732);
   U14330 : XOR2_X1 port map( A1 => n4904, A2 => n4905, Z => n4903);
   U14331 : XOR2_X1 port map( A1 => n16875, A2 => n1318, Z => n4904);
   U14332 : XOR2_X1 port map( A1 => n25582, A2 => n16958, Z => n4905);
   U14336 : NAND3_X2 port map( A1 => n15972, A2 => n9110, A3 => n9111, ZN => 
                           n8378);
   U14343 : XOR2_X1 port map( A1 => n19542, A2 => n4919, Z => n4918);
   U14347 : XOR2_X1 port map( A1 => n4922, A2 => n4921, Z => n17183);
   U14348 : XOR2_X1 port map( A1 => n15214, A2 => n15215, Z => n4921);
   U14353 : NAND2_X1 port map( A1 => n9280, A2 => n850, ZN => n7537);
   U14354 : XOR2_X1 port map( A1 => Plaintext(44), A2 => Key(44), Z => n9437);
   U14355 : OAI21_X1 port map( A1 => n10768, A2 => n16811, B => n4940, ZN => 
                           n16815);
   U14357 : XOR2_X1 port map( A1 => n13761, A2 => n9055, Z => n4943);
   U14362 : XOR2_X1 port map( A1 => n7200, A2 => n20602, Z => n4949);
   U14363 : INV_X2 port map( I => n4950, ZN => n11354);
   U14366 : NOR2_X1 port map( A1 => n26645, A2 => n4953, ZN => n13663);
   U14368 : XOR2_X1 port map( A1 => n7257, A2 => n13200, Z => n4956);
   U14372 : XOR2_X1 port map( A1 => n12816, A2 => n1311, Z => n4964);
   U14374 : NOR2_X1 port map( A1 => n21970, A2 => n23744, ZN => n12693);
   U14376 : XOR2_X1 port map( A1 => n24255, A2 => n7027, Z => n14085);
   U14379 : NAND2_X2 port map( A1 => n4661, A2 => n1177, ZN => n6827);
   U14382 : XOR2_X1 port map( A1 => n4988, A2 => n4985, Z => n6624);
   U14384 : XOR2_X1 port map( A1 => n2265, A2 => n21683, Z => n4986);
   U14385 : XOR2_X1 port map( A1 => n15256, A2 => n8880, Z => n4987);
   U14386 : OAI21_X1 port map( A1 => n21969, A2 => n13613, B => n16339, ZN => 
                           n13588);
   U14390 : XOR2_X1 port map( A1 => n23369, A2 => n23750, Z => n4992);
   U14391 : NOR2_X2 port map( A1 => n10397, A2 => n16675, ZN => n5379);
   U14392 : XOR2_X1 port map( A1 => n16989, A2 => n14572, Z => n4994);
   U14394 : XOR2_X1 port map( A1 => n28263, A2 => n22381, Z => n4995);
   U14395 : XOR2_X1 port map( A1 => n13064, A2 => n18128, Z => n4996);
   U14398 : XOR2_X1 port map( A1 => n5001, A2 => n21419, Z => Ciphertext(128));
   U14401 : XOR2_X1 port map( A1 => Plaintext(125), A2 => Key(125), Z => n8264)
                           ;
   U14405 : XOR2_X1 port map( A1 => n5013, A2 => n5010, Z => n12653);
   U14406 : XOR2_X1 port map( A1 => n5011, A2 => n5012, Z => n5010);
   U14407 : XOR2_X1 port map( A1 => n27604, A2 => n14643, Z => n5011);
   U14408 : XOR2_X1 port map( A1 => n21373, A2 => n10339, Z => n5012);
   U14409 : XOR2_X1 port map( A1 => n19352, A2 => n19451, Z => n19407);
   U14410 : NAND2_X1 port map( A1 => n16375, A2 => n3470, ZN => n15631);
   U14414 : XOR2_X1 port map( A1 => n13410, A2 => n5025, Z => n5024);
   U14415 : XOR2_X1 port map( A1 => n4558, A2 => n22512, Z => n5025);
   U14428 : XOR2_X1 port map( A1 => n5619, A2 => n5043, Z => n21728);
   U14429 : NAND2_X1 port map( A1 => n24576, A2 => n4122, ZN => n5044);
   U14433 : NAND2_X1 port map( A1 => n12482, A2 => n14137, ZN => n5060);
   U14436 : XOR2_X1 port map( A1 => n5064, A2 => n1142, Z => n5063);
   U14437 : XOR2_X1 port map( A1 => n11417, A2 => n5740, Z => n5064);
   U14443 : NAND4_X1 port map( A1 => n28545, A2 => n14721, A3 => n13494, A4 => 
                           n5070, ZN => n13015);
   U14444 : NAND2_X2 port map( A1 => n5075, A2 => n5072, ZN => n16455);
   U14446 : NOR2_X1 port map( A1 => n26371, A2 => n7235, ZN => n5074);
   U14448 : OAI21_X1 port map( A1 => n9217, A2 => n6022, B => n13687, ZN => 
                           n17197);
   U14449 : XOR2_X1 port map( A1 => n6675, A2 => n14637, Z => n5079);
   U14451 : XOR2_X1 port map( A1 => n1198, A2 => n18237, Z => n9736);
   U14455 : NOR2_X1 port map( A1 => n27010, A2 => n27129, ZN => n20080);
   U14457 : NAND3_X1 port map( A1 => n25130, A2 => n24028, A3 => n11413, ZN => 
                           n5776);
   U14459 : XOR2_X1 port map( A1 => n5086, A2 => n5083, Z => n7706);
   U14460 : XOR2_X1 port map( A1 => n5084, A2 => n5085, Z => n5083);
   U14461 : XOR2_X1 port map( A1 => n23156, A2 => n920, Z => n5084);
   U14462 : XOR2_X1 port map( A1 => n36, A2 => n20448, Z => n5085);
   U14466 : AOI22_X2 port map( A1 => n10717, A2 => n11073, B1 => n20193, B2 => 
                           n20192, ZN => n21376);
   U14472 : INV_X2 port map( I => n9022, ZN => n5541);
   U14473 : XOR2_X1 port map( A1 => n1638, A2 => n27589, Z => n9582);
   U14474 : XOR2_X1 port map( A1 => n20565, A2 => n1638, Z => n20412);
   U14475 : XOR2_X1 port map( A1 => n12468, A2 => n1638, Z => n19725);
   U14476 : XNOR2_X1 port map( A1 => Plaintext(52), A2 => Key(52), ZN => n5095)
                           ;
   U14477 : INV_X1 port map( I => n7175, ZN => n5096);
   U14478 : XOR2_X1 port map( A1 => n13761, A2 => n21373, Z => n5097);
   U14479 : XOR2_X1 port map( A1 => n9981, A2 => n5097, Z => n8671);
   U14480 : INV_X2 port map( I => n12695, ZN => n19819);
   U14484 : XOR2_X1 port map( A1 => n19350, A2 => n20919, Z => n5105);
   U14488 : NAND2_X2 port map( A1 => n16385, A2 => n16384, ZN => n16897);
   U14490 : INV_X1 port map( I => n5122, ZN => n16633);
   U14493 : NAND2_X1 port map( A1 => n14137, A2 => n16619, ZN => n5124);
   U14498 : NOR2_X1 port map( A1 => n16557, A2 => n26396, ZN => n11195);
   U14500 : INV_X2 port map( I => n5140, ZN => n14695);
   U14503 : XOR2_X1 port map( A1 => n5142, A2 => n5144, Z => n15225);
   U14504 : XOR2_X1 port map( A1 => n12604, A2 => n5143, Z => n5142);
   U14509 : NAND2_X2 port map( A1 => n5228, A2 => n18765, ZN => n11552);
   U14514 : NOR2_X1 port map( A1 => n9734, A2 => n11497, ZN => n5153);
   U14519 : XOR2_X1 port map( A1 => n19188, A2 => n9335, Z => n5168);
   U14520 : XOR2_X1 port map( A1 => n14876, A2 => n1320, Z => n5547);
   U14524 : XOR2_X1 port map( A1 => n18237, A2 => n18168, Z => n18273);
   U14525 : NAND2_X2 port map( A1 => n17836, A2 => n17835, ZN => n18168);
   U14528 : OR2_X1 port map( A1 => n13756, A2 => n11467, Z => n10371);
   U14532 : AND2_X1 port map( A1 => n563, A2 => n16274, Z => n8812);
   U14537 : XOR2_X1 port map( A1 => n5186, A2 => n14479, Z => Ciphertext(143));
   U14546 : INV_X1 port map( I => n18863, ZN => n5189);
   U14550 : NAND2_X2 port map( A1 => n19104, A2 => n19103, ZN => n19210);
   U14553 : XOR2_X1 port map( A1 => n8788, A2 => n5194, Z => n8786);
   U14555 : OR2_X1 port map( A1 => n6433, A2 => n7319, Z => n13517);
   U14563 : NAND2_X2 port map( A1 => n16478, A2 => n14122, ZN => n17088);
   U14564 : AOI22_X2 port map( A1 => n12450, A2 => n17182, B1 => n8367, B2 => 
                           n17184, ZN => n17726);
   U14567 : AOI21_X1 port map( A1 => n12096, A2 => n24190, B => n27252, ZN => 
                           n13059);
   U14573 : NAND2_X1 port map( A1 => n15959, A2 => n8922, ZN => n7662);
   U14575 : NAND2_X1 port map( A1 => n24286, A2 => n18602, ZN => n8354);
   U14578 : XOR2_X1 port map( A1 => n5210, A2 => n19477, Z => n19314);
   U14579 : XOR2_X1 port map( A1 => n19536, A2 => n23480, Z => n5210);
   U14582 : XOR2_X1 port map( A1 => n11672, A2 => n11630, Z => n7589);
   U14583 : NAND2_X1 port map( A1 => n23225, A2 => n5216, ZN => n5215);
   U14584 : NAND2_X1 port map( A1 => n7299, A2 => n15378, ZN => n5216);
   U14587 : XOR2_X1 port map( A1 => n20060, A2 => n20445, Z => n20061);
   U14593 : XOR2_X1 port map( A1 => n16818, A2 => n8178, Z => n8177);
   U14600 : INV_X2 port map( I => n5226, ZN => n18557);
   U14604 : XOR2_X1 port map( A1 => n21890, A2 => n10676, Z => n6638);
   U14607 : OR2_X1 port map( A1 => n10126, A2 => n1699, Z => n12373);
   U14609 : NAND3_X1 port map( A1 => n14038, A2 => n25327, A3 => n12139, ZN => 
                           n5228);
   U14615 : INV_X2 port map( I => n11491, ZN => n5253);
   U14619 : XOR2_X1 port map( A1 => n12533, A2 => n10352, Z => n6060);
   U14620 : NAND2_X1 port map( A1 => n16528, A2 => n15203, ZN => n5240);
   U14622 : NAND2_X2 port map( A1 => n19670, A2 => n5234, ZN => n20277);
   U14624 : OR2_X1 port map( A1 => n20875, A2 => n11869, Z => n7827);
   U14627 : INV_X1 port map( I => n14533, ZN => n5978);
   U14634 : AND2_X1 port map( A1 => n17578, A2 => n2895, Z => n6389);
   U14635 : NAND3_X1 port map( A1 => n10797, A2 => n27403, A3 => n952, ZN => 
                           n10174);
   U14636 : AND2_X1 port map( A1 => n16278, A2 => n12507, Z => n10740);
   U14643 : XOR2_X1 port map( A1 => n18167, A2 => n12361, Z => n9025);
   U14648 : NAND2_X2 port map( A1 => n7629, A2 => n7628, ZN => n16619);
   U14653 : AOI21_X2 port map( A1 => n8940, A2 => n7357, B => n5254, ZN => 
                           n8939);
   U14657 : XNOR2_X1 port map( A1 => n13916, A2 => n20396, ZN => n10855);
   U14668 : XOR2_X1 port map( A1 => n5268, A2 => n6866, Z => n19891);
   U14669 : XOR2_X1 port map( A1 => n6808, A2 => n9071, Z => n5268);
   U14675 : NAND2_X1 port map( A1 => n20146, A2 => n20197, ZN => n5271);
   U14679 : OR2_X1 port map( A1 => n17460, A2 => n5605, Z => n17462);
   U14682 : XOR2_X1 port map( A1 => n5272, A2 => n7713, Z => n8948);
   U14683 : XOR2_X1 port map( A1 => n20531, A2 => n20530, Z => n5272);
   U14689 : INV_X2 port map( I => n5277, ZN => n7370);
   U14693 : XOR2_X1 port map( A1 => n22760, A2 => n25098, Z => n19294);
   U14695 : XOR2_X1 port map( A1 => n12099, A2 => n27378, Z => n20554);
   U14704 : XOR2_X1 port map( A1 => n28460, A2 => n658, Z => n7425);
   U14705 : XOR2_X1 port map( A1 => n5287, A2 => n22820, Z => n9214);
   U14707 : OAI21_X2 port map( A1 => n13781, A2 => n15833, B => n15919, ZN => 
                           n16250);
   U14709 : XOR2_X1 port map( A1 => n18251, A2 => n18250, Z => n5289);
   U14727 : OR2_X1 port map( A1 => n17506, A2 => n9021, Z => n5300);
   U14728 : XOR2_X1 port map( A1 => n617, A2 => n17115, Z => n11762);
   U14730 : NAND2_X1 port map( A1 => n13988, A2 => n21998, ZN => n7381);
   U14731 : NAND2_X2 port map( A1 => n12837, A2 => n15838, ZN => n12839);
   U14733 : XOR2_X1 port map( A1 => n5303, A2 => n14544, Z => Ciphertext(39));
   U14737 : XOR2_X1 port map( A1 => n5304, A2 => n20807, Z => Ciphertext(41));
   U14739 : XOR2_X1 port map( A1 => n5492, A2 => n13750, Z => n14852);
   U14741 : NAND2_X2 port map( A1 => n28545, A2 => n14721, ZN => n19167);
   U14745 : NOR2_X1 port map( A1 => n13764, A2 => n11839, ZN => n13763);
   U14749 : XOR2_X1 port map( A1 => n18035, A2 => n27451, Z => n7792);
   U14750 : XOR2_X1 port map( A1 => n18355, A2 => n18113, Z => n18035);
   U14754 : XOR2_X1 port map( A1 => n16889, A2 => n16834, Z => n6276);
   U14756 : XOR2_X1 port map( A1 => n19406, A2 => n28263, Z => n8675);
   U14757 : OR2_X1 port map( A1 => n19160, A2 => n22237, Z => n9032);
   U14764 : NOR2_X1 port map( A1 => n10580, A2 => n25374, ZN => n10725);
   U14768 : XOR2_X1 port map( A1 => n11644, A2 => n9876, Z => n5613);
   U14771 : XOR2_X1 port map( A1 => n6706, A2 => n626, Z => n6703);
   U14774 : NAND3_X1 port map( A1 => n15701, A2 => n16475, A3 => n16151, ZN => 
                           n16152);
   U14775 : XOR2_X1 port map( A1 => n5597, A2 => n14650, Z => n10786);
   U14776 : OR2_X1 port map( A1 => n13885, A2 => n13886, Z => n5325);
   U14779 : XOR2_X1 port map( A1 => n5819, A2 => n5820, Z => n16935);
   U14781 : XOR2_X1 port map( A1 => n19529, A2 => n14325, Z => n5328);
   U14784 : OR2_X1 port map( A1 => n15986, A2 => n16145, Z => n15825);
   U14785 : XOR2_X1 port map( A1 => Plaintext(67), A2 => Key(67), Z => n15526);
   U14787 : XOR2_X1 port map( A1 => Plaintext(23), A2 => Key(23), Z => n5333);
   U14789 : XOR2_X1 port map( A1 => n12803, A2 => n12783, Z => n10063);
   U14791 : XOR2_X1 port map( A1 => n20440, A2 => n5335, Z => n5334);
   U14803 : INV_X1 port map( I => n20363, ZN => n7975);
   U14804 : NAND2_X1 port map( A1 => n12795, A2 => n24574, ZN => n5344);
   U14810 : OR2_X1 port map( A1 => n17715, A2 => n17623, Z => n5349);
   U14815 : XOR2_X1 port map( A1 => n18186, A2 => n12902, Z => n18187);
   U14817 : NAND2_X1 port map( A1 => n19816, A2 => n960, ZN => n12632);
   U14819 : XOR2_X1 port map( A1 => n21302, A2 => n20552, Z => n20531);
   U14823 : NAND2_X1 port map( A1 => n21267, A2 => n21498, ZN => n5355);
   U14825 : NAND2_X1 port map( A1 => n19876, A2 => n19842, ZN => n5357);
   U14830 : OR2_X1 port map( A1 => n19806, A2 => n13863, Z => n19543);
   U14832 : OR2_X1 port map( A1 => n20663, A2 => n20658, Z => n15580);
   U14835 : AND2_X1 port map( A1 => n7977, A2 => n8215, Z => n6804);
   U14840 : NAND2_X1 port map( A1 => n7955, A2 => n7954, ZN => n20854);
   U14843 : OAI21_X1 port map( A1 => n22536, A2 => n6323, B => n27375, ZN => 
                           n7913);
   U14845 : XOR2_X1 port map( A1 => n22771, A2 => n14623, Z => n10974);
   U14847 : XOR2_X1 port map( A1 => n5369, A2 => n14572, Z => Ciphertext(83));
   U14848 : OAI22_X1 port map( A1 => n21051, A2 => n21050, B1 => n21053, B2 => 
                           n9421, ZN => n5369);
   U14855 : XOR2_X1 port map( A1 => n9123, A2 => n14404, Z => n9803);
   U14862 : NAND2_X2 port map( A1 => n19963, A2 => n19964, ZN => n20280);
   U14864 : NAND2_X1 port map( A1 => n7565, A2 => n19147, ZN => n10315);
   U14877 : NAND2_X1 port map( A1 => n943, A2 => n9377, ZN => n15702);
   U14878 : INV_X2 port map( I => n5401, ZN => n5797);
   U14881 : AND2_X1 port map( A1 => n5680, A2 => n16207, Z => n5569);
   U14886 : XOR2_X1 port map( A1 => n18336, A2 => n5912, Z => n5911);
   U14887 : XOR2_X1 port map( A1 => n5412, A2 => n14535, Z => Ciphertext(179));
   U14890 : XOR2_X1 port map( A1 => n9524, A2 => n13225, Z => n5417);
   U14899 : XOR2_X1 port map( A1 => n6759, A2 => n6760, Z => n6860);
   U14903 : NAND2_X1 port map( A1 => n5656, A2 => n28543, ZN => n5655);
   U14911 : NAND2_X1 port map( A1 => n21566, A2 => n27118, ZN => n13128);
   U14918 : XOR2_X1 port map( A1 => n11511, A2 => n11513, Z => n19584);
   U14933 : OR2_X1 port map( A1 => n10393, A2 => n6843, Z => n10392);
   U14934 : NOR2_X1 port map( A1 => n13327, A2 => n23488, ZN => n5491);
   U14941 : INV_X2 port map( I => n5448, ZN => n15981);
   U14942 : XNOR2_X1 port map( A1 => Plaintext(57), A2 => Key(57), ZN => n5448)
                           ;
   U14943 : INV_X2 port map( I => n5450, ZN => n21586);
   U14946 : XOR2_X1 port map( A1 => n5454, A2 => n24840, Z => Ciphertext(158));
   U14950 : XOR2_X1 port map( A1 => n16744, A2 => n21613, Z => n10684);
   U14951 : NAND2_X2 port map( A1 => n5456, A2 => n8815, ZN => n8740);
   U14952 : NAND2_X2 port map( A1 => n6483, A2 => n6484, ZN => n8882);
   U14954 : XOR2_X1 port map( A1 => n16820, A2 => n16836, Z => n17102);
   U14956 : NOR2_X1 port map( A1 => n27671, A2 => n6504, ZN => n6503);
   U14961 : INV_X2 port map( I => n5463, ZN => n13564);
   U14964 : XOR2_X1 port map( A1 => n5755, A2 => n5468, Z => n5752);
   U14965 : XOR2_X1 port map( A1 => n12182, A2 => n15022, Z => n5468);
   U14973 : AOI21_X1 port map( A1 => n15165, A2 => n15333, B => n15164, ZN => 
                           n15163);
   U14978 : XOR2_X1 port map( A1 => n7221, A2 => n16910, Z => n5474);
   U14979 : NAND2_X2 port map( A1 => n6967, A2 => n18177, ZN => n19019);
   U14980 : XOR2_X1 port map( A1 => n5479, A2 => n6871, Z => n21270);
   U14981 : XOR2_X1 port map( A1 => n10084, A2 => n20532, Z => n5479);
   U14984 : XOR2_X1 port map( A1 => n13314, A2 => n18352, Z => n5481);
   U14990 : INV_X1 port map( I => n19693, ZN => n9401);
   U14994 : NAND2_X1 port map( A1 => n21605, A2 => n21608, ZN => n5486);
   U14996 : XOR2_X1 port map( A1 => n5490, A2 => n1096, Z => n6597);
   U14998 : INV_X1 port map( I => n14089, ZN => n8699);
   U14999 : XOR2_X1 port map( A1 => n18900, A2 => n24532, Z => n5494);
   U15000 : NOR2_X1 port map( A1 => n7817, A2 => n6968, ZN => n18599);
   U15010 : XOR2_X1 port map( A1 => n18106, A2 => n11502, Z => n18210);
   U15013 : NOR2_X1 port map( A1 => n10428, A2 => n15560, ZN => n11206);
   U15015 : NAND2_X2 port map( A1 => n18816, A2 => n18815, ZN => n13812);
   U15019 : OR2_X1 port map( A1 => n8430, A2 => n5535, Z => n8348);
   U15020 : INV_X2 port map( I => n5505, ZN => n10289);
   U15027 : XOR2_X1 port map( A1 => n21255, A2 => n20880, Z => n10277);
   U15028 : NAND2_X2 port map( A1 => n9955, A2 => n9957, ZN => n21255);
   U15047 : NAND2_X2 port map( A1 => n21445, A2 => n5519, ZN => n21446);
   U15049 : INV_X2 port map( I => n5521, ZN => n7682);
   U15050 : INV_X1 port map( I => n6799, ZN => n6877);
   U15051 : XOR2_X1 port map( A1 => n5522, A2 => n6296, Z => n6625);
   U15053 : XOR2_X1 port map( A1 => n6106, A2 => n6105, Z => n7067);
   U15057 : XOR2_X1 port map( A1 => n6059, A2 => n6060, Z => n5524);
   U15059 : XOR2_X1 port map( A1 => n5379, A2 => n23053, Z => n16852);
   U15064 : XOR2_X1 port map( A1 => n5530, A2 => n5531, Z => n13727);
   U15066 : OAI21_X1 port map( A1 => n20868, A2 => n20866, B => n5532, ZN => 
                           n20760);
   U15075 : NAND2_X1 port map( A1 => n6466, A2 => n13934, ZN => n6465);
   U15080 : XOR2_X1 port map( A1 => n19171, A2 => n19184, Z => n6220);
   U15081 : XOR2_X1 port map( A1 => n5867, A2 => n6739, Z => n20735);
   U15084 : XOR2_X1 port map( A1 => n5543, A2 => n655, Z => n10704);
   U15087 : OR2_X1 port map( A1 => n18780, A2 => n10579, Z => n5545);
   U15089 : XNOR2_X1 port map( A1 => n21336, A2 => n11097, ZN => n7267);
   U15096 : INV_X2 port map( I => n5550, ZN => n13188);
   U15099 : NAND2_X1 port map( A1 => n11873, A2 => n5554, ZN => n10203);
   U15102 : INV_X2 port map( I => n16691, ZN => n5558);
   U15109 : XNOR2_X1 port map( A1 => Plaintext(56), A2 => Key(56), ZN => n5580)
                           ;
   U15116 : NAND2_X1 port map( A1 => n17711, A2 => n5584, ZN => n10983);
   U15120 : XOR2_X1 port map( A1 => n5589, A2 => n19409, Z => n5588);
   U15121 : XOR2_X1 port map( A1 => n7346, A2 => n19560, Z => n5589);
   U15123 : XOR2_X1 port map( A1 => n5593, A2 => n5591, Z => n5590);
   U15124 : XOR2_X1 port map( A1 => n12959, A2 => n5592, Z => n5591);
   U15130 : XOR2_X1 port map( A1 => n18112, A2 => n5601, Z => n5600);
   U15133 : INV_X2 port map( I => n5605, ZN => n9898);
   U15139 : INV_X2 port map( I => n15632, ZN => n5612);
   U15144 : NAND2_X1 port map( A1 => n16267, A2 => n16268, ZN => n5617);
   U15145 : XOR2_X1 port map( A1 => n14700, A2 => n14699, Z => n20555);
   U15146 : XOR2_X1 port map( A1 => n14372, A2 => n9964, Z => n5619);
   U15148 : XOR2_X1 port map( A1 => n27437, A2 => n20741, Z => n20716);
   U15149 : XOR2_X1 port map( A1 => n5623, A2 => n21426, Z => n21427);
   U15150 : XOR2_X1 port map( A1 => n5623, A2 => n7011, Z => n8807);
   U15152 : NOR2_X1 port map( A1 => n21395, A2 => n14759, ZN => n5627);
   U15160 : XOR2_X1 port map( A1 => n20547, A2 => n5647, Z => n5646);
   U15161 : XOR2_X1 port map( A1 => n20581, A2 => n20692, Z => n5647);
   U15168 : NOR2_X1 port map( A1 => n21050, A2 => n9421, ZN => n5663);
   U15172 : AND2_X1 port map( A1 => n23474, A2 => n24089, Z => n5666);
   U15175 : INV_X2 port map( I => n14677, ZN => n5675);
   U15176 : XOR2_X1 port map( A1 => Plaintext(21), A2 => Key(21), Z => n14433);
   U15178 : XOR2_X1 port map( A1 => n5682, A2 => n14624, Z => n21306);
   U15179 : XOR2_X1 port map( A1 => n5446, A2 => n5682, Z => n20440);
   U15184 : XOR2_X1 port map( A1 => n21301, A2 => n5687, Z => n5686);
   U15185 : XOR2_X1 port map( A1 => n23849, A2 => n1279, Z => n5687);
   U15186 : INV_X2 port map( I => n5689, ZN => n11426);
   U15187 : NAND2_X1 port map( A1 => n822, A2 => n23713, ZN => n5691);
   U15190 : NOR2_X1 port map( A1 => n7854, A2 => n5707, ZN => n5706);
   U15192 : XOR2_X1 port map( A1 => n5712, A2 => n21683, Z => Ciphertext(178));
   U15200 : XOR2_X1 port map( A1 => n20725, A2 => n14273, Z => n5727);
   U15202 : INV_X2 port map( I => n10447, ZN => n5740);
   U15203 : XOR2_X1 port map( A1 => n25166, A2 => n21039, Z => n5741);
   U15206 : XOR2_X1 port map( A1 => n5742, A2 => n21037, Z => n17823);
   U15208 : NAND2_X2 port map( A1 => n7074, A2 => n8708, ZN => n5742);
   U15209 : XOR2_X1 port map( A1 => n9559, A2 => n9558, Z => n18414);
   U15210 : NOR2_X1 port map( A1 => n18456, A2 => n11426, ZN => n5748);
   U15212 : INV_X2 port map( I => n5752, ZN => n15021);
   U15213 : INV_X2 port map( I => n5797, ZN => n7535);
   U15217 : XOR2_X1 port map( A1 => n7044, A2 => n1092, Z => n12182);
   U15218 : OR2_X1 port map( A1 => n26154, A2 => n10764, Z => n5762);
   U15219 : OR2_X1 port map( A1 => n17587, A2 => n27424, Z => n5763);
   U15229 : XOR2_X1 port map( A1 => n8861, A2 => n17135, Z => n5783);
   U15230 : XOR2_X1 port map( A1 => n16993, A2 => n17070, Z => n17135);
   U15231 : NAND2_X2 port map( A1 => n5786, A2 => n5784, ZN => n14213);
   U15232 : INV_X1 port map( I => n19639, ZN => n5786);
   U15235 : XOR2_X1 port map( A1 => n20438, A2 => n5793, Z => n5792);
   U15236 : XOR2_X1 port map( A1 => n20423, A2 => n24840, Z => n5793);
   U15241 : OAI21_X1 port map( A1 => n7017, A2 => n18005, B => n1780, ZN => 
                           n14317);
   U15244 : XOR2_X1 port map( A1 => Plaintext(109), A2 => Key(109), Z => n6603)
                           ;
   U15245 : NAND2_X1 port map( A1 => n5805, A2 => n28160, ZN => n18777);
   U15246 : XOR2_X1 port map( A1 => n19528, A2 => n595, Z => n8428);
   U15247 : XOR2_X1 port map( A1 => n19528, A2 => n603, Z => n9360);
   U15249 : XNOR2_X1 port map( A1 => n5808, A2 => n5809, ZN => n5807);
   U15251 : XOR2_X1 port map( A1 => n9279, A2 => n13195, Z => n5809);
   U15256 : XOR2_X1 port map( A1 => n17072, A2 => n5821, Z => n5820);
   U15257 : XOR2_X1 port map( A1 => n10999, A2 => n7355, Z => n5821);
   U15262 : AOI21_X2 port map( A1 => n21827, A2 => n13238, B => n5825, ZN => 
                           n18012);
   U15264 : XOR2_X1 port map( A1 => n22839, A2 => n18081, Z => n8955);
   U15265 : XOR2_X1 port map( A1 => n18238, A2 => n22673, Z => n7625);
   U15266 : XOR2_X1 port map( A1 => n19431, A2 => n5833, Z => n6349);
   U15267 : XOR2_X1 port map( A1 => n19406, A2 => n13001, Z => n19431);
   U15269 : XOR2_X1 port map( A1 => n19481, A2 => n5834, Z => n5833);
   U15270 : XOR2_X1 port map( A1 => n12612, A2 => n1314, Z => n5834);
   U15274 : NAND4_X1 port map( A1 => n10249, A2 => n8385, A3 => n12323, A4 => 
                           n8384, ZN => n5840);
   U15277 : INV_X2 port map( I => n5853, ZN => n16270);
   U15280 : XOR2_X1 port map( A1 => n26141, A2 => n20369, Z => n17119);
   U15281 : AND2_X1 port map( A1 => n14649, A2 => n24525, Z => n5860);
   U15286 : XOR2_X1 port map( A1 => n20422, A2 => n21926, Z => n5867);
   U15290 : XOR2_X1 port map( A1 => n5872, A2 => n5871, Z => n5870);
   U15298 : OAI21_X1 port map( A1 => n8045, A2 => n1166, B => n23844, ZN => 
                           n8044);
   U15305 : XOR2_X1 port map( A1 => n18103, A2 => n23186, Z => n5912);
   U15310 : INV_X2 port map( I => n18718, ZN => n13372);
   U15311 : INV_X2 port map( I => n5927, ZN => n16335);
   U15313 : XNOR2_X1 port map( A1 => Plaintext(145), A2 => Key(145), ZN => 
                           n5927);
   U15314 : XOR2_X1 port map( A1 => n17094, A2 => n16943, Z => n16779);
   U15316 : NAND2_X1 port map( A1 => n13614, A2 => n5931, ZN => n6693);
   U15317 : NAND2_X1 port map( A1 => n5934, A2 => n20186, ZN => n6692);
   U15324 : XOR2_X1 port map( A1 => n7751, A2 => n14549, Z => n5940);
   U15327 : INV_X2 port map( I => n5946, ZN => n17548);
   U15331 : XOR2_X1 port map( A1 => n12042, A2 => n5949, Z => n8489);
   U15332 : XOR2_X1 port map( A1 => n28521, A2 => n5949, Z => n15472);
   U15333 : XOR2_X1 port map( A1 => n23314, A2 => n5949, Z => n15015);
   U15334 : OAI21_X1 port map( A1 => n9855, A2 => n891, B => n5956, ZN => n5953
                           );
   U15335 : OR3_X1 port map( A1 => n9344, A2 => n891, A3 => n18101, Z => n5952)
                           ;
   U15339 : XOR2_X1 port map( A1 => n5963, A2 => n5965, Z => n5962);
   U15340 : XOR2_X1 port map( A1 => n17059, A2 => n27936, Z => n5963);
   U15341 : XOR2_X1 port map( A1 => n25386, A2 => n15669, Z => n5965);
   U15346 : NAND2_X2 port map( A1 => n6841, A2 => n6839, ZN => n6838);
   U15347 : NAND2_X1 port map( A1 => n5974, A2 => n25966, ZN => n13498);
   U15355 : NAND2_X1 port map( A1 => n18417, A2 => n875, ZN => n5981);
   U15357 : XOR2_X1 port map( A1 => n18280, A2 => n918, Z => n5988);
   U15359 : XOR2_X1 port map( A1 => Plaintext(142), A2 => Key(142), Z => n13417
                           );
   U15363 : XOR2_X1 port map( A1 => n20485, A2 => n19966, Z => n6001);
   U15372 : INV_X2 port map( I => n6014, ZN => n18556);
   U15375 : XOR2_X1 port map( A1 => n6123, A2 => n14652, Z => n6015);
   U15380 : XOR2_X1 port map( A1 => n1193, A2 => n27654, Z => n8203);
   U15381 : XOR2_X1 port map( A1 => n6024, A2 => n11555, Z => n11687);
   U15386 : INV_X2 port map( I => n7870, ZN => n10639);
   U15390 : NOR2_X1 port map( A1 => n23653, A2 => n6046, ZN => n13912);
   U15394 : NAND2_X1 port map( A1 => n754, A2 => n19750, ZN => n19762);
   U15400 : NAND3_X1 port map( A1 => n22824, A2 => n21292, A3 => n26913, ZN => 
                           n6091);
   U15401 : NAND2_X1 port map( A1 => n6066, A2 => n13888, ZN => n6065);
   U15403 : XOR2_X1 port map( A1 => n5224, A2 => n14491, Z => n6068);
   U15404 : XOR2_X1 port map( A1 => n9650, A2 => n6287, Z => n6071);
   U15411 : NAND2_X1 port map( A1 => n21989, A2 => n20151, ZN => n19817);
   U15416 : OAI22_X2 port map( A1 => n902, A2 => n17085, B1 => n5718, B2 => 
                           n14168, ZN => n6137);
   U15420 : XOR2_X1 port map( A1 => n27084, A2 => n14526, Z => n11972);
   U15421 : XOR2_X1 port map( A1 => n27084, A2 => n14633, Z => n13633);
   U15422 : INV_X2 port map( I => n7067, ZN => n10210);
   U15423 : XOR2_X1 port map( A1 => n6107, A2 => n6660, Z => n6106);
   U15424 : XOR2_X1 port map( A1 => n13071, A2 => n6652, Z => n6107);
   U15425 : NAND2_X2 port map( A1 => n6119, A2 => n6117, ZN => n16644);
   U15429 : XOR2_X1 port map( A1 => n16854, A2 => n16795, Z => n14336);
   U15431 : XOR2_X1 port map( A1 => n20376, A2 => n21642, Z => n6126);
   U15437 : XOR2_X1 port map( A1 => Plaintext(107), A2 => Key(107), Z => n6140)
                           ;
   U15438 : XOR2_X1 port map( A1 => n6135, A2 => n15684, Z => n6134);
   U15441 : XOR2_X1 port map( A1 => n13661, A2 => n12363, Z => n6138);
   U15442 : INV_X2 port map( I => n6140, ZN => n15330);
   U15444 : XOR2_X1 port map( A1 => n6148, A2 => n543, Z => n17414);
   U15445 : XOR2_X1 port map( A1 => n17033, A2 => n17034, Z => n6148);
   U15446 : NAND2_X1 port map( A1 => n21684, A2 => n2777, ZN => n6152);
   U15447 : NAND2_X1 port map( A1 => n6152, A2 => n2778, ZN => n6149);
   U15448 : XOR2_X1 port map( A1 => n6535, A2 => n20535, Z => n6154);
   U15451 : XOR2_X1 port map( A1 => n6158, A2 => n19250, Z => n6157);
   U15454 : NAND2_X1 port map( A1 => n20031, A2 => n20171, ZN => n6162);
   U15456 : XOR2_X1 port map( A1 => n8293, A2 => n14876, Z => n9598);
   U15458 : NAND3_X1 port map( A1 => n25927, A2 => n9567, A3 => n953, ZN => 
                           n8765);
   U15459 : XOR2_X1 port map( A1 => n6168, A2 => n25351, Z => n6288);
   U15460 : XOR2_X1 port map( A1 => n18331, A2 => n6289, Z => n6168);
   U15464 : XOR2_X1 port map( A1 => n6176, A2 => n16583, Z => n6175);
   U15465 : XOR2_X1 port map( A1 => n28373, A2 => n20707, Z => n6176);
   U15466 : INV_X1 port map( I => Plaintext(105), ZN => n6177);
   U15467 : XOR2_X1 port map( A1 => n6177, A2 => Key(105), Z => n6434);
   U15469 : NOR2_X1 port map( A1 => n21653, A2 => n6182, ZN => n8753);
   U15470 : XOR2_X1 port map( A1 => n7752, A2 => n6186, Z => n19024);
   U15472 : INV_X2 port map( I => n15884, ZN => n16189);
   U15474 : AOI21_X1 port map( A1 => n20609, A2 => n842, B => n6247, ZN => 
                           n6925);
   U15480 : XOR2_X1 port map( A1 => n1134, A2 => n19434, Z => n6218);
   U15481 : INV_X2 port map( I => n6457, ZN => n6219);
   U15484 : OAI22_X1 port map( A1 => n9836, A2 => n27471, B1 => n27407, B2 => 
                           n8771, ZN => n15520);
   U15490 : INV_X2 port map( I => n6229, ZN => n14423);
   U15495 : XOR2_X1 port map( A1 => n7050, A2 => n14587, Z => n8195);
   U15501 : INV_X2 port map( I => n6259, ZN => n15586);
   U15506 : XOR2_X1 port map( A1 => n28407, A2 => n1297, Z => n6271);
   U15508 : XOR2_X1 port map( A1 => n6274, A2 => n6679, Z => n6678);
   U15510 : INV_X1 port map( I => n11984, ZN => n6277);
   U15514 : NAND2_X2 port map( A1 => n7447, A2 => n7450, ZN => n9051);
   U15521 : XOR2_X1 port map( A1 => n6298, A2 => n6297, Z => n6296);
   U15522 : XOR2_X1 port map( A1 => n16991, A2 => n21703, Z => n6297);
   U15523 : XOR2_X1 port map( A1 => n13852, A2 => n16993, Z => n6298);
   U15525 : NAND2_X1 port map( A1 => n18912, A2 => n26645, ZN => n14201);
   U15529 : AOI21_X1 port map( A1 => n22910, A2 => n6837, B => n16266, ZN => 
                           n16268);
   U15533 : NAND2_X1 port map( A1 => n21387, A2 => n22421, ZN => n6319);
   U15538 : XOR2_X1 port map( A1 => n18050, A2 => n13978, Z => n18773);
   U15539 : XOR2_X1 port map( A1 => n7338, A2 => n20671, Z => n18049);
   U15556 : XOR2_X1 port map( A1 => n19421, A2 => n6275, Z => n18519);
   U15562 : NAND3_X1 port map( A1 => n9379, A2 => n23096, A3 => n24334, ZN => 
                           n9111);
   U15565 : XOR2_X1 port map( A1 => n20384, A2 => n13288, Z => n6377);
   U15567 : XOR2_X1 port map( A1 => n6380, A2 => n6382, Z => n6379);
   U15568 : XOR2_X1 port map( A1 => n23137, A2 => n6381, Z => n6380);
   U15569 : XOR2_X1 port map( A1 => n19551, A2 => n6385, Z => n6384);
   U15570 : XOR2_X1 port map( A1 => n19392, A2 => n21077, Z => n6385);
   U15571 : XOR2_X1 port map( A1 => n5351, A2 => n8657, Z => n19551);
   U15572 : XOR2_X1 port map( A1 => n19183, A2 => n6387, Z => n6386);
   U15573 : XNOR2_X1 port map( A1 => n25166, A2 => n25376, ZN => n6387);
   U15584 : XOR2_X1 port map( A1 => n26029, A2 => n21153, Z => n20720);
   U15588 : XOR2_X1 port map( A1 => Plaintext(111), A2 => Key(111), Z => n16288
                           );
   U15591 : NOR2_X1 port map( A1 => n4315, A2 => n22764, ZN => n6432);
   U15592 : INV_X2 port map( I => n6434, ZN => n15885);
   U15596 : NOR2_X1 port map( A1 => n821, A2 => n15623, ZN => n6442);
   U15601 : XOR2_X1 port map( A1 => n19503, A2 => n6453, Z => n6452);
   U15602 : XOR2_X1 port map( A1 => n4175, A2 => n21733, Z => n6453);
   U15604 : XOR2_X1 port map( A1 => n9900, A2 => n6456, Z => n7385);
   U15605 : XOR2_X1 port map( A1 => n19529, A2 => n19559, Z => n19434);
   U15606 : AOI21_X2 port map( A1 => n6463, A2 => n8473, B => n6460, ZN => 
                           n6459);
   U15608 : NAND2_X2 port map( A1 => n766, A2 => n28025, ZN => n17468);
   U15611 : XOR2_X1 port map( A1 => n12202, A2 => n5147, Z => n6475);
   U15612 : NAND2_X2 port map( A1 => n12421, A2 => n13586, ZN => n6562);
   U15615 : NAND2_X2 port map( A1 => n6789, A2 => n6786, ZN => n6485);
   U15621 : XOR2_X1 port map( A1 => n8424, A2 => n16856, Z => n6500);
   U15622 : NAND2_X1 port map( A1 => n7750, A2 => n6501, ZN => n11229);
   U15629 : XOR2_X1 port map( A1 => n16874, A2 => n16752, Z => n6515);
   U15632 : NOR2_X1 port map( A1 => n28499, A2 => n12111, ZN => n14036);
   U15635 : XOR2_X1 port map( A1 => n6528, A2 => n4076, Z => n13785);
   U15636 : XOR2_X1 port map( A1 => n6528, A2 => n24121, Z => n18951);
   U15637 : INV_X1 port map( I => n19861, ZN => n6529);
   U15641 : XOR2_X1 port map( A1 => n8983, A2 => n6536, Z => n9860);
   U15642 : XOR2_X1 port map( A1 => n24577, A2 => n10339, Z => n6536);
   U15643 : XOR2_X1 port map( A1 => n6539, A2 => n6541, Z => n8736);
   U15644 : XOR2_X1 port map( A1 => n22123, A2 => n5147, Z => n6541);
   U15650 : INV_X2 port map( I => n15696, ZN => n6547);
   U15651 : XOR2_X1 port map( A1 => n12322, A2 => n6550, Z => n7303);
   U15652 : XOR2_X1 port map( A1 => n11124, A2 => n16938, Z => n6550);
   U15655 : XOR2_X1 port map( A1 => n6554, A2 => n925, Z => n10311);
   U15656 : XOR2_X1 port map( A1 => n6554, A2 => n18234, Z => n18235);
   U15659 : XOR2_X1 port map( A1 => n19352, A2 => n19521, Z => n19460);
   U15661 : NAND3_X1 port map( A1 => n24078, A2 => n20516, A3 => n28016, ZN => 
                           n8700);
   U15665 : MUX2_X1 port map( I0 => n14671, I1 => n24997, S => n19630, Z => 
                           n6561);
   U15666 : XOR2_X1 port map( A1 => n25306, A2 => n14630, Z => n6563);
   U15667 : NOR2_X2 port map( A1 => n21622, A2 => n21621, ZN => n21626);
   U15671 : INV_X2 port map( I => n6574, ZN => n17324);
   U15677 : XOR2_X1 port map( A1 => n19333, A2 => n8322, Z => n19039);
   U15686 : XOR2_X1 port map( A1 => n4833, A2 => n28186, Z => n6594);
   U15687 : XOR2_X1 port map( A1 => n3390, A2 => n21261, Z => n6595);
   U15688 : INV_X1 port map( I => n20376, ZN => n20508);
   U15696 : XOR2_X1 port map( A1 => n18273, A2 => n8329, Z => n6614);
   U15697 : XOR2_X1 port map( A1 => n18274, A2 => n18272, Z => n6615);
   U15700 : NAND2_X1 port map( A1 => n9051, A2 => n23072, ZN => n6621);
   U15701 : NOR2_X1 port map( A1 => n17722, A2 => n17723, ZN => n6630);
   U15706 : XNOR2_X1 port map( A1 => n6638, A2 => n16885, ZN => n6637);
   U15708 : INV_X2 port map( I => n6640, ZN => n8968);
   U15709 : XOR2_X1 port map( A1 => n12242, A2 => n12771, Z => n19548);
   U15711 : XOR2_X1 port map( A1 => n27438, A2 => n20383, Z => n15711);
   U15713 : NAND2_X2 port map( A1 => n15722, A2 => n16828, ZN => n17992);
   U15718 : XOR2_X1 port map( A1 => n22792, A2 => n14614, Z => n6660);
   U15722 : INV_X2 port map( I => n9001, ZN => n20868);
   U15727 : NAND2_X1 port map( A1 => n1109, A2 => n23120, ZN => n10227);
   U15729 : XOR2_X1 port map( A1 => n17106, A2 => n21820, Z => n6673);
   U15730 : XOR2_X1 port map( A1 => n27564, A2 => n1283, Z => n8954);
   U15731 : XOR2_X1 port map( A1 => n6675, A2 => n1295, Z => n10996);
   U15732 : XOR2_X1 port map( A1 => n27564, A2 => n18290, Z => n18291);
   U15733 : XOR2_X1 port map( A1 => n280, A2 => n27564, Z => n12601);
   U15736 : INV_X2 port map( I => n6678, ZN => n14671);
   U15737 : XOR2_X1 port map( A1 => n19202, A2 => n6680, Z => n6679);
   U15738 : XOR2_X1 port map( A1 => n13906, A2 => n19522, Z => n6680);
   U15742 : XOR2_X1 port map( A1 => n16959, A2 => n11684, Z => n16848);
   U15743 : XOR2_X1 port map( A1 => n16959, A2 => n12204, Z => n17153);
   U15747 : OAI21_X2 port map( A1 => n10532, A2 => n21512, B => n6700, ZN => 
                           n21342);
   U15749 : INV_X2 port map( I => n6703, ZN => n12225);
   U15750 : XOR2_X1 port map( A1 => n17141, A2 => n1319, Z => n6704);
   U15755 : AOI22_X1 port map( A1 => n17598, A2 => n17981, B1 => n26076, B2 => 
                           n23963, ZN => n17599);
   U15756 : XOR2_X1 port map( A1 => n18215, A2 => n14596, Z => n10754);
   U15763 : XOR2_X1 port map( A1 => n6737, A2 => n10179, Z => n6736);
   U15764 : XOR2_X1 port map( A1 => n6941, A2 => n20421, Z => n6739);
   U15767 : XOR2_X1 port map( A1 => n18047, A2 => n6745, Z => n18322);
   U15775 : XOR2_X1 port map( A1 => n15639, A2 => n1061, Z => n6748);
   U15777 : XOR2_X1 port map( A1 => n6753, A2 => n6752, Z => n6751);
   U15778 : XOR2_X1 port map( A1 => n19512, A2 => n13787, Z => n6752);
   U15781 : INV_X1 port map( I => n24639, ZN => n6758);
   U15783 : XOR2_X1 port map( A1 => n21373, A2 => n9397, Z => n20454);
   U15785 : NAND3_X2 port map( A1 => n11210, A2 => n11691, A3 => n20184, ZN => 
                           n21373);
   U15786 : NAND2_X1 port map( A1 => n16678, A2 => n6763, ZN => n13881);
   U15794 : INV_X1 port map( I => n9920, ZN => n6775);
   U15800 : NOR2_X1 port map( A1 => n6780, A2 => n19734, ZN => n13722);
   U15802 : MUX2_X1 port map( I0 => n11902, I1 => n13250, S => n10031, Z => 
                           n6789);
   U15803 : XOR2_X1 port map( A1 => n10839, A2 => n6790, Z => n10838);
   U15804 : XOR2_X1 port map( A1 => n6791, A2 => n6792, Z => n6790);
   U15805 : XOR2_X1 port map( A1 => n14744, A2 => n767, Z => n6791);
   U15806 : XOR2_X1 port map( A1 => n24885, A2 => n14340, Z => n6792);
   U15807 : XOR2_X1 port map( A1 => n4501, A2 => n21262, Z => n21263);
   U15808 : XOR2_X1 port map( A1 => n6795, A2 => n21533, Z => Ciphertext(148));
   U15810 : NAND2_X1 port map( A1 => n10763, A2 => n6803, ZN => n13169);
   U15812 : NOR2_X1 port map( A1 => n12016, A2 => n6803, ZN => n7347);
   U15813 : AOI21_X1 port map( A1 => n21710, A2 => n13718, B => n6803, ZN => 
                           n15705);
   U15814 : NOR2_X2 port map( A1 => n6805, A2 => n6804, ZN => n8672);
   U15815 : XOR2_X1 port map( A1 => n2507, A2 => n19346, Z => n10615);
   U15816 : NAND2_X1 port map( A1 => n20219, A2 => n27010, ZN => n20053);
   U15820 : INV_X2 port map( I => n6822, ZN => n6861);
   U15822 : XOR2_X1 port map( A1 => n11460, A2 => n13512, Z => n6823);
   U15824 : NAND2_X1 port map( A1 => n17312, A2 => n14578, ZN => n6825);
   U15825 : INV_X1 port map( I => n6826, ZN => n7784);
   U15826 : NAND2_X1 port map( A1 => n17419, A2 => n15529, ZN => n6826);
   U15833 : NOR2_X2 port map( A1 => n6858, A2 => n6857, ZN => n11819);
   U15835 : NAND2_X1 port map( A1 => n6487, A2 => n19155, ZN => n18908);
   U15836 : XOR2_X1 port map( A1 => n21179, A2 => n6864, Z => n10927);
   U15837 : NOR2_X1 port map( A1 => n18590, A2 => n1011, ZN => n13765);
   U15838 : XOR2_X1 port map( A1 => n19504, A2 => n12015, Z => n6866);
   U15839 : XOR2_X1 port map( A1 => n6868, A2 => n6869, Z => n6870);
   U15841 : XOR2_X1 port map( A1 => n17051, A2 => n554, Z => n6869);
   U15843 : XOR2_X1 port map( A1 => n27624, A2 => n13001, Z => n8216);
   U15844 : XOR2_X1 port map( A1 => n27624, A2 => n19563, Z => n12110);
   U15845 : XOR2_X1 port map( A1 => n27396, A2 => n21305, Z => n20532);
   U15846 : XOR2_X1 port map( A1 => n20568, A2 => n11071, Z => n6871);
   U15852 : XNOR2_X1 port map( A1 => Plaintext(18), A2 => Key(18), ZN => n6886)
                           ;
   U15854 : NAND2_X2 port map( A1 => n17001, A2 => n17000, ZN => n17917);
   U15855 : NAND2_X2 port map( A1 => n6894, A2 => n6893, ZN => n20222);
   U15856 : NAND2_X2 port map( A1 => n20138, A2 => n19999, ZN => n20223);
   U15857 : NAND3_X1 port map( A1 => n11805, A2 => n25279, A3 => n19941, ZN => 
                           n6895);
   U15859 : NOR2_X1 port map( A1 => n6898, A2 => n16679, ZN => n16048);
   U15869 : XOR2_X1 port map( A1 => n6921, A2 => n20727, Z => Ciphertext(4));
   U15877 : XOR2_X1 port map( A1 => n14980, A2 => n18312, Z => n6943);
   U15878 : XOR2_X1 port map( A1 => n25391, A2 => n15494, Z => n6944);
   U15886 : XOR2_X1 port map( A1 => n7762, A2 => n6951, Z => n17446);
   U15890 : NOR2_X1 port map( A1 => n21535, A2 => n21531, ZN => n6957);
   U15891 : XOR2_X1 port map( A1 => n6960, A2 => n14851, Z => n14848);
   U15892 : XOR2_X1 port map( A1 => n8664, A2 => n15385, Z => n8663);
   U15896 : NAND2_X1 port map( A1 => n21535, A2 => n21534, ZN => n6972);
   U15899 : NAND3_X1 port map( A1 => n10210, A2 => n14666, A3 => n20865, ZN => 
                           n20464);
   U15900 : XOR2_X1 port map( A1 => n18069, A2 => n18070, Z => n18347);
   U15901 : AOI21_X2 port map( A1 => n17995, A2 => n17994, B => n11283, ZN => 
                           n18069);
   U15902 : INV_X1 port map( I => n16214, ZN => n7968);
   U15903 : AND2_X1 port map( A1 => n11175, A2 => n19822, Z => n10761);
   U15910 : XOR2_X1 port map( A1 => n17063, A2 => n6984, Z => n6983);
   U15912 : NOR2_X1 port map( A1 => n10585, A2 => n13933, ZN => n13932);
   U15915 : XOR2_X1 port map( A1 => n19549, A2 => n6986, Z => n6985);
   U15917 : XOR2_X1 port map( A1 => n12410, A2 => n1300, Z => n11312);
   U15920 : NAND2_X1 port map( A1 => n11847, A2 => n11846, ZN => n8894);
   U15921 : NAND2_X1 port map( A1 => n8894, A2 => n20149, ZN => n8893);
   U15929 : XOR2_X1 port map( A1 => n6997, A2 => n15149, Z => Ciphertext(21));
   U15931 : NAND3_X1 port map( A1 => n9728, A2 => n27923, A3 => n27416, ZN => 
                           n7000);
   U15934 : OAI21_X2 port map( A1 => n9677, A2 => n8419, B => n21070, ZN => 
                           n8069);
   U15939 : XOR2_X1 port map( A1 => n9749, A2 => n18210, Z => n9745);
   U15940 : NOR2_X1 port map( A1 => n25363, A2 => n27631, ZN => n8624);
   U15941 : XOR2_X1 port map( A1 => n15795, A2 => Key(177), Z => n10035);
   U15943 : NOR2_X1 port map( A1 => n21668, A2 => n21667, ZN => n11760);
   U15944 : AOI21_X1 port map( A1 => n16317, A2 => n16321, B => n7007, ZN => 
                           n7219);
   U15948 : XOR2_X1 port map( A1 => n10056, A2 => n20208, Z => n13890);
   U15950 : OR2_X1 port map( A1 => n10610, A2 => n20593, Z => n9564);
   U15953 : XOR2_X1 port map( A1 => n18059, A2 => n12302, Z => n7010);
   U15956 : NOR2_X1 port map( A1 => n18627, A2 => n820, ZN => n14300);
   U15962 : OAI22_X2 port map( A1 => n8088, A2 => n8087, B1 => n15686, B2 => 
                           n16139, ZN => n8084);
   U15966 : XOR2_X1 port map( A1 => n10319, A2 => n10317, Z => n19741);
   U15967 : NAND2_X1 port map( A1 => n8702, A2 => n11047, ZN => n15600);
   U15976 : XOR2_X1 port map( A1 => n11176, A2 => n11178, Z => n7025);
   U15979 : NAND3_X1 port map( A1 => n13444, A2 => n25342, A3 => n21116, ZN => 
                           n21121);
   U15981 : XOR2_X1 port map( A1 => n18226, A2 => n18225, Z => n7027);
   U15983 : INV_X2 port map( I => n7029, ZN => n9896);
   U15989 : XOR2_X1 port map( A1 => n17082, A2 => n13633, Z => n7031);
   U15990 : NOR2_X1 port map( A1 => n8717, A2 => n14393, ZN => n7036);
   U15991 : XOR2_X1 port map( A1 => n10995, A2 => n10997, Z => n14414);
   U15993 : XOR2_X1 port map( A1 => n19387, A2 => n13624, Z => n9545);
   U16002 : AND2_X1 port map( A1 => n10894, A2 => n21765, Z => n10693);
   U16008 : NAND2_X1 port map( A1 => n12212, A2 => n12211, ZN => n12210);
   U16012 : XOR2_X1 port map( A1 => n10933, A2 => n10935, Z => n15344);
   U16019 : NOR2_X1 port map( A1 => n21501, A2 => n14634, ZN => n7116);
   U16020 : AND3_X2 port map( A1 => n21550, A2 => n21552, A3 => n21551, Z => 
                           n7085);
   U16022 : NAND2_X2 port map( A1 => n10385, A2 => n24574, ZN => n12270);
   U16023 : OR2_X1 port map( A1 => n2813, A2 => n361, Z => n7088);
   U16026 : NAND2_X2 port map( A1 => n7090, A2 => n9735, ZN => n18063);
   U16028 : NOR2_X1 port map( A1 => n13198, A2 => n12765, ZN => n13197);
   U16034 : XOR2_X1 port map( A1 => n21819, A2 => n16803, Z => n7097);
   U16035 : XOR2_X1 port map( A1 => n11644, A2 => n7106, Z => n9129);
   U16044 : XOR2_X1 port map( A1 => n21238, A2 => n13114, Z => n13113);
   U16046 : OR2_X1 port map( A1 => n17530, A2 => n17196, Z => n7363);
   U16049 : XOR2_X1 port map( A1 => n9998, A2 => n16848, Z => n16851);
   U16056 : XOR2_X1 port map( A1 => n16764, A2 => n545, Z => n8238);
   U16057 : OAI22_X1 port map( A1 => n11741, A2 => n21473, B1 => n6517, B2 => 
                           n10833, ZN => n10832);
   U16059 : XOR2_X1 port map( A1 => n7145, A2 => n1061, Z => Ciphertext(145));
   U16064 : XOR2_X1 port map( A1 => n11787, A2 => n21707, Z => n14775);
   U16069 : NOR2_X1 port map( A1 => n15295, A2 => n19872, ZN => n11474);
   U16072 : XOR2_X1 port map( A1 => n18351, A2 => n7154, Z => n13818);
   U16073 : XOR2_X1 port map( A1 => n7338, A2 => n8332, Z => n7154);
   U16082 : XNOR2_X1 port map( A1 => n12823, A2 => n18121, ZN => n7170);
   U16085 : XOR2_X1 port map( A1 => n15708, A2 => n7397, Z => n8042);
   U16097 : XOR2_X1 port map( A1 => n7717, A2 => n7170, Z => n14369);
   U16101 : AND2_X1 port map( A1 => n2952, A2 => n27699, Z => n17616);
   U16102 : INV_X1 port map( I => n27573, ZN => n7878);
   U16103 : OR2_X1 port map( A1 => n14126, A2 => n10046, Z => n7798);
   U16114 : NAND2_X1 port map( A1 => n10000, A2 => n20684, ZN => n20688);
   U16115 : XNOR2_X1 port map( A1 => n5379, A2 => n20880, ZN => n13404);
   U16116 : XOR2_X1 port map( A1 => Plaintext(4), A2 => Key(4), Z => n15892);
   U16117 : NAND2_X2 port map( A1 => n7185, A2 => n10652, ZN => n13548);
   U16118 : INV_X2 port map( I => n7189, ZN => n12699);
   U16120 : NOR2_X1 port map( A1 => n11011, A2 => n11012, ZN => n7193);
   U16130 : XOR2_X1 port map( A1 => n8825, A2 => n7203, Z => n8824);
   U16131 : XOR2_X1 port map( A1 => n7204, A2 => n19039, Z => n7203);
   U16141 : OAI21_X2 port map( A1 => n699, A2 => n16819, B => n9542, ZN => 
                           n8089);
   U16146 : XOR2_X1 port map( A1 => n7218, A2 => n17058, Z => n7482);
   U16149 : XOR2_X1 port map( A1 => n18273, A2 => n823, Z => n7222);
   U16150 : AOI22_X2 port map( A1 => n20892, A2 => n20893, B1 => n21025, B2 => 
                           n20891, ZN => n20917);
   U16151 : XOR2_X1 port map( A1 => n7223, A2 => n20909, Z => Ciphertext(56));
   U16154 : XOR2_X1 port map( A1 => n15043, A2 => n7224, Z => n13223);
   U16155 : XOR2_X1 port map( A1 => n17084, A2 => n7225, Z => n7224);
   U16159 : INV_X1 port map( I => n8151, ZN => n7443);
   U16162 : XOR2_X1 port map( A1 => n23053, A2 => n14556, Z => n7231);
   U16167 : XOR2_X1 port map( A1 => n8800, A2 => n8331, Z => n7240);
   U16170 : INV_X2 port map( I => n7242, ZN => n10150);
   U16175 : XOR2_X1 port map( A1 => n19536, A2 => n27352, Z => n7250);
   U16179 : XOR2_X1 port map( A1 => n9981, A2 => n686, Z => n14715);
   U16180 : XOR2_X1 port map( A1 => n11838, A2 => n7252, Z => n8637);
   U16185 : NAND2_X1 port map( A1 => n16036, A2 => n25017, ZN => n7255);
   U16186 : INV_X2 port map( I => n10914, ZN => n18293);
   U16189 : XOR2_X1 port map( A1 => n7258, A2 => n11288, Z => Ciphertext(6));
   U16190 : AOI22_X1 port map( A1 => n20613, A2 => n20612, B1 => n4820, B2 => 
                           n20628, ZN => n7258);
   U16191 : NAND2_X1 port map( A1 => n21622, A2 => n14406, ZN => n13096);
   U16194 : INV_X1 port map( I => n9759, ZN => n16729);
   U16197 : OR2_X1 port map( A1 => n16407, A2 => n265, Z => n11495);
   U16199 : XOR2_X1 port map( A1 => Plaintext(148), A2 => Key(148), Z => n8406)
                           ;
   U16200 : XOR2_X1 port map( A1 => n16907, A2 => n560, Z => n7264);
   U16201 : OAI22_X1 port map( A1 => n15348, A2 => n14423, B1 => n19694, B2 => 
                           n12256, ZN => n19639);
   U16206 : XOR2_X1 port map( A1 => n2505, A2 => n19511, Z => n7268);
   U16213 : CLKBUF_X2 port map( I => Key(161), Z => n20877);
   U16216 : INV_X2 port map( I => n15431, ZN => n18352);
   U16218 : INV_X1 port map( I => n7271, ZN => n10531);
   U16219 : AOI21_X1 port map( A1 => n8340, A2 => n14908, B => n16731, ZN => 
                           n7271);
   U16220 : OR2_X1 port map( A1 => n14183, A2 => n14666, Z => n20867);
   U16224 : NAND2_X2 port map( A1 => n14182, A2 => n20870, ZN => n20879);
   U16225 : OAI21_X1 port map( A1 => n8021, A2 => n16455, B => n7237, ZN => 
                           n12483);
   U16238 : NAND3_X1 port map( A1 => n9319, A2 => n27411, A3 => n21655, ZN => 
                           n9318);
   U16242 : AOI21_X1 port map( A1 => n20280, A2 => n22786, B => n7749, ZN => 
                           n7930);
   U16243 : NAND2_X2 port map( A1 => n7819, A2 => n7294, ZN => n20165);
   U16249 : XOR2_X1 port map( A1 => n11279, A2 => n11276, Z => n7301);
   U16252 : XOR2_X1 port map( A1 => n7305, A2 => n24711, Z => Ciphertext(36));
   U16253 : AOI22_X1 port map( A1 => n20793, A2 => n11147, B1 => n22536, B2 => 
                           n20792, ZN => n7305);
   U16255 : OR2_X1 port map( A1 => n20142, A2 => n20107, Z => n12801);
   U16256 : INV_X2 port map( I => n7307, ZN => n14745);
   U16261 : XOR2_X1 port map( A1 => n21428, A2 => n21427, Z => n7315);
   U16262 : XOR2_X1 port map( A1 => n13557, A2 => n7317, Z => n17193);
   U16263 : XOR2_X1 port map( A1 => n16747, A2 => n16748, Z => n7317);
   U16267 : XOR2_X1 port map( A1 => n10364, A2 => n7320, Z => n10363);
   U16269 : XOR2_X1 port map( A1 => n10075, A2 => n17135, Z => n11845);
   U16275 : NOR2_X1 port map( A1 => n12272, A2 => n10866, ZN => n10865);
   U16279 : NAND2_X1 port map( A1 => n10230, A2 => n14520, ZN => n7332);
   U16280 : NOR2_X1 port map( A1 => n12598, A2 => n21020, ZN => n10661);
   U16281 : XOR2_X1 port map( A1 => n7336, A2 => n22512, Z => Ciphertext(13));
   U16289 : XOR2_X1 port map( A1 => n21418, A2 => n7339, Z => n13180);
   U16290 : XOR2_X1 port map( A1 => n12181, A2 => n21302, Z => n7339);
   U16295 : XOR2_X1 port map( A1 => n7346, A2 => n19302, Z => n19058);
   U16296 : INV_X2 port map( I => n13022, ZN => n10558);
   U16297 : XOR2_X1 port map( A1 => n684, A2 => n9860, Z => n13022);
   U16302 : INV_X1 port map( I => n16272, ZN => n10427);
   U16314 : NOR2_X1 port map( A1 => n16067, A2 => n9768, ZN => n10507);
   U16315 : AND2_X1 port map( A1 => n15003, A2 => n20777, Z => n10350);
   U16316 : XOR2_X1 port map( A1 => n17123, A2 => n17154, Z => n12342);
   U16323 : OAI21_X1 port map( A1 => n16617, A2 => n15813, B => n11005, ZN => 
                           n15816);
   U16330 : OAI21_X1 port map( A1 => n13774, A2 => n11767, B => n11764, ZN => 
                           n12788);
   U16335 : XOR2_X1 port map( A1 => n18330, A2 => n14506, Z => n7375);
   U16338 : XNOR2_X1 port map( A1 => n16817, A2 => n17070, ZN => n10195);
   U16343 : OAI21_X1 port map( A1 => n16488, A2 => n25875, B => n24089, ZN => 
                           n8532);
   U16345 : NOR3_X1 port map( A1 => n21032, A2 => n21031, A3 => n21045, ZN => 
                           n21034);
   U16349 : INV_X2 port map( I => n14348, ZN => n21275);
   U16350 : OAI21_X1 port map( A1 => n21217, A2 => n22027, B => n12394, ZN => 
                           n21219);
   U16355 : NOR2_X1 port map( A1 => n7460, A2 => n921, ZN => n7398);
   U16356 : AND2_X1 port map( A1 => n5425, A2 => n12257, Z => n11410);
   U16358 : OAI21_X1 port map( A1 => n11490, A2 => n21590, B => n14679, ZN => 
                           n21442);
   U16359 : OR2_X1 port map( A1 => n10851, A2 => n27431, Z => n13974);
   U16361 : OAI21_X2 port map( A1 => n9965, A2 => n13282, B => n13957, ZN => 
                           n7652);
   U16368 : NAND2_X1 port map( A1 => n9050, A2 => n11485, ZN => n7420);
   U16371 : XOR2_X1 port map( A1 => n7425, A2 => n611, Z => n7424);
   U16374 : XOR2_X1 port map( A1 => n14675, A2 => n21900, Z => n7435);
   U16375 : NAND2_X2 port map( A1 => n19839, A2 => n756, ZN => n19675);
   U16377 : INV_X2 port map( I => n12220, ZN => n8254);
   U16378 : XOR2_X1 port map( A1 => n22780, A2 => n13669, Z => n8597);
   U16381 : OR2_X1 port map( A1 => n7265, A2 => n26039, Z => n7466);
   U16382 : XOR2_X1 port map( A1 => n7467, A2 => n9582, Z => n7588);
   U16383 : XOR2_X1 port map( A1 => n11550, A2 => n11549, Z => n7471);
   U16385 : XOR2_X1 port map( A1 => n7475, A2 => n18108, Z => n7474);
   U16389 : AND2_X1 port map( A1 => n18091, A2 => n28105, Z => n9222);
   U16391 : XNOR2_X1 port map( A1 => Plaintext(27), A2 => Key(27), ZN => n7486)
                           ;
   U16392 : NOR2_X1 port map( A1 => n7487, A2 => n14137, ZN => n15813);
   U16407 : NAND2_X1 port map( A1 => n7515, A2 => n20750, ZN => n7513);
   U16408 : AOI21_X1 port map( A1 => n20711, A2 => n12416, B => n20749, ZN => 
                           n7514);
   U16411 : NAND3_X1 port map( A1 => n19227, A2 => n18826, A3 => n19451, ZN => 
                           n7522);
   U16416 : XOR2_X1 port map( A1 => n370, A2 => n24312, Z => n7529);
   U16417 : OR2_X1 port map( A1 => n5990, A2 => n23772, Z => n10735);
   U16418 : NOR2_X2 port map( A1 => n8086, A2 => n8085, ZN => n16699);
   U16421 : INV_X2 port map( I => n10078, ZN => n16910);
   U16422 : NAND2_X2 port map( A1 => n7543, A2 => n7541, ZN => n10078);
   U16425 : XOR2_X1 port map( A1 => n26719, A2 => n18076, Z => n7545);
   U16427 : XOR2_X1 port map( A1 => n7244, A2 => n1296, Z => n7547);
   U16429 : XOR2_X1 port map( A1 => n12816, A2 => n7552, Z => n11450);
   U16430 : XOR2_X1 port map( A1 => n12042, A2 => n27366, Z => n7552);
   U16431 : NAND2_X1 port map( A1 => n21706, A2 => n6802, ZN => n9910);
   U16432 : OAI21_X1 port map( A1 => n9065, A2 => n3325, B => n20873, ZN => 
                           n7554);
   U16433 : NAND2_X1 port map( A1 => n7557, A2 => n7556, ZN => n7555);
   U16434 : NOR2_X1 port map( A1 => n3325, A2 => n20873, ZN => n7556);
   U16435 : INV_X1 port map( I => n9065, ZN => n7557);
   U16436 : XOR2_X1 port map( A1 => n9063, A2 => n14638, Z => n13579);
   U16439 : XOR2_X1 port map( A1 => n7563, A2 => n20354, Z => n7560);
   U16441 : NAND2_X2 port map( A1 => n7565, A2 => n18426, ZN => n9642);
   U16442 : OAI21_X2 port map( A1 => n9604, A2 => n10116, B => n10929, ZN => 
                           n18426);
   U16443 : XOR2_X1 port map( A1 => Plaintext(46), A2 => Key(46), Z => n16120);
   U16447 : INV_X2 port map( I => n7571, ZN => n17479);
   U16450 : XNOR2_X1 port map( A1 => n7583, A2 => n10945, ZN => n7582);
   U16451 : XOR2_X1 port map( A1 => n19488, A2 => n12623, Z => n7583);
   U16458 : OR3_X1 port map( A1 => n8120, A2 => n14457, A3 => n8121, Z => n7595
                           );
   U16460 : NAND2_X2 port map( A1 => n7596, A2 => n9562, ZN => n10337);
   U16463 : XOR2_X1 port map( A1 => n16873, A2 => n13945, Z => n7605);
   U16467 : NAND2_X2 port map( A1 => n7616, A2 => n7613, ZN => n18142);
   U16468 : INV_X1 port map( I => n12809, ZN => n15554);
   U16477 : INV_X2 port map( I => n7638, ZN => n10588);
   U16478 : XOR2_X1 port map( A1 => n17970, A2 => n7408, Z => n8689);
   U16479 : XOR2_X1 port map( A1 => n7640, A2 => n7639, Z => n14302);
   U16485 : XOR2_X1 port map( A1 => n7655, A2 => n20352, Z => n7654);
   U16486 : XOR2_X1 port map( A1 => n22756, A2 => n28278, Z => n7655);
   U16487 : XOR2_X1 port map( A1 => n7658, A2 => n7660, Z => n19757);
   U16490 : NAND2_X1 port map( A1 => n9979, A2 => n10512, ZN => n7663);
   U16491 : XOR2_X1 port map( A1 => n17046, A2 => n7665, Z => n7664);
   U16492 : XOR2_X1 port map( A1 => n7786, A2 => n21607, Z => n7665);
   U16502 : XOR2_X1 port map( A1 => n7386, A2 => n11183, Z => n13348);
   U16505 : XOR2_X1 port map( A1 => n19503, A2 => n19502, Z => n7679);
   U16507 : OAI21_X1 port map( A1 => n14557, A2 => n16314, B => n16316, ZN => 
                           n15783);
   U16508 : AOI22_X1 port map( A1 => n16239, A2 => n16315, B1 => n16316, B2 => 
                           n16241, ZN => n8687);
   U16510 : OAI22_X2 port map( A1 => n7695, A2 => n7693, B1 => n10141, B2 => 
                           n7694, ZN => n17757);
   U16511 : XOR2_X1 port map( A1 => n7697, A2 => n7696, Z => n7760);
   U16512 : XOR2_X1 port map( A1 => n14203, A2 => n21613, Z => n7696);
   U16513 : XOR2_X1 port map( A1 => n11261, A2 => n13840, Z => n7697);
   U16517 : INV_X2 port map( I => n7700, ZN => n17403);
   U16518 : XOR2_X1 port map( A1 => n7707, A2 => n17085, Z => n7709);
   U16522 : XOR2_X1 port map( A1 => n17064, A2 => n7711, Z => n7710);
   U16523 : XOR2_X1 port map( A1 => n26038, A2 => n10294, Z => n7711);
   U16525 : XOR2_X1 port map( A1 => n20532, A2 => n7714, Z => n7713);
   U16526 : XOR2_X1 port map( A1 => n5082, A2 => n11152, Z => n7714);
   U16528 : XOR2_X1 port map( A1 => n698, A2 => n14215, Z => n18119);
   U16531 : INV_X1 port map( I => n15894, ZN => n16338);
   U16532 : XOR2_X1 port map( A1 => n22829, A2 => n21313, Z => n7723);
   U16534 : XOR2_X1 port map( A1 => n7726, A2 => n7727, Z => n7725);
   U16537 : NOR2_X1 port map( A1 => n14975, A2 => n20294, ZN => n7731);
   U16539 : NOR2_X1 port map( A1 => n7735, A2 => n14858, ZN => n7835);
   U16540 : NAND2_X1 port map( A1 => n26147, A2 => n7735, ZN => n11828);
   U16543 : INV_X1 port map( I => Plaintext(147), ZN => n7748);
   U16545 : XOR2_X1 port map( A1 => n7751, A2 => n18125, Z => n12854);
   U16546 : AND2_X1 port map( A1 => n7756, A2 => n16705, Z => n7754);
   U16547 : XOR2_X1 port map( A1 => n24000, A2 => n27848, Z => n7816);
   U16549 : OR2_X1 port map( A1 => n7370, A2 => n26615, Z => n7757);
   U16553 : XOR2_X1 port map( A1 => n8663, A2 => n7760, Z => n18452);
   U16554 : XOR2_X1 port map( A1 => n16869, A2 => n16870, Z => n7762);
   U16555 : XOR2_X1 port map( A1 => n7764, A2 => n21085, Z => n17934);
   U16556 : XOR2_X1 port map( A1 => n15237, A2 => n7764, Z => n14996);
   U16557 : XOR2_X1 port map( A1 => n7764, A2 => n14007, Z => n10947);
   U16559 : XOR2_X1 port map( A1 => n13007, A2 => n642, Z => n15362);
   U16562 : INV_X2 port map( I => n16065, ZN => n16316);
   U16564 : XOR2_X1 port map( A1 => n7776, A2 => n14650, Z => n19198);
   U16565 : XOR2_X1 port map( A1 => n19328, A2 => n7776, Z => n14105);
   U16568 : INV_X1 port map( I => n7784, ZN => n7780);
   U16572 : XOR2_X1 port map( A1 => n7803, A2 => n18235, Z => n13647);
   U16573 : XOR2_X1 port map( A1 => n7804, A2 => n27348, Z => n7803);
   U16577 : XOR2_X1 port map( A1 => n16939, A2 => n7816, Z => n7815);
   U16578 : XOR2_X1 port map( A1 => n7824, A2 => n12122, Z => n10876);
   U16579 : XOR2_X1 port map( A1 => n7824, A2 => n13133, Z => n13132);
   U16583 : NOR2_X1 port map( A1 => n11868, A2 => n27468, ZN => n7836);
   U16584 : XOR2_X1 port map( A1 => n7837, A2 => n20871, Z => Ciphertext(48));
   U16587 : XOR2_X1 port map( A1 => n18115, A2 => n7844, Z => n7843);
   U16588 : XOR2_X1 port map( A1 => n14026, A2 => n18352, Z => n7844);
   U16592 : NAND2_X1 port map( A1 => n8512, A2 => n8722, ZN => n7850);
   U16593 : INV_X2 port map( I => n7852, ZN => n15425);
   U16595 : XOR2_X1 port map( A1 => n7598, A2 => n21594, Z => n10688);
   U16596 : XOR2_X1 port map( A1 => n7858, A2 => n7857, Z => n7856);
   U16597 : XOR2_X1 port map( A1 => n14753, A2 => n25358, Z => n7858);
   U16599 : OR2_X1 port map( A1 => n11733, A2 => n28231, Z => n7864);
   U16605 : NAND2_X2 port map( A1 => n7873, A2 => n10163, ZN => n15057);
   U16606 : XOR2_X1 port map( A1 => n7875, A2 => n1190, Z => n7874);
   U16607 : INV_X1 port map( I => n16120, ZN => n13256);
   U16610 : XOR2_X1 port map( A1 => n25946, A2 => n1301, Z => n7883);
   U16611 : XOR2_X1 port map( A1 => n20577, A2 => n20429, Z => n7886);
   U16612 : XOR2_X1 port map( A1 => n5224, A2 => n1295, Z => n7887);
   U16614 : NAND2_X1 port map( A1 => n7890, A2 => n13769, ZN => n11850);
   U16615 : XOR2_X1 port map( A1 => n7902, A2 => n8524, Z => n7903);
   U16616 : INV_X2 port map( I => n7903, ZN => n10537);
   U16621 : NAND2_X1 port map( A1 => n3223, A2 => n22786, ZN => n10818);
   U16624 : NOR2_X1 port map( A1 => n17323, A2 => n7912, ZN => n17265);
   U16625 : NOR2_X1 port map( A1 => n20801, A2 => n27375, ZN => n13365);
   U16629 : NAND3_X2 port map( A1 => n14865, A2 => n16152, A3 => n14864, ZN => 
                           n16826);
   U16630 : XOR2_X1 port map( A1 => n16890, A2 => n12293, Z => n7916);
   U16632 : AOI21_X1 port map( A1 => n16213, A2 => n1266, B => n27240, ZN => 
                           n16214);
   U16635 : XOR2_X1 port map( A1 => n19289, A2 => n9926, Z => n7922);
   U16637 : XOR2_X1 port map( A1 => n19460, A2 => n9925, Z => n7923);
   U16643 : OAI21_X1 port map( A1 => n10851, A2 => n7944, B => n12508, ZN => 
                           n7945);
   U16644 : XOR2_X1 port map( A1 => n7949, A2 => n7947, Z => n7950);
   U16646 : INV_X2 port map( I => n7950, ZN => n14944);
   U16648 : XOR2_X1 port map( A1 => n4076, A2 => n20652, Z => n15683);
   U16658 : NAND2_X1 port map( A1 => n7980, A2 => n6999, ZN => n18905);
   U16659 : NAND2_X1 port map( A1 => n13347, A2 => n7980, ZN => n13346);
   U16662 : NOR2_X1 port map( A1 => n845, A2 => n26422, ZN => n7999);
   U16666 : XOR2_X1 port map( A1 => n9274, A2 => n13860, Z => n8002);
   U16669 : INV_X2 port map( I => n8011, ZN => n19850);
   U16670 : XOR2_X1 port map( A1 => n8018, A2 => n8019, Z => n10220);
   U16671 : XOR2_X1 port map( A1 => n17031, A2 => n10737, Z => n8016);
   U16672 : XOR2_X1 port map( A1 => n17124, A2 => n10195, Z => n8017);
   U16673 : XOR2_X1 port map( A1 => n16907, A2 => n16807, Z => n8019);
   U16676 : XOR2_X1 port map( A1 => n15537, A2 => n22784, Z => n8024);
   U16678 : NAND2_X1 port map( A1 => n14303, A2 => n8031, ZN => n15862);
   U16686 : NOR2_X1 port map( A1 => n20901, A2 => n28552, ZN => n20900);
   U16687 : INV_X2 port map( I => n8051, ZN => n10554);
   U16689 : INV_X2 port map( I => n8064, ZN => n11992);
   U16690 : XOR2_X1 port map( A1 => n9842, A2 => n9841, Z => n8064);
   U16698 : XOR2_X1 port map( A1 => n16778, A2 => n12523, Z => n8080);
   U16700 : XOR2_X1 port map( A1 => n8089, A2 => n16906, Z => n12555);
   U16701 : XOR2_X1 port map( A1 => n8089, A2 => n11972, Z => n9541);
   U16706 : XOR2_X1 port map( A1 => n11999, A2 => n13648, Z => n8112);
   U16713 : NOR2_X2 port map( A1 => n15677, A2 => n11242, ZN => n13371);
   U16715 : NAND2_X1 port map( A1 => n12221, A2 => n8254, ZN => n8123);
   U16717 : NAND2_X1 port map( A1 => n8126, A2 => n18570, ZN => n18499);
   U16725 : XOR2_X1 port map( A1 => n8140, A2 => n21247, Z => n8139);
   U16727 : XOR2_X1 port map( A1 => n10516, A2 => n17130, Z => n8143);
   U16728 : XOR2_X1 port map( A1 => n20546, A2 => n20544, Z => n8149);
   U16735 : NOR2_X1 port map( A1 => n9661, A2 => n22865, ZN => n9948);
   U16736 : INV_X2 port map( I => n8793, ZN => n8165);
   U16739 : XOR2_X1 port map( A1 => n21311, A2 => n21216, Z => n20388);
   U16750 : XOR2_X1 port map( A1 => n19383, A2 => n8195, Z => n8194);
   U16754 : XOR2_X1 port map( A1 => n18347, A2 => n8201, Z => n8200);
   U16755 : XOR2_X1 port map( A1 => n18290, A2 => n14492, Z => n8201);
   U16756 : XOR2_X1 port map( A1 => n18208, A2 => n8203, Z => n8202);
   U16759 : AOI22_X2 port map( A1 => n8211, A2 => n15579, B1 => n9393, B2 => 
                           n16229, ZN => n10393);
   U16760 : XOR2_X1 port map( A1 => n8216, A2 => n13155, Z => n13154);
   U16766 : XOR2_X1 port map( A1 => n8274, A2 => n17015, Z => n16763);
   U16767 : XOR2_X1 port map( A1 => n7302, A2 => n922, Z => n8242);
   U16770 : NAND2_X1 port map( A1 => n996, A2 => n14271, ZN => n10618);
   U16776 : NOR2_X1 port map( A1 => n8262, A2 => n23231, ZN => n12334);
   U16782 : NOR2_X1 port map( A1 => n9175, A2 => n11756, ZN => n8267);
   U16784 : NOR2_X2 port map( A1 => n10376, A2 => n8272, ZN => n8271);
   U16785 : XOR2_X1 port map( A1 => n8274, A2 => n20873, Z => n16720);
   U16787 : NAND2_X2 port map( A1 => n11042, A2 => n12822, ZN => n8274);
   U16789 : XOR2_X1 port map( A1 => n8293, A2 => n20771, Z => n20514);
   U16792 : AND3_X1 port map( A1 => n1257, A2 => n15701, A3 => n9759, Z => 
                           n9059);
   U16793 : NAND2_X1 port map( A1 => n17352, A2 => n17479, ZN => n10416);
   U16797 : XOR2_X1 port map( A1 => n8309, A2 => n10684, Z => n8308);
   U16800 : NAND2_X1 port map( A1 => n20752, A2 => n8311, ZN => n20753);
   U16802 : NAND2_X1 port map( A1 => n7910, A2 => n16005, ZN => n15210);
   U16804 : XOR2_X1 port map( A1 => n9597, A2 => n15651, Z => n8316);
   U16806 : XOR2_X1 port map( A1 => n20772, A2 => n20394, Z => n8318);
   U16813 : NAND2_X2 port map( A1 => n8346, A2 => n8345, ZN => n8344);
   U16814 : XOR2_X1 port map( A1 => n22839, A2 => n1281, Z => n8329);
   U16815 : INV_X1 port map( I => n10378, ZN => n8332);
   U16822 : XOR2_X1 port map( A1 => n8807, A2 => n8342, Z => n8341);
   U16823 : XOR2_X1 port map( A1 => n14421, A2 => n1317, Z => n8342);
   U16825 : NAND2_X1 port map( A1 => n12809, A2 => n25314, ZN => n8351);
   U16828 : NOR2_X1 port map( A1 => n8357, A2 => n18493, ZN => n8781);
   U16831 : AOI21_X2 port map( A1 => n19675, A2 => n8358, B => n15117, ZN => 
                           n20156);
   U16834 : OR2_X1 port map( A1 => n17335, A2 => n17563, Z => n8367);
   U16835 : INV_X2 port map( I => n8370, ZN => n10666);
   U16837 : NOR2_X1 port map( A1 => n8373, A2 => n9314, ZN => n16593);
   U16838 : NOR2_X1 port map( A1 => n27381, A2 => n8373, ZN => n16594);
   U16839 : MUX2_X1 port map( I0 => n8373, I1 => n6843, S => n9314, Z => n16420
                           );
   U16842 : XOR2_X1 port map( A1 => n8378, A2 => n14587, Z => n16905);
   U16843 : INV_X1 port map( I => n15969, ZN => n15967);
   U16844 : XOR2_X1 port map( A1 => Plaintext(6), A2 => Key(6), Z => n13418);
   U16846 : INV_X1 port map( I => n19652, ZN => n8390);
   U16847 : NOR2_X1 port map( A1 => n1519, A2 => n16516, ZN => n16375);
   U16852 : OAI22_X1 port map( A1 => n8925, A2 => n8398, B1 => n1269, B2 => 
                           n13677, ZN => n15978);
   U16853 : OAI21_X1 port map( A1 => n15976, A2 => n8398, B => n15959, ZN => 
                           n15962);
   U16855 : XOR2_X1 port map( A1 => n5740, A2 => n21707, Z => n19502);
   U16856 : XOR2_X1 port map( A1 => n5740, A2 => n13678, Z => n12635);
   U16857 : INV_X4 port map( I => n14211, ZN => n18101);
   U16858 : NAND2_X1 port map( A1 => n13983, A2 => n994, ZN => n8401);
   U16859 : XOR2_X1 port map( A1 => Plaintext(149), A2 => Key(149), Z => n8408)
                           ;
   U16862 : NAND3_X2 port map( A1 => n10850, A2 => n17933, A3 => n10849, ZN => 
                           n18359);
   U16863 : XOR2_X1 port map( A1 => n9125, A2 => n8405, Z => n9058);
   U16865 : XOR2_X1 port map( A1 => n20402, A2 => n14589, Z => n8405);
   U16868 : XOR2_X1 port map( A1 => Plaintext(146), A2 => Key(146), Z => n16104
                           );
   U16869 : XOR2_X1 port map( A1 => n8413, A2 => n10934, Z => n10933);
   U16872 : XOR2_X1 port map( A1 => n13514, A2 => n9833, Z => n8422);
   U16876 : XOR2_X1 port map( A1 => n19526, A2 => n10400, Z => n8429);
   U16877 : INV_X2 port map( I => n8430, ZN => n14126);
   U16878 : XOR2_X1 port map( A1 => n18171, A2 => n920, Z => n8431);
   U16879 : OR2_X1 port map( A1 => n8651, A2 => n18685, Z => n8433);
   U16883 : XOR2_X1 port map( A1 => n8438, A2 => n981, Z => n15754);
   U16884 : INV_X2 port map( I => n8439, ZN => n19499);
   U16885 : XOR2_X1 port map( A1 => n8441, A2 => n10766, Z => n8440);
   U16889 : XOR2_X1 port map( A1 => n8451, A2 => n18279, Z => n8450);
   U16890 : XOR2_X1 port map( A1 => n28287, A2 => n20919, Z => n8451);
   U16893 : AOI21_X2 port map( A1 => n8470, A2 => n7274, B => n8469, ZN => 
                           n20654);
   U16894 : NOR3_X2 port map( A1 => n8479, A2 => n8478, A3 => n8477, ZN => 
                           n21254);
   U16895 : XOR2_X1 port map( A1 => n9952, A2 => n9159, Z => n8484);
   U16898 : NOR2_X2 port map( A1 => n9164, A2 => n8501, ZN => n11364);
   U16900 : XOR2_X1 port map( A1 => n5698, A2 => n19285, Z => n19485);
   U16903 : XOR2_X1 port map( A1 => n19486, A2 => n610, Z => n8504);
   U16904 : XOR2_X1 port map( A1 => n10056, A2 => n21077, Z => n8505);
   U16905 : NOR2_X1 port map( A1 => n18927, A2 => n19160, ZN => n8516);
   U16910 : XOR2_X1 port map( A1 => n580, A2 => n11970, Z => n8524);
   U16911 : NOR2_X1 port map( A1 => n1550, A2 => n10537, ZN => n13612);
   U16913 : NAND2_X2 port map( A1 => n9180, A2 => n8528, ZN => n17868);
   U16914 : INV_X2 port map( I => n8529, ZN => n19870);
   U16922 : INV_X2 port map( I => n8545, ZN => n10978);
   U16924 : XOR2_X1 port map( A1 => n17096, A2 => n8551, Z => n8548);
   U16926 : XOR2_X1 port map( A1 => n17139, A2 => n21090, Z => n8551);
   U16927 : NAND3_X1 port map( A1 => n20659, A2 => n20664, A3 => n8559, ZN => 
                           n20660);
   U16929 : INV_X2 port map( I => n15619, ZN => n19720);
   U16931 : XOR2_X1 port map( A1 => n8570, A2 => n8569, Z => n8568);
   U16932 : XOR2_X1 port map( A1 => n2265, A2 => n21262, Z => n8569);
   U16933 : XOR2_X1 port map( A1 => n13101, A2 => n16868, Z => n8570);
   U16942 : XOR2_X1 port map( A1 => n7065, A2 => n21454, Z => n8582);
   U16945 : NAND2_X1 port map( A1 => n8586, A2 => n8585, ZN => n8584);
   U16948 : XOR2_X1 port map( A1 => n8596, A2 => n8595, Z => n10401);
   U16949 : XOR2_X1 port map( A1 => n21366, A2 => n8597, Z => n8596);
   U16950 : XOR2_X1 port map( A1 => n10529, A2 => n11261, Z => n8600);
   U16952 : XOR2_X1 port map( A1 => n8608, A2 => n23731, Z => n11887);
   U16953 : INV_X1 port map( I => n8610, ZN => n9305);
   U16954 : NOR2_X1 port map( A1 => n7299, A2 => n24538, ZN => n12294);
   U16955 : NOR2_X1 port map( A1 => n7299, A2 => n13424, ZN => n11977);
   U16956 : NAND2_X1 port map( A1 => n21457, A2 => n7299, ZN => n21458);
   U16957 : NOR2_X1 port map( A1 => n12074, A2 => n12073, ZN => n12072);
   U16958 : INV_X2 port map( I => n19932, ZN => n19750);
   U16965 : XOR2_X1 port map( A1 => n8636, A2 => n21613, Z => n19175);
   U16966 : INV_X2 port map( I => n8637, ZN => n10985);
   U16967 : OAI22_X2 port map( A1 => n8641, A2 => n8639, B1 => n8638, B2 => 
                           n28160, ZN => n19160);
   U16968 : NOR2_X1 port map( A1 => n8640, A2 => n18776, ZN => n8639);
   U16970 : NAND2_X1 port map( A1 => n8645, A2 => n15041, ZN => n18820);
   U16972 : XOR2_X1 port map( A1 => Key(88), A2 => Plaintext(88), Z => n8648);
   U16974 : NAND3_X1 port map( A1 => n1059, A2 => n16027, A3 => n8647, ZN => 
                           n15847);
   U16976 : XOR2_X1 port map( A1 => n634, A2 => n8650, Z => n8649);
   U16979 : INV_X2 port map( I => n8654, ZN => n8717);
   U16980 : XOR2_X1 port map( A1 => n27357, A2 => n21557, Z => n14266);
   U16983 : MUX2_X1 port map( I0 => n15965, I1 => n16338, S => n16339, Z => 
                           n8665);
   U16984 : XOR2_X1 port map( A1 => n27360, A2 => n21164, Z => n8669);
   U16985 : XOR2_X1 port map( A1 => n25313, A2 => n10339, Z => n8670);
   U16991 : XOR2_X1 port map( A1 => n18323, A2 => n15057, Z => n8681);
   U16992 : XOR2_X1 port map( A1 => n18322, A2 => n18325, Z => n8682);
   U16995 : OAI21_X2 port map( A1 => n16312, A2 => n8687, B => n8686, ZN => 
                           n16567);
   U16996 : XOR2_X1 port map( A1 => n8691, A2 => n8688, Z => n18418);
   U16997 : XOR2_X1 port map( A1 => n8690, A2 => n8689, Z => n8688);
   U16998 : XOR2_X1 port map( A1 => n9722, A2 => n25371, Z => n8690);
   U16999 : XOR2_X1 port map( A1 => n18257, A2 => n18322, Z => n8691);
   U17000 : OR2_X1 port map( A1 => n1166, A2 => n18908, Z => n8694);
   U17001 : INV_X1 port map( I => n8696, ZN => n16105);
   U17003 : XOR2_X1 port map( A1 => n21247, A2 => n20423, Z => n20509);
   U17004 : NAND2_X2 port map( A1 => n8699, A2 => n8698, ZN => n21247);
   U17006 : INV_X1 port map( I => n18556, ZN => n8703);
   U17007 : XOR2_X1 port map( A1 => n11708, A2 => n1277, Z => n19142);
   U17008 : XOR2_X1 port map( A1 => n63, A2 => n19507, Z => n19183);
   U17012 : NAND2_X2 port map( A1 => n1127, A2 => n8717, ZN => n12982);
   U17024 : NAND2_X1 port map( A1 => n8741, A2 => n21484, ZN => n21460);
   U17032 : INV_X1 port map( I => n8760, ZN => n20846);
   U17034 : OAI21_X1 port map( A1 => n8760, A2 => n28213, B => n20843, ZN => 
                           n20844);
   U17035 : NOR2_X2 port map( A1 => n8763, A2 => n8762, ZN => n16572);
   U17041 : XOR2_X1 port map( A1 => n8776, A2 => n12481, Z => n16762);
   U17044 : NAND2_X2 port map( A1 => n17699, A2 => n17698, ZN => n18021);
   U17048 : NOR2_X1 port map( A1 => n8798, A2 => n16455, ZN => n8797);
   U17051 : INV_X2 port map( I => n8805, ZN => n21723);
   U17056 : XOR2_X1 port map( A1 => n8819, A2 => n16943, Z => n8900);
   U17058 : XOR2_X1 port map( A1 => n19492, A2 => n10214, Z => n8822);
   U17059 : XOR2_X1 port map( A1 => n10671, A2 => n558, Z => n8825);
   U17064 : XOR2_X1 port map( A1 => n8832, A2 => n26473, Z => Ciphertext(185));
   U17065 : OAI21_X1 port map( A1 => n8853, A2 => n8854, B => n8851, ZN => 
                           n12021);
   U17066 : XNOR2_X1 port map( A1 => n8857, A2 => n8858, ZN => n8855);
   U17068 : XOR2_X1 port map( A1 => n12601, A2 => n18089, Z => n8858);
   U17069 : OR2_X1 port map( A1 => n10389, A2 => n1284, Z => n8860);
   U17070 : XOR2_X1 port map( A1 => n14753, A2 => n20650, Z => n8861);
   U17077 : NOR2_X1 port map( A1 => n4122, A2 => n24576, ZN => n8875);
   U17079 : XOR2_X1 port map( A1 => n3, A2 => n21411, Z => n11867);
   U17083 : OAI21_X1 port map( A1 => n21208, A2 => n21324, B => n9131, ZN => 
                           n12097);
   U17087 : XOR2_X1 port map( A1 => n16990, A2 => n8904, Z => n8902);
   U17088 : NAND2_X1 port map( A1 => n15000, A2 => n14128, ZN => n8921);
   U17089 : NOR3_X1 port map( A1 => n26252, A2 => n28151, A3 => n22224, ZN => 
                           n8929);
   U17093 : INV_X1 port map( I => n13247, ZN => n13623);
   U17096 : INV_X2 port map( I => n8948, ZN => n21027);
   U17099 : XOR2_X1 port map( A1 => n8954, A2 => n8955, Z => n8953);
   U17104 : XOR2_X1 port map( A1 => Plaintext(60), A2 => Key(60), Z => n10573);
   U17110 : XOR2_X1 port map( A1 => n4585, A2 => n8965, Z => n8964);
   U17111 : XOR2_X1 port map( A1 => n1912, A2 => n14560, Z => n8965);
   U17113 : NAND2_X2 port map( A1 => n11533, A2 => n11532, ZN => n13530);
   U17114 : XOR2_X1 port map( A1 => n5026, A2 => n556, Z => n8984);
   U17120 : XOR2_X1 port map( A1 => n8992, A2 => n8993, Z => n8991);
   U17121 : XOR2_X1 port map( A1 => n19489, A2 => n14489, Z => n8993);
   U17125 : XOR2_X1 port map( A1 => n11339, A2 => n11867, Z => n9006);
   U17126 : XOR2_X1 port map( A1 => n617, A2 => n9008, Z => n9007);
   U17127 : XOR2_X1 port map( A1 => n16916, A2 => n26053, Z => n9008);
   U17128 : XOR2_X1 port map( A1 => n9013, A2 => n9016, Z => n9779);
   U17132 : XOR2_X1 port map( A1 => n9017, A2 => n19193, Z => n9016);
   U17137 : XOR2_X1 port map( A1 => n9025, A2 => n9024, Z => n18456);
   U17144 : XOR2_X1 port map( A1 => n19523, A2 => n9036, Z => n9035);
   U17145 : XOR2_X1 port map( A1 => n5653, A2 => n1290, Z => n9036);
   U17146 : XOR2_X1 port map( A1 => n19250, A2 => n19522, Z => n9038);
   U17152 : NAND2_X1 port map( A1 => n11214, A2 => n7364, ZN => n20300);
   U17157 : NOR2_X1 port map( A1 => n9047, A2 => n12061, ZN => n21678);
   U17158 : NAND2_X1 port map( A1 => n9047, A2 => n12061, ZN => n21684);
   U17160 : NAND2_X1 port map( A1 => n2777, A2 => n9047, ZN => n21675);
   U17162 : XOR2_X1 port map( A1 => n20761, A2 => n27391, Z => n13504);
   U17166 : XOR2_X1 port map( A1 => n19527, A2 => n19500, Z => n19394);
   U17167 : OAI21_X2 port map( A1 => n12627, A2 => n9060, B => n12138, ZN => 
                           n19500);
   U17170 : XOR2_X1 port map( A1 => n9316, A2 => n7302, Z => n9071);
   U17171 : INV_X1 port map( I => n9072, ZN => n16811);
   U17172 : NAND3_X2 port map( A1 => n9386, A2 => n10510, A3 => n10508, ZN => 
                           n18360);
   U17173 : XOR2_X1 port map( A1 => n13807, A2 => n9081, Z => n9080);
   U17174 : XOR2_X1 port map( A1 => n24363, A2 => n18072, Z => n13807);
   U17178 : XOR2_X1 port map( A1 => n19516, A2 => n1289, Z => n9096);
   U17180 : AOI21_X1 port map( A1 => n11766, A2 => n7944, B => n11765, ZN => 
                           n11764);
   U17181 : NAND2_X1 port map( A1 => n20165, A2 => n4858, ZN => n11256);
   U17185 : NAND2_X2 port map( A1 => n12389, A2 => n14689, ZN => n20269);
   U17188 : MUX2_X1 port map( I0 => n9472, I1 => n24336, S => n28224, Z => 
                           n9121);
   U17189 : XOR2_X1 port map( A1 => n20576, A2 => n20353, Z => n9124);
   U17190 : XOR2_X1 port map( A1 => n9670, A2 => n11866, Z => n9130);
   U17191 : XOR2_X1 port map( A1 => n9414, A2 => n20877, Z => n9137);
   U17194 : NAND3_X1 port map( A1 => n16409, A2 => n16648, A3 => n9139, ZN => 
                           n15382);
   U17196 : XOR2_X1 port map( A1 => n15001, A2 => n18010, Z => n9145);
   U17198 : INV_X2 port map( I => n9147, ZN => n19883);
   U17200 : XOR2_X1 port map( A1 => n19281, A2 => n18831, Z => n9148);
   U17201 : XOR2_X1 port map( A1 => n9774, A2 => n26038, Z => n9154);
   U17209 : XNOR2_X1 port map( A1 => Plaintext(159), A2 => Key(159), ZN => 
                           n9173);
   U17210 : XOR2_X1 port map( A1 => Plaintext(161), A2 => Key(161), Z => n9218)
                           ;
   U17217 : XOR2_X1 port map( A1 => n28293, A2 => n25337, Z => n15293);
   U17218 : NAND2_X1 port map( A1 => n25389, A2 => n10810, ZN => n9191);
   U17220 : XOR2_X1 port map( A1 => n9063, A2 => n20369, Z => n9197);
   U17222 : INV_X2 port map( I => n15225, ZN => n21507);
   U17225 : XOR2_X1 port map( A1 => n18199, A2 => n9201, Z => n10711);
   U17226 : XOR2_X1 port map( A1 => n7951, A2 => n6562, Z => n9201);
   U17229 : OAI21_X2 port map( A1 => n13550, A2 => n13549, B => n18956, ZN => 
                           n13046);
   U17230 : NAND2_X2 port map( A1 => n11361, A2 => n19776, ZN => n20490);
   U17236 : XOR2_X1 port map( A1 => n9229, A2 => n12713, Z => Ciphertext(80));
   U17237 : XOR2_X1 port map( A1 => n15743, A2 => n17765, Z => n9230);
   U17239 : OAI21_X1 port map( A1 => n16107, A2 => n22801, B => n9432, ZN => 
                           n9431);
   U17241 : XOR2_X1 port map( A1 => n17784, A2 => n9242, Z => n9241);
   U17243 : XOR2_X1 port map( A1 => n9244, A2 => n17008, Z => n17012);
   U17248 : XOR2_X1 port map( A1 => n9257, A2 => n9254, Z => n19901);
   U17249 : XOR2_X1 port map( A1 => n9256, A2 => n9255, Z => n9254);
   U17250 : XOR2_X1 port map( A1 => n19406, A2 => n14491, Z => n9255);
   U17257 : XOR2_X1 port map( A1 => n9274, A2 => n17627, Z => n17628);
   U17258 : XOR2_X1 port map( A1 => n7130, A2 => n10544, Z => n9279);
   U17265 : XOR2_X1 port map( A1 => n11493, A2 => n19384, Z => n9284);
   U17270 : NOR3_X1 port map( A1 => n9946, A2 => n24524, A3 => n27647, ZN => 
                           n9743);
   U17275 : NAND2_X1 port map( A1 => n9323, A2 => n18621, ZN => n12306);
   U17276 : XOR2_X1 port map( A1 => n19331, A2 => n9325, Z => n9742);
   U17277 : XOR2_X1 port map( A1 => n19333, A2 => n8777, Z => n9325);
   U17281 : NAND2_X1 port map( A1 => n26639, A2 => n27433, ZN => n18402);
   U17283 : XOR2_X1 port map( A1 => Plaintext(37), A2 => Key(37), Z => n11835);
   U17284 : XOR2_X1 port map( A1 => n19536, A2 => n20906, Z => n9335);
   U17285 : OR2_X1 port map( A1 => n23408, A2 => n7908, Z => n9337);
   U17286 : XOR2_X1 port map( A1 => n9338, A2 => n19222, Z => n19223);
   U17294 : AND2_X1 port map( A1 => n9561, A2 => n19820, Z => n9367);
   U17298 : XOR2_X1 port map( A1 => n23352, A2 => n13524, Z => n16740);
   U17299 : XOR2_X1 port map( A1 => n17114, A2 => n27705, Z => n16770);
   U17300 : XOR2_X1 port map( A1 => n17069, A2 => n27705, Z => n15594);
   U17303 : XOR2_X1 port map( A1 => n19401, A2 => n9384, Z => n9383);
   U17304 : XOR2_X1 port map( A1 => n8912, A2 => n5653, Z => n9384);
   U17305 : INV_X1 port map( I => n7355, ZN => n21517);
   U17306 : XOR2_X1 port map( A1 => n28233, A2 => n7355, Z => n17746);
   U17307 : AOI21_X2 port map( A1 => n9394, A2 => n16270, B => n10321, ZN => 
                           n16517);
   U17309 : XOR2_X1 port map( A1 => n27858, A2 => n9397, Z => n21241);
   U17311 : INV_X2 port map( I => n9411, ZN => n18445);
   U17313 : NAND3_X1 port map( A1 => n20312, A2 => n9417, A3 => n10167, ZN => 
                           n13551);
   U17314 : INV_X1 port map( I => Plaintext(157), ZN => n9420);
   U17315 : XOR2_X1 port map( A1 => n9420, A2 => Key(157), Z => n9557);
   U17318 : NAND2_X2 port map( A1 => n10257, A2 => n10258, ZN => n17895);
   U17324 : XOR2_X1 port map( A1 => n15711, A2 => n20320, Z => n9451);
   U17326 : NAND3_X1 port map( A1 => n21739, A2 => n14350, A3 => n9458, ZN => 
                           n14060);
   U17328 : XOR2_X1 port map( A1 => n36, A2 => n918, Z => n9463);
   U17335 : INV_X2 port map( I => n4618, ZN => n9477);
   U17340 : XOR2_X1 port map( A1 => n9489, A2 => n18018, Z => n10614);
   U17341 : XOR2_X1 port map( A1 => n18016, A2 => n9490, Z => n9489);
   U17343 : NOR2_X1 port map( A1 => n7039, A2 => n9494, ZN => n14901);
   U17345 : XOR2_X1 port map( A1 => n18171, A2 => n9499, Z => n9498);
   U17347 : XOR2_X1 port map( A1 => n9505, A2 => n548, Z => n9504);
   U17348 : XOR2_X1 port map( A1 => n19509, A2 => n19508, Z => n15213);
   U17351 : XOR2_X1 port map( A1 => n9513, A2 => n9511, Z => n9510);
   U17352 : XOR2_X1 port map( A1 => n22792, A2 => n9512, Z => n9511);
   U17353 : XOR2_X1 port map( A1 => n9531, A2 => n9529, Z => n9535);
   U17354 : XOR2_X1 port map( A1 => n17124, A2 => n9530, Z => n9529);
   U17355 : XOR2_X1 port map( A1 => n9532, A2 => n17126, Z => n9531);
   U17356 : XOR2_X1 port map( A1 => n9536, A2 => n14999, Z => n9532);
   U17357 : INV_X2 port map( I => n9535, ZN => n10559);
   U17360 : XOR2_X1 port map( A1 => n10378, A2 => n21216, Z => n9543);
   U17371 : INV_X2 port map( I => n9557, ZN => n16244);
   U17376 : XOR2_X1 port map( A1 => n16822, A2 => n26566, Z => n9574);
   U17377 : XOR2_X1 port map( A1 => n9576, A2 => n12916, Z => Ciphertext(147));
   U17378 : XOR2_X1 port map( A1 => n9580, A2 => n10063, Z => n10062);
   U17379 : XOR2_X1 port map( A1 => n18305, A2 => n9581, Z => n9580);
   U17380 : XOR2_X1 port map( A1 => n761, A2 => n24258, Z => n9581);
   U17381 : XOR2_X1 port map( A1 => Key(47), A2 => Plaintext(47), Z => n11722);
   U17383 : XOR2_X1 port map( A1 => n9656, A2 => n21839, Z => n9585);
   U17387 : XOR2_X1 port map( A1 => n9791, A2 => n9345, Z => n19469);
   U17388 : XOR2_X1 port map( A1 => Key(120), A2 => n9596, Z => n14311);
   U17389 : INV_X1 port map( I => Plaintext(120), ZN => n9596);
   U17391 : NOR2_X1 port map( A1 => n1223, A2 => n10577, ZN => n9609);
   U17393 : XOR2_X1 port map( A1 => n6123, A2 => n14633, Z => n9613);
   U17394 : XOR2_X1 port map( A1 => n10641, A2 => n13332, Z => n9620);
   U17400 : XOR2_X1 port map( A1 => n136, A2 => n21554, Z => n9638);
   U17401 : XOR2_X1 port map( A1 => n13855, A2 => n27364, Z => n9640);
   U17402 : INV_X2 port map( I => n9641, ZN => n18645);
   U17407 : XOR2_X1 port map( A1 => n27245, A2 => n9663, Z => n9662);
   U17409 : XOR2_X1 port map( A1 => n9063, A2 => n19285, Z => n12261);
   U17410 : XOR2_X1 port map( A1 => n9063, A2 => n21449, Z => n9771);
   U17414 : XOR2_X1 port map( A1 => n28483, A2 => n21742, Z => n9680);
   U17415 : XOR2_X1 port map( A1 => n13300, A2 => n10751, Z => n9682);
   U17418 : NOR2_X1 port map( A1 => n11968, A2 => n9691, ZN => n17931);
   U17421 : XOR2_X1 port map( A1 => n9708, A2 => n9710, Z => n9707);
   U17422 : XOR2_X1 port map( A1 => n19406, A2 => n9709, Z => n9708);
   U17423 : XOR2_X1 port map( A1 => n982, A2 => n13001, Z => n9710);
   U17424 : XOR2_X1 port map( A1 => n11990, A2 => n19242, Z => n9711);
   U17425 : XOR2_X1 port map( A1 => n12343, A2 => n9724, Z => n9723);
   U17426 : NAND2_X2 port map( A1 => n15136, A2 => n17988, ZN => n18088);
   U17428 : XOR2_X1 port map( A1 => Plaintext(151), A2 => Key(151), Z => n10064
                           );
   U17432 : XOR2_X1 port map( A1 => n9741, A2 => n9740, Z => n9739);
   U17433 : XOR2_X1 port map( A1 => n19201, A2 => n14492, Z => n9740);
   U17434 : XOR2_X1 port map( A1 => n14608, A2 => n19430, Z => n9741);
   U17436 : XOR2_X1 port map( A1 => n9750, A2 => n9747, Z => n9746);
   U17437 : XOR2_X1 port map( A1 => n18211, A2 => n9748, Z => n9747);
   U17438 : XOR2_X1 port map( A1 => n18209, A2 => n14489, Z => n9749);
   U17440 : INV_X2 port map( I => n15156, ZN => n14319);
   U17442 : NOR2_X1 port map( A1 => n5502, A2 => n9759, ZN => n9801);
   U17444 : NAND3_X1 port map( A1 => n18583, A2 => n7190, A3 => n18507, ZN => 
                           n18342);
   U17446 : NAND2_X1 port map( A1 => n1253, A2 => n905, ZN => n9764);
   U17449 : INV_X1 port map( I => n22741, ZN => n13513);
   U17450 : XOR2_X1 port map( A1 => n19248, A2 => n9771, Z => n11479);
   U17452 : XOR2_X1 port map( A1 => n9774, A2 => n20381, Z => n11655);
   U17454 : INV_X2 port map( I => n9779, ZN => n12502);
   U17455 : XOR2_X1 port map( A1 => n18087, A2 => n14995, Z => n9780);
   U17458 : AND2_X1 port map( A1 => n15981, A2 => n15924, Z => n9787);
   U17459 : XOR2_X1 port map( A1 => n3390, A2 => n15731, Z => n15730);
   U17460 : XOR2_X1 port map( A1 => n9791, A2 => n20908, Z => n19262);
   U17462 : NOR2_X1 port map( A1 => n9794, A2 => n15828, ZN => n9793);
   U17468 : XOR2_X1 port map( A1 => n9802, A2 => n7365, Z => n18030);
   U17481 : XOR2_X1 port map( A1 => n9846, A2 => n21643, Z => Ciphertext(166));
   U17483 : XOR2_X1 port map( A1 => n27858, A2 => n1061, Z => n9858);
   U17484 : XOR2_X1 port map( A1 => n20580, A2 => n13342, Z => n9859);
   U17486 : XOR2_X1 port map( A1 => n9862, A2 => n13787, Z => Ciphertext(84));
   U17487 : NAND4_X1 port map( A1 => n9866, A2 => n15479, A3 => n21057, A4 => 
                           n10687, ZN => n9868);
   U17495 : NAND2_X2 port map( A1 => n12024, A2 => n12019, ZN => n21711);
   U17499 : XOR2_X1 port map( A1 => n14608, A2 => n14432, Z => n9920);
   U17501 : INV_X2 port map( I => n9924, ZN => n19744);
   U17502 : XOR2_X1 port map( A1 => n19333, A2 => n27444, Z => n9925);
   U17503 : XOR2_X1 port map( A1 => n19562, A2 => n923, Z => n9926);
   U17504 : XOR2_X1 port map( A1 => n9928, A2 => n9927, Z => Ciphertext(180));
   U17505 : INV_X1 port map( I => n21703, ZN => n9927);
   U17508 : XOR2_X1 port map( A1 => n11643, A2 => n11010, Z => n9932);
   U17516 : XOR2_X1 port map( A1 => n7284, A2 => n10277, Z => n9964);
   U17518 : OAI21_X1 port map( A1 => n21664, A2 => n11263, B => n10984, ZN => 
                           n9972);
   U17519 : NAND2_X1 port map( A1 => n766, A2 => n10580, ZN => n9975);
   U17521 : XOR2_X1 port map( A1 => n3663, A2 => n20406, Z => n9983);
   U17525 : XOR2_X1 port map( A1 => n94, A2 => n9999, Z => n9998);
   U17528 : XOR2_X1 port map( A1 => Plaintext(176), A2 => Key(176), Z => n16228
                           );
   U17529 : XOR2_X1 port map( A1 => n27365, A2 => n19042, Z => n10004);
   U17530 : NAND3_X1 port map( A1 => n22570, A2 => n1256, A3 => n10597, ZN => 
                           n12336);
   U17531 : NAND2_X1 port map( A1 => n17403, A2 => n26198, ZN => n17405);
   U17532 : INV_X1 port map( I => n10217, ZN => n21221);
   U17534 : INV_X1 port map( I => n17422, ZN => n17530);
   U17539 : XOR2_X1 port map( A1 => n699, A2 => n1064, Z => n10122);
   U17540 : XOR2_X1 port map( A1 => n18175, A2 => n18138, Z => n18139);
   U17541 : NAND2_X1 port map( A1 => n10030, A2 => n13819, ZN => n13826);
   U17542 : INV_X2 port map( I => n10032, ZN => n11110);
   U17543 : XOR2_X1 port map( A1 => n10852, A2 => n596, Z => n10033);
   U17544 : AOI21_X1 port map( A1 => n14177, A2 => n16461, B => n3479, ZN => 
                           n10034);
   U17545 : XOR2_X1 port map( A1 => n22793, A2 => n19490, Z => n10944);
   U17546 : AND2_X1 port map( A1 => n10040, A2 => n10174, Z => n15498);
   U17550 : XOR2_X1 port map( A1 => n16785, A2 => n10048, Z => n10047);
   U17551 : XOR2_X1 port map( A1 => n13524, A2 => n1288, Z => n10048);
   U17553 : XOR2_X1 port map( A1 => n11261, A2 => n18215, Z => n10051);
   U17555 : XOR2_X1 port map( A1 => n5529, A2 => n21033, Z => n10053);
   U17561 : NAND2_X2 port map( A1 => n14615, A2 => n10066, ZN => n17952);
   U17562 : OAI21_X1 port map( A1 => n1224, A2 => n24406, B => n10067, ZN => 
                           n10066);
   U17563 : AOI21_X1 port map( A1 => n1224, A2 => n1036, B => n21785, ZN => 
                           n10067);
   U17566 : XOR2_X1 port map( A1 => n10071, A2 => n19196, Z => n10070);
   U17569 : NAND3_X2 port map( A1 => n11231, A2 => n11230, A3 => n20094, ZN => 
                           n20424);
   U17572 : INV_X2 port map( I => n19399, ZN => n19931);
   U17575 : XOR2_X1 port map( A1 => n23950, A2 => n18078, Z => n17779);
   U17576 : NAND2_X1 port map( A1 => n15981, A2 => n16136, ZN => n15928);
   U17581 : XOR2_X1 port map( A1 => n17069, A2 => n10123, Z => n12091);
   U17582 : XOR2_X1 port map( A1 => n16750, A2 => n10123, Z => n14428);
   U17584 : XOR2_X1 port map( A1 => Key(81), A2 => Plaintext(81), Z => n14607);
   U17585 : INV_X2 port map( I => n10144, ZN => n15490);
   U17587 : NAND2_X2 port map( A1 => n15499, A2 => n15500, ZN => n21659);
   U17588 : XOR2_X1 port map( A1 => n10146, A2 => n14457, Z => Ciphertext(173))
                           ;
   U17591 : NOR2_X2 port map( A1 => n21668, A2 => n21629, ZN => n12615);
   U17592 : INV_X2 port map( I => n15476, ZN => n21668);
   U17597 : XOR2_X1 port map( A1 => n14215, A2 => n20989, Z => n10179);
   U17602 : XOR2_X1 port map( A1 => n26848, A2 => n25840, Z => n15402);
   U17605 : XOR2_X1 port map( A1 => Plaintext(20), A2 => Key(20), Z => n10204);
   U17606 : INV_X2 port map( I => n10204, ZN => n16207);
   U17607 : NOR2_X1 port map( A1 => n10303, A2 => n16207, ZN => n15756);
   U17610 : XOR2_X1 port map( A1 => n12114, A2 => n12327, Z => n10213);
   U17611 : XOR2_X1 port map( A1 => n13357, A2 => n11275, Z => n10214);
   U17615 : XOR2_X1 port map( A1 => n10494, A2 => n14596, Z => n10234);
   U17616 : XOR2_X1 port map( A1 => n534, A2 => n10236, Z => n10431);
   U17617 : XOR2_X1 port map( A1 => n16792, A2 => n10237, Z => n10236);
   U17622 : OAI21_X2 port map( A1 => n10254, A2 => n10253, B => n12252, ZN => 
                           n12251);
   U17623 : INV_X2 port map( I => n10255, ZN => n19846);
   U17627 : AOI21_X1 port map( A1 => n21221, A2 => n10268, B => n12430, ZN => 
                           n21217);
   U17628 : XNOR2_X1 port map( A1 => Plaintext(139), A2 => Key(139), ZN => 
                           n10269);
   U17632 : OAI21_X1 port map( A1 => n20623, A2 => n25318, B => n22766, ZN => 
                           n10275);
   U17633 : INV_X1 port map( I => n20620, ZN => n10276);
   U17637 : XOR2_X1 port map( A1 => n668, A2 => n12515, Z => n11220);
   U17640 : XOR2_X1 port map( A1 => n10294, A2 => n20692, Z => n16834);
   U17641 : OR2_X1 port map( A1 => n10579, A2 => n7966, Z => n10297);
   U17643 : XNOR2_X1 port map( A1 => Plaintext(22), A2 => Key(22), ZN => n10303
                           );
   U17646 : XOR2_X1 port map( A1 => n10313, A2 => n10310, Z => n10638);
   U17647 : XOR2_X1 port map( A1 => n10312, A2 => n10311, Z => n10310);
   U17648 : INV_X1 port map( I => n12585, ZN => n10314);
   U17649 : NAND2_X1 port map( A1 => n780, A2 => n10315, ZN => n10316);
   U17651 : XOR2_X1 port map( A1 => n10318, A2 => n18857, Z => n10317);
   U17652 : XOR2_X1 port map( A1 => n22784, A2 => n20877, Z => n10320);
   U17655 : XOR2_X1 port map( A1 => n18113, A2 => n21733, Z => n10327);
   U17657 : XOR2_X1 port map( A1 => n20540, A2 => n20404, Z => n21438);
   U17659 : INV_X2 port map( I => n10332, ZN => n13424);
   U17660 : XOR2_X1 port map( A1 => n10335, A2 => n20321, Z => Ciphertext(97));
   U17663 : INV_X1 port map( I => n14558, ZN => n15798);
   U17667 : AOI21_X2 port map( A1 => n11356, A2 => n19934, B => n11355, ZN => 
                           n21190);
   U17668 : XOR2_X1 port map( A1 => n5351, A2 => n21602, Z => n13512);
   U17669 : XOR2_X1 port map( A1 => n10358, A2 => n21090, Z => n19308);
   U17671 : XOR2_X1 port map( A1 => n18327, A2 => n10365, Z => n10364);
   U17672 : XOR2_X1 port map( A1 => n15472, A2 => n21385, Z => n10369);
   U17673 : XOR2_X1 port map( A1 => n10370, A2 => n14593, Z => Ciphertext(129))
                           ;
   U17674 : XOR2_X1 port map( A1 => n21235, A2 => n25642, Z => n10373);
   U17675 : XOR2_X1 port map( A1 => n27408, A2 => n1286, Z => n10374);
   U17680 : XOR2_X1 port map( A1 => n18314, A2 => n14600, Z => n10382);
   U17681 : XOR2_X1 port map( A1 => n21438, A2 => n13590, Z => n10383);
   U17683 : XOR2_X1 port map( A1 => n19556, A2 => n19557, Z => n10390);
   U17686 : OAI21_X1 port map( A1 => n21891, A2 => n23096, B => n24334, ZN => 
                           n16596);
   U17687 : XOR2_X1 port map( A1 => n22749, A2 => n24528, Z => n10400);
   U17689 : XOR2_X1 port map( A1 => n10413, A2 => n10412, Z => n10499);
   U17690 : XOR2_X1 port map( A1 => n19389, A2 => n14741, Z => n10412);
   U17693 : NAND2_X1 port map( A1 => n18545, A2 => n27739, ZN => n18538);
   U17695 : XOR2_X1 port map( A1 => n3477, A2 => n23839, Z => n10441);
   U17696 : XOR2_X1 port map( A1 => n11074, A2 => n11014, Z => n10442);
   U17698 : XOR2_X1 port map( A1 => n1709, A2 => n11918, Z => n11917);
   U17699 : XOR2_X1 port map( A1 => n1709, A2 => n12481, Z => n11524);
   U17700 : XOR2_X1 port map( A1 => n1709, A2 => n13285, Z => n13284);
   U17705 : NAND3_X1 port map( A1 => n26031, A2 => n18666, A3 => n24297, ZN => 
                           n10455);
   U17707 : XOR2_X1 port map( A1 => n18249, A2 => n10456, Z => n18315);
   U17708 : XOR2_X1 port map( A1 => n11364, A2 => n10456, Z => n17827);
   U17712 : INV_X2 port map( I => n10465, ZN => n10591);
   U17713 : XOR2_X1 port map( A1 => n20549, A2 => n10467, Z => n10466);
   U17714 : XOR2_X1 port map( A1 => n7848, A2 => n20871, Z => n10467);
   U17715 : XOR2_X1 port map( A1 => n10475, A2 => n14610, Z => Ciphertext(38));
   U17718 : NOR2_X1 port map( A1 => n10050, A2 => n20799, ZN => n10478);
   U17719 : OAI21_X2 port map( A1 => n11637, A2 => n11636, B => n10479, ZN => 
                           n19090);
   U17720 : XOR2_X1 port map( A1 => n21299, A2 => n10481, Z => n14273);
   U17721 : INV_X1 port map( I => n20727, ZN => n10481);
   U17722 : NOR2_X2 port map( A1 => n10486, A2 => n15175, ZN => n11627);
   U17727 : XOR2_X1 port map( A1 => n19555, A2 => n19266, Z => n10495);
   U17728 : INV_X2 port map( I => n10497, ZN => n14528);
   U17737 : XNOR2_X1 port map( A1 => n10906, A2 => n11408, ZN => n10516);
   U17739 : OAI21_X1 port map( A1 => n19796, A2 => n8255, B => n26120, ZN => 
                           n10521);
   U17740 : NOR2_X1 port map( A1 => n13247, A2 => n14103, ZN => n12720);
   U17744 : XOR2_X1 port map( A1 => n10527, A2 => n10526, Z => n10525);
   U17745 : XOR2_X1 port map( A1 => n27145, A2 => n21709, Z => n10526);
   U17746 : XOR2_X1 port map( A1 => n18161, A2 => n15237, Z => n10527);
   U17749 : NOR3_X1 port map( A1 => n12060, A2 => n12197, A3 => n20890, ZN => 
                           n10530);
   U17754 : AOI21_X1 port map( A1 => n18606, A2 => n25803, B => n18688, ZN => 
                           n14099);
   U17755 : INV_X1 port map( I => n18688, ZN => n12912);
   U17759 : INV_X1 port map( I => n15909, ZN => n16234);
   U17765 : NAND2_X1 port map( A1 => n17852, A2 => n4508, ZN => n15311);
   U17771 : INV_X1 port map( I => n19357, ZN => n14469);
   U17772 : INV_X1 port map( I => n14550, ZN => n13624);
   U17780 : INV_X2 port map( I => n13420, ZN => n15936);
   U17782 : NOR2_X1 port map( A1 => n561, A2 => n16201, ZN => n16029);
   U17783 : NAND2_X1 port map( A1 => n15885, A2 => n24271, ZN => n14682);
   U17785 : NOR2_X1 port map( A1 => n6688, A2 => n16571, ZN => n12050);
   U17789 : INV_X1 port map( I => n12639, ZN => n11893);
   U17794 : NOR3_X1 port map( A1 => n21798, A2 => n17486, A3 => n17487, ZN => 
                           n15063);
   U17801 : INV_X1 port map( I => n12735, ZN => n11476);
   U17818 : NOR2_X1 port map( A1 => n166, A2 => n18779, ZN => n14829);
   U17823 : NAND2_X1 port map( A1 => n19952, A2 => n19951, ZN => n11464);
   U17829 : NOR2_X1 port map( A1 => n968, A2 => n23977, ZN => n11062);
   U17833 : INV_X1 port map( I => n14854, ZN => n11860);
   U17836 : NAND2_X1 port map( A1 => n12830, A2 => n19974, ZN => n12829);
   U17837 : INV_X2 port map( I => n14529, ZN => n21441);
   U17838 : NOR2_X1 port map( A1 => n13847, A2 => n7904, ZN => n13843);
   U17841 : INV_X1 port map( I => n13600, ZN => n12945);
   U17848 : INV_X1 port map( I => n16331, ZN => n15937);
   U17849 : NOR2_X1 port map( A1 => n16284, A2 => n14218, ZN => n11294);
   U17850 : NOR2_X1 port map( A1 => n11293, A2 => n16278, ZN => n11292);
   U17856 : NAND2_X1 port map( A1 => n16241, A2 => n14557, ZN => n14941);
   U17857 : NOR2_X1 port map( A1 => n21873, A2 => n10970, ZN => n11396);
   U17860 : NAND2_X1 port map( A1 => n16728, A2 => n14364, ZN => n16435);
   U17861 : NAND2_X1 port map( A1 => n14857, A2 => n15930, ZN => n11830);
   U17863 : INV_X1 port map( I => n16656, ZN => n11204);
   U17864 : NAND2_X1 port map( A1 => n16013, A2 => n16011, ZN => n12358);
   U17866 : NOR2_X1 port map( A1 => n14682, A2 => n3298, ZN => n14681);
   U17867 : NAND3_X1 port map( A1 => n10830, A2 => n14306, A3 => n7460, ZN => 
                           n10792);
   U17868 : OAI21_X1 port map( A1 => n14435, A2 => n16271, B => n14434, ZN => 
                           n16079);
   U17869 : NAND2_X1 port map( A1 => n24591, A2 => n21873, ZN => n15269);
   U17870 : NOR2_X1 port map( A1 => n22454, A2 => n24227, ZN => n16085);
   U17872 : NOR2_X1 port map( A1 => n16117, A2 => n8925, ZN => n14267);
   U17876 : NAND2_X1 port map( A1 => n16029, A2 => n3874, ZN => n15596);
   U17879 : NOR2_X1 port map( A1 => n12786, A2 => n1241, ZN => n12785);
   U17883 : NAND2_X1 port map( A1 => n1252, A2 => n8344, ZN => n16382);
   U17885 : NOR2_X1 port map( A1 => n23105, A2 => n8263, ZN => n12193);
   U17889 : NAND2_X1 port map( A1 => n17510, A2 => n17513, ZN => n11943);
   U17892 : NAND3_X1 port map( A1 => n11761, A2 => n12692, A3 => n14103, ZN => 
                           n17218);
   U17895 : NOR2_X1 port map( A1 => n17513, A2 => n24585, ZN => n13933);
   U17898 : NOR2_X1 port map( A1 => n17211, A2 => n11992, ZN => n12397);
   U17901 : OAI21_X1 port map( A1 => n11893, A2 => n11892, B => n14592, ZN => 
                           n12638);
   U17902 : NOR2_X1 port map( A1 => n23276, A2 => n14528, ZN => n11892);
   U17908 : NOR2_X1 port map( A1 => n17416, A2 => n717, ZN => n11571);
   U17909 : OAI21_X1 port map( A1 => n17473, A2 => n11857, B => n13339, ZN => 
                           n17246);
   U17910 : OAI21_X1 port map( A1 => n831, A2 => n1232, B => n22620, ZN => 
                           n14863);
   U17912 : NOR2_X1 port map( A1 => n15592, A2 => n14859, ZN => n14963);
   U17916 : NOR2_X1 port map( A1 => n26939, A2 => n1219, ZN => n14931);
   U17923 : NOR2_X1 port map( A1 => n1175, A2 => n18537, ZN => n18545);
   U17925 : INV_X1 port map( I => n12736, ZN => n11475);
   U17927 : NAND2_X1 port map( A1 => n25592, A2 => n781, ZN => n18992);
   U17928 : AOI21_X1 port map( A1 => n15416, A2 => n10569, B => n18693, ZN => 
                           n12911);
   U17931 : OAI21_X1 port map( A1 => n28542, A2 => n18620, B => n27887, ZN => 
                           n18055);
   U17934 : NAND2_X1 port map( A1 => n18176, A2 => n14245, ZN => n14244);
   U17940 : NOR2_X1 port map( A1 => n6725, A2 => n10924, ZN => n14419);
   U17951 : NAND2_X1 port map( A1 => n25339, A2 => n19006, ZN => n14440);
   U17952 : INV_X1 port map( I => n19643, ZN => n11315);
   U17956 : INV_X1 port map( I => n15118, ZN => n15114);
   U17962 : NOR2_X1 port map( A1 => n19931, A2 => n19930, ZN => n15648);
   U17966 : NAND2_X1 port map( A1 => n19950, A2 => n14651, ZN => n11465);
   U17968 : NAND2_X1 port map( A1 => n974, A2 => n19948, ZN => n14690);
   U17970 : NAND2_X1 port map( A1 => n20317, A2 => n20316, ZN => n13837);
   U17974 : OAI21_X1 port map( A1 => n12287, A2 => n21175, B => n14260, ZN => 
                           n13388);
   U17977 : NOR3_X1 port map( A1 => n10963, A2 => n20225, A3 => n20474, ZN => 
                           n12241);
   U17980 : NOR2_X1 port map( A1 => n22919, A2 => n612, ZN => n20882);
   U17984 : INV_X1 port map( I => n24575, ZN => n20637);
   U17987 : NOR2_X1 port map( A1 => n10558, A2 => n10730, ZN => n20969);
   U17991 : NAND2_X1 port map( A1 => n951, A2 => n11490, ZN => n21509);
   U17993 : NOR2_X1 port map( A1 => n11439, A2 => n20658, ZN => n11438);
   U17995 : NOR2_X1 port map( A1 => n20879, A2 => n20875, ZN => n12728);
   U17996 : INV_X1 port map( I => n21484, ZN => n11739);
   U17997 : NAND2_X1 port map( A1 => n21484, A2 => n21481, ZN => n10833);
   U18002 : NAND2_X1 port map( A1 => n27926, A2 => n13990, ZN => n15134);
   U18003 : AOI21_X1 port map( A1 => n16333, A2 => n7152, B => n14385, ZN => 
                           n15135);
   U18004 : NOR2_X1 port map( A1 => n16307, A2 => n16196, ZN => n16198);
   U18005 : NOR2_X1 port map( A1 => n6237, A2 => n16127, ZN => n15932);
   U18006 : NOR2_X1 port map( A1 => n14442, A2 => n795, ZN => n12875);
   U18007 : INV_X1 port map( I => n14910, ZN => n14907);
   U18010 : NAND2_X1 port map( A1 => n26665, A2 => n15525, ZN => n15987);
   U18011 : NOR2_X1 port map( A1 => n16072, A2 => n16234, ZN => n15633);
   U18012 : AOI22_X1 port map( A1 => n16259, A2 => n14347, B1 => n16236, B2 => 
                           n16258, ZN => n15634);
   U18014 : NAND2_X1 port map( A1 => n15025, A2 => n11024, ZN => n14884);
   U18018 : NAND2_X1 port map( A1 => n12777, A2 => n12776, ZN => n12775);
   U18019 : AOI21_X1 port map( A1 => n16220, A2 => n16253, B => n15812, ZN => 
                           n12776);
   U18023 : NAND2_X1 port map( A1 => n16021, A2 => n16017, ZN => n16018);
   U18025 : NOR2_X1 port map( A1 => n14557, A2 => n16315, ZN => n15074);
   U18026 : NOR2_X1 port map( A1 => n14831, A2 => n16299, ZN => n14830);
   U18029 : OAI21_X1 port map( A1 => n10552, A2 => n14684, B => n16338, ZN => 
                           n11125);
   U18030 : NAND2_X1 port map( A1 => n16333, A2 => n13417, ZN => n14943);
   U18031 : OAI21_X1 port map( A1 => n16145, A2 => n16144, B => n14530, ZN => 
                           n15510);
   U18034 : NAND2_X1 port map( A1 => n16170, A2 => n13742, ZN => n14328);
   U18036 : NAND2_X1 port map( A1 => n1059, A2 => n15611, ZN => n12977);
   U18042 : NAND2_X1 port map( A1 => n7300, A2 => n16196, ZN => n13914);
   U18047 : NAND3_X1 port map( A1 => n13283, A2 => n23880, A3 => n14309, ZN => 
                           n13207);
   U18048 : NAND2_X1 port map( A1 => n26298, A2 => n16677, ZN => n13283);
   U18052 : NAND2_X1 port map( A1 => n10546, A2 => n1224, ZN => n13063);
   U18053 : NAND2_X1 port map( A1 => n900, A2 => n5612, ZN => n11030);
   U18057 : NAND2_X1 port map( A1 => n17738, A2 => n17737, ZN => n12027);
   U18061 : NAND2_X1 port map( A1 => n11716, A2 => n10577, ZN => n11699);
   U18064 : INV_X1 port map( I => n17647, ZN => n15390);
   U18065 : OAI21_X1 port map( A1 => n827, A2 => n8075, B => n14255, ZN => 
                           n14265);
   U18066 : NAND2_X1 port map( A1 => n17473, A2 => n11857, ZN => n15492);
   U18069 : NAND3_X1 port map( A1 => n12964, A2 => n23231, A3 => n28118, ZN => 
                           n17819);
   U18070 : NOR2_X1 port map( A1 => n17262, A2 => n28501, ZN => n11945);
   U18073 : NAND2_X1 port map( A1 => n17981, A2 => n26076, ZN => n17878);
   U18074 : NAND2_X1 port map( A1 => n14707, A2 => n1219, ZN => n14934);
   U18076 : NOR2_X1 port map( A1 => n831, A2 => n1232, ZN => n10954);
   U18081 : NOR2_X1 port map( A1 => n786, A2 => n24175, ZN => n12002);
   U18082 : NOR2_X1 port map( A1 => n5425, A2 => n17757, ZN => n13861);
   U18084 : INV_X1 port map( I => n14589, ZN => n10853);
   U18085 : INV_X1 port map( I => n14544, ZN => n11191);
   U18086 : NAND2_X1 port map( A1 => n11432, A2 => n23926, ZN => n11431);
   U18099 : NAND2_X1 port map( A1 => n13184, A2 => n13532, ZN => n10960);
   U18100 : NOR2_X1 port map( A1 => n166, A2 => n288, ZN => n15000);
   U18102 : NAND2_X1 port map( A1 => n10672, A2 => n18453, ZN => n11387);
   U18104 : NOR2_X1 port map( A1 => n18743, A2 => n10640, ZN => n18405);
   U18108 : NOR3_X1 port map( A1 => n18620, A2 => n1006, A3 => n1187, ZN => 
                           n12379);
   U18110 : NAND2_X1 port map( A1 => n19008, A2 => n736, ZN => n18952);
   U18112 : NAND2_X1 port map( A1 => n13946, A2 => n13873, ZN => n18730);
   U18114 : NAND2_X1 port map( A1 => n18388, A2 => n18390, ZN => n14922);
   U18115 : INV_X1 port map( I => n15266, ZN => n13483);
   U18116 : INV_X1 port map( I => n11983, ZN => n11826);
   U18118 : NAND2_X1 port map( A1 => n26036, A2 => n18728, ZN => n11618);
   U18119 : NOR2_X1 port map( A1 => n18690, A2 => n13646, ZN => n18691);
   U18122 : NOR2_X1 port map( A1 => n18873, A2 => n23305, ZN => n12576);
   U18123 : NOR2_X1 port map( A1 => n3057, A2 => n19062, ZN => n11117);
   U18125 : NOR2_X1 port map( A1 => n992, A2 => n7084, ZN => n15530);
   U18129 : NOR2_X1 port map( A1 => n1164, A2 => n14358, ZN => n11626);
   U18131 : INV_X1 port map( I => n19233, ZN => n19338);
   U18132 : NOR2_X1 port map( A1 => n27026, A2 => n18556, ZN => n15243);
   U18133 : INV_X1 port map( I => n26962, ZN => n15230);
   U18134 : NAND2_X1 port map( A1 => n15250, A2 => n19793, ZN => n15277);
   U18139 : NOR3_X1 port map( A1 => n19857, A2 => n19858, A3 => n1119, ZN => 
                           n11985);
   U18141 : NOR2_X1 port map( A1 => n11936, A2 => n10562, ZN => n11901);
   U18143 : NAND2_X1 port map( A1 => n14740, A2 => n20189, ZN => n19361);
   U18144 : INV_X1 port map( I => n12594, ZN => n12593);
   U18146 : NOR2_X1 port map( A1 => n15268, A2 => n19822, ZN => n12440);
   U18147 : NOR2_X1 port map( A1 => n20194, A2 => n20294, ZN => n14974);
   U18151 : INV_X1 port map( I => n20323, ZN => n19962);
   U18153 : NOR2_X1 port map( A1 => n7767, A2 => n19808, ZN => n12159);
   U18158 : INV_X1 port map( I => n15117, ZN => n15115);
   U18159 : INV_X1 port map( I => n19673, ZN => n15116);
   U18161 : OAI22_X1 port map( A1 => n15146, A2 => n10770, B1 => n26807, B2 => 
                           n23065, ZN => n15145);
   U18162 : NAND2_X1 port map( A1 => n12267, A2 => n12266, ZN => n12264);
   U18167 : NAND2_X1 port map( A1 => n19682, A2 => n15067, ZN => n11856);
   U18171 : NAND2_X1 port map( A1 => n20292, A2 => n13252, ZN => n11541);
   U18172 : NAND2_X1 port map( A1 => n25843, A2 => n23592, ZN => n13098);
   U18175 : NOR2_X1 port map( A1 => n22295, A2 => n22776, ZN => n12491);
   U18176 : INV_X1 port map( I => n21059, ZN => n15721);
   U18181 : NAND2_X1 port map( A1 => n21058, A2 => n14341, ZN => n11017);
   U18189 : INV_X1 port map( I => n11166, ZN => n11165);
   U18190 : OAI22_X1 port map( A1 => n21043, A2 => n21050, B1 => n9422, B2 => 
                           n21042, ZN => n12073);
   U18191 : INV_X1 port map( I => n15169, ZN => n11031);
   U18192 : OAI21_X1 port map( A1 => n21698, A2 => n21697, B => n21696, ZN => 
                           n12019);
   U18195 : NAND2_X1 port map( A1 => n20998, A2 => n21000, ZN => n12082);
   U18199 : OAI21_X1 port map( A1 => n12046, A2 => n12045, B => n12044, ZN => 
                           n12540);
   U18201 : OAI22_X1 port map( A1 => n1515, A2 => n21713, B1 => n8757, B2 => 
                           n15706, ZN => n12752);
   U18202 : NAND2_X1 port map( A1 => n13879, A2 => n20895, ZN => n13878);
   U18203 : NOR2_X1 port map( A1 => n20895, A2 => n20899, ZN => n12126);
   U18206 : INV_X1 port map( I => n7516, ZN => n12417);
   U18207 : INV_X1 port map( I => n20785, ZN => n20738);
   U18213 : NAND2_X1 port map( A1 => n13846, A2 => n27512, ZN => n13841);
   U18214 : INV_X1 port map( I => n14460, ZN => n13846);
   U18215 : NAND2_X1 port map( A1 => n21203, A2 => n13424, ZN => n10928);
   U18216 : NAND2_X1 port map( A1 => n3549, A2 => n13772, ZN => n14539);
   U18217 : NAND2_X1 port map( A1 => n14873, A2 => n21396, ZN => n12652);
   U18218 : AOI21_X1 port map( A1 => n13790, A2 => n26505, B => n12296, ZN => 
                           n12295);
   U18223 : OAI21_X1 port map( A1 => n21593, A2 => n951, B => n12900, ZN => 
                           n21551);
   U18228 : AOI21_X1 port map( A1 => n21546, A2 => n13426, B => n11201, ZN => 
                           n11200);
   U18229 : NAND2_X1 port map( A1 => n13103, A2 => n16082, ZN => n12777);
   U18231 : INV_X1 port map( I => n12529, ZN => n15347);
   U18233 : INV_X1 port map( I => n16550, ZN => n15548);
   U18242 : OAI22_X1 port map( A1 => n15983, A2 => n15984, B1 => n16021, B2 => 
                           n14530, ZN => n15827);
   U18250 : INV_X1 port map( I => n23505, ZN => n12223);
   U18255 : NAND3_X1 port map( A1 => n1257, A2 => n26993, A3 => n794, ZN => 
                           n14864);
   U18260 : NAND2_X1 port map( A1 => n14802, A2 => n15061, ZN => n14801);
   U18269 : NAND3_X1 port map( A1 => n16605, A2 => n4060, A3 => n16055, ZN => 
                           n15370);
   U18274 : AOI21_X1 port map( A1 => n5062, A2 => n16632, B => n718, ZN => 
                           n12212);
   U18276 : NOR2_X1 port map( A1 => n17516, A2 => n3545, ZN => n11590);
   U18277 : NOR2_X1 port map( A1 => n17517, A2 => n15037, ZN => n11591);
   U18279 : OAI21_X1 port map( A1 => n899, A2 => n242, B => n17185, ZN => 
                           n12506);
   U18280 : INV_X1 port map( I => n18088, ZN => n18329);
   U18283 : INV_X1 port map( I => n17906, ZN => n17948);
   U18285 : NAND2_X1 port map( A1 => n17800, A2 => n9772, ZN => n14112);
   U18286 : NAND2_X1 port map( A1 => n17880, A2 => n17597, ZN => n14111);
   U18290 : NAND2_X1 port map( A1 => n7358, A2 => n17783, ZN => n15533);
   U18305 : INV_X1 port map( I => n14659, ZN => n10784);
   U18308 : NAND2_X1 port map( A1 => n17744, A2 => n25929, ZN => n12166);
   U18315 : NOR2_X1 port map( A1 => n14446, A2 => n17927, ZN => n12516);
   U18316 : NAND3_X1 port map( A1 => n17986, A2 => n12611, A3 => n17751, ZN => 
                           n17705);
   U18319 : NOR2_X1 port map( A1 => n4802, A2 => n12257, ZN => n13862);
   U18322 : INV_X1 port map( I => n17887, ZN => n17972);
   U18323 : INV_X1 port map( I => n18180, ZN => n12824);
   U18324 : OAI21_X1 port map( A1 => n17906, A2 => n17694, B => n25724, ZN => 
                           n11281);
   U18325 : INV_X1 port map( I => n17645, ZN => n11282);
   U18326 : INV_X1 port map( I => n11559, ZN => n19205);
   U18327 : INV_X1 port map( I => n25006, ZN => n14325);
   U18328 : NAND2_X1 port map( A1 => n13946, A2 => n19134, ZN => n18822);
   U18329 : NOR2_X1 port map( A1 => n18959, A2 => n27043, ZN => n15202);
   U18331 : INV_X1 port map( I => n14095, ZN => n13886);
   U18332 : INV_X1 port map( I => n18771, ZN => n13885);
   U18336 : NAND3_X1 port map( A1 => n8714, A2 => n11718, A3 => n19033, ZN => 
                           n18864);
   U18343 : NAND3_X1 port map( A1 => n18619, A2 => n18617, A3 => n18618, ZN => 
                           n12772);
   U18344 : INV_X1 port map( I => n13045, ZN => n12227);
   U18345 : INV_X1 port map( I => n13046, ZN => n12226);
   U18346 : NAND2_X1 port map( A1 => n23017, A2 => n7390, ZN => n12495);
   U18347 : NOR2_X1 port map( A1 => n19052, A2 => n24061, ZN => n13972);
   U18349 : INV_X1 port map( I => n14479, ZN => n12327);
   U18350 : NAND2_X1 port map( A1 => n19133, A2 => n12113, ZN => n12138);
   U18353 : NOR2_X1 port map( A1 => n18392, A2 => n19152, ZN => n18394);
   U18360 : INV_X1 port map( I => n14779, ZN => n18935);
   U18363 : NAND2_X1 port map( A1 => n19989, A2 => n13248, ZN => n20019);
   U18368 : INV_X1 port map( I => n14855, ZN => n11859);
   U18369 : NAND2_X1 port map( A1 => n14217, A2 => n14216, ZN => n15281);
   U18370 : NAND2_X1 port map( A1 => n15276, A2 => n12570, ZN => n14216);
   U18371 : NOR2_X1 port map( A1 => n15278, A2 => n15277, ZN => n15276);
   U18372 : NOR2_X1 port map( A1 => n23592, A2 => n8032, ZN => n13091);
   U18374 : INV_X1 port map( I => n20019, ZN => n11670);
   U18378 : NAND2_X1 port map( A1 => n20323, A2 => n1731, ZN => n20496);
   U18379 : OR2_X1 port map( A1 => n20328, A2 => n4738, Z => n10741);
   U18380 : INV_X1 port map( I => n15151, ZN => n15150);
   U18381 : INV_X1 port map( I => n25362, ZN => n15651);
   U18387 : NAND2_X1 port map( A1 => n20224, A2 => n20059, ZN => n10938);
   U18390 : NAND2_X1 port map( A1 => n19985, A2 => n20338, ZN => n14497);
   U18391 : INV_X1 port map( I => n20431, ZN => n20201);
   U18393 : NAND2_X1 port map( A1 => n855, A2 => n4225, ZN => n15369);
   U18394 : NOR2_X1 port map( A1 => n11757, A2 => n12477, ZN => n14063);
   U18395 : NOR2_X1 port map( A1 => n11372, A2 => n20165, ZN => n12922);
   U18396 : NAND2_X1 port map( A1 => n15320, A2 => n11052, ZN => n14262);
   U18401 : OAI21_X1 port map( A1 => n14153, A2 => n675, B => n14481, ZN => 
                           n14952);
   U18403 : NAND3_X1 port map( A1 => n12712, A2 => n20323, A3 => n1731, ZN => 
                           n19998);
   U18406 : NAND2_X1 port map( A1 => n27630, A2 => n183, ZN => n13074);
   U18407 : NAND3_X1 port map( A1 => n15334, A2 => n22779, A3 => n1114, ZN => 
                           n15333);
   U18411 : INV_X1 port map( I => n14811, ZN => n14810);
   U18412 : NAND2_X1 port map( A1 => n22745, A2 => n26710, ZN => n11073);
   U18414 : NAND2_X1 port map( A1 => n10666, A2 => n20642, ZN => n15325);
   U18415 : INV_X1 port map( I => n20000, ZN => n11926);
   U18416 : NAND2_X1 port map( A1 => n20184, A2 => n15193, ZN => n15192);
   U18417 : NAND2_X1 port map( A1 => n10616, A2 => n20183, ZN => n13233);
   U18422 : NAND2_X1 port map( A1 => n1105, A2 => n11747, ZN => n11746);
   U18424 : NAND3_X1 port map( A1 => n14292, A2 => n20210, A3 => n20209, ZN => 
                           n20037);
   U18425 : INV_X1 port map( I => n13585, ZN => n13599);
   U18427 : INV_X1 port map( I => n27877, ZN => n16095);
   U18429 : NAND2_X1 port map( A1 => n14385, A2 => n16334, ZN => n13989);
   U18431 : NOR2_X1 port map( A1 => n12056, A2 => n12055, ZN => n12054);
   U18432 : NOR2_X1 port map( A1 => n21457, A2 => n26505, ZN => n11978);
   U18434 : NAND2_X1 port map( A1 => n1077, A2 => n21620, ZN => n11736);
   U18436 : NAND2_X1 port map( A1 => n21669, A2 => n10591, ZN => n15483);
   U18438 : NOR2_X1 port map( A1 => n22794, A2 => n21413, ZN => n11467);
   U18439 : NAND2_X1 port map( A1 => n21173, A2 => n21172, ZN => n15653);
   U18440 : NAND2_X1 port map( A1 => n13768, A2 => n15524, ZN => n21163);
   U18443 : NOR2_X1 port map( A1 => n10878, A2 => n11622, ZN => n11865);
   U18445 : NOR2_X1 port map( A1 => n803, A2 => n7009, ZN => n21639);
   U18447 : NAND2_X1 port map( A1 => n20847, A2 => n20850, ZN => n11321);
   U18449 : OAI21_X1 port map( A1 => n800, A2 => n22536, B => n20798, ZN => 
                           n20793);
   U18450 : INV_X1 port map( I => n25360, ZN => n20837);
   U18452 : OAI21_X1 port map( A1 => n10608, A2 => n14860, B => n10031, ZN => 
                           n13106);
   U18456 : NOR2_X1 port map( A1 => n11850, A2 => n11849, ZN => n11848);
   U18457 : NOR2_X1 port map( A1 => n23579, A2 => n10851, ZN => n11766);
   U18462 : INV_X1 port map( I => n21659, ZN => n21653);
   U18463 : NAND2_X1 port map( A1 => n21405, A2 => n12650, ZN => n21402);
   U18464 : NAND2_X1 port map( A1 => n20874, A2 => n20876, ZN => n12684);
   U18465 : INV_X1 port map( I => n14645, ZN => n15195);
   U18470 : INV_X1 port map( I => n20999, ZN => n12538);
   U18471 : INV_X1 port map( I => n14436, ZN => n13082);
   U18472 : NAND2_X1 port map( A1 => n20749, A2 => n6051, ZN => n14242);
   U18474 : INV_X1 port map( I => n21000, ZN => n12188);
   U18475 : NAND2_X1 port map( A1 => n21165, A2 => n21168, ZN => n12845);
   U18480 : OAI21_X1 port map( A1 => n27404, A2 => n10674, B => n12399, ZN => 
                           n21596);
   U18481 : NAND2_X1 port map( A1 => n21648, A2 => n438, ZN => n15426);
   U18482 : INV_X1 port map( I => n14637, ZN => n15519);
   U18484 : NOR2_X1 port map( A1 => n8173, A2 => n13613, ZN => n10552);
   U18486 : INV_X1 port map( I => n10359, ZN => n10878);
   U18487 : XNOR2_X1 port map( A1 => n10948, A2 => n10946, ZN => n10570);
   U18488 : AND2_X1 port map( A1 => n721, A2 => n22821, Z => n10576);
   U18489 : AND2_X1 port map( A1 => n20338, A2 => n20152, Z => n10582);
   U18496 : XNOR2_X1 port map( A1 => n16993, A2 => n1308, ZN => n10612);
   U18497 : INV_X1 port map( I => n13738, ZN => n13093);
   U18502 : NOR2_X1 port map( A1 => n20263, A2 => n13600, ZN => n10623);
   U18511 : XNOR2_X1 port map( A1 => n22741, A2 => n20766, ZN => n10646);
   U18512 : XNOR2_X1 port map( A1 => n20350, A2 => n20349, ZN => n10647);
   U18513 : XNOR2_X1 port map( A1 => n20356, A2 => n20357, ZN => n10648);
   U18520 : AND2_X1 port map( A1 => n940, A2 => n21608, Z => n10664);
   U18524 : XNOR2_X1 port map( A1 => n6878, A2 => n25358, ZN => n10676);
   U18525 : AND2_X1 port map( A1 => n18668, A2 => n18432, Z => n10677);
   U18527 : XNOR2_X1 port map( A1 => n18046, A2 => n18045, ZN => n10678);
   U18529 : XNOR2_X1 port map( A1 => n21357, A2 => n18258, ZN => n10680);
   U18531 : OR2_X1 port map( A1 => n6892, A2 => n24564, Z => n10691);
   U18533 : AND2_X1 port map( A1 => n11668, A2 => n10898, Z => n10695);
   U18534 : NOR2_X1 port map( A1 => n15347, A2 => n13435, ZN => n10697);
   U18535 : NAND2_X1 port map( A1 => n28525, A2 => n20200, ZN => n10701);
   U18539 : XNOR2_X1 port map( A1 => n19432, A2 => n14526, ZN => n10713);
   U18540 : XNOR2_X1 port map( A1 => n15754, A2 => n19517, ZN => n10715);
   U18541 : XNOR2_X1 port map( A1 => n20347, A2 => n20346, ZN => n10716);
   U18543 : INV_X1 port map( I => n20816, ZN => n20593);
   U18546 : XOR2_X1 port map( A1 => n1197, A2 => n23354, Z => n10729);
   U18551 : INV_X1 port map( I => n17924, ZN => n17584);
   U18552 : XNOR2_X1 port map( A1 => n18161, A2 => n21642, ZN => n10734);
   U18555 : XNOR2_X1 port map( A1 => n6490, A2 => n21210, ZN => n10737);
   U18558 : INV_X1 port map( I => n14886, ZN => n16305);
   U18559 : XOR2_X1 port map( A1 => n23849, A2 => n23554, Z => n10747);
   U18560 : XNOR2_X1 port map( A1 => n19388, A2 => n14560, ZN => n10749);
   U18561 : XNOR2_X1 port map( A1 => n21318, A2 => n20404, ZN => n10751);
   U18562 : XNOR2_X1 port map( A1 => n27661, A2 => n14550, ZN => n10752);
   U18565 : INV_X1 port map( I => n17180, ZN => n17567);
   U18566 : INV_X1 port map( I => n18914, ZN => n19041);
   U18568 : INV_X1 port map( I => n15848, ZN => n16201);
   U18571 : XNOR2_X1 port map( A1 => n22757, A2 => n21476, ZN => n10766);
   U18573 : INV_X1 port map( I => n14414, ZN => n11160);
   U18576 : INV_X2 port map( I => n15344, ZN => n14103);
   U18580 : XNOR2_X1 port map( A1 => n94, A2 => n21707, ZN => n10772);
   U18581 : INV_X1 port map( I => n15506, ZN => n15149);
   U18582 : INV_X1 port map( I => n21683, ZN => n11181);
   U18583 : INV_X1 port map( I => n14572, ZN => n15271);
   U18587 : INV_X1 port map( I => n14457, ZN => n13746);
   U18588 : INV_X1 port map( I => n14535, ZN => n15680);
   U18589 : INV_X1 port map( I => n20671, ZN => n11918);
   U18590 : INV_X1 port map( I => n7409, ZN => n12769);
   U18591 : INV_X1 port map( I => n7387, ZN => n11152);
   U18592 : INV_X1 port map( I => n21705, ZN => n13285);
   U18593 : INV_X1 port map( I => n14540, ZN => n13200);
   U18594 : INV_X1 port map( I => n20396, ZN => n21048);
   U18595 : INV_X1 port map( I => n21010, ZN => n14007);
   U18597 : INV_X1 port map( I => n7365, ZN => n13678);
   U18598 : INV_X1 port map( I => n20321, ZN => n15669);
   U18599 : INV_X1 port map( I => Key(59), ZN => n13738);
   U18602 : INV_X1 port map( I => n21554, ZN => n12813);
   U18604 : INV_X1 port map( I => n21039, ZN => n12713);
   U18606 : INV_X1 port map( I => n20873, ZN => n11975);
   U18607 : XOR2_X1 port map( A1 => n10773, A2 => n16965, Z => n11935);
   U18608 : NAND3_X1 port map( A1 => n12260, A2 => n19198, A3 => n12259, ZN => 
                           n10774);
   U18611 : OAI21_X1 port map( A1 => n7180, A2 => n26734, B => n10777, ZN => 
                           n15179);
   U18615 : XOR2_X1 port map( A1 => n10785, A2 => n10783, Z => n10787);
   U18616 : XOR2_X1 port map( A1 => n22774, A2 => n10784, Z => n10783);
   U18617 : XOR2_X1 port map( A1 => n10786, A2 => n7244, Z => n10785);
   U18621 : OAI21_X1 port map( A1 => n21359, A2 => n10547, B => n26651, ZN => 
                           n21362);
   U18622 : NAND2_X1 port map( A1 => n713, A2 => n2895, ZN => n17861);
   U18626 : OAI21_X1 port map( A1 => n1065, A2 => n26647, B => n14350, ZN => 
                           n21735);
   U18629 : INV_X2 port map( I => n10813, ZN => n14306);
   U18630 : INV_X2 port map( I => n10815, ZN => n13184);
   U18636 : NOR2_X1 port map( A1 => n9916, A2 => n11089, ZN => n10829);
   U18638 : XOR2_X1 port map( A1 => n13253, A2 => n14633, Z => n14668);
   U18642 : INV_X2 port map( I => n10838, ZN => n14859);
   U18643 : XOR2_X1 port map( A1 => n17132, A2 => n16779, Z => n10839);
   U18646 : NAND2_X1 port map( A1 => n10844, A2 => n12463, ZN => n11849);
   U18648 : XOR2_X1 port map( A1 => Plaintext(76), A2 => Key(76), Z => n12271);
   U18649 : INV_X1 port map( I => n20070, ZN => n15178);
   U18656 : XOR2_X1 port map( A1 => n17150, A2 => n10855, Z => n10854);
   U18659 : AOI21_X1 port map( A1 => n20998, A2 => n10858, B => n12179, ZN => 
                           n11345);
   U18670 : XOR2_X1 port map( A1 => n11405, A2 => n17721, Z => n10880);
   U18673 : OAI21_X1 port map( A1 => n12934, A2 => n12935, B => n15503, ZN => 
                           n10889);
   U18674 : NOR2_X1 port map( A1 => n24188, A2 => n25984, ZN => n18960);
   U18676 : AOI21_X1 port map( A1 => n16077, A2 => n27123, B => n10905, ZN => 
                           n15968);
   U18677 : XOR2_X1 port map( A1 => n10906, A2 => n16944, Z => n16945);
   U18680 : XOR2_X1 port map( A1 => n26058, A2 => n14463, Z => n10917);
   U18681 : XOR2_X1 port map( A1 => n10950, A2 => n10922, Z => n10921);
   U18682 : XOR2_X1 port map( A1 => n20584, A2 => n21435, Z => n10922);
   U18683 : XOR2_X1 port map( A1 => n16744, A2 => n11680, Z => n10968);
   U18684 : XOR2_X1 port map( A1 => n11680, A2 => n17141, Z => n16947);
   U18685 : XOR2_X1 port map( A1 => n11680, A2 => n17097, Z => n16865);
   U18687 : XOR2_X1 port map( A1 => n21180, A2 => n11153, Z => n10926);
   U18689 : XOR2_X1 port map( A1 => n4877, A2 => n20607, Z => n10934);
   U18691 : INV_X2 port map( I => n10570, ZN => n10941);
   U18693 : XOR2_X1 port map( A1 => n10641, A2 => n10947, Z => n10946);
   U18694 : XOR2_X1 port map( A1 => n18210, A2 => n18056, Z => n10948);
   U18696 : XOR2_X1 port map( A1 => n6932, A2 => n16937, Z => n17130);
   U18698 : NAND2_X1 port map( A1 => n51, A2 => n9308, ZN => n12105);
   U18699 : OAI21_X1 port map( A1 => n16338, A2 => n9308, B => n16339, ZN => 
                           n12106);
   U18701 : XOR2_X1 port map( A1 => n13064, A2 => n9876, Z => n11034);
   U18706 : XOR2_X1 port map( A1 => n11678, A2 => n10968, Z => n11677);
   U18707 : XOR2_X1 port map( A1 => Plaintext(3), A2 => Key(3), Z => n11395);
   U18710 : XOR2_X1 port map( A1 => n16965, A2 => n14619, Z => n16966);
   U18716 : XOR2_X1 port map( A1 => n18330, A2 => n18088, Z => n10998);
   U18721 : XOR2_X1 port map( A1 => n17008, A2 => n12291, Z => n11003);
   U18722 : XOR2_X1 port map( A1 => n27425, A2 => n1273, Z => n11010);
   U18723 : INV_X1 port map( I => n25342, ZN => n21126);
   U18724 : AND2_X1 port map( A1 => n21118, A2 => n21120, Z => n11012);
   U18725 : XOR2_X1 port map( A1 => n18061, A2 => n21557, Z => n11014);
   U18730 : XOR2_X1 port map( A1 => n11022, A2 => n14598, Z => n18199);
   U18731 : XOR2_X1 port map( A1 => n11022, A2 => n21631, Z => n18287);
   U18732 : XOR2_X1 port map( A1 => Key(97), A2 => Plaintext(97), Z => n11024);
   U18733 : NOR2_X1 port map( A1 => n22800, A2 => n25304, ZN => n11032);
   U18736 : XOR2_X1 port map( A1 => n6765, A2 => n17055, Z => n11038);
   U18737 : NOR2_X2 port map( A1 => n11039, A2 => n12785, ZN => n17055);
   U18739 : XOR2_X1 port map( A1 => n11046, A2 => n12816, Z => n14840);
   U18740 : XOR2_X1 port map( A1 => n11046, A2 => n20763, Z => n20384);
   U18742 : NOR2_X1 port map( A1 => n26154, A2 => n11052, ZN => n14261);
   U18743 : NAND2_X2 port map( A1 => n11976, A2 => n21458, ZN => n21484);
   U18745 : INV_X2 port map( I => n13491, ZN => n21730);
   U18748 : AND2_X1 port map( A1 => n16217, A2 => n11080, Z => n11084);
   U18751 : XOR2_X1 port map( A1 => n14669, A2 => n14668, Z => n11090);
   U18757 : NOR2_X1 port map( A1 => n27368, A2 => n12191, ZN => n11108);
   U18762 : XOR2_X1 port map( A1 => n23314, A2 => n20459, Z => n11141);
   U18764 : XOR2_X1 port map( A1 => n6996, A2 => n21703, Z => n11153);
   U18765 : NOR2_X1 port map( A1 => n21347, A2 => n2447, ZN => n14079);
   U18766 : NOR3_X1 port map( A1 => n2447, A2 => n21355, A3 => n21344, ZN => 
                           n21335);
   U18767 : NOR2_X1 port map( A1 => n21340, A2 => n2447, ZN => n21338);
   U18768 : AOI21_X1 port map( A1 => n21348, A2 => n2447, B => n21347, ZN => 
                           n21349);
   U18771 : NAND2_X2 port map( A1 => n21393, A2 => n11163, ZN => n13741);
   U18774 : XOR2_X1 port map( A1 => n4020, A2 => n11177, Z => n11176);
   U18775 : XOR2_X1 port map( A1 => n26962, A2 => n19451, Z => n11177);
   U18776 : XOR2_X1 port map( A1 => n11174, A2 => n19452, Z => n11178);
   U18777 : XOR2_X1 port map( A1 => n11179, A2 => n20382, Z => n20816);
   U18778 : XOR2_X1 port map( A1 => n13458, A2 => n11180, Z => n11179);
   U18779 : XOR2_X1 port map( A1 => n14421, A2 => n20603, Z => n11180);
   U18783 : XOR2_X1 port map( A1 => n18132, A2 => n11191, Z => n11190);
   U18787 : INV_X1 port map( I => n21622, ZN => n11201);
   U18789 : NAND2_X1 port map( A1 => n12712, A2 => n26485, ZN => n11214);
   U18790 : XOR2_X1 port map( A1 => n28265, A2 => n23375, Z => n11222);
   U18791 : OAI22_X1 port map( A1 => n18822, A2 => n28507, B1 => n1159, B2 => 
                           n13946, ZN => n18823);
   U18792 : XOR2_X1 port map( A1 => n13513, A2 => n11234, Z => n11233);
   U18794 : XOR2_X1 port map( A1 => n28488, A2 => n21594, Z => n11244);
   U18795 : XOR2_X1 port map( A1 => n19071, A2 => n5147, Z => n11245);
   U18796 : XOR2_X1 port map( A1 => n11247, A2 => n11246, Z => n11287);
   U18797 : XOR2_X1 port map( A1 => n19404, A2 => n10615, Z => n11246);
   U18799 : NAND2_X2 port map( A1 => n28554, A2 => n11251, ZN => n21636);
   U18800 : NAND4_X1 port map( A1 => n28554, A2 => n11250, A3 => n11249, A4 => 
                           n11251, ZN => n21640);
   U18801 : XOR2_X1 port map( A1 => n28527, A2 => n20650, Z => n11253);
   U18803 : XOR2_X1 port map( A1 => n20434, A2 => n27447, Z => n11900);
   U18805 : NAND2_X1 port map( A1 => n11262, A2 => n14427, ZN => n18726);
   U18807 : XOR2_X1 port map( A1 => n11278, A2 => n13504, Z => n11277);
   U18810 : INV_X1 port map( I => n20614, ZN => n11288);
   U18816 : XOR2_X1 port map( A1 => n9455, A2 => n20949, Z => n13729);
   U18818 : OAI21_X1 port map( A1 => n20844, A2 => n20850, B => n11320, ZN => 
                           n20845);
   U18821 : XOR2_X1 port map( A1 => n19292, A2 => n18790, Z => n11322);
   U18822 : XOR2_X1 port map( A1 => n19559, A2 => n13825, Z => n19292);
   U18824 : XOR2_X1 port map( A1 => n3506, A2 => n20508, Z => n20455);
   U18825 : INV_X2 port map( I => n11326, ZN => n21501);
   U18827 : XOR2_X1 port map( A1 => n17019, A2 => n11337, Z => n11336);
   U18835 : OAI21_X1 port map( A1 => n3954, A2 => n11353, B => n19696, ZN => 
                           n19663);
   U18836 : NAND2_X1 port map( A1 => n19784, A2 => n19661, ZN => n11353);
   U18839 : INV_X2 port map( I => n12549, ZN => n14592);
   U18843 : XOR2_X1 port map( A1 => n28263, A2 => n19201, Z => n18900);
   U18844 : XOR2_X1 port map( A1 => n13996, A2 => n13285, Z => n13648);
   U18845 : XOR2_X1 port map( A1 => n18263, A2 => n13996, Z => n11525);
   U18846 : XOR2_X1 port map( A1 => n12246, A2 => n6535, Z => n12355);
   U18847 : INV_X1 port map( I => n11373, ZN => n17505);
   U18849 : NAND2_X1 port map( A1 => n11378, A2 => n11377, ZN => n15160);
   U18852 : OAI21_X2 port map( A1 => n867, A2 => n19915, B => n19575, ZN => 
                           n19097);
   U18857 : NAND2_X1 port map( A1 => n11390, A2 => n11424, ZN => n16449);
   U18859 : XOR2_X1 port map( A1 => n16950, A2 => n21553, Z => n11397);
   U18860 : INV_X2 port map( I => n11404, ZN => n18665);
   U18861 : XOR2_X1 port map( A1 => n18215, A2 => n5890, Z => n11405);
   U18865 : XOR2_X1 port map( A1 => n11417, A2 => n20621, Z => n19239);
   U18866 : MUX2_X1 port map( I0 => n19937, I1 => n12617, S => n7176, Z => 
                           n19604);
   U18867 : NAND2_X1 port map( A1 => n13572, A2 => n16530, ZN => n11422);
   U18869 : XOR2_X1 port map( A1 => n19240, A2 => n10646, Z => n11427);
   U18870 : XOR2_X1 port map( A1 => n24885, A2 => n14637, Z => n11430);
   U18874 : NAND2_X1 port map( A1 => n3948, A2 => n16380, ZN => n16177);
   U18875 : NAND2_X1 port map( A1 => n11453, A2 => n14097, ZN => n18690);
   U18876 : NAND2_X1 port map( A1 => n18385, A2 => n18687, ZN => n11452);
   U18877 : NOR2_X1 port map( A1 => n18608, A2 => n11453, ZN => n18606);
   U18879 : MUX2_X1 port map( I0 => n18693, I1 => n10569, S => n18687, Z => 
                           n15718);
   U18880 : INV_X1 port map( I => n21413, ZN => n12650);
   U18881 : NAND3_X1 port map( A1 => n21409, A2 => n13741, A3 => n21408, ZN => 
                           n11456);
   U18882 : NAND2_X1 port map( A1 => n11458, A2 => n21412, ZN => n11457);
   U18883 : NOR2_X1 port map( A1 => n21413, A2 => n13741, ZN => n11458);
   U18884 : NAND2_X1 port map( A1 => n15461, A2 => n11871, ZN => n11463);
   U18889 : XOR2_X1 port map( A1 => n19528, A2 => n11481, Z => n11480);
   U18890 : XOR2_X1 port map( A1 => n27422, A2 => n25376, Z => n11481);
   U18894 : INV_X1 port map( I => n18913, ZN => n11486);
   U18897 : INV_X2 port map( I => n15636, ZN => n21499);
   U18898 : NAND2_X1 port map( A1 => n7941, A2 => n27467, ZN => n21467);
   U18899 : NAND2_X2 port map( A1 => n14100, A2 => n14099, ZN => n14098);
   U18903 : XOR2_X1 port map( A1 => n3291, A2 => n20603, Z => n11512);
   U18904 : XOR2_X1 port map( A1 => n19173, A2 => n18928, Z => n11513);
   U18908 : NAND2_X1 port map( A1 => n11522, A2 => n21110, ZN => n13011);
   U18915 : XOR2_X1 port map( A1 => n7200, A2 => n25808, Z => n11535);
   U18917 : XOR2_X1 port map( A1 => n9455, A2 => n16875, Z => n11539);
   U18919 : NAND2_X2 port map( A1 => n11545, A2 => n16352, ZN => n16571);
   U18920 : NAND2_X2 port map( A1 => n18733, A2 => n18732, ZN => n19375);
   U18922 : XOR2_X1 port map( A1 => n11555, A2 => n14436, Z => n18014);
   U18924 : NAND2_X1 port map( A1 => n14826, A2 => n24570, ZN => n17999);
   U18925 : NOR2_X2 port map( A1 => n11566, A2 => n14681, ZN => n16516);
   U18926 : XOR2_X1 port map( A1 => n25317, A2 => n9123, Z => n11574);
   U18933 : XOR2_X1 port map( A1 => n1097, A2 => n15537, Z => n11592);
   U18936 : XOR2_X1 port map( A1 => n11601, A2 => n14418, Z => Ciphertext(95));
   U18937 : XOR2_X1 port map( A1 => Plaintext(172), A2 => Key(172), Z => n11628
                           );
   U18939 : NAND2_X1 port map( A1 => n12949, A2 => n1253, ZN => n12423);
   U18942 : AOI21_X1 port map( A1 => n17871, A2 => n12983, B => n17872, ZN => 
                           n17704);
   U18946 : INV_X1 port map( I => n19804, ZN => n15278);
   U18948 : NAND3_X1 port map( A1 => n19644, A2 => n19866, A3 => n19643, ZN => 
                           n12184);
   U18954 : INV_X1 port map( I => n13320, ZN => n17540);
   U18957 : NAND2_X1 port map( A1 => n20816, A2 => n20817, ZN => n13287);
   U18961 : NAND3_X1 port map( A1 => n9661, A2 => n8165, A3 => n17509, ZN => 
                           n13218);
   U18962 : NAND2_X1 port map( A1 => n27241, A2 => n18454, ZN => n18380);
   U18964 : NAND2_X1 port map( A1 => n28300, A2 => n9005, ZN => n11802);
   U18965 : INV_X1 port map( I => n25306, ZN => n13468);
   U18977 : NOR2_X1 port map( A1 => n14909, A2 => n21764, ZN => n13220);
   U18981 : NAND2_X1 port map( A1 => n20842, A2 => n13056, ZN => n20835);
   U18983 : INV_X1 port map( I => Key(40), ZN => n15506);
   U18985 : INV_X1 port map( I => n18600, ZN => n18412);
   U18988 : AOI21_X1 port map( A1 => n26435, A2 => n13979, B => n23991, ZN => 
                           n11735);
   U18999 : XOR2_X1 port map( A1 => Plaintext(170), A2 => Key(170), Z => n11813
                           );
   U19001 : AOI21_X1 port map( A1 => n21484, A2 => n694, B => n11622, ZN => 
                           n11623);
   U19004 : NAND2_X1 port map( A1 => n11817, A2 => n13532, ZN => n15084);
   U19006 : AOI21_X1 port map( A1 => n11627, A2 => n22789, B => n21564, ZN => 
                           n12904);
   U19008 : NAND2_X2 port map( A1 => n16091, A2 => n16090, ZN => n16534);
   U19011 : OR2_X1 port map( A1 => n13943, A2 => n21703, Z => n11645);
   U19012 : XOR2_X1 port map( A1 => n11649, A2 => n11648, Z => n11714);
   U19013 : XOR2_X1 port map( A1 => n25328, A2 => n14593, Z => n11648);
   U19018 : XOR2_X1 port map( A1 => n17035, A2 => n11671, Z => n14143);
   U19019 : XOR2_X1 port map( A1 => n25006, A2 => n11676, Z => n11675);
   U19022 : XOR2_X1 port map( A1 => n5890, A2 => n15271, Z => n11682);
   U19024 : XOR2_X1 port map( A1 => n11684, A2 => n15162, Z => n17034);
   U19027 : XOR2_X1 port map( A1 => n5904, A2 => n11226, Z => n20483);
   U19028 : XOR2_X1 port map( A1 => n5904, A2 => n14620, Z => n20322);
   U19029 : NAND3_X1 port map( A1 => n12177, A2 => n20183, A3 => n13719, ZN => 
                           n11691);
   U19030 : NAND2_X2 port map( A1 => n28326, A2 => n13719, ZN => n20184);
   U19031 : NOR2_X1 port map( A1 => n12149, A2 => n17894, ZN => n11694);
   U19035 : XOR2_X1 port map( A1 => n12382, A2 => n21373, Z => n11701);
   U19036 : NAND2_X1 port map( A1 => n27160, A2 => n27344, ZN => n15128);
   U19038 : NOR2_X1 port map( A1 => n22385, A2 => n11983, ZN => n11705);
   U19039 : XOR2_X1 port map( A1 => n22749, A2 => n11708, Z => n11707);
   U19048 : XOR2_X1 port map( A1 => n11728, A2 => n14587, Z => Ciphertext(140))
                           ;
   U19049 : INV_X1 port map( I => n12599, ZN => n17648);
   U19054 : NAND2_X1 port map( A1 => n11743, A2 => n21397, ZN => n12651);
   U19057 : XOR2_X1 port map( A1 => n11752, A2 => n11753, Z => n15557);
   U19058 : XOR2_X1 port map( A1 => n15088, A2 => n20348, Z => n11753);
   U19059 : NAND2_X1 port map( A1 => n24179, A2 => n11756, ZN => n11757);
   U19060 : XOR2_X1 port map( A1 => n27352, A2 => n20989, Z => n19172);
   U19061 : XOR2_X1 port map( A1 => n16918, A2 => n14590, Z => n11769);
   U19064 : XOR2_X1 port map( A1 => n11780, A2 => n16798, Z => n16799);
   U19067 : AOI21_X1 port map( A1 => n13597, A2 => n23575, B => n19124, ZN => 
                           n13596);
   U19069 : NAND2_X1 port map( A1 => n15623, A2 => n12699, ZN => n12724);
   U19070 : INV_X2 port map( I => n11795, ZN => n21578);
   U19071 : XNOR2_X1 port map( A1 => n11799, A2 => n11796, ZN => n11795);
   U19072 : XOR2_X1 port map( A1 => n11798, A2 => n11797, Z => n11796);
   U19073 : XOR2_X1 port map( A1 => n22788, A2 => n12816, Z => n11797);
   U19074 : XOR2_X1 port map( A1 => n20434, A2 => n12925, Z => n11798);
   U19075 : XOR2_X1 port map( A1 => n21238, A2 => n10755, Z => n11799);
   U19085 : INV_X2 port map( I => n11835, ZN => n15686);
   U19086 : XOR2_X1 port map( A1 => n6123, A2 => n13164, Z => n12135);
   U19087 : NOR2_X1 port map( A1 => n22783, A2 => n25342, ZN => n14939);
   U19089 : XOR2_X1 port map( A1 => n14675, A2 => n10612, Z => n11838);
   U19093 : XOR2_X1 port map( A1 => n11845, A2 => n11843, Z => n17137);
   U19094 : INV_X2 port map( I => n11852, ZN => n17301);
   U19096 : INV_X2 port map( I => n17137, ZN => n11857);
   U19100 : OAI21_X1 port map( A1 => n11622, A2 => n21481, B => n24213, ZN => 
                           n21479);
   U19101 : XOR2_X1 port map( A1 => n6867, A2 => n20871, Z => n11866);
   U19102 : NOR2_X1 port map( A1 => n22753, A2 => n27468, ZN => n20874);
   U19104 : AOI22_X1 port map( A1 => n17797, A2 => n8070, B1 => n7985, B2 => 
                           n9772, ZN => n17675);
   U19105 : XOR2_X1 port map( A1 => n12742, A2 => n25946, Z => n13497);
   U19106 : OAI21_X1 port map( A1 => n17953, A2 => n17757, B => n22834, ZN => 
                           n17758);
   U19109 : XOR2_X1 port map( A1 => n18326, A2 => n11887, Z => n11886);
   U19111 : XOR2_X1 port map( A1 => n11898, A2 => n11897, Z => n11896);
   U19112 : XOR2_X1 port map( A1 => n20550, A2 => n20433, Z => n11897);
   U19114 : INV_X1 port map( I => n20558, ZN => n11904);
   U19115 : XOR2_X1 port map( A1 => n11912, A2 => n14564, Z => Ciphertext(113))
                           ;
   U19121 : XOR2_X1 port map( A1 => n11935, A2 => n11934, Z => n11933);
   U19122 : XOR2_X1 port map( A1 => n16941, A2 => n1317, Z => n11934);
   U19124 : AOI21_X1 port map( A1 => n4604, A2 => n20963, B => n705, ZN => 
                           n20958);
   U19125 : XOR2_X1 port map( A1 => n2462, A2 => n4793, Z => n13118);
   U19128 : OAI21_X1 port map( A1 => n12941, A2 => n11369, B => n19914, ZN => 
                           n11950);
   U19129 : MUX2_X1 port map( I0 => n11955, I1 => n11954, S => n13301, Z => 
                           n11953);
   U19132 : XOR2_X1 port map( A1 => n13803, A2 => n20768, Z => n11965);
   U19134 : XOR2_X1 port map( A1 => n18077, A2 => n18113, Z => n11970);
   U19135 : XOR2_X1 port map( A1 => n14659, A2 => n11975, Z => n11974);
   U19141 : NOR2_X2 port map( A1 => n11986, A2 => n11985, ZN => n19989);
   U19142 : XOR2_X1 port map( A1 => n11990, A2 => n18897, Z => n11989);
   U19144 : XOR2_X1 port map( A1 => n19285, A2 => n14624, Z => n11995);
   U19146 : MUX2_X1 port map( I0 => n15864, I1 => n121, S => n12010, Z => 
                           n15867);
   U19147 : INV_X2 port map( I => n15989, ZN => n12010);
   U19149 : XOR2_X1 port map( A1 => Plaintext(36), A2 => Key(36), Z => n12059);
   U19150 : XOR2_X1 port map( A1 => n14608, A2 => n1286, Z => n12015);
   U19157 : OAI21_X1 port map( A1 => n16083, A2 => n12035, B => n16082, ZN => 
                           n14710);
   U19158 : XOR2_X1 port map( A1 => n18058, A2 => n12037, Z => n12036);
   U19160 : XOR2_X1 port map( A1 => n6108, A2 => n18243, Z => n17967);
   U19161 : XNOR2_X1 port map( A1 => n12041, A2 => n13493, ZN => n12040);
   U19162 : XOR2_X1 port map( A1 => n16977, A2 => n10772, Z => n12041);
   U19168 : INV_X2 port map( I => n12059, ZN => n14520);
   U19169 : INV_X1 port map( I => n21055, ZN => n12067);
   U19172 : XOR2_X1 port map( A1 => n4966, A2 => n21313, Z => n12069);
   U19174 : INV_X1 port map( I => n19234, ZN => n19402);
   U19175 : XOR2_X1 port map( A1 => n12072, A2 => n1064, Z => Ciphertext(81));
   U19183 : XOR2_X1 port map( A1 => n13916, A2 => n24000, Z => n12089);
   U19186 : XOR2_X1 port map( A1 => n18272, A2 => n18207, Z => n12093);
   U19187 : INV_X2 port map( I => n24978, ZN => n21328);
   U19190 : XOR2_X1 port map( A1 => Plaintext(78), A2 => Key(78), Z => n12125);
   U19192 : XOR2_X1 port map( A1 => n12110, A2 => n12109, Z => n12108);
   U19193 : XOR2_X1 port map( A1 => n7302, A2 => n22673, Z => n12109);
   U19195 : NAND2_X1 port map( A1 => n12112, A2 => n12234, ZN => n12888);
   U19197 : XOR2_X1 port map( A1 => n15038, A2 => n7431, Z => n12120);
   U19198 : XOR2_X1 port map( A1 => n17116, A2 => n21199, Z => n12122);
   U19200 : NAND2_X1 port map( A1 => n14975, A2 => n20195, ZN => n12130);
   U19201 : NAND2_X1 port map( A1 => n19958, A2 => n860, ZN => n12131);
   U19202 : XOR2_X1 port map( A1 => n7302, A2 => n20702, Z => n19408);
   U19206 : XOR2_X1 port map( A1 => n18208, A2 => n13165, Z => n12136);
   U19212 : INV_X1 port map( I => n13573, ZN => n19129);
   U19214 : AND2_X1 port map( A1 => n17906, A2 => n25724, Z => n12170);
   U19217 : NAND2_X1 port map( A1 => n12179, A2 => n928, ZN => n20988);
   U19218 : AOI22_X2 port map( A1 => n20247, A2 => n20246, B1 => n20248, B2 => 
                           n20249, ZN => n20423);
   U19221 : XOR2_X1 port map( A1 => n24357, A2 => n14587, Z => n13150);
   U19223 : XOR2_X1 port map( A1 => n24357, A2 => n9250, Z => n18149);
   U19226 : XOR2_X1 port map( A1 => n12209, A2 => n20961, Z => n19256);
   U19228 : XOR2_X1 port map( A1 => n28517, A2 => n21216, Z => n16805);
   U19229 : XOR2_X1 port map( A1 => n28517, A2 => n16938, Z => n15097);
   U19231 : XOR2_X1 port map( A1 => n22820, A2 => n21434, Z => n14372);
   U19232 : NAND2_X2 port map( A1 => n15163, A2 => n20083, ZN => n21434);
   U19233 : NAND2_X2 port map( A1 => n13046, A2 => n13045, ZN => n19490);
   U19236 : XOR2_X1 port map( A1 => n12230, A2 => n21227, Z => n15253);
   U19237 : XOR2_X1 port map( A1 => n12230, A2 => n1275, Z => n13332);
   U19238 : XOR2_X1 port map( A1 => n7280, A2 => n12230, Z => n13008);
   U19240 : XOR2_X1 port map( A1 => n2873, A2 => n18068, Z => n12233);
   U19241 : NAND2_X1 port map( A1 => n25324, A2 => n12235, ZN => n13373);
   U19243 : MUX2_X1 port map( I0 => n20685, I1 => n12235, S => n10534, Z => 
                           n20673);
   U19245 : XOR2_X1 port map( A1 => n17013, A2 => n21141, Z => n12249);
   U19246 : NOR2_X1 port map( A1 => n12254, A2 => n21208, ZN => n12253);
   U19247 : XOR2_X1 port map( A1 => n12246, A2 => n20519, Z => n12957);
   U19248 : XOR2_X1 port map( A1 => n12246, A2 => n20989, Z => n20106);
   U19250 : XOR2_X1 port map( A1 => n15817, A2 => Key(77), Z => n16012);
   U19251 : NAND2_X1 port map( A1 => n20323, A2 => n8299, ZN => n19960);
   U19252 : XOR2_X1 port map( A1 => n12278, A2 => n10747, Z => n12277);
   U19254 : XOR2_X1 port map( A1 => n12283, A2 => n12282, Z => n12281);
   U19255 : XOR2_X1 port map( A1 => n19562, A2 => n14573, Z => n12282);
   U19256 : XOR2_X1 port map( A1 => n13852, A2 => n26793, Z => n12291);
   U19258 : INV_X1 port map( I => n16881, ZN => n12285);
   U19261 : XOR2_X1 port map( A1 => n12410, A2 => n22890, Z => n12293);
   U19262 : INV_X1 port map( I => n13790, ZN => n14902);
   U19264 : XOR2_X1 port map( A1 => n18106, A2 => n11181, Z => n12300);
   U19265 : NAND2_X2 port map( A1 => n12306, A2 => n12304, ZN => n19045);
   U19266 : NAND2_X1 port map( A1 => n18620, A2 => n28542, ZN => n12305);
   U19269 : INV_X1 port map( I => n12314, ZN => n20472);
   U19271 : XOR2_X1 port map( A1 => n21198, A2 => n21288, Z => n12316);
   U19274 : XOR2_X1 port map( A1 => n28058, A2 => n20872, Z => n12322);
   U19278 : XOR2_X1 port map( A1 => n8293, A2 => n21649, Z => n14368);
   U19281 : NAND2_X1 port map( A1 => n21539, A2 => n21667, ZN => n12352);
   U19282 : XOR2_X1 port map( A1 => n8912, A2 => n20807, Z => n12354);
   U19284 : XOR2_X1 port map( A1 => n10535, A2 => n14506, Z => n12363);
   U19286 : XOR2_X1 port map( A1 => n12365, A2 => n21613, Z => n12733);
   U19287 : XOR2_X1 port map( A1 => n12365, A2 => n21436, Z => n13589);
   U19288 : XOR2_X1 port map( A1 => n9678, A2 => n12365, Z => n14978);
   U19290 : XOR2_X1 port map( A1 => n27378, A2 => n12365, Z => n13189);
   U19292 : XOR2_X1 port map( A1 => n17131, A2 => n12381, Z => n12380);
   U19293 : XOR2_X1 port map( A1 => n17133, A2 => n14604, Z => n12381);
   U19295 : XOR2_X1 port map( A1 => n25332, A2 => n24682, Z => n15691);
   U19297 : INV_X2 port map( I => n12396, ZN => n13049);
   U19304 : XOR2_X1 port map( A1 => n24197, A2 => n1277, Z => n12405);
   U19307 : XOR2_X1 port map( A1 => n17156, A2 => n17155, Z => n13320);
   U19308 : OAI21_X1 port map( A1 => n13622, A2 => n22766, B => n13085, ZN => 
                           n13084);
   U19309 : XOR2_X1 port map( A1 => n24094, A2 => n7011, Z => n21189);
   U19312 : XOR2_X1 port map( A1 => n18283, A2 => n13464, Z => n12414);
   U19314 : NAND2_X1 port map( A1 => n12417, A2 => n25325, ZN => n12416);
   U19319 : MUX2_X1 port map( I0 => n11870, I1 => n22835, S => n3525, Z => 
                           n12830);
   U19320 : NOR2_X1 port map( A1 => n13475, A2 => n15709, ZN => n13023);
   U19326 : XOR2_X1 port map( A1 => n22792, A2 => n20713, Z => n12437);
   U19331 : INV_X1 port map( I => n18013, ZN => n14066);
   U19333 : NAND3_X1 port map( A1 => n12446, A2 => n15498, A3 => n15499, ZN => 
                           n21655);
   U19334 : NAND2_X1 port map( A1 => n13349, A2 => n23017, ZN => n12451);
   U19337 : XOR2_X1 port map( A1 => n17088, A2 => n14123, Z => n12454);
   U19340 : XOR2_X1 port map( A1 => n14227, A2 => n22806, Z => n12457);
   U19341 : XOR2_X1 port map( A1 => n15161, A2 => n12458, Z => n19692);
   U19342 : XOR2_X1 port map( A1 => n15691, A2 => n19514, Z => n12458);
   U19346 : NAND2_X1 port map( A1 => n14926, A2 => n12493, ZN => n12721);
   U19347 : INV_X1 port map( I => n12930, ZN => n17985);
   U19351 : XOR2_X1 port map( A1 => n17100, A2 => n17101, Z => n17104);
   U19358 : OAI21_X1 port map( A1 => n18912, A2 => n25367, B => n14201, ZN => 
                           n18869);
   U19371 : NAND2_X1 port map( A1 => n20836, A2 => n13057, ZN => n13073);
   U19372 : NAND2_X1 port map( A1 => n20992, A2 => n26712, ZN => n20995);
   U19375 : NOR2_X1 port map( A1 => n15179, A2 => n5558, ZN => n15649);
   U19376 : NAND2_X1 port map( A1 => n11382, A2 => n15674, ZN => n12989);
   U19378 : XOR2_X1 port map( A1 => n13695, A2 => n13773, Z => n12515);
   U19379 : XOR2_X1 port map( A1 => n6309, A2 => n19489, Z => n18938);
   U19380 : XOR2_X1 port map( A1 => n20458, A2 => n21033, Z => n20354);
   U19381 : XOR2_X1 port map( A1 => Plaintext(156), A2 => Key(156), Z => n12534
                           );
   U19383 : XOR2_X1 port map( A1 => n13458, A2 => n13459, Z => n12522);
   U19387 : XOR2_X1 port map( A1 => Plaintext(1), A2 => Key(1), Z => n12529);
   U19391 : INV_X2 port map( I => n12534, ZN => n16273);
   U19392 : NAND2_X1 port map( A1 => n12542, A2 => n19101, ZN => n19203);
   U19399 : XOR2_X1 port map( A1 => n17131, A2 => n12565, Z => n12564);
   U19400 : XOR2_X1 port map( A1 => n16910, A2 => n14573, Z => n12565);
   U19402 : XOR2_X1 port map( A1 => n22879, A2 => n15506, Z => n18193);
   U19403 : XOR2_X1 port map( A1 => n12572, A2 => n18081, Z => n18024);
   U19404 : XOR2_X1 port map( A1 => n13299, A2 => n12202, Z => n12574);
   U19409 : XOR2_X1 port map( A1 => n18088, A2 => n18236, Z => n12602);
   U19410 : OAI21_X1 port map( A1 => n27454, A2 => n27679, B => n12603, ZN => 
                           n20039);
   U19414 : XOR2_X1 port map( A1 => n7302, A2 => n14473, Z => n19282);
   U19416 : XOR2_X1 port map( A1 => n2508, A2 => n21454, Z => n12906);
   U19417 : XOR2_X1 port map( A1 => n22768, A2 => n20707, Z => n12623);
   U19418 : NOR2_X1 port map( A1 => n12625, A2 => n21529, ZN => n21520);
   U19419 : AOI21_X1 port map( A1 => n21528, A2 => n12625, B => n21530, ZN => 
                           n21532);
   U19420 : XOR2_X1 port map( A1 => n452, A2 => n14432, Z => n16982);
   U19422 : NOR2_X1 port map( A1 => n20151, A2 => n20338, ZN => n12631);
   U19424 : NAND2_X1 port map( A1 => n14059, A2 => n12643, ZN => n20127);
   U19426 : XOR2_X1 port map( A1 => n12646, A2 => n12645, Z => n13296);
   U19427 : XOR2_X1 port map( A1 => n15604, A2 => n25980, Z => n12645);
   U19428 : NAND2_X1 port map( A1 => n7539, A2 => n12647, ZN => n16603);
   U19429 : NAND2_X2 port map( A1 => n12652, A2 => n12651, ZN => n21413);
   U19430 : INV_X1 port map( I => n14679, ZN => n12654);
   U19431 : INV_X2 port map( I => n12655, ZN => n13693);
   U19433 : NAND2_X1 port map( A1 => n15199, A2 => n27412, ZN => n15198);
   U19438 : INV_X2 port map( I => n13679, ZN => n14343);
   U19440 : XOR2_X1 port map( A1 => n10529, A2 => n21090, Z => n13959);
   U19441 : XOR2_X1 port map( A1 => n27348, A2 => n10529, Z => n15385);
   U19443 : OR2_X1 port map( A1 => n24550, A2 => n16565, Z => n12700);
   U19446 : XOR2_X1 port map( A1 => n18269, A2 => n12715, Z => n12714);
   U19447 : XOR2_X1 port map( A1 => n22829, A2 => n27589, Z => n12715);
   U19449 : XOR2_X1 port map( A1 => n13354, A2 => n19512, Z => n12717);
   U19451 : NAND2_X1 port map( A1 => n17390, A2 => n15504, ZN => n12719);
   U19453 : NAND2_X1 port map( A1 => n17386, A2 => n24368, ZN => n14253);
   U19454 : XOR2_X1 port map( A1 => n14743, A2 => n4876, Z => n16439);
   U19455 : INV_X1 port map( I => n12732, ZN => n18711);
   U19465 : XOR2_X1 port map( A1 => n28407, A2 => n21419, Z => n18122);
   U19466 : XOR2_X1 port map( A1 => n12532, A2 => n11679, Z => n12778);
   U19467 : XOR2_X1 port map( A1 => n12926, A2 => n22778, Z => n12779);
   U19469 : OAI21_X1 port map( A1 => n15345, A2 => n13986, B => n12784, ZN => 
                           n13798);
   U19470 : XOR2_X1 port map( A1 => n12788, A2 => n21454, Z => Ciphertext(136))
                           ;
   U19475 : NAND2_X1 port map( A1 => n21568, A2 => n12797, ZN => n21569);
   U19476 : XOR2_X1 port map( A1 => n28355, A2 => n14573, Z => n12803);
   U19478 : INV_X2 port map( I => n12926, ZN => n12925);
   U19479 : OR2_X1 port map( A1 => n13032, A2 => n21109, Z => n13031);
   U19480 : XOR2_X1 port map( A1 => Plaintext(123), A2 => Key(123), Z => n13420
                           );
   U19481 : NOR2_X1 port map( A1 => n1191, A2 => n18344, ZN => n12821);
   U19482 : XOR2_X1 port map( A1 => n14026, A2 => n12824, Z => n12823);
   U19486 : NAND2_X1 port map( A1 => n7017, A2 => n18005, ZN => n17711);
   U19487 : XOR2_X1 port map( A1 => n18357, A2 => n12854, Z => n12853);
   U19490 : XOR2_X1 port map( A1 => n17139, A2 => n12831, Z => n12857);
   U19491 : XOR2_X1 port map( A1 => n4866, A2 => n20514, Z => n12860);
   U19494 : XOR2_X1 port map( A1 => n25387, A2 => n1309, Z => n12862);
   U19496 : AOI22_X1 port map( A1 => n13533, A2 => n16280, B1 => n16279, B2 => 
                           n11291, ZN => n15941);
   U19503 : NAND2_X1 port map( A1 => n16273, A2 => n8867, ZN => n12874);
   U19505 : NOR2_X1 port map( A1 => n21901, A2 => n17687, ZN => n13730);
   U19509 : XOR2_X1 port map( A1 => n12903, A2 => n12813, Z => Ciphertext(151))
                           ;
   U19511 : XOR2_X1 port map( A1 => n19547, A2 => n12906, Z => n12907);
   U19512 : XOR2_X1 port map( A1 => n19510, A2 => n19312, Z => n19547);
   U19514 : XOR2_X1 port map( A1 => n22792, A2 => n12916, Z => n12915);
   U19515 : INV_X1 port map( I => n14506, ZN => n12916);
   U19516 : XOR2_X1 port map( A1 => n12932, A2 => n17671, Z => n17672);
   U19519 : XOR2_X1 port map( A1 => n36, A2 => n14650, Z => n21251);
   U19521 : XOR2_X1 port map( A1 => n12958, A2 => n12957, Z => n12956);
   U19526 : XOR2_X1 port map( A1 => n21364, A2 => n25642, Z => n21365);
   U19527 : XOR2_X1 port map( A1 => n13092, A2 => n25642, Z => n21429);
   U19528 : XOR2_X1 port map( A1 => n18057, A2 => n18068, Z => n13000);
   U19531 : NOR2_X1 port map( A1 => n829, A2 => n13129, ZN => n17816);
   U19539 : NOR2_X1 port map( A1 => n17227, A2 => n17346, ZN => n13054);
   U19542 : XOR2_X1 port map( A1 => n5529, A2 => n20602, Z => n13077);
   U19543 : XOR2_X1 port map( A1 => n18020, A2 => n13079, Z => n13078);
   U19544 : XOR2_X1 port map( A1 => n25306, A2 => n21784, Z => n13079);
   U19546 : AND2_X1 port map( A1 => n22766, A2 => n20625, Z => n13081);
   U19547 : INV_X1 port map( I => n18392, ZN => n18395);
   U19548 : NOR3_X1 port map( A1 => n13095, A2 => n20804, A3 => n20803, ZN => 
                           n20796);
   U19549 : NAND2_X1 port map( A1 => n20799, A2 => n13095, ZN => n20791);
   U19555 : XOR2_X1 port map( A1 => n26082, A2 => n14610, Z => n16389);
   U19558 : XOR2_X1 port map( A1 => n20763, A2 => n21314, Z => n13114);
   U19559 : XOR2_X1 port map( A1 => n20563, A2 => n15064, Z => n13115);
   U19561 : XOR2_X1 port map( A1 => n19405, A2 => n20396, Z => n13117);
   U19563 : XOR2_X1 port map( A1 => n19406, A2 => n14463, Z => n18831);
   U19564 : XOR2_X1 port map( A1 => n25312, A2 => n13122, Z => n13153);
   U19567 : XOR2_X1 port map( A1 => n13131, A2 => n13134, Z => n13130);
   U19568 : XOR2_X1 port map( A1 => n147, A2 => n16916, Z => n13133);
   U19569 : XOR2_X1 port map( A1 => n13916, A2 => n23021, Z => n13134);
   U19571 : NAND2_X1 port map( A1 => n25415, A2 => n6110, ZN => n13137);
   U19574 : XOR2_X1 port map( A1 => n18066, A2 => n18112, Z => n13151);
   U19575 : XOR2_X1 port map( A1 => n18035, A2 => n13153, Z => n13152);
   U19576 : XOR2_X1 port map( A1 => n14608, A2 => n1281, Z => n13155);
   U19578 : NAND2_X2 port map( A1 => n19030, A2 => n19029, ZN => n19481);
   U19579 : OAI21_X1 port map( A1 => n15469, A2 => n21606, B => n15470, ZN => 
                           n13161);
   U19582 : XOR2_X1 port map( A1 => n446, A2 => n14581, Z => n21316);
   U19584 : INV_X2 port map( I => n13170, ZN => n21702);
   U19585 : NAND2_X1 port map( A1 => n13170, A2 => n773, ZN => n13172);
   U19586 : XOR2_X1 port map( A1 => n22768, A2 => n22837, Z => n15361);
   U19587 : XOR2_X1 port map( A1 => n7130, A2 => n1302, Z => n13178);
   U19588 : XOR2_X1 port map( A1 => n24197, A2 => n4137, Z => n13179);
   U19589 : XOR2_X1 port map( A1 => n21153, A2 => n20511, Z => n21418);
   U19590 : NAND2_X2 port map( A1 => n13340, A2 => n15102, ZN => n18182);
   U19592 : XOR2_X1 port map( A1 => n20410, A2 => n25362, Z => n13190);
   U19596 : OAI21_X1 port map( A1 => n15424, A2 => n14582, B => n12648, ZN => 
                           n15054);
   U19597 : XOR2_X1 port map( A1 => n21305, A2 => n7044, Z => n13195);
   U19601 : XOR2_X1 port map( A1 => n13201, A2 => n20555, Z => n21068);
   U19605 : NAND2_X1 port map( A1 => n7354, A2 => n20979, ZN => n20811);
   U19607 : XOR2_X1 port map( A1 => n17154, A2 => n546, Z => n17155);
   U19608 : XOR2_X1 port map( A1 => n16913, A2 => n16816, Z => n17154);
   U19609 : XOR2_X1 port map( A1 => n18241, A2 => n10907, Z => n13225);
   U19612 : XOR2_X1 port map( A1 => n17839, A2 => n13228, Z => n18642);
   U19613 : XOR2_X1 port map( A1 => n17837, A2 => n17838, Z => n13228);
   U19614 : CLKBUF_X2 port map( I => Key(107), Z => n16961);
   U19615 : NAND2_X1 port map( A1 => n17764, A2 => n1025, ZN => n13238);
   U19616 : XNOR2_X1 port map( A1 => n8879, A2 => n13787, ZN => n13288);
   U19619 : INV_X1 port map( I => n17847, ZN => n14976);
   U19620 : NAND2_X1 port map( A1 => n20869, A2 => n20868, ZN => n14182);
   U19621 : NAND2_X1 port map( A1 => n14190, A2 => n14189, ZN => n15408);
   U19622 : XOR2_X1 port map( A1 => n13300, A2 => n14368, Z => n20460);
   U19626 : NAND2_X1 port map( A1 => n18499, A2 => n22977, ZN => n14206);
   U19628 : NAND2_X2 port map( A1 => n20135, A2 => n13267, ZN => n21116);
   U19630 : XOR2_X1 port map( A1 => n20351, A2 => n10647, Z => n14567);
   U19640 : NOR2_X1 port map( A1 => n15565, A2 => n15909, ZN => n16236);
   U19641 : NAND2_X2 port map( A1 => n13295, A2 => n21322, ZN => n21355);
   U19645 : NOR3_X1 port map( A1 => n24646, A2 => n11908, A3 => n14137, ZN => 
                           n16546);
   U19658 : INV_X2 port map( I => n13337, ZN => n14858);
   U19659 : XOR2_X1 port map( A1 => Plaintext(38), A2 => Key(38), Z => n13337);
   U19663 : INV_X2 port map( I => n13343, ZN => n13613);
   U19664 : XOR2_X1 port map( A1 => Plaintext(15), A2 => Key(15), Z => n13343);
   U19665 : INV_X2 port map( I => n11487, ZN => n20262);
   U19669 : XOR2_X1 port map( A1 => n13348, A2 => n15148, Z => n13433);
   U19670 : NAND2_X1 port map( A1 => n19960, A2 => n26738, ZN => n19961);
   U19672 : XOR2_X1 port map( A1 => n13344, A2 => n16768, Z => n16769);
   U19677 : XOR2_X1 port map( A1 => n13364, A2 => n15253, Z => n13810);
   U19678 : OAI21_X1 port map( A1 => n16704, A2 => n12839, B => n14344, ZN => 
                           n16154);
   U19680 : XOR2_X1 port map( A1 => n13449, A2 => n21554, Z => n13450);
   U19682 : XOR2_X1 port map( A1 => n18264, A2 => n18265, Z => n13370);
   U19683 : AOI21_X1 port map( A1 => n20685, A2 => n13373, B => n28176, ZN => 
                           n20687);
   U19686 : XOR2_X1 port map( A1 => Plaintext(163), A2 => Key(163), Z => n13407
                           );
   U19690 : XOR2_X1 port map( A1 => n982, A2 => n15126, Z => n13938);
   U19691 : NAND2_X1 port map( A1 => n16398, A2 => n16731, ZN => n14246);
   U19695 : NOR2_X2 port map( A1 => n14924, A2 => n14923, ZN => n14926);
   U19703 : XOR2_X1 port map( A1 => n16947, A2 => n13404, Z => n13403);
   U19706 : INV_X2 port map( I => n13407, ZN => n16258);
   U19707 : OR2_X1 port map( A1 => n14908, A2 => n1257, Z => n14865);
   U19708 : NOR2_X1 port map( A1 => n21639, A2 => n15219, ZN => n15218);
   U19709 : XOR2_X1 port map( A1 => n14402, A2 => n19607, Z => n14248);
   U19710 : XOR2_X1 port map( A1 => n20456, A2 => n20455, Z => n13412);
   U19713 : XOR2_X1 port map( A1 => Plaintext(175), A2 => Key(175), Z => n15491
                           );
   U19715 : INV_X1 port map( I => n16902, ZN => n14687);
   U19716 : XOR2_X1 port map( A1 => n13425, A2 => n14469, Z => n19661);
   U19719 : OAI21_X1 port map( A1 => n13977, A2 => n7944, B => n13976, ZN => 
                           n13975);
   U19720 : XOR2_X1 port map( A1 => n13433, A2 => n15138, Z => n15642);
   U19722 : OR2_X1 port map( A1 => n4428, A2 => n21116, Z => n13436);
   U19725 : NAND2_X1 port map( A1 => n24951, A2 => n13444, ZN => n13474);
   U19728 : XOR2_X1 port map( A1 => n25313, A2 => n21679, Z => n13459);
   U19729 : XOR2_X1 port map( A1 => n14962, A2 => n13579, Z => n13466);
   U19730 : XOR2_X1 port map( A1 => n13466, A2 => n13580, Z => n19472);
   U19731 : XOR2_X1 port map( A1 => n13470, A2 => n14463, Z => Ciphertext(99));
   U19732 : INV_X2 port map( I => n13475, ZN => n13600);
   U19734 : MUX2_X1 port map( I0 => n25224, I1 => n21873, S => n13435, Z => 
                           n15890);
   U19737 : INV_X2 port map( I => n13507, ZN => n20732);
   U19739 : XOR2_X1 port map( A1 => n13856, A2 => n16905, Z => n13510);
   U19740 : XOR2_X1 port map( A1 => n17123, A2 => n17034, Z => n13511);
   U19741 : MUX2_X1 port map( I0 => n16383, I1 => n16381, S => n10261, Z => 
                           n16385);
   U19744 : XOR2_X1 port map( A1 => n13524, A2 => n21367, Z => n16870);
   U19745 : MUX2_X1 port map( I0 => n18003, I1 => n18002, S => n13530, Z => 
                           n18004);
   U19748 : NAND2_X2 port map( A1 => n16098, A2 => n16097, ZN => n14632);
   U19749 : XOR2_X1 port map( A1 => n27969, A2 => n27243, Z => n16835);
   U19750 : XOR2_X1 port map( A1 => n17147, A2 => n27848, Z => n17148);
   U19752 : INV_X2 port map( I => n26702, ZN => n16196);
   U19753 : XOR2_X1 port map( A1 => n15843, A2 => Key(95), Z => n16306);
   U19758 : XOR2_X1 port map( A1 => n13561, A2 => n13560, Z => n19755);
   U19759 : XOR2_X1 port map( A1 => n19343, A2 => n19178, Z => n13560);
   U19760 : NAND2_X1 port map( A1 => n14763, A2 => n13562, ZN => n14787);
   U19763 : OR3_X1 port map( A1 => n18600, A2 => n18599, A3 => n18602, Z => 
                           n15132);
   U19767 : XOR2_X1 port map( A1 => n21434, A2 => n21435, Z => n13590);
   U19769 : NAND2_X1 port map( A1 => n12465, A2 => n15724, ZN => n20810);
   U19774 : INV_X1 port map( I => n13622, ZN => n20619);
   U19775 : NOR3_X1 port map( A1 => n21618, A2 => n27023, A3 => n26435, ZN => 
                           n13625);
   U19776 : XOR2_X1 port map( A1 => n17083, A2 => n13632, Z => n13631);
   U19777 : XOR2_X1 port map( A1 => n17084, A2 => n17085, Z => n13632);
   U19778 : NAND2_X1 port map( A1 => n15209, A2 => n22421, ZN => n21205);
   U19780 : XOR2_X1 port map( A1 => n13644, A2 => n23156, Z => n13643);
   U19781 : XOR2_X1 port map( A1 => n14144, A2 => n21247, Z => n13644);
   U19783 : XOR2_X1 port map( A1 => n15081, A2 => n13647, Z => n18410);
   U19784 : XOR2_X1 port map( A1 => Plaintext(182), A2 => Key(182), Z => n14515
                           );
   U19786 : XOR2_X1 port map( A1 => n18120, A2 => n13676, Z => n13832);
   U19788 : MUX2_X1 port map( I0 => n16148, I1 => n13677, S => n15960, Z => 
                           n15961);
   U19790 : OR2_X2 port map( A1 => n16458, A2 => n16459, Z => n15708);
   U19794 : XOR2_X1 port map( A1 => n13702, A2 => n13699, Z => n21502);
   U19795 : XOR2_X1 port map( A1 => n13701, A2 => n13700, Z => n13699);
   U19796 : XOR2_X1 port map( A1 => n21257, A2 => n14556, Z => n13700);
   U19797 : XOR2_X1 port map( A1 => n21255, A2 => n21254, Z => n13701);
   U19802 : XOR2_X1 port map( A1 => n21651, A2 => n22749, Z => n13711);
   U19806 : NOR2_X1 port map( A1 => n13717, A2 => n16144, ZN => n15826);
   U19809 : XOR2_X1 port map( A1 => Plaintext(69), A2 => Key(69), Z => n15525);
   U19810 : NOR2_X1 port map( A1 => n13545, A2 => n730, ZN => n16309);
   U19813 : NOR2_X1 port map( A1 => n13565, A2 => n17871, ZN => n13735);
   U19814 : XOR2_X1 port map( A1 => n18087, A2 => n13737, Z => n14856);
   U19815 : NOR2_X1 port map( A1 => n22794, A2 => n13741, ZN => n13743);
   U19818 : XOR2_X1 port map( A1 => n14980, A2 => n28148, Z => n13747);
   U19819 : XOR2_X1 port map( A1 => n25337, A2 => n16938, Z => n13749);
   U19820 : XOR2_X1 port map( A1 => n21365, A2 => n13751, Z => n13750);
   U19821 : XOR2_X1 port map( A1 => n15226, A2 => n21363, Z => n13751);
   U19822 : NAND3_X1 port map( A1 => n27569, A2 => n1163, A3 => n19190, ZN => 
                           n18618);
   U19828 : OR2_X1 port map( A1 => n20223, A2 => n23374, Z => n13762);
   U19829 : NAND2_X1 port map( A1 => n14017, A2 => n13772, ZN => n14873);
   U19830 : XOR2_X1 port map( A1 => n14570, A2 => n19338, Z => n13773);
   U19832 : XOR2_X1 port map( A1 => n22760, A2 => n6540, Z => n13777);
   U19833 : XOR2_X1 port map( A1 => n19538, A2 => n13785, Z => n13784);
   U19835 : XOR2_X1 port map( A1 => Plaintext(137), A2 => Key(137), Z => n14224
                           );
   U19836 : XOR2_X1 port map( A1 => n21187, A2 => n21302, Z => n15477);
   U19840 : XOR2_X1 port map( A1 => n21153, A2 => n7365, Z => n13802);
   U19850 : XOR2_X1 port map( A1 => n13832, A2 => n18183, Z => n15694);
   U19851 : INV_X2 port map( I => n13833, ZN => n16123);
   U19852 : XNOR2_X1 port map( A1 => Plaintext(50), A2 => Key(50), ZN => n13833
                           );
   U19857 : INV_X1 port map( I => n15604, ZN => n18057);
   U19858 : XOR2_X1 port map( A1 => n18262, A2 => n13859, Z => n13858);
   U19860 : INV_X2 port map( I => n13863, ZN => n14193);
   U19861 : XOR2_X1 port map( A1 => n22756, A2 => n21683, Z => n20055);
   U19865 : OAI21_X1 port map( A1 => n13888, A2 => n21290, B => n21279, ZN => 
                           n21282);
   U19868 : XOR2_X1 port map( A1 => n14699, A2 => n446, Z => n13892);
   U19870 : XOR2_X1 port map( A1 => n8150, A2 => n10680, Z => n13894);
   U19871 : INV_X2 port map( I => n13896, ZN => n14424);
   U19873 : NAND2_X1 port map( A1 => n15401, A2 => n17421, ZN => n13903);
   U19874 : NAND2_X1 port map( A1 => n20901, A2 => n25629, ZN => n20902);
   U19876 : NOR2_X2 port map( A1 => n14304, A2 => n26623, ZN => n14752);
   U19877 : OR3_X1 port map( A1 => n21605, A2 => n15475, A3 => n21603, Z => 
                           n13921);
   U19878 : XOR2_X1 port map( A1 => n19376, A2 => n13923, Z => n14758);
   U19879 : XOR2_X1 port map( A1 => n12739, A2 => n21010, Z => n13923);
   U19881 : NAND2_X1 port map( A1 => n16513, A2 => n14320, ZN => n14483);
   U19882 : XOR2_X1 port map( A1 => n13929, A2 => n1286, Z => Ciphertext(135));
   U19883 : XOR2_X1 port map( A1 => n22847, A2 => n19316, Z => n13930);
   U19885 : XOR2_X1 port map( A1 => n24312, A2 => n14614, Z => n13936);
   U19887 : NOR2_X1 port map( A1 => n8049, A2 => n27813, ZN => n13983);
   U19888 : XOR2_X1 port map( A1 => n16875, A2 => n15162, Z => n13945);
   U19889 : XOR2_X1 port map( A1 => n18313, A2 => n13959, Z => n13958);
   U19890 : XOR2_X1 port map( A1 => n13342, A2 => n21191, Z => n15723);
   U19891 : XOR2_X1 port map( A1 => n9678, A2 => n21258, Z => n13965);
   U19892 : AOI22_X1 port map( A1 => n15345, A2 => n12508, B1 => n13986, B2 => 
                           n21455, ZN => n13977);
   U19893 : XOR2_X1 port map( A1 => n27371, A2 => n14540, Z => n13971);
   U19894 : XOR2_X1 port map( A1 => n13975, A2 => n21450, Z => Ciphertext(134))
                           ;
   U19896 : XOR2_X1 port map( A1 => n14006, A2 => n20727, Z => n16750);
   U19897 : XOR2_X1 port map( A1 => n14006, A2 => n14007, Z => n15466);
   U19898 : XOR2_X1 port map( A1 => n13996, A2 => n698, Z => n18261);
   U19899 : XOR2_X1 port map( A1 => n13999, A2 => n13998, Z => n16722);
   U19900 : XOR2_X1 port map( A1 => n14000, A2 => n16666, Z => n13998);
   U19901 : XOR2_X1 port map( A1 => n14023, A2 => n17108, Z => n13999);
   U19902 : XOR2_X1 port map( A1 => n14002, A2 => n19271, Z => n14001);
   U19905 : XOR2_X1 port map( A1 => n14011, A2 => n14010, Z => n14009);
   U19906 : XOR2_X1 port map( A1 => n19305, A2 => n15503, Z => n14010);
   U19907 : NAND2_X1 port map( A1 => n21645, A2 => n932, ZN => n15427);
   U19909 : XOR2_X1 port map( A1 => n17088, A2 => n26132, Z => n14014);
   U19910 : XOR2_X1 port map( A1 => n17087, A2 => n17089, Z => n14015);
   U19911 : XOR2_X1 port map( A1 => n19512, A2 => n21143, Z => n14021);
   U19913 : NAND2_X1 port map( A1 => n21279, A2 => n21292, ZN => n14024);
   U19916 : NAND2_X1 port map( A1 => n19942, A2 => n3226, ZN => n14044);
   U19919 : XOR2_X1 port map( A1 => n28292, A2 => n14526, Z => n14047);
   U19920 : XOR2_X1 port map( A1 => n18330, A2 => n18237, Z => n14048);
   U19925 : XOR2_X1 port map( A1 => n24384, A2 => n15271, Z => n18518);
   U19928 : XOR2_X1 port map( A1 => n17142, A2 => n14581, Z => n14073);
   U19930 : NAND2_X1 port map( A1 => n21353, A2 => n21342, ZN => n14078);
   U19931 : AOI21_X2 port map( A1 => n21331, A2 => n15463, B => n21330, ZN => 
                           n21347);
   U19935 : XOR2_X1 port map( A1 => n7244, A2 => n21449, Z => n18338);
   U19936 : INV_X2 port map( I => n14094, ZN => n20897);
   U19938 : BUF_X2 port map( I => n21502, Z => n14525);
   U19939 : AOI21_X1 port map( A1 => n21516, A2 => n21529, B => n21515, ZN => 
                           n14268);
   U19940 : NAND2_X1 port map( A1 => n15607, A2 => n15565, ZN => n15803);
   U19941 : XOR2_X1 port map( A1 => n14105, A2 => n14266, Z => n19329);
   U19942 : BUF_X2 port map( I => n16331, Z => n14107);
   U19943 : OR2_X1 port map( A1 => n7985, A2 => n14255, Z => n14110);
   U19944 : XNOR2_X1 port map( A1 => n18223, A2 => n18222, ZN => n14208);
   U19945 : INV_X1 port map( I => n17800, ZN => n14114);
   U19948 : INV_X1 port map( I => n14311, ZN => n16330);
   U19952 : INV_X2 port map( I => n14132, ZN => n17353);
   U19953 : NAND2_X1 port map( A1 => n12206, A2 => n25418, ZN => n14134);
   U19954 : XOR2_X1 port map( A1 => Plaintext(41), A2 => Key(41), Z => n14174);
   U19956 : XOR2_X1 port map( A1 => n14136, A2 => n21216, Z => Ciphertext(109))
                           ;
   U19958 : OAI22_X1 port map( A1 => n21514, A2 => n27389, B1 => n21525, B2 => 
                           n21536, ZN => n21515);
   U19960 : XOR2_X1 port map( A1 => n14151, A2 => n10715, Z => n14685);
   U19966 : NAND2_X1 port map( A1 => n20141, A2 => n20082, ZN => n20083);
   U19972 : AOI22_X1 port map( A1 => n15554, A2 => n721, B1 => n15553, B2 => 
                           n21682, ZN => n15552);
   U19983 : NOR2_X1 port map( A1 => n5434, A2 => n18377, ZN => n18378);
   U19986 : INV_X2 port map( I => n14202, ZN => n15025);
   U19987 : XOR2_X1 port map( A1 => n15856, A2 => Key(99), Z => n14202);
   U19988 : XOR2_X1 port map( A1 => n18224, A2 => n14208, Z => n14383);
   U19991 : OAI21_X1 port map( A1 => n21680, A2 => n10576, B => n15552, ZN => 
                           n15551);
   U19993 : NAND2_X1 port map( A1 => n16035, A2 => n719, ZN => n14214);
   U19995 : INV_X2 port map( I => n14220, ZN => n15565);
   U19996 : XOR2_X1 port map( A1 => Plaintext(165), A2 => Key(165), Z => n14220
                           );
   U19998 : INV_X1 port map( I => n20219, ZN => n14235);
   U19999 : XOR2_X1 port map( A1 => Plaintext(169), A2 => Key(169), Z => n14655
                           );
   U20004 : INV_X1 port map( I => n16475, ZN => n15528);
   U20007 : NAND2_X1 port map( A1 => n13371, A2 => n19134, ZN => n19136);
   U20009 : XNOR2_X1 port map( A1 => n27366, A2 => n21210, ZN => n15064);
   U20010 : XOR2_X1 port map( A1 => n16819, A2 => n15506, Z => n16855);
   U20012 : XOR2_X1 port map( A1 => Plaintext(134), A2 => Key(134), Z => n15354
                           );
   U20014 : XOR2_X1 port map( A1 => n14268, A2 => n21517, Z => Ciphertext(144))
                           ;
   U20017 : XOR2_X1 port map( A1 => n19059, A2 => n19058, Z => n19067);
   U20019 : INV_X1 port map( I => n21529, ZN => n21526);
   U20020 : XOR2_X1 port map( A1 => n23186, A2 => n18337, Z => n14956);
   U20021 : NAND2_X1 port map( A1 => n22581, A2 => n2023, ZN => n14292);
   U20024 : INV_X2 port map( I => n14305, ZN => n15209);
   U20025 : XOR2_X1 port map( A1 => n20062, A2 => n20061, Z => n14305);
   U20032 : XOR2_X1 port map( A1 => Plaintext(135), A2 => Key(135), Z => n14425
                           );
   U20036 : XOR2_X1 port map( A1 => Plaintext(116), A2 => Key(116), Z => n14814
                           );
   U20043 : XOR2_X1 port map( A1 => Plaintext(160), A2 => Key(160), Z => n16107
                           );
   U20045 : NAND2_X1 port map( A1 => n18643, A2 => n24701, ZN => n14375);
   U20048 : INV_X2 port map( I => n14383, ZN => n18466);
   U20052 : AND2_X1 port map( A1 => n21058, A2 => n28139, Z => n20560);
   U20053 : XOR2_X1 port map( A1 => n10705, A2 => n17086, Z => n16867);
   U20054 : XOR2_X1 port map( A1 => n28222, A2 => n21523, Z => n14402);
   U20058 : INV_X2 port map( I => n14416, ZN => n20894);
   U20062 : NAND2_X1 port map( A1 => n10001, A2 => n16271, ZN => n14434);
   U20063 : XNOR2_X1 port map( A1 => n22788, A2 => n21147, ZN => n15356);
   U20065 : NOR2_X1 port map( A1 => n15236, A2 => n15235, ZN => n15988);
   U20067 : INV_X1 port map( I => n21347, ZN => n21352);
   U20068 : XOR2_X1 port map( A1 => n20106, A2 => n20548, Z => n14455);
   U20069 : NAND2_X1 port map( A1 => n14401, A2 => n27372, ZN => n14969);
   U20072 : NAND2_X1 port map( A1 => n20948, A2 => n23088, ZN => n14465);
   U20076 : NAND2_X1 port map( A1 => n18643, A2 => n18747, ZN => n14484);
   U20078 : XOR2_X1 port map( A1 => n17828, A2 => n14487, Z => n18569);
   U20079 : XOR2_X1 port map( A1 => n18114, A2 => n17827, Z => n14487);
   U20081 : INV_X1 port map( I => n12431, ZN => n19625);
   U20082 : XOR2_X1 port map( A1 => n14495, A2 => n14758, Z => n14757);
   U20083 : XOR2_X1 port map( A1 => n25098, A2 => n20433, Z => n14496);
   U20089 : INV_X2 port map( I => n14515, ZN => n16266);
   U20091 : XNOR2_X1 port map( A1 => n21195, A2 => n21194, ZN => n14529);
   U20092 : XOR2_X1 port map( A1 => n16968, A2 => n16967, Z => n17003);
   U20094 : XOR2_X1 port map( A1 => n14534, A2 => n15340, Z => n21323);
   U20095 : XOR2_X1 port map( A1 => n21187, A2 => n21186, Z => n14534);
   U20096 : XOR2_X1 port map( A1 => n19310, A2 => n19292, Z => n19296);
   U20098 : XOR2_X1 port map( A1 => n28269, A2 => n21170, Z => n18333);
   U20099 : XOR2_X1 port map( A1 => n16734, A2 => n16735, Z => n16742);
   U20103 : XOR2_X1 port map( A1 => n28483, A2 => n20919, Z => n20724);
   U20105 : OR2_X1 port map( A1 => n14364, A2 => n16728, Z => n16475);
   U20107 : OR2_X1 port map( A1 => n21780, A2 => n24209, Z => n15291);
   U20108 : XOR2_X1 port map( A1 => n14605, A2 => n20851, Z => Ciphertext(47));
   U20111 : AND2_X1 port map( A1 => n15873, A2 => n14636, Z => n14635);
   U20112 : INV_X2 port map( I => n21016, ZN => n21096);
   U20113 : INV_X2 port map( I => n14655, ZN => n16088);
   U20115 : XOR2_X1 port map( A1 => n14659, A2 => n14782, Z => n14781);
   U20116 : OAI21_X1 port map( A1 => n24570, A2 => n18091, B => n14662, ZN => 
                           n18092);
   U20117 : XOR2_X1 port map( A1 => n18168, A2 => n1298, Z => n14670);
   U20119 : XOR2_X1 port map( A1 => n14678, A2 => n10716, Z => n14677);
   U20121 : INV_X2 port map( I => n14685, ZN => n19603);
   U20123 : NAND2_X1 port map( A1 => n14960, A2 => n25894, ZN => n18617);
   U20124 : XOR2_X1 port map( A1 => n20489, A2 => n20488, Z => n14700);
   U20125 : XOR2_X1 port map( A1 => n18071, A2 => n18226, Z => n14701);
   U20126 : NOR2_X1 port map( A1 => n6725, A2 => n19033, ZN => n14702);
   U20127 : XOR2_X1 port map( A1 => n28233, A2 => n14631, Z => n14704);
   U20128 : INV_X2 port map( I => n18686, ZN => n18605);
   U20131 : NAND2_X1 port map( A1 => n14720, A2 => n27044, ZN => n14719);
   U20132 : NOR2_X1 port map( A1 => n19167, A2 => n5990, ZN => n14720);
   U20133 : XOR2_X1 port map( A1 => n15844, A2 => Key(94), Z => n15188);
   U20135 : XOR2_X1 port map( A1 => n20449, A2 => n21476, Z => n20451);
   U20136 : XOR2_X1 port map( A1 => n979, A2 => n14640, Z => n14741);
   U20138 : XOR2_X1 port map( A1 => n22774, A2 => n18113, Z => n14746);
   U20142 : XOR2_X1 port map( A1 => n16918, A2 => n21631, Z => n16919);
   U20143 : XOR2_X1 port map( A1 => n23480, A2 => n21705, Z => n18591);
   U20147 : AOI21_X1 port map( A1 => n20043, A2 => n20044, B => n28519, ZN => 
                           n15193);
   U20157 : XOR2_X1 port map( A1 => n16778, A2 => n20702, Z => n15556);
   U20158 : XOR2_X1 port map( A1 => n18353, A2 => n21164, Z => n14813);
   U20166 : XOR2_X1 port map( A1 => n9678, A2 => n22777, Z => n14850);
   U20167 : XOR2_X1 port map( A1 => n21371, A2 => n21434, Z => n14851);
   U20170 : NAND3_X1 port map( A1 => n21444, A2 => n21445, A3 => n21931, ZN => 
                           n15094);
   U20171 : NAND2_X1 port map( A1 => n15282, A2 => n16334, ZN => n14880);
   U20175 : INV_X2 port map( I => n14893, ZN => n15918);
   U20176 : XOR2_X1 port map( A1 => n20385, A2 => n21247, Z => n20368);
   U20177 : INV_X2 port map( I => n17806, ZN => n18262);
   U20180 : NAND2_X1 port map( A1 => n14636, A2 => n21773, ZN => n14909);
   U20181 : NAND2_X1 port map( A1 => n16130, A2 => n838, ZN => n14911);
   U20183 : XOR2_X1 port map( A1 => n20442, A2 => n20076, Z => n14915);
   U20185 : OR2_X1 port map( A1 => n21343, A2 => n2448, Z => n14927);
   U20186 : NAND2_X1 port map( A1 => n21355, A2 => n21342, ZN => n14928);
   U20187 : NAND3_X1 port map( A1 => n14934, A2 => n890, A3 => n7961, ZN => 
                           n14933);
   U20190 : NOR2_X1 port map( A1 => n15981, A2 => n15155, ZN => n15829);
   U20192 : XOR2_X1 port map( A1 => n25946, A2 => n14956, Z => n14955);
   U20197 : XOR2_X1 port map( A1 => n14978, A2 => n21155, Z => n21156);
   U20199 : NAND2_X1 port map( A1 => n14993, A2 => n25141, ZN => n14992);
   U20200 : NAND2_X1 port map( A1 => n11259, A2 => n22374, ZN => n14993);
   U20201 : XOR2_X1 port map( A1 => n28269, A2 => n19346, Z => n14995);
   U20202 : MUX2_X1 port map( I0 => n19982, I1 => n19983, S => n20413, Z => 
                           n19984);
   U20210 : XOR2_X1 port map( A1 => n15387, A2 => n20412, Z => n15017);
   U20211 : XOR2_X1 port map( A1 => n20511, A2 => n21651, Z => n15022);
   U20212 : AOI21_X1 port map( A1 => n20946, A2 => n15023, B => n20945, ZN => 
                           n20947);
   U20213 : XOR2_X1 port map( A1 => n24258, A2 => n21141, Z => n17602);
   U20214 : XOR2_X1 port map( A1 => n24258, A2 => n14593, Z => n18222);
   U20217 : XOR2_X1 port map( A1 => n21192, A2 => n20451, Z => n15039);
   U20219 : XOR2_X1 port map( A1 => n10535, A2 => n15044, Z => n15043);
   U20221 : MUX2_X1 port map( I0 => n15900, I1 => n15901, S => n15970, Z => 
                           n15903);
   U20225 : INV_X2 port map( I => n15432, ZN => n17487);
   U20226 : XOR2_X1 port map( A1 => n24153, A2 => n19886, Z => n15069);
   U20229 : NAND2_X1 port map( A1 => n18976, A2 => n15435, ZN => n15078);
   U20230 : XOR2_X1 port map( A1 => n15782, A2 => Key(150), Z => n16064);
   U20232 : INV_X2 port map( I => n16064, ZN => n16314);
   U20233 : XOR2_X1 port map( A1 => n15090, A2 => n20603, Z => Ciphertext(1));
   U20235 : NOR2_X1 port map( A1 => n8996, A2 => n14509, ZN => n15099);
   U20238 : XOR2_X1 port map( A1 => n24197, A2 => n14591, Z => n20006);
   U20239 : XOR2_X1 port map( A1 => n15119, A2 => n1297, Z => n20370);
   U20240 : XOR2_X1 port map( A1 => n23010, A2 => n14564, Z => n19557);
   U20241 : XOR2_X1 port map( A1 => n16768, A2 => n16746, Z => n16748);
   U20244 : AND2_X1 port map( A1 => n1009, A2 => n18752, Z => n15144);
   U20246 : XOR2_X1 port map( A1 => n20713, A2 => n15149, Z => n15148);
   U20247 : NAND2_X2 port map( A1 => n15153, A2 => n15152, ZN => n21606);
   U20248 : XOR2_X1 port map( A1 => n17113, A2 => n17112, Z => n17250);
   U20251 : XOR2_X1 port map( A1 => n15160, A2 => n21631, Z => Ciphertext(162))
                           ;
   U20255 : XOR2_X1 port map( A1 => n18186, A2 => n15174, Z => n15173);
   U20258 : XOR2_X1 port map( A1 => n19534, A2 => n19216, Z => n15201);
   U20259 : XOR2_X1 port map( A1 => n21158, A2 => n21010, Z => n15183);
   U20260 : INV_X1 port map( I => n21640, ZN => n21634);
   U20261 : XOR2_X1 port map( A1 => n17072, A2 => n17071, Z => n17076);
   U20263 : OR2_X1 port map( A1 => n20184, A2 => n20237, Z => n15194);
   U20265 : XOR2_X1 port map( A1 => n17141, A2 => n14564, Z => n15214);
   U20266 : XOR2_X1 port map( A1 => n16809, A2 => n6932, Z => n15215);
   U20267 : XOR2_X1 port map( A1 => n22829, A2 => n14555, Z => n15221);
   U20269 : OAI21_X1 port map( A1 => n15982, A2 => n26665, B => n14530, ZN => 
                           n15235);
   U20270 : INV_X1 port map( I => n15987, ZN => n15236);
   U20271 : XOR2_X1 port map( A1 => n15237, A2 => n14645, Z => n17658);
   U20272 : XOR2_X1 port map( A1 => n19344, A2 => n19477, Z => n15244);
   U20275 : NOR2_X2 port map( A1 => n21714, A2 => n20642, ZN => n20588);
   U20276 : NOR2_X1 port map( A1 => n16217, A2 => n11080, ZN => n15309);
   U20281 : XOR2_X1 port map( A1 => n17092, A2 => n17091, Z => n15272);
   U20282 : INV_X2 port map( I => n15273, ZN => n17362);
   U20284 : XOR2_X1 port map( A1 => n15293, A2 => n16933, Z => n15292);
   U20285 : XOR2_X1 port map( A1 => n19504, A2 => n10713, Z => n15303);
   U20288 : XOR2_X1 port map( A1 => n20567, A2 => n15319, Z => n15318);
   U20289 : XOR2_X1 port map( A1 => n5446, A2 => n20621, Z => n15319);
   U20291 : XOR2_X1 port map( A1 => n12739, A2 => n21642, Z => n15332);
   U20293 : XOR2_X1 port map( A1 => n24258, A2 => n14614, Z => n18089);
   U20294 : XOR2_X1 port map( A1 => n21184, A2 => n15341, Z => n15340);
   U20295 : XOR2_X1 port map( A1 => n21183, A2 => n21247, Z => n15341);
   U20296 : XNOR2_X1 port map( A1 => Plaintext(28), A2 => Key(28), ZN => n15342
                           );
   U20297 : XOR2_X1 port map( A1 => n19328, A2 => n7050, Z => n19199);
   U20304 : NAND2_X1 port map( A1 => n950, A2 => n20931, ZN => n15365);
   U20309 : INV_X2 port map( I => n15386, ZN => n20736);
   U20310 : XOR2_X1 port map( A1 => n21432, A2 => n20459, Z => n15392);
   U20311 : XOR2_X1 port map( A1 => n24193, A2 => n16855, Z => n15400);
   U20312 : XOR2_X1 port map( A1 => Key(104), A2 => Plaintext(104), Z => n15884
                           );
   U20316 : INV_X1 port map( I => n16434, ZN => n15421);
   U20317 : OR2_X1 port map( A1 => n21646, A2 => n21647, Z => n15428);
   U20318 : NAND2_X1 port map( A1 => n16130, A2 => n15440, ZN => n15842);
   U20320 : XOR2_X1 port map( A1 => n18317, A2 => n20741, Z => n18318);
   U20321 : XOR2_X1 port map( A1 => n27858, A2 => n21106, Z => n15455);
   U20324 : NAND2_X1 port map( A1 => n15469, A2 => n15475, ZN => n15468);
   U20325 : XOR2_X1 port map( A1 => Plaintext(187), A2 => Key(187), Z => n15904
                           );
   U20326 : XOR2_X1 port map( A1 => n14006, A2 => n14609, Z => n16473);
   U20327 : XOR2_X1 port map( A1 => n19461, A2 => n589, Z => n15493);
   U20328 : XOR2_X1 port map( A1 => Plaintext(63), A2 => Key(63), Z => n15872);
   U20329 : XOR2_X1 port map( A1 => n14203, A2 => n14616, Z => n15494);
   U20331 : XOR2_X1 port map( A1 => n25332, A2 => n21104, Z => n19179);
   U20332 : XOR2_X1 port map( A1 => n15734, A2 => n1298, Z => n20409);
   U20333 : NAND2_X2 port map( A1 => n15511, A2 => n15510, ZN => n16731);
   U20334 : INV_X2 port map( I => n15525, ZN => n16021);
   U20335 : NAND2_X1 port map( A1 => n16729, A2 => n1257, ZN => n15527);
   U20340 : XOR2_X1 port map( A1 => n15551, A2 => n14633, Z => Ciphertext(177))
                           ;
   U20341 : XOR2_X1 port map( A1 => n18234, A2 => n20769, Z => n15558);
   U20342 : INV_X2 port map( I => n15559, ZN => n16253);
   U20343 : XNOR2_X1 port map( A1 => Plaintext(186), A2 => Key(186), ZN => 
                           n15559);
   U20344 : INV_X2 port map( I => n15573, ZN => n19808);
   U20345 : XOR2_X1 port map( A1 => n15578, A2 => n15577, Z => n15576);
   U20346 : XOR2_X1 port map( A1 => n16929, A2 => n10544, Z => n15577);
   U20347 : XOR2_X1 port map( A1 => n16930, A2 => n17015, Z => n15578);
   U20348 : OAI21_X1 port map( A1 => n16229, A2 => n10001, B => n16271, ZN => 
                           n15579);
   U20349 : OAI21_X1 port map( A1 => n4739, A2 => n4738, B => n15583, ZN => 
                           n15582);
   U20353 : XOR2_X1 port map( A1 => n19341, A2 => n19342, Z => n15589);
   U20354 : XOR2_X1 port map( A1 => n20481, A2 => n25310, Z => n20461);
   U20355 : XOR2_X1 port map( A1 => n15594, A2 => n16960, Z => n15593);
   U20359 : XOR2_X1 port map( A1 => n3372, A2 => n14620, Z => n19277);
   U20360 : XOR2_X1 port map( A1 => n3372, A2 => n14535, Z => n19320);
   U20364 : XOR2_X1 port map( A1 => n19392, A2 => n19507, Z => n19356);
   U20367 : INV_X2 port map( I => n15670, ZN => n21389);
   U20370 : XOR2_X1 port map( A1 => Key(118), A2 => Plaintext(118), Z => n16184
                           );
   U20374 : AOI21_X1 port map( A1 => n15676, A2 => n16262, B => n16259, ZN => 
                           n15805);
   U20375 : XOR2_X1 port map( A1 => n19419, A2 => n19420, Z => n19426);
   U20376 : INV_X2 port map( I => n15688, ZN => n20739);
   U20377 : XOR2_X1 port map( A1 => n21380, A2 => n20425, Z => n15690);
   U20378 : INV_X2 port map( I => n15698, ZN => n15699);
   U20379 : XOR2_X1 port map( A1 => Plaintext(59), A2 => Key(59), Z => n15923);
   U20380 : MUX2_X1 port map( I0 => n23719, I1 => n24952, S => n1251, Z => 
                           n16463);
   U20383 : INV_X2 port map( I => n15738, ZN => n19798);
   U20384 : XOR2_X1 port map( A1 => n15740, A2 => n15739, Z => n15738);
   U20388 : NAND2_X1 port map( A1 => n25324, A2 => n20685, ZN => n20679);
   U20392 : CLKBUF_X2 port map( I => Key(111), Z => n21707);
   U20394 : NOR2_X1 port map( A1 => n21161, A2 => n21160, ZN => n20557);
   U20395 : INV_X1 port map( I => n16498, ZN => n16397);
   U20396 : NOR2_X2 port map( A1 => n16092, A2 => n10696, ZN => n16098);
   U20406 : BUF_X2 port map( I => Key(163), Z => n21631);
   U20407 : XOR2_X1 port map( A1 => Key(33), A2 => Plaintext(33), Z => n16343);
   U20408 : XOR2_X1 port map( A1 => Key(34), A2 => Plaintext(34), Z => n15922);
   U20409 : XOR2_X1 port map( A1 => Key(31), A2 => Plaintext(31), Z => n16342);
   U20410 : INV_X1 port map( I => Plaintext(14), ZN => n15757);
   U20411 : XOR2_X1 port map( A1 => n15757, A2 => Key(14), Z => n15894);
   U20412 : XOR2_X1 port map( A1 => Key(17), A2 => Plaintext(17), Z => n15758);
   U20413 : INV_X1 port map( I => Plaintext(16), ZN => n15759);
   U20414 : XOR2_X1 port map( A1 => n15759, A2 => Key(16), Z => n16209);
   U20415 : INV_X1 port map( I => Plaintext(39), ZN => n15762);
   U20416 : XOR2_X1 port map( A1 => n15762, A2 => Key(39), Z => n15929);
   U20418 : INV_X1 port map( I => Plaintext(49), ZN => n15763);
   U20419 : XOR2_X1 port map( A1 => n15763, A2 => Key(49), Z => n15869);
   U20420 : XOR2_X1 port map( A1 => Key(48), A2 => Plaintext(48), Z => n16128);
   U20421 : INV_X1 port map( I => Plaintext(53), ZN => n15764);
   U20422 : XOR2_X1 port map( A1 => n15764, A2 => Key(53), Z => n16126);
   U20423 : NOR2_X1 port map( A1 => n15869, A2 => n16123, ZN => n15767);
   U20425 : NOR2_X1 port map( A1 => n16115, A2 => n14644, ZN => n15769);
   U20426 : XOR2_X1 port map( A1 => Key(58), A2 => Plaintext(58), Z => n15924);
   U20429 : XOR2_X1 port map( A1 => Key(42), A2 => Plaintext(42), Z => n15957);
   U20430 : INV_X1 port map( I => Plaintext(45), ZN => n15773);
   U20431 : XOR2_X1 port map( A1 => n15773, A2 => Key(45), Z => n15958);
   U20432 : INV_X1 port map( I => Plaintext(43), ZN => n15774);
   U20433 : XOR2_X1 port map( A1 => n15774, A2 => Key(43), Z => n15934);
   U20434 : XOR2_X1 port map( A1 => Key(62), A2 => Plaintext(62), Z => n16131);
   U20435 : NAND2_X1 port map( A1 => n21773, A2 => n7235, ZN => n15775);
   U20437 : INV_X1 port map( I => Plaintext(155), ZN => n15779);
   U20439 : INV_X1 port map( I => Plaintext(154), ZN => n15781);
   U20440 : XOR2_X1 port map( A1 => n15781, A2 => Key(154), Z => n16066);
   U20441 : XOR2_X1 port map( A1 => Key(153), A2 => Plaintext(153), Z => n16068
                           );
   U20442 : INV_X1 port map( I => Plaintext(150), ZN => n15782);
   U20445 : INV_X1 port map( I => Plaintext(131), ZN => n15786);
   U20446 : XOR2_X1 port map( A1 => n15786, A2 => Key(131), Z => n16325);
   U20451 : XOR2_X1 port map( A1 => Key(133), A2 => Plaintext(133), Z => n16158
                           );
   U20452 : XOR2_X1 port map( A1 => Key(132), A2 => Plaintext(132), Z => n16159
                           );
   U20453 : NAND2_X1 port map( A1 => n16159, A2 => n16158, ZN => n16156);
   U20454 : INV_X1 port map( I => n16156, ZN => n15793);
   U20455 : NAND2_X1 port map( A1 => n15793, A2 => n25135, ZN => n15794);
   U20456 : INV_X1 port map( I => Plaintext(177), ZN => n15795);
   U20457 : XOR2_X1 port map( A1 => Key(179), A2 => Plaintext(179), Z => n15796
                           );
   U20458 : XOR2_X1 port map( A1 => Key(2), A2 => Plaintext(2), Z => n15889);
   U20460 : NAND3_X1 port map( A1 => n15892, A2 => n21873, A3 => n7374, ZN => 
                           n15799);
   U20461 : XOR2_X1 port map( A1 => Key(166), A2 => Plaintext(166), Z => n16093
                           );
   U20462 : INV_X1 port map( I => Plaintext(167), ZN => n15800);
   U20463 : XOR2_X1 port map( A1 => n15800, A2 => Key(167), Z => n16260);
   U20464 : INV_X2 port map( I => n16260, ZN => n16231);
   U20465 : INV_X1 port map( I => Plaintext(162), ZN => n15801);
   U20467 : XOR2_X1 port map( A1 => Key(164), A2 => Plaintext(164), Z => n15909
                           );
   U20469 : XOR2_X1 port map( A1 => Key(185), A2 => Plaintext(185), Z => n15806
                           );
   U20470 : XOR2_X1 port map( A1 => Key(184), A2 => Plaintext(184), Z => n16227
                           );
   U20471 : NOR2_X1 port map( A1 => n16266, A2 => n16080, ZN => n15811);
   U20473 : XOR2_X1 port map( A1 => Key(171), A2 => Plaintext(171), Z => n16274
                           );
   U20474 : NOR2_X1 port map( A1 => n13577, A2 => n14763, ZN => n15814);
   U20475 : INV_X1 port map( I => Plaintext(77), ZN => n15817);
   U20477 : INV_X1 port map( I => Plaintext(73), ZN => n15819);
   U20482 : XOR2_X1 port map( A1 => Key(82), A2 => Plaintext(82), Z => n15834);
   U20484 : XOR2_X1 port map( A1 => Key(68), A2 => Plaintext(68), Z => n16143);
   U20485 : INV_X1 port map( I => Plaintext(71), ZN => n15824);
   U20486 : XOR2_X1 port map( A1 => n15824, A2 => Key(71), Z => n15835);
   U20488 : XOR2_X1 port map( A1 => Key(86), A2 => Plaintext(86), Z => n15832);
   U20489 : NOR2_X1 port map( A1 => n16203, A2 => n8684, ZN => n15833);
   U20490 : XOR2_X1 port map( A1 => Key(85), A2 => Plaintext(85), Z => n15848);
   U20491 : NAND2_X1 port map( A1 => n16147, A2 => n15986, ZN => n15838);
   U20493 : INV_X1 port map( I => Plaintext(95), ZN => n15843);
   U20494 : INV_X1 port map( I => Plaintext(94), ZN => n15844);
   U20495 : INV_X1 port map( I => Plaintext(93), ZN => n15845);
   U20496 : XOR2_X1 port map( A1 => n15845, A2 => Key(93), Z => n15917);
   U20497 : INV_X1 port map( I => n16012, ZN => n16009);
   U20498 : INV_X1 port map( I => Plaintext(115), ZN => n15850);
   U20499 : XOR2_X1 port map( A1 => n15850, A2 => Key(115), Z => n16166);
   U20500 : XOR2_X1 port map( A1 => Key(117), A2 => Plaintext(117), Z => n16165
                           );
   U20501 : INV_X1 port map( I => Plaintext(114), ZN => n15851);
   U20502 : XOR2_X1 port map( A1 => Key(101), A2 => Plaintext(101), Z => n15881
                           );
   U20503 : INV_X1 port map( I => Plaintext(99), ZN => n15856);
   U20505 : XOR2_X1 port map( A1 => Key(96), A2 => Plaintext(96), Z => n16006);
   U20507 : XOR2_X1 port map( A1 => Key(106), A2 => Plaintext(106), Z => n16190
                           );
   U20508 : XOR2_X1 port map( A1 => Key(103), A2 => Plaintext(103), Z => n16187
                           );
   U20509 : XOR2_X1 port map( A1 => Key(113), A2 => Plaintext(113), Z => n15859
                           );
   U20510 : XOR2_X1 port map( A1 => Key(124), A2 => Plaintext(124), Z => n16331
                           );
   U20512 : NOR2_X1 port map( A1 => n16011, A2 => n16009, ZN => n15865);
   U20515 : INV_X1 port map( I => n15869, ZN => n16127);
   U20518 : NAND2_X1 port map( A1 => n15983, A2 => n15982, ZN => n15875);
   U20520 : NAND2_X1 port map( A1 => n13343, A2 => n22623, ZN => n15897);
   U20522 : NAND2_X1 port map( A1 => n16080, A2 => n22910, ZN => n15901);
   U20523 : INV_X1 port map( I => n15904, ZN => n16255);
   U20524 : NAND2_X1 port map( A1 => n15685, A2 => n15796, ZN => n15908);
   U20525 : NOR2_X1 port map( A1 => n14306, A2 => n14171, ZN => n15914);
   U20526 : MUX2_X1 port map( I0 => n15914, I1 => n15913, S => n7460, Z => 
                           n15915);
   U20527 : NAND2_X1 port map( A1 => n15924, A2 => n15923, ZN => n16133);
   U20528 : NOR3_X1 port map( A1 => n5095, A2 => n15995, A3 => n16123, ZN => 
                           n16697);
   U20532 : INV_X1 port map( I => n15957, ZN => n16119);
   U20534 : NAND2_X1 port map( A1 => n21773, A2 => n14386, ZN => n15974);
   U20539 : NAND3_X1 port map( A1 => n15998, A2 => n14584, A3 => n13731, ZN => 
                           n15999);
   U20543 : NAND2_X1 port map( A1 => n16639, A2 => n16597, ZN => n16025);
   U20545 : NAND2_X1 port map( A1 => n16034, A2 => n16304, ZN => n16035);
   U20549 : NOR2_X1 port map( A1 => n16064, A2 => n16240, ZN => n16067);
   U20550 : INV_X1 port map( I => n24872, ZN => n16315);
   U20551 : NOR2_X1 port map( A1 => n16258, A2 => n16095, ZN => n16070);
   U20552 : NOR2_X1 port map( A1 => n16071, A2 => n16070, ZN => n16075);
   U20553 : NAND2_X1 port map( A1 => n16264, A2 => n16072, ZN => n16074);
   U20554 : NAND2_X1 port map( A1 => n16231, A2 => n16230, ZN => n16073);
   U20555 : NAND3_X1 port map( A1 => n2814, A2 => n1032, A3 => n14861, ZN => 
                           n16358);
   U20557 : OAI21_X1 port map( A1 => n16089, A2 => n16275, B => n13577, ZN => 
                           n16090);
   U20558 : INV_X1 port map( I => n16093, ZN => n16263);
   U20559 : NOR2_X1 port map( A1 => n16263, A2 => n16258, ZN => n16096);
   U20560 : AOI21_X1 port map( A1 => n16096, A2 => n16095, B => n16094, ZN => 
                           n16097);
   U20565 : AOI21_X1 port map( A1 => n16160, A2 => n12509, B => n16321, ZN => 
                           n16161);
   U20566 : NOR2_X2 port map( A1 => n16162, A2 => n16161, ZN => n16526);
   U20567 : NOR2_X1 port map( A1 => n16287, A2 => n16292, ZN => n16163);
   U20569 : AOI21_X1 port map( A1 => n4751, A2 => n14559, B => n16168, ZN => 
                           n16169);
   U20571 : AOI21_X1 port map( A1 => n16685, A2 => n16176, B => n10261, ZN => 
                           n16178);
   U20572 : NAND2_X1 port map( A1 => n28032, A2 => n577, ZN => n16181);
   U20573 : NAND2_X1 port map( A1 => n16182, A2 => n16292, ZN => n16183);
   U20574 : INV_X1 port map( I => n16187, ZN => n16301);
   U20575 : NOR2_X1 port map( A1 => n16573, A2 => n16513, ZN => n16204);
   U20579 : NAND2_X1 port map( A1 => n16657, A2 => n2391, ZN => n16221);
   U20581 : OAI22_X1 port map( A1 => n16221, A2 => n24580, B1 => n16563, B2 => 
                           n16561, ZN => n16222);
   U20583 : NOR2_X1 port map( A1 => n16234, A2 => n16263, ZN => n16235);
   U20584 : OAI21_X1 port map( A1 => n16236, A2 => n16235, B => n16264, ZN => 
                           n16237);
   U20586 : NAND4_X1 port map( A1 => n10767, A2 => n26659, A3 => n16251, A4 => 
                           n16250, ZN => n16249);
   U20587 : NAND2_X1 port map( A1 => n15565, A2 => n16258, ZN => n16265);
   U20589 : NAND2_X1 port map( A1 => n14452, A2 => n26982, ZN => n16285);
   U20592 : OAI21_X1 port map( A1 => n16351, A2 => n21873, B => n10970, ZN => 
                           n16352);
   U20593 : NAND3_X1 port map( A1 => n23227, A2 => n26161, A3 => n1032, ZN => 
                           n16356);
   U20594 : NOR2_X1 port map( A1 => n4630, A2 => n23505, ZN => n16366);
   U20597 : AOI21_X1 port map( A1 => n16609, A2 => n27019, B => n4644, ZN => 
                           n16379);
   U20598 : NAND2_X1 port map( A1 => n16685, A2 => n16380, ZN => n16381);
   U20601 : AOI21_X1 port map( A1 => n16644, A2 => n14968, B => n27372, ZN => 
                           n16402);
   U20602 : NOR2_X1 port map( A1 => n26262, A2 => n16699, ZN => n16407);
   U20603 : NAND2_X1 port map( A1 => n1045, A2 => n16715, ZN => n16415);
   U20604 : XOR2_X1 port map( A1 => n17038, A2 => n14623, Z => n16417);
   U20606 : NAND3_X1 port map( A1 => n22660, A2 => n7378, A3 => n16574, ZN => 
                           n16441);
   U20607 : NAND2_X1 port map( A1 => n16518, A2 => n1052, ZN => n16443);
   U20608 : NAND3_X1 port map( A1 => n16447, A2 => n16446, A3 => n16445, ZN => 
                           n16448);
   U20612 : NOR2_X1 port map( A1 => n16455, A2 => n16651, ZN => n16457);
   U20613 : XOR2_X1 port map( A1 => n16913, A2 => n14624, Z => n16464);
   U20617 : XOR2_X1 port map( A1 => n16817, A2 => n20941, Z => n16501);
   U20618 : XOR2_X1 port map( A1 => n23369, A2 => n14596, Z => n16520);
   U20620 : NOR2_X1 port map( A1 => n4938, A2 => n16810, ZN => n16528);
   U20622 : NAND2_X1 port map( A1 => n16587, A2 => n25255, ZN => n16589);
   U20626 : NAND3_X1 port map( A1 => n16621, A2 => n718, A3 => n16620, ZN => 
                           n16623);
   U20628 : OR2_X1 port map( A1 => n16634, A2 => n1051, Z => n16635);
   U20630 : XOR2_X1 port map( A1 => n25159, A2 => n19218, Z => n16666);
   U20632 : NOR2_X1 port map( A1 => n15701, A2 => n16728, ZN => n16719);
   U20633 : NOR2_X1 port map( A1 => n794, A2 => n1257, ZN => n16718);
   U20635 : INV_X1 port map( I => n16722, ZN => n17486);
   U20636 : NAND2_X1 port map( A1 => n14968, A2 => n1241, ZN => n16737);
   U20637 : XOR2_X1 port map( A1 => n2266, A2 => n21422, Z => n16739);
   U20639 : XOR2_X1 port map( A1 => n16801, A2 => n21436, Z => n16745);
   U20640 : XOR2_X1 port map( A1 => n17116, A2 => n24000, Z => n16749);
   U20641 : XOR2_X1 port map( A1 => n16957, A2 => n20621, Z => n16752);
   U20642 : XOR2_X1 port map( A1 => n16881, A2 => n16755, Z => n16756);
   U20646 : XOR2_X1 port map( A1 => n17102, A2 => n16769, Z => n16773);
   U20647 : XOR2_X1 port map( A1 => n6345, A2 => n14489, Z => n16771);
   U20649 : XOR2_X1 port map( A1 => n17147, A2 => n16924, Z => n16960);
   U20651 : XOR2_X1 port map( A1 => n23779, A2 => n16944, Z => n16781);
   U20653 : XOR2_X1 port map( A1 => n23779, A2 => n16861, Z => n16783);
   U20654 : XOR2_X1 port map( A1 => n17125, A2 => n21384, Z => n16787);
   U20655 : XOR2_X1 port map( A1 => n16788, A2 => n16787, Z => n16789);
   U20656 : XOR2_X1 port map( A1 => n16975, A2 => n20674, Z => n16793);
   U20657 : XOR2_X1 port map( A1 => n17028, A2 => n3001, Z => n16794);
   U20658 : XOR2_X1 port map( A1 => n16818, A2 => n9902, Z => n16795);
   U20663 : XOR2_X1 port map( A1 => n6932, A2 => n14549, Z => n16808);
   U20664 : NAND3_X1 port map( A1 => n16815, A2 => n16812, A3 => n16814, ZN => 
                           n16816);
   U20668 : XOR2_X1 port map( A1 => n17085, A2 => n10535, Z => n16830);
   U20670 : INV_X1 port map( I => n16846, ZN => n17509);
   U20671 : XOR2_X1 port map( A1 => n17150, A2 => n16835, Z => n16839);
   U20672 : XOR2_X1 port map( A1 => n25933, A2 => n2266, Z => n16838);
   U20675 : XOR2_X1 port map( A1 => n17141, A2 => n14405, Z => n16840);
   U20677 : XOR2_X1 port map( A1 => n16929, A2 => n17077, Z => n16849);
   U20678 : XOR2_X1 port map( A1 => n25683, A2 => n16849, Z => n16850);
   U20679 : XOR2_X1 port map( A1 => n16851, A2 => n16850, Z => n17422);
   U20680 : XOR2_X1 port map( A1 => n16910, A2 => n14436, Z => n16860);
   U20681 : XOR2_X1 port map( A1 => n16865, A2 => n16864, Z => n16866);
   U20683 : XOR2_X1 port map( A1 => n26082, A2 => n14638, Z => n16873);
   U20684 : NAND2_X1 port map( A1 => n17447, A2 => n17381, ZN => n16878);
   U20685 : XOR2_X1 port map( A1 => n12410, A2 => n20617, Z => n16876);
   U20687 : XOR2_X1 port map( A1 => n16883, A2 => n14360, Z => n16884);
   U20688 : XOR2_X1 port map( A1 => n17126, A2 => n16884, Z => n16885);
   U20689 : XOR2_X1 port map( A1 => n16931, A2 => n14335, Z => n16898);
   U20690 : XOR2_X1 port map( A1 => n27969, A2 => n14597, Z => n16900);
   U20691 : XOR2_X1 port map( A1 => n16899, A2 => n16900, Z => n16901);
   U20692 : AOI21_X1 port map( A1 => n17391, A2 => n9252, B => n15504, ZN => 
                           n16902);
   U20693 : XOR2_X1 port map( A1 => n17094, A2 => n14652, Z => n16906);
   U20695 : INV_X1 port map( I => n17088, ZN => n16912);
   U20696 : XOR2_X1 port map( A1 => n6878, A2 => n17044, Z => n16920);
   U20697 : XOR2_X1 port map( A1 => n16920, A2 => n16919, Z => n16921);
   U20699 : XOR2_X1 port map( A1 => n14123, A2 => n20967, Z => n16928);
   U20700 : XOR2_X1 port map( A1 => n12410, A2 => n20989, Z => n16933);
   U20703 : INV_X1 port map( I => n19346, ZN => n21533);
   U20705 : XOR2_X1 port map( A1 => n10538, A2 => n16961, Z => n16962);
   U20707 : XOR2_X1 port map( A1 => n17055, A2 => n16975, Z => n16976);
   U20711 : XOR2_X1 port map( A1 => n17009, A2 => n17010, Z => n17011);
   U20712 : XOR2_X1 port map( A1 => n17012, A2 => n17011, Z => n17469);
   U20713 : XOR2_X1 port map( A1 => n17017, A2 => n17018, Z => n17293);
   U20714 : XOR2_X1 port map( A1 => n6345, A2 => n21642, Z => n17019);
   U20715 : OAI21_X1 port map( A1 => n17318, A2 => n22840, B => n6624, ZN => 
                           n17021);
   U20716 : NAND3_X1 port map( A1 => n17286, A2 => n17317, A3 => n17318, ZN => 
                           n17023);
   U20719 : XOR2_X1 port map( A1 => n17109, A2 => n21037, Z => n17030);
   U20720 : XOR2_X1 port map( A1 => n17038, A2 => n17098, Z => n17041);
   U20721 : XOR2_X1 port map( A1 => n17039, A2 => n14645, Z => n17040);
   U20722 : XOR2_X1 port map( A1 => n17041, A2 => n17040, Z => n17042);
   U20725 : XOR2_X1 port map( A1 => n17056, A2 => n17055, Z => n17057);
   U20726 : XOR2_X1 port map( A1 => n2266, A2 => n17065, Z => n17066);
   U20727 : XOR2_X1 port map( A1 => n17070, A2 => n21033, Z => n17071);
   U20729 : XOR2_X1 port map( A1 => n1237, A2 => n14457, Z => n17089);
   U20730 : XOR2_X1 port map( A1 => n17098, A2 => n20961, Z => n17101);
   U20733 : XOR2_X1 port map( A1 => n12410, A2 => n21650, Z => n17110);
   U20734 : XOR2_X1 port map( A1 => n5499, A2 => n17117, Z => n17120);
   U20735 : XOR2_X1 port map( A1 => n17120, A2 => n17119, Z => n17122);
   U20736 : XOR2_X1 port map( A1 => n12831, A2 => n21649, Z => n17128);
   U20739 : NAND2_X1 port map( A1 => n17163, A2 => n17286, ZN => n17164);
   U20743 : NOR2_X1 port map( A1 => n23571, A2 => n17526, ZN => n17195);
   U20754 : OAI21_X1 port map( A1 => n3376, A2 => n10568, B => n24070, ZN => 
                           n17259);
   U20757 : NAND3_X1 port map( A1 => n10015, A2 => n17530, A3 => n17421, ZN => 
                           n17272);
   U20760 : MUX2_X1 port map( I0 => n9865, I1 => n17036, S => n17204, Z => 
                           n17288);
   U20763 : NAND2_X1 port map( A1 => n7275, A2 => n17513, ZN => n17300);
   U20764 : NAND2_X1 port map( A1 => n17302, A2 => n17301, ZN => n17305);
   U20765 : MUX2_X1 port map( I0 => n17305, I1 => n17304, S => n17306, Z => 
                           n17310);
   U20767 : AOI21_X1 port map( A1 => n27947, A2 => n17962, B => n1025, ZN => 
                           n17333);
   U20768 : NAND3_X1 port map( A1 => n7361, A2 => n17567, A3 => n8593, ZN => 
                           n17340);
   U20771 : XOR2_X1 port map( A1 => n28265, A2 => n22165, Z => n17351);
   U20772 : XOR2_X1 port map( A1 => n18316, A2 => n17351, Z => n17399);
   U20773 : OAI21_X1 port map( A1 => n17479, A2 => n17353, B => n26418, ZN => 
                           n17354);
   U20781 : NAND2_X1 port map( A1 => n24517, A2 => n10546, ZN => n17380);
   U20782 : XOR2_X1 port map( A1 => n18182, A2 => n7368, Z => n17396);
   U20783 : XOR2_X1 port map( A1 => n17397, A2 => n17396, Z => n17398);
   U20785 : NAND2_X1 port map( A1 => n25380, A2 => n12225, ZN => n17424);
   U20789 : MUX2_X1 port map( I0 => n17450, I1 => n17518, S => n27959, Z => 
                           n17451);
   U20795 : INV_X1 port map( I => n7102, ZN => n17504);
   U20797 : INV_X1 port map( I => n17538, ZN => n17539);
   U20798 : NAND2_X1 port map( A1 => n17541, A2 => n17540, ZN => n17550);
   U20802 : MUX2_X1 port map( I0 => n17565, I1 => n17563, S => n17735, Z => 
                           n17568);
   U20803 : NAND2_X1 port map( A1 => n24304, A2 => n5218, ZN => n17587);
   U20806 : XOR2_X1 port map( A1 => n18110, A2 => n18142, Z => n17601);
   U20807 : XOR2_X1 port map( A1 => n17602, A2 => n17601, Z => n17603);
   U20809 : NAND2_X1 port map( A1 => n9485, A2 => n18005, ZN => n17606);
   U20812 : XOR2_X1 port map( A1 => n18179, A2 => n15669, Z => n17627);
   U20814 : XOR2_X1 port map( A1 => n17659, A2 => n17658, Z => n17660);
   U20818 : NOR2_X1 port map( A1 => n21898, A2 => n885, ZN => n17669);
   U20819 : XOR2_X1 port map( A1 => n28393, A2 => n20702, Z => n17671);
   U20823 : NAND2_X1 port map( A1 => n413, A2 => n17694, ZN => n17695);
   U20827 : XOR2_X1 port map( A1 => n18179, A2 => n18352, Z => n17707);
   U20833 : XOR2_X1 port map( A1 => n14203, A2 => n20807, Z => n17721);
   U20834 : NOR2_X1 port map( A1 => n17724, A2 => n17726, ZN => n17725);
   U20836 : INV_X1 port map( I => n17733, ZN => n17734);
   U20837 : NAND2_X1 port map( A1 => n17734, A2 => n26308, ZN => n17738);
   U20838 : NAND2_X1 port map( A1 => n26308, A2 => n17735, ZN => n17737);
   U20839 : NAND2_X1 port map( A1 => n18665, A2 => n14510, ZN => n17747);
   U20841 : XOR2_X1 port map( A1 => n18012, A2 => n20766, Z => n17765);
   U20843 : NAND2_X1 port map( A1 => n17773, A2 => n4812, ZN => n17776);
   U20844 : XOR2_X1 port map( A1 => n20727, A2 => n18211, Z => n17778);
   U20845 : XOR2_X1 port map( A1 => n17779, A2 => n17778, Z => n17780);
   U20848 : NAND2_X1 port map( A1 => n13621, A2 => n12815, ZN => n17805);
   U20849 : NAND2_X1 port map( A1 => n18741, A2 => n27715, ZN => n17815);
   U20850 : XOR2_X1 port map( A1 => n18119, A2 => n17823, Z => n17828);
   U20851 : XOR2_X1 port map( A1 => n18246, A2 => n18021, Z => n18114);
   U20852 : XOR2_X1 port map( A1 => n27384, A2 => n18168, Z => n18219);
   U20853 : XOR2_X1 port map( A1 => n18274, A2 => n18219, Z => n17839);
   U20854 : XOR2_X1 port map( A1 => n18063, A2 => n18070, Z => n17838);
   U20855 : XOR2_X1 port map( A1 => n18022, A2 => n14518, Z => n17837);
   U20859 : INV_X1 port map( I => n18569, ZN => n18643);
   U20860 : INV_X1 port map( I => n18066, ZN => n17884);
   U20861 : NAND2_X1 port map( A1 => n17887, A2 => n22646, ZN => n17885);
   U20862 : XOR2_X1 port map( A1 => n18280, A2 => n7387, Z => n17909);
   U20866 : INV_X1 port map( I => n9636, ZN => n17937);
   U20869 : NAND2_X1 port map( A1 => n14342, A2 => n17989, ZN => n17990);
   U20871 : XOR2_X1 port map( A1 => n18097, A2 => n21143, Z => n18009);
   U20872 : XOR2_X1 port map( A1 => n18074, A2 => n1061, Z => n18010);
   U20873 : XOR2_X1 port map( A1 => n25901, A2 => n7409, Z => n18017);
   U20874 : XOR2_X1 port map( A1 => n13410, A2 => n18017, Z => n18018);
   U20875 : XOR2_X1 port map( A1 => n22126, A2 => n13686, Z => n18020);
   U20876 : XOR2_X1 port map( A1 => n18022, A2 => n14404, Z => n18023);
   U20877 : XOR2_X1 port map( A1 => n18024, A2 => n18023, Z => n18025);
   U20878 : XOR2_X1 port map( A1 => n18147, A2 => n21553, Z => n18033);
   U20881 : XOR2_X1 port map( A1 => n18135, A2 => n1305, Z => n18045);
   U20882 : XOR2_X1 port map( A1 => n13464, A2 => n18049, Z => n18050);
   U20883 : XOR2_X1 port map( A1 => n18132, A2 => n14604, Z => n18052);
   U20884 : XOR2_X1 port map( A1 => n18053, A2 => n18052, Z => n18054);
   U20886 : XOR2_X1 port map( A1 => n18209, A2 => n18226, Z => n18073);
   U20887 : XOR2_X1 port map( A1 => n18074, A2 => n14488, Z => n18075);
   U20889 : XOR2_X1 port map( A1 => n25892, A2 => n20467, Z => n18083);
   U20891 : XOR2_X1 port map( A1 => n18241, A2 => n20912, Z => n18108);
   U20893 : XOR2_X1 port map( A1 => n18301, A2 => n13686, Z => n18118);
   U20894 : XOR2_X1 port map( A1 => n18120, A2 => n20692, Z => n18121);
   U20895 : INV_X1 port map( I => n18225, ZN => n18134);
   U20896 : XOR2_X1 port map( A1 => n18137, A2 => n14418, Z => n18138);
   U20897 : INV_X1 port map( I => n18146, ZN => n18377);
   U20898 : XOR2_X1 port map( A1 => n18147, A2 => n20614, Z => n18148);
   U20899 : XOR2_X1 port map( A1 => n25312, A2 => n23186, Z => n18150);
   U20900 : XOR2_X1 port map( A1 => n18149, A2 => n18150, Z => n18154);
   U20901 : XOR2_X1 port map( A1 => n18171, A2 => n20674, Z => n18151);
   U20902 : XOR2_X1 port map( A1 => n18152, A2 => n18151, Z => n18153);
   U20904 : XOR2_X1 port map( A1 => n14066, A2 => n20952, Z => n18157);
   U20905 : XOR2_X1 port map( A1 => n18158, A2 => n18157, Z => n18159);
   U20906 : XOR2_X1 port map( A1 => n18160, A2 => n18159, Z => n18601);
   U20907 : NAND2_X1 port map( A1 => n18472, A2 => n18458, ZN => n18176);
   U20908 : NAND3_X1 port map( A1 => n18412, A2 => n14408, A3 => n376, ZN => 
                           n18177);
   U20909 : XOR2_X1 port map( A1 => n18182, A2 => n20872, Z => n18183);
   U20910 : XOR2_X1 port map( A1 => n1194, A2 => n14640, Z => n18185);
   U20911 : XOR2_X1 port map( A1 => n18184, A2 => n18185, Z => n18188);
   U20912 : XOR2_X1 port map( A1 => n18187, A2 => n18188, Z => n18609);
   U20917 : XOR2_X1 port map( A1 => n18206, A2 => n14432, Z => n18207);
   U20918 : XOR2_X1 port map( A1 => n280, A2 => n18221, Z => n18223);
   U20919 : XOR2_X1 port map( A1 => n18227, A2 => n1292, Z => n18228);
   U20922 : XOR2_X1 port map( A1 => n18263, A2 => n18249, Z => n18251);
   U20923 : XOR2_X1 port map( A1 => n698, A2 => n20617, Z => n18250);
   U20924 : XOR2_X1 port map( A1 => n14215, A2 => n21476, Z => n18260);
   U20925 : XOR2_X1 port map( A1 => n18261, A2 => n18260, Z => n18266);
   U20926 : XOR2_X1 port map( A1 => n26486, A2 => n18262, Z => n18265);
   U20930 : XOR2_X1 port map( A1 => n18288, A2 => n18287, Z => n18289);
   U20932 : XOR2_X1 port map( A1 => n18307, A2 => n14558, Z => n18308);
   U20936 : XOR2_X1 port map( A1 => n27348, A2 => n14581, Z => n18325);
   U20937 : NAND3_X1 port map( A1 => n18377, A2 => n14494, A3 => n5434, ZN => 
                           n18343);
   U20938 : XOR2_X1 port map( A1 => n28393, A2 => n14491, Z => n18345);
   U20939 : XOR2_X1 port map( A1 => n18346, A2 => n18345, Z => n18350);
   U20941 : INV_X1 port map( I => n18360, ZN => n18361);
   U20942 : NOR2_X1 port map( A1 => n18581, A2 => n18531, ZN => n18372);
   U20948 : AOI21_X1 port map( A1 => n18419, A2 => n18739, B => n26894, ZN => 
                           n18421);
   U20950 : NAND3_X1 port map( A1 => n24207, A2 => n14140, A3 => n18428, ZN => 
                           n18429);
   U20951 : XOR2_X1 port map( A1 => n19430, A2 => n14633, Z => n18436);
   U20952 : XOR2_X1 port map( A1 => n19315, A2 => n18436, Z => n18437);
   U20955 : NAND2_X1 port map( A1 => n18610, A2 => n18697, ZN => n18453);
   U20957 : NAND2_X1 port map( A1 => n18556, A2 => n6800, ZN => n18464);
   U20958 : NOR2_X1 port map( A1 => n26880, A2 => n18697, ZN => n18469);
   U20961 : NAND2_X1 port map( A1 => n14332, A2 => n18666, ZN => n18480);
   U20962 : INV_X1 port map( I => n23841, ZN => n18493);
   U20963 : NOR2_X1 port map( A1 => n18653, A2 => n18493, ZN => n18494);
   U20968 : XOR2_X1 port map( A1 => n18521, A2 => n18520, Z => n19863);
   U20970 : NAND2_X1 port map( A1 => n11685, A2 => n18589, ZN => n18528);
   U20971 : NAND3_X1 port map( A1 => n18540, A2 => n18539, A3 => n18538, ZN => 
                           n18544);
   U20974 : NAND2_X1 port map( A1 => n14376, A2 => n18749, ZN => n18571);
   U20975 : NOR2_X1 port map( A1 => n19123, A2 => n12583, ZN => n18577);
   U20978 : NOR2_X1 port map( A1 => n26277, A2 => n4661, ZN => n18592);
   U20979 : NAND3_X1 port map( A1 => n28106, A2 => n26277, A3 => n28481, ZN => 
                           n18595);
   U20981 : INV_X1 port map( I => n14959, ZN => n18603);
   U20982 : NAND2_X1 port map( A1 => n18603, A2 => n18949, ZN => n18619);
   U20983 : NOR2_X1 port map( A1 => n18610, A2 => n18609, ZN => n18611);
   U20986 : NAND3_X1 port map( A1 => n18769, A2 => n18770, A3 => n8576, ZN => 
                           n18635);
   U20991 : NOR2_X1 port map( A1 => n18673, A2 => n24672, ZN => n18676);
   U20995 : NAND2_X1 port map( A1 => n18715, A2 => n13372, ZN => n18717);
   U20996 : NAND2_X1 port map( A1 => n18720, A2 => n1184, ZN => n18721);
   U20997 : INV_X1 port map( I => n19135, ZN => n18731);
   U20999 : MUX2_X1 port map( I0 => n12139, I1 => n18760, S => n18971, Z => 
                           n18765);
   U21002 : NAND2_X1 port map( A1 => n18798, A2 => n18799, ZN => n18801);
   U21005 : INV_X1 port map( I => n18813, ZN => n18818);
   U21006 : INV_X1 port map( I => n18814, ZN => n18817);
   U21007 : NAND2_X1 port map( A1 => n19225, A2 => n18871, ZN => n18826);
   U21008 : NAND2_X1 port map( A1 => n18932, A2 => n18828, ZN => n18830);
   U21012 : XOR2_X1 port map( A1 => n19220, A2 => n21553, Z => n18857);
   U21016 : NOR2_X1 port map( A1 => n18995, A2 => n23546, ZN => n18903);
   U21018 : XOR2_X1 port map( A1 => n25098, A2 => n20871, Z => n18916);
   U21019 : XOR2_X1 port map( A1 => n2467, A2 => n21482, Z => n18937);
   U21023 : NOR2_X1 port map( A1 => n12521, A2 => n19073, ZN => n18976);
   U21025 : OAI21_X1 port map( A1 => n27465, A2 => n997, B => n19086, ZN => 
                           n19000);
   U21030 : NAND2_X1 port map( A1 => n19053, A2 => n28372, ZN => n19054);
   U21032 : XOR2_X1 port map( A1 => n24501, A2 => n14598, Z => n19065);
   U21033 : XOR2_X1 port map( A1 => n6539, A2 => n19065, Z => n19066);
   U21035 : XOR2_X1 port map( A1 => n27362, A2 => n14555, Z => n19072);
   U21036 : XOR2_X1 port map( A1 => n19317, A2 => n19072, Z => n19084);
   U21037 : NAND2_X1 port map( A1 => n25559, A2 => n15429, ZN => n19078);
   U21039 : NOR2_X1 port map( A1 => n1125, A2 => n669, ZN => n19153);
   U21041 : XOR2_X1 port map( A1 => n11328, A2 => n7346, Z => n19174);
   U21042 : XOR2_X1 port map( A1 => n4768, A2 => n14488, Z => n19178);
   U21043 : XOR2_X1 port map( A1 => n19368, A2 => n14544, Z => n19182);
   U21044 : XOR2_X1 port map( A1 => n12739, A2 => n20727, Z => n19193);
   U21045 : XOR2_X1 port map( A1 => n27362, A2 => n14574, Z => n19195);
   U21047 : XOR2_X1 port map( A1 => n19421, A2 => n20851, Z => n19202);
   U21048 : INV_X1 port map( I => n19210, ZN => n19209);
   U21049 : INV_X1 port map( I => n20602, ZN => n19208);
   U21050 : INV_X1 port map( I => n19203, ZN => n19204);
   U21051 : NOR3_X1 port map( A1 => n19205, A2 => n20602, A3 => n19204, ZN => 
                           n19207);
   U21052 : AOI22_X1 port map( A1 => n19209, A2 => n19208, B1 => n19207, B2 => 
                           n19206, ZN => n19213);
   U21053 : NAND3_X1 port map( A1 => n19211, A2 => n19210, A3 => n20602, ZN => 
                           n19212);
   U21054 : XOR2_X1 port map( A1 => n6309, A2 => n14597, Z => n19216);
   U21055 : XOR2_X1 port map( A1 => n28488, A2 => n21703, Z => n19222);
   U21056 : NAND2_X1 port map( A1 => n19225, A2 => n996, ZN => n19226);
   U21059 : XOR2_X1 port map( A1 => n23691, A2 => n19500, Z => n19327);
   U21061 : XOR2_X1 port map( A1 => n19478, A2 => n21597, Z => n19235);
   U21062 : NAND2_X1 port map( A1 => n19763, A2 => n23868, ZN => n19247);
   U21065 : XOR2_X1 port map( A1 => n14558, A2 => n19562, Z => n19242);
   U21066 : NAND2_X1 port map( A1 => n19930, A2 => n7238, ZN => n19243);
   U21067 : XOR2_X1 port map( A1 => n5653, A2 => n14581, Z => n19251);
   U21068 : XOR2_X1 port map( A1 => n19492, A2 => n19251, Z => n19252);
   U21069 : XOR2_X1 port map( A1 => n19488, A2 => n19256, Z => n19257);
   U21071 : XOR2_X1 port map( A1 => n13904, A2 => n14445, Z => n19266);
   U21072 : XOR2_X1 port map( A1 => n19366, A2 => n19267, Z => n19268);
   U21073 : INV_X1 port map( I => n16961, ZN => n19270);
   U21074 : XOR2_X1 port map( A1 => n19496, A2 => n19270, Z => n19271);
   U21076 : XOR2_X1 port map( A1 => n28464, A2 => n20692, Z => n19284);
   U21077 : XOR2_X1 port map( A1 => n7397, A2 => n7050, Z => n19286);
   U21078 : XOR2_X1 port map( A1 => n19294, A2 => n19293, Z => n19295);
   U21079 : XOR2_X1 port map( A1 => n19296, A2 => n19295, Z => n19905);
   U21082 : XOR2_X1 port map( A1 => n27374, A2 => n14622, Z => n19304);
   U21083 : XOR2_X1 port map( A1 => n8912, A2 => n19306, Z => n19307);
   U21084 : XOR2_X1 port map( A1 => n984, A2 => n19500, Z => n19316);
   U21086 : XOR2_X1 port map( A1 => n22381, A2 => n14589, Z => n19335);
   U21088 : XOR2_X1 port map( A1 => n13904, A2 => n14549, Z => n19342);
   U21090 : XOR2_X1 port map( A1 => n19430, A2 => n19368, Z => n19370);
   U21091 : XOR2_X1 port map( A1 => n14340, A2 => n19482, Z => n19369);
   U21092 : XOR2_X1 port map( A1 => n19370, A2 => n19369, Z => n19371);
   U21093 : XOR2_X1 port map( A1 => n11054, A2 => n15669, Z => n19372);
   U21094 : INV_X1 port map( I => n19377, ZN => n19378);
   U21095 : XOR2_X1 port map( A1 => n26545, A2 => n21422, Z => n19379);
   U21096 : XOR2_X1 port map( A1 => n19446, A2 => n20584, Z => n19384);
   U21097 : XOR2_X1 port map( A1 => n28464, A2 => n21679, Z => n19390);
   U21098 : XOR2_X1 port map( A1 => n19446, A2 => n21357, Z => n19401);
   U21100 : XOR2_X1 port map( A1 => n28464, A2 => n21554, Z => n19418);
   U21104 : XOR2_X1 port map( A1 => n27448, A2 => n20605, Z => n19429);
   U21105 : XOR2_X1 port map( A1 => n15126, A2 => n14506, Z => n19433);
   U21106 : XOR2_X1 port map( A1 => n7346, A2 => n20614, Z => n19436);
   U21108 : XOR2_X1 port map( A1 => n19487, A2 => n7387, Z => n19440);
   U21109 : XOR2_X1 port map( A1 => n19447, A2 => n22770, Z => n19448);
   U21110 : XOR2_X1 port map( A1 => n19540, A2 => n21141, Z => n19452);
   U21111 : XOR2_X1 port map( A1 => n26469, A2 => n14619, Z => n19454);
   U21112 : XOR2_X1 port map( A1 => n19455, A2 => n19454, Z => n19456);
   U21119 : XOR2_X1 port map( A1 => n19480, A2 => n19481, Z => n19484);
   U21121 : INV_X1 port map( I => n21085, ZN => n19495);
   U21122 : XOR2_X1 port map( A1 => n19510, A2 => n21227, Z => n19511);
   U21123 : XOR2_X1 port map( A1 => n19513, A2 => n19512, Z => n19514);
   U21124 : XOR2_X1 port map( A1 => n19516, A2 => n7368, Z => n19517);
   U21125 : XOR2_X1 port map( A1 => n19552, A2 => n27149, Z => n19539);
   U21126 : XOR2_X1 port map( A1 => n19540, A2 => n1283, Z => n19541);
   U21127 : INV_X1 port map( I => n19543, ZN => n19545);
   U21133 : XOR2_X1 port map( A1 => n26329, A2 => n21183, Z => n19607);
   U21135 : NAND2_X1 port map( A1 => n3317, A2 => n13926, ZN => n19608);
   U21136 : NAND3_X1 port map( A1 => n19824, A2 => n19823, A3 => n28378, ZN => 
                           n19610);
   U21139 : NOR2_X1 port map( A1 => n27823, A2 => n12393, ZN => n19616);
   U21141 : NAND2_X1 port map( A1 => n14343, A2 => n10978, ZN => n19619);
   U21144 : XOR2_X1 port map( A1 => n21153, A2 => n27169, Z => n19628);
   U21146 : INV_X1 port map( I => n19642, ZN => n19644);
   U21147 : NOR2_X1 port map( A1 => n23857, A2 => n13278, ZN => n19647);
   U21148 : NAND2_X1 port map( A1 => n14565, A2 => n19658, ZN => n19659);
   U21151 : INV_X1 port map( I => n19672, ZN => n19878);
   U21160 : XOR2_X1 port map( A1 => n14436, A2 => n21237, Z => n19701);
   U21163 : NOR2_X1 port map( A1 => n28377, A2 => n14304, ZN => n19722);
   U21164 : INV_X1 port map( I => n19721, ZN => n19724);
   U21165 : INV_X1 port map( I => n19722, ZN => n19723);
   U21169 : INV_X1 port map( I => n19765, ZN => n19767);
   U21173 : MUX2_X1 port map( I0 => n19813, I1 => n19812, S => n5048, Z => 
                           n19815);
   U21174 : NOR2_X1 port map( A1 => n11920, A2 => n1366, ZN => n19816);
   U21175 : NOR2_X1 port map( A1 => n19817, A2 => n20152, ZN => n20341);
   U21176 : XOR2_X1 port map( A1 => n21257, A2 => n20038, Z => n19818);
   U21181 : NOR2_X1 port map( A1 => n20110, A2 => n978, ZN => n19859);
   U21183 : INV_X1 port map( I => n19865, ZN => n19867);
   U21189 : NAND2_X1 port map( A1 => n19883, A2 => n19882, ZN => n19884);
   U21190 : XOR2_X1 port map( A1 => n14616, A2 => n21435, Z => n19886);
   U21195 : NAND2_X1 port map( A1 => n22140, A2 => n9401, ZN => n19942);
   U21197 : NOR2_X1 port map( A1 => n20194, A2 => n20291, ZN => n19958);
   U21198 : XOR2_X1 port map( A1 => n11389, A2 => n12769, Z => n19966);
   U21200 : NOR2_X1 port map( A1 => n22758, A2 => n1105, ZN => n19972);
   U21203 : XOR2_X1 port map( A1 => n20385, A2 => n22755, Z => n20007);
   U21209 : NAND3_X1 port map( A1 => n20087, A2 => n20050, A3 => n22000, ZN => 
                           n20036);
   U21213 : XOR2_X1 port map( A1 => n25361, A2 => n9678, Z => n20047);
   U21215 : NAND2_X1 port map( A1 => n10721, A2 => n20050, ZN => n20051);
   U21216 : NAND2_X1 port map( A1 => n20073, A2 => n20072, ZN => n20074);
   U21218 : XOR2_X1 port map( A1 => n20488, A2 => n14418, Z => n20076);
   U21219 : XOR2_X1 port map( A1 => n21257, A2 => n21434, Z => n20442);
   U21220 : OAI22_X1 port map( A1 => n20201, A2 => n20101, B1 => n20102, B2 => 
                           n12503, ZN => n20091);
   U21221 : NOR2_X1 port map( A1 => n20432, A2 => n20091, ZN => n20092);
   U21224 : NAND2_X1 port map( A1 => n20286, A2 => n23906, ZN => n20116);
   U21225 : XOR2_X1 port map( A1 => n20581, A2 => n20435, Z => n20119);
   U21227 : NAND2_X1 port map( A1 => n26650, A2 => n21208, ZN => n20133);
   U21229 : NAND3_X1 port map( A1 => n20133, A2 => n21325, A3 => n21327, ZN => 
                           n20135);
   U21231 : XOR2_X1 port map( A1 => n20650, A2 => n22791, Z => n20148);
   U21233 : NOR2_X1 port map( A1 => n9450, A2 => n20162, ZN => n20161);
   U21234 : NAND2_X1 port map( A1 => n20309, A2 => n9264, ZN => n20163);
   U21235 : NAND3_X1 port map( A1 => n20163, A2 => n26355, A3 => n20162, ZN => 
                           n20164);
   U21237 : NAND2_X1 port map( A1 => n20197, A2 => n13252, ZN => n20198);
   U21238 : NOR3_X1 port map( A1 => n13294, A2 => n20219, A3 => n12143, ZN => 
                           n20220);
   U21242 : XOR2_X1 port map( A1 => n26029, A2 => n21302, Z => n20241);
   U21244 : XOR2_X1 port map( A1 => n20552, A2 => n22755, Z => n20250);
   U21247 : XOR2_X1 port map( A1 => n21258, A2 => n14549, Z => n20283);
   U21248 : NAND3_X1 port map( A1 => n858, A2 => n7927, A3 => n20280, ZN => 
                           n20281);
   U21251 : INV_X1 port map( I => n20496, ZN => n20303);
   U21252 : NOR2_X1 port map( A1 => n334, A2 => n12712, ZN => n20301);
   U21253 : NAND2_X1 port map( A1 => n8300, A2 => n12712, ZN => n20298);
   U21254 : OAI22_X1 port map( A1 => n20301, A2 => n20300, B1 => n26738, B2 => 
                           n20298, ZN => n20302);
   U21255 : AOI21_X1 port map( A1 => n20303, A2 => n21772, B => n20302, ZN => 
                           n20304);
   U21256 : XOR2_X1 port map( A1 => n20550, A2 => n14550, Z => n20320);
   U21257 : INV_X1 port map( I => Key(188), ZN => n20321);
   U21260 : XOR2_X1 port map( A1 => n27396, A2 => n14638, Z => n20335);
   U21261 : OAI22_X1 port map( A1 => n20340, A2 => n11920, B1 => n3290, B2 => 
                           n20337, ZN => n20342);
   U21262 : NOR2_X1 port map( A1 => n20342, A2 => n20341, ZN => n20343);
   U21263 : XOR2_X1 port map( A1 => n27673, A2 => n28502, Z => n20347);
   U21264 : XOR2_X1 port map( A1 => n20488, A2 => n21712, Z => n20346);
   U21267 : XOR2_X1 port map( A1 => n11389, A2 => n7011, Z => n20350);
   U21268 : XOR2_X1 port map( A1 => n20452, A2 => n21597, Z => n20349);
   U21269 : XOR2_X1 port map( A1 => n13834, A2 => n21607, Z => n20352);
   U21271 : XOR2_X1 port map( A1 => n21197, A2 => n20404, Z => n20357);
   U21272 : XOR2_X1 port map( A1 => n20404, A2 => n20851, Z => n20358);
   U21274 : XOR2_X1 port map( A1 => n26884, A2 => n21256, Z => n20359);
   U21276 : XOR2_X1 port map( A1 => n21191, A2 => n11918, Z => n20362);
   U21277 : XOR2_X1 port map( A1 => n20363, A2 => n20362, Z => n20364);
   U21279 : XOR2_X1 port map( A1 => n21151, A2 => n20368, Z => n20373);
   U21280 : XOR2_X1 port map( A1 => n13585, A2 => n5082, Z => n20371);
   U21283 : OAI22_X1 port map( A1 => n21624, A2 => n21627, B1 => n21622, B2 => 
                           n14406, ZN => n20374);
   U21284 : XOR2_X1 port map( A1 => n20379, A2 => n136, Z => n20380);
   U21285 : XOR2_X1 port map( A1 => n20501, A2 => n20380, Z => n20382);
   U21286 : XOR2_X1 port map( A1 => n27396, A2 => n20908, Z => n20387);
   U21287 : NAND2_X1 port map( A1 => n28553, A2 => n27416, ZN => n20401);
   U21288 : NOR2_X1 port map( A1 => n23913, A2 => n9264, ZN => n20392);
   U21291 : XOR2_X1 port map( A1 => n20771, A2 => n14588, Z => n20394);
   U21292 : XOR2_X1 port map( A1 => n23648, A2 => n21048, Z => n20398);
   U21294 : NAND2_X1 port map( A1 => n28017, A2 => n10666, ZN => n20403);
   U21295 : XOR2_X1 port map( A1 => n20452, A2 => n7368, Z => n20406);
   U21297 : NAND2_X1 port map( A1 => n20414, A2 => n4738, ZN => n20418);
   U21298 : OAI21_X1 port map( A1 => n20416, A2 => n20415, B => n4739, ZN => 
                           n20417);
   U21299 : NAND2_X1 port map( A1 => n20418, A2 => n20417, ZN => n21426);
   U21301 : XOR2_X1 port map( A1 => n22806, A2 => n20707, Z => n20421);
   U21303 : XOR2_X1 port map( A1 => n20511, A2 => n21218, Z => n20425);
   U21304 : AOI21_X1 port map( A1 => n20739, A2 => n20781, B => n15689, ZN => 
                           n20426);
   U21305 : OAI21_X1 port map( A1 => n20781, A2 => n13188, B => n20426, ZN => 
                           n20427);
   U21308 : NOR2_X1 port map( A1 => n20691, A2 => n20696, ZN => n20465);
   U21309 : XOR2_X1 port map( A1 => n20580, A2 => n20450, Z => n21192);
   U21315 : XOR2_X1 port map( A1 => n20552, A2 => n21449, Z => n20476);
   U21316 : XOR2_X1 port map( A1 => n20477, A2 => n20476, Z => n20478);
   U21321 : INV_X1 port map( I => n14489, ZN => n20499);
   U21322 : XOR2_X1 port map( A1 => n9161, A2 => n20499, Z => n20500);
   U21323 : INV_X1 port map( I => n20733, ZN => n20504);
   U21324 : NAND2_X1 port map( A1 => n20504, A2 => n25145, ZN => n20505);
   U21326 : XOR2_X1 port map( A1 => n27087, A2 => n14479, Z => n20515);
   U21328 : XOR2_X1 port map( A1 => n13808, A2 => n21517, Z => n20525);
   U21330 : NAND3_X1 port map( A1 => n14341, A2 => n20972, A3 => n20561, ZN => 
                           n20562);
   U21331 : XOR2_X1 port map( A1 => n14144, A2 => n20566, Z => n20567);
   U21333 : INV_X1 port map( I => n20570, ZN => n20572);
   U21334 : OAI22_X1 port map( A1 => n20574, A2 => n20573, B1 => n20572, B2 => 
                           n20571, ZN => n20575);
   U21336 : XOR2_X1 port map( A1 => n21434, A2 => n13746, Z => n20578);
   U21337 : INV_X1 port map( I => n20584, ZN => n20585);
   U21338 : NOR2_X1 port map( A1 => n20685, A2 => n25324, ZN => n20592);
   U21340 : NAND2_X1 port map( A1 => n20667, A2 => n13234, ZN => n20595);
   U21341 : NAND3_X1 port map( A1 => n14750, A2 => n22764, A3 => n7319, ZN => 
                           n20601);
   U21342 : NAND2_X1 port map( A1 => n20608, A2 => n22764, ZN => n20600);
   U21345 : OAI21_X1 port map( A1 => n8935, A2 => n20609, B => n20608, ZN => 
                           n20610);
   U21346 : OAI21_X1 port map( A1 => n20618, A2 => n939, B => n20623, ZN => 
                           n20612);
   U21347 : INV_X1 port map( I => n20618, ZN => n20628);
   U21348 : NAND2_X1 port map( A1 => n939, A2 => n20623, ZN => n20615);
   U21349 : AOI21_X1 port map( A1 => n14146, A2 => n20625, B => n20624, ZN => 
                           n20629);
   U21350 : OAI22_X1 port map( A1 => n20629, A2 => n24597, B1 => n20627, B2 => 
                           n20628, ZN => n20630);
   U21351 : XOR2_X1 port map( A1 => n20630, A2 => n14549, Z => Ciphertext(11));
   U21353 : OR2_X1 port map( A1 => n20739, A2 => n20633, Z => n20636);
   U21354 : NAND2_X1 port map( A1 => n20633, A2 => n20786, ZN => n20634);
   U21355 : NAND3_X1 port map( A1 => n20637, A2 => n13188, A3 => n20736, ZN => 
                           n20638);
   U21356 : NAND2_X1 port map( A1 => n20656, A2 => n848, ZN => n20649);
   U21357 : NAND3_X1 port map( A1 => n20663, A2 => n848, A3 => n20658, ZN => 
                           n20648);
   U21358 : INV_X1 port map( I => n4934, ZN => n20664);
   U21359 : INV_X1 port map( I => n14581, ZN => n20666);
   U21364 : AOI21_X1 port map( A1 => n20688, A2 => n13234, B => n20687, ZN => 
                           n20689);
   U21365 : XOR2_X1 port map( A1 => n20689, A2 => n1290, Z => Ciphertext(23));
   U21367 : NAND2_X1 port map( A1 => n20696, A2 => n20695, ZN => n20700);
   U21369 : XOR2_X1 port map( A1 => n20767, A2 => n21077, Z => n20719);
   U21370 : XOR2_X1 port map( A1 => n20720, A2 => n20719, Z => n20721);
   U21372 : NAND2_X1 port map( A1 => n24575, A2 => n20736, ZN => n20737);
   U21373 : NOR2_X1 port map( A1 => n25325, A2 => n20751, ZN => n20740);
   U21374 : XOR2_X1 port map( A1 => n20742, A2 => n22890, Z => Ciphertext(31));
   U21376 : NAND2_X1 port map( A1 => n20899, A2 => n20894, ZN => n20758);
   U21377 : XOR2_X1 port map( A1 => n20767, A2 => n20766, Z => n20768);
   U21378 : XOR2_X1 port map( A1 => n20773, A2 => n7284, Z => n20774);
   U21379 : XOR2_X1 port map( A1 => n27423, A2 => n21482, Z => n20775);
   U21380 : NAND2_X1 port map( A1 => n14647, A2 => n20786, ZN => n20784);
   U21381 : NOR2_X1 port map( A1 => n24575, A2 => n20786, ZN => n20788);
   U21383 : NAND2_X1 port map( A1 => n20791, A2 => n10477, ZN => n20792);
   U21388 : OAI21_X1 port map( A1 => n28213, A2 => n25360, B => n20833, ZN => 
                           n20824);
   U21391 : NAND2_X1 port map( A1 => n20979, A2 => n20887, ZN => n20812);
   U21392 : NAND3_X1 port map( A1 => n11319, A2 => n11318, A3 => n20847, ZN => 
                           n20822);
   U21394 : NAND2_X1 port map( A1 => n20822, A2 => n20843, ZN => n20823);
   U21395 : AOI21_X1 port map( A1 => n20824, A2 => n20827, B => n20823, ZN => 
                           n20825);
   U21396 : XOR2_X1 port map( A1 => n20825, A2 => n924, Z => Ciphertext(42));
   U21397 : NAND2_X1 port map( A1 => n20842, A2 => n20827, ZN => n20828);
   U21398 : INV_X1 port map( I => n14488, ZN => n21243);
   U21399 : XOR2_X1 port map( A1 => n20829, A2 => n21243, Z => Ciphertext(43));
   U21402 : OR2_X1 port map( A1 => n20833, A2 => n20827, Z => n20840);
   U21403 : NAND3_X1 port map( A1 => n20846, A2 => n20837, A3 => n20842, ZN => 
                           n20838);
   U21404 : XOR2_X1 port map( A1 => n20845, A2 => n21422, Z => Ciphertext(46));
   U21406 : NAND2_X1 port map( A1 => n20857, A2 => n20899, ZN => n20858);
   U21407 : NOR2_X1 port map( A1 => n20868, A2 => n20862, ZN => n20863);
   U21408 : NAND2_X1 port map( A1 => n20867, A2 => n20866, ZN => n20869);
   U21409 : NAND2_X1 port map( A1 => n20888, A2 => n12598, ZN => n20889);
   U21410 : NAND2_X1 port map( A1 => n21029, A2 => n1083, ZN => n20892);
   U21413 : NAND3_X1 port map( A1 => n22803, A2 => n20910, A3 => n20911, ZN => 
                           n20905);
   U21414 : NAND2_X1 port map( A1 => n20913, A2 => n1071, ZN => n20903);
   U21415 : XOR2_X1 port map( A1 => n20907, A2 => n20906, Z => Ciphertext(55));
   U21419 : NAND2_X1 port map( A1 => n15545, A2 => n10558, ZN => n20922);
   U21422 : NAND3_X1 port map( A1 => n20938, A2 => n25610, A3 => n10639, ZN => 
                           n20939);
   U21423 : XOR2_X1 port map( A1 => n20943, A2 => n23657, Z => Ciphertext(60));
   U21424 : OAI21_X1 port map( A1 => n22738, A2 => n23088, B => n20944, ZN => 
                           n20946);
   U21425 : XOR2_X1 port map( A1 => n20947, A2 => n14619, Z => Ciphertext(61));
   U21428 : NAND2_X1 port map( A1 => n20958, A2 => n20957, ZN => n20959);
   U21429 : NAND2_X1 port map( A1 => n20960, A2 => n20959, ZN => n20962);
   U21430 : XOR2_X1 port map( A1 => n20962, A2 => n20961, Z => Ciphertext(64));
   U21431 : AOI21_X1 port map( A1 => n20964, A2 => n20963, B => n4604, ZN => 
                           n20966);
   U21440 : NAND2_X1 port map( A1 => n21040, A2 => n10635, ZN => n21023);
   U21442 : NOR3_X1 port map( A1 => n21050, A2 => n21030, A3 => n21040, ZN => 
                           n21031);
   U21443 : XOR2_X1 port map( A1 => n21034, A2 => n1316, Z => Ciphertext(78));
   U21446 : AOI21_X1 port map( A1 => n27392, A2 => n10635, B => n22797, ZN => 
                           n21053);
   U21448 : NAND2_X1 port map( A1 => n21070, A2 => n7904, ZN => n21071);
   U21450 : NOR2_X1 port map( A1 => n13476, A2 => n21078, ZN => n21073);
   U21451 : INV_X1 port map( I => n14600, ZN => n21075);
   U21456 : NAND3_X1 port map( A1 => n26462, A2 => n4277, A3 => n13021, ZN => 
                           n21105);
   U21460 : OAI21_X1 port map( A1 => n23976, A2 => n13472, B => n21124, ZN => 
                           n21125);
   U21461 : AOI22_X1 port map( A1 => n21127, A2 => n21116, B1 => n21126, B2 => 
                           n21125, ZN => n21128);
   U21462 : XOR2_X1 port map( A1 => n21128, A2 => n6287, Z => Ciphertext(101));
   U21463 : NAND3_X1 port map( A1 => n13447, A2 => n26554, A3 => n21275, ZN => 
                           n21131);
   U21464 : NOR2_X1 port map( A1 => n26773, A2 => n14260, ZN => n21134);
   U21466 : XOR2_X1 port map( A1 => n21145, A2 => n21144, Z => n21147);
   U21467 : XOR2_X1 port map( A1 => n15680, A2 => n21435, Z => n21155);
   U21469 : XOR2_X1 port map( A1 => n21182, A2 => n21557, Z => n21184);
   U21470 : XOR2_X1 port map( A1 => n4137, A2 => n21185, Z => n21186);
   U21471 : XOR2_X1 port map( A1 => n21189, A2 => n21188, Z => n21195);
   U21472 : XNOR2_X1 port map( A1 => n21190, A2 => n21191, ZN => n21193);
   U21473 : XOR2_X1 port map( A1 => n21192, A2 => n21193, Z => n21194);
   U21474 : XOR2_X1 port map( A1 => n21198, A2 => n27423, Z => n21200);
   U21475 : OAI21_X1 port map( A1 => n13791, A2 => n21202, B => n14529, ZN => 
                           n21203);
   U21477 : NOR2_X1 port map( A1 => n25307, A2 => n21213, ZN => n21214);
   U21478 : XOR2_X1 port map( A1 => n21219, A2 => n21218, Z => Ciphertext(110))
                           ;
   U21479 : MUX2_X1 port map( I0 => n21457, I1 => n13791, S => n21441, Z => 
                           n21232);
   U21480 : NAND2_X1 port map( A1 => n21232, A2 => n13424, ZN => n21233);
   U21481 : NAND2_X2 port map( A1 => n21234, A2 => n21233, ZN => n21292);
   U21484 : XOR2_X1 port map( A1 => n21243, A2 => n12382, Z => n21244);
   U21486 : XOR2_X1 port map( A1 => n21249, A2 => n5082, Z => n21250);
   U21487 : XOR2_X1 port map( A1 => n21251, A2 => n21250, Z => n21252);
   U21488 : XOR2_X1 port map( A1 => n21253, A2 => n21252, Z => n21266);
   U21489 : XOR2_X1 port map( A1 => n21261, A2 => n1097, Z => n21264);
   U21490 : XOR2_X1 port map( A1 => n21264, A2 => n21263, Z => n21265);
   U21491 : INV_X1 port map( I => n21500, ZN => n21463);
   U21492 : NOR2_X1 port map( A1 => n14409, A2 => n9378, ZN => n21272);
   U21493 : NAND2_X1 port map( A1 => n15375, A2 => n22824, ZN => n21280);
   U21494 : XOR2_X1 port map( A1 => n21285, A2 => n1283, Z => Ciphertext(117));
   U21495 : XOR2_X1 port map( A1 => n21289, A2 => n21288, Z => Ciphertext(118))
                           ;
   U21496 : XOR2_X1 port map( A1 => n21294, A2 => n14616, Z => Ciphertext(119))
                           ;
   U21497 : MUX2_X1 port map( I0 => n5519, I1 => n21395, S => n21445, Z => 
                           n21297);
   U21498 : XOR2_X1 port map( A1 => n21305, A2 => n21304, Z => n21307);
   U21499 : XOR2_X1 port map( A1 => n21307, A2 => n21306, Z => n21308);
   U21501 : NAND3_X1 port map( A1 => n14525, A2 => n27442, A3 => n21464, ZN => 
                           n21322);
   U21508 : INV_X1 port map( I => n14652, ZN => n21363);
   U21509 : INV_X1 port map( I => n14596, ZN => n21570);
   U21511 : XOR2_X1 port map( A1 => n5446, A2 => n21707, Z => n21379);
   U21512 : XOR2_X1 port map( A1 => n21380, A2 => n21379, Z => n21381);
   U21513 : XOR2_X1 port map( A1 => n21432, A2 => n21384, Z => n21385);
   U21515 : NAND3_X1 port map( A1 => n13756, A2 => n7199, A3 => n21415, ZN => 
                           n21399);
   U21516 : NOR2_X1 port map( A1 => n21445, A2 => n21395, ZN => n21396);
   U21517 : NAND3_X1 port map( A1 => n21415, A2 => n21405, A3 => n21413, ZN => 
                           n21398);
   U21518 : XOR2_X1 port map( A1 => n21401, A2 => n14555, Z => Ciphertext(126))
                           ;
   U21519 : NOR2_X1 port map( A1 => n7199, A2 => n21408, ZN => n21403);
   U21521 : XOR2_X1 port map( A1 => n21404, A2 => n14643, Z => Ciphertext(127))
                           ;
   U21522 : AOI21_X1 port map( A1 => n22794, A2 => n21413, B => n21412, ZN => 
                           n21414);
   U21524 : XOR2_X1 port map( A1 => n26329, A2 => n21419, Z => n21420);
   U21526 : AOI21_X1 port map( A1 => n13987, A2 => n7944, B => n23579, ZN => 
                           n21452);
   U21527 : INV_X1 port map( I => n21547, ZN => n21621);
   U21529 : NAND2_X1 port map( A1 => n21460, A2 => n21477, ZN => n21471);
   U21532 : INV_X1 port map( I => n21481, ZN => n21468);
   U21533 : NAND3_X1 port map( A1 => n21473, A2 => n694, A3 => n21468, ZN => 
                           n21469);
   U21537 : NOR2_X1 port map( A1 => n21481, A2 => n21484, ZN => n21488);
   U21539 : OAI21_X1 port map( A1 => n21485, A2 => n21484, B => n21483, ZN => 
                           n21491);
   U21540 : OAI21_X1 port map( A1 => n21489, A2 => n21488, B => n21487, ZN => 
                           n21490);
   U21543 : NAND3_X1 port map( A1 => n7941, A2 => n21499, A3 => n21498, ZN => 
                           n21504);
   U21544 : OAI21_X1 port map( A1 => n21531, A2 => n770, B => n21528, ZN => 
                           n21516);
   U21545 : NAND2_X1 port map( A1 => n21531, A2 => n770, ZN => n21519);
   U21547 : OAI21_X1 port map( A1 => n27389, A2 => n21534, B => n21531, ZN => 
                           n21527);
   U21548 : NOR2_X1 port map( A1 => n21668, A2 => n21539, ZN => n21540);
   U21549 : INV_X1 port map( I => n21702, ZN => n21542);
   U21550 : NAND2_X1 port map( A1 => n21549, A2 => n11490, ZN => n21550);
   U21556 : INV_X1 port map( I => n5721, ZN => n21690);
   U21560 : AOI21_X1 port map( A1 => n22848, A2 => n6181, B => n21656, ZN => 
                           n21658);
   U21562 : MUX2_X1 port map( I0 => n21667, I1 => n21666, S => n5675, Z => 
                           n21670);
   U21564 : OAI21_X1 port map( A1 => n721, A2 => n21685, B => n25314, ZN => 
                           n21680);
   U21566 : INV_X1 port map( I => n21707, ZN => n21708);
   U770 : INV_X2 port map( I => n12834, ZN => n17515);
   U12416 : INV_X4 port map( I => n27905, ZN => n15667);
   U731 : NOR2_X2 port map( A1 => n1033, A2 => n17519, ZN => n17321);
   U18272 : OAI21_X2 port map( A1 => n15815, A2 => n10643, B => n23134, ZN => 
                           n13203);
   U4282 : NOR2_X2 port map( A1 => n17975, A2 => n23577, ZN => n13943);
   U540 : INV_X2 port map( I => n643, ZN => n18602);
   U7631 : NOR2_X2 port map( A1 => n14027, A2 => n17702, ZN => n18062);
   U1568 : NAND2_X2 port map( A1 => n16280, A2 => n21787, ZN => n16186);
   U6389 : NAND2_X2 port map( A1 => n8576, A2 => n7791, ZN => n18439);
   U132 : INV_X4 port map( I => n21578, ZN => n13432);
   U4778 : INV_X4 port map( I => n18344, ZN => n881);
   U7624 : INV_X2 port map( I => n2437, ZN => n2436);
   U639 : INV_X4 port map( I => n713, ZN => n1203);
   U517 : INV_X2 port map( I => n12221, ZN => n14308);
   U7015 : INV_X2 port map( I => n10444, ZN => n7341);
   U7094 : AOI21_X2 port map( A1 => n14838, A2 => n858, B => n7796, ZN => n7795
                           );
   U4213 : INV_X2 port map( I => n21295, ZN => n14281);
   U718 : INV_X2 port map( I => n17193, ZN => n17307);
   U882 : INV_X4 port map( I => n14906, ZN => n13211);
   U4927 : NOR2_X2 port map( A1 => n15486, A2 => n18940, ZN => n19026);
   U5337 : OAI21_X2 port map( A1 => n12668, A2 => n16561, B => n16654, ZN => 
                           n8207);
   U4006 : INV_X2 port map( I => n17607, ZN => n12676);
   U888 : INV_X4 port map( I => n13025, ZN => n1048);
   U345 : INV_X2 port map( I => n14302, ZN => n19801);
   U4482 : BUF_X2 port map( I => n17336, Z => n7361);
   U6950 : NOR2_X2 port map( A1 => n26684, A2 => n15627, ZN => n12024);
   U102 : INV_X2 port map( I => n10605, ZN => n21729);
   U5468 : NAND2_X2 port map( A1 => n13924, A2 => n20288, ZN => n6285);
   U4533 : NAND2_X2 port map( A1 => n25629, A2 => n22767, ZN => n20809);
   U8043 : OAI21_X2 port map( A1 => n5382, A2 => n16564, B => n434, ZN => 
                           n12337);
   U9748 : AOI22_X2 port map( A1 => n7821, A2 => n25576, B1 => n6592, B2 => 
                           n7822, ZN => n4469);
   U597 : NAND2_X2 port map( A1 => n6435, A2 => n17683, ZN => n17715);
   U5044 : AOI21_X2 port map( A1 => n16481, A2 => n15107, B => n14965, ZN => 
                           n14964);
   U854 : NAND2_X2 port map( A1 => n16679, A2 => n6763, ZN => n6939);
   U717 : INV_X2 port map( I => n10046, ZN => n1038);
   U30 : INV_X2 port map( I => n13987, ZN => n13986);
   U343 : INV_X4 port map( I => n8968, ZN => n1127);
   U616 : NAND2_X2 port map( A1 => n443, A2 => n17984, ZN => n12913);
   U518 : INV_X2 port map( I => n18654, ZN => n18741);
   U946 : INV_X2 port map( I => n15342, ZN => n840);
   U1281 : NAND2_X2 port map( A1 => n17482, A2 => n17483, ZN => n8940);
   U55 : NAND2_X2 port map( A1 => n11515, A2 => n7645, ZN => n21638);
   U526 : NOR2_X2 port map( A1 => n11919, A2 => n18613, ZN => n18470);
   U364 : INV_X2 port map( I => n24275, ZN => n19444);
   U45 : NAND3_X2 port map( A1 => n7105, A2 => n7537, A3 => n10394, ZN => n9458
                           );
   U1270 : INV_X1 port map( I => n14748, ZN => n14142);
   U5008 : NAND2_X2 port map( A1 => n25926, A2 => n17969, ZN => n17651);
   U4545 : NAND3_X2 port map( A1 => n20056, A2 => n15369, A3 => n20071, ZN => 
                           n15368);
   U886 : INV_X4 port map( I => n16562, ZN => n16654);
   U6073 : OAI21_X2 port map( A1 => n10686, A2 => n27674, B => n20016, ZN => 
                           n1914);
   U10223 : OAI21_X2 port map( A1 => n2118, A2 => n26853, B => n2116, ZN => 
                           n16542);
   U370 : NAND3_X2 port map( A1 => n12807, A2 => n18997, A3 => n12806, ZN => 
                           n19521);
   U15515 : OR2_X1 port map( A1 => n6286, A2 => n6264, Z => n6284);
   U18553 : INV_X1 port map( I => n15917, ZN => n16307);
   U7024 : NAND2_X2 port map( A1 => n20728, A2 => n28553, ZN => n20733);
   U347 : INV_X2 port map( I => n19194, ZN => n19529);
   U4842 : BUF_X2 port map( I => n15869, Z => n15998);
   U279 : NAND2_X2 port map( A1 => n8073, A2 => n9583, ZN => n10488);
   U6443 : OAI21_X2 port map( A1 => n14312, A2 => n17987, B => n12611, ZN => 
                           n6170);
   U5658 : AOI21_X2 port map( A1 => n23002, A2 => n17984, B => n12590, ZN => 
                           n14312);
   U6565 : OAI21_X2 port map( A1 => n15504, A2 => n10942, B => n7073, ZN => 
                           n12445);
   U870 : NAND2_X2 port map( A1 => n912, A2 => n24167, ZN => n2760);
   U8277 : NOR2_X2 port map( A1 => n7270, A2 => n13731, ZN => n16125);
   U1750 : NAND2_X2 port map( A1 => n9891, A2 => n5244, ZN => n53);
   U5429 : INV_X2 port map( I => n21667, ZN => n5673);
   U3690 : INV_X2 port map( I => n11024, ZN => n14989);
   U4228 : AOI21_X2 port map( A1 => n20496, A2 => n20495, B => n20494, ZN => 
                           n21235);
   U5344 : NAND2_X2 port map( A1 => n9314, A2 => n14906, ZN => n16673);
   U5702 : INV_X2 port map( I => n2901, ZN => n3875);
   U338 : INV_X2 port map( I => n7004, ZN => n19630);
   U7994 : NAND2_X2 port map( A1 => n8519, A2 => n8518, ZN => n9276);
   U3738 : NOR2_X2 port map( A1 => n13853, A2 => n20237, ZN => n20239);
   U7187 : OAI21_X2 port map( A1 => n11315, A2 => n11314, B => n34, ZN => 
                           n11313);
   U934 : NAND2_X2 port map( A1 => n16280, A2 => n16278, ZN => n16284);
   U461 : NAND2_X2 port map( A1 => n15598, A2 => n15600, ZN => n19101);
   U283 : NOR2_X2 port map( A1 => n3954, A2 => n19781, ZN => n8048);
   U892 : NAND2_X2 port map( A1 => n13402, A2 => n15794, ZN => n12726);
   U5017 : INV_X2 port map( I => n7156, ZN => n829);
   U813 : AOI21_X2 port map( A1 => n16724, A2 => n16723, B => n14264, ZN => 
                           n16727);
   U335 : INV_X2 port map( I => n606, ZN => n19866);
   U6701 : AOI21_X2 port map( A1 => n6270, A2 => n7759, B => n11505, ZN => 
                           n6269);
   U5754 : NAND2_X2 port map( A1 => n7430, A2 => n913, ZN => n6270);
   U5110 : INV_X2 port map( I => n15021, ZN => n1085);
   U4574 : BUF_X2 port map( I => n19593, Z => n19731);
   U196 : INV_X2 port map( I => n20142, ZN => n14153);
   U954 : BUF_X4 port map( I => n15758, Z => n16339);
   U8254 : INV_X4 port map( I => n16086, ZN => n1267);
   U785 : INV_X4 port map( I => n17497, ZN => n8180);
   U4887 : OAI21_X2 port map( A1 => n20142, A2 => n5047, B => n1932, ZN => 
                           n20207);
   U10 : INV_X2 port map( I => n12784, ZN => n12508);
   U443 : NAND2_X2 port map( A1 => n18548, A2 => n10083, ZN => n2728);
   U5137 : INV_X4 port map( I => n15067, ZN => n810);
   U327 : BUF_X4 port map( I => n13121, Z => n13110);
   U4362 : AOI21_X2 port map( A1 => n23125, A2 => n1383, B => n5994, ZN => 
                           n5993);
   U222 : NAND2_X2 port map( A1 => n6855, A2 => n1933, ZN => n8135);
   U4490 : NAND2_X2 port map( A1 => n1413, A2 => n12092, ZN => n16608);
   U357 : NAND2_X2 port map( A1 => n979, A2 => n2462, ZN => n2466);
   U4144 : OR2_X1 port map( A1 => n2232, A2 => n2447, Z => n11156);
   U5338 : INV_X2 port map( I => n16572, ZN => n16574);
   U5083 : INV_X2 port map( I => n15923, ZN => n16134);
   U1125 : INV_X2 port map( I => n2284, ZN => n15199);
   U9265 : NAND3_X2 port map( A1 => n12452, A2 => n12451, A3 => n27941, ZN => 
                           n12255);
   U16769 : INV_X2 port map( I => n15258, ZN => n20817);
   U9995 : OAI21_X2 port map( A1 => n12499, A2 => n17321, B => n636, ZN => 
                           n2757);
   U7843 : NAND2_X2 port map( A1 => n17321, A2 => n17431, ZN => n4875);
   U6211 : INV_X2 port map( I => n19784, ZN => n19697);
   U6647 : NAND2_X2 port map( A1 => n16246, A2 => n16428, ZN => n14853);
   U4627 : NOR2_X2 port map( A1 => n6293, A2 => n17460, ZN => n17464);
   U1488 : NAND2_X2 port map( A1 => n7180, A2 => n26814, ZN => n5917);
   U15198 : NOR2_X2 port map( A1 => n855, A2 => n22735, ZN => n13271);
   U7113 : OAI21_X2 port map( A1 => n7935, A2 => n13315, B => n23253, ZN => 
                           n7934);
   U9017 : NAND2_X2 port map( A1 => n464, A2 => n14790, ZN => n12749);
   U5335 : OAI21_X2 port map( A1 => n6077, A2 => n11342, B => n7759, ZN => 
                           n11341);
   U735 : NOR2_X2 port map( A1 => n11113, A2 => n17318, ZN => n17163);
   U4392 : NAND2_X2 port map( A1 => n13578, A2 => n27347, ZN => n10436);
   U826 : NOR2_X2 port map( A1 => n16572, A2 => n7378, ZN => n14618);
   U4197 : NOR2_X2 port map( A1 => n21026, A2 => n21025, ZN => n12056);
   U344 : INV_X2 port map( I => n2458, ZN => n12863);
   U10353 : INV_X4 port map( I => n9261, ZN => n2976);
   U19042 : INV_X1 port map( I => n13274, ZN => n16287);
   U4563 : INV_X2 port map( I => n1127, ZN => n8952);
   U8131 : INV_X4 port map( I => n16731, ZN => n1257);
   U9 : INV_X2 port map( I => n20911, ZN => n1071);
   U12097 : INV_X4 port map( I => n2654, ZN => n16220);
   U4280 : NAND2_X2 port map( A1 => n12371, A2 => n9328, ZN => n13122);
   U14301 : NAND2_X2 port map( A1 => n20428, A2 => n20427, ZN => n4860);
   U7928 : INV_X4 port map( I => n22865, ZN => n4715);
   U889 : INV_X2 port map( I => n16567, ZN => n1052);
   U6426 : AOI22_X2 port map( A1 => n12144, A2 => n17830, B1 => n100, B2 => 
                           n18101, ZN => n5125);
   U9759 : AOI21_X2 port map( A1 => n17762, A2 => n5826, B => n6109, ZN => 
                           n5825);
   U494 : OAI21_X2 port map( A1 => n24666, A2 => n18475, B => n6512, ZN => 
                           n7484);
   U5063 : NAND2_X2 port map( A1 => n6480, A2 => n16301, ZN => n6479);
   U4781 : INV_X2 port map( I => n18110, ZN => n1198);
   U4084 : OR2_X1 port map( A1 => n13693, A2 => n15359, Z => n17214);
   U476 : AOI21_X2 port map( A1 => n18716, A2 => n18717, B => n1014, ZN => 
                           n11242);
   U10600 : BUF_X2 port map( I => n13833, Z => n7270);
   U16217 : NAND2_X1 port map( A1 => n8287, A2 => n16124, ZN => n8286);
   U339 : INV_X2 port map( I => n8824, ZN => n12941);
   U6377 : NAND2_X2 port map( A1 => n18774, A2 => n14648, ZN => n18624);
   U57 : OAI21_X2 port map( A1 => n8767, A2 => n9134, B => n3299, ZN => n8766);
   U8394 : BUF_X2 port map( I => Key(178), Z => n14491);
   U185 : NAND2_X2 port map( A1 => n10681, A2 => n10436, ZN => n11880);
   U8693 : BUF_X2 port map( I => n20631, Z => n21720);
   U15134 : INV_X1 port map( I => n1835, ZN => n5967);
   U4878 : INV_X2 port map( I => n13308, ZN => n8757);
   U148 : NOR2_X2 port map( A1 => n11544, A2 => n11543, ZN => n13253);
   U5292 : INV_X2 port map( I => n7269, ZN => n14861);
   U1324 : INV_X2 port map( I => n10126, ZN => n11263);
   U4986 : OAI21_X2 port map( A1 => n17785, A2 => n10823, B => n17958, ZN => 
                           n9062);
   U6410 : INV_X2 port map( I => n15366, ZN => n1189);
   U7 : INV_X2 port map( I => n4860, ZN => n8388);
   U1176 : OAI21_X1 port map( A1 => n12364, A2 => n20290, B => n7933, ZN => 
                           n7932);
   U4791 : NAND3_X2 port map( A1 => n17864, A2 => n23564, A3 => n739, ZN => 
                           n17865);
   U4606 : OAI21_X2 port map( A1 => n9331, A2 => n24586, B => n11391, ZN => 
                           n9328);
   U4806 : INV_X2 port map( I => n17919, ZN => n763);
   U4967 : NAND2_X2 port map( A1 => n18344, A2 => n13564, ZN => n12820);
   U4463 : INV_X2 port map( I => n7834, ZN => n1207);
   U5709 : INV_X2 port map( I => n15317, ZN => n17363);
   U63 : INV_X1 port map( I => n27460, ZN => n21681);
   U10677 : BUF_X2 port map( I => Key(99), Z => n14650);
   U830 : NOR2_X2 port map( A1 => n4556, A2 => n4555, ZN => n15751);
   U18028 : OAI21_X2 port map( A1 => n16139, A2 => n14857, B => n16138, ZN => 
                           n11461);
   U961 : INV_X2 port map( I => n8406, ZN => n16062);
   U7964 : AOI21_X2 port map( A1 => n11605, A2 => n11604, B => n16559, ZN => 
                           n1373);
   U6798 : OAI21_X2 port map( A1 => n16140, A2 => n796, B => n15930, ZN => 
                           n13362);
   U951 : NAND2_X2 port map( A1 => n4485, A2 => n25266, ZN => n15358);
   U15897 : INV_X1 port map( I => n21486, ZN => n21489);
   U4651 : OAI21_X2 port map( A1 => n838, A2 => n26371, B => n15358, ZN => 
                           n15973);
   U4053 : OR2_X1 port map( A1 => n735, A2 => n15478, Z => n7895);
   U655 : INV_X2 port map( I => n2910, ZN => n11967);
   U6849 : BUF_X2 port map( I => n13209, Z => n4751);
   U10517 : NOR2_X1 port map( A1 => n16125, A2 => n15995, ZN => n8287);
   U20472 : INV_X2 port map( I => n16266, ZN => n15809);
   U4796 : INV_X1 port map( I => n17894, ZN => n828);
   U18038 : OAI21_X2 port map( A1 => n15810, A2 => n15811, B => n6315, ZN => 
                           n13102);
   U4403 : OAI21_X2 port map( A1 => n11516, A2 => n19652, B => n19800, ZN => 
                           n9453);
   U5356 : INV_X4 port map( I => n4462, ZN => n4281);
   U7929 : BUF_X2 port map( I => n14844, Z => n1701);
   U9213 : NOR2_X2 port map( A1 => n11445, A2 => n9873, ZN => n5560);
   U6503 : NAND2_X2 port map( A1 => n7524, A2 => n17226, ZN => n2324);
   U4621 : INV_X2 port map( I => n14548, ZN => n7834);
   U5721 : INV_X2 port map( I => n5506, ZN => n15317);
   U10607 : BUF_X2 port map( I => n15872, Z => n16130);
   U10669 : CLKBUF_X2 port map( I => Key(71), Z => n14597);
   U549 : INV_X4 port map( I => n13538, ZN => n1010);
   U5389 : NOR2_X2 port map( A1 => n6315, A2 => n16266, ZN => n5744);
   U2803 : OR2_X2 port map( A1 => n564, A2 => n6886, Z => n16122);
   U10541 : NOR2_X2 port map( A1 => n4750, A2 => n6647, ZN => n4881);
   U12030 : INV_X2 port map( I => n2544, ZN => n2670);
   U9926 : NAND2_X1 port map( A1 => n15112, A2 => n17441, ZN => n15111);
   U5169 : INV_X2 port map( I => n26623, ZN => n13926);
   U18632 : OAI22_X2 port map( A1 => n14035, A2 => n10823, B1 => n24003, B2 => 
                           n14034, ZN => n17960);
   U5764 : NOR2_X2 port map( A1 => n8157, A2 => n8156, ZN => n12884);
   U18033 : NAND2_X1 port map( A1 => n12483, A2 => n26039, ZN => n12214);
   U8065 : NAND2_X2 port map( A1 => n16647, A2 => n16681, ZN => n9889);
   U11927 : NOR2_X2 port map( A1 => n795, A2 => n16273, ZN => n12535);
   U13758 : OAI21_X2 port map( A1 => n18379, A2 => n4158, B => n881, ZN => 
                           n6732);
   U6212 : NAND2_X2 port map( A1 => n4443, A2 => n4442, ZN => n11551);
   U6738 : NAND2_X2 port map( A1 => n6239, A2 => n1865, ZN => n5197);
   U5647 : NAND2_X2 port map( A1 => n4104, A2 => n4103, ZN => n4100);
   U1529 : AOI21_X2 port map( A1 => n12503, A2 => n20287, B => n6801, ZN => 
                           n10329);
   U8032 : AOI21_X2 port map( A1 => n9482, A2 => n16733, B => n9202, ZN => 
                           n7755);
   U15947 : INV_X1 port map( I => n7182, ZN => n19702);
   U5628 : INV_X4 port map( I => n13564, ZN => n4158);
   U4569 : INV_X2 port map( I => n14391, ZN => n12395);
   U8984 : NAND2_X2 port map( A1 => n2553, A2 => n12431, ZN => n13651);
   U6818 : INV_X1 port map( I => n561, ZN => n1059);
   U871 : BUF_X4 port map( I => n16538, Z => n145);
   U6687 : NOR3_X2 port map( A1 => n23719, A2 => n22542, A3 => n25772, ZN => 
                           n9753);
   U9387 : INV_X2 port map( I => n9073, ZN => n11602);
   U524 : INV_X2 port map( I => n18454, ZN => n3554);
   U11963 : INV_X4 port map( I => n2525, ZN => n5931);
   U5410 : INV_X4 port map( I => n15822, ZN => n799);
   U8380 : BUF_X2 port map( I => Key(141), Z => n14638);
   U4642 : NAND2_X2 port map( A1 => n16654, A2 => n2391, ZN => n16656);
   U5803 : INV_X2 port map( I => n15929, ZN => n8620);
   U18256 : AOI22_X2 port map( A1 => n16412, A2 => n16496, B1 => n23048, B2 => 
                           n16611, ZN => n14841);
   U2493 : BUF_X4 port map( I => n23083, Z => n891);
   U460 : INV_X4 port map( I => n19006, ZN => n18956);
   U6795 : NAND2_X2 port map( A1 => n9970, A2 => n9969, ZN => n4954);
   U679 : NOR2_X2 port map( A1 => n4805, A2 => n4803, ZN => n5425);
   U10988 : INV_X2 port map( I => n2277, ZN => n14639);
   U19199 : INV_X2 port map( I => n12125, ZN => n12528);
   U15060 : NAND2_X2 port map( A1 => n27878, A2 => n574, ZN => n15969);
   U10229 : NOR2_X1 port map( A1 => n2301, A2 => n2300, ZN => n2299);
   U7958 : OAI22_X2 port map( A1 => n16430, A2 => n25973, B1 => n24183, B2 => 
                           n1802, ZN => n15650);
   U5325 : NAND2_X2 port map( A1 => n8915, A2 => n8916, ZN => n8846);
   U9164 : INV_X1 port map( I => n19850, ZN => n19681);
   U7792 : AOI21_X2 port map( A1 => n7016, A2 => n5416, B => n15515, ZN => 
                           n13503);
   U8965 : OAI21_X2 port map( A1 => n19601, A2 => n19600, B => n8145, ZN => 
                           n19602);
   U18557 : INV_X2 port map( I => n16711, ZN => n11505);
   U8354 : BUF_X2 port map( I => Key(55), Z => n14622);
   U6439 : NAND2_X1 port map( A1 => n12983, A2 => n21768, ZN => n3141);
   U6872 : BUF_X2 port map( I => Key(128), Z => n14619);
   U7316 : INV_X4 port map( I => n12256, ZN => n977);
   U19450 : NAND3_X2 port map( A1 => n731, A2 => n1090, A3 => n22737, ZN => 
                           n12849);
   U14112 : INV_X2 port map( I => n4610, ZN => n17822);
   U33 : INV_X2 port map( I => n102, ZN => n929);
   U8994 : NOR2_X1 port map( A1 => n5316, A2 => n5315, ZN => n7236);
   U1418 : OAI22_X2 port map( A1 => n9564, A2 => n9179, B1 => n9567, B2 => n953
                           , ZN => n9565);
   U467 : INV_X1 port map( I => n18540, ZN => n469);
   U20050 : NOR2_X2 port map( A1 => n9967, A2 => n15809, ZN => n15810);
   U8120 : OAI21_X2 port map( A1 => n11660, A2 => n460, B => n8315, ZN => n8763
                           );
   U326 : INV_X4 port map( I => n19499, ZN => n811);
   U10004 : NAND2_X2 port map( A1 => n2835, A2 => n14357, ZN => n3847);
   U8033 : AOI22_X2 port map( A1 => n10584, A2 => n1256, B1 => n12318, B2 => 
                           n22570, ZN => n12317);
   U1431 : NOR2_X2 port map( A1 => n18919, A2 => n12196, ZN => n18840);
   U20336 : INV_X2 port map( I => n15540, ZN => n18687);
   U3554 : NOR2_X2 port map( A1 => n7261, A2 => n9089, ZN => n9180);
   U19536 : NAND2_X1 port map( A1 => n13034, A2 => n929, ZN => n13033);
   U874 : NOR2_X2 port map( A1 => n27381, A2 => n9314, ZN => n16491);
   U5217 : AOI21_X2 port map( A1 => n17893, A2 => n8126, B => n17892, ZN => 
                           n18939);
   U5788 : NAND2_X2 port map( A1 => n16140, A2 => n11423, ZN => n2343);
   U5540 : INV_X1 port map( I => n8627, ZN => n10121);
   U6836 : INV_X2 port map( I => n21773, ZN => n8303);
   U9766 : NAND2_X2 port map( A1 => n8994, A2 => n1021, ZN => n1905);
   U6116 : INV_X1 port map( I => n22000, ZN => n12124);
   U3713 : INV_X2 port map( I => n18710, ZN => n14207);
   U16112 : AOI21_X2 port map( A1 => n1101, A2 => n13754, B => n8480, ZN => 
                           n8479);
   U12846 : INV_X2 port map( I => n4801, ZN => n4800);
   U13587 : OAI21_X2 port map( A1 => n17478, A2 => n25608, B => n23275, ZN => 
                           n4801);
   U2156 : NAND2_X1 port map( A1 => n751, A2 => n287, ZN => n4655);
   U5123 : BUF_X2 port map( I => n11603, Z => n8864);
   U4537 : BUF_X2 port map( I => n5721, Z => n2569);
   U7444 : OAI22_X1 port map( A1 => n18935, A2 => n11331, B1 => n14779, B2 => 
                           n19019, ZN => n5711);
   U106 : NAND2_X2 port map( A1 => n21713, A2 => n14334, ZN => n13174);
   U948 : INV_X2 port map( I => n15526, ZN => n15982);
   U5631 : INV_X2 port map( I => n18124, ZN => n18516);
   U17246 : INV_X4 port map( I => n9252, ZN => n11761);
   U3693 : INV_X2 port map( I => n16646, ZN => n16681);
   U6790 : NAND2_X2 port map( A1 => n1263, A2 => n8873, ZN => n8872);
   U6756 : OAI21_X2 port map( A1 => n6240, A2 => n6713, B => n9526, ZN => n6239
                           );
   U1581 : AOI21_X2 port map( A1 => n3867, A2 => n23920, B => n3386, ZN => 
                           n3866);
   U6325 : OAI21_X2 port map( A1 => n5116, A2 => n5115, B => n23966, ZN => 
                           n5113);
   U4321 : INV_X4 port map( I => n12884, ZN => n14177);
   U2096 : NOR2_X2 port map( A1 => n6701, A2 => n21361, ZN => n6700);
   U3993 : AND3_X1 port map( A1 => n16577, A2 => n16576, A3 => n1253, Z => 
                           n16579);
   U6420 : INV_X2 port map( I => n9076, ZN => n14345);
   U1889 : NAND2_X1 port map( A1 => n76, A2 => n75, ZN => n74);
   U5542 : INV_X2 port map( I => n11551, ZN => n1134);
   U19321 : OAI21_X1 port map( A1 => n23011, A2 => n17927, B => n12429, ZN => 
                           n17744);
   U3217 : OR2_X1 port map( A1 => n8666, A2 => n12025, Z => n4969);
   U5133 : NAND2_X2 port map( A1 => n24421, A2 => n734, ZN => n20571);
   U9812 : NOR2_X1 port map( A1 => n14931, A2 => n9751, ZN => n14932);
   U99 : BUF_X4 port map( I => n20815, Z => n7518);
   U450 : INV_X2 port map( I => n8467, ZN => n13946);
   U11021 : INV_X2 port map( I => n15228, ZN => n19586);
   U3710 : NOR3_X2 port map( A1 => n2238, A2 => n2285, A3 => n25903, ZN => 
                           n1464);
   U7040 : INV_X2 port map( I => n4064, ZN => n10444);
   U9984 : NAND2_X1 port map( A1 => n6369, A2 => n1037, ZN => n6362);
   U5157 : OAI21_X2 port map( A1 => n24478, A2 => n19747, B => n1125, ZN => 
                           n2035);
   U8770 : NAND3_X1 port map( A1 => n13259, A2 => n5575, A3 => n5577, ZN => 
                           n11231);
   U6961 : NAND2_X2 port map( A1 => n9676, A2 => n6676, ZN => n21057);
   U682 : OAI21_X1 port map( A1 => n27670, A2 => n10141, B => n17241, ZN => 
                           n7695);
   U9990 : AOI21_X2 port map( A1 => n10634, A2 => n17381, B => n7433, ZN => 
                           n11773);
   U2794 : INV_X4 port map( I => n15930, ZN => n7525);
   U531 : NAND2_X1 port map( A1 => n7100, A2 => n7099, ZN => n247);
   U13998 : NOR2_X2 port map( A1 => n4281, A2 => n28231, ZN => n15496);
   U4237 : NOR3_X1 port map( A1 => n13213, A2 => n7167, A3 => n964, ZN => 
                           n13688);
   U8593 : OAI21_X1 port map( A1 => n1080, A2 => n21702, B => n15208, ZN => 
                           n12402);
   U14868 : NAND3_X1 port map( A1 => n20636, A2 => n20634, A3 => n20635, ZN => 
                           n6734);
   U7649 : NAND2_X1 port map( A1 => n17782, A2 => n9105, ZN => n6622);
   U16801 : OAI21_X2 port map( A1 => n23676, A2 => n28408, B => n744, ZN => 
                           n13485);
   U281 : INV_X2 port map( I => n4246, ZN => n19831);
   U7298 : INV_X1 port map( I => n10704, ZN => n19774);
   U274 : INV_X1 port map( I => n3600, ZN => n1129);
   U8157 : AOI22_X2 port map( A1 => n16150, A2 => n8398, B1 => n8925, B2 => 
                           n8926, ZN => n5007);
   U12370 : NAND2_X2 port map( A1 => n3981, A2 => n2976, ZN => n4168);
   U4968 : INV_X1 port map( I => n27737, ZN => n760);
   U6110 : OR2_X1 port map( A1 => n14472, A2 => n9190, Z => n9189);
   U822 : NAND2_X1 port map( A1 => n10891, A2 => n8021, ZN => n125);
   U12584 : NAND2_X1 port map( A1 => n11927, A2 => n12106, ZN => n3158);
   U5065 : NOR2_X2 port map( A1 => n15712, A2 => n16345, ZN => n11962);
   U5843 : BUF_X2 port map( I => Key(28), Z => n14593);
   U5841 : BUF_X2 port map( I => Key(112), Z => n14492);
   U8323 : BUF_X2 port map( I => Key(184), Z => n21141);
   U5845 : BUF_X2 port map( I => Key(73), Z => n20650);
   U4345 : CLKBUF_X2 port map( I => Key(66), Z => n14445);
   U6870 : BUF_X2 port map( I => Key(100), Z => n14614);
   U10656 : BUF_X2 port map( I => Key(16), Z => n14652);
   U5834 : BUF_X2 port map( I => Key(13), Z => n20433);
   U8398 : BUF_X2 port map( I => Key(102), Z => n21649);
   U5088 : CLKBUF_X2 port map( I => Key(88), Z => n14543);
   U6871 : BUF_X2 port map( I => Key(30), Z => n20851);
   U4342 : CLKBUF_X2 port map( I => Key(51), Z => n21523);
   U6859 : BUF_X2 port map( I => Key(133), Z => n20871);
   U4346 : CLKBUF_X2 port map( I => Key(106), Z => n20607);
   U10681 : CLKBUF_X2 port map( I => Key(29), Z => n21085);
   U8369 : BUF_X2 port map( I => Key(42), Z => n14620);
   U4850 : CLKBUF_X2 port map( I => Key(1), Z => n14537);
   U10714 : CLKBUF_X2 port map( I => Key(179), Z => n20396);
   U4510 : CLKBUF_X2 port map( I => Key(54), Z => n14405);
   U5403 : BUF_X2 port map( I => n15923, Z => n15878);
   U19523 : INV_X1 port map( I => n573, ZN => n13430);
   U10597 : BUF_X2 port map( I => n15834, Z => n14171);
   U10611 : BUF_X2 port map( I => n15848, Z => n15919);
   U8310 : INV_X1 port map( I => n4990, ZN => n8173);
   U5402 : BUF_X2 port map( I => n9437, Z => n4926);
   U943 : INV_X2 port map( I => n15981, ZN => n15979);
   U10555 : BUF_X2 port map( I => n15958, Z => n14546);
   U2633 : NAND2_X1 port map( A1 => n15980, A2 => n16136, ZN => n15927);
   U17123 : OR2_X1 port map( A1 => n14832, A2 => n3298, Z => n9000);
   U10503 : INV_X1 port map( I => n4380, ZN => n4231);
   U20561 : NAND2_X1 port map( A1 => n16100, A2 => n16241, ZN => n16102);
   U10396 : NAND2_X1 port map( A1 => n9085, A2 => n9084, ZN => n7333);
   U10374 : INV_X1 port map( I => n3199, ZN => n4490);
   U2346 : CLKBUF_X2 port map( I => n16618, Z => n173);
   U4829 : INV_X2 port map( I => n13721, ZN => n16513);
   U8016 : AOI21_X1 port map( A1 => n14891, A2 => n1257, B => n14820, ZN => 
                           n15336);
   U10292 : INV_X1 port map( I => n16360, ZN => n2709);
   U1946 : NOR2_X1 port map( A1 => n16551, A2 => n92, ZN => n5773);
   U7980 : NAND2_X1 port map( A1 => n16554, A2 => n4737, ZN => n16367);
   U10200 : INV_X1 port map( I => n11598, ZN => n10193);
   U10137 : INV_X1 port map( I => n16744, ZN => n17097);
   U10144 : INV_X1 port map( I => n4776, ZN => n5625);
   U6628 : CLKBUF_X4 port map( I => n17334, Z => n10539);
   U6640 : CLKBUF_X4 port map( I => n17250, Z => n14509);
   U16390 : INV_X2 port map( I => n7482, ZN => n10081);
   U10113 : BUF_X2 port map( I => n17221, Z => n14062);
   U11968 : NAND2_X1 port map( A1 => n2863, A2 => n2527, ZN => n2862);
   U18838 : OR2_X1 port map( A1 => n12639, A2 => n14592, Z => n14771);
   U20769 : NAND2_X1 port map( A1 => n17338, A2 => n347, ZN => n17339);
   U6533 : INV_X1 port map( I => n10821, ZN => n3342);
   U4060 : INV_X2 port map( I => n17724, ZN => n14230);
   U631 : INV_X2 port map( I => n14269, ZN => n17915);
   U12728 : OAI21_X1 port map( A1 => n11514, A2 => n22734, B => n3235, ZN => 
                           n11939);
   U1034 : INV_X1 port map( I => n18095, ZN => n1480);
   U3111 : CLKBUF_X1 port map( I => n643, Z => n376);
   U2685 : CLKBUF_X2 port map( I => n18649, Z => n277);
   U1913 : INV_X1 port map( I => n18753, ZN => n1009);
   U13034 : NOR2_X1 port map( A1 => n11070, A2 => n277, ZN => n3388);
   U17223 : NAND2_X1 port map( A1 => n9248, A2 => n9198, ZN => n9249);
   U505 : NOR2_X1 port map( A1 => n23666, A2 => n15227, ZN => n18028);
   U7498 : NAND2_X1 port map( A1 => n4198, A2 => n18454, ZN => n1502);
   U967 : INV_X2 port map( I => n18719, ZN => n18491);
   U12231 : OR2_X1 port map( A1 => n9348, A2 => n2783, Z => n2782);
   U9546 : INV_X1 port map( I => n18648, ZN => n11703);
   U5586 : BUF_X2 port map( I => n18794, Z => n7084);
   U428 : INV_X2 port map( I => n14098, ZN => n19190);
   U18359 : NAND2_X1 port map( A1 => n24743, A2 => n26762, ZN => n11118);
   U4748 : BUF_X2 port map( I => n28384, Z => n14257);
   U7438 : NAND2_X1 port map( A1 => n1163, A2 => n22981, ZN => n12428);
   U9377 : INV_X1 port map( I => n8301, ZN => n6602);
   U21027 : NAND2_X1 port map( A1 => n19028, A2 => n24055, ZN => n19029);
   U12418 : NAND2_X1 port map( A1 => n18787, A2 => n3009, ZN => n3015);
   U1832 : CLKBUF_X2 port map( I => n8704, Z => n63);
   U9190 : INV_X1 port map( I => n11054, ZN => n4048);
   U330 : CLKBUF_X4 port map( I => n19949, Z => n14651);
   U4055 : INV_X2 port map( I => n2076, ZN => n15478);
   U7312 : CLKBUF_X2 port map( I => n19399, Z => n7238);
   U7317 : BUF_X2 port map( I => n14039, Z => n2925);
   U1107 : NAND2_X1 port map( A1 => n10041, A2 => n14109, ZN => n9418);
   U21152 : NAND2_X1 port map( A1 => n6861, A2 => n19730, ZN => n19677);
   U9051 : NAND2_X1 port map( A1 => n19543, A2 => n6263, ZN => n6262);
   U5171 : INV_X2 port map( I => n6219, ZN => n19823);
   U270 : INV_X1 port map( I => n19913, ZN => n8227);
   U7217 : NAND2_X1 port map( A1 => n775, A2 => n777, ZN => n8325);
   U324 : INV_X2 port map( I => n19802, ZN => n969);
   U3734 : NAND2_X1 port map( A1 => n19763, A2 => n10041, ZN => n11094);
   U8974 : NAND2_X1 port map( A1 => n19695, A2 => n9361, ZN => n6893);
   U1124 : INV_X2 port map( I => n9899, ZN => n20188);
   U8836 : INV_X1 port map( I => n4269, ZN => n5856);
   U160 : NAND2_X1 port map( A1 => n4655, A2 => n4654, ZN => n4653);
   U7106 : NAND3_X1 port map( A1 => n26140, A2 => n20073, A3 => n4225, ZN => 
                           n20058);
   U8804 : NAND2_X1 port map( A1 => n6313, A2 => n957, ZN => n4370);
   U7077 : NAND2_X1 port map( A1 => n20149, A2 => n11870, ZN => n2974);
   U8834 : INV_X1 port map( I => n20097, ZN => n6820);
   U17552 : INV_X1 port map( I => n23825, ZN => n20383);
   U19977 : INV_X2 port map( I => n14183, ZN => n20865);
   U5997 : BUF_X2 port map( I => n21266, Z => n21500);
   U6994 : NOR2_X1 port map( A1 => n20853, A2 => n20979, ZN => n15603);
   U8640 : NAND3_X1 port map( A1 => n15616, A2 => n21666, A3 => n4623, ZN => 
                           n15482);
   U18905 : NAND3_X1 port map( A1 => n12353, A2 => n12352, A3 => n23999, ZN => 
                           n11515);
   U8592 : INV_X1 port map( I => n5261, ZN => n13446);
   U7002 : INV_X1 port map( I => n1739, ZN => n1738);
   U12703 : NAND2_X1 port map( A1 => n14612, A2 => n14613, ZN => n3221);
   U6938 : NAND2_X1 port map( A1 => n15742, A2 => n20911, ZN => n4345);
   U19053 : NAND2_X1 port map( A1 => n22844, A2 => n6517, ZN => n11741);
   U21557 : AOI21_X1 port map( A1 => n21612, A2 => n15475, B => n12517, ZN => 
                           n21595);
   U8395 : BUF_X2 port map( I => Key(130), Z => n14526);
   U6865 : BUF_X2 port map( I => Key(115), Z => n21384);
   U4661 : CLKBUF_X2 port map( I => Key(127), Z => n14574);
   U8370 : CLKBUF_X2 port map( I => Key(134), Z => n20617);
   U16779 : INV_X2 port map( I => n8264, ZN => n16167);
   U10627 : CLKBUF_X2 port map( I => n16143, Z => n14530);
   U6783 : NOR2_X1 port map( A1 => n16293, A2 => n16182, ZN => n5790);
   U8182 : AOI21_X1 port map( A1 => n15977, A2 => n13677, B => n15976, ZN => 
                           n13813);
   U10441 : OAI21_X1 port map( A1 => n4405, A2 => n16305, B => n3771, ZN => 
                           n16311);
   U8181 : AOI21_X1 port map( A1 => n9364, A2 => n4456, B => n25017, ZN => 
                           n3199);
   U1441 : NAND2_X1 port map( A1 => n16813, A2 => n16810, ZN => n16553);
   U10109 : BUF_X2 port map( I => n13320, Z => n6977);
   U10100 : INV_X1 port map( I => n10563, ZN => n8252);
   U6621 : INV_X2 port map( I => n4127, ZN => n8125);
   U758 : CLKBUF_X4 port map( I => n17180, Z => n17335);
   U10070 : OAI22_X1 port map( A1 => n540, A2 => n613, B1 => n28353, B2 => 
                           n23777, ZN => n2863);
   U10053 : NAND2_X1 port map( A1 => n17407, A2 => n17312, ZN => n8253);
   U15928 : NAND2_X1 port map( A1 => n10821, A2 => n14998, ZN => n13767);
   U6445 : NAND2_X1 port map( A1 => n5955, A2 => n18101, ZN => n7825);
   U15349 : AOI21_X1 port map( A1 => n11264, A2 => n22781, B => n8323, ZN => 
                           n9735);
   U9736 : INV_X1 port map( I => n11661, ZN => n4015);
   U4990 : NAND2_X1 port map( A1 => n10817, A2 => n9675, ZN => n10137);
   U7702 : OAI21_X1 port map( A1 => n7615, A2 => n23056, B => n7614, ZN => 
                           n7613);
   U514 : INV_X1 port map( I => n6029, ZN => n18780);
   U529 : BUF_X2 port map( I => n7383, Z => n4639);
   U20947 : NAND2_X1 port map( A1 => n18470, A2 => n18696, ZN => n18407);
   U3630 : NOR2_X1 port map( A1 => n18028, A2 => n18786, ZN => n18031);
   U434 : CLKBUF_X4 port map( I => n6598, Z => n1152);
   U5175 : CLKBUF_X1 port map( I => n19397, Z => n14109);
   U18140 : NOR2_X1 port map( A1 => n19730, A2 => n7326, ZN => n11334);
   U4731 : NAND2_X1 port map( A1 => n15383, A2 => n7376, ZN => n19519);
   U7263 : NAND2_X1 port map( A1 => n3006, A2 => n27401, ZN => n19646);
   U17948 : OAI21_X1 port map( A1 => n19743, A2 => n9812, B => n14507, ZN => 
                           n19745);
   U21310 : OR2_X1 port map( A1 => n20462, A2 => n14666, Z => n20463);
   U15610 : NAND2_X1 port map( A1 => n9868, A2 => n6473, ZN => n9867);
   U10692 : CLKBUF_X2 port map( I => Key(49), Z => n14575);
   U10676 : CLKBUF_X2 port map( I => Key(43), Z => n21104);
   U8386 : CLKBUF_X2 port map( I => Key(180), Z => n20807);
   U6803 : NOR3_X1 port map( A1 => n719, A2 => n16330, A3 => n720, ZN => n4488)
                           ;
   U5774 : AOI21_X1 port map( A1 => n5615, A2 => n15938, B => n16302, ZN => 
                           n5614);
   U20659 : INV_X1 port map( I => n16897, ZN => n16798);
   U1611 : CLKBUF_X2 port map( I => n9027, Z => n3);
   U3832 : CLKBUF_X1 port map( I => n17193, Z => n7055);
   U19501 : NAND2_X1 port map( A1 => n17556, A2 => n24299, ZN => n12871);
   U12257 : OAI21_X1 port map( A1 => n831, A2 => n22620, B => n2901, ZN => 
                           n2815);
   U20708 : OAI21_X1 port map( A1 => n17400, A2 => n17401, B => n8692, ZN => 
                           n16995);
   U18090 : NOR2_X1 port map( A1 => n17467, A2 => n25796, ZN => n17404);
   U7775 : INV_X1 port map( I => n22781, ZN => n17623);
   U3849 : CLKBUF_X2 port map( I => n13205, Z => n6690);
   U17734 : NOR2_X1 port map( A1 => n10816, A2 => n10513, ZN => n10817);
   U17556 : INV_X2 port map( I => n10061, ZN => n14342);
   U9756 : CLKBUF_X2 port map( I => n17731, Z => n5890);
   U4768 : INV_X1 port map( I => n10206, ZN => n5338);
   U20399 : BUF_X2 port map( I => n17983, Z => n18674);
   U4595 : NAND2_X1 port map( A1 => n18752, A2 => n14287, ZN => n6755);
   U456 : INV_X2 port map( I => n23060, ZN => n2070);
   U9385 : NAND2_X1 port map( A1 => n22809, A2 => n19101, ZN => n18906);
   U6307 : INV_X2 port map( I => n11906, ZN => n874);
   U7403 : NAND2_X1 port map( A1 => n10083, A2 => n2726, ZN => n9408);
   U7342 : NOR2_X1 port map( A1 => n19061, A2 => n19062, ZN => n13595);
   U3927 : INV_X1 port map( I => n9612, ZN => n9812);
   U8571 : NAND2_X1 port map( A1 => n5045, A2 => n5044, ZN => n2622);
   U19088 : AOI21_X1 port map( A1 => n4428, A2 => n21116, B => n25342, ZN => 
                           n13471);
   U18204 : OAI21_X1 port map( A1 => n14146, A2 => n20625, B => n24597, ZN => 
                           n13080);
   U7609 : BUF_X4 port map( I => n18442, Z => n12375);
   U10252 : NAND3_X2 port map( A1 => n7864, A2 => n7862, A3 => n16681, ZN => 
                           n16002);
   U10019 : OAI21_X2 port map( A1 => n5409, A2 => n894, B => n5408, ZN => 
                           n17236);
   U3143 : NAND2_X2 port map( A1 => n19007, A2 => n19006, ZN => n13045);
   U13999 : INV_X4 port map( I => n17479, ZN => n10141);
   U10106 : BUF_X2 port map( I => n17198, Z => n17433);
   U8299 : BUF_X2 port map( I => n16068, Z => n16240);
   U8285 : INV_X2 port map( I => n10269, ZN => n16332);
   U10551 : INV_X2 port map( I => n16339, ZN => n8191);
   U5390 : INV_X2 port map( I => n15330, ZN => n16300);
   U20537 : NOR2_X1 port map( A1 => n12272, A2 => n16013, ZN => n15990);
   U17844 : OAI21_X1 port map( A1 => n16314, A2 => n16240, B => n9768, ZN => 
                           n15106);
   U20533 : NOR2_X1 port map( A1 => n16119, A2 => n14546, ZN => n15976);
   U17858 : NOR2_X1 port map( A1 => n25224, A2 => n13435, ZN => n14252);
   U15834 : NAND2_X1 port map( A1 => n16082, A2 => n16253, ZN => n16257);
   U8159 : NOR3_X1 port map( A1 => n15885, A2 => n24271, A3 => n16300, ZN => 
                           n6304);
   U20005 : NOR2_X1 port map( A1 => n14857, A2 => n14858, ZN => n15931);
   U4501 : NOR2_X1 port map( A1 => n14557, A2 => n16064, ZN => n16313);
   U2688 : AOI21_X1 port map( A1 => n16082, A2 => n16220, B => n15559, ZN => 
                           n6064);
   U6800 : NAND2_X1 port map( A1 => n12918, A2 => n798, ZN => n14384);
   U10490 : NAND2_X1 port map( A1 => n3794, A2 => n4532, ZN => n3793);
   U18016 : NAND2_X1 port map( A1 => n22454, A2 => n1267, ZN => n16445);
   U10489 : AOI21_X1 port map( A1 => n799, A2 => n4115, B => n4114, ZN => n4113
                           );
   U6760 : AOI21_X1 port map( A1 => n15878, A2 => n9787, B => n15770, ZN => 
                           n9786);
   U8156 : NOR2_X1 port map( A1 => n15262, A2 => n15261, ZN => n15260);
   U4318 : INV_X2 port map( I => n16468, ZN => n4295);
   U2513 : BUF_X4 port map( I => n15239, Z => n15061);
   U3666 : INV_X1 port map( I => n16419, ZN => n3913);
   U18986 : NAND2_X1 port map( A1 => n8344, A2 => n479, ZN => n14069);
   U8051 : NAND2_X1 port map( A1 => n16483, A2 => n7395, ZN => n7416);
   U20609 : NAND2_X1 port map( A1 => n16450, A2 => n16654, ZN => n16453);
   U12863 : NOR2_X1 port map( A1 => n1051, A2 => n173, ZN => n16547);
   U1877 : AOI21_X1 port map( A1 => n13211, A2 => n16672, B => n571, ZN => 
                           n10397);
   U7999 : NAND2_X1 port map( A1 => n6939, A2 => n6937, ZN => n6936);
   U824 : INV_X1 port map( I => n25875, ZN => n908);
   U5041 : NAND3_X1 port map( A1 => n24580, A2 => n16563, A3 => n12026, ZN => 
                           n3063);
   U20599 : NAND3_X1 port map( A1 => n16383, A2 => n16687, A3 => n16382, ZN => 
                           n16384);
   U14666 : OAI21_X1 port map( A1 => n5324, A2 => n5266, B => n5265, ZN => 
                           n16179);
   U1856 : NOR2_X1 port map( A1 => n2760, A2 => n1793, ZN => n2761);
   U10236 : AOI21_X1 port map( A1 => n16547, A2 => n14337, B => n16546, ZN => 
                           n12213);
   U2957 : INV_X1 port map( I => n16868, ZN => n10279);
   U803 : INV_X1 port map( I => n26576, ZN => n15162);
   U5717 : BUF_X2 port map( I => n17217, Z => n10942);
   U746 : INV_X2 port map( I => n17324, ZN => n7912);
   U7824 : NOR3_X1 port map( A1 => n17510, A2 => n4832, A3 => n5489, ZN => 
                           n9410);
   U6546 : OAI21_X1 port map( A1 => n1892, A2 => n24774, B => n14658, ZN => 
                           n16548);
   U12540 : INV_X1 port map( I => n613, ZN => n8273);
   U11269 : INV_X2 port map( I => n636, ZN => n17431);
   U737 : NAND2_X1 port map( A1 => n8996, A2 => n14509, ZN => n17485);
   U2315 : NOR2_X1 port map( A1 => n2901, A2 => n1232, ZN => n1966);
   U6609 : NOR3_X1 port map( A1 => n11761, A2 => n14103, A3 => n12692, ZN => 
                           n15735);
   U695 : NOR2_X1 port map( A1 => n13693, A2 => n11857, ZN => n15394);
   U10066 : OR2_X1 port map( A1 => n12549, A2 => n17475, Z => n17538);
   U704 : NOR2_X1 port map( A1 => n9358, A2 => n22918, ZN => n9987);
   U10038 : INV_X1 port map( I => n2934, ZN => n12553);
   U12270 : NAND3_X1 port map( A1 => n2831, A2 => n8273, A3 => n23778, ZN => 
                           n7715);
   U20788 : NAND3_X1 port map( A1 => n17444, A2 => n17443, A3 => n27168, ZN => 
                           n17445);
   U10016 : NAND2_X1 port map( A1 => n4172, A2 => n3624, ZN => n3623);
   U7876 : INV_X1 port map( I => n23276, ZN => n4798);
   U5290 : NOR2_X1 port map( A1 => n25013, A2 => n9879, ZN => n6330);
   U7771 : INV_X1 port map( I => n24127, ZN => n17904);
   U6461 : NOR2_X1 port map( A1 => n17676, A2 => n9330, ZN => n9329);
   U6484 : CLKBUF_X2 port map( I => n13530, Z => n5238);
   U2100 : NAND2_X1 port map( A1 => n1217, A2 => n10513, ZN => n17612);
   U5644 : INV_X1 port map( I => n17702, ZN => n2562);
   U14286 : NAND2_X1 port map( A1 => n4828, A2 => n9105, ZN => n17860);
   U15699 : NAND3_X1 port map( A1 => n17523, A2 => n18130, A3 => n6620, ZN => 
                           n9356);
   U18317 : INV_X1 port map( I => n25312, ZN => n14322);
   U20280 : INV_X1 port map( I => n18482, ZN => n18663);
   U2269 : INV_X1 port map( I => n12023, ZN => n14332);
   U12039 : NOR3_X1 port map( A1 => n18769, A2 => n18770, A3 => n8576, ZN => 
                           n2602);
   U17926 : NAND2_X1 port map( A1 => n288, A2 => n14128, ZN => n14828);
   U18094 : NAND2_X1 port map( A1 => n14022, A2 => n5115, ZN => n10873);
   U4767 : INV_X1 port map( I => n5338, ZN => n1167);
   U6311 : NOR2_X1 port map( A1 => n8623, A2 => n6438, ZN => n2735);
   U17812 : NOR2_X1 port map( A1 => n27457, A2 => n18505, ZN => n11704);
   U6326 : AOI21_X1 port map( A1 => n18628, A2 => n18546, B => n3416, ZN => 
                           n8270);
   U7542 : INV_X1 port map( I => n6827, ZN => n7687);
   U4589 : OAI21_X1 port map( A1 => n15143, A2 => n5320, B => n15142, ZN => 
                           n19147);
   U9478 : OR2_X1 port map( A1 => n18464, A2 => n8113, Z => n14721);
   U1556 : INV_X1 port map( I => n18947, ZN => n757);
   U6294 : INV_X1 port map( I => n4953, ZN => n18912);
   U4428 : NAND2_X1 port map( A1 => n10205, A2 => n18828, ZN => n3315);
   U6257 : NAND2_X1 port map( A1 => n9376, A2 => n11696, ZN => n6599);
   U9349 : NAND2_X1 port map( A1 => n22882, A2 => n19157, ZN => n9881);
   U7399 : NOR2_X1 port map( A1 => n22019, A2 => n14358, ZN => n13869);
   U12140 : INV_X2 port map( I => n19623, ZN => n19790);
   U5534 : NAND2_X1 port map( A1 => n19743, A2 => n19744, ZN => n14507);
   U4248 : INV_X2 port map( I => n11175, ZN => n13771);
   U5161 : INV_X1 port map( I => n19614, ZN => n19888);
   U5533 : INV_X1 port map( I => n5253, ZN => n15295);
   U21161 : NOR2_X1 port map( A1 => n26654, A2 => n19586, ZN => n19706);
   U19051 : NAND2_X1 port map( A1 => n11213, A2 => n9762, ZN => n15046);
   U308 : CLKBUF_X2 port map( I => n19870, Z => n463);
   U21150 : NAND2_X1 port map( A1 => n23864, A2 => n26767, ZN => n19668);
   U12096 : NOR2_X1 port map( A1 => n14282, A2 => n19918, ZN => n11317);
   U7220 : NAND2_X1 port map( A1 => n5308, A2 => n8952, ZN => n7037);
   U4730 : OAI21_X1 port map( A1 => n19624, A2 => n19623, B => n2320, ZN => 
                           n6954);
   U9009 : NOR2_X1 port map( A1 => n7037, A2 => n7036, ZN => n9193);
   U11948 : NOR2_X1 port map( A1 => n2656, A2 => n5616, ZN => n10721);
   U8854 : NAND2_X1 port map( A1 => n20029, A2 => n14059, ZN => n11255);
   U6093 : INV_X1 port map( I => n20156, ZN => n1109);
   U5477 : INV_X1 port map( I => n20138, ZN => n6471);
   U12145 : INV_X1 port map( I => n23817, ZN => n20197);
   U18377 : NAND2_X1 port map( A1 => n20491, A2 => n12712, ZN => n20492);
   U15694 : NAND2_X1 port map( A1 => n20165, A2 => n24862, ZN => n20128);
   U16000 : AOI21_X1 port map( A1 => n20126, A2 => n20309, B => n14063, ZN => 
                           n14157);
   U8715 : INV_X1 port map( I => n8879, ZN => n2770);
   U94 : INV_X1 port map( I => n21931, ZN => n13772);
   U18225 : AOI21_X1 port map( A1 => n22800, A2 => n13432, B => n8668, ZN => 
                           n13431);
   U6995 : NAND2_X1 port map( A1 => n20977, A2 => n3125, ZN => n10351);
   U14352 : NOR2_X1 port map( A1 => n22828, A2 => n850, ZN => n20590);
   U5442 : NAND2_X1 port map( A1 => n22828, A2 => n24576, ZN => n4086);
   U14700 : NOR2_X1 port map( A1 => n21328, A2 => n15463, ZN => n10253);
   U21389 : INV_X1 port map( I => n27332, ZN => n20855);
   U5899 : INV_X1 port map( I => n20879, ZN => n20876);
   U8505 : NAND2_X1 port map( A1 => n940, A2 => n12517, ZN => n13830);
   U19 : NAND2_X1 port map( A1 => n3972, A2 => n7811, ZN => n22753);
   U43 : NOR2_X1 port map( A1 => n21175, A2 => n20263, ZN => n22208);
   U54 : NAND2_X1 port map( A1 => n15315, A2 => n20644, ZN => n23323);
   U60 : OAI21_X1 port map( A1 => n14647, A2 => n20786, B => n20781, ZN => 
                           n9333);
   U79 : NAND2_X1 port map( A1 => n11248, A2 => n15378, ZN => n23226);
   U81 : NAND2_X1 port map( A1 => n21273, A2 => n3530, ZN => n20063);
   U85 : NOR2_X1 port map( A1 => n27406, A2 => n850, ZN => n21727);
   U90 : NOR2_X1 port map( A1 => n14647, A2 => n20739, ZN => n23870);
   U125 : BUF_X2 port map( I => n20735, Z => n15689);
   U134 : NAND2_X1 port map( A1 => n21723, A2 => n21699, ZN => n22652);
   U174 : NAND3_X1 port map( A1 => n23700, A2 => n5934, A3 => n20186, ZN => 
                           n11556);
   U191 : INV_X1 port map( I => n5616, ZN => n22581);
   U294 : NAND2_X1 port map( A1 => n28199, A2 => n8756, ZN => n22213);
   U431 : INV_X1 port map( I => n11417, ZN => n22866);
   U449 : NOR2_X1 port map( A1 => n3312, A2 => n15041, ZN => n24332);
   U464 : NAND3_X1 port map( A1 => n24062, A2 => n6145, A3 => n28136, ZN => 
                           n3010);
   U507 : OR2_X1 port map( A1 => n19159, A2 => n22345, Z => n21918);
   U552 : NOR2_X1 port map( A1 => n28491, A2 => n4199, ZN => n24472);
   U566 : INV_X2 port map( I => n19148, ZN => n19009);
   U588 : NOR2_X1 port map( A1 => n736, A2 => n18426, ZN => n1577);
   U592 : NAND2_X1 port map( A1 => n19163, A2 => n19161, ZN => n24382);
   U619 : INV_X2 port map( I => n18396, ZN => n180);
   U692 : NAND2_X1 port map( A1 => n737, A2 => n9730, ZN => n22035);
   U703 : NAND2_X1 port map( A1 => n24243, A2 => n2072, ZN => n22339);
   U706 : NOR2_X1 port map( A1 => n15623, A2 => n27631, ZN => n18387);
   U722 : NAND2_X1 port map( A1 => n11382, A2 => n9248, ZN => n12048);
   U723 : NOR2_X1 port map( A1 => n26292, A2 => n15423, ZN => n18484);
   U726 : NAND2_X1 port map( A1 => n14510, A2 => n1018, ZN => n7577);
   U773 : INV_X1 port map( I => n18219, ZN => n24295);
   U807 : NAND3_X1 port map( A1 => n18101, A2 => n22739, A3 => n891, ZN => 
                           n8222);
   U837 : NAND2_X1 port map( A1 => n17606, A2 => n11579, ZN => n23030);
   U839 : NAND2_X1 port map( A1 => n4507, A2 => n12951, ZN => n22599);
   U845 : NAND2_X1 port map( A1 => n6794, A2 => n11112, ZN => n10587);
   U850 : NOR3_X1 port map( A1 => n4590, A2 => n890, A3 => n17349, ZN => n9751)
                           ;
   U883 : NOR2_X1 port map( A1 => n2952, A2 => n4914, ZN => n17615);
   U893 : INV_X1 port map( I => n8075, ZN => n23856);
   U926 : AND2_X1 port map( A1 => n7447, A2 => n7450, Z => n22734);
   U944 : NAND2_X1 port map( A1 => n4414, A2 => n13043, ZN => n8849);
   U998 : NOR2_X1 port map( A1 => n17192, A2 => n1629, ZN => n22498);
   U1008 : OAI22_X1 port map( A1 => n17209, A2 => n26198, B1 => n7003, B2 => 
                           n1222, ZN => n24453);
   U1010 : NAND2_X1 port map( A1 => n17519, A2 => n636, ZN => n23012);
   U1015 : NOR2_X1 port map( A1 => n17313, A2 => n14578, ZN => n6902);
   U1025 : NAND3_X1 port map( A1 => n8263, A2 => n17519, A3 => n23105, ZN => 
                           n9856);
   U1043 : INV_X1 port map( I => n3300, ZN => n10546);
   U1045 : NOR2_X1 port map( A1 => n17313, A2 => n14533, ZN => n17407);
   U1071 : NAND2_X1 port map( A1 => n17336, A2 => n17564, ZN => n16973);
   U1095 : INV_X1 port map( I => n23053, ZN => n23860);
   U1102 : AND2_X1 port map( A1 => n22838, A2 => n24089, Z => n1856);
   U1126 : AND2_X1 port map( A1 => n8373, A2 => n9314, Z => n2658);
   U1130 : INV_X1 port map( I => n16638, ZN => n22929);
   U1140 : OR2_X1 port map( A1 => n10155, A2 => n12331, Z => n1665);
   U1150 : NOR2_X1 port map( A1 => n1046, A2 => n1048, ZN => n23861);
   U1158 : AND2_X1 port map( A1 => n24552, A2 => n1052, Z => n10584);
   U1160 : NAND3_X1 port map( A1 => n14967, A2 => n14969, A3 => n1681, ZN => 
                           n14966);
   U1161 : NOR3_X1 port map( A1 => n10597, A2 => n1256, A3 => n22570, ZN => 
                           n3330);
   U1193 : AND2_X1 port map( A1 => n12331, A2 => n913, Z => n6077);
   U1194 : INV_X1 port map( I => n16455, ZN => n16648);
   U1209 : INV_X2 port map( I => n12331, ZN => n833);
   U1227 : NAND2_X1 port map( A1 => n15973, A2 => n14386, ZN => n5075);
   U1231 : NAND2_X1 port map( A1 => n15973, A2 => n14636, ZN => n15241);
   U1247 : INV_X1 port map( I => n16136, ZN => n15155);
   U1249 : OAI21_X1 port map( A1 => n11568, A2 => n16298, B => n16300, ZN => 
                           n23525);
   U1250 : OR2_X1 port map( A1 => n15930, A2 => n25873, Z => n7158);
   U1252 : OR2_X1 port map( A1 => n14293, A2 => n14644, Z => n21814);
   U1311 : NOR2_X2 port map( A1 => n4940, A2 => n4518, ZN => n11932);
   U1350 : OAI21_X2 port map( A1 => n24491, A2 => n11442, B => n19819, ZN => 
                           n23395);
   U1406 : NOR2_X2 port map( A1 => n6892, A2 => n4898, ZN => n17918);
   U1407 : NAND2_X2 port map( A1 => n11497, A2 => n2549, ZN => n17630);
   U1408 : NAND2_X2 port map( A1 => n18959, A2 => n19143, ZN => n5138);
   U1411 : NOR2_X2 port map( A1 => n934, A2 => n4860, ZN => n20696);
   U1414 : OAI21_X2 port map( A1 => n19875, A2 => n11670, B => n11631, ZN => 
                           n22533);
   U1422 : NAND2_X2 port map( A1 => n14891, A2 => n9759, ZN => n8519);
   U1456 : NAND2_X2 port map( A1 => n28299, A2 => n27647, ZN => n87);
   U1458 : INV_X2 port map( I => n26570, ZN => n5285);
   U1497 : NAND2_X1 port map( A1 => n10477, A2 => n6371, ZN => n22017);
   U1511 : OAI21_X1 port map( A1 => n7913, A2 => n10478, B => n22015, ZN => 
                           n10475);
   U1514 : NAND2_X1 port map( A1 => n21064, A2 => n27426, ZN => n11069);
   U1531 : NAND3_X1 port map( A1 => n21079, A2 => n21078, A3 => n25952, ZN => 
                           n11924);
   U1548 : AOI21_X1 port map( A1 => n13477, A2 => n23748, B => n19843, ZN => 
                           n2004);
   U1551 : AOI21_X1 port map( A1 => n10197, A2 => n21332, B => n4143, ZN => 
                           n5261);
   U1558 : NOR2_X1 port map( A1 => n8452, A2 => n26410, ZN => n6005);
   U1577 : NOR2_X1 port map( A1 => n19082, A2 => n11983, ZN => n18983);
   U1601 : AOI21_X1 port map( A1 => n800, A2 => n20804, B => n935, ZN => n22016
                           );
   U1619 : NOR2_X1 port map( A1 => n2484, A2 => n19045, ZN => n13887);
   U1625 : OAI21_X1 port map( A1 => n17912, A2 => n13061, B => n4508, ZN => 
                           n4507);
   U1633 : NOR2_X1 port map( A1 => n11380, A2 => n7009, ZN => n11379);
   U1637 : CLKBUF_X2 port map( I => n20804, Z => n22536);
   U1654 : NAND2_X1 port map( A1 => n20852, A2 => n20982, ZN => n3125);
   U1659 : INV_X1 port map( I => n11671, ZN => n7187);
   U1669 : NOR2_X1 port map( A1 => n5768, A2 => n7971, ZN => n10763);
   U1678 : NOR2_X1 port map( A1 => n6630, A2 => n25144, ZN => n23510);
   U1700 : NAND2_X1 port map( A1 => n15061, A2 => n24374, ZN => n7862);
   U1712 : AOI21_X1 port map( A1 => n11069, A2 => n9377, B => n944, ZN => n6849
                           );
   U1725 : NAND3_X1 port map( A1 => n4703, A2 => n15041, A3 => n4705, ZN => 
                           n5702);
   U1733 : BUF_X2 port map( I => n21120, Z => n4428);
   U1741 : OAI21_X1 port map( A1 => n2756, A2 => n17520, B => n14917, ZN => 
                           n12194);
   U1761 : NAND2_X1 port map( A1 => n7266, A2 => n15282, ZN => n15940);
   U1767 : AOI21_X1 port map( A1 => n16333, A2 => n769, B => n7266, ZN => 
                           n10270);
   U1780 : AOI21_X1 port map( A1 => n21387, A2 => n21275, B => n21389, ZN => 
                           n14613);
   U1781 : OAI21_X1 port map( A1 => n13447, A2 => n13448, B => n28428, ZN => 
                           n6321);
   U1787 : INV_X1 port map( I => n9619, ZN => n10702);
   U1840 : OAI21_X1 port map( A1 => n19129, A2 => n12111, B => n12139, ZN => 
                           n9060);
   U1859 : NOR2_X1 port map( A1 => n4022, A2 => n22828, ZN => n5045);
   U1879 : NOR2_X1 port map( A1 => n15869, A2 => n14370, ZN => n15994);
   U1934 : NOR2_X1 port map( A1 => n12748, A2 => n17522, ZN => n12554);
   U1958 : AOI21_X1 port map( A1 => n8050, A2 => n8051, B => n21024, ZN => 
                           n22881);
   U1968 : NAND2_X1 port map( A1 => n22033, A2 => n1460, ZN => n1520);
   U2001 : NOR2_X1 port map( A1 => n21083, A2 => n6473, ZN => n21088);
   U2004 : NOR2_X1 port map( A1 => n8968, A2 => n8717, ZN => n8951);
   U2007 : INV_X2 port map( I => n20998, ZN => n928);
   U2044 : NAND2_X1 port map( A1 => n21086, A2 => n21083, ZN => n21078);
   U2053 : AOI21_X1 port map( A1 => n740, A2 => n6681, B => n14453, ZN => n1661
                           );
   U2074 : OAI22_X1 port map( A1 => n14302, A2 => n1459, B1 => n19802, B2 => 
                           n10057, ZN => n22033);
   U2144 : NAND3_X1 port map( A1 => n16338, A2 => n22357, A3 => n15897, ZN => 
                           n15898);
   U2152 : NOR2_X1 port map( A1 => n19, A2 => n23212, ZN => n22417);
   U2167 : NAND3_X1 port map( A1 => n27404, A2 => n21612, A3 => n15469, ZN => 
                           n22427);
   U2169 : INV_X2 port map( I => n7464, ZN => n14279);
   U2177 : NOR2_X1 port map( A1 => n22799, A2 => n18728, ZN => n13369);
   U2194 : NOR2_X1 port map( A1 => n8507, A2 => n12206, ZN => n3217);
   U2195 : INV_X2 port map( I => n14554, ZN => n12206);
   U2196 : NAND2_X1 port map( A1 => n10614, A2 => n24032, ZN => n18563);
   U2203 : INV_X1 port map( I => n14352, ZN => n20744);
   U2214 : NAND2_X1 port map( A1 => n10183, A2 => n12340, ZN => n4577);
   U2221 : INV_X1 port map( I => n576, ZN => n9967);
   U2232 : INV_X1 port map( I => n19140, ZN => n996);
   U2241 : INV_X1 port map( I => n23744, ZN => n1047);
   U2248 : NOR3_X1 port map( A1 => n1519, A2 => n12637, A3 => n16557, ZN => 
                           n4337);
   U2283 : NAND2_X1 port map( A1 => n6373, A2 => n3297, ZN => n16505);
   U2293 : OR2_X1 port map( A1 => n11961, A2 => n11048, Z => n2878);
   U2307 : INV_X1 port map( I => n15728, ZN => n21062);
   U2316 : NAND2_X1 port map( A1 => n3979, A2 => n16426, ZN => n11606);
   U2337 : NOR2_X1 port map( A1 => n19872, A2 => n19873, ZN => n22688);
   U2342 : NAND2_X1 port map( A1 => n11419, A2 => n4898, ZN => n6206);
   U2344 : INV_X1 port map( I => n4898, ZN => n24403);
   U2361 : INV_X1 port map( I => n3729, ZN => n4595);
   U2362 : NAND2_X1 port map( A1 => n16403, A2 => n458, ZN => n16404);
   U2377 : INV_X1 port map( I => n14194, ZN => n5434);
   U2380 : INV_X2 port map( I => n4719, ZN => n17994);
   U2385 : OR3_X1 port map( A1 => n27044, A2 => n27432, A3 => n12978, Z => 
                           n21756);
   U2388 : INV_X2 port map( I => n6047, ZN => n22140);
   U2402 : OAI22_X2 port map( A1 => n3815, A2 => n20207, B1 => n4138, B2 => 
                           n20206, ZN => n4137);
   U2403 : XNOR2_X1 port map( A1 => n21197, A2 => n21357, ZN => n21760);
   U2404 : NAND2_X2 port map( A1 => n1606, A2 => n1607, ZN => n22830);
   U2411 : AND3_X2 port map( A1 => n27414, A2 => n15076, A3 => n20245, Z => 
                           n21761);
   U2438 : NAND2_X1 port map( A1 => n19122, A2 => n19124, ZN => n2091);
   U2471 : OAI22_X1 port map( A1 => n16561, A2 => n8181, B1 => n16449, B2 => 
                           n16448, ZN => n16450);
   U2478 : INV_X1 port map( I => n14320, ZN => n16514);
   U2501 : CLKBUF_X12 port map( I => n13665, Z => n13660);
   U2508 : NAND2_X1 port map( A1 => n14566, A2 => n20244, ZN => n23306);
   U2551 : CLKBUF_X12 port map( I => n21916, Z => n6393);
   U2586 : AOI21_X1 port map( A1 => n7251, A2 => n13771, B => n11110, ZN => 
                           n11111);
   U2587 : NAND3_X1 port map( A1 => n11110, A2 => n15560, A3 => n10293, ZN => 
                           n6666);
   U2684 : NAND2_X1 port map( A1 => n17474, A2 => n26754, ZN => n17531);
   U2702 : INV_X1 port map( I => n11680, ZN => n8547);
   U2704 : INV_X1 port map( I => n14744, ZN => n14743);
   U2725 : INV_X1 port map( I => n9314, ZN => n742);
   U2741 : NAND2_X1 port map( A1 => n5324, A2 => n479, ZN => n16383);
   U2749 : INV_X1 port map( I => n17757, ZN => n786);
   U2760 : OAI21_X1 port map( A1 => n9051, A2 => n27146, B => n23072, ZN => 
                           n22584);
   U2780 : AND2_X1 port map( A1 => n21268, A2 => n5355, Z => n22824);
   U2790 : NAND2_X1 port map( A1 => n21392, A2 => n24538, ZN => n11560);
   U2791 : NOR2_X1 port map( A1 => n24817, A2 => n21387, ZN => n22511);
   U2807 : INV_X1 port map( I => n136, ZN => n23426);
   U2813 : NAND2_X1 port map( A1 => n27484, A2 => n20413, ZN => n23929);
   U2816 : NOR2_X1 port map( A1 => n26154, A2 => n27484, ZN => n5760);
   U2824 : NAND3_X1 port map( A1 => n24408, A2 => n24407, A3 => n23450, ZN => 
                           n22696);
   U2826 : NOR2_X1 port map( A1 => n9446, A2 => n23913, ZN => n23912);
   U2828 : CLKBUF_X1 port map( I => n9899, Z => n22224);
   U2833 : CLKBUF_X2 port map( I => n20065, Z => n22295);
   U2849 : NAND2_X1 port map( A1 => n22748, A2 => n19753, ZN => n22288);
   U2854 : NOR2_X1 port map( A1 => n12431, A2 => n866, ZN => n22056);
   U2861 : AND3_X1 port map( A1 => n12433, A2 => n28527, A3 => n12432, Z => 
                           n21912);
   U2917 : INV_X2 port map( I => n10545, ZN => n21777);
   U2922 : INV_X2 port map( I => n7751, ZN => n884);
   U2943 : NAND2_X1 port map( A1 => n14342, A2 => n17847, ZN => n23020);
   U2961 : NOR3_X1 port map( A1 => n4590, A2 => n23633, A3 => n3621, ZN => 
                           n14708);
   U2994 : NAND2_X1 port map( A1 => n16121, A2 => n9830, ZN => n23261);
   U3009 : NAND2_X1 port map( A1 => n15875, A2 => n13717, ZN => n24270);
   U3014 : OAI21_X1 port map( A1 => n21122, A2 => n4428, B => n21123, ZN => 
                           n22377);
   U3017 : AND2_X1 port map( A1 => n705, A2 => n20964, Z => n23662);
   U3036 : NOR2_X1 port map( A1 => n10666, A2 => n20642, ZN => n23678);
   U3039 : NAND2_X1 port map( A1 => n21666, A2 => n21667, ZN => n15167);
   U3045 : NOR2_X1 port map( A1 => n21266, A2 => n14525, ZN => n23213);
   U3050 : OR2_X1 port map( A1 => n2882, A2 => n10332, Z => n21392);
   U3051 : OR2_X1 port map( A1 => n1381, A2 => n15512, Z => n15129);
   U3066 : NAND2_X1 port map( A1 => n956, A2 => n9087, ZN => n22012);
   U3082 : OAI21_X1 port map( A1 => n23993, A2 => n14059, B => n8610, ZN => 
                           n11356);
   U3089 : OR2_X1 port map( A1 => n12203, A2 => n12124, Z => n12009);
   U3099 : NOR2_X1 port map( A1 => n1835, A2 => n22224, ZN => n8932);
   U3115 : AND2_X1 port map( A1 => n8299, A2 => n11215, Z => n21882);
   U3122 : NOR2_X1 port map( A1 => n19678, A2 => n19587, ZN => n23886);
   U3123 : NAND2_X1 port map( A1 => n19667, A2 => n19790, ZN => n23215);
   U3196 : NOR2_X1 port map( A1 => n3276, A2 => n8611, ZN => n3275);
   U3198 : NOR2_X1 port map( A1 => n24062, A2 => n19010, ZN => n18787);
   U3214 : AND2_X1 port map( A1 => n23302, A2 => n23428, Z => n22809);
   U3238 : NAND2_X1 port map( A1 => n18646, A2 => n24032, ZN => n12870);
   U3243 : AND2_X2 port map( A1 => n4268, A2 => n10097, Z => n8604);
   U3247 : CLKBUF_X2 port map( I => n18773, Z => n13390);
   U3274 : INV_X2 port map( I => n18019, ZN => n21784);
   U3275 : INV_X1 port map( I => n17332, ZN => n23893);
   U3278 : CLKBUF_X2 port map( I => n10107, Z => n23950);
   U3289 : NOR2_X1 port map( A1 => n17712, A2 => n17867, ZN => n22111);
   U3299 : OAI21_X1 port map( A1 => n22851, A2 => n22781, B => n17682, ZN => 
                           n1429);
   U3303 : NAND2_X1 port map( A1 => n18100, A2 => n25192, ZN => n17760);
   U3305 : NOR2_X1 port map( A1 => n17947, A2 => n23441, ZN => n24064);
   U3313 : AOI21_X1 port map( A1 => n21792, A2 => n14180, B => n24397, ZN => 
                           n7601);
   U3319 : OR2_X1 port map( A1 => n17665, A2 => n17694, Z => n17947);
   U3322 : AND2_X1 port map( A1 => n11112, A2 => n17969, Z => n21886);
   U3342 : NAND2_X1 port map( A1 => n3376, A2 => n10568, ZN => n23494);
   U3344 : INV_X1 port map( I => n24649, ZN => n15055);
   U3346 : CLKBUF_X2 port map( I => n1473, Z => n23863);
   U3348 : NAND2_X1 port map( A1 => n23346, A2 => n23345, ZN => n2362);
   U3349 : NAND2_X1 port map( A1 => n2490, A2 => n2576, ZN => n23346);
   U3358 : NAND2_X1 port map( A1 => n16471, A2 => n11932, ZN => n16812);
   U3373 : BUF_X1 port map( I => n10393, Z => n23096);
   U3376 : AND2_X1 port map( A1 => n14766, A2 => n14878, Z => n21800);
   U3379 : OAI22_X1 port map( A1 => n11567, A2 => n16189, B1 => n6359, B2 => 
                           n7022, ZN => n11566);
   U3380 : CLKBUF_X2 port map( I => n13739, Z => n22542);
   U3385 : NOR3_X1 port map( A1 => n516, A2 => n14303, A3 => n16167, ZN => 
                           n12767);
   U3391 : INV_X4 port map( I => n16271, ZN => n21786);
   U3400 : NOR2_X1 port map( A1 => n13080, A2 => n13081, ZN => n23938);
   U3406 : AOI21_X1 port map( A1 => n13436, A2 => n10724, B => n22377, ZN => 
                           n10335);
   U3407 : NAND2_X1 port map( A1 => n7342, A2 => n20592, ZN => n15036);
   U3414 : AOI22_X1 port map( A1 => n705, A2 => n22525, B1 => n4605, B2 => 
                           n4604, ZN => n23980);
   U3426 : INV_X2 port map( I => n13009, ZN => n4277);
   U3429 : NOR2_X1 port map( A1 => n20963, A2 => n22526, ZN => n22525);
   U3435 : CLKBUF_X1 port map( I => n20665, Z => n23119);
   U3436 : AND3_X1 port map( A1 => n3855, A2 => n10040, A3 => n10174, Z => 
                           n22848);
   U3453 : INV_X1 port map( I => n11069, ZN => n23157);
   U3467 : AND2_X1 port map( A1 => n21697, A2 => n15307, Z => n21843);
   U3469 : NOR2_X1 port map( A1 => n15167, A2 => n23999, ZN => n22484);
   U3471 : OR3_X1 port map( A1 => n20928, A2 => n12465, A3 => n20979, Z => 
                           n20929);
   U3472 : AND2_X1 port map( A1 => n12849, A2 => n15335, Z => n23247);
   U3493 : NOR2_X1 port map( A1 => n2569, A2 => n2813, ZN => n22925);
   U3498 : CLKBUF_X4 port map( I => n20777, Z => n20979);
   U3499 : CLKBUF_X2 port map( I => n687, Z => n23991);
   U3520 : BUF_X2 port map( I => n21931, Z => n23802);
   U3522 : CLKBUF_X2 port map( I => n13325, Z => n22364);
   U3525 : BUF_X4 port map( I => n20526, Z => n21024);
   U3540 : CLKBUF_X2 port map( I => n20447, Z => n23156);
   U3552 : CLKBUF_X2 port map( I => n20458, Z => n23173);
   U3555 : NOR2_X1 port map( A1 => n21869, A2 => n22302, ZN => n10967);
   U3566 : AND2_X1 port map( A1 => n11786, A2 => n5198, Z => n21869);
   U3576 : NOR2_X1 port map( A1 => n11557, A2 => n20186, ZN => n24173);
   U3592 : NAND2_X1 port map( A1 => n20416, A2 => n20413, ZN => n7048);
   U3598 : INV_X2 port map( I => n13853, ZN => n20016);
   U3600 : NAND2_X1 port map( A1 => n20313, A2 => n25455, ZN => n22025);
   U3612 : AOI21_X1 port map( A1 => n2373, A2 => n20018, B => n11259, ZN => 
                           n22596);
   U3621 : AND2_X1 port map( A1 => n11871, A2 => n22835, Z => n9921);
   U3631 : AND2_X1 port map( A1 => n20280, A2 => n7749, Z => n14838);
   U3641 : CLKBUF_X1 port map( I => n3223, Z => n23416);
   U3653 : AND2_X1 port map( A1 => n19788, A2 => n19623, Z => n3391);
   U3658 : NAND2_X1 port map( A1 => n7042, A2 => n7040, ZN => n9992);
   U3674 : OR2_X1 port map( A1 => n2320, A2 => n19623, Z => n21860);
   U3685 : NOR2_X1 port map( A1 => n19519, A2 => n45, ZN => n9188);
   U3691 : NAND2_X1 port map( A1 => n14531, A2 => n19666, ZN => n19788);
   U3705 : NAND2_X1 port map( A1 => n1122, A2 => n14671, ZN => n6451);
   U3723 : NAND2_X1 port map( A1 => n174, A2 => n6976, ZN => n21946);
   U3724 : AND2_X1 port map( A1 => n863, A2 => n19819, Z => n2316);
   U3736 : CLKBUF_X2 port map( I => n19692, Z => n7376);
   U3752 : CLKBUF_X2 port map( I => n735, Z => n22174);
   U3755 : CLKBUF_X2 port map( I => n19806, Z => n24135);
   U3787 : AND2_X1 port map( A1 => n25081, A2 => n9584, Z => n10700);
   U3789 : BUF_X4 port map( I => n10550, Z => n814);
   U3791 : NOR2_X1 port map( A1 => n12030, A2 => n21912, ZN => n12031);
   U3799 : INV_X1 port map( I => n7204, ZN => n22694);
   U3806 : INV_X1 port map( I => n22731, ZN => n22750);
   U3809 : INV_X1 port map( I => n11552, ZN => n4441);
   U3835 : INV_X1 port map( I => n19198, ZN => n22266);
   U3837 : INV_X1 port map( I => n19350, ZN => n1140);
   U3848 : AOI21_X1 port map( A1 => n4224, A2 => n10265, B => n23970, ZN => 
                           n10264);
   U3864 : NAND2_X1 port map( A1 => n8695, A2 => n19025, ZN => n23467);
   U3865 : INV_X1 port map( I => n22346, ZN => n19038);
   U3887 : NAND3_X1 port map( A1 => n19082, A2 => n27258, A3 => n11983, ZN => 
                           n13212);
   U3919 : NOR2_X1 port map( A1 => n14271, A2 => n7533, ZN => n1329);
   U3920 : AND2_X1 port map( A1 => n1716, A2 => n23871, Z => n1376);
   U3921 : INV_X2 port map( I => n9538, ZN => n10801);
   U3956 : NAND2_X1 port map( A1 => n18031, A2 => n18629, ZN => n22559);
   U3962 : NAND2_X1 port map( A1 => n22073, A2 => n18665, ZN => n2109);
   U3971 : INV_X1 port map( I => n7799, ZN => n24460);
   U3981 : NOR2_X1 port map( A1 => n18620, A2 => n18621, ZN => n12245);
   U3986 : INV_X1 port map( I => n18658, ZN => n22450);
   U3989 : NAND2_X1 port map( A1 => n22239, A2 => n10594, ZN => n22238);
   U3994 : NAND2_X1 port map( A1 => n18770, A2 => n457, ZN => n23740);
   U3998 : BUF_X2 port map( I => n18753, Z => n24429);
   U4009 : INV_X1 port map( I => n9150, ZN => n23006);
   U4010 : BUF_X2 port map( I => n12220, Z => n7446);
   U4014 : CLKBUF_X2 port map( I => n12023, Z => n24297);
   U4028 : INV_X1 port map( I => n4505, ZN => n22600);
   U4032 : INV_X1 port map( I => n25865, ZN => n22886);
   U4037 : NAND2_X1 port map( A1 => n23031, A2 => n23030, ZN => n17609);
   U4043 : AOI21_X1 port map( A1 => n23233, A2 => n21943, B => n17783, ZN => 
                           n4505);
   U4049 : NAND2_X1 port map( A1 => n12170, A2 => n17947, ZN => n9079);
   U4057 : NOR2_X1 port map( A1 => n7990, A2 => n23391, ZN => n24307);
   U4061 : NOR2_X1 port map( A1 => n17591, A2 => n3347, ZN => n24076);
   U4065 : INV_X1 port map( I => n23311, ZN => n17966);
   U4066 : NAND2_X1 port map( A1 => n14110, A2 => n14265, ZN => n17674);
   U4072 : BUF_X2 port map( I => n17895, Z => n24479);
   U4082 : OR2_X1 port map( A1 => n13547, A2 => n23696, Z => n10895);
   U4089 : AND2_X1 port map( A1 => n14976, A2 => n17989, Z => n21888);
   U4108 : CLKBUF_X2 port map( I => n18002, Z => n22594);
   U4131 : NOR2_X1 port map( A1 => n16969, A2 => n10568, ZN => n23974);
   U4148 : INV_X1 port map( I => n23797, ZN => n17319);
   U4149 : NAND2_X1 port map( A1 => n17519, A2 => n6608, ZN => n22531);
   U4152 : NAND2_X1 port map( A1 => n23012, A2 => n24038, ZN => n5513);
   U4154 : NAND2_X1 port map( A1 => n17554, A2 => n17222, ZN => n22242);
   U4159 : INV_X1 port map( I => n17435, ZN => n9466);
   U4163 : NAND2_X1 port map( A1 => n14453, A2 => n17557, ZN => n23327);
   U4167 : NAND2_X1 port map( A1 => n14861, A2 => n17569, ZN => n14354);
   U4188 : CLKBUF_X2 port map( I => n8546, Z => n24159);
   U4195 : INV_X2 port map( I => n27662, ZN => n1037);
   U4204 : BUF_X2 port map( I => n28293, Z => n24033);
   U4224 : INV_X1 port map( I => n16857, ZN => n3039);
   U4235 : NAND2_X1 port map( A1 => n23244, A2 => n16615, ZN => n14842);
   U4240 : NAND2_X1 port map( A1 => n5227, A2 => n11204, ZN => n10990);
   U4247 : AND2_X1 port map( A1 => n15061, A2 => n28231, Z => n21831);
   U4254 : CLKBUF_X2 port map( I => n23907, Z => n22201);
   U4256 : OAI21_X1 port map( A1 => n14739, A2 => n5438, B => n9917, ZN => 
                           n22277);
   U4265 : INV_X1 port map( I => n16394, ZN => n22411);
   U4285 : BUF_X4 port map( I => n23128, Z => n7759);
   U4308 : CLKBUF_X2 port map( I => n6617, Z => n24028);
   U4324 : NOR2_X1 port map( A1 => n10091, A2 => n10090, ZN => n24405);
   U4350 : NOR2_X1 port map( A1 => n23221, A2 => n5788, ZN => n23220);
   U4354 : NAND2_X1 port map( A1 => n5790, A2 => n5789, ZN => n23219);
   U4359 : NAND2_X1 port map( A1 => n21786, A2 => n9986, ZN => n10440);
   U4361 : NAND3_X1 port map( A1 => n9892, A2 => n15155, A3 => n15979, ZN => 
                           n8345);
   U4365 : NAND2_X1 port map( A1 => n14684, A2 => n21969, ZN => n22357);
   U4370 : CLKBUF_X2 port map( I => n13435, Z => n24227);
   U4379 : CLKBUF_X2 port map( I => n4990, Z => n21969);
   U4384 : INV_X1 port map( I => n21557, ZN => n23168);
   U4385 : INV_X1 port map( I => n21106, ZN => n24121);
   U4386 : CLKBUF_X2 port map( I => n2799, Z => n24216);
   U4398 : INV_X1 port map( I => Plaintext(84), ZN => n23845);
   U4408 : INV_X1 port map( I => n15936, ZN => n720);
   U4414 : CLKBUF_X2 port map( I => n576, Z => n22910);
   U4423 : OAI21_X1 port map( A1 => n16271, A2 => n23104, B => n15685, ZN => 
                           n16272);
   U4424 : INV_X1 port map( I => n3651, ZN => n23837);
   U4425 : NOR2_X1 port map( A1 => n16274, A2 => n14763, ZN => n11877);
   U4426 : NOR3_X1 port map( A1 => n4751, A2 => n6647, A3 => n16326, ZN => 
                           n23875);
   U4427 : NOR2_X1 port map( A1 => n16181, A2 => n12678, ZN => n5788);
   U4429 : NOR2_X1 port map( A1 => n12116, A2 => n263, ZN => n15765);
   U4430 : OAI21_X1 port map( A1 => n1263, A2 => n14442, B => n841, ZN => n7117
                           );
   U4444 : INV_X2 port map( I => n16207, ZN => n23270);
   U4449 : OAI21_X1 port map( A1 => n14171, A2 => n15822, B => n7540, ZN => 
                           n4116);
   U4452 : NAND2_X1 port map( A1 => n12694, A2 => n21970, ZN => n24341);
   U4460 : INV_X1 port map( I => n8373, ZN => n16672);
   U4462 : NAND2_X1 port map( A1 => n22614, A2 => n6399, ZN => n23277);
   U4483 : OAI21_X1 port map( A1 => n9484, A2 => n835, B => n5081, ZN => n92);
   U4505 : NAND2_X1 port map( A1 => n16408, A2 => n24844, ZN => n16392);
   U4513 : INV_X1 port map( I => n16951, ZN => n22190);
   U4516 : CLKBUF_X4 port map( I => n14878, Z => n23758);
   U4517 : NOR2_X1 port map( A1 => n16488, A2 => n24089, ZN => n22496);
   U4521 : NAND2_X1 port map( A1 => n14739, A2 => n912, ZN => n10112);
   U4524 : AOI21_X1 port map( A1 => n16553, A2 => n12224, B => n4938, ZN => 
                           n7806);
   U4544 : INV_X1 port map( I => n17531, ZN => n21942);
   U4557 : INV_X1 port map( I => n7385, ZN => n6455);
   U4568 : NOR2_X1 port map( A1 => n4465, A2 => n13740, ZN => n3343);
   U4576 : NAND2_X1 port map( A1 => n10821, A2 => n13740, ZN => n14396);
   U4596 : NOR2_X1 port map( A1 => n14861, A2 => n3875, ZN => n23563);
   U4599 : NAND2_X1 port map( A1 => n10563, A2 => n27161, ZN => n5697);
   U4624 : CLKBUF_X2 port map( I => n7108, Z => n23633);
   U4637 : NOR3_X1 port map( A1 => n6425, A2 => n765, A3 => n24509, ZN => n6627
                           );
   U4643 : INV_X1 port map( I => n26614, ZN => n7694);
   U4654 : CLKBUF_X2 port map( I => n9285, Z => n22851);
   U4665 : NOR2_X1 port map( A1 => n17929, A2 => n17635, ZN => n13112);
   U4667 : NOR2_X1 port map( A1 => n17630, A2 => n2068, ZN => n1411);
   U4672 : INV_X1 port map( I => n22253, ZN => n12149);
   U4675 : NAND2_X1 port map( A1 => n23979, A2 => n27947, ZN => n22175);
   U4691 : INV_X1 port map( I => n13478, ZN => n22113);
   U4694 : NAND2_X1 port map( A1 => n4593, A2 => n26939, ZN => n4592);
   U4706 : INV_X1 port map( I => n15488, ZN => n22504);
   U4733 : NAND2_X1 port map( A1 => n10594, A2 => n3062, ZN => n4389);
   U4734 : NAND2_X1 port map( A1 => n6827, A2 => n26277, ZN => n4981);
   U4746 : NAND2_X1 port map( A1 => n26292, A2 => n18661, ZN => n18664);
   U4760 : NAND3_X1 port map( A1 => n11618, A2 => n10116, A3 => n18479, ZN => 
                           n142);
   U4784 : OAI21_X1 port map( A1 => n8944, A2 => n8943, B => n18779, ZN => 
                           n23613);
   U4785 : INV_X1 port map( I => n19145, ZN => n24466);
   U4794 : INV_X1 port map( I => n23559, ZN => n18893);
   U4802 : NAND2_X1 port map( A1 => n2617, A2 => n12584, ZN => n19044);
   U4812 : NOR2_X1 port map( A1 => n23305, A2 => n18794, ZN => n1924);
   U4836 : NAND2_X1 port map( A1 => n18896, A2 => n2541, ZN => n2540);
   U4843 : NAND2_X1 port map( A1 => n18889, A2 => n19062, ZN => n13401);
   U4852 : NAND2_X1 port map( A1 => n4080, A2 => n7970, ZN => n3618);
   U4871 : INV_X2 port map( I => n28446, ZN => n19506);
   U4876 : INV_X1 port map( I => n26833, ZN => n22726);
   U4885 : NOR2_X1 port map( A1 => n754, A2 => n19931, ZN => n9718);
   U4889 : NOR2_X1 port map( A1 => n9812, A2 => n19744, ZN => n150);
   U4901 : INV_X1 port map( I => n19749, ZN => n23462);
   U4903 : NAND2_X1 port map( A1 => n15575, A2 => n19878, ZN => n10243);
   U4904 : NOR2_X1 port map( A1 => n19730, A2 => n6861, ZN => n19595);
   U4913 : CLKBUF_X2 port map( I => n15156, Z => n24196);
   U4924 : CLKBUF_X2 port map( I => n11220, Z => n23977);
   U4925 : NAND2_X1 port map( A1 => n13926, A2 => n14304, ZN => n24390);
   U4941 : AOI21_X1 port map( A1 => n19624, A2 => n19623, B => n12444, ZN => 
                           n23682);
   U4943 : AOI21_X1 port map( A1 => n11454, A2 => n674, B => n1129, ZN => n4395
                           );
   U4948 : INV_X1 port map( I => n976, ZN => n19871);
   U4950 : AOI21_X1 port map( A1 => n9813, A2 => n9812, B => n26625, ZN => 
                           n9811);
   U4995 : INV_X2 port map( I => n20057, ZN => n4225);
   U5004 : INV_X1 port map( I => n14957, ZN => n10399);
   U5029 : AND2_X1 port map( A1 => n19, A2 => n20073, Z => n21865);
   U5050 : INV_X1 port map( I => n20280, ZN => n774);
   U5072 : OAI21_X1 port map( A1 => n9343, A2 => n5, B => n958, ZN => n9342);
   U5100 : NOR2_X1 port map( A1 => n21699, A2 => n21725, ZN => n22654);
   U5103 : NAND2_X1 port map( A1 => n723, A2 => n10588, ZN => n15324);
   U5115 : NAND2_X1 port map( A1 => n3096, A2 => n14679, ZN => n10884);
   U5158 : INV_X1 port map( I => n20964, ZN => n22526);
   U5166 : NAND3_X1 port map( A1 => n21724, A2 => n21721, A3 => n21696, ZN => 
                           n20486);
   U5167 : NOR2_X1 port map( A1 => n23678, A2 => n10588, ZN => n23677);
   U5179 : AOI21_X1 port map( A1 => n20633, A2 => n5540, B => n5806, ZN => 
                           n10087);
   U5184 : NAND2_X1 port map( A1 => n5215, A2 => n5214, ZN => n21234);
   U5190 : AND2_X1 port map( A1 => n934, A2 => n20703, Z => n21872);
   U5193 : NAND3_X1 port map( A1 => n10530, A2 => n12057, A3 => n12054, ZN => 
                           n21042);
   U5206 : AND2_X1 port map( A1 => n23679, A2 => n8742, Z => n22844);
   U5240 : CLKBUF_X1 port map( I => Key(11), Z => n20912);
   U5241 : INV_X1 port map( I => n18003, ZN => n14885);
   U5255 : OR2_X1 port map( A1 => n4630, A2 => n4938, Z => n21799);
   U5265 : AND2_X1 port map( A1 => n1135, A2 => n11444, Z => n21804);
   U5275 : AND2_X1 port map( A1 => n23083, A2 => n14986, Z => n21807);
   U5278 : AND2_X1 port map( A1 => n19631, A2 => n9896, Z => n21812);
   U5283 : XNOR2_X1 port map( A1 => n2515, A2 => n21709, ZN => n21816);
   U5286 : XNOR2_X1 port map( A1 => n21373, A2 => n21037, ZN => n21818);
   U5287 : XNOR2_X1 port map( A1 => n16801, A2 => n14445, ZN => n21819);
   U5293 : XNOR2_X1 port map( A1 => n13469, A2 => n7368, ZN => n21820);
   U5297 : XNOR2_X1 port map( A1 => n3701, A2 => n20967, ZN => n21821);
   U5299 : AND2_X1 port map( A1 => n6314, A2 => n16086, Z => n21822);
   U5310 : AND2_X1 port map( A1 => n7113, A2 => n21800, Z => n21830);
   U5312 : AND2_X1 port map( A1 => n1033, A2 => n1701, Z => n21832);
   U5320 : XNOR2_X1 port map( A1 => n20607, A2 => n22939, ZN => n21838);
   U5343 : OR2_X1 port map( A1 => n3549, A2 => n21445, Z => n21848);
   U5346 : AND2_X1 port map( A1 => n9887, A2 => n5008, Z => n21850);
   U5351 : OR2_X1 port map( A1 => n4639, A2 => n5434, Z => n21852);
   U5360 : XNOR2_X1 port map( A1 => n14006, A2 => n21533, ZN => n21855);
   U5361 : XOR2_X1 port map( A1 => n19462, A2 => n13093, Z => n21856);
   U5363 : XNOR2_X1 port map( A1 => n11794, A2 => n26473, ZN => n21857);
   U5366 : OR2_X1 port map( A1 => n891, A2 => n22396, Z => n21859);
   U5385 : AND2_X1 port map( A1 => n8303, A2 => n14386, Z => n21867);
   U5386 : XOR2_X1 port map( A1 => n20038, A2 => n20538, Z => n21868);
   U5397 : XOR2_X1 port map( A1 => Plaintext(64), A2 => Key(64), Z => n21874);
   U5414 : OR2_X1 port map( A1 => n9653, A2 => n12056, Z => n21875);
   U5423 : XOR2_X1 port map( A1 => Plaintext(30), A2 => Key(30), Z => n21876);
   U5428 : NOR2_X1 port map( A1 => n14611, A2 => n20090, ZN => n21879);
   U5430 : AND2_X1 port map( A1 => n17818, A2 => n8262, Z => n21881);
   U5435 : XNOR2_X1 port map( A1 => Plaintext(10), A2 => Key(10), ZN => n21885)
                           ;
   U5449 : OR2_X1 port map( A1 => n12264, A2 => n12263, Z => n21892);
   U5465 : XNOR2_X1 port map( A1 => n26575, A2 => n21742, ZN => n21894);
   U5469 : NAND4_X1 port map( A1 => n7897, A2 => n7899, A3 => n7900, A4 => 
                           n7898, ZN => n21896);
   U5470 : XNOR2_X1 port map( A1 => n17035, A2 => n26141, ZN => n21897);
   U5475 : INV_X1 port map( I => n10220, ZN => n17268);
   U5480 : XNOR2_X1 port map( A1 => n3751, A2 => n9455, ZN => n21899);
   U5481 : INV_X1 port map( I => n17555, ZN => n14453);
   U5482 : INV_X1 port map( I => n24509, ZN => n17385);
   U5484 : INV_X1 port map( I => n21774, ZN => n17352);
   U5485 : XNOR2_X1 port map( A1 => n9534, A2 => n21336, ZN => n21900);
   U5487 : XNOR2_X1 port map( A1 => n25892, A2 => n14620, ZN => n21902);
   U5488 : XNOR2_X1 port map( A1 => n12532, A2 => n11408, ZN => n21903);
   U5497 : XNOR2_X1 port map( A1 => n6745, A2 => n14588, ZN => n21906);
   U5503 : XNOR2_X1 port map( A1 => n18172, A2 => n20906, ZN => n21908);
   U5505 : XNOR2_X1 port map( A1 => n27816, A2 => n1291, ZN => n21909);
   U5520 : XNOR2_X1 port map( A1 => n19307, A2 => n19308, ZN => n21914);
   U5525 : XNOR2_X1 port map( A1 => n27425, A2 => n14622, ZN => n21917);
   U5547 : XOR2_X1 port map( A1 => n14187, A2 => n21262, Z => n21920);
   U5550 : XNOR2_X1 port map( A1 => n19363, A2 => n14588, ZN => n21922);
   U5552 : XNOR2_X1 port map( A1 => n5913, A2 => n5911, ZN => n21923);
   U5556 : INV_X1 port map( I => n12468, ZN => n10341);
   U5559 : XNOR2_X1 port map( A1 => n13761, A2 => n20435, ZN => n21927);
   U5566 : XNOR2_X1 port map( A1 => n20763, A2 => n20941, ZN => n21928);
   U5569 : XNOR2_X1 port map( A1 => n21241, A2 => n20119, ZN => n21930);
   U5570 : XNOR2_X1 port map( A1 => n13821, A2 => n21156, ZN => n21931);
   U5573 : INV_X1 port map( I => n21502, ZN => n7941);
   U5575 : XNOR2_X1 port map( A1 => n5102, A2 => n1667, ZN => n21934);
   U5579 : XNOR2_X1 port map( A1 => n12320, A2 => n23021, ZN => n21937);
   U5585 : XNOR2_X1 port map( A1 => n17078, A2 => n21039, ZN => n21938);
   U5594 : XOR2_X1 port map( A1 => n17049, A2 => n23779, Z => n21940);
   U5596 : INV_X2 port map( I => n21941, ZN => n8423);
   U5598 : XOR2_X1 port map( A1 => n19176, A2 => n19281, Z => n7520);
   U5611 : OAI21_X2 port map( A1 => n7174, A2 => n19094, B => n7570, ZN => 
                           n24312);
   U5613 : NAND2_X2 port map( A1 => n21944, A2 => n10931, ZN => n14957);
   U5623 : NOR2_X1 port map( A1 => n21946, A2 => n26061, ZN => n21945);
   U5624 : NAND2_X1 port map( A1 => n26758, A2 => n23026, ZN => n15348);
   U5639 : NAND2_X2 port map( A1 => n7788, A2 => n7787, ZN => n19107);
   U5640 : XOR2_X1 port map( A1 => n21948, A2 => n20674, Z => Ciphertext(20));
   U5643 : NAND2_X1 port map( A1 => n23573, A2 => n22466, ZN => n21948);
   U5653 : XOR2_X1 port map( A1 => n20718, A2 => n13803, Z => n5808);
   U5655 : XOR2_X1 port map( A1 => n20424, A2 => n21304, Z => n20718);
   U5664 : XOR2_X1 port map( A1 => n28466, A2 => n6867, Z => n7830);
   U5666 : AOI21_X2 port map( A1 => n6249, A2 => n5558, B => n21949, ZN => 
                           n17094);
   U5690 : XOR2_X1 port map( A1 => n19187, A2 => n21804, Z => n19554);
   U5735 : OAI21_X2 port map( A1 => n15952, A2 => n2523, B => n21959, ZN => 
                           n21958);
   U5748 : NOR2_X1 port map( A1 => n4915, A2 => n4917, ZN => n2779);
   U5752 : NAND2_X2 port map( A1 => n1530, A2 => n21962, ZN => n2016);
   U5753 : NOR2_X2 port map( A1 => n22987, A2 => n21963, ZN => n2710);
   U5757 : XOR2_X1 port map( A1 => n19552, A2 => n3243, Z => n10208);
   U5865 : NAND2_X1 port map( A1 => n23278, A2 => n26638, ZN => n19832);
   U5870 : INV_X1 port map( I => n12693, ZN => n22876);
   U5873 : NAND2_X2 port map( A1 => n8665, A2 => n4969, ZN => n21970);
   U5886 : XOR2_X1 port map( A1 => n3807, A2 => n3809, Z => n17173);
   U5888 : XOR2_X1 port map( A1 => Plaintext(13), A2 => Key(13), Z => n4990);
   U5889 : XOR2_X1 port map( A1 => n4965, A2 => n23589, Z => n15636);
   U5900 : XOR2_X1 port map( A1 => n7709, A2 => n17014, Z => n24060);
   U5933 : OR2_X1 port map( A1 => n11287, A2 => n3953, Z => n19696);
   U5943 : XOR2_X1 port map( A1 => n18109, A2 => n18107, Z => n7476);
   U5952 : NAND2_X2 port map( A1 => n110, A2 => n3627, ZN => n12846);
   U5953 : XOR2_X1 port map( A1 => n9552, A2 => n9620, Z => n9619);
   U5954 : XOR2_X1 port map( A1 => n6101, A2 => n14744, Z => n16854);
   U5956 : XOR2_X1 port map( A1 => n19430, A2 => n19521, Z => n13089);
   U5957 : OAI21_X2 port map( A1 => n13905, A2 => n18923, B => n18435, ZN => 
                           n19430);
   U6006 : AOI22_X2 port map( A1 => n21983, A2 => n9378, B1 => n1541, B2 => 
                           n21064, ZN => n11209);
   U6013 : XOR2_X1 port map( A1 => n22538, A2 => n11040, Z => n5264);
   U6019 : XOR2_X1 port map( A1 => n5499, A2 => n20694, Z => n11037);
   U6023 : NAND3_X2 port map( A1 => n15441, A2 => n8001, A3 => n14028, ZN => 
                           n5499);
   U6032 : XOR2_X1 port map( A1 => n18011, A2 => n17909, Z => n21984);
   U6034 : XOR2_X1 port map( A1 => n18297, A2 => n17910, Z => n21985);
   U6041 : XOR2_X1 port map( A1 => n18008, A2 => n18205, Z => n18163);
   U6050 : INV_X2 port map( I => n6968, ZN => n24286);
   U6062 : XOR2_X1 port map( A1 => n23608, A2 => n6823, Z => n6822);
   U6069 : NAND3_X1 port map( A1 => n21622, A2 => n21627, A3 => n21624, ZN => 
                           n21580);
   U6075 : XOR2_X1 port map( A1 => n19231, A2 => n27358, Z => n21988);
   U6080 : NAND3_X2 port map( A1 => n14772, A2 => n14771, A3 => n13356, ZN => 
                           n17976);
   U6084 : XOR2_X1 port map( A1 => n7948, A2 => n544, Z => n7947);
   U6130 : NAND2_X2 port map( A1 => n23891, A2 => n23283, ZN => n22839);
   U6131 : INV_X1 port map( I => n21994, ZN => n21993);
   U6141 : NAND2_X2 port map( A1 => n10395, A2 => n16362, ZN => n11124);
   U6154 : NOR2_X1 port map( A1 => n8377, A2 => n19079, ZN => n21999);
   U6175 : OAI21_X2 port map( A1 => n18963, A2 => n18964, B => n22001, ZN => 
                           n14272);
   U6192 : INV_X2 port map( I => n20625, ZN => n939);
   U6194 : NAND2_X2 port map( A1 => n20486, A2 => n10284, ZN => n20625);
   U6200 : XOR2_X1 port map( A1 => n8132, A2 => n22005, Z => n589);
   U6201 : INV_X1 port map( I => n14616, ZN => n22005);
   U6206 : XOR2_X1 port map( A1 => n11990, A2 => n9656, Z => n4262);
   U6223 : XOR2_X1 port map( A1 => n22008, A2 => n919, Z => Ciphertext(33));
   U6232 : XOR2_X1 port map( A1 => n21181, A2 => n11574, Z => n22010);
   U6251 : INV_X2 port map( I => n22018, ZN => n22840);
   U6256 : XOR2_X1 port map( A1 => n8902, A2 => n8903, Z => n22018);
   U6261 : XOR2_X1 port map( A1 => n6085, A2 => n23414, Z => n24010);
   U6308 : XOR2_X1 port map( A1 => n18162, A2 => n18302, Z => n15109);
   U6316 : OAI21_X2 port map( A1 => n8090, A2 => n7687, B => n22022, ZN => 
                           n3312);
   U6347 : XOR2_X1 port map( A1 => n4833, A2 => n21533, Z => n22102);
   U6383 : XOR2_X1 port map( A1 => n3830, A2 => n23818, Z => n22647);
   U6384 : INV_X1 port map( I => n6756, ZN => n10936);
   U6385 : NAND2_X1 port map( A1 => n6756, A2 => n22027, ZN => n6832);
   U6396 : XOR2_X1 port map( A1 => n19272, A2 => n980, Z => n19322);
   U6455 : INV_X2 port map( I => n12046, ZN => n20997);
   U6457 : XOR2_X1 port map( A1 => n22036, A2 => n21708, Z => Ciphertext(182));
   U6486 : XOR2_X1 port map( A1 => n19379, A2 => n19376, Z => n23717);
   U6488 : XOR2_X1 port map( A1 => n13918, A2 => n19532, Z => n19376);
   U6492 : AOI21_X2 port map( A1 => n22040, A2 => n20789, B => n20788, ZN => 
                           n20803);
   U6495 : NOR2_X1 port map( A1 => n19889, A2 => n7240, ZN => n3986);
   U6497 : XOR2_X1 port map( A1 => n22041, A2 => n21705, Z => Ciphertext(181));
   U6498 : OAI22_X1 port map( A1 => n8444, A2 => n9267, B1 => n21704, B2 => 
                           n21706, ZN => n22041);
   U6513 : XOR2_X1 port map( A1 => n5971, A2 => n5972, Z => n22178);
   U6514 : NAND2_X1 port map( A1 => n2730, A2 => n9875, ZN => n8772);
   U6524 : XOR2_X1 port map( A1 => n4996, A2 => n22044, Z => n12208);
   U6525 : XOR2_X1 port map( A1 => n27430, A2 => n6563, Z => n22044);
   U6540 : NAND2_X2 port map( A1 => n22051, A2 => n25411, ZN => n1416);
   U6549 : NAND2_X2 port map( A1 => n1418, A2 => n24294, ZN => n22051);
   U6566 : NAND2_X1 port map( A1 => n18785, A2 => n25331, ZN => n7095);
   U6570 : NAND2_X2 port map( A1 => n13042, A2 => n13655, ZN => n14663);
   U6585 : NAND2_X2 port map( A1 => n11611, A2 => n11613, ZN => n19560);
   U6586 : XOR2_X1 port map( A1 => n22055, A2 => n918, Z => Ciphertext(26));
   U6593 : INV_X4 port map( I => n5909, ZN => n20338);
   U6595 : NAND2_X2 port map( A1 => n22575, A2 => n9719, ZN => n5909);
   U6601 : XOR2_X1 port map( A1 => n7103, A2 => n25333, Z => n22500);
   U6613 : INV_X1 port map( I => n9840, ZN => n23001);
   U6631 : AOI22_X1 port map( A1 => n13861, A2 => n27359, B1 => n13862, B2 => 
                           n17952, ZN => n15102);
   U6653 : OR2_X1 port map( A1 => n10704, A2 => n8717, Z => n19638);
   U6688 : NOR2_X1 port map( A1 => n2023, A2 => n13147, ZN => n12479);
   U6697 : XOR2_X1 port map( A1 => n22069, A2 => n10056, Z => n12222);
   U6740 : OAI21_X2 port map( A1 => n17491, A2 => n830, B => n7456, ZN => 
                           n22085);
   U6775 : XOR2_X1 port map( A1 => n8608, A2 => n18105, Z => n22077);
   U6785 : XOR2_X1 port map( A1 => n22080, A2 => n2105, Z => n23576);
   U6786 : XOR2_X1 port map( A1 => n22081, A2 => n25941, Z => n22080);
   U6787 : NAND2_X1 port map( A1 => n22082, A2 => n14282, ZN => n23822);
   U6804 : NAND2_X1 port map( A1 => n23150, A2 => n18409, ZN => n18368);
   U6807 : NAND3_X1 port map( A1 => n4780, A2 => n26277, A3 => n4661, ZN => 
                           n23150);
   U6817 : XOR2_X1 port map( A1 => n18218, A2 => n8505, Z => n3582);
   U6883 : OR2_X1 port map( A1 => n23842, A2 => n14228, Z => n16121);
   U6922 : NAND3_X2 port map( A1 => n12164, A2 => n12561, A3 => n3207, ZN => 
                           n10149);
   U6932 : NAND2_X2 port map( A1 => n19574, A2 => n11369, ZN => n19095);
   U6934 : NOR2_X2 port map( A1 => n867, A2 => n12941, ZN => n19574);
   U6944 : XOR2_X1 port map( A1 => n2306, A2 => n21370, Z => n5406);
   U6952 : NAND2_X2 port map( A1 => n3972, A2 => n7811, ZN => n3971);
   U6956 : NAND2_X2 port map( A1 => n9402, A2 => n21025, ZN => n3972);
   U6965 : NOR2_X2 port map( A1 => n18243, A2 => n7705, ZN => n3557);
   U6967 : NAND3_X1 port map( A1 => n8181, A2 => n27914, A3 => n26578, ZN => 
                           n16451);
   U6975 : XOR2_X1 port map( A1 => n5022, A2 => n5021, Z => n5020);
   U6978 : XOR2_X1 port map( A1 => n20438, A2 => n23500, Z => n22091);
   U6982 : OAI21_X1 port map( A1 => n28499, A2 => n19133, B => n18970, ZN => 
                           n7232);
   U7021 : XOR2_X1 port map( A1 => n6616, A2 => n4500, Z => n3594);
   U7026 : OR2_X1 port map( A1 => n14860, A2 => n11905, Z => n12426);
   U7032 : XOR2_X1 port map( A1 => n27371, A2 => n21090, Z => n2477);
   U7038 : NOR2_X2 port map( A1 => n4739, A2 => n24315, ZN => n5830);
   U7056 : XOR2_X1 port map( A1 => n20385, A2 => n14144, Z => n20764);
   U7059 : OAI21_X2 port map( A1 => n13100, A2 => n20473, B => n13099, ZN => 
                           n20385);
   U7062 : NOR2_X1 port map( A1 => n22097, A2 => n5736, ZN => n22946);
   U7063 : AOI21_X1 port map( A1 => n8162, A2 => n8163, B => n6037, ZN => 
                           n22097);
   U7074 : NOR2_X1 port map( A1 => n13763, A2 => n13866, ZN => n13865);
   U7084 : NAND2_X1 port map( A1 => n8057, A2 => n20164, ZN => n22099);
   U7105 : XOR2_X1 port map( A1 => n21157, A2 => n22102, Z => n1613);
   U7121 : XOR2_X1 port map( A1 => n6946, A2 => n18278, Z => n3331);
   U7124 : XOR2_X1 port map( A1 => n8448, A2 => n3869, Z => n2750);
   U7154 : XOR2_X1 port map( A1 => n27087, A2 => n7408, Z => n22108);
   U7157 : AND2_X1 port map( A1 => n13467, A2 => n5523, Z => n18688);
   U7174 : NAND2_X1 port map( A1 => n2254, A2 => n4934, ZN => n22579);
   U7175 : NAND2_X2 port map( A1 => n3825, A2 => n23765, ZN => n2254);
   U7181 : NOR3_X1 port map( A1 => n7498, A2 => n10081, A3 => n10985, ZN => 
                           n24059);
   U7194 : OAI21_X2 port map( A1 => n13688, A2 => n11206, B => n19713, ZN => 
                           n6511);
   U7199 : XOR2_X1 port map( A1 => n11684, A2 => n14591, Z => n17056);
   U7233 : NAND3_X1 port map( A1 => n13597, A2 => n2617, A3 => n19122, ZN => 
                           n22115);
   U7243 : XOR2_X1 port map( A1 => n1019, A2 => n698, Z => n24134);
   U7252 : NAND2_X2 port map( A1 => n16595, A2 => n16596, ZN => n16924);
   U7253 : INV_X2 port map( I => n22116, ZN => n21388);
   U7260 : NOR2_X1 port map( A1 => n18763, A2 => n5115, ZN => n22118);
   U7270 : NAND2_X1 port map( A1 => n27367, A2 => n12726, ZN => n4869);
   U7271 : NAND2_X2 port map( A1 => n15777, A2 => n15778, ZN => n11238);
   U7274 : XOR2_X1 port map( A1 => n23704, A2 => n8431, Z => n22121);
   U7279 : INV_X2 port map( I => n22122, ZN => n9131);
   U7321 : INV_X2 port map( I => n17840, ZN => n22126);
   U7338 : XOR2_X1 port map( A1 => n9802, A2 => n10056, Z => n17718);
   U7349 : XOR2_X1 port map( A1 => n6595, A2 => n6594, Z => n22130);
   U7362 : OR2_X1 port map( A1 => n10627, A2 => n7085, Z => n21568);
   U7364 : NAND2_X1 port map( A1 => n22203, A2 => n23455, ZN => n24138);
   U7370 : AOI21_X2 port map( A1 => n13788, A2 => n3009, B => n24062, ZN => 
                           n3033);
   U7372 : NOR2_X2 port map( A1 => n8816, A2 => n8817, ZN => n10851);
   U7379 : NAND2_X1 port map( A1 => n22184, A2 => n21608, ZN => n13889);
   U7381 : OAI22_X2 port map( A1 => n18394, A2 => n18393, B1 => n19151, B2 => 
                           n18395, ZN => n19290);
   U7455 : XOR2_X1 port map( A1 => n11681, A2 => n22139, Z => n18482);
   U7456 : XOR2_X1 port map( A1 => n17753, A2 => n3640, Z => n22139);
   U7480 : NAND2_X1 port map( A1 => n9381, A2 => n8459, ZN => n22142);
   U7482 : NAND2_X2 port map( A1 => n11614, A2 => n22143, ZN => n12331);
   U7483 : NAND2_X1 port map( A1 => n7427, A2 => n14277, ZN => n22143);
   U7501 : NAND2_X2 port map( A1 => n22707, A2 => n22144, ZN => n13925);
   U7504 : AND2_X1 port map( A1 => n27734, A2 => n9978, Z => n10111);
   U7512 : XOR2_X1 port map( A1 => n16856, A2 => n11917, Z => n22146);
   U7525 : AOI21_X2 port map( A1 => n2139, A2 => n9827, B => n2138, ZN => 
                           n10920);
   U7532 : NAND2_X2 port map( A1 => n5586, A2 => n5585, ZN => n14237);
   U7555 : OAI21_X2 port map( A1 => n3203, A2 => n15633, B => n15634, ZN => 
                           n5118);
   U7559 : NAND2_X1 port map( A1 => n12584, A2 => n23575, ZN => n18573);
   U7594 : NAND2_X1 port map( A1 => n13247, A2 => n14103, ZN => n17391);
   U7596 : XOR2_X1 port map( A1 => n10524, A2 => n16898, Z => n13247);
   U7602 : NOR2_X1 port map( A1 => n9683, A2 => n5118, ZN => n14739);
   U7603 : XNOR2_X1 port map( A1 => n27384, A2 => n18236, ZN => n22265);
   U7622 : XOR2_X1 port map( A1 => n16829, A2 => n15062, Z => n22158);
   U7629 : BUF_X4 port map( I => n10533, Z => n6022);
   U7637 : INV_X1 port map( I => n9758, ZN => n22163);
   U7663 : NAND3_X1 port map( A1 => n1255, A2 => n458, A3 => n3729, ZN => 
                           n23804);
   U7665 : OAI21_X2 port map( A1 => n2709, A2 => n9288, B => n2708, ZN => 
                           n23053);
   U7690 : NOR2_X2 port map( A1 => n12629, A2 => n20341, ZN => n20038);
   U7697 : OAI22_X2 port map( A1 => n13656, A2 => n5584, B1 => n5583, B2 => 
                           n13657, ZN => n18125);
   U7712 : XOR2_X1 port map( A1 => n15662, A2 => n15661, Z => n7658);
   U7722 : NAND2_X1 port map( A1 => n13990, A2 => n27926, ZN => n22171);
   U7730 : NAND2_X1 port map( A1 => n13989, A2 => n16332, ZN => n22172);
   U7745 : NAND2_X2 port map( A1 => n22176, A2 => n22175, ZN => n11126);
   U7757 : XOR2_X1 port map( A1 => n19562, A2 => n15126, Z => n19315);
   U7760 : XOR2_X1 port map( A1 => n24325, A2 => n22761, Z => n14669);
   U7761 : XOR2_X1 port map( A1 => n5969, A2 => n22178, Z => n5985);
   U7802 : NAND2_X2 port map( A1 => n23679, A2 => n8742, ZN => n11622);
   U7804 : INV_X1 port map( I => n15474, ZN => n22184);
   U7805 : NAND2_X1 port map( A1 => n15470, A2 => n9611, ZN => n15474);
   U7811 : XOR2_X1 port map( A1 => n10986, A2 => n21368, Z => n5144);
   U7817 : NAND2_X2 port map( A1 => n10168, A2 => n15368, ZN => n11815);
   U7821 : OAI21_X2 port map( A1 => n22272, A2 => n13289, B => n22185, ZN => 
                           n18791);
   U7831 : AND2_X2 port map( A1 => n22446, A2 => n22819, Z => n5759);
   U7832 : XOR2_X1 port map( A1 => n16991, A2 => n22190, Z => n10490);
   U7833 : AND2_X1 port map( A1 => n16100, A2 => n9768, Z => n10505);
   U7872 : NAND2_X2 port map( A1 => n22194, A2 => n15172, ZN => n15429);
   U7874 : NAND2_X2 port map( A1 => n21863, A2 => n5573, ZN => n20154);
   U7880 : XOR2_X1 port map( A1 => n22196, A2 => n23572, Z => n6327);
   U7890 : NAND2_X1 port map( A1 => n993, A2 => n9268, ZN => n23175);
   U7898 : INV_X2 port map( I => n7599, ZN => n22197);
   U7902 : OAI21_X2 port map( A1 => n2696, A2 => n2695, B => n10187, ZN => 
                           n2694);
   U7925 : XOR2_X1 port map( A1 => n28521, A2 => n14576, Z => n10755);
   U7939 : XOR2_X1 port map( A1 => n19551, A2 => n15220, Z => n22198);
   U7946 : XOR2_X1 port map( A1 => n26848, A2 => n20344, Z => n15456);
   U7982 : XOR2_X1 port map( A1 => n20285, A2 => n20284, Z => n24331);
   U7989 : XOR2_X1 port map( A1 => n16826, A2 => n12481, Z => n16964);
   U7997 : NAND2_X2 port map( A1 => n12213, A2 => n12210, ZN => n12481);
   U8006 : NOR2_X2 port map( A1 => n12357, A2 => n10720, ZN => n11027);
   U8036 : AND2_X1 port map( A1 => n17868, A2 => n17867, Z => n23357);
   U8046 : INV_X1 port map( I => n6909, ZN => n22205);
   U8055 : AND2_X1 port map( A1 => n17710, A2 => n12943, Z => n22206);
   U8069 : INV_X2 port map( I => n21388, ZN => n22212);
   U8070 : AND2_X1 port map( A1 => n4143, A2 => n22212, Z => n6320);
   U8077 : NAND2_X1 port map( A1 => n13775, A2 => n19774, ZN => n22214);
   U8113 : NOR2_X2 port map( A1 => n22290, A2 => n2735, ZN => n6725);
   U8162 : OAI21_X2 port map( A1 => n21807, A2 => n7247, B => n9344, ZN => 
                           n18102);
   U8168 : AOI21_X2 port map( A1 => n17666, A2 => n8614, B => n25508, ZN => 
                           n8613);
   U8179 : XOR2_X1 port map( A1 => n1142, A2 => n9063, Z => n7329);
   U8186 : OAI21_X1 port map( A1 => n23274, A2 => n21110, B => n13021, ZN => 
                           n3576);
   U8187 : XOR2_X1 port map( A1 => n22226, A2 => n21635, Z => Ciphertext(163));
   U8191 : AOI22_X1 port map( A1 => n23069, A2 => n21632, B1 => n21637, B2 => 
                           n21634, ZN => n22226);
   U8226 : XOR2_X1 port map( A1 => n4618, A2 => n28287, Z => n10312);
   U8267 : AOI21_X2 port map( A1 => n780, A2 => n1165, B => n22240, ZN => n3325
                           );
   U8268 : OAI22_X2 port map( A1 => n22241, A2 => n23510, B1 => n17320, B2 => 
                           n1617, ZN => n12094);
   U8271 : NAND3_X2 port map( A1 => n22289, A2 => n8517, A3 => n22242, ZN => 
                           n17887);
   U8274 : INV_X2 port map( I => n16155, ZN => n9095);
   U8288 : XOR2_X1 port map( A1 => n9023, A2 => Key(136), Z => n16155);
   U8294 : XOR2_X1 port map( A1 => n23928, A2 => n21191, Z => n20501);
   U8303 : AOI21_X2 port map( A1 => n4371, A2 => n13732, B => n21834, ZN => 
                           n23928);
   U8405 : BUF_X2 port map( I => n24525, Z => n166);
   U8415 : XOR2_X1 port map( A1 => n20511, A2 => n5682, Z => n20034);
   U8419 : AOI21_X2 port map( A1 => n9192, A2 => n14957, B => n3728, ZN => 
                           n20511);
   U8422 : XOR2_X1 port map( A1 => n18116, A2 => n18305, Z => n18026);
   U8423 : AOI22_X2 port map( A1 => n4071, A2 => n17789, B1 => n18330, B2 => 
                           n4288, ZN => n18305);
   U8424 : XOR2_X1 port map( A1 => n18104, A2 => n10327, Z => n5913);
   U8425 : XOR2_X1 port map( A1 => n14659, A2 => n18029, Z => n18104);
   U8429 : AOI22_X2 port map( A1 => n22247, A2 => n47, B1 => n23564, B2 => 
                           n6389, ZN => n6388);
   U8432 : NAND2_X2 port map( A1 => n8928, A2 => n8927, ZN => n9123);
   U8443 : NAND2_X2 port map( A1 => n22252, A2 => n6400, ZN => n17070);
   U8458 : NAND2_X1 port map( A1 => n3576, A2 => n929, ZN => n22256);
   U8485 : NAND2_X1 port map( A1 => n7148, A2 => n11329, ZN => n7294);
   U8494 : XNOR2_X1 port map( A1 => n11501, A2 => n19524, ZN => n22731);
   U8504 : NOR2_X2 port map( A1 => n22259, A2 => n82, ZN => n21609);
   U8506 : NAND2_X2 port map( A1 => n9734, A2 => n13819, ZN => n17676);
   U8525 : XOR2_X1 port map( A1 => n17009, A2 => n16797, Z => n5782);
   U8527 : XOR2_X1 port map( A1 => n16853, A2 => n22818, Z => n17009);
   U8534 : INV_X2 port map( I => n20395, ZN => n20730);
   U8550 : INV_X2 port map( I => n20665, ZN => n848);
   U8553 : NAND3_X2 port map( A1 => n6735, A2 => n6734, A3 => n20638, ZN => 
                           n20665);
   U8566 : XOR2_X1 port map( A1 => n14046, A2 => n22264, Z => n5523);
   U8567 : XOR2_X1 port map( A1 => n22265, A2 => n22773, Z => n22264);
   U8575 : XOR2_X1 port map( A1 => n6272, A2 => n18104, Z => n22267);
   U8599 : AOI21_X1 port map( A1 => n9702, A2 => n21692, B => n9057, ZN => 
                           n7977);
   U8613 : NAND2_X2 port map( A1 => n22273, A2 => n5518, ZN => n12626);
   U8623 : NAND2_X2 port map( A1 => n7023, A2 => n7553, ZN => n17750);
   U8625 : XOR2_X1 port map( A1 => n19539, A2 => n7250, Z => n2551);
   U8629 : XOR2_X1 port map( A1 => n21304, A2 => n1301, Z => n521);
   U8630 : NAND2_X2 port map( A1 => n11228, A2 => n11229, ZN => n21304);
   U8637 : AND2_X1 port map( A1 => n27044, A2 => n1772, Z => n22649);
   U8648 : NAND2_X1 port map( A1 => n23926, A2 => n17241, ZN => n22274);
   U8674 : NAND2_X2 port map( A1 => n11854, A2 => n20224, ZN => n20136);
   U8694 : OAI21_X2 port map( A1 => n15523, A2 => n14361, B => n1184, ZN => 
                           n22282);
   U8710 : XOR2_X1 port map( A1 => n19464, A2 => n21856, Z => n24529);
   U8733 : XOR2_X1 port map( A1 => n12717, A2 => n27400, Z => n7976);
   U8741 : XOR2_X1 port map( A1 => n15726, A2 => n19628, Z => n13359);
   U8744 : XOR2_X1 port map( A1 => n22287, A2 => n19462, Z => n22423);
   U8747 : OR2_X1 port map( A1 => n8423, A2 => n17293, Z => n6462);
   U8749 : OAI21_X1 port map( A1 => n19044, A2 => n12583, B => n24239, ZN => 
                           n2639);
   U8753 : NAND2_X2 port map( A1 => n5570, A2 => n22288, ZN => n7057);
   U8759 : NOR2_X2 port map( A1 => n23867, A2 => n22961, ZN => n15290);
   U8782 : XOR2_X1 port map( A1 => n1364, A2 => n1363, Z => n7463);
   U8793 : XOR2_X1 port map( A1 => n3038, A2 => n21877, Z => n22927);
   U8794 : XOR2_X1 port map( A1 => n3456, A2 => n4178, Z => n8564);
   U8795 : XNOR2_X1 port map( A1 => n17030, A2 => n11189, ZN => n22440);
   U8796 : NAND2_X1 port map( A1 => n13050, A2 => n4064, ZN => n13250);
   U8808 : XOR2_X1 port map( A1 => n1742, A2 => n13777, Z => n1741);
   U8825 : OR2_X1 port map( A1 => n10251, A2 => n18633, Z => n3454);
   U8831 : NAND2_X1 port map( A1 => n20225, A2 => n11854, ZN => n22303);
   U8838 : NAND2_X1 port map( A1 => n22306, A2 => n22305, ZN => n17870);
   U8859 : OAI22_X1 port map( A1 => n7193, A2 => n13471, B1 => n13474, B2 => 
                           n4057, ZN => n13470);
   U8868 : OR2_X1 port map( A1 => n26578, A2 => n8181, Z => n3070);
   U8889 : INV_X2 port map( I => n22314, ZN => n16136);
   U8891 : XNOR2_X1 port map( A1 => Plaintext(55), A2 => Key(55), ZN => n22314)
                           ;
   U8893 : XOR2_X1 port map( A1 => n19522, A2 => n22315, Z => n600);
   U8895 : INV_X1 port map( I => n14556, ZN => n22315);
   U8896 : NAND2_X2 port map( A1 => n1815, A2 => n1819, ZN => n19522);
   U8898 : AND2_X1 port map( A1 => n16678, A2 => n23107, Z => n12525);
   U8909 : NAND2_X2 port map( A1 => n7911, A2 => n2563, ZN => n22345);
   U8941 : INV_X2 port map( I => n9053, ZN => n17559);
   U8972 : XOR2_X1 port map( A1 => n23500, A2 => n20718, Z => n20722);
   U8973 : NAND3_X1 port map( A1 => n14409, A2 => n944, A3 => n20180, ZN => 
                           n6852);
   U8975 : XOR2_X1 port map( A1 => n22322, A2 => n19433, Z => n13107);
   U8976 : XOR2_X1 port map( A1 => n22169, A2 => n19432, Z => n22322);
   U8983 : XOR2_X1 port map( A1 => n21311, A2 => n23928, Z => n20533);
   U8986 : NOR2_X2 port map( A1 => n6850, A2 => n6849, ZN => n21083);
   U9024 : NAND2_X2 port map( A1 => n23431, A2 => n19015, ZN => n18808);
   U9040 : XOR2_X1 port map( A1 => n20420, A2 => n22331, Z => n8343);
   U9041 : XOR2_X1 port map( A1 => n27604, A2 => n21426, Z => n22331);
   U9059 : NAND3_X1 port map( A1 => n5009, A2 => n21507, A3 => n951, ZN => 
                           n5509);
   U9083 : NOR2_X2 port map( A1 => n22333, A2 => n15915, ZN => n16426);
   U9090 : OR2_X1 port map( A1 => n14894, A2 => n7668, Z => n23537);
   U9094 : NAND2_X1 port map( A1 => n13011, A2 => n102, ZN => n22589);
   U9095 : AOI21_X2 port map( A1 => n22937, A2 => n12426, B => n13525, ZN => 
                           n102);
   U9098 : OR2_X1 port map( A1 => n14792, A2 => n4898, Z => n6209);
   U9117 : NOR2_X2 port map( A1 => n9312, A2 => n9311, ZN => n4175);
   U9120 : INV_X2 port map( I => n22335, ZN => n24070);
   U9121 : XOR2_X1 port map( A1 => n8685, A2 => n536, Z => n22335);
   U9142 : NOR2_X1 port map( A1 => n26059, A2 => n10217, ZN => n23823);
   U9158 : NAND2_X2 port map( A1 => n10250, A2 => n22339, ZN => n10249);
   U9177 : XOR2_X1 port map( A1 => n21854, A2 => n3880, Z => n22341);
   U9181 : XOR2_X1 port map( A1 => n15647, A2 => n3107, Z => n5517);
   U9193 : OAI21_X1 port map( A1 => n12145, A2 => n14282, B => n10593, ZN => 
                           n11822);
   U9221 : XOR2_X1 port map( A1 => n21903, A2 => n14073, Z => n22347);
   U9236 : XOR2_X1 port map( A1 => n6308, A2 => n21920, Z => n22354);
   U9247 : INV_X4 port map( I => n16429, ZN => n22614);
   U9252 : NAND3_X1 port map( A1 => n17424, A2 => n21754, A3 => n1231, ZN => 
                           n22658);
   U9268 : NAND2_X2 port map( A1 => n22358, A2 => n14294, ZN => n1791);
   U9275 : NAND2_X1 port map( A1 => n23771, A2 => n27454, ZN => n19362);
   U9290 : OAI21_X2 port map( A1 => n22319, A2 => n24702, B => n16226, ZN => 
                           n11878);
   U9313 : XOR2_X1 port map( A1 => n7284, A2 => n5547, Z => n11021);
   U9347 : NAND2_X2 port map( A1 => n22371, A2 => n22370, ZN => n2523);
   U9380 : NAND2_X2 port map( A1 => n2753, A2 => n2752, ZN => n17894);
   U9381 : NAND4_X2 port map( A1 => n7716, A2 => n4770, A3 => n7715, A4 => 
                           n22380, ZN => n7108);
   U9402 : NAND2_X2 port map( A1 => n22383, A2 => n9599, ZN => n6089);
   U9412 : AOI21_X2 port map( A1 => n727, A2 => n2895, B => n713, ZN => n17691)
                           ;
   U9448 : NAND2_X2 port map( A1 => n2218, A2 => n28442, ZN => n22386);
   U9470 : INV_X2 port map( I => n24373, ZN => n17447);
   U9473 : XOR2_X1 port map( A1 => n21908, A2 => n17707, Z => n22392);
   U9490 : XOR2_X1 port map( A1 => n22393, A2 => n14955, Z => n15366);
   U9544 : INV_X2 port map( I => n20065, ZN => n22398);
   U9554 : XOR2_X1 port map( A1 => n22401, A2 => n7315, Z => n687);
   U9563 : XOR2_X1 port map( A1 => n15402, A2 => n15403, Z => n22401);
   U9579 : XOR2_X1 port map( A1 => n3869, A2 => n1354, Z => n22402);
   U9591 : INV_X2 port map( I => n22404, ZN => n4143);
   U9592 : XNOR2_X1 port map( A1 => n10328, A2 => n385, ZN => n22404);
   U9598 : XOR2_X1 port map( A1 => n16751, A2 => n22405, Z => n2964);
   U9603 : XOR2_X1 port map( A1 => n2225, A2 => n21164, Z => n22405);
   U9609 : OAI21_X2 port map( A1 => n1169, A2 => n650, B => n8703, ZN => n4445)
                           ;
   U9662 : INV_X2 port map( I => n14914, ZN => n21325);
   U9713 : NOR2_X2 port map( A1 => n20393, A2 => n9440, ZN => n21318);
   U9746 : OAI21_X2 port map( A1 => n24627, A2 => n22418, B => n8901, ZN => 
                           n11600);
   U9754 : NAND2_X2 port map( A1 => n21276, A2 => n3221, ZN => n6066);
   U9768 : INV_X2 port map( I => n4140, ZN => n22421);
   U9777 : NAND3_X2 port map( A1 => n12337, A2 => n10743, A3 => n12336, ZN => 
                           n16929);
   U9778 : NAND2_X1 port map( A1 => n22000, A2 => n2890, ZN => n13146);
   U9789 : XOR2_X1 port map( A1 => n5417, A2 => n22424, Z => n18772);
   U9790 : XOR2_X1 port map( A1 => n18079, A2 => n638, Z => n22424);
   U9798 : NAND2_X2 port map( A1 => n5176, A2 => n790, ZN => n22425);
   U9802 : INV_X4 port map( I => n14595, ZN => n23968);
   U9803 : XOR2_X1 port map( A1 => n12091, A2 => n16473, Z => n12090);
   U9836 : XOR2_X1 port map( A1 => n27447, A2 => n1638, Z => n4314);
   U9849 : XOR2_X1 port map( A1 => n7914, A2 => n7916, Z => n6574);
   U9859 : NAND2_X2 port map( A1 => n8206, A2 => n8207, ZN => n16858);
   U9864 : INV_X2 port map( I => n20761, ZN => n24325);
   U9867 : NAND2_X2 port map( A1 => n10288, A2 => n10287, ZN => n20761);
   U9897 : XOR2_X1 port map( A1 => n16809, A2 => n17088, Z => n17140);
   U9898 : INV_X1 port map( I => n14611, ZN => n20101);
   U9916 : XOR2_X1 port map( A1 => n7812, A2 => n10320, Z => n6202);
   U9932 : XOR2_X1 port map( A1 => n22487, A2 => n14996, Z => n22432);
   U9949 : INV_X4 port map( I => n8988, ZN => n13502);
   U9956 : XOR2_X1 port map( A1 => n19431, A2 => n19542, Z => n8863);
   U9968 : NOR2_X2 port map( A1 => n22439, A2 => n18000, ZN => n11555);
   U9972 : XOR2_X1 port map( A1 => n10826, A2 => n22440, Z => n23448);
   U10026 : XOR2_X1 port map( A1 => n5772, A2 => n22444, Z => n5771);
   U10027 : XOR2_X1 port map( A1 => n21182, A2 => n12021, Z => n22444);
   U10030 : NOR2_X2 port map( A1 => n22445, A2 => n11771, ZN => n17898);
   U10034 : NOR2_X1 port map( A1 => n12719, A2 => n12720, ZN => n22445);
   U10068 : OAI21_X2 port map( A1 => n4291, A2 => n4292, B => n22449, ZN => 
                           n19163);
   U10080 : NAND2_X2 port map( A1 => n22451, A2 => n13020, ZN => n13021);
   U10093 : NAND2_X1 port map( A1 => n20473, A2 => n20472, ZN => n12020);
   U10112 : AOI22_X2 port map( A1 => n22460, A2 => n15471, B1 => n6262, B2 => 
                           n28095, ZN => n20234);
   U10148 : XOR2_X1 port map( A1 => n22463, A2 => n4372, Z => n3157);
   U10163 : XOR2_X1 port map( A1 => n13443, A2 => n11680, Z => n6705);
   U10165 : NAND2_X1 port map( A1 => n20673, A2 => n7698, ZN => n22466);
   U10194 : XOR2_X1 port map( A1 => n10234, A2 => n8, Z => n22470);
   U10209 : NAND2_X2 port map( A1 => n2094, A2 => n2093, ZN => n2095);
   U10214 : NAND2_X2 port map( A1 => n22475, A2 => n28501, ZN => n10258);
   U10215 : NAND2_X2 port map( A1 => n11944, A2 => n11943, ZN => n22475);
   U10238 : INV_X2 port map( I => n22478, ZN => n11089);
   U10245 : OAI21_X1 port map( A1 => n15189, A2 => n17489, B => n1039, ZN => 
                           n13198);
   U10271 : NAND2_X2 port map( A1 => n18747, A2 => n18639, ZN => n22482);
   U10273 : NOR2_X1 port map( A1 => n4538, A2 => n4540, ZN => n22944);
   U10287 : NAND2_X1 port map( A1 => n438, A2 => n21640, ZN => n15219);
   U10305 : NOR2_X1 port map( A1 => n21630, A2 => n21666, ZN => n22483);
   U10321 : NOR2_X2 port map( A1 => n17950, A2 => n17757, ZN => n23978);
   U10347 : AOI21_X1 port map( A1 => n22544, A2 => n7298, B => n1026, ZN => 
                           n1569);
   U10348 : NAND2_X2 port map( A1 => n5696, A2 => n22489, ZN => n3438);
   U10358 : INV_X2 port map( I => n22490, ZN => n9252);
   U10362 : XOR2_X1 port map( A1 => n16901, A2 => n11762, Z => n22490);
   U10370 : OR2_X2 port map( A1 => n6459, A2 => n4610, Z => n17933);
   U10371 : XOR2_X1 port map( A1 => n9514, A2 => n9510, Z => n15501);
   U10372 : NOR2_X2 port map( A1 => n7331, A2 => n7333, ZN => n23842);
   U10380 : NOR2_X2 port map( A1 => n23256, A2 => n14626, ZN => n23255);
   U10394 : AND2_X1 port map( A1 => n13896, A2 => n18549, Z => n10152);
   U10398 : XOR2_X1 port map( A1 => n8077, A2 => n8079, Z => n10923);
   U10404 : XOR2_X1 port map( A1 => n22493, A2 => n10466, Z => n10465);
   U10409 : XOR2_X1 port map( A1 => n21179, A2 => n10248, Z => n22493);
   U10443 : INV_X2 port map( I => n9979, ZN => n20598);
   U10483 : XOR2_X1 port map( A1 => n22500, A2 => n2649, Z => n2648);
   U10502 : OR2_X1 port map( A1 => n25959, A2 => n287, Z => n484);
   U10510 : NAND2_X2 port map( A1 => n754, A2 => n5889, ZN => n19749);
   U10554 : OR2_X1 port map( A1 => n8554, A2 => n18921, Z => n23742);
   U10569 : XOR2_X1 port map( A1 => n20241, A2 => n22508, Z => n20252);
   U10571 : XOR2_X1 port map( A1 => n20233, A2 => n4137, Z => n22508);
   U10595 : AND2_X1 port map( A1 => n2068, A2 => n9330, Z => n24518);
   U10708 : NOR2_X1 port map( A1 => n13205, A2 => n24127, ZN => n17411);
   U10718 : XOR2_X1 port map( A1 => n12147, A2 => n22512, Z => n16807);
   U10722 : NAND2_X2 port map( A1 => n11546, A2 => n11548, ZN => n12147);
   U10731 : XOR2_X1 port map( A1 => n20531, A2 => n20764, Z => n7809);
   U10740 : OR2_X1 port map( A1 => n16585, A2 => n23907, Z => n7112);
   U10742 : NAND2_X2 port map( A1 => n22515, A2 => n19735, ZN => n19592);
   U10745 : NAND2_X1 port map( A1 => n21719, A2 => n21699, ZN => n22516);
   U10749 : NAND2_X2 port map( A1 => n800, A2 => n6371, ZN => n20797);
   U10767 : OAI21_X2 port map( A1 => n3255, A2 => n22563, B => n813, ZN => 
                           n8190);
   U10773 : INV_X4 port map( I => n14442, ZN => n8873);
   U10776 : AOI21_X1 port map( A1 => n14658, A2 => n9018, B => n3961, ZN => 
                           n3350);
   U10778 : INV_X1 port map( I => n3963, ZN => n3961);
   U10779 : XOR2_X1 port map( A1 => n12489, A2 => n578, Z => n3963);
   U10795 : NAND2_X2 port map( A1 => n5015, A2 => n22523, ZN => n17969);
   U10796 : AOI22_X1 port map( A1 => n6762, A2 => n17317, B1 => n11113, B2 => 
                           n17318, ZN => n22523);
   U10797 : XOR2_X1 port map( A1 => n22524, A2 => n18163, Z => n23720);
   U10824 : XOR2_X1 port map( A1 => n18014, A2 => n12135, Z => n22604);
   U10835 : XOR2_X1 port map( A1 => n6241, A2 => n18019, Z => n18197);
   U10840 : NOR2_X2 port map( A1 => n17201, A2 => n7982, ZN => n18019);
   U10842 : OAI21_X2 port map( A1 => n12840, A2 => n730, B => n13876, ZN => 
                           n3443);
   U10843 : OAI22_X2 port map( A1 => n21832, A2 => n22531, B1 => n23739, B2 => 
                           n17519, ZN => n10856);
   U10846 : XOR2_X1 port map( A1 => n11015, A2 => n10442, Z => n18612);
   U10856 : XOR2_X1 port map( A1 => n17013, A2 => n10535, Z => n16764);
   U10857 : NAND2_X2 port map( A1 => n9870, A2 => n9871, ZN => n10535);
   U10869 : NAND2_X2 port map( A1 => n14617, A2 => n14793, ZN => n16646);
   U10872 : XOR2_X1 port map( A1 => n12816, A2 => n25356, Z => n11898);
   U10885 : OAI21_X2 port map( A1 => n8006, A2 => n8007, B => n12698, ZN => 
                           n18804);
   U10891 : XOR2_X1 port map( A1 => n11038, A2 => n11037, Z => n22538);
   U10896 : XOR2_X1 port map( A1 => n26029, A2 => n20437, Z => n22540);
   U10901 : NAND2_X2 port map( A1 => n3764, A2 => n3762, ZN => n8554);
   U10902 : XOR2_X1 port map( A1 => n6702, A2 => n6744, Z => n22541);
   U10915 : NOR2_X2 port map( A1 => n8872, A2 => n250, ZN => n22936);
   U10936 : XOR2_X1 port map( A1 => n18079, A2 => n21909, Z => n24520);
   U10938 : XOR2_X1 port map( A1 => n18225, A2 => n11502, Z => n18079);
   U10954 : XOR2_X1 port map( A1 => n1199, A2 => n27145, Z => n18095);
   U10960 : XOR2_X1 port map( A1 => n22552, A2 => n9594, Z => n13580);
   U10963 : XOR2_X1 port map( A1 => n19506, A2 => n4175, Z => n22552);
   U10964 : INV_X2 port map( I => n22554, ZN => n1711);
   U10971 : AOI21_X2 port map( A1 => n15380, A2 => n14332, B => n15379, ZN => 
                           n22626);
   U10974 : XOR2_X1 port map( A1 => n24493, A2 => n12696, Z => n21054);
   U10985 : AND3_X1 port map( A1 => n5575, A2 => n20255, A3 => n22830, Z => 
                           n23621);
   U10993 : AND2_X1 port map( A1 => n23184, A2 => n6991, Z => n7074);
   U10999 : XOR2_X1 port map( A1 => n8671, A2 => n3355, Z => n12585);
   U11006 : NOR2_X2 port map( A1 => n17583, A2 => n14403, ZN => n14659);
   U11007 : XOR2_X1 port map( A1 => n280, A2 => n18236, Z => n18116);
   U11019 : NAND2_X2 port map( A1 => n14157, A2 => n3138, ZN => n22806);
   U11020 : NAND2_X1 port map( A1 => n22574, A2 => n5002, ZN => n5001);
   U11024 : AND2_X1 port map( A1 => n24579, A2 => n13194, Z => n14043);
   U11029 : XOR2_X1 port map( A1 => n22567, A2 => n15292, Z => n5605);
   U11030 : XOR2_X1 port map( A1 => n12691, A2 => n9497, Z => n22567);
   U11031 : OR2_X1 port map( A1 => n20280, A2 => n7749, Z => n7750);
   U11042 : INV_X2 port map( I => n22568, ZN => n22799);
   U11048 : XOR2_X1 port map( A1 => n1385, A2 => n22571, Z => n1381);
   U11049 : XOR2_X1 port map( A1 => n27399, A2 => n21937, Z => n22571);
   U11054 : XNOR2_X1 port map( A1 => n17039, A2 => n14640, ZN => n6573);
   U11065 : INV_X2 port map( I => n19447, ZN => n22577);
   U11076 : OAI21_X1 port map( A1 => n848, A2 => n4934, B => n22579, ZN => 
                           n20653);
   U11084 : OR2_X1 port map( A1 => n12203, A2 => n22581, Z => n22679);
   U11087 : AOI22_X2 port map( A1 => n8976, A2 => n11880, B1 => n20045, B2 => 
                           n28524, ZN => n22777);
   U11092 : OR2_X1 port map( A1 => n21275, A2 => n4143, Z => n14612);
   U11093 : INV_X2 port map( I => n6066, ZN => n749);
   U11095 : XOR2_X1 port map( A1 => n28464, A2 => n26469, Z => n4045);
   U11096 : AND2_X1 port map( A1 => n15526, A2 => n26665, Z => n16147);
   U11099 : XOR2_X1 port map( A1 => n18153, A2 => n18154, Z => n18341);
   U11130 : XNOR2_X1 port map( A1 => Plaintext(54), A2 => Key(54), ZN => n22590
                           );
   U11131 : XOR2_X1 port map( A1 => n22591, A2 => n4582, Z => n4950);
   U11136 : OR2_X1 port map( A1 => n17941, A2 => n10513, Z => n8917);
   U11138 : XOR2_X1 port map( A1 => n22592, A2 => n7222, Z => n23622);
   U11160 : NOR2_X1 port map( A1 => n10498, A2 => n10601, ZN => n10470);
   U11161 : XOR2_X1 port map( A1 => n10500, A2 => n10501, Z => n22978);
   U11165 : XOR2_X1 port map( A1 => n19536, A2 => n3243, Z => n19415);
   U11179 : XOR2_X1 port map( A1 => n19393, A2 => n19392, Z => n19427);
   U11180 : NOR2_X2 port map( A1 => n15207, A2 => n14239, ZN => n19393);
   U11181 : NAND2_X2 port map( A1 => n22600, A2 => n22599, ZN => n823);
   U11195 : OAI22_X2 port map( A1 => n18708, A2 => n27701, B1 => n14289, B2 => 
                           n14288, ZN => n19405);
   U11199 : INV_X2 port map( I => n4271, ZN => n5115);
   U11204 : XOR2_X1 port map( A1 => n12136, A2 => n22604, Z => n4271);
   U11213 : NAND2_X2 port map( A1 => n22605, A2 => n18478, ZN => n19306);
   U11214 : XOR2_X1 port map( A1 => n2071, A2 => n13078, Z => n7087);
   U11233 : XOR2_X1 port map( A1 => n22607, A2 => n14620, Z => Ciphertext(131))
                           ;
   U11240 : NOR2_X1 port map( A1 => n277, A2 => n25331, ZN => n22609);
   U11242 : XOR2_X1 port map( A1 => n20047, A2 => n386, Z => n385);
   U11243 : NOR2_X2 port map( A1 => n1988, A2 => n22612, ZN => n20044);
   U11255 : XOR2_X1 port map( A1 => n2476, A2 => n20539, Z => n22613);
   U11276 : OAI21_X2 port map( A1 => n12296, A2 => n9715, B => n7299, ZN => 
                           n9714);
   U11294 : XOR2_X1 port map( A1 => n10299, A2 => n22619, Z => n15138);
   U11296 : XOR2_X1 port map( A1 => n10352, A2 => n21237, Z => n22619);
   U11297 : INV_X2 port map( I => n21277, ZN => n21208);
   U11298 : XOR2_X1 port map( A1 => n14455, A2 => n21930, Z => n21277);
   U11313 : XOR2_X1 port map( A1 => n4970, A2 => n14345, Z => n18015);
   U11318 : XOR2_X1 port map( A1 => n22777, A2 => n22624, Z => n386);
   U11319 : INV_X1 port map( I => n20807, ZN => n22624);
   U11322 : NAND3_X1 port map( A1 => n13478, A2 => n9854, A3 => n7002, ZN => 
                           n7411);
   U11346 : AOI21_X2 port map( A1 => n762, A2 => n24175, B => n26681, ZN => 
                           n22630);
   U11352 : XOR2_X1 port map( A1 => n2614, A2 => n16965, Z => n22631);
   U11358 : XOR2_X1 port map( A1 => n18202, A2 => n18315, Z => n17709);
   U11359 : XOR2_X1 port map( A1 => n18062, A2 => n18021, Z => n18202);
   U11363 : NAND2_X1 port map( A1 => n22632, A2 => n1166, ZN => n5903);
   U11364 : AOI21_X1 port map( A1 => n6889, A2 => n22634, B => n22633, ZN => 
                           n22632);
   U11371 : NAND2_X2 port map( A1 => n24447, A2 => n23840, ZN => n23641);
   U11377 : NOR2_X2 port map( A1 => n3658, A2 => n3448, ZN => n21290);
   U11379 : NAND2_X1 port map( A1 => n935, A2 => n23753, ZN => n20795);
   U11395 : OAI21_X2 port map( A1 => n15416, A2 => n11453, B => n13467, ZN => 
                           n11197);
   U11407 : NAND2_X2 port map( A1 => n10058, A2 => n17847, ZN => n14788);
   U11408 : OAI21_X2 port map( A1 => n6410, A2 => n14665, B => n22641, ZN => 
                           n14352);
   U11409 : AOI22_X2 port map( A1 => n20864, A2 => n20865, B1 => n14666, B2 => 
                           n12887, ZN => n22641);
   U11413 : NAND2_X2 port map( A1 => n14803, A2 => n14801, ZN => n15256);
   U11414 : AND2_X1 port map( A1 => n11454, A2 => n19689, Z => n1804);
   U11416 : XOR2_X1 port map( A1 => n24048, A2 => n22642, Z => n14673);
   U11419 : XOR2_X1 port map( A1 => n8413, A2 => n8177, Z => n22642);
   U11423 : NAND2_X2 port map( A1 => n22645, A2 => n23945, ZN => n20312);
   U11425 : OAI21_X2 port map( A1 => n10140, A2 => n10139, B => n7238, ZN => 
                           n22645);
   U11427 : NAND2_X1 port map( A1 => n9041, A2 => n23538, ZN => n18736);
   U11435 : XOR2_X1 port map( A1 => n19187, A2 => n22647, Z => n4317);
   U11436 : NAND3_X1 port map( A1 => n15324, A2 => n15325, A3 => n21714, ZN => 
                           n24136);
   U11439 : XOR2_X1 port map( A1 => n11479, A2 => n11480, Z => n11491);
   U11447 : XOR2_X1 port map( A1 => n24094, A2 => n27360, Z => n21245);
   U11449 : NOR2_X2 port map( A1 => n15066, A2 => n15065, ZN => n24094);
   U11466 : OAI21_X1 port map( A1 => n5889, A2 => n19931, B => n27452, ZN => 
                           n19572);
   U11478 : XOR2_X1 port map( A1 => n27470, A2 => n19042, Z => n4425);
   U11486 : OAI21_X1 port map( A1 => n2703, A2 => n516, B => n4456, ZN => 
                           n16036);
   U11487 : NAND3_X2 port map( A1 => n19702, A2 => n27202, A3 => n3861, ZN => 
                           n14845);
   U11493 : NAND2_X1 port map( A1 => n22654, A2 => n28027, ZN => n22653);
   U11510 : NAND3_X2 port map( A1 => n10883, A2 => n10884, A3 => n21459, ZN => 
                           n11053);
   U11516 : INV_X2 port map( I => n22659, ZN => n18370);
   U11526 : NOR2_X1 port map( A1 => n21455, A2 => n23579, ZN => n13774);
   U11528 : AND2_X1 port map( A1 => n6821, A2 => n3525, Z => n6819);
   U11576 : NAND2_X2 port map( A1 => n9405, A2 => n22666, ZN => n9261);
   U11578 : AOI22_X1 port map( A1 => n15765, A2 => n14512, B1 => n15768, B2 => 
                           n15995, ZN => n22666);
   U11590 : AND2_X1 port map( A1 => n3729, A2 => n16640, Z => n3218);
   U11591 : XOR2_X1 port map( A1 => n12246, A2 => n20453, Z => n3748);
   U11594 : INV_X2 port map( I => n23454, ZN => n11198);
   U11615 : AOI21_X2 port map( A1 => n3929, A2 => n3234, B => n17594, ZN => 
                           n17595);
   U11621 : NAND2_X2 port map( A1 => n22671, A2 => n15231, ZN => n5616);
   U11626 : NAND2_X2 port map( A1 => n5069, A2 => n5068, ZN => n5082);
   U11630 : OR2_X1 port map( A1 => n18344, A2 => n4679, Z => n12703);
   U11635 : XOR2_X1 port map( A1 => n452, A2 => n22673, Z => n537);
   U11646 : XOR2_X1 port map( A1 => n22674, A2 => n13948, Z => n23582);
   U11651 : XOR2_X1 port map( A1 => n21364, A2 => n2655, Z => n11279);
   U11654 : OAI21_X2 port map( A1 => n14952, A2 => n5048, B => n14951, ZN => 
                           n21364);
   U11657 : NAND2_X2 port map( A1 => n15072, A2 => n22676, ZN => n16612);
   U11658 : OAI21_X2 port map( A1 => n16302, A2 => n9595, B => n14107, ZN => 
                           n22676);
   U11670 : OAI21_X2 port map( A1 => n10037, A2 => n16271, B => n22678, ZN => 
                           n10036);
   U11671 : NAND3_X2 port map( A1 => n16229, A2 => n16271, A3 => n10001, ZN => 
                           n22678);
   U11688 : INV_X2 port map( I => n8118, ZN => n7061);
   U11689 : OAI21_X2 port map( A1 => n23079, A2 => n4395, B => n4394, ZN => 
                           n8118);
   U11692 : XOR2_X1 port map( A1 => n22684, A2 => n21314, Z => n23248);
   U11702 : NAND2_X2 port map( A1 => n22898, A2 => n22687, ZN => n11871);
   U11742 : OAI21_X2 port map( A1 => n11503, A2 => n16433, B => n22296, ZN => 
                           n7429);
   U11785 : AND2_X1 port map( A1 => n25374, A2 => n10580, Z => n17168);
   U11799 : NAND2_X2 port map( A1 => n7783, A2 => n7780, ZN => n6098);
   U11804 : OAI21_X2 port map( A1 => n21670, A2 => n4623, B => n22695, ZN => 
                           n2777);
   U11809 : NOR2_X2 port map( A1 => n10454, A2 => n17748, ZN => n19154);
   U11814 : XOR2_X1 port map( A1 => n27104, A2 => n16910, Z => n22698);
   U11817 : AND2_X1 port map( A1 => n18794, A2 => n19056, Z => n23794);
   U11824 : XOR2_X1 port map( A1 => n7403, A2 => n22837, Z => n8992);
   U11826 : XOR2_X1 port map( A1 => n21150, A2 => n15455, Z => n3219);
   U11842 : XOR2_X1 port map( A1 => n22700, A2 => n22699, Z => n24418);
   U11845 : XOR2_X1 port map( A1 => n18046, A2 => n4457, Z => n22699);
   U11846 : XOR2_X1 port map( A1 => n18334, A2 => n1557, Z => n22700);
   U11858 : INV_X2 port map( I => n24558, ZN => n13278);
   U11869 : NOR2_X1 port map( A1 => n16598, A2 => n26008, ZN => n12879);
   U11875 : NAND2_X2 port map( A1 => n22704, A2 => n2862, ZN => n7298);
   U11884 : XOR2_X1 port map( A1 => n10787, A2 => n12222, Z => n3105);
   U11902 : AOI21_X2 port map( A1 => n15326, A2 => n15480, B => n18977, ZN => 
                           n4546);
   U11910 : XOR2_X1 port map( A1 => n5724, A2 => n22709, Z => n5721);
   U11911 : XOR2_X1 port map( A1 => n21303, A2 => n20335, Z => n22709);
   U11918 : XOR2_X1 port map( A1 => n23440, A2 => n22711, Z => n14392);
   U11934 : NOR2_X2 port map( A1 => n11597, A2 => n11598, ZN => n16918);
   U11935 : OAI22_X2 port map( A1 => n16421, A2 => n7115, B1 => n14008, B2 => 
                           n16587, ZN => n11597);
   U11942 : XOR2_X1 port map( A1 => n22716, A2 => n1298, Z => Ciphertext(165));
   U11945 : NOR2_X1 port map( A1 => n15218, A2 => n15217, ZN => n22716);
   U11951 : XOR2_X1 port map( A1 => n1918, A2 => n1916, Z => n5473);
   U11985 : OAI22_X2 port map( A1 => n2825, A2 => n14107, B1 => n2824, B2 => 
                           n516, ZN => n13739);
   U11995 : XOR2_X1 port map( A1 => n22719, A2 => n5524, Z => n5841);
   U12004 : XOR2_X1 port map( A1 => n20725, A2 => n20055, Z => n20062);
   U12018 : XOR2_X1 port map( A1 => n19093, A2 => n7592, Z => n23325);
   U12025 : OR2_X1 port map( A1 => n20087, A2 => n22000, Z => n12008);
   U12054 : XOR2_X1 port map( A1 => n6416, A2 => n22726, Z => n22725);
   U12072 : AND2_X1 port map( A1 => n4151, A2 => n4150, Z => n23);
   U12098 : INV_X4 port map( I => n21764, ZN => n838);
   U12116 : NAND2_X2 port map( A1 => n21324, A2 => n21277, ZN => n21327);
   U12131 : NAND2_X1 port map( A1 => n13219, A2 => n23784, ZN => n24112);
   U12146 : INV_X1 port map( I => n8237, ZN => n24022);
   U12147 : NAND2_X1 port map( A1 => n5781, A2 => n13432, ZN => n12063);
   U12170 : INV_X1 port map( I => n22728, ZN => n22729);
   U12172 : NAND2_X1 port map( A1 => n20308, A2 => n20156, ZN => n15542);
   U12174 : INV_X2 port map( I => n15103, ZN => n948);
   U12175 : OR2_X2 port map( A1 => n2183, A2 => n2181, Z => n22730);
   U12180 : NAND2_X1 port map( A1 => n910, A2 => n16493, ZN => n6147);
   U12190 : INV_X1 port map( I => n16826, ZN => n17059);
   U12191 : OR2_X1 port map( A1 => n4543, A2 => n4546, Z => n22795);
   U12197 : NOR3_X1 port map( A1 => n5853, A2 => n9986, A3 => n23104, ZN => 
                           n10090);
   U12207 : NAND2_X1 port map( A1 => n4190, A2 => n22776, ZN => n23808);
   U12226 : NOR2_X1 port map( A1 => n19106, A2 => n23546, ZN => n7551);
   U12230 : CLKBUF_X1 port map( I => n19273, Z => n22810);
   U12237 : INV_X2 port map( I => n7940, ZN => n14450);
   U12245 : OAI21_X1 port map( A1 => n1956, A2 => n20073, B => n23212, ZN => 
                           n1954);
   U12253 : INV_X1 port map( I => n10401, ZN => n9728);
   U12255 : NAND2_X1 port map( A1 => n15239, A2 => n3553, ZN => n9891);
   U12258 : NAND2_X1 port map( A1 => n9294, A2 => n23295, ZN => n8098);
   U12267 : OR2_X1 port map( A1 => n2254, A2 => n20658, Z => n4933);
   U12280 : NAND3_X1 port map( A1 => n10588, A2 => n20598, A3 => n20642, ZN => 
                           n20487);
   U12283 : NAND2_X1 port map( A1 => n5222, A2 => n17567, ZN => n12450);
   U12288 : NAND3_X1 port map( A1 => n885, A2 => n17822, A3 => n21898, ZN => 
                           n4611);
   U12292 : OAI21_X1 port map( A1 => n21898, A2 => n23110, B => n17931, ZN => 
                           n10849);
   U12293 : OAI21_X1 port map( A1 => n21898, A2 => n13329, B => n825, ZN => 
                           n17670);
   U12302 : INV_X1 port map( I => n10543, ZN => n16653);
   U12303 : OAI22_X1 port map( A1 => n12700, A2 => n1256, B1 => n4983, B2 => 
                           n10597, ZN => n16569);
   U12312 : NAND2_X1 port map( A1 => n11854, A2 => n10963, ZN => n10964);
   U12314 : INV_X1 port map( I => n20868, ZN => n22736);
   U12322 : INV_X2 port map( I => n15454, ZN => n21175);
   U12323 : NAND2_X1 port map( A1 => n2484, A2 => n19045, ZN => n15640);
   U12328 : AOI22_X1 port map( A1 => n9296, A2 => n865, B1 => n5008, B2 => 
                           n14356, ZN => n23295);
   U12330 : OR2_X1 port map( A1 => n14679, A2 => n15646, Z => n21552);
   U12340 : NAND2_X1 port map( A1 => n7405, A2 => n9990, ZN => n22739);
   U12341 : NAND2_X1 port map( A1 => n3530, A2 => n21387, ZN => n21129);
   U12342 : NOR2_X1 port map( A1 => n21638, A2 => n21641, ZN => n22740);
   U12357 : NAND2_X1 port map( A1 => n17560, A2 => n23269, ZN => n24386);
   U12369 : INV_X1 port map( I => n13248, ZN => n15733);
   U12375 : AOI21_X2 port map( A1 => n12962, A2 => n12960, B => n15530, ZN => 
                           n22741);
   U12381 : AOI21_X1 port map( A1 => n12962, A2 => n12960, B => n15530, ZN => 
                           n19550);
   U12386 : NOR2_X1 port map( A1 => n27386, A2 => n22762, ZN => n22743);
   U12399 : OR2_X2 port map( A1 => n3006, A2 => n12952, Z => n22744);
   U12400 : INV_X2 port map( I => n23871, ZN => n11576);
   U12411 : AOI21_X1 port map( A1 => n18795, A2 => n19057, B => n12781, ZN => 
                           n14020);
   U12413 : OR3_X1 port map( A1 => n22745, A2 => n13104, A3 => n25340, Z => 
                           n11668);
   U12417 : BUF_X2 port map( I => n13610, Z => n12465);
   U12422 : NOR2_X1 port map( A1 => n20802, A2 => n8990, ZN => n7147);
   U12424 : NAND2_X1 port map( A1 => n16730, A2 => n12117, ZN => n8518);
   U12445 : NOR2_X1 port map( A1 => n3060, A2 => n23146, ZN => n6782);
   U12453 : NAND2_X1 port map( A1 => n13146, A2 => n20209, ZN => n24230);
   U12454 : INV_X1 port map( I => n18084, ZN => n23581);
   U12485 : AND2_X1 port map( A1 => n2820, A2 => n9117, Z => n24201);
   U12490 : NOR2_X1 port map( A1 => n731, A2 => n7904, ZN => n8419);
   U12496 : AND2_X1 port map( A1 => n15458, A2 => n11622, Z => n11624);
   U12512 : AOI22_X1 port map( A1 => n11841, A2 => n11840, B1 => n19092, B2 => 
                           n19090, ZN => n22749);
   U12515 : NAND2_X1 port map( A1 => n11160, A2 => n13968, ZN => n24049);
   U12516 : INV_X1 port map( I => n11107, ZN => n22751);
   U12519 : INV_X2 port map( I => n11107, ZN => n936);
   U12526 : INV_X2 port map( I => n9140, ZN => n14437);
   U12544 : NAND2_X1 port map( A1 => n20392, A2 => n20309, ZN => n23914);
   U12549 : INV_X1 port map( I => n20757, ZN => n14628);
   U12566 : NAND2_X1 port map( A1 => n23023, A2 => n3326, ZN => n13981);
   U12602 : INV_X4 port map( I => n14858, ZN => n796);
   U12611 : OAI21_X1 port map( A1 => n22809, A2 => n27704, B => n12359, ZN => 
                           n18708);
   U12617 : AND2_X1 port map( A1 => n20177, A2 => n20176, Z => n22759);
   U12631 : NAND2_X2 port map( A1 => n5995, A2 => n5993, ZN => n22762);
   U12640 : NAND2_X1 port map( A1 => n7330, A2 => n10610, ZN => n1880);
   U12646 : NAND3_X1 port map( A1 => n14113, A2 => n7807, A3 => n7330, ZN => 
                           n8764);
   U12648 : OR3_X2 port map( A1 => n5462, A2 => n8510, A3 => n5461, Z => n22763
                           );
   U12650 : OR3_X2 port map( A1 => n5462, A2 => n8510, A3 => n5461, Z => n22764
                           );
   U12652 : NAND2_X2 port map( A1 => n16518, A2 => n24550, ZN => n16652);
   U12660 : OAI21_X1 port map( A1 => n1091, A2 => n27450, B => n948, ZN => 
                           n8876);
   U12677 : NAND2_X1 port map( A1 => n4899, A2 => n26308, ZN => n22765);
   U12682 : AND2_X2 port map( A1 => n2623, A2 => n2624, Z => n22766);
   U12697 : INV_X1 port map( I => n19085, ZN => n4080);
   U12698 : NAND2_X1 port map( A1 => n5815, A2 => n6052, ZN => n24072);
   U12715 : NAND2_X1 port map( A1 => n23401, A2 => n20213, ZN => n23180);
   U12716 : NAND3_X1 port map( A1 => n13422, A2 => n23120, A3 => n20213, ZN => 
                           n20005);
   U12731 : INV_X1 port map( I => n18070, ZN => n13164);
   U12740 : NAND2_X1 port map( A1 => n1573, A2 => n1572, ZN => n12366);
   U12743 : XOR2_X1 port map( A1 => n823, A2 => n18238, Z => n22773);
   U12751 : INV_X1 port map( I => n18359, ZN => n531);
   U12753 : NAND2_X1 port map( A1 => n20308, A2 => n26009, ZN => n20216);
   U12770 : NAND2_X1 port map( A1 => n19788, A2 => n19790, ZN => n15079);
   U12771 : NAND2_X1 port map( A1 => n1153, A2 => n11982, ZN => n23937);
   U12779 : NAND2_X1 port map( A1 => n28539, A2 => n26198, ZN => n23102);
   U12780 : NOR2_X1 port map( A1 => n18005, A2 => n9485, ZN => n12001);
   U12781 : INV_X1 port map( I => n18005, ZN => n22896);
   U12782 : OR2_X2 port map( A1 => n23018, A2 => n21761, Z => n22780);
   U12786 : INV_X1 port map( I => n664, ZN => n19935);
   U12789 : INV_X1 port map( I => n21303, ZN => n8372);
   U12793 : NAND2_X1 port map( A1 => n24616, A2 => n23602, ZN => n22781);
   U12799 : NAND2_X1 port map( A1 => n6211, A2 => n15478, ZN => n1948);
   U12801 : NAND2_X1 port map( A1 => n2252, A2 => n2251, ZN => n22784);
   U12802 : NAND2_X1 port map( A1 => n15118, A2 => n19673, ZN => n8358);
   U12804 : NAND3_X2 port map( A1 => n18871, A2 => n24442, A3 => n10618, ZN => 
                           n12661);
   U12807 : NAND2_X1 port map( A1 => n5664, A2 => n25455, ZN => n14566);
   U12827 : BUF_X2 port map( I => n19791, Z => n2320);
   U12828 : NAND2_X1 port map( A1 => n21020, A2 => n7228, ZN => n24468);
   U12831 : INV_X2 port map( I => n15639, ZN => n19443);
   U12837 : NAND2_X1 port map( A1 => n5748, A2 => n14683, ZN => n322);
   U12844 : INV_X1 port map( I => n2321, ZN => n2939);
   U12847 : NOR2_X1 port map( A1 => n2321, A2 => n20704, ZN => n20691);
   U12852 : NAND2_X1 port map( A1 => n10931, A2 => n27235, ZN => n24408);
   U12857 : AOI21_X1 port map( A1 => n20609, A2 => n22764, B => n25315, ZN => 
                           n20604);
   U12859 : INV_X2 port map( I => n22763, ZN => n8935);
   U12869 : NOR2_X1 port map( A1 => n18622, A2 => n1187, ZN => n5250);
   U12874 : OR2_X1 port map( A1 => n21638, A2 => n21641, Z => n21632);
   U12882 : NAND2_X1 port map( A1 => n18588, A2 => n10437, ZN => n2786);
   U12888 : NAND2_X1 port map( A1 => n22212, A2 => n22421, ZN => n23786);
   U12903 : NOR2_X1 port map( A1 => n961, A2 => n24998, ZN => n22983);
   U12909 : AND2_X1 port map( A1 => n11861, A2 => n12594, Z => n22790);
   U12910 : INV_X2 port map( I => n20658, ZN => n844);
   U12912 : NAND2_X1 port map( A1 => n3824, A2 => n20658, ZN => n20662);
   U12920 : AND2_X1 port map( A1 => n5573, A2 => n22830, Z => n1605);
   U12943 : NAND2_X1 port map( A1 => n13740, A2 => n17352, ZN => n17240);
   U12944 : NOR2_X1 port map( A1 => n20245, A2 => n26741, ZN => n20247);
   U12957 : NAND2_X1 port map( A1 => n860, A2 => n20291, ZN => n7734);
   U12959 : NAND2_X2 port map( A1 => n8928, A2 => n8927, ZN => n22792);
   U12970 : NAND2_X2 port map( A1 => n24437, A2 => n4515, ZN => n22794);
   U12971 : NAND2_X1 port map( A1 => n24437, A2 => n4515, ZN => n21394);
   U12972 : NAND2_X2 port map( A1 => n4514, A2 => n4512, ZN => n24437);
   U12987 : NOR2_X1 port map( A1 => n19918, A2 => n10593, ZN => n11314);
   U12988 : NOR2_X1 port map( A1 => n4198, A2 => n1015, ZN => n7277);
   U13001 : OAI21_X1 port map( A1 => n14628, A2 => n20899, B => n14627, ZN => 
                           n23512);
   U13002 : XNOR2_X1 port map( A1 => n10248, A2 => n15710, ZN => n2855);
   U13004 : NOR2_X1 port map( A1 => n3312, A2 => n24181, ZN => n656);
   U13008 : OAI21_X1 port map( A1 => n6264, A2 => n27454, B => n20188, ZN => 
                           n6282);
   U13014 : NAND2_X1 port map( A1 => n2960, A2 => n17301, ZN => n16999);
   U13015 : OAI21_X1 port map( A1 => n7055, A2 => n1629, B => n17301, ZN => 
                           n229);
   U13017 : INV_X1 port map( I => n6746, ZN => n24494);
   U13038 : NOR2_X1 port map( A1 => n21099, A2 => n12309, ZN => n13018);
   U13045 : NAND2_X2 port map( A1 => n17866, A2 => n17865, ZN => n22802);
   U13048 : AOI22_X1 port map( A1 => n3935, A2 => n3350, B1 => n3961, B2 => 
                           n3936, ZN => n3934);
   U13058 : NOR2_X1 port map( A1 => n772, A2 => n15513, ZN => n22864);
   U13062 : OAI22_X1 port map( A1 => n22782, A2 => n15279, B1 => n860, B2 => 
                           n20146, ZN => n12673);
   U13083 : NAND3_X1 port map( A1 => n10545, A2 => n23624, A3 => n18633, ZN => 
                           n18634);
   U13093 : XOR2_X1 port map( A1 => n20389, A2 => n3356, Z => n22811);
   U13096 : INV_X1 port map( I => n1191, ZN => n22869);
   U13099 : NOR2_X1 port map( A1 => n21538, A2 => n27389, ZN => n14229);
   U13102 : AND2_X2 port map( A1 => n2566, A2 => n2567, Z => n22812);
   U13108 : AND2_X2 port map( A1 => n16288, A2 => n13274, Z => n16182);
   U13117 : CLKBUF_X12 port map( I => Key(19), Z => n14590);
   U13122 : NAND3_X1 port map( A1 => n102, A2 => n21111, A3 => n4277, ZN => 
                           n13030);
   U13130 : NOR2_X1 port map( A1 => n22974, A2 => n27889, ZN => n3655);
   U13131 : NOR2_X1 port map( A1 => n10562, A2 => n11936, ZN => n22974);
   U13132 : NOR2_X1 port map( A1 => n22813, A2 => n11487, ZN => n1451);
   U13139 : XOR2_X1 port map( A1 => n7546, A2 => n7545, Z => n22814);
   U13149 : NAND3_X2 port map( A1 => n19702, A2 => n19836, A3 => n815, ZN => 
                           n19620);
   U13157 : NAND3_X1 port map( A1 => n18101, A2 => n25192, A3 => n100, ZN => 
                           n14984);
   U13161 : AND2_X2 port map( A1 => n3982, A2 => n9261, Z => n16661);
   U13168 : INV_X1 port map( I => n19478, ZN => n15684);
   U13173 : OAI22_X2 port map( A1 => n21831, A2 => n24067, B1 => n24066, B2 => 
                           n15481, ZN => n22818);
   U13176 : OAI22_X1 port map( A1 => n21831, A2 => n24067, B1 => n24066, B2 => 
                           n15481, ZN => n16857);
   U13181 : INV_X1 port map( I => n13351, ZN => n24108);
   U13183 : NAND2_X1 port map( A1 => n4662, A2 => n1048, ZN => n6564);
   U13198 : OAI21_X1 port map( A1 => n21501, A2 => n21499, B => n14450, ZN => 
                           n6081);
   U13200 : OAI21_X1 port map( A1 => n14450, A2 => n7941, B => n21499, ZN => 
                           n4516);
   U13201 : OAI21_X1 port map( A1 => n21500, A2 => n21499, B => n14450, ZN => 
                           n4513);
   U13214 : INV_X1 port map( I => n7168, ZN => n4780);
   U13222 : OR2_X1 port map( A1 => n21487, A2 => n11622, Z => n21474);
   U13224 : XOR2_X1 port map( A1 => n1888, A2 => n3985, Z => n22825);
   U13230 : XOR2_X1 port map( A1 => n5560, A2 => n1359, Z => n22826);
   U13237 : INV_X2 port map( I => n14291, ZN => n18627);
   U13245 : NOR3_X1 port map( A1 => n13255, A2 => n2185, A3 => n4274, ZN => 
                           n3885);
   U13261 : INV_X2 port map( I => n23916, ZN => n808);
   U13263 : NOR2_X1 port map( A1 => n23916, A2 => n20273, ZN => n12826);
   U13273 : NAND2_X1 port map( A1 => n23916, A2 => n20273, ZN => n24407);
   U13282 : OAI22_X1 port map( A1 => n1046, A2 => n5310, B1 => n4644, B2 => 
                           n5874, ZN => n4662);
   U13292 : NAND3_X2 port map( A1 => n12164, A2 => n12561, A3 => n3207, ZN => 
                           n22829);
   U13296 : OAI21_X1 port map( A1 => n15894, A2 => n16209, B => n16339, ZN => 
                           n23879);
   U13309 : NAND2_X1 port map( A1 => n8487, A2 => n12218, ZN => n23169);
   U13311 : AOI21_X1 port map( A1 => n12218, A2 => n19883, B => n2049, ZN => 
                           n4241);
   U13319 : INV_X1 port map( I => n9772, ZN => n17880);
   U13324 : NOR3_X1 port map( A1 => n26960, A2 => n26741, A3 => n22779, ZN => 
                           n15164);
   U13325 : AND3_X1 port map( A1 => n5395, A2 => n12335, A3 => n5394, Z => 
                           n22831);
   U13333 : NAND2_X1 port map( A1 => n21174, A2 => n21166, ZN => n3642);
   U13339 : OAI21_X1 port map( A1 => n12226, A2 => n12227, B => n12209, ZN => 
                           n1834);
   U13355 : AOI21_X2 port map( A1 => n4800, A2 => n4799, B => n23188, ZN => 
                           n22834);
   U13372 : XOR2_X1 port map( A1 => n18132, A2 => n18081, Z => n22836);
   U13377 : INV_X1 port map( I => n12675, ZN => n1067);
   U13378 : NAND2_X2 port map( A1 => n10965, A2 => n12255, ZN => n22837);
   U13383 : OAI21_X1 port map( A1 => n3204, A2 => n3205, B => n22762, ZN => 
                           n23455);
   U13387 : NAND2_X1 port map( A1 => n21621, A2 => n20365, ZN => n11286);
   U13390 : OAI22_X2 port map( A1 => n23259, A2 => n24008, B1 => n14071, B2 => 
                           n796, ZN => n22838);
   U13406 : NOR2_X1 port map( A1 => n1156, A2 => n27465, ZN => n8313);
   U13415 : XOR2_X1 port map( A1 => n5065, A2 => n5063, Z => n22842);
   U13423 : NOR2_X1 port map( A1 => n18799, A2 => n7018, ZN => n11554);
   U13424 : NOR2_X1 port map( A1 => n14437, A2 => n9047, ZN => n15553);
   U13425 : INV_X1 port map( I => n8673, ZN => n8997);
   U13426 : INV_X2 port map( I => n2359, ZN => n21685);
   U13427 : NAND3_X1 port map( A1 => n2778, A2 => n25314, A3 => n2359, ZN => 
                           n21676);
   U13431 : NAND2_X1 port map( A1 => n3960, A2 => n8290, ZN => n1497);
   U13432 : XOR2_X1 port map( A1 => n26496, A2 => n22123, Z => n22846);
   U13433 : INV_X1 port map( I => n9422, ZN => n21030);
   U13437 : OAI21_X1 port map( A1 => n1519, A2 => n3470, B => n14478, ZN => 
                           n9668);
   U13444 : INV_X1 port map( I => n19968, ZN => n20278);
   U13448 : NOR2_X1 port map( A1 => n13009, A2 => n11522, ZN => n11751);
   U13456 : NOR2_X1 port map( A1 => n20188, A2 => n8100, ZN => n190);
   U13457 : OAI21_X1 port map( A1 => n20188, A2 => n27454, B => n8100, ZN => 
                           n12723);
   U13478 : XOR2_X1 port map( A1 => n17117, A2 => n11671, Z => n16874);
   U13480 : OAI21_X2 port map( A1 => n1858, A2 => n2789, B => n1854, ZN => 
                           n11671);
   U13485 : OR2_X1 port map( A1 => n22825, A2 => n10971, Z => n9150);
   U13487 : NAND2_X1 port map( A1 => n17891, A2 => n18498, ZN => n18570);
   U13492 : INV_X1 port map( I => n23359, ZN => n23142);
   U13512 : INV_X2 port map( I => n10638, ZN => n22856);
   U13516 : AOI21_X2 port map( A1 => n16140, A2 => n14520, B => n7525, ZN => 
                           n23259);
   U13522 : NAND2_X2 port map( A1 => n9459, A2 => n17457, ZN => n2835);
   U13527 : XOR2_X1 port map( A1 => n6295, A2 => n15576, Z => n17457);
   U13538 : NAND2_X2 port map( A1 => n4899, A2 => n26308, ZN => n4898);
   U13542 : AOI22_X2 port map( A1 => n16503, A2 => n913, B1 => n11894, B2 => 
                           n11503, ZN => n11343);
   U13553 : OAI21_X2 port map( A1 => n22864, A2 => n22863, B => n21713, ZN => 
                           n5995);
   U13557 : OAI21_X1 port map( A1 => n23793, A2 => n23794, B => n12571, ZN => 
                           n4675);
   U13563 : INV_X2 port map( I => n5391, ZN => n22865);
   U13567 : XOR2_X1 port map( A1 => n22741, A2 => n22866, Z => n19248);
   U13570 : XOR2_X1 port map( A1 => n22868, A2 => n9145, Z => n24525);
   U13574 : XOR2_X1 port map( A1 => n9144, A2 => n23581, Z => n22868);
   U13579 : NAND3_X1 port map( A1 => n27386, A2 => n6182, A3 => n22762, ZN => 
                           n1634);
   U13599 : NAND2_X2 port map( A1 => n13601, A2 => n24423, ZN => n11224);
   U13601 : XNOR2_X1 port map( A1 => n2681, A2 => n2679, ZN => n10536);
   U13620 : OR2_X1 port map( A1 => n10220, A2 => n542, Z => n17386);
   U13625 : XOR2_X1 port map( A1 => n27444, A2 => n19430, Z => n19542);
   U13632 : OAI21_X2 port map( A1 => n22876, A2 => n24215, B => n24341, ZN => 
                           n2061);
   U13633 : XOR2_X1 port map( A1 => n22877, A2 => n8568, Z => n17336);
   U13640 : OAI21_X2 port map( A1 => n22881, A2 => n8060, B => n22880, ZN => 
                           n20964);
   U13654 : OAI21_X2 port map( A1 => n18404, A2 => n13455, B => n11478, ZN => 
                           n23060);
   U13655 : XOR2_X1 port map( A1 => Plaintext(72), A2 => Key(72), Z => n24311);
   U13670 : XNOR2_X1 port map( A1 => n19305, A2 => n19261, ZN => n19240);
   U13673 : AOI22_X2 port map( A1 => n18919, A2 => n6708, B1 => n1415, B2 => 
                           n11577, ZN => n22887);
   U13678 : INV_X2 port map( I => n22889, ZN => n13467);
   U13680 : INV_X1 port map( I => n20741, ZN => n22890);
   U13684 : NAND2_X2 port map( A1 => n13224, A2 => n3112, ZN => n15639);
   U13688 : NOR2_X2 port map( A1 => n24603, A2 => n1720, ZN => n22893);
   U13699 : NOR2_X2 port map( A1 => n24091, A2 => n24090, ZN => n5204);
   U13703 : XOR2_X1 port map( A1 => n3925, A2 => n22926, Z => n24098);
   U13731 : XOR2_X1 port map( A1 => n19214, A2 => n22795, Z => n19255);
   U13734 : NAND2_X2 port map( A1 => n22900, A2 => n3934, ZN => n11391);
   U13735 : NAND2_X1 port map( A1 => n3118, A2 => n14658, ZN => n22900);
   U13741 : NAND2_X1 port map( A1 => n10620, A2 => n13385, ZN => n17254);
   U13742 : NAND2_X2 port map( A1 => n19635, A2 => n21813, ZN => n2553);
   U13744 : NAND2_X2 port map( A1 => n22902, A2 => n13498, ZN => n23418);
   U13745 : NAND2_X2 port map( A1 => n2285, A2 => n2238, ZN => n22902);
   U13751 : XOR2_X1 port map( A1 => n4020, A2 => n19281, Z => n4019);
   U13753 : NOR2_X2 port map( A1 => n20319, A2 => n20318, ZN => n12812);
   U13760 : INV_X1 port map( I => n22751, ZN => n23919);
   U13762 : XOR2_X1 port map( A1 => n19220, A2 => n19435, Z => n19359);
   U13784 : OR2_X1 port map( A1 => n19490, A2 => n12209, Z => n22913);
   U13785 : NAND2_X2 port map( A1 => n13617, A2 => n22914, ZN => n15502);
   U13795 : AOI22_X1 port map( A1 => n18580, A2 => n13612, B1 => n10537, B2 => 
                           n23062, ZN => n22914);
   U13796 : NAND3_X1 port map( A1 => n21896, A2 => n16639, A3 => n16640, ZN => 
                           n23840);
   U13830 : XOR2_X1 port map( A1 => n16932, A2 => n16931, Z => n6295);
   U13840 : XOR2_X1 port map( A1 => n16944, A2 => n26449, Z => n23659);
   U13852 : AND2_X1 port map( A1 => n3850, A2 => n16203, Z => n10575);
   U13853 : INV_X2 port map( I => n22927, ZN => n17230);
   U13858 : OAI21_X2 port map( A1 => n716, A2 => n17867, B => n14167, ZN => 
                           n17772);
   U13860 : NAND2_X2 port map( A1 => n19585, A2 => n10698, ZN => n20065);
   U13868 : XOR2_X1 port map( A1 => n21418, A2 => n21420, Z => n22931);
   U13875 : NOR2_X1 port map( A1 => n15986, A2 => n15987, ZN => n22932);
   U13891 : INV_X2 port map( I => n18314, ZN => n22938);
   U13910 : XOR2_X1 port map( A1 => n22944, A2 => n14638, Z => Ciphertext(104))
                           ;
   U13946 : XOR2_X1 port map( A1 => n22946, A2 => n5734, Z => Ciphertext(49));
   U13969 : XOR2_X1 port map( A1 => n11555, A2 => n18142, Z => n18191);
   U13971 : NAND3_X2 port map( A1 => n9152, A2 => n7232, A3 => n19022, ZN => 
                           n19451);
   U13978 : NOR2_X1 port map( A1 => n23650, A2 => n15705, ZN => n8832);
   U13980 : XOR2_X1 port map( A1 => Plaintext(181), A2 => Key(181), Z => n576);
   U13985 : XOR2_X1 port map( A1 => n20092, A2 => n5949, Z => n2889);
   U14009 : NAND2_X1 port map( A1 => n23042, A2 => n7358, ZN => n22956);
   U14028 : AOI21_X2 port map( A1 => n16078, A2 => n10427, B => n10036, ZN => 
                           n23128);
   U14030 : NAND2_X2 port map( A1 => n12062, A2 => n12064, ZN => n12061);
   U14044 : XOR2_X1 port map( A1 => n3510, A2 => n22960, Z => n10301);
   U14053 : AOI21_X2 port map( A1 => n4788, A2 => n14579, B => n16484, ZN => 
                           n14122);
   U14054 : NOR2_X2 port map( A1 => n7517, A2 => n16525, ZN => n4788);
   U14056 : AND2_X2 port map( A1 => n1902, A2 => n23486, Z => n23023);
   U14060 : XOR2_X1 port map( A1 => n20546, A2 => n20498, Z => n3996);
   U14062 : XOR2_X1 port map( A1 => n20480, A2 => n4501, Z => n20498);
   U14067 : NAND2_X2 port map( A1 => n24430, A2 => n7458, ZN => n20336);
   U14070 : AOI22_X1 port map( A1 => n17279, A2 => n13421, B1 => n17278, B2 => 
                           n14278, ZN => n22962);
   U14089 : NOR3_X2 port map( A1 => n7457, A2 => n5910, A3 => n7618, ZN => 
                           n22965);
   U14091 : NOR2_X1 port map( A1 => n21110, A2 => n11522, ZN => n11521);
   U14094 : OR2_X1 port map( A1 => n12726, A2 => n16707, Z => n16709);
   U14105 : NOR2_X1 port map( A1 => n27492, A2 => n19163, ZN => n22967);
   U14138 : INV_X1 port map( I => n22974, ZN => n10346);
   U14161 : XOR2_X1 port map( A1 => n15487, A2 => n4398, Z => n1370);
   U14169 : XOR2_X1 port map( A1 => n12204, A2 => n21419, Z => n11193);
   U14184 : AOI21_X1 port map( A1 => n27630, A2 => n961, B => n22983, ZN => 
                           n6449);
   U14190 : AOI21_X2 port map( A1 => n23864, A2 => n12444, B => n19623, ZN => 
                           n9878);
   U14195 : XOR2_X1 port map( A1 => n12626, A2 => n14544, Z => n7221);
   U14207 : XOR2_X1 port map( A1 => n18276, A2 => n22988, Z => n3351);
   U14225 : XOR2_X1 port map( A1 => n7861, A2 => n3615, Z => n3614);
   U14252 : XOR2_X1 port map( A1 => n22994, A2 => n20433, Z => Ciphertext(168))
                           ;
   U14253 : NAND2_X1 port map( A1 => n1635, A2 => n1633, ZN => n22994);
   U14255 : OAI21_X2 port map( A1 => n974, A2 => n19830, B => n22995, ZN => 
                           n19946);
   U14265 : XOR2_X1 port map( A1 => n16765, A2 => n14797, Z => n14796);
   U14270 : NAND2_X2 port map( A1 => n22996, A2 => n23722, ZN => n24181);
   U14272 : XOR2_X1 port map( A1 => n16959, A2 => n21602, Z => n3411);
   U14282 : INV_X1 port map( I => n12625, ZN => n21524);
   U14294 : XOR2_X1 port map( A1 => n6024, A2 => n14, Z => n18133);
   U14296 : XOR2_X1 port map( A1 => n11233, A2 => n8339, Z => n8338);
   U14308 : INV_X4 port map( I => n23002, ZN => n13389);
   U14311 : OR2_X1 port map( A1 => n20852, A2 => n20982, Z => n15005);
   U14312 : INV_X2 port map( I => n1381, ZN => n15513);
   U14321 : NAND2_X1 port map( A1 => n3984, A2 => n10289, ZN => n23005);
   U14324 : XOR2_X1 port map( A1 => n20762, A2 => n21928, Z => n23007);
   U14333 : XOR2_X1 port map( A1 => n16992, A2 => n16786, Z => n4272);
   U14339 : INV_X2 port map( I => n4814, ZN => n23011);
   U14344 : XOR2_X1 port map( A1 => n26576, A2 => n20908, Z => n16616);
   U14346 : XOR2_X1 port map( A1 => n23013, A2 => n14015, Z => n14132);
   U14349 : XOR2_X1 port map( A1 => n17086, A2 => n14014, Z => n23013);
   U14371 : XOR2_X1 port map( A1 => n20252, A2 => n23014, Z => n21092);
   U14375 : OR2_X1 port map( A1 => n18426, A2 => n19148, Z => n18434);
   U14399 : OR2_X1 port map( A1 => n841, A2 => n9557, Z => n23910);
   U14403 : INV_X1 port map( I => n23064, ZN => n12951);
   U14411 : NAND2_X2 port map( A1 => n13232, A2 => n7082, ZN => n23064);
   U14417 : NAND2_X1 port map( A1 => n899, A2 => n16406, ZN => n23019);
   U14421 : XOR2_X1 port map( A1 => n8601, A2 => n8600, Z => n3005);
   U14423 : OR2_X1 port map( A1 => n22840, A2 => n10209, Z => n6654);
   U14424 : XOR2_X1 port map( A1 => n698, A2 => n2604, Z => n23022);
   U14426 : NAND3_X1 port map( A1 => n15348, A2 => n2102, A3 => n977, ZN => 
                           n11150);
   U14441 : XOR2_X1 port map( A1 => n6108, A2 => n21784, Z => n7106);
   U14442 : XOR2_X1 port map( A1 => n12351, A2 => n19371, Z => n23026);
   U14465 : XOR2_X1 port map( A1 => n2176, A2 => n2174, Z => n3490);
   U14471 : OR2_X1 port map( A1 => n23907, A2 => n25693, Z => n16588);
   U14481 : AND3_X1 port map( A1 => n22776, A2 => n22398, A3 => n9525, Z => 
                           n23205);
   U14505 : NOR2_X2 port map( A1 => n9322, A2 => n18956, ZN => n12357);
   U14510 : NAND2_X2 port map( A1 => n13563, A2 => n25099, ZN => n9322);
   U14534 : XOR2_X1 port map( A1 => n5937, A2 => n1134, Z => n23047);
   U14547 : NAND2_X1 port map( A1 => n9003, A2 => n9005, ZN => n23054);
   U14565 : XOR2_X1 port map( A1 => n4633, A2 => n2376, Z => n2375);
   U14566 : XOR2_X1 port map( A1 => n18212, A2 => n21893, Z => n5989);
   U14568 : XOR2_X1 port map( A1 => n16773, A2 => n23103, Z => n14533);
   U14586 : NAND2_X2 port map( A1 => n23066, A2 => n14353, ZN => n17867);
   U14588 : OAI21_X1 port map( A1 => n2137, A2 => n21161, B => n10031, ZN => 
                           n23067);
   U14596 : NAND3_X2 port map( A1 => n23071, A2 => n13581, A3 => n9337, ZN => 
                           n13855);
   U14598 : AND2_X1 port map( A1 => n26491, A2 => n23072, Z => n9108);
   U14602 : XOR2_X1 port map( A1 => n18036, A2 => n18262, Z => n23074);
   U14610 : XOR2_X1 port map( A1 => n9104, A2 => n8310, Z => n5432);
   U14637 : XNOR2_X1 port map( A1 => n8132, A2 => n21649, ZN => n23764);
   U14646 : XNOR2_X1 port map( A1 => n23127, A2 => n2020, ZN => n23081);
   U14654 : INV_X1 port map( I => n6205, ZN => n23652);
   U14660 : XOR2_X1 port map( A1 => n19239, A2 => n19240, Z => n23086);
   U14678 : OAI21_X1 port map( A1 => n12046, A2 => n12045, B => n2514, ZN => 
                           n1825);
   U14688 : INV_X2 port map( I => n23094, ZN => n9986);
   U14690 : XOR2_X1 port map( A1 => Plaintext(178), A2 => Key(178), Z => n23094
                           );
   U14691 : INV_X1 port map( I => n10093, ZN => n23165);
   U14702 : NAND2_X1 port map( A1 => n242, A2 => n17576, ZN => n17503);
   U14703 : INV_X2 port map( I => n1964, ZN => n14501);
   U14710 : XOR2_X1 port map( A1 => n1649, A2 => n1648, Z => n1964);
   U14711 : NAND2_X2 port map( A1 => n23097, A2 => n7548, ZN => n8399);
   U14712 : NOR2_X2 port map( A1 => n1783, A2 => n1785, ZN => n19140);
   U14721 : XOR2_X1 port map( A1 => n16770, A2 => n16771, Z => n23103);
   U14726 : INV_X2 port map( I => n624, ZN => n23105);
   U14744 : AND2_X1 port map( A1 => n19107, A2 => n14836, Z => n3670);
   U14746 : INV_X2 port map( I => n23109, ZN => n1458);
   U14747 : NAND2_X2 port map( A1 => n11664, A2 => n18102, ZN => n23186);
   U14765 : XOR2_X1 port map( A1 => n23111, A2 => n9063, Z => n13712);
   U14767 : INV_X2 port map( I => n19393, ZN => n23111);
   U14777 : NAND2_X2 port map( A1 => n15514, A2 => n10046, ZN => n2037);
   U14778 : XOR2_X1 port map( A1 => n23116, A2 => n3404, Z => n6549);
   U14793 : AOI21_X2 port map( A1 => n12790, A2 => n26243, B => n12789, ZN => 
                           n2437);
   U14800 : NAND2_X2 port map( A1 => n8320, A2 => n6581, ZN => n8322);
   U14802 : XOR2_X1 port map( A1 => n3134, A2 => n9148, Z => n9147);
   U14820 : XOR2_X1 port map( A1 => n2019, A2 => n2018, Z => n23127);
   U14831 : XOR2_X1 port map( A1 => n13458, A2 => n6154, Z => n1518);
   U14854 : XOR2_X1 port map( A1 => n23139, A2 => n15017, Z => n15386);
   U14856 : XOR2_X1 port map( A1 => n15016, A2 => n15015, Z => n23139);
   U14863 : XOR2_X1 port map( A1 => n23142, A2 => n602, Z => n1888);
   U14871 : NOR2_X1 port map( A1 => n16196, A2 => n15917, ZN => n2283);
   U14892 : XOR2_X1 port map( A1 => n19387, A2 => n19302, Z => n3022);
   U14893 : NAND2_X2 port map( A1 => n905, A2 => n12726, ZN => n16576);
   U14922 : OAI22_X2 port map( A1 => n23158, A2 => n23157, B1 => n2062, B2 => 
                           n12310, ZN => n11107);
   U14924 : NAND2_X2 port map( A1 => n9286, A2 => n23160, ZN => n9285);
   U14959 : XOR2_X1 port map( A1 => n792, A2 => n23168, Z => n303);
   U14969 : OR2_X1 port map( A1 => n15282, A2 => n14843, Z => n1931);
   U14970 : XOR2_X1 port map( A1 => n12099, A2 => n14405, Z => n20356);
   U14972 : NAND2_X2 port map( A1 => n10967, A2 => n12239, ZN => n12099);
   U14976 : AOI21_X2 port map( A1 => n24620, A2 => n23171, B => n23170, ZN => 
                           n7622);
   U15003 : NAND3_X2 port map( A1 => n23175, A2 => n19105, A3 => n2356, ZN => 
                           n14833);
   U15023 : INV_X2 port map( I => n23178, ZN => n574);
   U15024 : XNOR2_X1 port map( A1 => Plaintext(9), A2 => Key(9), ZN => n23178);
   U15030 : NAND4_X2 port map( A1 => n23181, A2 => n20003, A3 => n20005, A4 => 
                           n23180, ZN => n15119);
   U15039 : XOR2_X1 port map( A1 => n11074, A2 => n18030, Z => n1648);
   U15044 : NAND2_X2 port map( A1 => n1587, A2 => n9356, ZN => n11074);
   U15058 : NAND2_X2 port map( A1 => n2853, A2 => n2852, ZN => n2850);
   U15069 : INV_X2 port map( I => n23185, ZN => n12256);
   U15070 : XNOR2_X1 port map( A1 => n9044, A2 => n23717, ZN => n23185);
   U15071 : AOI21_X2 port map( A1 => n4749, A2 => n24330, B => n17848, ZN => 
                           n23187);
   U15082 : OAI22_X2 port map( A1 => n17538, A2 => n1035, B1 => n4798, B2 => 
                           n4797, ZN => n23188);
   U15086 : XOR2_X1 port map( A1 => n24582, A2 => n12249, Z => n3779);
   U15091 : AOI21_X1 port map( A1 => n12433, A2 => n12432, B => n28527, ZN => 
                           n12030);
   U15094 : NOR2_X1 port map( A1 => n13391, A2 => n16457, ZN => n16458);
   U15095 : OAI21_X2 port map( A1 => n19062, A2 => n23643, B => n19061, ZN => 
                           n23191);
   U15106 : XOR2_X1 port map( A1 => n17672, A2 => n24116, Z => n18725);
   U15125 : INV_X1 port map( I => n27390, ZN => n843);
   U15131 : NAND2_X2 port map( A1 => n1520, A2 => n9390, ZN => n11048);
   U15132 : NAND2_X2 port map( A1 => n15507, A2 => n15969, ZN => n16630);
   U15137 : NAND2_X1 port map( A1 => n24628, A2 => n4532, ZN => n23992);
   U15140 : NOR2_X1 port map( A1 => n1113, A2 => n22295, ZN => n4190);
   U15153 : INV_X2 port map( I => n23202, ZN => n9670);
   U15154 : INV_X2 port map( I => n23203, ZN => n18442);
   U15166 : XOR2_X1 port map( A1 => n23211, A2 => n1295, Z => Ciphertext(3));
   U15169 : OAI21_X2 port map( A1 => n17234, A2 => n894, B => n27788, ZN => 
                           n17235);
   U15170 : NAND2_X2 port map( A1 => n23322, A2 => n866, ZN => n19669);
   U15177 : NAND2_X2 port map( A1 => n23220, A2 => n23219, ZN => n16497);
   U15180 : INV_X1 port map( I => n16183, ZN => n23221);
   U15222 : NAND2_X2 port map( A1 => n4416, A2 => n3034, ZN => n4414);
   U15226 : XOR2_X1 port map( A1 => n12209, A2 => n25372, Z => n3733);
   U15233 : NOR2_X1 port map( A1 => n23227, A2 => n17188, ZN => n10694);
   U15237 : XOR2_X1 port map( A1 => n21240, A2 => n23228, Z => n23834);
   U15240 : XOR2_X1 port map( A1 => n21149, A2 => n23426, Z => n23228);
   U15250 : XOR2_X1 port map( A1 => n2016, A2 => n15149, Z => n4889);
   U15263 : NAND2_X1 port map( A1 => n1863, A2 => n1864, ZN => n23232);
   U15279 : INV_X1 port map( I => n26076, ZN => n827);
   U15282 : OR2_X1 port map( A1 => n26076, A2 => n6098, Z => n17798);
   U15285 : OR2_X1 port map( A1 => n24316, A2 => n23072, Z => n24462);
   U15288 : NAND2_X1 port map( A1 => n24120, A2 => n14917, ZN => n6608);
   U15299 : NOR2_X1 port map( A1 => n2818, A2 => n22237, ZN => n2817);
   U15304 : XOR2_X1 port map( A1 => n6746, A2 => n16893, Z => n23238);
   U15307 : OAI21_X2 port map( A1 => n10693, A2 => n13229, B => n23597, ZN => 
                           n23239);
   U15320 : XOR2_X1 port map( A1 => n14601, A2 => n14610, Z => n20233);
   U15344 : OAI22_X1 port map( A1 => n16611, A2 => n16493, B1 => n1243, B2 => 
                           n25698, ZN => n23244);
   U15366 : XOR2_X1 port map( A1 => n16987, A2 => n16805, Z => n7712);
   U15376 : NAND2_X2 port map( A1 => n26635, A2 => n27227, ZN => n14448);
   U15387 : NAND2_X2 port map( A1 => n14447, A2 => n2347, ZN => n20480);
   U15388 : INV_X1 port map( I => n6842, ZN => n15971);
   U15391 : NAND2_X1 port map( A1 => n15806, A2 => n14515, ZN => n6842);
   U15396 : AND2_X1 port map( A1 => n19873, A2 => n19870, Z => n13226);
   U15397 : INV_X2 port map( I => n23258, ZN => n21456);
   U15410 : NOR2_X1 port map( A1 => n11816, A2 => n13184, ZN => n10962);
   U15428 : OAI21_X1 port map( A1 => n10276, A2 => n22766, B => n10275, ZN => 
                           n23260);
   U15430 : NOR3_X2 port map( A1 => n26363, A2 => n24406, A3 => n17547, ZN => 
                           n13062);
   U15450 : NAND2_X2 port map( A1 => n12570, A2 => n19793, ZN => n23817);
   U15452 : NAND2_X2 port map( A1 => n15079, A2 => n12443, ZN => n12570);
   U15453 : XOR2_X1 port map( A1 => n9002, A2 => n19453, Z => n19537);
   U15476 : XOR2_X1 port map( A1 => n3506, A2 => n20543, Z => n20497);
   U15491 : XOR2_X1 port map( A1 => n12102, A2 => n15719, Z => n8601);
   U15494 : NAND2_X2 port map( A1 => n12619, A2 => n12618, ZN => n18137);
   U15497 : INV_X2 port map( I => n3003, ZN => n18633);
   U15519 : INV_X2 port map( I => n23284, ZN => n8468);
   U15526 : INV_X2 port map( I => n15997, ZN => n12116);
   U15531 : XOR2_X1 port map( A1 => n2959, A2 => Key(51), Z => n15997);
   U15544 : XOR2_X1 port map( A1 => n3580, A2 => n23285, Z => n3579);
   U15547 : XOR2_X1 port map( A1 => n17876, A2 => n21821, Z => n23285);
   U15554 : XOR2_X1 port map( A1 => n5594, A2 => n5590, Z => n14759);
   U15560 : XOR2_X1 port map( A1 => n18034, A2 => n14781, Z => n14780);
   U15561 : XOR2_X1 port map( A1 => n18061, A2 => n5413, Z => n18034);
   U15574 : NAND2_X1 port map( A1 => n19580, A2 => n19843, ZN => n23445);
   U15578 : XOR2_X1 port map( A1 => n9544, A2 => n19264, Z => n5937);
   U15579 : XOR2_X1 port map( A1 => n8343, A2 => n8341, Z => n20783);
   U15580 : XNOR2_X1 port map( A1 => n19383, A2 => n550, ZN => n23312);
   U15589 : XOR2_X1 port map( A1 => n17127, A2 => n6137, Z => n23294);
   U15597 : AOI22_X1 port map( A1 => n21537, A2 => n21525, B1 => n21519, B2 => 
                           n21520, ZN => n7145);
   U15599 : NAND2_X2 port map( A1 => n23301, A2 => n308, ZN => n17015);
   U15627 : INV_X2 port map( I => n23304, ZN => n14178);
   U15628 : XOR2_X1 port map( A1 => Key(74), A2 => Plaintext(74), Z => n23304);
   U15630 : XOR2_X1 port map( A1 => n16763, A2 => n11041, Z => n11040);
   U15646 : XOR2_X1 port map( A1 => n4658, A2 => n12281, Z => n23307);
   U15685 : OAI21_X2 port map( A1 => n7774, A2 => n23315, B => n17448, ZN => 
                           n7156);
   U15689 : OAI22_X1 port map( A1 => n1224, A2 => n21785, B1 => n17548, B2 => 
                           n10546, ZN => n23315);
   U15695 : INV_X4 port map( I => n23318, ZN => n7180);
   U15704 : NOR2_X2 port map( A1 => n13704, A2 => n15309, ZN => n23318);
   U15710 : XOR2_X1 port map( A1 => n22207, A2 => n18027, Z => n18229);
   U15723 : XNOR2_X1 port map( A1 => n10494, A2 => n19350, ZN => n3464);
   U15752 : XOR2_X1 port map( A1 => n23325, A2 => n6530, Z => n19861);
   U15768 : XOR2_X1 port map( A1 => n6507, A2 => n10752, Z => n12501);
   U15770 : NOR2_X2 port map( A1 => n17519, A2 => n14917, ZN => n17432);
   U15771 : INV_X2 port map( I => n12473, ZN => n14917);
   U15772 : XOR2_X1 port map( A1 => n11002, A2 => n11003, Z => n12473);
   U15789 : XOR2_X1 port map( A1 => n23411, A2 => n4285, Z => n23329);
   U15797 : AND2_X1 port map( A1 => n15760, A2 => n10905, Z => n10632);
   U15801 : AND2_X1 port map( A1 => n9772, A2 => n26076, Z => n14025);
   U15818 : NOR2_X1 port map( A1 => n8584, A2 => n23333, ZN => n23492);
   U15821 : AOI21_X1 port map( A1 => n8588, A2 => n20620, B => n24597, ZN => 
                           n23333);
   U15831 : NAND2_X2 port map( A1 => n23335, A2 => n24444, ZN => n12559);
   U15842 : XOR2_X1 port map( A1 => n23336, A2 => n4637, Z => n2864);
   U15848 : XOR2_X1 port map( A1 => n4636, A2 => n4635, Z => n23336);
   U15863 : XOR2_X1 port map( A1 => Plaintext(108), A2 => Key(108), Z => n13274
                           );
   U15865 : AND2_X1 port map( A1 => n18055, A2 => n18774, Z => n24440);
   U15871 : OR2_X1 port map( A1 => n28542, A2 => n14648, Z => n12244);
   U15879 : XOR2_X1 port map( A1 => n5688, A2 => n5686, Z => n10104);
   U15880 : INV_X2 port map( I => n23341, ZN => n577);
   U15881 : XNOR2_X1 port map( A1 => Plaintext(112), A2 => Key(112), ZN => 
                           n23341);
   U15888 : XOR2_X1 port map( A1 => n13748, A2 => n23347, Z => n10640);
   U15918 : INV_X1 port map( I => n21650, ZN => n23354);
   U15925 : XNOR2_X1 port map( A1 => n11222, A2 => n8111, ZN => n97);
   U15933 : NOR2_X1 port map( A1 => n28302, A2 => n17868, ZN => n23356);
   U15960 : XOR2_X1 port map( A1 => n24098, A2 => n16797, Z => n23393);
   U15963 : XOR2_X1 port map( A1 => n16881, A2 => n17032, Z => n16797);
   U15965 : XOR2_X1 port map( A1 => n2994, A2 => n2225, Z => n16856);
   U15970 : NAND2_X1 port map( A1 => n17887, A2 => n22817, ZN => n23365);
   U16016 : NAND2_X2 port map( A1 => n15113, A2 => n15115, ZN => n20213);
   U16017 : XOR2_X1 port map( A1 => n16993, A2 => n16853, Z => n4094);
   U16018 : OAI21_X2 port map( A1 => n6397, A2 => n6396, B => n6395, ZN => 
                           n16993);
   U16031 : XOR2_X1 port map( A1 => n21857, A2 => n17054, Z => n23373);
   U16033 : XOR2_X1 port map( A1 => n12099, A2 => n21255, Z => n13300);
   U16036 : AND2_X1 port map( A1 => n977, A2 => n11225, Z => n19695);
   U16061 : INV_X2 port map( I => n23713, ZN => n2478);
   U16066 : XOR2_X1 port map( A1 => n1651, A2 => n10443, Z => n14000);
   U16080 : OR2_X1 port map( A1 => n22811, A2 => n5807, Z => n9648);
   U16086 : XOR2_X1 port map( A1 => n23383, A2 => n11226, Z => Ciphertext(107))
                           ;
   U16092 : AOI21_X2 port map( A1 => n17915, A2 => n17783, B => n7358, ZN => 
                           n23386);
   U16099 : NOR2_X1 port map( A1 => n10539, A2 => n17183, ZN => n9767);
   U16122 : XOR2_X1 port map( A1 => n23393, A2 => n14082, Z => n16406);
   U16127 : XOR2_X1 port map( A1 => n27573, A2 => n14575, Z => n3925);
   U16140 : NOR2_X1 port map( A1 => n5866, A2 => n17411, ZN => n5865);
   U16144 : NAND2_X2 port map( A1 => n17292, A2 => n14367, ZN => n17402);
   U16152 : XOR2_X1 port map( A1 => n20537, A2 => n21197, Z => n21256);
   U16157 : NAND2_X2 port map( A1 => n12827, A2 => n12829, ZN => n21197);
   U16166 : INV_X4 port map( I => n17513, ZN => n24018);
   U16188 : XOR2_X1 port map( A1 => n9707, A2 => n9711, Z => n19399);
   U16198 : NAND3_X2 port map( A1 => n9686, A2 => n9684, A3 => n13673, ZN => 
                           n17665);
   U16209 : INV_X1 port map( I => n23407, ZN => n9518);
   U16210 : NAND3_X1 port map( A1 => n23408, A2 => n7908, A3 => n7927, ZN => 
                           n23407);
   U16212 : XOR2_X1 port map( A1 => n853, A2 => n8655, Z => n23858);
   U16223 : XOR2_X1 port map( A1 => n19278, A2 => n19277, Z => n23409);
   U16227 : XOR2_X1 port map( A1 => n23198, A2 => n9161, Z => n23411);
   U16229 : NAND2_X1 port map( A1 => n23413, A2 => n15918, ZN => n12083);
   U16230 : XOR2_X1 port map( A1 => n20714, A2 => n21301, Z => n7590);
   U16231 : NAND2_X2 port map( A1 => n13646, A2 => n18687, ZN => n7799);
   U16234 : OAI21_X1 port map( A1 => n1258, A2 => n14989, B => n11940, ZN => 
                           n23413);
   U16235 : XOR2_X1 port map( A1 => n6087, A2 => n21922, Z => n23414);
   U16237 : NAND2_X1 port map( A1 => n9359, A2 => n9991, ZN => n9990);
   U16260 : XOR2_X1 port map( A1 => n27415, A2 => n4768, Z => n10852);
   U16288 : NOR2_X1 port map( A1 => n6354, A2 => n25829, ZN => n23419);
   U16298 : INV_X2 port map( I => n23420, ZN => n1460);
   U16300 : OAI21_X2 port map( A1 => n21012, A2 => n21135, B => n27266, ZN => 
                           n21015);
   U16301 : OAI21_X2 port map( A1 => n874, A2 => n19033, B => n23422, ZN => 
                           n9971);
   U16304 : NAND3_X1 port map( A1 => n19720, A2 => n12467, A3 => n6219, ZN => 
                           n23423);
   U16307 : XOR2_X1 port map( A1 => n4422, A2 => n23429, Z => n4420);
   U16317 : NAND2_X1 port map( A1 => n23433, A2 => n427, ZN => n23432);
   U16319 : NAND2_X1 port map( A1 => n24294, A2 => n25411, ZN => n23433);
   U16320 : NAND2_X2 port map( A1 => n23435, A2 => n4032, ZN => n3914);
   U16340 : NAND2_X1 port map( A1 => n11736, A2 => n11735, ZN => n23438);
   U16342 : INV_X2 port map( I => n4274, ZN => n20253);
   U16351 : NAND2_X1 port map( A1 => n4378, A2 => n4379, ZN => n10819);
   U16363 : AOI21_X2 port map( A1 => n23453, A2 => n18621, B => n13390, ZN => 
                           n12453);
   U16370 : INV_X4 port map( I => n3982, ZN => n13758);
   U16446 : OR3_X1 port map( A1 => n11391, A2 => n14180, A3 => n27658, Z => 
                           n9457);
   U16455 : XOR2_X1 port map( A1 => n4866, A2 => n4865, Z => n20411);
   U16469 : NAND3_X2 port map( A1 => n5395, A2 => n12335, A3 => n5394, ZN => 
                           n6745);
   U16474 : OR2_X1 port map( A1 => n8604, A2 => n18715, Z => n4291);
   U16476 : XOR2_X1 port map( A1 => n23478, A2 => n6944, Z => n6945);
   U16480 : XOR2_X1 port map( A1 => n18175, A2 => n6943, Z => n23478);
   U16484 : AOI21_X1 port map( A1 => n13505, A2 => n22811, B => n8594, ZN => 
                           n2536);
   U16533 : XOR2_X1 port map( A1 => n23482, A2 => n4696, Z => n6259);
   U16541 : NAND3_X1 port map( A1 => n18930, A2 => n2484, A3 => n6216, ZN => 
                           n3032);
   U16569 : NOR2_X2 port map( A1 => n1968, A2 => n6661, ZN => n3179);
   U16571 : XOR2_X1 port map( A1 => n2367, A2 => n23485, Z => n20469);
   U16580 : XOR2_X1 port map( A1 => n2366, A2 => n2365, Z => n23485);
   U16602 : AOI21_X2 port map( A1 => n7591, A2 => n26036, B => n10555, ZN => 
                           n9604);
   U16604 : XOR2_X1 port map( A1 => n6745, A2 => n12674, Z => n18085);
   U16609 : XOR2_X1 port map( A1 => n23492, A2 => n13738, Z => Ciphertext(10));
   U16633 : NOR2_X2 port map( A1 => n17191, A2 => n23497, ZN => n17724);
   U16668 : INV_X1 port map( I => n21327, ZN => n23499);
   U16677 : INV_X2 port map( I => n3224, ZN => n23500);
   U16683 : INV_X2 port map( I => n25384, ZN => n15331);
   U16691 : XOR2_X1 port map( A1 => Plaintext(129), A2 => Key(129), Z => n13209
                           );
   U16692 : INV_X2 port map( I => n24568, ZN => n9041);
   U16718 : INV_X2 port map( I => n23504, ZN => n7326);
   U16729 : XOR2_X1 port map( A1 => n13156, A2 => n13154, Z => n23504);
   U16738 : NAND2_X2 port map( A1 => n16250, A2 => n16251, ZN => n124);
   U16741 : INV_X2 port map( I => n1496, ZN => n11054);
   U16742 : NAND2_X2 port map( A1 => n1495, A2 => n1493, ZN => n1496);
   U16744 : NAND2_X2 port map( A1 => n10491, A2 => n10492, ZN => n14654);
   U16746 : XOR2_X1 port map( A1 => n23508, A2 => n20617, Z => Ciphertext(7));
   U16747 : OAI22_X1 port map( A1 => n20627, A2 => n4820, B1 => n20616, B2 => 
                           n20615, ZN => n23508);
   U16751 : XOR2_X1 port map( A1 => n8957, A2 => n12114, Z => n19420);
   U16757 : NOR2_X1 port map( A1 => n19955, A2 => n19827, ZN => n19466);
   U16771 : XOR2_X1 port map( A1 => n14950, A2 => n4179, Z => n11189);
   U16778 : XOR2_X1 port map( A1 => n23515, A2 => n20554, Z => n14916);
   U16780 : XOR2_X1 port map( A1 => n20771, A2 => n20537, Z => n23515);
   U16799 : NAND2_X2 port map( A1 => n9433, A2 => n9431, ZN => n16565);
   U16811 : XOR2_X1 port map( A1 => n1526, A2 => n1525, Z => n23518);
   U16819 : OR2_X1 port map( A1 => n5368, A2 => n5317, Z => n11732);
   U16832 : XNOR2_X1 port map( A1 => n22802, A2 => n20961, ZN => n9081);
   U16845 : XOR2_X1 port map( A1 => n19424, A2 => n19423, Z => n19425);
   U16897 : XOR2_X1 port map( A1 => n23528, A2 => n17042, Z => n17412);
   U16917 : NAND2_X1 port map( A1 => n11286, A2 => n22364, ZN => n3401);
   U16925 : INV_X2 port map( I => n23535, ZN => n17302);
   U16930 : XNOR2_X1 port map( A1 => n6515, A2 => n6513, ZN => n23535);
   U16934 : NAND2_X2 port map( A1 => n23536, A2 => n2415, ZN => n21111);
   U16961 : NAND2_X2 port map( A1 => n17306, A2 => n17302, ZN => n16996);
   U16962 : NAND2_X1 port map( A1 => n20624, A2 => n939, ZN => n8588);
   U16975 : NOR2_X1 port map( A1 => n16326, A2 => n14326, ZN => n16170);
   U16986 : XOR2_X1 port map( A1 => n18040, A2 => n13449, Z => n13410);
   U16990 : XOR2_X1 port map( A1 => n10088, A2 => n9038, Z => n9037);
   U17025 : NOR2_X2 port map( A1 => n24045, A2 => n23544, ZN => n19144);
   U17027 : XOR2_X1 port map( A1 => n18313, A2 => n18310, Z => n2159);
   U17030 : NOR2_X2 port map( A1 => n10681, A2 => n4710, ZN => n23548);
   U17036 : NOR2_X2 port map( A1 => n19660, A2 => n9193, ZN => n23916);
   U17047 : OAI22_X2 port map( A1 => n17759, A2 => n788, B1 => n17758, B2 => 
                           n23978, ZN => n18061);
   U17052 : NAND2_X2 port map( A1 => n23836, A2 => n3590, ZN => n13927);
   U17061 : AOI22_X2 port map( A1 => n23552, A2 => n19830, B1 => n19946, B2 => 
                           n7376, ZN => n20059);
   U17062 : NAND2_X2 port map( A1 => n23553, A2 => n14977, ZN => n14401);
   U17072 : XOR2_X1 port map( A1 => n18330, A2 => n23554, Z => n9242);
   U17074 : INV_X1 port map( I => n14340, ZN => n23554);
   U17081 : NOR3_X1 port map( A1 => n19981, A2 => n4021, A3 => n20023, ZN => 
                           n3271);
   U17084 : XOR2_X1 port map( A1 => n16826, A2 => n4179, Z => n16751);
   U17097 : OR2_X1 port map( A1 => n16707, A2 => n7132, Z => n7054);
   U17098 : AND2_X1 port map( A1 => n899, A2 => n17345, Z => n17574);
   U17102 : NAND2_X1 port map( A1 => n5134, A2 => n14070, ZN => n5133);
   U17116 : NAND2_X2 port map( A1 => n2632, A2 => n14595, ZN => n11044);
   U17118 : NAND2_X2 port map( A1 => n24661, A2 => n451, ZN => n4353);
   U17130 : NOR2_X1 port map( A1 => n1459, A2 => n1460, ZN => n523);
   U17156 : XOR2_X1 port map( A1 => n23686, A2 => n23849, Z => n13948);
   U17164 : NAND2_X1 port map( A1 => n20672, A2 => n7342, ZN => n23573);
   U17168 : XOR2_X1 port map( A1 => n14775, A2 => n17884, Z => n23574);
   U17182 : OAI21_X1 port map( A1 => n13986, A2 => n21455, B => n6080, ZN => 
                           n7946);
   U17242 : NAND3_X2 port map( A1 => n1706, A2 => n3716, A3 => n3717, ZN => 
                           n10456);
   U17247 : NOR2_X2 port map( A1 => n1378, A2 => n1377, ZN => n23871);
   U17256 : XOR2_X1 port map( A1 => n21238, A2 => n4964, Z => n23589);
   U17261 : AOI21_X2 port map( A1 => n14519, A2 => n14178, B => n12272, ZN => 
                           n15821);
   U17264 : XOR2_X1 port map( A1 => n7604, A2 => n7605, Z => n24373);
   U17271 : NAND2_X1 port map( A1 => n24553, A2 => n20269, ZN => n23593);
   U17282 : NAND2_X1 port map( A1 => n14132, A2 => n21774, ZN => n14998);
   U17288 : XOR2_X1 port map( A1 => n15177, A2 => n10525, Z => n14194);
   U17292 : XOR2_X1 port map( A1 => n23601, A2 => n20666, Z => Ciphertext(17));
   U17293 : AOI22_X1 port map( A1 => n8482, A2 => n23119, B1 => n8481, B2 => 
                           n20664, ZN => n23601);
   U17296 : NAND2_X2 port map( A1 => n3329, A2 => n5690, ZN => n13757);
   U17330 : NAND2_X2 port map( A1 => n7661, A2 => n7662, ZN => n3982);
   U17338 : NAND2_X2 port map( A1 => n15111, A2 => n17445, ZN => n13129);
   U17339 : XOR2_X1 port map( A1 => n19534, A2 => n23607, Z => n663);
   U17342 : XOR2_X1 port map( A1 => n10038, A2 => n2389, Z => n23607);
   U17369 : NAND2_X2 port map( A1 => n5859, A2 => n23613, ZN => n18947);
   U17372 : XOR2_X1 port map( A1 => n23614, A2 => n25840, Z => Ciphertext(73));
   U17385 : AOI22_X2 port map( A1 => n14765, A2 => n17670, B1 => n28401, B2 => 
                           n17669, ZN => n18038);
   U17397 : INV_X2 port map( I => n23622, ZN => n10251);
   U17403 : INV_X2 port map( I => n26639, ZN => n23624);
   U17435 : INV_X2 port map( I => n24672, ZN => n18757);
   U17443 : NAND2_X1 port map( A1 => n15992, A2 => n4281, ZN => n23630);
   U17448 : XOR2_X1 port map( A1 => n17039, A2 => n23352, Z => n17150);
   U17453 : XNOR2_X1 port map( A1 => n10378, A2 => n18314, ZN => n5022);
   U17456 : OAI21_X2 port map( A1 => n14234, A2 => n11782, B => n11781, ZN => 
                           n18314);
   U17457 : AOI21_X1 port map( A1 => n6798, A2 => n21532, B => n23634, ZN => 
                           n6795);
   U17465 : XOR2_X1 port map( A1 => n13982, A2 => n12049, Z => n10500);
   U17466 : XOR2_X1 port map( A1 => n16818, A2 => n4876, Z => n17131);
   U17469 : NAND2_X2 port map( A1 => n16485, A2 => n7855, ZN => n16818);
   U17470 : NAND2_X2 port map( A1 => n23635, A2 => n15241, ZN => n15239);
   U17471 : XOR2_X1 port map( A1 => n23637, A2 => n4903, Z => n2712);
   U17477 : INV_X2 port map( I => n23638, ZN => n14962);
   U17490 : NAND2_X2 port map( A1 => n12083, A2 => n15858, ZN => n12224);
   U17491 : XOR2_X1 port map( A1 => n19484, A2 => n19483, Z => n489);
   U17500 : AND2_X1 port map( A1 => n17548, A2 => n24517, Z => n24371);
   U17511 : XOR2_X1 port map( A1 => n23646, A2 => n21265, Z => n11326);
   U17523 : XOR2_X1 port map( A1 => n10208, A2 => n26726, Z => n8788);
   U17536 : INV_X1 port map( I => n23647, ZN => n1927);
   U17558 : XOR2_X1 port map( A1 => n20521, A2 => n20522, Z => n11862);
   U17571 : INV_X2 port map( I => n12759, ZN => n23648);
   U17583 : NAND2_X2 port map( A1 => n14255, A2 => n9772, ZN => n17799);
   U17586 : NOR2_X1 port map( A1 => n9267, A2 => n12018, ZN => n23650);
   U17594 : INV_X2 port map( I => n21716, ZN => n23653);
   U17599 : NOR2_X1 port map( A1 => n18530, A2 => n18581, ZN => n13360);
   U17603 : XOR2_X1 port map( A1 => n18198, A2 => n23656, Z => n6174);
   U17608 : XOR2_X1 port map( A1 => n5529, A2 => n23657, Z => n23656);
   U17612 : INV_X1 port map( I => n20941, ZN => n23657);
   U17614 : OR2_X1 port map( A1 => n19021, A2 => n28499, Z => n9152);
   U17619 : AOI21_X2 port map( A1 => n9651, A2 => n2037, B => n8093, ZN => 
                           n2036);
   U17634 : XNOR2_X1 port map( A1 => n19385, A2 => n19386, ZN => n24279);
   U17638 : XOR2_X1 port map( A1 => n13658, A2 => n16976, Z => n13493);
   U17654 : NAND3_X1 port map( A1 => n1040, A2 => n24585, A3 => n5639, ZN => 
                           n5766);
   U17664 : INV_X1 port map( I => n7087, ZN => n23666);
   U17678 : OR2_X1 port map( A1 => n12670, A2 => n22253, Z => n8148);
   U17679 : XOR2_X1 port map( A1 => n12114, A2 => n9283, Z => n23667);
   U17701 : XOR2_X1 port map( A1 => n23668, A2 => n17603, Z => n18427);
   U17716 : NAND2_X1 port map( A1 => n26081, A2 => n17510, ZN => n17262);
   U17723 : NOR2_X1 port map( A1 => n814, A2 => n6976, ZN => n2315);
   U17726 : NAND2_X1 port map( A1 => n21508, A2 => n8721, ZN => n23671);
   U17729 : NAND3_X1 port map( A1 => n10173, A2 => n22848, A3 => n15199, ZN => 
                           n9317);
   U17748 : NAND2_X2 port map( A1 => n14088, A2 => n23680, ZN => n24324);
   U17770 : NAND2_X2 port map( A1 => n8630, A2 => n23683, ZN => n21311);
   U17775 : XOR2_X1 port map( A1 => n337, A2 => n11679, Z => n17051);
   U17778 : NAND2_X2 port map( A1 => n14853, A2 => n16247, ZN => n11679);
   U17779 : INV_X2 port map( I => n23684, ZN => n17474);
   U17799 : NOR2_X2 port map( A1 => n1035, A2 => n17477, ZN => n14275);
   U17802 : XOR2_X1 port map( A1 => n16439, A2 => n23694, Z => n13276);
   U17803 : XOR2_X1 port map( A1 => n4877, A2 => n26656, Z => n23694);
   U17813 : XOR2_X1 port map( A1 => n23697, A2 => n1725, Z => n12596);
   U17815 : XOR2_X1 port map( A1 => n22926, A2 => n17044, Z => n23697);
   U17819 : XOR2_X1 port map( A1 => n23698, A2 => n23816, Z => Ciphertext(53));
   U17820 : NOR2_X1 port map( A1 => n8161, A2 => n8160, ZN => n23698);
   U17851 : XOR2_X1 port map( A1 => n7244, A2 => n13122, Z => n23704);
   U17852 : AND2_X1 port map( A1 => n10952, A2 => n17372, Z => n23853);
   U17875 : AOI22_X2 port map( A1 => n7499, A2 => n11685, B1 => n7500, B2 => 
                           n14308, ZN => n7911);
   U17894 : XOR2_X1 port map( A1 => n16940, A2 => n14733, Z => n4601);
   U17905 : NAND2_X2 port map( A1 => n4212, A2 => n9050, ZN => n18904);
   U17919 : XOR2_X1 port map( A1 => n6535, A2 => n22512, Z => n20025);
   U17922 : NAND2_X2 port map( A1 => n23716, A2 => n1380, ZN => n1716);
   U17930 : OR2_X1 port map( A1 => n8534, A2 => n23474, Z => n23718);
   U17936 : NOR3_X1 port map( A1 => n16704, A2 => n3443, A3 => n10868, ZN => 
                           n1424);
   U17957 : NAND2_X2 port map( A1 => n2623, A2 => n2624, ZN => n4822);
   U17958 : OAI21_X1 port map( A1 => n5816, A2 => n25314, B => n23726, ZN => 
                           n1583);
   U17959 : XOR2_X1 port map( A1 => n8808, A2 => n23727, Z => n8805);
   U17960 : XOR2_X1 port map( A1 => n8807, A2 => n21818, Z => n23727);
   U17969 : NAND2_X1 port map( A1 => n540, A2 => n28353, ZN => n17342);
   U17975 : NOR2_X2 port map( A1 => n858, A2 => n14663, ZN => n7796);
   U17983 : XOR2_X1 port map( A1 => n23730, A2 => n11141, Z => n11105);
   U17989 : XOR2_X1 port map( A1 => n13808, A2 => n23731, Z => n23730);
   U17994 : INV_X1 port map( I => n21336, ZN => n23731);
   U18037 : XOR2_X1 port map( A1 => n23735, A2 => n155, Z => n5946);
   U18044 : NOR2_X2 port map( A1 => n14019, A2 => n14020, ZN => n19478);
   U18055 : OAI21_X2 port map( A1 => n23736, A2 => n17900, B => n17769, ZN => 
                           n24363);
   U18056 : NOR2_X2 port map( A1 => n10659, A2 => n17768, ZN => n23736);
   U18059 : XOR2_X1 port map( A1 => n16911, A2 => n26713, Z => n23737);
   U18142 : NAND2_X2 port map( A1 => n6907, A2 => n247, ZN => n6906);
   U18164 : NAND3_X2 port map( A1 => n6732, A2 => n6733, A3 => n6731, ZN => 
                           n4953);
   U18165 : OAI21_X1 port map( A1 => n10663, A2 => n14939, B => n13444, ZN => 
                           n5482);
   U18183 : XOR2_X1 port map( A1 => n16767, A2 => n8309, Z => n6868);
   U18187 : XOR2_X1 port map( A1 => n9477, A2 => n7150, Z => n12289);
   U18205 : XOR2_X1 port map( A1 => n23755, A2 => n22826, Z => n3155);
   U18208 : XOR2_X1 port map( A1 => n8396, A2 => n19443, Z => n23755);
   U18212 : XOR2_X1 port map( A1 => n20006, A2 => n20007, Z => n20008);
   U18230 : INV_X4 port map( I => n10289, ZN => n23761);
   U18235 : NAND2_X1 port map( A1 => n23757, A2 => n23879, ZN => n16212);
   U18239 : OR2_X1 port map( A1 => n11518, A2 => n16339, Z => n23757);
   U18240 : AND2_X1 port map( A1 => n27460, A2 => n9140, Z => n5715);
   U18253 : NAND2_X1 port map( A1 => n18538, A2 => n18539, ZN => n23760);
   U18268 : NAND2_X2 port map( A1 => n6303, A2 => n9000, ZN => n13721);
   U18289 : XOR2_X1 port map( A1 => n2667, A2 => n2668, Z => n2666);
   U18367 : NAND2_X2 port map( A1 => n4226, A2 => n6057, ZN => n20057);
   U18410 : AOI21_X1 port map( A1 => n10210, A2 => n22736, B => n27380, ZN => 
                           n23784);
   U18428 : XOR2_X1 port map( A1 => n2742, A2 => n23788, Z => n9612);
   U18435 : NAND2_X1 port map( A1 => n10775, A2 => n10774, ZN => n23788);
   U18483 : XOR2_X1 port map( A1 => n18173, A2 => n14215, Z => n12633);
   U18491 : NOR2_X2 port map( A1 => n24126, A2 => n17820, ZN => n14215);
   U18500 : INV_X1 port map( I => n10338, ZN => n16241);
   U18504 : XOR2_X1 port map( A1 => n15779, A2 => Key(155), Z => n10338);
   U18518 : OAI21_X2 port map( A1 => n12154, A2 => n12153, B => n23798, ZN => 
                           n12637);
   U18522 : XOR2_X1 port map( A1 => n8776, A2 => n9774, Z => n17108);
   U18547 : NAND2_X2 port map( A1 => n13110, A2 => n19650, ZN => n19735);
   U18567 : XOR2_X1 port map( A1 => n11787, A2 => n1371, Z => n4398);
   U18609 : NOR2_X1 port map( A1 => n24351, A2 => n16654, ZN => n11068);
   U18614 : NAND2_X1 port map( A1 => n3099, A2 => n13383, ZN => n23812);
   U18624 : XOR2_X1 port map( A1 => n19421, A2 => n23816, Z => n19423);
   U18627 : INV_X1 port map( I => n20880, ZN => n23816);
   U18633 : XNOR2_X1 port map( A1 => n20404, A2 => n12365, ZN => n24153);
   U18645 : NAND2_X2 port map( A1 => n6443, A2 => n6444, ZN => n6445);
   U18651 : NOR2_X1 port map( A1 => n11440, A2 => n11438, ZN => n23820);
   U18653 : INV_X1 port map( I => n8892, ZN => n23824);
   U18662 : XOR2_X1 port map( A1 => n19024, A2 => n15244, Z => n23827);
   U18663 : NAND2_X2 port map( A1 => n20623, A2 => n15287, ZN => n20620);
   U18667 : NAND2_X2 port map( A1 => n10919, A2 => n10918, ZN => n11580);
   U18679 : XOR2_X1 port map( A1 => n12681, A2 => n18109, Z => n4133);
   U18686 : OAI22_X2 port map( A1 => n4001, A2 => n1558, B1 => n1412, B2 => 
                           n6708, ZN => n18637);
   U18692 : XOR2_X1 port map( A1 => n4094, A2 => n4093, Z => n23829);
   U18705 : XOR2_X1 port map( A1 => n23830, A2 => n18350, Z => n18578);
   U18713 : XOR2_X1 port map( A1 => n18347, A2 => n18348, Z => n23830);
   U18715 : OAI21_X2 port map( A1 => n24162, A2 => n17358, B => n8609, ZN => 
                           n23831);
   U18718 : NAND2_X2 port map( A1 => n9425, A2 => n25352, ZN => n21043);
   U18744 : XOR2_X1 port map( A1 => n17142, A2 => n27387, Z => n17054);
   U18753 : AND2_X1 port map( A1 => n14724, A2 => n1032, Z => n17191);
   U18755 : XOR2_X1 port map( A1 => n8748, A2 => n12344, Z => n2064);
   U18756 : XOR2_X1 port map( A1 => n12925, A2 => n23839, Z => n15387);
   U18758 : INV_X1 port map( I => n14598, ZN => n23839);
   U18760 : AOI21_X2 port map( A1 => n17410, A2 => n27970, B => n15305, ZN => 
                           n24127);
   U18784 : XOR2_X1 port map( A1 => n19321, A2 => n13117, Z => n13116);
   U18785 : XOR2_X1 port map( A1 => n4626, A2 => n2507, Z => n19321);
   U18842 : NOR3_X2 port map( A1 => n15302, A2 => n15301, A3 => n16204, ZN => 
                           n16836);
   U18848 : OAI21_X2 port map( A1 => n23853, A2 => n23852, B => n17374, ZN => 
                           n17957);
   U18850 : INV_X4 port map( I => n24181, ZN => n15041);
   U18871 : XOR2_X1 port map( A1 => n23858, A2 => n12733, Z => n6164);
   U18872 : NAND2_X2 port map( A1 => n23859, A2 => n6226, ZN => n7987);
   U18878 : XOR2_X1 port map( A1 => n16944, A2 => n23860, Z => n16841);
   U18893 : NOR2_X1 port map( A1 => n3572, A2 => n16287, ZN => n15860);
   U18902 : NAND2_X1 port map( A1 => n15255, A2 => n17530, ZN => n9359);
   U18929 : INV_X1 port map( I => n10105, ZN => n23868);
   U18944 : XOR2_X1 port map( A1 => n17053, A2 => n12831, Z => n16893);
   U18951 : NOR2_X1 port map( A1 => n23948, A2 => n14512, ZN => n23946);
   U18971 : NAND3_X1 port map( A1 => n25795, A2 => n4537, A3 => n20171, ZN => 
                           n3933);
   U18973 : AOI22_X2 port map( A1 => n11602, A2 => n23672, B1 => n19103, B2 => 
                           n11554, ZN => n5433);
   U18984 : OAI22_X1 port map( A1 => n19790, A2 => n2320, B1 => n19624, B2 => 
                           n23322, ZN => n12401);
   U19000 : XOR2_X1 port map( A1 => n23873, A2 => n20912, Z => Ciphertext(58));
   U19002 : INV_X2 port map( I => n23874, ZN => n4634);
   U19005 : XOR2_X1 port map( A1 => Plaintext(126), A2 => Key(126), Z => n23874
                           );
   U19016 : XOR2_X1 port map( A1 => n11999, A2 => n14813, Z => n4222);
   U19020 : XOR2_X1 port map( A1 => n5212, A2 => n21855, Z => n16955);
   U19023 : INV_X1 port map( I => n18417, ZN => n13327);
   U19037 : NAND2_X2 port map( A1 => n5995, A2 => n5993, ZN => n2284);
   U19041 : NAND2_X1 port map( A1 => n12006, A2 => n13147, ZN => n12005);
   U19043 : NOR2_X1 port map( A1 => n20187, A2 => n26970, ZN => n23877);
   U19050 : AOI21_X1 port map( A1 => n10101, A2 => n21565, B => n28308, ZN => 
                           n10100);
   U19068 : NAND2_X1 port map( A1 => n11719, A2 => n9618, ZN => n14070);
   U19077 : NAND2_X2 port map( A1 => n5632, A2 => n17651, ZN => n5631);
   U19084 : NOR3_X1 port map( A1 => n8947, A2 => n8946, A3 => n20802, ZN => 
                           n24118);
   U19091 : XOR2_X1 port map( A1 => n23881, A2 => n637, Z => n9024);
   U19092 : XOR2_X1 port map( A1 => n28393, A2 => n28355, Z => n23881);
   U19098 : NAND2_X1 port map( A1 => n23883, A2 => n12519, ZN => n20672);
   U19127 : XOR2_X1 port map( A1 => n18317, A2 => n21679, Z => n23888);
   U19145 : INV_X1 port map( I => n17082, ZN => n24163);
   U19151 : NOR2_X2 port map( A1 => n23893, A2 => n23892, ZN => n23891);
   U19153 : NOR2_X1 port map( A1 => n17764, A2 => n17963, ZN => n23892);
   U19180 : INV_X2 port map( I => n23895, ZN => n2654);
   U19188 : XOR2_X1 port map( A1 => Plaintext(189), A2 => Key(189), Z => n23895
                           );
   U19194 : NAND2_X2 port map( A1 => n23897, A2 => n12775, ZN => n12482);
   U19203 : NAND2_X1 port map( A1 => n11006, A2 => n11007, ZN => n23897);
   U19209 : XOR2_X1 port map( A1 => n6126, A2 => n20377, Z => n23898);
   U19211 : NOR2_X1 port map( A1 => n13032, A2 => n26462, ZN => n8542);
   U19213 : AOI21_X2 port map( A1 => n1961, A2 => n1960, B => n23899, ZN => 
                           n19516);
   U19225 : XOR2_X1 port map( A1 => n13152, A2 => n23903, Z => n15343);
   U19235 : XOR2_X1 port map( A1 => n13150, A2 => n13151, Z => n23903);
   U19242 : XOR2_X1 port map( A1 => n10076, A2 => n23904, Z => n17202);
   U19249 : XOR2_X1 port map( A1 => n10490, A2 => n11397, Z => n23904);
   U19257 : XOR2_X1 port map( A1 => n11899, A2 => n11896, Z => n20709);
   U19259 : XOR2_X1 port map( A1 => n9339, A2 => n19304, Z => n3020);
   U19263 : NAND2_X2 port map( A1 => n23910, A2 => n23908, ZN => n16058);
   U19275 : OAI21_X2 port map( A1 => n24388, A2 => n7229, B => n15497, ZN => 
                           n16447);
   U19300 : OAI21_X2 port map( A1 => n24996, A2 => n24844, B => n23918, ZN => 
                           n16247);
   U19303 : XOR2_X1 port map( A1 => n4833, A2 => n1715, Z => n15088);
   U19306 : OR2_X1 port map( A1 => n4634, A2 => n25384, Z => n23922);
   U19313 : XOR2_X1 port map( A1 => n10445, A2 => n22780, Z => n11278);
   U19323 : XOR2_X1 port map( A1 => n20533, A2 => n20454, Z => n6759);
   U19348 : AOI21_X2 port map( A1 => n15376, A2 => n19599, B => n23934, ZN => 
                           n11148);
   U19352 : XOR2_X1 port map( A1 => n10360, A2 => n23940, Z => n3313);
   U19365 : XOR2_X1 port map( A1 => n491, A2 => n26634, Z => n4716);
   U19366 : NAND2_X1 port map( A1 => n26625, A2 => n9924, ZN => n14163);
   U19395 : NOR2_X2 port map( A1 => n4715, A2 => n23863, ZN => n622);
   U19415 : AND2_X1 port map( A1 => n2762, A2 => n16695, Z => n23958);
   U19444 : INV_X2 port map( I => n21082, ZN => n13476);
   U19464 : XOR2_X1 port map( A1 => n19524, A2 => n23691, Z => n19508);
   U19468 : XOR2_X1 port map( A1 => n9125, A2 => n12915, Z => n23967);
   U19483 : XOR2_X1 port map( A1 => n23969, A2 => n1276, Z => Ciphertext(142));
   U19484 : NOR2_X1 port map( A1 => n10834, A2 => n10832, ZN => n23969);
   U19493 : NOR2_X1 port map( A1 => n5978, A2 => n25013, ZN => n23971);
   U19495 : XOR2_X1 port map( A1 => n4358, A2 => n4360, Z => n7383);
   U19498 : NOR2_X1 port map( A1 => n15457, A2 => n23748, ZN => n4499);
   U19499 : XOR2_X1 port map( A1 => n2015, A2 => n4497, Z => n2941);
   U19517 : XOR2_X1 port map( A1 => n18244, A2 => n2140, Z => n24122);
   U19520 : INV_X2 port map( I => n16989, ZN => n1237);
   U19524 : NOR2_X2 port map( A1 => n24051, A2 => n5997, ZN => n16989);
   U19529 : INV_X2 port map( I => n20107, ZN => n5048);
   U19534 : XOR2_X1 port map( A1 => n12181, A2 => n4137, Z => n20510);
   U19535 : NOR2_X2 port map( A1 => n9768, A2 => n16316, ZN => n7631);
   U19537 : NAND2_X1 port map( A1 => n24309, A2 => n14156, ZN => n15091);
   U19545 : NOR2_X2 port map( A1 => n1016, A2 => n8254, ZN => n10009);
   U19553 : XOR2_X1 port map( A1 => n17108, A2 => n23986, Z => n17113);
   U19554 : XOR2_X1 port map( A1 => n25386, A2 => n2225, Z => n23986);
   U19560 : OAI22_X2 port map( A1 => n3948, A2 => n16685, B1 => n16176, B2 => 
                           n1252, ZN => n60);
   U19562 : AOI21_X2 port map( A1 => n11436, A2 => n11435, B => n24607, ZN => 
                           n11434);
   U19580 : NOR2_X1 port map( A1 => n20312, A2 => n2525, ZN => n5354);
   U19595 : XOR2_X1 port map( A1 => n3176, A2 => n23996, Z => n11852);
   U19598 : XOR2_X1 port map( A1 => n16759, A2 => n24584, Z => n23996);
   U19604 : XOR2_X1 port map( A1 => n16829, A2 => n16793, Z => n23998);
   U19617 : NAND2_X2 port map( A1 => n7192, A2 => n7672, ZN => n20685);
   U19623 : NAND2_X1 port map( A1 => n9946, A2 => n24524, ZN => n6504);
   U19625 : XOR2_X1 port map( A1 => n15609, A2 => n4179, Z => n4525);
   U19635 : XOR2_X1 port map( A1 => n21375, A2 => n21927, Z => n24004);
   U19643 : XOR2_X1 port map( A1 => n4310, A2 => n27904, Z => n18288);
   U19644 : AOI21_X2 port map( A1 => n13326, A2 => n1260, B => n16182, ZN => 
                           n16044);
   U19661 : NOR2_X1 port map( A1 => n12145, A2 => n19918, ZN => n19733);
   U19662 : NOR2_X2 port map( A1 => n24009, A2 => n3822, ZN => n3828);
   U19668 : XOR2_X1 port map( A1 => n8902, A2 => n8903, Z => n5516);
   U19675 : INV_X2 port map( I => n24010, ZN => n13824);
   U19699 : XOR2_X1 port map( A1 => n16897, A2 => n16914, Z => n24287);
   U19704 : XOR2_X1 port map( A1 => n24013, A2 => n17058, Z => n12549);
   U19726 : AND2_X1 port map( A1 => n1634, A2 => n14032, Z => n1633);
   U19751 : NAND2_X2 port map( A1 => n12766, A2 => n10609, ZN => n16471);
   U19762 : OAI21_X2 port map( A1 => n4086, A2 => n4087, B => n4084, ZN => 
                           n20658);
   U19800 : XOR2_X1 port map( A1 => n5929, A2 => n5930, Z => n6457);
   U19803 : XOR2_X1 port map( A1 => n2350, A2 => n2348, Z => n8430);
   U19804 : XOR2_X1 port map( A1 => n8821, A2 => n8822, Z => n5209);
   U19816 : OAI21_X2 port map( A1 => n24036, A2 => n12126, B => n13878, ZN => 
                           n7516);
   U19823 : AOI21_X2 port map( A1 => n6646, A2 => n3508, B => n24208, ZN => 
                           n7065);
   U19827 : NOR2_X1 port map( A1 => n12008, A2 => n20050, ZN => n12007);
   U19842 : NOR2_X1 port map( A1 => n25493, A2 => n7120, ZN => n12562);
   U19848 : XOR2_X1 port map( A1 => n12620, A2 => n16985, Z => n4764);
   U19875 : NAND2_X2 port map( A1 => n22823, A2 => n6547, ZN => n5683);
   U19903 : XOR2_X1 port map( A1 => n13930, A2 => n9360, Z => n7340);
   U19923 : XOR2_X1 port map( A1 => n2710, A2 => n8885, Z => n21239);
   U19926 : XOR2_X1 port map( A1 => n16486, A2 => n537, Z => n24048);
   U19934 : XOR2_X1 port map( A1 => n16946, A2 => n16852, Z => n10396);
   U19947 : INV_X2 port map( I => n24052, ZN => n1637);
   U19949 : XOR2_X1 port map( A1 => Plaintext(32), A2 => Key(32), Z => n24052);
   U19951 : AND2_X1 port map( A1 => n26616, A2 => n5541, Z => n3544);
   U19955 : XOR2_X1 port map( A1 => n24582, A2 => n16887, Z => n10935);
   U19957 : OR2_X1 port map( A1 => n14792, A2 => n14397, Z => n15096);
   U19968 : OR2_X1 port map( A1 => n18966, A2 => n14272, Z => n5110);
   U19971 : XNOR2_X1 port map( A1 => n16820, A2 => n17116, ZN => n3268);
   U19974 : NAND2_X2 port map( A1 => n14842, A2 => n14841, ZN => n17116);
   U19992 : NAND2_X2 port map( A1 => n15638, A2 => n10727, ZN => n15717);
   U20001 : XOR2_X1 port map( A1 => n24080, A2 => n21384, Z => Ciphertext(18));
   U20002 : NAND2_X1 port map( A1 => n20288, A2 => n20200, ZN => n12757);
   U20011 : XOR2_X1 port map( A1 => n7385, A2 => n24060, Z => n9527);
   U20037 : NAND2_X2 port map( A1 => n25161, A2 => n19160, ZN => n2218);
   U20044 : OAI22_X2 port map( A1 => n4839, A2 => n16525, B1 => n4840, B2 => 
                           n3537, ZN => n14313);
   U20085 : OAI21_X2 port map( A1 => n24374, A2 => n15061, B => n26463, ZN => 
                           n24067);
   U20101 : INV_X2 port map( I => n5034, ZN => n9472);
   U20104 : XOR2_X1 port map( A1 => n5036, A2 => n21914, Z => n5034);
   U20129 : XOR2_X1 port map( A1 => n18249, A2 => n22191, Z => n5021);
   U20139 : XOR2_X1 port map( A1 => n8115, A2 => n10441, Z => n2374);
   U20146 : NAND2_X2 port map( A1 => n12761, A2 => n12763, ZN => n16810);
   U20150 : NAND2_X2 port map( A1 => n9888, A2 => n16359, ZN => n8605);
   U20156 : XOR2_X1 port map( A1 => n12664, A2 => n6765, Z => n17058);
   U20165 : XOR2_X1 port map( A1 => n12321, A2 => n18173, Z => n24079);
   U20168 : OAI22_X1 port map( A1 => n15927, A2 => n15926, B1 => n16133, B2 => 
                           n16132, ZN => n8086);
   U20182 : OAI22_X1 port map( A1 => n20669, A2 => n13234, B1 => n20668, B2 => 
                           n28165, ZN => n24080);
   U20191 : NOR2_X1 port map( A1 => n14196, A2 => n17966, ZN => n14195);
   U20209 : AOI21_X1 port map( A1 => n21082, A2 => n21086, B => n21088, ZN => 
                           n1339);
   U20224 : XOR2_X1 port map( A1 => n2520, A2 => n20353, Z => n12080);
   U20249 : XOR2_X1 port map( A1 => n15447, A2 => n11734, Z => n24088);
   U20250 : NAND2_X1 port map( A1 => n8408, A2 => n8406, ZN => n15946);
   U20256 : OAI21_X2 port map( A1 => n12928, A2 => n5839, B => n5838, ZN => 
                           n5837);
   U20257 : XOR2_X1 port map( A1 => n27387, A2 => n25347, Z => n2274);
   U20268 : NAND2_X1 port map( A1 => n27662, A2 => n6185, ZN => n24090);
   U20273 : OAI21_X2 port map( A1 => n2817, A2 => n2816, B => n18856, ZN => 
                           n1436);
   U20286 : INV_X1 port map( I => n3268, ZN => n16871);
   U20303 : NAND3_X2 port map( A1 => n22319, A2 => n7868, A3 => n14786, ZN => 
                           n24093);
   U20319 : OAI22_X2 port map( A1 => n2759, A2 => n361, B1 => n2570, B2 => 
                           n1079, ZN => n10040);
   U20322 : INV_X2 port map( I => n24097, ZN => n1699);
   U20338 : NOR2_X1 port map( A1 => n1618, A2 => n27710, ZN => n650);
   U20365 : NAND2_X2 port map( A1 => n17733, A2 => n347, ZN => n4899);
   U20366 : XOR2_X1 port map( A1 => n17100, A2 => n21816, Z => n24254);
   U20405 : XOR2_X1 port map( A1 => n1481, A2 => n1480, Z => n24115);
   U20538 : NOR2_X1 port map( A1 => n6442, A2 => n6512, ZN => n24117);
   U20542 : XOR2_X1 port map( A1 => n24118, A2 => n12769, Z => Ciphertext(37));
   U20576 : INV_X2 port map( I => n24120, ZN => n636);
   U20578 : NAND2_X1 port map( A1 => n13039, A2 => n8223, ZN => n13040);
   U20600 : XOR2_X1 port map( A1 => n25159, A2 => n24121, Z => n10736);
   U20611 : INV_X2 port map( I => n15652, ZN => n16677);
   U20614 : NAND2_X2 port map( A1 => n24320, A2 => n13870, ZN => n15652);
   U20616 : XOR2_X1 port map( A1 => n2690, A2 => n24122, Z => n2871);
   U20661 : NAND2_X1 port map( A1 => n8908, A2 => n25056, ZN => n24130);
   U20666 : AND2_X1 port map( A1 => n21609, A2 => n8271, Z => n21605);
   U20676 : XOR2_X1 port map( A1 => n24138, A2 => n21651, Z => Ciphertext(170))
                           ;
   U20694 : XOR2_X1 port map( A1 => n7923, A2 => n7922, Z => n9924);
   U20724 : OAI21_X2 port map( A1 => n1807, A2 => n13246, B => n19954, ZN => 
                           n24145);
   U20728 : BUF_X2 port map( I => n19400, Z => n24146);
   U20741 : XOR2_X1 port map( A1 => n17116, A2 => n6345, Z => n24148);
   U20748 : NOR2_X1 port map( A1 => n24150, A2 => n20796, ZN => n7527);
   U20749 : NOR2_X1 port map( A1 => n20798, A2 => n11147, ZN => n24150);
   U20755 : XOR2_X1 port map( A1 => n24153, A2 => n10950, Z => n24152);
   U20761 : XOR2_X1 port map( A1 => n16987, A2 => n24154, Z => n2124);
   U20794 : XOR2_X1 port map( A1 => n13851, A2 => n15604, Z => n17811);
   U20801 : INV_X2 port map( I => n24160, ZN => n14183);
   U20805 : XOR2_X1 port map( A1 => n20461, A2 => n20460, Z => n24160);
   U20811 : INV_X2 port map( I => n6490, ZN => n24166);
   U20815 : NAND2_X2 port map( A1 => n7754, A2 => n24168, ZN => n7786);
   U20821 : AND2_X1 port map( A1 => n18101, A2 => n8155, Z => n12144);
   U20830 : NAND3_X2 port map( A1 => n19095, A2 => n19097, A3 => n19096, ZN => 
                           n20043);
   U20840 : XOR2_X1 port map( A1 => n6774, A2 => n19541, Z => n4920);
   U20867 : XOR2_X1 port map( A1 => n19493, A2 => n659, Z => n24176);
   U20880 : XOR2_X1 port map( A1 => n19177, A2 => n24177, Z => n13561);
   U20890 : XOR2_X1 port map( A1 => n24275, A2 => n19477, Z => n24177);
   U20928 : AND2_X1 port map( A1 => n20745, A2 => n11820, Z => n24178);
   U20960 : XOR2_X1 port map( A1 => n7776, A2 => n19550, Z => n19503);
   U20967 : NAND3_X1 port map( A1 => n21475, A2 => n7349, A3 => n21486, ZN => 
                           n24356);
   U20993 : INV_X2 port map( I => n24199, ZN => n540);
   U21003 : INV_X1 port map( I => n10561, ZN => n18770);
   U21004 : NAND2_X1 port map( A1 => n3003, A2 => n10561, ZN => n12682);
   U21009 : XOR2_X1 port map( A1 => n10252, A2 => n7792, Z => n10561);
   U21017 : XOR2_X1 port map( A1 => n6271, A2 => n11074, Z => n24202);
   U21057 : NOR2_X2 port map( A1 => n4228, A2 => n4227, ZN => n20073);
   U21058 : INV_X1 port map( I => n13057, ZN => n20849);
   U21063 : NAND2_X1 port map( A1 => n11319, A2 => n20850, ZN => n13057);
   U21081 : XOR2_X1 port map( A1 => n1651, A2 => n12813, Z => n24205);
   U21085 : XOR2_X1 port map( A1 => n24206, A2 => n4096, Z => n19778);
   U21087 : XOR2_X1 port map( A1 => n19319, A2 => n19320, Z => n24206);
   U21101 : OAI21_X1 port map( A1 => n4967, A2 => n16625, B => n25670, ZN => 
                           n16626);
   U21114 : XOR2_X1 port map( A1 => n13949, A2 => n27415, Z => n19538);
   U21128 : OR2_X1 port map( A1 => n3984, A2 => n18578, Z => n1786);
   U21130 : AND2_X1 port map( A1 => n1643, A2 => n24210, Z => n24439);
   U21132 : NAND3_X1 port map( A1 => n5573, A2 => n20155, A3 => n22830, ZN => 
                           n24210);
   U21142 : AND2_X1 port map( A1 => n4738, A2 => n24315, Z => n24464);
   U21149 : AND2_X1 port map( A1 => n11835, A2 => n12059, Z => n7735);
   U21166 : NAND2_X1 port map( A1 => n21474, A2 => n24212, ZN => n21475);
   U21180 : INV_X1 port map( I => n24213, ZN => n24212);
   U21196 : XOR2_X1 port map( A1 => n16374, A2 => n24220, Z => n2586);
   U21202 : XOR2_X1 port map( A1 => n1235, A2 => n16937, Z => n24220);
   U21207 : INV_X2 port map( I => n24223, ZN => n13509);
   U21214 : XOR2_X1 port map( A1 => n21158, A2 => n12320, Z => n12992);
   U21241 : XOR2_X1 port map( A1 => n24231, A2 => n20602, Z => Ciphertext(0));
   U21243 : NAND2_X2 port map( A1 => n24232, A2 => n15799, ZN => n11908);
   U21245 : INV_X1 port map( I => n21043, ZN => n9424);
   U21258 : NAND2_X1 port map( A1 => n24462, A2 => n24461, ZN => n33);
   U21275 : OR2_X1 port map( A1 => n2013, A2 => n10548, Z => n2012);
   U21307 : XOR2_X1 port map( A1 => n13937, A2 => n24241, Z => n13386);
   U21317 : XOR2_X1 port map( A1 => n24242, A2 => n13936, Z => n24241);
   U21319 : XNOR2_X1 port map( A1 => n16977, A2 => n566, ZN => n24264);
   U21320 : XOR2_X1 port map( A1 => n6327, A2 => n10683, Z => n24244);
   U21360 : NAND2_X2 port map( A1 => n24248, A2 => n5917, ZN => n6397);
   U21361 : OAI21_X2 port map( A1 => n6399, A2 => n7180, B => n5557, ZN => 
                           n24248);
   U21375 : XOR2_X1 port map( A1 => n24249, A2 => n6932, Z => n2276);
   U21382 : XOR2_X1 port map( A1 => n7257, A2 => n14616, Z => n24249);
   U21433 : NAND2_X1 port map( A1 => n21773, A2 => n21764, ZN => n15839);
   U21436 : XOR2_X1 port map( A1 => Plaintext(65), A2 => Key(65), Z => n569);
   U21444 : XOR2_X1 port map( A1 => n24253, A2 => n13200, Z => Ciphertext(35));
   U21445 : AOI22_X1 port map( A1 => n20754, A2 => n12417, B1 => n25334, B2 => 
                           n20753, ZN => n24253);
   U21458 : XOR2_X1 port map( A1 => n653, A2 => n9230, Z => n18740);
   U21483 : NAND2_X1 port map( A1 => n12066, A2 => n2093, ZN => n24259);
   U21502 : NAND2_X2 port map( A1 => n11415, A2 => n8575, ZN => n19143);
   U21504 : XOR2_X1 port map( A1 => n18311, A2 => n24263, Z => n7285);
   U21506 : XOR2_X1 port map( A1 => n13840, A2 => n14445, Z => n24263);
   U21534 : XOR2_X1 port map( A1 => n6288, A2 => n590, Z => n24266);
   U21536 : XOR2_X1 port map( A1 => n1372, A2 => n2691, Z => n9842);
   U21568 : XOR2_X1 port map( A1 => n18181, A2 => n9543, Z => n6306);
   U21570 : NAND3_X1 port map( A1 => n23441, A2 => n25724, A3 => n728, ZN => 
                           n3173);
   U21573 : XOR2_X1 port map( A1 => n24276, A2 => n20990, Z => Ciphertext(67));
   U21575 : XOR2_X1 port map( A1 => n24277, A2 => n20967, Z => Ciphertext(65));
   U21576 : OAI22_X1 port map( A1 => n15023, A2 => n21880, B1 => n20966, B2 => 
                           n705, ZN => n24277);
   U21578 : XOR2_X1 port map( A1 => n15303, A2 => n24279, Z => n664);
   U21580 : NAND2_X1 port map( A1 => n20980, A2 => n20979, ZN => n24280);
   U21581 : XOR2_X1 port map( A1 => n24281, A2 => n20771, Z => n9549);
   U21587 : NAND2_X2 port map( A1 => n14068, A2 => n14067, ZN => n16685);
   U21588 : XOR2_X1 port map( A1 => n24284, A2 => n2586, Z => n17345);
   U21589 : XOR2_X1 port map( A1 => n2585, A2 => n6707, Z => n24284);
   U21591 : XOR2_X1 port map( A1 => n16753, A2 => n24287, Z => n6513);
   U21593 : XOR2_X1 port map( A1 => n2220, A2 => n2219, Z => n5169);
   U21596 : INV_X2 port map( I => n24289, ZN => n24509);
   U21604 : XOR2_X1 port map( A1 => n22836, A2 => n24295, Z => n18224);
   U21607 : XOR2_X1 port map( A1 => n6867, A2 => n11022, Z => n12037);
   U21608 : NAND2_X2 port map( A1 => n5920, A2 => n4100, ZN => n11022);
   U21612 : OR2_X1 port map( A1 => n13662, A2 => n6800, Z => n3745);
   U21615 : NAND2_X2 port map( A1 => n24302, A2 => n4983, ZN => n5999);
   U21616 : AOI21_X1 port map( A1 => n25329, A2 => n20695, B => n27429, ZN => 
                           n20466);
   U21621 : INV_X2 port map( I => n24308, ZN => n17556);
   U21625 : XOR2_X1 port map( A1 => n16440, A2 => n13276, Z => n14117);
   U21627 : XOR2_X1 port map( A1 => n18258, A2 => n18047, Z => n18164);
   U21628 : XOR2_X1 port map( A1 => n16755, A2 => n17070, Z => n17008);
   U21631 : NOR2_X2 port map( A1 => n4828, A2 => n9105, ZN => n9052);
   U21633 : INV_X4 port map( I => n16531, ZN => n13964);
   U21637 : INV_X2 port map( I => n24311, ZN => n15989);
   U21638 : INV_X1 port map( I => n24321, ZN => n24320);
   U21639 : OAI21_X1 port map( A1 => n13142, A2 => n16280, B => n16050, ZN => 
                           n24321);
   U21640 : OAI21_X2 port map( A1 => n24322, A2 => n15714, B => n13188, ZN => 
                           n15713);
   U21641 : NOR2_X1 port map( A1 => n15688, A2 => n15689, ZN => n24322);
   U21642 : INV_X4 port map( I => n24324, ZN => n20237);
   U21644 : XOR2_X1 port map( A1 => n24325, A2 => n3868, Z => n21366);
   U21646 : OAI22_X2 port map( A1 => n13098, A2 => n20068, B1 => n20033, B2 => 
                           n20032, ZN => n14144);
   U21647 : XOR2_X1 port map( A1 => n24328, A2 => n15690, Z => n15688);
   U21648 : XOR2_X1 port map( A1 => n20509, A2 => n1506, Z => n24328);
   U21649 : INV_X2 port map( I => n24329, ZN => n10548);
   U21652 : XOR2_X1 port map( A1 => n884, A2 => n18234, Z => n8664);
   U21660 : OAI21_X2 port map( A1 => n7835, A2 => n2345, B => n2344, ZN => 
                           n12694);
   U21662 : NAND2_X1 port map( A1 => n16563, A2 => n16657, ZN => n16216);
   U21672 : XOR2_X1 port map( A1 => n94, A2 => n16958, Z => n2665);
   U21673 : OAI21_X2 port map( A1 => n24387, A2 => n17559, B => n24349, ZN => 
                           n11533);
   U21675 : INV_X1 port map( I => n5578, ZN => n6247);
   U21686 : XOR2_X1 port map( A1 => n24356, A2 => n21476, Z => Ciphertext(139))
                           ;
   U21687 : XOR2_X1 port map( A1 => n10670, A2 => n24358, Z => n11723);
   U21688 : XOR2_X1 port map( A1 => n28278, A2 => n1304, Z => n24358);
   U21691 : NAND3_X1 port map( A1 => n20795, A2 => n20797, A3 => n10050, ZN => 
                           n7526);
   U21692 : XOR2_X1 port map( A1 => n19504, A2 => n19335, Z => n19336);
   U21698 : OAI21_X2 port map( A1 => n4841, A2 => n16149, B => n5007, ZN => 
                           n14364);
   U21700 : XOR2_X1 port map( A1 => n3390, A2 => n20377, Z => n4896);
   U21701 : XOR2_X1 port map( A1 => n9598, A2 => n21154, Z => n13821);
   U21703 : NOR2_X2 port map( A1 => n13309, A2 => n7323, ZN => n17117);
   U21705 : NAND2_X2 port map( A1 => n10007, A2 => n2706, ZN => n15544);
   U21716 : OAI22_X2 port map( A1 => n8881, A2 => n13796, B1 => n4642, B2 => 
                           n14219, ZN => n10362);
   U21724 : XOR2_X1 port map( A1 => n12341, A2 => n12342, Z => n3363);
   U21730 : XOR2_X1 port map( A1 => n24399, A2 => n14630, Z => Ciphertext(24));
   U21732 : XOR2_X1 port map( A1 => n18082, A2 => n18083, Z => n2441);
   U21735 : XOR2_X1 port map( A1 => n23648, A2 => n21411, Z => n20348);
   U21737 : XOR2_X1 port map( A1 => n24415, A2 => n2463, Z => n2049);
   U21738 : XOR2_X1 port map( A1 => n21371, A2 => n20343, Z => n10950);
   U21740 : INV_X2 port map( I => n7108, ZN => n17349);
   U21741 : XOR2_X1 port map( A1 => n15237, A2 => n11502, Z => n18046);
   U21743 : INV_X2 port map( I => n24416, ZN => n12692);
   U21746 : INV_X2 port map( I => n24418, ZN => n1018);
   U21749 : INV_X2 port map( I => n19864, ZN => n19917);
   U21752 : XOR2_X1 port map( A1 => n12107, A2 => n7209, Z => n24427);
   U21753 : OAI21_X2 port map( A1 => n16179, A2 => n16178, B => n16177, ZN => 
                           n17147);
   U21755 : INV_X2 port map( I => n7745, ZN => n7338);
   U21756 : NAND2_X2 port map( A1 => n6214, A2 => n6213, ZN => n7745);
   U21759 : XOR2_X1 port map( A1 => n19347, A2 => n19184, Z => n1833);
   U21761 : OAI21_X1 port map( A1 => n21601, A2 => n21608, B => n24432, ZN => 
                           n5454);
   U21768 : INV_X2 port map( I => n616, ZN => n15189);
   U21771 : XNOR2_X1 port map( A1 => n18280, A2 => n1397, ZN => n257);
   U21773 : XOR2_X1 port map( A1 => n24438, A2 => n3816, Z => n20471);
   U21774 : XOR2_X1 port map( A1 => n21179, A2 => n3818, Z => n24438);
   U21775 : NAND2_X2 port map( A1 => n24439, A2 => n1642, ZN => n1638);
   U21780 : AND2_X1 port map( A1 => n12559, A2 => n12836, Z => n20992);
   U21786 : XOR2_X1 port map( A1 => n19324, A2 => n6528, Z => n19177);
   U21790 : NAND2_X1 port map( A1 => n15980, A2 => n16136, ZN => n14948);
   U21791 : NAND2_X1 port map( A1 => n6351, A2 => n28240, ZN => n24450);
   U21792 : INV_X2 port map( I => n24451, ZN => n24513);
   U21793 : XOR2_X1 port map( A1 => n7506, A2 => n7507, Z => n24451);
   U21797 : NOR2_X1 port map( A1 => n13194, A2 => n19941, ZN => n9310);
   U21799 : XOR2_X1 port map( A1 => n19321, A2 => n19322, Z => n4625);
   U21802 : XOR2_X1 port map( A1 => n19366, A2 => n5804, Z => n4708);
   U21806 : OAI22_X1 port map( A1 => n860, A2 => n20196, B1 => n14975, B2 => 
                           n20195, ZN => n20292);
   U21808 : NAND2_X2 port map( A1 => n14728, A2 => n16285, ZN => n16496);
   U21813 : NAND2_X1 port map( A1 => n24469, A2 => n24468, ZN => n20974);
   U21814 : NAND2_X1 port map( A1 => n7904, A2 => n24470, ZN => n24469);
   U21816 : OAI21_X2 port map( A1 => n24473, A2 => n24472, B => n18807, ZN => 
                           n3906);
   U21818 : NOR2_X1 port map( A1 => n9930, A2 => n845, ZN => n9929);
   U21824 : NAND3_X2 port map( A1 => n10977, A2 => n10976, A3 => n24476, ZN => 
                           n6699);
   U21825 : NAND3_X1 port map( A1 => n7970, A2 => n75, A3 => n27464, ZN => 
                           n24476);
   U21827 : XOR2_X1 port map( A1 => n17080, A2 => n21938, Z => n24477);
   U21829 : INV_X2 port map( I => n22744, ZN => n24478);
   U21831 : XOR2_X1 port map( A1 => n18181, A2 => n18284, Z => n15675);
   U21832 : XOR2_X1 port map( A1 => n6307, A2 => n6306, Z => n9761);
   U21833 : NAND2_X2 port map( A1 => n24480, A2 => n11125, ZN => n14906);
   U21835 : NAND2_X2 port map( A1 => n11316, A2 => n11313, ZN => n13853);
   U21840 : NOR2_X1 port map( A1 => n27460, A2 => n2777, ZN => n12810);
   U21842 : XOR2_X1 port map( A1 => n16804, A2 => n7097, Z => n24487);
   U21845 : XOR2_X1 port map( A1 => n24494, A2 => n12725, Z => n5525);
   U21852 : INV_X2 port map( I => n11968, ZN => n825);
   U21853 : NAND2_X2 port map( A1 => n5229, A2 => n8667, ZN => n11968);
   U21854 : OAI21_X1 port map( A1 => n11839, A2 => n14580, B => n24497, ZN => 
                           n18655);
   U21857 : XOR2_X1 port map( A1 => n12564, A2 => n24499, Z => n3527);
   U21859 : XOR2_X1 port map( A1 => n16537, A2 => n21897, Z => n1916);
   U21861 : NOR2_X2 port map( A1 => n17292, A2 => n14367, ZN => n24502);
   U21864 : NAND2_X1 port map( A1 => n1728, A2 => n1731, ZN => n1727);
   U21868 : XOR2_X1 port map( A1 => n5595, A2 => n18060, Z => n24506);
   U21872 : NOR3_X1 port map( A1 => n26615, A2 => n7370, A3 => n17196, ZN => 
                           n7778);
   U21873 : INV_X4 port map( I => n15699, ZN => n1030);
   U21876 : OR2_X1 port map( A1 => n13997, A2 => n3225, Z => n24514);
   U21884 : OR2_X2 port map( A1 => n6783, A2 => n6784, Z => n24528);
   U21886 : INV_X2 port map( I => n8564, ZN => n10549);
   U21887 : XNOR2_X1 port map( A1 => n7302, A2 => n14637, ZN => n24532);
   U21891 : XNOR2_X1 port map( A1 => n21309, A2 => n11701, ZN => n24536);
   U4503 : NAND2_X2 port map( A1 => n9393, A2 => n23104, ZN => n16078);
   U97 : NOR2_X2 port map( A1 => n21780, A2 => n8757, ZN => n22961);
   U852 : NAND2_X2 port map( A1 => n11374, A2 => n16574, ZN => n13604);
   U2476 : OAI21_X2 port map( A1 => n14320, A2 => n13721, B => n8999, ZN => 
                           n11374);
   U12775 : AND2_X2 port map( A1 => n7817, A2 => n18457, Z => n18600);
   U1186 : OAI22_X2 port map( A1 => n23758, A2 => n26244, B1 => n16587, B2 => 
                           n9725, ZN => n11776);
   U12035 : NAND2_X2 port map( A1 => n902, A2 => n5716, ZN => n2597);
   U2234 : AOI22_X2 port map( A1 => n5709, A2 => n25554, B1 => n25670, B2 => 
                           n907, ZN => n5708);
   U4209 : BUF_X4 port map( I => n20366, Z => n21624);
   U3130 : NAND2_X2 port map( A1 => n23424, A2 => n23423, ZN => n12895);
   U15488 : INV_X2 port map( I => n7987, ZN => n17981);
   U8705 : BUF_X2 port map( I => n21295, Z => n5519);
   U16796 : INV_X2 port map( I => n11369, ZN => n12614);
   U151 : BUF_X4 port map( I => n5841, Z => n3549);
   U1203 : INV_X4 port map( I => n23842, ZN => n14254);
   U12044 : AOI21_X1 port map( A1 => n13693, A2 => n11857, B => n17213, ZN => 
                           n2610);
   U2101 : OAI21_X2 port map( A1 => n21879, A2 => n13924, B => n6285, ZN => 
                           n6283);
   U8790 : INV_X2 port map( I => n14144, ZN => n1099);
   U13340 : NAND3_X2 port map( A1 => n18980, A2 => n19068, A3 => n22338, ZN => 
                           n15517);
   U12575 : OAI21_X2 port map( A1 => n26699, A2 => n8022, B => n4392, ZN => 
                           n18555);
   U12821 : NAND2_X2 port map( A1 => n23267, A2 => n26345, ZN => n13616);
   U4810 : OAI21_X2 port map( A1 => n13563, A2 => n2070, B => n23268, ZN => 
                           n23267);
   U972 : NOR2_X2 port map( A1 => n23987, A2 => n622, ZN => n7447);
   U433 : INV_X2 port map( I => n9002, ZN => n23818);
   U7388 : OAI21_X2 port map( A1 => n19190, A2 => n19191, B => n7995, ZN => 
                           n18990);
   U12404 : OAI21_X2 port map( A1 => n24460, A2 => n24459, B => n18463, ZN => 
                           n14100);
   U4740 : NOR2_X2 port map( A1 => n11196, A2 => n18605, ZN => n24459);
   U7971 : NAND2_X2 port map( A1 => n4164, A2 => n14177, ZN => n4163);
   U1716 : OAI21_X2 port map( A1 => n818, A2 => n4705, B => n8645, ZN => n8054)
                           ;
   U1555 : OAI21_X2 port map( A1 => n6320, A2 => n21387, B => n6319, ZN => 
                           n6318);
   U6181 : INV_X4 port map( I => n12502, ZN => n864);
   U3108 : OAI21_X2 port map( A1 => n13379, A2 => n23368, B => n13378, ZN => 
                           n11228);
   U633 : NAND2_X2 port map( A1 => n3889, A2 => n18677, ZN => n18999);
   U21839 : BUF_X4 port map( I => n7608, Z => n24485);
   U2413 : INV_X2 port map( I => n20405, ZN => n20642);
   U5595 : NOR2_X2 port map( A1 => n18583, A2 => n18586, ZN => n7741);
   U2866 : INV_X2 port map( I => n9761, ZN => n18586);
   U905 : NAND2_X2 port map( A1 => n16079, A2 => n10439, ZN => n11658);
   U466 : INV_X2 port map( I => n23905, ZN => n782);
   U20929 : INV_X2 port map( I => n14586, ZN => n24179);
   U799 : OAI21_X2 port map( A1 => n26658, A2 => n22285, B => n22594, ZN => 
                           n17611);
   U19834 : INV_X2 port map( I => n21323, ZN => n13791);
   U20301 : INV_X2 port map( I => n15359, ZN => n17534);
   U1457 : INV_X1 port map( I => n26993, ZN => n23163);
   U26 : INV_X2 port map( I => n12846, ZN => n21172);
   U1542 : INV_X2 port map( I => n14260, ZN => n5141);
   U18298 : AOI21_X2 port map( A1 => n25493, A2 => n7120, B => n12791, ZN => 
                           n12790);
   U940 : INV_X2 port map( I => n18101, ZN => n1202);
   U2134 : NAND2_X2 port map( A1 => n26643, A2 => n17894, ZN => n17701);
   U20223 : INV_X2 port map( I => n16066, ZN => n16312);
   U9229 : INV_X2 port map( I => n19260, ZN => n3243);
   U4004 : OAI22_X2 port map( A1 => n9521, A2 => n9520, B1 => n774, B2 => 
                           n13378, ZN => n9519);
   U4303 : INV_X2 port map( I => n5535, ZN => n10046);
   U2526 : INV_X2 port map( I => n4308, ZN => n14017);
   U669 : OAI21_X2 port map( A1 => n14308, A2 => n1016, B => n7446, ZN => 
                           n23745);
   U10472 : OAI21_X2 port map( A1 => n15906, A2 => n16347, B => n13705, ZN => 
                           n13704);
   U12480 : NOR2_X2 port map( A1 => n18101, A2 => n9344, ZN => n4461);
   U146 : INV_X2 port map( I => n9056, ZN => n9737);
   U3712 : NOR2_X2 port map( A1 => n25697, A2 => n17969, ZN => n6813);
   U2108 : NOR2_X2 port map( A1 => n19890, A2 => n8330, ZN => n23689);
   U1182 : INV_X2 port map( I => n16689, ZN => n16387);
   U305 : OAI21_X2 port map( A1 => n4069, A2 => n3920, B => n810, ZN => n22387)
                           ;
   U5920 : NOR3_X2 port map( A1 => n12894, A2 => n14752, A3 => n3317, ZN => 
                           n12893);
   U2381 : INV_X2 port map( I => n22429, ZN => n18124);
   U928 : NAND2_X2 port map( A1 => n23979, A2 => n787, ZN => n17332);
   U144 : NOR2_X2 port map( A1 => n21091, A2 => n25309, ZN => n1541);
   U1921 : INV_X2 port map( I => n17991, ZN => n4749);
   U1110 : INV_X2 port map( I => n19532, ZN => n2389);
   U5511 : NAND2_X2 port map( A1 => n22307, A2 => n7321, ZN => n17771);
   U15362 : INV_X2 port map( I => n17474, ZN => n23276);
   U2869 : OAI21_X2 port map( A1 => n6378, A2 => n24055, B => n19026, ZN => 
                           n19030);
   U851 : NOR2_X2 port map( A1 => n15061, A2 => n4281, ZN => n4280);
   U659 : INV_X2 port map( I => n10134, ZN => n8658);
   U8035 : OAI21_X2 port map( A1 => n9139, A2 => n16455, B => n16651, ZN => 
                           n5559);
   U3297 : NOR2_X2 port map( A1 => n6628, A2 => n5361, ZN => n22241);
   U10199 : INV_X2 port map( I => n3179, ZN => n2455);
   U945 : INV_X2 port map( I => n5095, ZN => n13731);
   U2113 : NAND3_X2 port map( A1 => n3773, A2 => n14456, A3 => n7300, ZN => 
                           n7483);
   U18299 : OAI21_X2 port map( A1 => n17842, A2 => n5238, B => n13051, ZN => 
                           n14474);
   U11185 : INV_X4 port map( I => n22602, ZN => n23002);
   U49 : OAI21_X2 port map( A1 => n12615, A2 => n15570, B => n15616, ZN => 
                           n23243);
   U1122 : AOI21_X2 port map( A1 => n2039, A2 => n1047, B => n24650, ZN => 
                           n6611);
   U867 : NAND2_X2 port map( A1 => n18101, A2 => n9344, ZN => n4306);
   U336 : NOR2_X2 port map( A1 => n4931, A2 => n7682, ZN => n19705);
   U3016 : INV_X2 port map( I => n21692, ZN => n10595);
   U204 : INV_X4 port map( I => n20237, ZN => n12177);
   U1060 : INV_X2 port map( I => n540, ZN => n23777);
   U5152 : INV_X2 port map( I => n13325, ZN => n13426);
   U1143 : OAI21_X2 port map( A1 => n26107, A2 => n16576, B => n16437, ZN => 
                           n2577);
   U7626 : NAND2_X2 port map( A1 => n11858, A2 => n1215, ZN => n17858);
   U9141 : NOR2_X2 port map( A1 => n19890, A2 => n12393, ZN => n4069);
   U4531 : INV_X2 port map( I => n8089, ZN => n24500);
   U17549 : AOI21_X2 port map( A1 => n250, A2 => n16273, B => n8873, ZN => 
                           n12605);
   U2971 : NOR2_X2 port map( A1 => n10464, A2 => n17229, ZN => n23066);
   U332 : INV_X2 port map( I => n12941, ZN => n1115);
   U4407 : NOR2_X2 port map( A1 => n16283, A2 => n21787, ZN => n11290);
   U19789 : INV_X2 port map( I => n15958, ZN => n13677);
   U319 : INV_X2 port map( I => n14039, ZN => n20110);
   U1303 : BUF_X2 port map( I => n7065, Z => n23198);
   U6160 : NAND2_X2 port map( A1 => n204, A2 => n4810, ZN => n14895);
   U367 : INV_X2 port map( I => n2941, ZN => n15457);
   U1698 : AOI22_X2 port map( A1 => n16276, A2 => n14786, B1 => n22319, B2 => 
                           n8812, ZN => n1794);
   U4519 : NAND2_X2 port map( A1 => n9116, A2 => n16651, ZN => n16456);
   U1485 : NOR2_X2 port map( A1 => n11743, A2 => n23802, ZN => n13770);
   U1907 : AOI21_X2 port map( A1 => n18541, A2 => n2012, B => n18543, ZN => 
                           n10278);
   U3518 : NAND2_X2 port map( A1 => n10414, A2 => n14396, ZN => n3283);
   U953 : INV_X2 port map( I => n27240, ZN => n7226);
   U2630 : NAND2_X2 port map( A1 => n24283, A2 => n7379, ZN => n20244);
   U661 : NAND2_X2 port map( A1 => n21790, A2 => n27871, ZN => n18764);
   U410 : NAND2_X2 port map( A1 => n7523, A2 => n7522, ZN => n19281);
   U139 : INV_X2 port map( I => n15512, ZN => n21713);
   U2729 : INV_X2 port map( I => n8656, ZN => n10126);
   U14172 : INV_X2 port map( I => n22991, ZN => n9223);
   U318 : NAND2_X2 port map( A1 => n28357, A2 => n19872, ZN => n22515);
   U2010 : OAI21_X2 port map( A1 => n27630, A2 => n961, B => n8723, ZN => n2833
                           );
   U277 : NAND2_X2 port map( A1 => n19709, A2 => n6394, ZN => n1606);
   U16271 : INV_X4 port map( I => n4410, ZN => n1017);
   U3795 : INV_X4 port map( I => n6617, ZN => n5081);
   U12915 : INV_X2 port map( I => n20154, ZN => n6254);
   U20160 : AOI22_X2 port map( A1 => n16189, A2 => n16188, B1 => n16298, B2 => 
                           n11568, ZN => n14832);
   U16318 : NAND2_X2 port map( A1 => n781, A2 => n25592, ZN => n8006);
   U638 : NOR2_X2 port map( A1 => n7799, A2 => n18463, ZN => n12969);
   U5013 : INV_X2 port map( I => n809, ZN => n11631);
   U2856 : AOI21_X2 port map( A1 => n2794, A2 => n2793, B => n23748, ZN => 
                           n2792);
   U7101 : NAND3_X2 port map( A1 => n5280, A2 => n10227, A3 => n10221, ZN => 
                           n10226);
   U1213 : INV_X2 port map( I => n16225, ZN => n14786);
   U2960 : NOR2_X2 port map( A1 => n25724, A2 => n17906, ZN => n5866);
   U340 : INV_X4 port map( I => n9584, ZN => n9701);
   U3161 : BUF_X2 port map( I => n19720, Z => n24392);
   U8760 : INV_X2 port map( I => n9918, ZN => n1097);
   U3177 : NAND2_X2 port map( A1 => n9971, A2 => n18942, ZN => n1495);
   U2312 : NAND2_X2 port map( A1 => n5489, A2 => n17510, ZN => n6199);
   U6847 : BUF_X4 port map( I => n11722, Z => n8926);
   U17366 : NAND2_X2 port map( A1 => n8191, A2 => n21969, ZN => n23610);
   U14042 : NOR2_X1 port map( A1 => n23070, A2 => n4337, ZN => n22959);
   U1671 : AND2_X2 port map( A1 => n18002, A2 => n18003, Z => n12104);
   U298 : INV_X2 port map( I => n19917, ZN => n12145);
   U1177 : NAND2_X2 port map( A1 => n9725, A2 => n23907, ZN => n16421);
   U7816 : AOI21_X2 port map( A1 => n7694, A2 => n13766, B => n790, ZN => n7693
                           );
   U3497 : INV_X2 port map( I => n22529, ZN => n906);
   U630 : INV_X2 port map( I => n25966, ZN => n9480);
   U4851 : NAND2_X2 port map( A1 => n133, A2 => n18997, ZN => n1961);
   U1181 : INV_X2 port map( I => n16517, ZN => n22570);
   U20506 : OAI21_X2 port map( A1 => n15857, A2 => n14108, B => n1258, ZN => 
                           n15858);
   U1243 : NOR3_X2 port map( A1 => n13406, A2 => n799, A3 => n7398, ZN => 
                           n22333);
   U1892 : AOI21_X2 port map( A1 => n16363, A2 => n27160, B => n5670, ZN => 
                           n5669);
   U18569 : INV_X2 port map( I => n18161, ZN => n10907);
   U12712 : INV_X2 port map( I => n16652, ZN => n24302);
   U1692 : BUF_X4 port map( I => n21055, Z => n12066);
   U979 : INV_X4 port map( I => n23023, ZN => n11182);
   U755 : INV_X2 port map( I => n10536, ZN => n1016);
   U512 : INV_X2 port map( I => n6999, ZN => n18943);
   U20194 : INV_X2 port map( I => n10730, ZN => n21099);
   U774 : INV_X2 port map( I => n10246, ZN => n17492);
   U2210 : BUF_X4 port map( I => n17745, Z => n7358);
   U14616 : NAND3_X2 port map( A1 => n12485, A2 => n25733, A3 => n17524, ZN => 
                           n11170);
   U2913 : OAI21_X2 port map( A1 => n10437, A2 => n18588, B => n18546, ZN => 
                           n10014);
   U13041 : INV_X2 port map( I => n19928, ZN => n15048);
   U6557 : NAND2_X2 port map( A1 => n13070, A2 => n1036, ZN => n7846);
   U7782 : NAND2_X2 port map( A1 => n17723, A2 => n25697, ZN => n6799);
   U8515 : NAND2_X1 port map( A1 => n6485, A2 => n21083, ZN => n6881);
   U714 : NAND2_X2 port map( A1 => n8269, A2 => n2445, ZN => n22912);
   U7254 : NAND2_X2 port map( A1 => n9646, A2 => n113, ZN => n6234);
   U1196 : NAND2_X2 port map( A1 => n16600, A2 => n5557, ZN => n24182);
   U19973 : INV_X4 port map( I => n14178, ZN => n16013);
   U3404 : INV_X2 port map( I => n26665, ZN => n16144);
   U1965 : NOR2_X2 port map( A1 => n9593, A2 => n17487, ZN => n13997);
   U16079 : NAND2_X2 port map( A1 => n15620, A2 => n15621, ZN => n11155);
   U6845 : BUF_X4 port map( I => n15889, Z => n16086);
   U6725 : INV_X2 port map( I => n16571, ZN => n1053);
   U12669 : OAI21_X2 port map( A1 => n361, A2 => n851, B => n21689, ZN => n2804
                           );
   U18746 : AOI21_X2 port map( A1 => n2147, A2 => n24485, B => n23837, ZN => 
                           n23836);
   U5708 : INV_X4 port map( I => n24517, ZN => n1036);
   U333 : OR2_X2 port map( A1 => n22978, A2 => n25308, Z => n19936);
   U14445 : OAI21_X2 port map( A1 => n15828, A2 => n21773, B => n15358, ZN => 
                           n5073);
   U955 : NAND2_X2 port map( A1 => n21901, A2 => n22646, ZN => n17971);
   U19045 : INV_X2 port map( I => n16516, ZN => n16558);
   U14938 : NOR2_X2 port map( A1 => n454, A2 => n951, ZN => n21506);
   U5713 : INV_X4 port map( I => n14126, ZN => n898);
   U1923 : NAND3_X2 port map( A1 => n14184, A2 => n20415, A3 => n14185, ZN => 
                           n14258);
   U6728 : INV_X2 port map( I => n16433, ZN => n7430);
   U2330 : OAI22_X2 port map( A1 => n18145, A2 => n18586, B1 => n15137, B2 => 
                           n18583, ZN => n18814);
   U16268 : NAND2_X2 port map( A1 => n1087, A2 => n8050, ZN => n21026);
   U7891 : NAND2_X2 port map( A1 => n832, A2 => n11113, ZN => n17161);
   U4277 : INV_X2 port map( I => n7966, ZN => n10556);
   U19205 : OAI21_X2 port map( A1 => n1263, A2 => n795, B => n9223, ZN => 
                           n16108);
   U17094 : NAND2_X2 port map( A1 => n26343, A2 => n12692, ZN => n17524);
   U18060 : INV_X2 port map( I => n13421, ZN => n17281);
   U8138 : OAI21_X2 port map( A1 => n12535, A2 => n12536, B => n24641, ZN => 
                           n9433);
   U2682 : NOR2_X2 port map( A1 => n669, A2 => n11114, ZN => n19747);
   U15942 : NAND2_X1 port map( A1 => n23362, A2 => n15631, ZN => n16377);
   U98 : NAND2_X2 port map( A1 => n12310, A2 => n28314, ZN => n11207);
   U6434 : NAND2_X2 port map( A1 => n3929, A2 => n17726, ZN => n17657);
   U1092 : BUF_X4 port map( I => n17446, Z => n21785);
   U930 : INV_X2 port map( I => n6886, ZN => n3735);
   U3181 : INV_X1 port map( I => n17694, ZN => n17905);
   U11291 : INV_X4 port map( I => n1879, ZN => n8512);
   U4437 : OAI21_X2 port map( A1 => n16148, A2 => n4926, B => n8926, ZN => 
                           n9258);
   U329 : OR2_X2 port map( A1 => n25354, A2 => n9147, Z => n19671);
   U710 : INV_X2 port map( I => n8109, ZN => n22325);
   U18853 : INV_X2 port map( I => n20043, ZN => n20181);
   U3359 : AOI21_X2 port map( A1 => n22163, A2 => n22162, B => n9799, ZN => 
                           n9797);
   U21764 : AOI21_X2 port map( A1 => n16014, A2 => n16013, B => n12272, ZN => 
                           n16015);
   U2506 : CLKBUF_X4 port map( I => n16131, Z => n14386);
   U15691 : OAI21_X2 port map( A1 => n14804, A2 => n12964, B => n28118, ZN => 
                           n6604);
   U13022 : NAND2_X2 port map( A1 => n7609, A2 => n997, ZN => n24361);
   U17967 : NAND3_X1 port map( A1 => n14690, A2 => n971, A3 => n14319, ZN => 
                           n14689);
   U7095 : OAI22_X2 port map( A1 => n13301, A2 => n25254, B1 => n21932, B2 => 
                           n22398, ZN => n5388);
   U545 : AOI22_X2 port map( A1 => n19008, A2 => n18953, B1 => n6089, B2 => 
                           n18426, ZN => n18923);
   U104 : INV_X4 port map( I => n10610, ZN => n953);
   U1804 : OAI21_X2 port map( A1 => n21626, A2 => n21624, B => n21623, ZN => 
                           n6568);
   U10660 : CLKBUF_X2 port map( I => Key(157), Z => n14630);
   U17900 : OAI21_X2 port map( A1 => n17482, A2 => n25733, B => n17483, ZN => 
                           n11771);
   U9163 : BUF_X2 port map( I => n19891, Z => n6865);
   U1132 : NOR3_X2 port map( A1 => n8530, A2 => n24089, A3 => n22838, ZN => 
                           n5670);
   U1695 : INV_X2 port map( I => n16619, ZN => n5062);
   U14623 : NAND3_X2 port map( A1 => n19668, A2 => n19669, A3 => n28425, ZN => 
                           n5234);
   U1955 : NAND3_X2 port map( A1 => n24674, A2 => n8256, A3 => n23968, ZN => 
                           n8152);
   U16011 : NAND2_X2 port map( A1 => n14103, A2 => n26343, ZN => n7073);
   U3069 : NAND2_X2 port map( A1 => n6097, A2 => n6096, ZN => n24208);
   U5574 : OR2_X1 port map( A1 => n27528, A2 => n15454, Z => n21933);
   U5236 : INV_X2 port map( I => n7817, ZN => n18473);
   U1075 : OAI21_X2 port map( A1 => n11416, A2 => n10545, B => n3454, ZN => 
                           n11415);
   U4525 : NOR2_X2 port map( A1 => n718, A2 => n11908, ZN => n10643);
   U246 : NOR2_X2 port map( A1 => n19835, A2 => n967, ZN => n4929);
   U1087 : INV_X2 port map( I => n2564, ZN => n10908);
   U224 : NAND3_X2 port map( A1 => n26730, A2 => n24534, A3 => n4710, ZN => 
                           n12872);
   U5183 : OAI21_X2 port map( A1 => n21013, A2 => n13600, B => n21175, ZN => 
                           n21014);
   U12390 : AOI21_X2 port map( A1 => n18641, A2 => n18746, B => n14362, ZN => 
                           n11637);
   U3749 : OR2_X2 port map( A1 => n25305, A2 => n24228, Z => n21813);
   U8346 : BUF_X2 port map( I => Key(45), Z => n20621);
   U484 : NAND2_X1 port map( A1 => n11890, A2 => n3902, ZN => n18540);
   U7476 : AOI21_X2 port map( A1 => n4389, A2 => n18489, B => n5037, ZN => 
                           n4388);
   U3213 : NOR2_X2 port map( A1 => n24611, A2 => n10649, ZN => n24104);
   U2909 : INV_X2 port map( I => n5759, ZN => n22218);
   U9903 : INV_X4 port map( I => n2895, ZN => n6076);
   U4417 : NOR2_X2 port map( A1 => n6861, A2 => n7326, ZN => n19848);
   U4120 : BUF_X4 port map( I => n8155, Z => n22396);
   U9945 : NOR2_X1 port map( A1 => n11945, A2 => n9410, ZN => n10257);
   U282 : OAI21_X2 port map( A1 => n24364, A2 => n11317, B => n27916, ZN => 
                           n11316);
   U2031 : NAND2_X2 port map( A1 => n14912, A2 => n13757, ZN => n19013);
   U317 : NAND2_X2 port map( A1 => n19839, A2 => n22422, ZN => n19621);
   U5374 : BUF_X4 port map( I => n6508, Z => n1617);
   U8827 : NAND2_X2 port map( A1 => n10399, A2 => n28071, ZN => n10287);
   U3881 : OAI21_X2 port map( A1 => n18904, A2 => n18943, B => n13346, ZN => 
                           n22954);
   U11712 : AOI21_X2 port map( A1 => n14888, A2 => n16200, B => n8241, ZN => 
                           n3854);
   U8533 : NAND2_X1 port map( A1 => n17254, A2 => n4536, ZN => n22263);
   U11924 : OAI21_X2 port map( A1 => n19921, A2 => n19748, B => n2492, ZN => 
                           n4774);
   U4828 : INV_X2 port map( I => n2391, ZN => n12026);
   U11522 : NOR2_X2 port map( A1 => n9179, A2 => n732, ZN => n8767);
   U2659 : INV_X4 port map( I => n819, ZN => n875);
   U733 : INV_X2 port map( I => n5523, ZN => n10569);
   U2999 : AOI22_X2 port map( A1 => n8980, A2 => n10604, B1 => n6909, B2 => 
                           n10636, ZN => n350);
   U2136 : OAI21_X2 port map( A1 => n357, A2 => n18590, B => n7446, ZN => n5342
                           );
   U14664 : INV_X2 port map( I => n5264, ZN => n10603);
   U21794 : OAI21_X2 port map( A1 => n806, A2 => n20174, B => n24554, ZN => 
                           n7418);
   U4339 : INV_X1 port map( I => n15891, ZN => n16350);
   U10661 : BUF_X2 port map( I => Key(150), Z => n14616);
   U8111 : NAND2_X2 port map( A1 => n124, A2 => n16649, ZN => n16393);
   U2028 : NOR2_X2 port map( A1 => n1835, A2 => n20234, ZN => n22921);
   U18912 : NAND2_X2 port map( A1 => n23236, A2 => n14562, ZN => n14259);
   U761 : INV_X2 port map( I => n24379, ZN => n1440);
   U2934 : INV_X2 port map( I => n5473, ZN => n12498);
   U15870 : NAND2_X1 port map( A1 => n23339, A2 => n24299, ZN => n23338);
   U4757 : INV_X2 port map( I => n18341, ZN => n18507);
   U7387 : OAI21_X2 port map( A1 => n12577, A2 => n12576, B => n26395, ZN => 
                           n3865);
   U7457 : NOR2_X2 port map( A1 => n7084, A2 => n12781, ZN => n12577);
   U18556 : INV_X1 port map( I => n18772, ZN => n18623);
   U4411 : OAI21_X2 port map( A1 => n10357, A2 => n5706, B => n1115, ZN => 
                           n6548);
   U20751 : OAI21_X2 port map( A1 => n309, A2 => n24162, B => n21824, ZN => 
                           n17252);
   U2048 : OR3_X1 port map( A1 => n20064, A2 => n9525, A3 => n22398, Z => 
                           n22517);
   U582 : INV_X2 port map( I => n28370, ZN => n2098);
   U18996 : NOR2_X2 port map( A1 => n18627, A2 => n235, ZN => n18626);
   U1679 : NOR2_X2 port map( A1 => n5370, A2 => n8883, ZN => n14468);
   U6539 : AOI22_X2 port map( A1 => n7621, A2 => n17181, B1 => n7620, B2 => 
                           n17565, ZN => n7619);
   U4311 : INV_X4 port map( I => n11238, ZN => n12949);
   U2505 : INV_X1 port map( I => n17745, ZN => n1216);
   U14137 : INV_X4 port map( I => n4634, ZN => n15787);
   U5724 : NOR3_X2 port map( A1 => n16574, A2 => n7378, A3 => n22660, ZN => 
                           n15302);
   U421 : NAND2_X2 port map( A1 => n13354, A2 => n19274, ZN => n13778);
   U12244 : OAI22_X2 port map( A1 => n18860, A2 => n2798, B1 => n14222, B2 => 
                           n18861, ZN => n15424);
   U14875 : AOI21_X2 port map( A1 => n14179, A2 => n9264, B => n9449, ZN => 
                           n23143);
   U14238 : INV_X4 port map( I => n15787, ZN => n13742);
   U10883 : NOR2_X2 port map( A1 => n12151, A2 => n12152, ZN => n23798);
   U439 : OAI21_X2 port map( A1 => n18931, A2 => n3014, B => n3032, ZN => n3031
                           );
   U228 : INV_X2 port map( I => n14663, ZN => n23408);
   U166 : BUF_X2 port map( I => n8366, Z => n446);
   U13078 : INV_X2 port map( I => n16988, ZN => n1235);
   U14511 : NAND2_X1 port map( A1 => n11651, A2 => n23044, ZN => n23043);
   U14971 : NAND2_X2 port map( A1 => n5830, A2 => n5762, ZN => n5761);
   U2160 : NAND3_X2 port map( A1 => n2390, A2 => n12026, A3 => n24580, ZN => 
                           n16452);
   U7752 : NOR2_X2 port map( A1 => n14230, A2 => n26610, ZN => n3234);
   U12813 : INV_X2 port map( I => n20516, ZN => n22785);
   U6896 : NOR2_X2 port map( A1 => n24307, A2 => n7991, ZN => n11781);
   U18995 : NAND2_X2 port map( A1 => n18627, A2 => n235, ZN => n11711);
   U853 : NOR3_X2 port map( A1 => n23979, A2 => n787, A3 => n11182, ZN => 
                           n22104);
   U2519 : BUF_X2 port map( I => n16325, Z => n14559);
   U1599 : INV_X1 port map( I => n4883, ZN => n18448);
   U8988 : AOI21_X2 port map( A1 => n19269, A2 => n5332, B => n11836, ZN => 
                           n8412);
   U2924 : NOR2_X2 port map( A1 => n24155, A2 => n24156, ZN => n21986);
   U4631 : OAI21_X2 port map( A1 => n7194, A2 => n10911, B => n17415, ZN => 
                           n5281);
   U13169 : AOI21_X2 port map( A1 => n4212, A2 => n1444, B => n1443, ZN => 
                           n1442);
   U1168 : OAI21_X2 port map( A1 => n21825, A2 => n26277, B => n28106, ZN => 
                           n273);
   U19176 : INV_X2 port map( I => n21035, ZN => n21050);
   U4692 : OAI21_X1 port map( A1 => n2955, A2 => n4914, B => n2953, ZN => n2956
                           );
   U6341 : NAND3_X1 port map( A1 => n2133, A2 => n18727, A3 => n18728, ZN => 
                           n2132);
   U452 : INV_X2 port map( I => n3030, ZN => n3014);
   U2641 : CLKBUF_X2 port map( I => n8118, Z => n260);
   U7844 : NAND3_X1 port map( A1 => n22279, A2 => n23032, A3 => n6722, ZN => 
                           n22192);
   U15982 : NAND3_X2 port map( A1 => n16589, A2 => n16588, A3 => n9725, ZN => 
                           n16590);
   U1760 : INV_X4 port map( I => n10613, ZN => n1119);
   U2744 : AND2_X1 port map( A1 => n22345, A2 => n15502, Z => n7445);
   U2227 : INV_X2 port map( I => n16494, ZN => n910);
   U1041 : NOR2_X2 port map( A1 => n627, A2 => n5447, ZN => n6214);
   U2379 : BUF_X4 port map( I => n13759, Z => n6264);
   U16369 : OR2_X1 port map( A1 => n12022, A2 => n7298, Z => n2524);
   U9055 : NAND2_X1 port map( A1 => n13760, A2 => n19360, ZN => n13736);
   U3903 : INV_X4 port map( I => n14654, ZN => n987);
   U18309 : NOR2_X2 port map( A1 => n4063, A2 => n26533, ZN => n13723);
   U171 : AND2_X2 port map( A1 => n9371, A2 => n7086, Z => n22756);
   U6502 : NAND2_X2 port map( A1 => n4814, A2 => n17927, ZN => n17640);
   U7563 : NAND2_X2 port map( A1 => n25499, A2 => n10537, ZN => n1974);
   U10685 : BUF_X2 port map( I => Key(63), Z => n14610);
   U911 : NOR2_X2 port map( A1 => n17332, A2 => n9905, ZN => n5447);
   U444 : AND2_X2 port map( A1 => n8043, A2 => n8044, Z => n21758);
   U9752 : NAND2_X2 port map( A1 => n8382, A2 => n17981, ZN => n8381);
   U2651 : BUF_X2 port map( I => n10144, Z => n265);
   U2719 : OAI22_X2 port map( A1 => n11789, A2 => n25710, B1 => n1110, B2 => 
                           n25254, ZN => n21963);
   U316 : INV_X2 port map( I => n7582, ZN => n19914);
   U8169 : NOR2_X2 port map( A1 => n13362, A2 => n15931, ZN => n8088);
   U4821 : NOR2_X2 port map( A1 => n26262, A2 => n8084, ZN => n16696);
   U7654 : NOR2_X1 port map( A1 => n14599, A2 => n17677, ZN => n2100);
   U9310 : NAND2_X1 port map( A1 => n9409, A2 => n9408, ZN => n6417);
   U12776 : AOI22_X2 port map( A1 => n2832, A2 => n183, B1 => n2833, B2 => 
                           n25722, ZN => n12468);
   U2717 : NAND2_X2 port map( A1 => n9725, A2 => n14879, ZN => n16360);
   U18039 : NOR2_X2 port map( A1 => n6316, A2 => n6315, ZN => n15807);
   U12276 : BUF_X4 port map( I => n10856, Z => n9105);
   U7130 : INV_X1 port map( I => n13759, ZN => n14740);
   U9201 : INV_X1 port map( I => n19407, ZN => n8678);
   U5178 : BUF_X4 port map( I => n12612, Z => n7302);
   U2511 : OAI21_X2 port map( A1 => n13215, A2 => n13214, B => n16175, ZN => 
                           n14803);
   U5122 : NOR2_X2 port map( A1 => n8864, A2 => n20474, ZN => n13100);
   U10356 : BUF_X4 port map( I => n16646, Z => n5244);
   U4584 : INV_X2 port map( I => n10580, ZN => n17292);
   U5768 : NAND3_X2 port map( A1 => n2343, A2 => n2342, A3 => n796, ZN => n2344
                           );
   U13595 : NOR2_X2 port map( A1 => n1499, A2 => n1500, ZN => n22996);
   U3007 : NAND2_X2 port map( A1 => n23781, A2 => n16311, ZN => n16494);
   U10659 : BUF_X2 port map( I => Key(89), Z => n14640);
   U5806 : BUF_X2 port map( I => n15188, Z => n1270);
   U18263 : NAND2_X1 port map( A1 => n15297, A2 => n24952, ZN => n15296);
   U18264 : OAI21_X1 port map( A1 => n25415, A2 => n28400, B => n15298, ZN => 
                           n15297);
   U6143 : NOR2_X2 port map( A1 => n8836, A2 => n978, ZN => n8835);
   U2188 : NAND2_X2 port map( A1 => n2891, A2 => n1133, ZN => n8836);
   U17724 : NOR2_X1 port map( A1 => n12397, A2 => n23974, ZN => n6483);
   U7823 : AOI21_X2 port map( A1 => n16996, A2 => n1631, B => n9481, ZN => 
                           n1630);
   U20517 : INV_X1 port map( I => n16130, ZN => n15873);
   U2931 : NOR2_X2 port map( A1 => n22492, A2 => n21888, ZN => n23616);
   U1351 : AOI21_X2 port map( A1 => n5760, A2 => n24315, B => n2545, ZN => 
                           n5182);
   U14153 : INV_X4 port map( I => n18639, ZN => n22977);
   U12961 : INV_X2 port map( I => n6076, ZN => n3346);
   U3589 : NOR2_X2 port map( A1 => n11072, A2 => n7703, ZN => n5068);
   U5551 : BUF_X4 port map( I => n20153, Z => n7618);
   U6856 : BUF_X2 port map( I => n10573, Z => n7235);
   U4495 : OAI21_X2 port map( A1 => n23530, A2 => n23531, B => n28257, ZN => 
                           n3380);
   U2507 : OAI22_X2 port map( A1 => n9168, A2 => n27494, B1 => n20314, B2 => 
                           n20244, ZN => n6421);
   U1024 : INV_X2 port map( I => n19782, ZN => n15028);
   U5196 : INV_X2 port map( I => n2484, ZN => n19046);
   U3381 : OAI21_X2 port map( A1 => n16308, A2 => n16309, B => n1270, ZN => 
                           n23781);
   U5120 : OAI21_X2 port map( A1 => n13924, A2 => n20288, B => n20430, ZN => 
                           n20289);
   U382 : NAND3_X2 port map( A1 => n2726, A2 => n11696, A3 => n1152, ZN => 
                           n6242);
   U12327 : NOR2_X2 port map( A1 => n21734, A2 => n6281, ZN => n21738);
   U985 : AOI21_X2 port map( A1 => n17195, A2 => n7363, B => n7778, ZN => n7783
                           );
   U981 : AOI21_X2 port map( A1 => n22979, A2 => n13035, B => n17432, ZN => 
                           n5512);
   U8207 : NAND2_X2 port map( A1 => n13783, A2 => n16027, ZN => n13782);
   U74 : INV_X2 port map( I => n21545, ZN => n21543);
   U4609 : OAI21_X2 port map( A1 => n1207, A2 => n13350, B => n28457, ZN => 
                           n1568);
   U18246 : AOI21_X2 port map( A1 => n16708, A2 => n16709, B => n1253, ZN => 
                           n16710);
   U1228 : OAI22_X2 port map( A1 => n10697, A2 => n22975, B1 => n16351, B2 => 
                           n16086, ZN => n24232);
   U10923 : NAND3_X1 port map( A1 => n25679, A2 => n1512, A3 => n4914, ZN => 
                           n6991);
   U1833 : NAND2_X2 port map( A1 => n242, A2 => n899, ZN => n17577);
   U4572 : BUF_X4 port map( I => n11354, Z => n9762);
   U17590 : NOR2_X2 port map( A1 => n14141, A2 => n26673, ZN => n23651);
   U3291 : AOI21_X2 port map( A1 => n17997, A2 => n17998, B => n14826, ZN => 
                           n22439);
   U2515 : NAND2_X2 port map( A1 => n16524, A2 => n3537, ZN => n2693);
   U18841 : AOI21_X2 port map( A1 => n13040, A2 => n12423, B => n26108, ZN => 
                           n12537);
   U6182 : INV_X4 port map( I => n9701, ZN => n9645);
   U9070 : NAND2_X1 port map( A1 => n13666, A2 => n19926, ZN => n14240);
   U21747 : BUF_X4 port map( I => n14997, Z => n24419);
   U6114 : NAND3_X2 port map( A1 => n3989, A2 => n26528, A3 => n3988, ZN => 
                           n3277);
   U3854 : OAI21_X2 port map( A1 => n2993, A2 => n23752, B => n19165, ZN => 
                           n10240);
   U4259 : OAI22_X2 port map( A1 => n4554, A2 => n7759, B1 => n4553, B2 => 
                           n26835, ZN => n22958);
   U800 : OAI21_X2 port map( A1 => n1021, A2 => n23811, B => n23810, ZN => 
                           n15664);
   U2647 : INV_X4 port map( I => n20171, ZN => n4782);
   U5802 : OAI21_X1 port map( A1 => n1853, A2 => n944, B => n1851, ZN => n23536
                           );
   U13199 : NOR2_X1 port map( A1 => n4014, A2 => n9344, ZN => n4013);
   U3345 : NOR2_X1 port map( A1 => n26989, A2 => n17493, ZN => n22164);
   U12081 : INV_X2 port map( I => n21636, ZN => n7009);
   U6770 : NAND2_X2 port map( A1 => n10793, A2 => n10792, ZN => n10791);
   U2496 : NAND2_X2 port map( A1 => n2120, A2 => n14649, ZN => n8384);
   U10317 : INV_X2 port map( I => n12974, ZN => n16055);
   U18579 : NOR3_X2 port map( A1 => n27171, A2 => n17881, A3 => n23806, ZN => 
                           n5370);
   U4121 : OAI21_X1 port map( A1 => n6589, A2 => n20744, B => n20749, ZN => 
                           n6053);
   U2995 : AOI22_X2 port map( A1 => n21891, A2 => n742, B1 => n741, B2 => 
                           n16361, ZN => n16362);
   U819 : NOR2_X2 port map( A1 => n13608, A2 => n4998, ZN => n4479);
   U6842 : AND2_X2 port map( A1 => n333, A2 => n15905, Z => n11693);
   U4682 : NOR2_X2 port map( A1 => n1213, A2 => n728, ZN => n9078);
   U15955 : NAND3_X1 port map( A1 => n15542, A2 => n20121, A3 => n23401, ZN => 
                           n7012);
   U68 : OAI21_X2 port map( A1 => n20729, A2 => n20731, B => n25145, ZN => 
                           n20734);
   U10381 : AOI22_X2 port map( A1 => n15966, A2 => n16348, B1 => n15969, B2 => 
                           n15968, ZN => n2660);
   U9178 : NAND3_X1 port map( A1 => n20678, A2 => n20679, A3 => n26557, ZN => 
                           n22343);
   U13174 : INV_X2 port map( I => n10830, ZN => n4532);
   U2942 : OAI21_X2 port map( A1 => n1870, A2 => n12677, B => n12676, ZN => 
                           n23833);
   U8769 : INV_X2 port map( I => n13271, ZN => n20056);
   U10242 : AOI21_X2 port map( A1 => n15419, A2 => n15418, B => n910, ZN => 
                           n12607);
   U1597 : INV_X2 port map( I => n18776, ZN => n4161);
   U17199 : NOR2_X1 port map( A1 => n9258, A2 => n9259, ZN => n8513);
   U21567 : OAI21_X1 port map( A1 => n10636, A2 => n22747, B => n21717, ZN => 
                           n21718);
   U1248 : NAND2_X2 port map( A1 => n8398, A2 => n4926, ZN => n15959);
   U5789 : NOR2_X2 port map( A1 => n8620, A2 => n14520, ZN => n13776);
   U938 : NAND2_X2 port map( A1 => n12507, A2 => n16279, ZN => n13142);
   U1386 : INV_X4 port map( I => n8926, ZN => n8398);
   U7547 : NOR2_X1 port map( A1 => n5705, A2 => n14417, ZN => n4786);
   U331 : INV_X1 port map( I => n19280, ZN => n2223);
   U16272 : AND2_X2 port map( A1 => n16379, A2 => n16378, Z => n7323);
   U3606 : INV_X2 port map( I => n16166, ZN => n16279);
   U16380 : AND2_X2 port map( A1 => n7464, A2 => n7463, Z => n10690);
   U121 : INV_X2 port map( I => n9756, ZN => n10031);
   U1509 : OR2_X1 port map( A1 => n24392, A2 => n19895, Z => n3336);
   U4330 : INV_X4 port map( I => n15885, ZN => n16299);
   U1795 : INV_X1 port map( I => n23344, ZN => n8500);
   U457 : NAND2_X2 port map( A1 => n427, A2 => n782, ZN => n12058);
   U489 : NAND2_X2 port map( A1 => n171, A2 => n820, ZN => n9012);
   U2911 : OAI22_X2 port map( A1 => n2445, A2 => n10437, B1 => n18588, B2 => 
                           n18628, ZN => n171);
   U5364 : OAI21_X2 port map( A1 => n6192, A2 => n7064, B => n16188, ZN => 
                           n4062);
   U1061 : INV_X4 port map( I => n14639, ZN => n24091);
   U18282 : NOR2_X2 port map( A1 => n23197, A2 => n21842, ZN => n17692);
   U908 : AOI21_X2 port map( A1 => n15878, A2 => n15770, B => n10451, ZN => 
                           n10450);
   U21788 : OR2_X2 port map( A1 => n27401, A2 => n19645, Z => n19925);
   U10945 : NOR3_X1 port map( A1 => n1376, A2 => n22551, A3 => n18895, ZN => 
                           n18638);
   U5084 : INV_X2 port map( I => n25225, ZN => n15497);
   U5637 : INV_X2 port map( I => n10640, ZN => n13619);
   U377 : INV_X2 port map( I => n4175, ZN => n19328);
   U1807 : INV_X2 port map( I => n1551, ZN => n18581);
   U3034 : OR2_X2 port map( A1 => n6850, A2 => n6849, Z => n22796);
   U13958 : INV_X4 port map( I => n26296, ZN => n11454);
   U5539 : INV_X2 port map( I => n10301, ZN => n12218);
   U17795 : INV_X1 port map( I => n24566, ZN => n17348);
   U1486 : BUF_X4 port map( I => n19863, Z => n19918);
   U14650 : INV_X2 port map( I => n16466, ZN => n16663);
   U5028 : INV_X2 port map( I => n14658, ZN => n17499);
   U6447 : AOI21_X1 port map( A1 => n17809, A2 => n1349, B => n7599, ZN => 
                           n8612);
   U1238 : OAI21_X2 port map( A1 => n1055, A2 => n13307, B => n14695, ZN => 
                           n22117);
   U2963 : INV_X2 port map( I => n4414, ZN => n1219);
   U4105 : NOR2_X2 port map( A1 => n198, A2 => n199, ZN => n13232);
   U7103 : OAI21_X2 port map( A1 => n14176, A2 => n25175, B => n25759, ZN => 
                           n9306);
   U4491 : INV_X2 port map( I => n8344, ZN => n5266);
   U859 : INV_X4 port map( I => n15029, ZN => n4630);
   U16153 : NAND3_X1 port map( A1 => n14163, A2 => n10272, A3 => n19765, ZN => 
                           n9689);
   U1890 : INV_X4 port map( I => n997, ZN => n75);
   U1170 : OAI21_X2 port map( A1 => n16656, A2 => n16657, B => n22280, ZN => 
                           n11067);
   U1911 : NAND3_X2 port map( A1 => n2692, A2 => n2693, A3 => n6911, ZN => 
                           n5159);
   U1118 : INV_X2 port map( I => n2577, ZN => n2490);
   U5773 : AOI21_X2 port map( A1 => n4784, A2 => n12734, B => n2557, ZN => 
                           n13402);
   U2121 : AOI22_X2 port map( A1 => n11674, A2 => n17302, B1 => n17307, B2 => 
                           n17306, ZN => n23160);
   U8052 : NAND2_X2 port map( A1 => n4166, A2 => n4165, ZN => n4164);
   U10682 : BUF_X2 port map( I => Key(166), Z => n14544);
   U7491 : NOR2_X2 port map( A1 => n18490, A2 => n26121, ZN => n9602);
   U4715 : INV_X1 port map( I => n25105, ZN => n2796);
   U1454 : NOR2_X2 port map( A1 => n5746, A2 => n25261, ZN => n5705);
   U20169 : INV_X1 port map( I => n22819, ZN => n822);
   U12419 : NAND2_X2 port map( A1 => n18771, A2 => n14095, ZN => n3030);
   U3095 : AOI21_X1 port map( A1 => n9087, A2 => n5906, B => n734, ZN => n11243
                           );
   U6317 : OAI21_X2 port map( A1 => n7741, A2 => n18378, B => n18585, ZN => 
                           n7740);
   U604 : NAND2_X2 port map( A1 => n26243, A2 => n12562, ZN => n12561);
   U6404 : INV_X1 port map( I => n22325, ZN => n15568);
   U7632 : NAND2_X2 port map( A1 => n794, A2 => n9759, ZN => n22162);
   U15546 : INV_X4 port map( I => n19937, ZN => n19785);
   U4816 : BUF_X4 port map( I => n16846, Z => n17436);
   U19432 : INV_X2 port map( I => n9906, ZN => n10161);
   U19434 : NAND2_X2 port map( A1 => n5681, A2 => n564, ZN => n9906);
   U9913 : OAI21_X2 port map( A1 => n9466, A2 => n9948, B => n28367, ZN => 
                           n6226);
   U5318 : INV_X2 port map( I => n25013, ZN => n17312);
   U9776 : NOR2_X2 port map( A1 => n5480, A2 => n1020, ZN => n3072);
   U1680 : NAND2_X2 port map( A1 => n25144, A2 => n6629, ZN => n22353);
   U1506 : AOI21_X2 port map( A1 => n19758, A2 => n19752, B => n19630, ZN => 
                           n6682);
   U17473 : INV_X2 port map( I => n304, ZN => n19752);
   U1469 : AOI21_X1 port map( A1 => n23649, A2 => n27926, B => n12919, ZN => 
                           n24423);
   U3797 : NAND2_X1 port map( A1 => n2675, A2 => n3469, ZN => n22093);
   U2464 : OAI21_X1 port map( A1 => n4753, A2 => n1987, B => n1985, ZN => 
                           n16047);
   U10998 : NAND3_X1 port map( A1 => n6892, A2 => n22244, A3 => n22337, ZN => 
                           n22558);
   U1286 : BUF_X2 port map( I => n9218, Z => n22801);
   U1860 : INV_X2 port map( I => n1037, ZN => n17172);
   U4755 : BUF_X2 port map( I => n2398, Z => n2177);
   U15760 : NOR2_X2 port map( A1 => n10161, A2 => n23270, ZN => n6730);
   U8356 : BUF_X2 port map( I => Key(57), Z => n14591);
   U13541 : OAI21_X1 port map( A1 => n14395, A2 => n18939, B => n6487, ZN => 
                           n22860);
   U10603 : INV_X2 port map( I => n840, ZN => n1268);
   U4412 : NOR2_X2 port map( A1 => n12272, A2 => n5362, ZN => n12274);
   U4383 : NOR2_X1 port map( A1 => n2472, A2 => n20238, ZN => n2471);
   U996 : INV_X2 port map( I => n1886, ZN => n13477);
   U16098 : AOI21_X2 port map( A1 => n26321, A2 => n879, B => n25935, ZN => 
                           n12348);
   U8921 : NAND3_X1 port map( A1 => n10011, A2 => n10012, A3 => n1016, ZN => 
                           n23884);
   U9255 : NAND2_X1 port map( A1 => n8321, A2 => n18820, ZN => n8320);
   U5261 : BUF_X4 port map( I => n7987, Z => n8070);
   U5409 : INV_X2 port map( I => n13417, ZN => n798);
   U21721 : OAI21_X1 port map( A1 => n24387, A2 => n27351, B => n24386, ZN => 
                           n17231);
   U4387 : NAND3_X1 port map( A1 => n6160, A2 => n15413, A3 => n22758, ZN => 
                           n6159);
   U16158 : OAI21_X2 port map( A1 => n11663, A2 => n18100, B => n25192, ZN => 
                           n11664);
   U8727 : INV_X2 port map( I => n20489, ZN => n11885);
   U10665 : BUF_X2 port map( I => Key(104), Z => n14600);
   U12243 : OAI21_X2 port map( A1 => n28240, A2 => n2798, B => n23597, ZN => 
                           n18961);
   U19692 : NAND2_X1 port map( A1 => n17490, A2 => n17362, ZN => n13385);
   U1205 : INV_X2 port map( I => n13927, ZN => n13690);
   U4994 : NOR2_X1 port map( A1 => n14708, A2 => n14706, ZN => n14705);
   U20300 : OAI21_X2 port map( A1 => n11878, A2 => n11877, B => n24093, ZN => 
                           n11876);
   U7936 : INV_X2 port map( I => n9362, ZN => n14578);
   U833 : NOR2_X1 port map( A1 => n17856, A2 => n26491, ZN => n22086);
   U14760 : NAND2_X1 port map( A1 => n20779, A2 => n27332, ZN => n9029);
   U5448 : NAND2_X2 port map( A1 => n15689, A2 => n20739, ZN => n20785);
   U8618 : OAI21_X1 port map( A1 => n20781, A2 => n20586, B => n9333, ZN => 
                           n20428);
   U14202 : OAI21_X1 port map( A1 => n11270, A2 => n17510, B => n23040, ZN => 
                           n22986);
   U2636 : INV_X1 port map( I => n13043, ZN => n7961);
   U9821 : NAND2_X1 port map( A1 => n15384, A2 => n3611, ZN => n17741);
   U10003 : INV_X1 port map( I => n17295, ZN => n3848);
   U1561 : NAND3_X2 port map( A1 => n10520, A2 => n978, A3 => n12395, ZN => 
                           n20111);
   U6494 : NOR2_X1 port map( A1 => n11738, A2 => n13291, ZN => n11737);
   U8255 : INV_X2 port map( I => n16088, ZN => n14763);
   U14549 : INV_X1 port map( I => n10569, ZN => n18385);
   U8026 : AOI21_X2 port map( A1 => n16491, A2 => n24334, B => n16490, ZN => 
                           n5518);
   U1595 : NAND2_X2 port map( A1 => n21332, A2 => n22212, ZN => n5251);
   U20621 : AOI21_X1 port map( A1 => n16653, A2 => n434, B => n16566, ZN => 
                           n16568);
   U3114 : BUF_X2 port map( I => n11215, Z => n23065);
   U5051 : INV_X2 port map( I => n5442, ZN => n1243);
   U6813 : NAND2_X2 port map( A1 => n11423, A2 => n15686, ZN => n2342);
   U6507 : INV_X1 port map( I => n26939, ZN => n14234);
   U14758 : INV_X4 port map( I => n6459, ZN => n23110);
   U777 : BUF_X4 port map( I => n16935, Z => n17518);
   U4397 : BUF_X2 port map( I => n21885, Z => n24132);
   U16682 : NOR2_X2 port map( A1 => n15331, A2 => n10707, ZN => n4647);
   U10439 : NAND2_X2 port map( A1 => n26186, A2 => n15919, ZN => n4032);
   U16918 : AND2_X2 port map( A1 => n652, A2 => n18385, Z => n23534);
   U12156 : OAI22_X2 port map( A1 => n6538, A2 => n13025, B1 => n1048, B2 => 
                           n16378, ZN => n13309);
   U4512 : CLKBUF_X2 port map( I => Key(81), Z => n7397);
   U3012 : BUF_X2 port map( I => Key(85), Z => n14360);
   U8388 : CLKBUF_X2 port map( I => Key(143), Z => n20683);
   U8366 : BUF_X2 port map( I => Key(93), Z => n21557);
   U6867 : BUF_X2 port map( I => Key(76), Z => n21044);
   U5846 : BUF_X2 port map( I => Key(186), Z => n14535);
   U8338 : BUF_X2 port map( I => Key(39), Z => n20949);
   U4341 : CLKBUF_X2 port map( I => Key(65), Z => n19346);
   U5837 : BUF_X2 port map( I => Key(118), Z => n14432);
   U6864 : BUF_X2 port map( I => Key(151), Z => n21033);
   U10639 : BUF_X2 port map( I => Key(120), Z => n20769);
   U3394 : BUF_X2 port map( I => Key(68), Z => n20692);
   U10643 : BUF_X2 port map( I => Key(148), Z => n14436);
   U8377 : CLKBUF_X2 port map( I => Key(113), Z => n21367);
   U8311 : INV_X1 port map( I => Key(136), ZN => n1283);
   U20391 : BUF_X2 port map( I => Key(116), Z => n21650);
   U5835 : BUF_X2 port map( I => Key(61), Z => n21336);
   U6861 : BUF_X2 port map( I => Key(82), Z => n20702);
   U10683 : BUF_X2 port map( I => Key(105), Z => n14624);
   U6873 : BUF_X2 port map( I => Key(60), Z => n21613);
   U10698 : BUF_X2 port map( I => Key(31), Z => n20614);
   U8392 : BUF_X2 port map( I => Key(190), Z => n14573);
   U6869 : BUF_X2 port map( I => Key(52), Z => n14589);
   U8360 : BUF_X2 port map( I => Key(174), Z => n14418);
   U5087 : BUF_X2 port map( I => Key(181), Z => n20602);
   U3011 : BUF_X2 port map( I => Key(162), Z => n14549);
   U10625 : CLKBUF_X2 port map( I => n11395, Z => n10970);
   U1828 : INV_X1 port map( I => n16141, ZN => n14857);
   U10476 : INV_X1 port map( I => n21436, ZN => n6287);
   U10585 : CLKBUF_X1 port map( I => n16274, Z => n13577);
   U2455 : CLKBUF_X4 port map( I => n569, Z => n21764);
   U20529 : NAND2_X1 port map( A1 => n15937, A2 => n16167, ZN => n15938);
   U1254 : NAND2_X1 port map( A1 => n14386, A2 => n13857, ZN => n9794);
   U1792 : NAND2_X1 port map( A1 => n3850, A2 => n15919, ZN => n14888);
   U10539 : BUF_X2 port map( I => n15330, Z => n3298);
   U8281 : OAI21_X1 port map( A1 => n7022, A2 => n15330, B => n16189, ZN => 
                           n6193);
   U18017 : INV_X1 port map( I => n16318, ZN => n12509);
   U8236 : NAND2_X1 port map( A1 => n14763, A2 => n14764, ZN => n7406);
   U2716 : OAI21_X1 port map( A1 => n15769, A2 => n15921, B => n16340, ZN => 
                           n3521);
   U10506 : INV_X1 port map( I => n16050, ZN => n15853);
   U14233 : NOR2_X1 port map( A1 => n4751, A2 => n15787, ZN => n4753);
   U21352 : NOR2_X1 port map( A1 => n22454, A2 => n24591, ZN => n24247);
   U15715 : NAND2_X1 port map( A1 => n14559, A2 => n6647, ZN => n15942);
   U10446 : NAND2_X1 port map( A1 => n13123, A2 => n15946, ZN => n8410);
   U16732 : AOI21_X1 port map( A1 => n15776, A2 => n7235, B => n14636, ZN => 
                           n8157);
   U4349 : NAND2_X1 port map( A1 => n24376, A2 => n13306, ZN => n11545);
   U10360 : CLKBUF_X2 port map( I => n11908, Z => n14337);
   U20943 : CLKBUF_X2 port map( I => n16691, Z => n24183);
   U3006 : BUF_X2 port map( I => n14137, Z => n23134);
   U1397 : INV_X2 port map( I => n7265, ZN => n16409);
   U14283 : AOI21_X1 port map( A1 => n14264, A2 => n6911, B => n1246, ZN => 
                           n16726);
   U11103 : NAND2_X1 port map( A1 => n4756, A2 => n3399, ZN => n24029);
   U2776 : NAND2_X1 port map( A1 => n16048, A2 => n26024, ZN => n300);
   U18271 : NAND2_X1 port map( A1 => n15442, A2 => n25487, ZN => n15441);
   U16634 : OAI22_X1 port map( A1 => n9764, A2 => n8223, B1 => n16705, B2 => 
                           n905, ZN => n7921);
   U18963 : NAND2_X1 port map( A1 => n16515, A2 => n16572, ZN => n13546);
   U18027 : INV_X1 port map( I => n16693, ZN => n12504);
   U18200 : INV_X1 port map( I => n16845, ZN => n23754);
   U1100 : INV_X1 port map( I => n12831, ZN => n23345);
   U14846 : CLKBUF_X2 port map( I => n16845, Z => n23137);
   U10110 : BUF_X2 port map( I => n17183, Z => n13358);
   U4192 : CLKBUF_X4 port map( I => n16998, Z => n17306);
   U10107 : INV_X2 port map( I => n11581, ZN => n2831);
   U1048 : CLKBUF_X4 port map( I => n2901, Z => n2814);
   U782 : INV_X2 port map( I => n17353, ZN => n13740);
   U1717 : INV_X2 port map( I => n24513, ZN => n17507);
   U728 : INV_X2 port map( I => n8996, ZN => n11284);
   U2984 : CLKBUF_X2 port map( I => n28538, Z => n23449);
   U19485 : NAND2_X1 port map( A1 => n23971, A2 => n1234, ZN => n5693);
   U4575 : INV_X1 port map( I => n4111, ZN => n1952);
   U19095 : NAND2_X1 port map( A1 => n17534, A2 => n11857, ZN => n13339);
   U13834 : CLKBUF_X2 port map( I => n7370, Z => n22918);
   U17915 : INV_X1 port map( I => n14862, ZN => n17229);
   U20022 : OAI21_X1 port map( A1 => n17307, A2 => n16999, B => n17176, ZN => 
                           n17179);
   U4147 : NOR2_X1 port map( A1 => n17576, A2 => n1228, ZN => n23724);
   U1028 : OAI21_X1 port map( A1 => n613, A2 => n23778, B => n12882, ZN => 
                           n13245);
   U4129 : CLKBUF_X2 port map( I => n2636, Z => n22724);
   U678 : CLKBUF_X2 port map( I => n13043, Z => n3621);
   U4475 : INV_X2 port map( I => n2897, ZN => n727);
   U4618 : INV_X1 port map( I => n4486, ZN => n14707);
   U7710 : INV_X2 port map( I => n14792, ZN => n6892);
   U10734 : INV_X2 port map( I => n17824, ZN => n1349);
   U7762 : BUF_X2 port map( I => n17897, Z => n7120);
   U6086 : NOR2_X1 port map( A1 => n7599, A2 => n17935, ZN => n17810);
   U17933 : OAI22_X1 port map( A1 => n17740, A2 => n14397, B1 => n6892, B2 => 
                           n17582, ZN => n14403);
   U14516 : INV_X2 port map( I => n7358, ZN => n23044);
   U2603 : NOR2_X1 port map( A1 => n23245, A2 => n26055, ZN => n9269);
   U19339 : NAND2_X1 port map( A1 => n17608, A2 => n12850, ZN => n14318);
   U12075 : AOI21_X1 port map( A1 => n1219, A2 => n22724, B => n23391, ZN => 
                           n15384);
   U18075 : NAND2_X1 port map( A1 => n17686, A2 => n27862, ZN => n14467);
   U9779 : OAI21_X1 port map( A1 => n24518, A2 => n5296, B => n6910, ZN => 
                           n5779);
   U18485 : NAND2_X1 port map( A1 => n17791, A2 => n11498, ZN => n17792);
   U7634 : INV_X1 port map( I => n4558, ZN => n8790);
   U12329 : INV_X2 port map( I => n2912, ZN => n11425);
   U768 : CLKBUF_X2 port map( I => n18574, Z => n14569);
   U9622 : CLKBUF_X2 port map( I => n18482, Z => n14420);
   U2996 : CLKBUF_X2 port map( I => n10570, Z => n348);
   U7620 : BUF_X2 port map( I => n13181, Z => n4661);
   U15938 : CLKBUF_X1 port map( I => n6144, Z => n23361);
   U16108 : AND2_X1 port map( A1 => n2912, A2 => n18456, Z => n9730);
   U3258 : CLKBUF_X2 port map( I => n6029, Z => n22973);
   U6380 : CLKBUF_X2 port map( I => n18612, Z => n9248);
   U18124 : CLKBUF_X4 port map( I => n10536, Z => n23743);
   U3244 : CLKBUF_X4 port map( I => n10614, Z => n21790);
   U19131 : CLKBUF_X2 port map( I => n1172, Z => n23889);
   U6399 : INV_X2 port map( I => n23004, ZN => n1004);
   U559 : INV_X2 port map( I => n12699, ZN => n12979);
   U3261 : CLKBUF_X1 port map( I => n18466, Z => n24054);
   U7570 : NOR2_X1 port map( A1 => n25500, A2 => n18454, ZN => n3763);
   U11828 : NOR2_X1 port map( A1 => n3903, A2 => n1010, ZN => n12189);
   U9596 : INV_X1 port map( I => n12325, ZN => n10250);
   U20956 : NAND2_X1 port map( A1 => n7770, A2 => n376, ZN => n18460);
   U20885 : NAND2_X1 port map( A1 => n18064, A2 => n7350, ZN => n18065);
   U17943 : NAND2_X1 port map( A1 => n18506, A2 => n11817, ZN => n11744);
   U3948 : OAI21_X1 port map( A1 => n7276, A2 => n7277, B => n5338, ZN => 
                           n23363);
   U16326 : OAI21_X1 port map( A1 => n21795, A2 => n23436, B => n11783, ZN => 
                           n23716);
   U3235 : INV_X1 port map( I => n18533, ZN => n24149);
   U17932 : NAND2_X1 port map( A1 => n18723, A2 => n18724, ZN => n15380);
   U7500 : INV_X2 port map( I => n18879, ZN => n999);
   U7445 : INV_X2 port map( I => n19150, ZN => n14925);
   U2891 : NAND3_X1 port map( A1 => n23742, A2 => n26778, A3 => n4549, ZN => 
                           n21962);
   U12680 : INV_X2 port map( I => n14836, ZN => n3619);
   U11365 : NOR2_X1 port map( A1 => n6889, A2 => n14237, ZN => n22633);
   U1668 : INV_X2 port map( I => n3932, ZN => n18895);
   U9384 : AND2_X1 port map( A1 => n12667, A2 => n19045, Z => n10709);
   U1636 : AOI22_X1 port map( A1 => n7551, A2 => n14836, B1 => n14545, B2 => 
                           n18903, ZN => n23097);
   U474 : OAI21_X1 port map( A1 => n26327, A2 => n19123, B => n2616, ZN => 
                           n22566);
   U15639 : NAND2_X1 port map( A1 => n12589, A2 => n6534, ZN => n6533);
   U21024 : NAND2_X1 port map( A1 => n19087, A2 => n19117, ZN => n19002);
   U3910 : NAND3_X1 port map( A1 => n12583, A2 => n23575, A3 => n19122, ZN => 
                           n24239);
   U16821 : NOR2_X1 port map( A1 => n816, A2 => n21765, ZN => n15299);
   U3838 : NAND2_X1 port map( A1 => n18851, A2 => n11576, ZN => n23434);
   U7395 : AOI21_X1 port map( A1 => n2746, A2 => n19120, B => n8740, ZN => 
                           n6783);
   U413 : INV_X1 port map( I => n19522, ZN => n9283);
   U21080 : INV_X1 port map( I => n19352, ZN => n19299);
   U9204 : INV_X1 port map( I => n27624, ZN => n9316);
   U9198 : INV_X1 port map( I => n19327, ZN => n4615);
   U18941 : INV_X1 port map( I => n19905, ZN => n19907);
   U1474 : CLKBUF_X4 port map( I => n11287, Z => n1121);
   U3168 : CLKBUF_X2 port map( I => n19905, Z => n24109);
   U11485 : BUF_X4 port map( I => n10057, Z => n11936);
   U14645 : INV_X2 port map( I => n23081, ZN => n669);
   U4255 : BUF_X2 port map( I => n19781, Z => n4480);
   U4244 : INV_X2 port map( I => n10978, ZN => n967);
   U2226 : NAND2_X1 port map( A1 => n9887, A2 => n19882, ZN => n8487);
   U342 : INV_X2 port map( I => n12863, ZN => n14282);
   U3059 : INV_X2 port map( I => n9361, ZN => n19599);
   U9020 : NAND2_X1 port map( A1 => n24679, A2 => n19597, ZN => n7584);
   U1898 : INV_X1 port map( I => n8487, ZN => n6571);
   U18150 : OAI21_X1 port map( A1 => n19623, A2 => n12431, B => n10411, ZN => 
                           n13002);
   U265 : INV_X1 port map( I => n815, ZN => n19838);
   U5491 : OAI21_X1 port map( A1 => n6571, A2 => n6570, B => n865, ZN => n13434
                           );
   U15287 : INV_X4 port map( I => n3101, ZN => n23253);
   U3118 : NOR2_X1 port map( A1 => n11303, A2 => n19574, ZN => n22617);
   U8903 : NAND2_X1 port map( A1 => n5047, A2 => n675, ZN => n14481);
   U5025 : INV_X2 port map( I => n20195, ZN => n733);
   U3110 : CLKBUF_X4 port map( I => n13248, Z => n23906);
   U17327 : NAND2_X1 port map( A1 => n960, A2 => n1366, ZN => n9462);
   U15726 : NAND2_X1 port map( A1 => n2599, A2 => n20308, ZN => n6670);
   U165 : AOI21_X1 port map( A1 => n8032, A2 => n20269, B => n10885, ZN => 
                           n10901);
   U6089 : INV_X2 port map( I => n2656, ZN => n13147);
   U7625 : NAND2_X1 port map( A1 => n5354, A2 => n959, ZN => n6097);
   U230 : BUF_X2 port map( I => n20338, Z => n3290);
   U8783 : NAND2_X1 port map( A1 => n8204, A2 => n9191, ZN => n3728);
   U8788 : NAND2_X1 port map( A1 => n13454, A2 => n20262, ZN => n13453);
   U8787 : INV_X2 port map( I => n1355, ZN => n3707);
   U8732 : INV_X1 port map( I => n21364, ZN => n3392);
   U3528 : BUF_X2 port map( I => n21270, Z => n9378);
   U3495 : CLKBUF_X2 port map( I => n4860, Z => n480);
   U16241 : NOR2_X1 port map( A1 => n10630, A2 => n20951, ZN => n20945);
   U8345 : BUF_X2 port map( I => Key(48), Z => n20584);
   U10653 : BUF_X2 port map( I => Key(108), Z => n14564);
   U10680 : CLKBUF_X2 port map( I => Key(74), Z => n7368);
   U8385 : CLKBUF_X2 port map( I => Key(103), Z => n14555);
   U3010 : BUF_X2 port map( I => n573, Z => n24271);
   U8315 : CLKBUF_X2 port map( I => n15904, Z => n16082);
   U3386 : OAI22_X1 port map( A1 => n1267, A2 => n16350, B1 => n15347, B2 => 
                           n10970, ZN => n24376);
   U17060 : NAND2_X1 port map( A1 => n12605, A2 => n12874, ZN => n8827);
   U10594 : BUF_X1 port map( I => n3443, Z => n22510);
   U12991 : OAI21_X1 port map( A1 => n834, A2 => n4295, B => n3361, ZN => 
                           n15442);
   U17788 : NAND2_X1 port map( A1 => n7265, A2 => n8021, ZN => n16454);
   U2993 : BUF_X2 port map( I => n17337, Z => n347);
   U4189 : BUF_X2 port map( I => n17555, Z => n24299);
   U18945 : NAND2_X1 port map( A1 => n9481, A2 => n17175, ZN => n17176);
   U5291 : AOI21_X1 port map( A1 => n1232, A2 => n831, B => n2814, ZN => n3624)
                           ;
   U5288 : NAND2_X1 port map( A1 => n13568, A2 => n765, ZN => n17545);
   U3250 : INV_X2 port map( I => n3292, ZN => n6709);
   U10946 : NOR2_X1 port map( A1 => n25738, A2 => n8882, ZN => n8884);
   U949 : BUF_X2 port map( I => n4414, Z => n4590);
   U6465 : OR2_X1 port map( A1 => n17968, A2 => n11112, Z => n10300);
   U2920 : BUF_X2 port map( I => n18663, Z => n24207);
   U1518 : INV_X1 port map( I => n1440, ZN => n18589);
   U5229 : INV_X2 port map( I => n18473, ZN => n18472);
   U17005 : INV_X1 port map( I => n8702, ZN => n18704);
   U15216 : INV_X1 port map( I => n8651, ZN => n10596);
   U20075 : AOI21_X1 port map( A1 => n18745, A2 => n14484, B => n18749, ZN => 
                           n17892);
   U9531 : NAND2_X1 port map( A1 => n18572, A2 => n18571, ZN => n14767);
   U9474 : NAND2_X1 port map( A1 => n11946, A2 => n18528, ZN => n2420);
   U3204 : CLKBUF_X2 port map( I => n8611, Z => n22920);
   U2896 : BUF_X2 port map( I => n14382, Z => n23405);
   U2888 : NAND2_X1 port map( A1 => n8226, A2 => n3619, ZN => n3671);
   U1489 : BUF_X2 port map( I => n19672, Z => n19876);
   U13747 : NAND2_X1 port map( A1 => n22903, A2 => n19889, ZN => n13353);
   U9008 : NOR2_X1 port map( A1 => n4439, A2 => n19759, ZN => n4438);
   U8899 : INV_X2 port map( I => n675, ZN => n5163);
   U6088 : INV_X1 port map( I => n21989, ZN => n22843);
   U5093 : INV_X2 port map( I => n21258, ZN => n14699);
   U2187 : NOR2_X2 port map( A1 => n2891, A2 => n11988, ZN => n19858);
   U2461 : OR2_X1 port map( A1 => n11722, A2 => n15960, Z => n3249);
   U15862 : INV_X4 port map( I => n6906, ZN => n9354);
   U4062 : NAND2_X2 port map( A1 => n2781, A2 => n4916, ZN => n2780);
   U3228 : AOI21_X2 port map( A1 => n7867, A2 => n235, B => n22457, ZN => n7865
                           );
   U10198 : NAND2_X2 port map( A1 => n9617, A2 => n9616, ZN => n9615);
   U6731 : NOR2_X2 port map( A1 => n3369, A2 => n13955, ZN => n13954);
   U5828 : INV_X1 port map( I => n16158, ZN => n16317);
   U2465 : NAND2_X1 port map( A1 => n1987, A2 => n23922, ZN => n1986);
   U8304 : INV_X1 port map( I => n16159, ZN => n16318);
   U14061 : NOR2_X1 port map( A1 => n14171, A2 => n4532, ZN => n13406);
   U8225 : NOR2_X1 port map( A1 => n9308, A2 => n16339, ZN => n8666);
   U5070 : NOR2_X1 port map( A1 => n14512, A2 => n16123, ZN => n6236);
   U3688 : INV_X2 port map( I => n16289, ZN => n1260);
   U8297 : INV_X1 port map( I => n15924, ZN => n15926);
   U6827 : INV_X1 port map( I => n7608, ZN => n2148);
   U19787 : AOI21_X1 port map( A1 => n16148, A2 => n13677, B => n16119, ZN => 
                           n16117);
   U5811 : NAND2_X1 port map( A1 => n15832, A2 => n8648, ZN => n15611);
   U10566 : NAND2_X1 port map( A1 => n16298, A2 => n24271, ZN => n13518);
   U20540 : INV_X1 port map( I => n16006, ZN => n16194);
   U5400 : CLKBUF_X2 port map( I => n14886, Z => n7300);
   U10545 : INV_X2 port map( I => n16013, ZN => n9443);
   U6831 : INV_X1 port map( I => n8867, ZN => n1259);
   U4841 : INV_X1 port map( I => n25763, ZN => n16259);
   U3692 : INV_X1 port map( I => n21885, ZN => n16348);
   U6771 : NAND3_X1 port map( A1 => n7022, A2 => n16299, A3 => n16188, ZN => 
                           n16171);
   U8231 : NOR2_X1 port map( A1 => n1260, A2 => n6427, ZN => n3571);
   U17076 : NOR2_X1 port map( A1 => n8873, A2 => n22801, ZN => n8868);
   U1251 : NOR2_X1 port map( A1 => n12116, A2 => n13731, ZN => n12115);
   U1257 : NOR2_X1 port map( A1 => n12918, A2 => n16332, ZN => n23649);
   U20564 : NAND2_X1 port map( A1 => n16320, A2 => n7311, ZN => n16160);
   U18022 : NOR2_X1 port map( A1 => n16017, A2 => n13717, ZN => n15837);
   U1018 : AOI21_X1 port map( A1 => n16298, A2 => n7022, B => n16300, ZN => 
                           n6477);
   U2256 : NOR2_X1 port map( A1 => n15610, A2 => n16027, ZN => n22712);
   U20546 : NAND3_X1 port map( A1 => n577, A2 => n16292, A3 => n3572, ZN => 
                           n16042);
   U1253 : NAND2_X1 port map( A1 => n6427, A2 => n16289, ZN => n16290);
   U11369 : NOR3_X1 port map( A1 => n13742, A2 => n10707, A3 => n1987, ZN => 
                           n16323);
   U1797 : NOR2_X1 port map( A1 => n3850, A2 => n24581, ZN => n12976);
   U10771 : NAND2_X1 port map( A1 => n1269, A2 => n14546, ZN => n16149);
   U8273 : NAND2_X1 port map( A1 => n16011, A2 => n16013, ZN => n15820);
   U10538 : NAND2_X1 port map( A1 => n799, A2 => n14415, ZN => n4287);
   U10486 : NOR2_X1 port map( A1 => n15974, A2 => n838, ZN => n8602);
   U8241 : NOR2_X1 port map( A1 => n2111, A2 => n16307, ZN => n16308);
   U14574 : NAND2_X1 port map( A1 => n3874, A2 => n24581, ZN => n5205);
   U19754 : NOR2_X1 port map( A1 => n14886, A2 => n26702, ZN => n16197);
   U11373 : NAND2_X1 port map( A1 => n4752, A2 => n1987, ZN => n1985);
   U13465 : AND2_X1 port map( A1 => n25365, A2 => n24581, Z => n13781);
   U20447 : NAND2_X1 port map( A1 => n14559, A2 => n13742, ZN => n15788);
   U4840 : NAND3_X1 port map( A1 => n914, A2 => n27240, A3 => n840, ZN => n2047
                           );
   U5915 : INV_X1 port map( I => n21970, ZN => n6612);
   U20514 : OAI21_X1 port map( A1 => n16125, A2 => n15868, B => n15995, ZN => 
                           n15871);
   U13566 : AOI21_X1 port map( A1 => n8603, A2 => n838, B => n8602, ZN => 
                           n23635);
   U8151 : NAND2_X1 port map( A1 => n16078, A2 => n8212, ZN => n8211);
   U10407 : NAND2_X1 port map( A1 => n10820, A2 => n10819, ZN => n4555);
   U1083 : NAND2_X1 port map( A1 => n14766, A2 => n25693, ZN => n14008);
   U10350 : NAND2_X1 port map( A1 => n10261, A2 => n8344, ZN => n10259);
   U20013 : INV_X2 port map( I => n16483, ZN => n14264);
   U11913 : NOR2_X1 port map( A1 => n14676, A2 => n9683, ZN => n2762);
   U8084 : NAND2_X1 port map( A1 => n10422, A2 => n22529, ZN => n4554);
   U3420 : INV_X1 port map( I => n14878, ZN => n16584);
   U8127 : INV_X1 port map( I => n16224, ZN => n16609);
   U2057 : INV_X1 port map( I => n12482, ZN => n1051);
   U10241 : NOR2_X1 port map( A1 => n1051, A2 => n5122, ZN => n5121);
   U18273 : NOR2_X1 port map( A1 => n16617, A2 => n5062, ZN => n15815);
   U6654 : NAND2_X1 port map( A1 => n16585, A2 => n23758, ZN => n7046);
   U1381 : NOR2_X1 port map( A1 => n24812, A2 => n16658, ZN => n22281);
   U3004 : CLKBUF_X2 port map( I => n16494, Z => n23048);
   U19698 : NAND2_X1 port map( A1 => n16456, A2 => n28083, ZN => n13391);
   U15463 : NAND2_X1 port map( A1 => n145, A2 => n5442, ZN => n15419);
   U2131 : NAND2_X1 port map( A1 => n24844, A2 => n8084, ZN => n16428);
   U857 : INV_X1 port map( I => n16691, ZN => n6399);
   U876 : INV_X1 port map( I => n7180, ZN => n16690);
   U5349 : INV_X1 port map( I => n25693, ZN => n14656);
   U13972 : NOR2_X1 port map( A1 => n12039, A2 => n6373, ZN => n14056);
   U10887 : NAND3_X1 port map( A1 => n8901, A2 => n13927, A3 => n793, ZN => 
                           n1465);
   U6661 : AOI21_X1 port map( A1 => n4869, A2 => n16707, B => n1253, ZN => 
                           n4870);
   U15283 : NAND2_X1 port map( A1 => n5917, A2 => n25973, ZN => n6249);
   U1162 : NOR2_X1 port map( A1 => n16575, A2 => n14887, ZN => n13606);
   U4309 : NAND3_X1 port map( A1 => n15186, A2 => n22614, A3 => n5558, ZN => 
                           n6346);
   U18657 : NAND2_X1 port map( A1 => n9829, A2 => n9830, ZN => n16552);
   U8001 : NAND3_X1 port map( A1 => n5235, A2 => n4938, A3 => n1597, ZN => 
                           n1596);
   U846 : OAI21_X1 port map( A1 => n16611, A2 => n23048, B => n25698, ZN => 
                           n2116);
   U20625 : NAND3_X1 port map( A1 => n173, A2 => n16617, A3 => n25287, ZN => 
                           n16624);
   U19922 : NOR2_X1 port map( A1 => n14056, A2 => n1053, ZN => n14055);
   U15984 : CLKBUF_X2 port map( I => n7257, Z => n23369);
   U1105 : BUF_X2 port map( I => n11408, Z => n9614);
   U1684 : INV_X1 port map( I => n17141, ZN => n9507);
   U10183 : INV_X1 port map( I => n4656, ZN => n2614);
   U5036 : INV_X2 port map( I => n901, ZN => n766);
   U15378 : INV_X2 port map( I => n13509, ZN => n6021);
   U12605 : AND2_X1 port map( A1 => n13727, A2 => n3963, Z => n17358);
   U16589 : NAND2_X1 port map( A1 => n24517, A2 => n17547, ZN => n7845);
   U752 : INV_X2 port map( I => n17362, ZN => n1039);
   U17361 : NOR2_X1 port map( A1 => n26255, A2 => n8093, ZN => n9556);
   U17463 : INV_X1 port map( I => n17412, ZN => n17204);
   U7883 : NAND2_X1 port map( A1 => n17175, A2 => n1629, ZN => n1631);
   U7795 : AOI21_X1 port map( A1 => n8154, A2 => n9661, B => n17508, ZN => 
                           n4160);
   U4613 : NAND2_X1 port map( A1 => n10461, A2 => n17492, ZN => n13779);
   U15228 : INV_X1 port map( I => n1232, ZN => n23227);
   U4600 : NAND2_X1 port map( A1 => n717, A2 => n17418, ZN => n3094);
   U14020 : NOR3_X1 port map( A1 => n3838, A2 => n6672, A3 => n25971, ZN => 
                           n3836);
   U15063 : INV_X1 port map( I => n14997, ZN => n23778);
   U2036 : NOR2_X1 port map( A1 => n10985, A2 => n11992, ZN => n2966);
   U12541 : OR2_X1 port map( A1 => n28538, A2 => n613, Z => n17311);
   U20775 : NAND2_X1 port map( A1 => n9593, A2 => n17486, ZN => n17365);
   U20776 : NAND2_X1 port map( A1 => n25983, A2 => n17561, ZN => n17364);
   U9927 : NAND2_X1 port map( A1 => n17468, A2 => n17467, ZN => n6463);
   U12358 : OAI21_X1 port map( A1 => n17560, A2 => n17559, B => n21798, ZN => 
                           n17562);
   U12234 : NOR2_X1 port map( A1 => n12882, A2 => n14997, ZN => n2790);
   U6608 : NOR2_X1 port map( A1 => n25983, A2 => n17561, ZN => n10432);
   U13336 : NAND3_X1 port map( A1 => n1032, A2 => n2814, A3 => n26161, ZN => 
                           n3625);
   U16623 : NOR2_X1 port map( A1 => n7912, A2 => n12225, ZN => n17521);
   U6521 : NOR2_X1 port map( A1 => n17417, A2 => n3094, ZN => n3093);
   U19461 : NOR2_X1 port map( A1 => n26655, A2 => n17490, ZN => n12765);
   U19914 : NAND2_X1 port map( A1 => n765, A2 => n12340, ZN => n17444);
   U16143 : NAND2_X1 port map( A1 => n17402, A2 => n17468, ZN => n17406);
   U5294 : NOR3_X1 port map( A1 => n1032, A2 => n17188, A3 => n831, ZN => 
                           n10464);
   U15585 : NOR2_X1 port map( A1 => n17199, A2 => n6425, ZN => n17200);
   U4141 : BUF_X4 port map( I => n22085, Z => n21792);
   U1905 : AOI21_X1 port map( A1 => n17492, A2 => n10461, B => n14944, ZN => 
                           n8107);
   U6508 : INV_X2 port map( I => n17992, ZN => n17605);
   U4797 : INV_X1 port map( I => n6098, ZN => n8075);
   U5267 : INV_X1 port map( I => n17898, ZN => n12983);
   U673 : INV_X1 port map( I => n17726, ZN => n1214);
   U887 : NAND2_X1 port map( A1 => n413, A2 => n17906, ZN => n17646);
   U18947 : NAND2_X1 port map( A1 => n2285, A2 => n22851, ZN => n12087);
   U9910 : INV_X1 port map( I => n7298, ZN => n1209);
   U4466 : INV_X1 port map( I => n17895, ZN => n725);
   U2754 : INV_X1 port map( I => n17855, ZN => n1215);
   U20003 : NAND2_X1 port map( A1 => n17904, A2 => n1213, ZN => n14982);
   U15753 : NOR2_X1 port map( A1 => n8070, A2 => n23963, ZN => n8186);
   U14647 : NOR3_X1 port map( A1 => n891, A2 => n18101, A3 => n22739, ZN => 
                           n24087);
   U7715 : NAND2_X1 port map( A1 => n13061, A2 => n17912, ZN => n15531);
   U9811 : NAND2_X1 port map( A1 => n17677, A2 => n25515, ZN => n2958);
   U9813 : NOR2_X1 port map( A1 => n825, A2 => n9691, ZN => n6481);
   U5252 : NOR2_X1 port map( A1 => n17801, A2 => n12815, ZN => n11808);
   U4116 : NAND2_X1 port map( A1 => n7984, A2 => n8070, ZN => n7983);
   U18294 : OAI21_X1 port map( A1 => n13061, A2 => n23044, B => n11653, ZN => 
                           n11652);
   U18927 : NOR2_X1 port map( A1 => n1210, A2 => n11579, ZN => n12677);
   U20820 : AOI21_X1 port map( A1 => n28239, A2 => n25, B => n5218, ZN => 
                           n17686);
   U16810 : NAND2_X1 port map( A1 => n2285, A2 => n25966, ZN => n17714);
   U18969 : NOR2_X1 port map( A1 => n17581, A2 => n11419, ZN => n17583);
   U6361 : NOR2_X1 port map( A1 => n8882, A2 => n25, ZN => n8883);
   U7628 : INV_X1 port map( I => n23186, ZN => n6744);
   U798 : INV_X1 port map( I => n13119, ZN => n18068);
   U2938 : INV_X1 port map( I => n18243, ZN => n23429);
   U13536 : NAND2_X1 port map( A1 => n18663, A2 => n14745, ZN => n18722);
   U12707 : INV_X2 port map( I => n14745, ZN => n1184);
   U7554 : NAND2_X1 port map( A1 => n18552, A2 => n738, ZN => n13192);
   U19773 : NAND3_X1 port map( A1 => n18743, A2 => n26228, A3 => n27457, ZN => 
                           n18744);
   U2950 : AOI21_X1 port map( A1 => n1015, A2 => n15010, B => n877, ZN => n3565
                           );
   U3687 : NAND2_X1 port map( A1 => n25382, A2 => n532, ZN => n4348);
   U17692 : NAND2_X1 port map( A1 => n3903, A2 => n10289, ZN => n11187);
   U9570 : INV_X1 port map( I => n8126, ZN => n18572);
   U7568 : NAND2_X1 port map( A1 => n12573, A2 => n1407, ZN => n6689);
   U712 : NOR2_X1 port map( A1 => n14371, A2 => n881, ZN => n23594);
   U12100 : INV_X2 port map( I => n18633, ZN => n18769);
   U724 : NOR2_X1 port map( A1 => n8022, A2 => n738, ZN => n18483);
   U18901 : NOR2_X1 port map( A1 => n10904, A2 => n18778, ZN => n18506);
   U4793 : AOI21_X1 port map( A1 => n18625, A2 => n8254, B => n10009, ZN => 
                           n10918);
   U11511 : OAI21_X1 port map( A1 => n18387, A2 => n12979, B => n7078, ZN => 
                           n12938);
   U1412 : NOR2_X1 port map( A1 => n18684, A2 => n18685, ZN => n5642);
   U698 : NOR2_X1 port map( A1 => n8022, A2 => n14420, ZN => n14361);
   U693 : NAND2_X1 port map( A1 => n5439, A2 => n1013, ZN => n23092);
   U4721 : NOR2_X1 port map( A1 => n27895, A2 => n6800, ZN => n15399);
   U7524 : NOR2_X1 port map( A1 => n18529, A2 => n23743, ZN => n11946);
   U7569 : INV_X1 port map( I => n18476, ZN => n6440);
   U17946 : NAND2_X1 port map( A1 => n1502, A2 => n3565, ZN => n23722);
   U14058 : NAND2_X1 port map( A1 => n5746, A2 => n737, ZN => n18415);
   U7538 : AOI21_X1 port map( A1 => n18413, A2 => n25712, B => n737, ZN => 
                           n18369);
   U1349 : OAI21_X1 port map( A1 => n18383, A2 => n18381, B => n3554, ZN => 
                           n18382);
   U4763 : AOI21_X1 port map( A1 => n759, A2 => n25769, B => n10537, ZN => 
                           n2418);
   U3234 : NAND3_X1 port map( A1 => n18533, A2 => n1017, A3 => n1005, ZN => 
                           n13005);
   U6335 : AOI22_X1 port map( A1 => n18529, A2 => n7446, B1 => n12832, B2 => 
                           n23743, ZN => n9470);
   U17445 : OAI21_X1 port map( A1 => n18583, A2 => n7190, B => n18507, ZN => 
                           n14219);
   U18955 : NAND3_X1 port map( A1 => n12305, A2 => n14648, A3 => n12375, ZN => 
                           n12304);
   U9497 : NOR2_X1 port map( A1 => n18415, A2 => n18604, ZN => n7771);
   U6298 : NOR2_X1 port map( A1 => n8877, A2 => n22518, ZN => n1872);
   U7523 : NOR2_X1 port map( A1 => n18491, A2 => n882, ZN => n4292);
   U3720 : INV_X2 port map( I => n25798, ZN => n19052);
   U21882 : INV_X1 port map( I => n19164, ZN => n3276);
   U6253 : NOR2_X1 port map( A1 => n4705, A2 => n15041, ZN => n3610);
   U1857 : NAND2_X1 port map( A1 => n15480, A2 => n18977, ZN => n22075);
   U12623 : NAND2_X1 port map( A1 => n12360, A2 => n18798, ZN => n12359);
   U440 : INV_X1 port map( I => n18996, ZN => n133);
   U13051 : NAND2_X1 port map( A1 => n12781, A2 => n7084, ZN => n12961);
   U498 : NOR2_X1 port map( A1 => n6598, A2 => n11696, ZN => n22096);
   U9397 : NAND2_X1 port map( A1 => n11331, A2 => n444, ZN => n18233);
   U15275 : NAND3_X1 port map( A1 => n987, A2 => n5840, A3 => n25559, ZN => 
                           n12132);
   U21715 : INV_X1 port map( I => n10362, ZN => n6708);
   U1887 : NAND2_X1 port map( A1 => n18910, A2 => n26345, ZN => n23057);
   U19165 : NOR2_X1 port map( A1 => n27175, A2 => n24801, ZN => n19037);
   U454 : INV_X2 port map( I => n4703, ZN => n18964);
   U15969 : OAI21_X1 port map( A1 => n25592, A2 => n18798, B => n18991, ZN => 
                           n18993);
   U17405 : NAND2_X1 port map( A1 => n18819, A2 => n4703, ZN => n9658);
   U7422 : NOR2_X1 port map( A1 => n2070, A2 => n13942, ZN => n13183);
   U2742 : NOR2_X1 port map( A1 => n9922, A2 => n22345, ZN => n7502);
   U4258 : NAND2_X1 port map( A1 => n19109, A2 => n2356, ZN => n13882);
   U9357 : NAND2_X1 port map( A1 => n12961, A2 => n23920, ZN => n12960);
   U385 : NAND2_X1 port map( A1 => n9233, A2 => n1165, ZN => n9232);
   U5978 : AOI21_X1 port map( A1 => n18895, A2 => n23905, B => n25411, ZN => 
                           n10812);
   U6252 : NAND2_X1 port map( A1 => n19052, A2 => n27868, ZN => n12452);
   U9340 : NOR3_X1 port map( A1 => n8554, A2 => n873, A3 => n25381, ZN => n8553
                           );
   U6246 : OAI21_X1 port map( A1 => n13942, A2 => n18948, B => n4206, ZN => 
                           n9327);
   U7329 : INV_X1 port map( I => n2016, ZN => n5804);
   U15352 : INV_X1 port map( I => n7659, ZN => n19432);
   U3020 : INV_X1 port map( I => n11220, ZN => n10291);
   U5535 : INV_X1 port map( I => n19744, ZN => n4132);
   U2918 : INV_X2 port map( I => n735, ZN => n724);
   U19915 : NOR2_X1 port map( A1 => n22140, A2 => n13194, ZN => n14042);
   U7315 : INV_X1 port map( I => n26633, ZN => n976);
   U7311 : NOR2_X1 port map( A1 => n19728, A2 => n1133, ZN => n19857);
   U334 : NAND2_X1 port map( A1 => n8754, A2 => n14393, ZN => n5308);
   U1495 : NOR2_X1 port map( A1 => n28357, A2 => n5253, ZN => n6142);
   U9123 : NOR2_X1 port map( A1 => n2631, A2 => n2632, ZN => n2633);
   U13901 : INV_X1 port map( I => n26625, ZN => n10557);
   U297 : NOR2_X1 port map( A1 => n14789, A2 => n19570, ZN => n19099);
   U18168 : NOR2_X1 port map( A1 => n19889, A2 => n19681, ZN => n19682);
   U4921 : NOR2_X1 port map( A1 => n14726, A2 => n1128, ZN => n14516);
   U363 : AOI21_X1 port map( A1 => n6393, A2 => n24579, B => n19597, ZN => 
                           n7585);
   U9013 : NAND2_X1 port map( A1 => n6875, A2 => n5707, ZN => n6874);
   U21140 : AOI22_X1 port map( A1 => n19616, A2 => n19890, B1 => n810, B2 => 
                           n23782, ZN => n19617);
   U3668 : INV_X1 port map( I => n14752, ZN => n19825);
   U5147 : NOR3_X1 port map( A1 => n8048, A2 => n15027, A3 => n7129, ZN => 
                           n19662);
   U7192 : NAND2_X1 port map( A1 => n4120, A2 => n45, ZN => n1608);
   U13134 : NAND2_X1 port map( A1 => n3657, A2 => n23046, ZN => n22813);
   U2721 : NAND2_X1 port map( A1 => n9525, A2 => n11947, ZN => n11499);
   U8822 : INV_X1 port map( I => n20049, ZN => n2512);
   U20090 : NAND2_X1 port map( A1 => n15732, A2 => n23906, ZN => n14521);
   U223 : NAND2_X1 port map( A1 => n4191, A2 => n25710, ZN => n5203);
   U12550 : NAND2_X1 port map( A1 => n19968, A2 => n7908, ZN => n7143);
   U7167 : NOR2_X1 port map( A1 => n20273, A2 => n25389, ZN => n8205);
   U13243 : INV_X1 port map( I => n2185, ZN => n20254);
   U19599 : INV_X1 port map( I => n20288, ZN => n20089);
   U231 : INV_X1 port map( I => n19989, ZN => n23229);
   U14910 : INV_X2 port map( I => n20324, ZN => n12712);
   U21603 : NAND2_X1 port map( A1 => n20151, A2 => n1366, ZN => n24293);
   U6058 : AOI21_X1 port map( A1 => n8462, A2 => n25390, B => n11786, ZN => 
                           n8461);
   U247 : NOR2_X1 port map( A1 => n22943, A2 => n27630, ZN => n22311);
   U1888 : NAND2_X1 port map( A1 => n13301, A2 => n22295, ZN => n13541);
   U6037 : NOR2_X1 port map( A1 => n4109, A2 => n3870, ZN => n1357);
   U1029 : INV_X1 port map( I => n6215, ZN => n9875);
   U13473 : INV_X1 port map( I => n3803, ZN => n20310);
   U21201 : NAND3_X1 port map( A1 => n20262, A2 => n9875, A3 => n183, ZN => 
                           n19979);
   U5456 : INV_X1 port map( I => n20328, ZN => n2545);
   U9732 : OAI21_X1 port map( A1 => n21865, A2 => n22417, B => n26140, ZN => 
                           n6070);
   U8799 : NOR2_X1 port map( A1 => n20040, A2 => n1835, ZN => n2198);
   U4007 : NAND2_X1 port map( A1 => n20136, A2 => n7122, ZN => n20473);
   U1385 : AOI21_X1 port map( A1 => n20921, A2 => n24539, B => n5797, ZN => 
                           n5799);
   U95 : INV_X2 port map( I => n10797, ZN => n15352);
   U17332 : OR2_X1 port map( A1 => n15728, A2 => n3746, Z => n21061);
   U6009 : NOR2_X1 port map( A1 => n21441, A2 => n13791, ZN => n9715);
   U100 : OAI21_X1 port map( A1 => n21699, A2 => n12290, B => n21724, ZN => 
                           n22655);
   U17262 : NOR2_X1 port map( A1 => n20591, A2 => n15103, ZN => n9280);
   U17981 : NAND2_X1 port map( A1 => n13308, A2 => n1699, ZN => n12374);
   U1157 : NOR2_X1 port map( A1 => n12253, A2 => n10809, ZN => n12252);
   U8651 : NAND2_X1 port map( A1 => n20784, A2 => n20785, ZN => n20789);
   U5561 : INV_X1 port map( I => n21325, ZN => n23514);
   U56 : OAI21_X1 port map( A1 => n27380, A2 => n20865, B => n13037, ZN => 
                           n13036);
   U8565 : NAND2_X1 port map( A1 => n13416, A2 => n10797, ZN => n1767);
   U3743 : NOR2_X1 port map( A1 => n21136, A2 => n20263, ZN => n21013);
   U8558 : NAND2_X1 port map( A1 => n3660, A2 => n15702, ZN => n3448);
   U6903 : NAND2_X1 port map( A1 => n10385, A2 => n22732, ZN => n10101);
   U4358 : INV_X1 port map( I => n2800, ZN => n721);
   U13 : OR2_X1 port map( A1 => n3042, A2 => n20911, Z => n2842);
   U21 : AND2_X1 port map( A1 => n21086, A2 => n6485, Z => n1338);
   U35 : AND2_X1 port map( A1 => n12251, A2 => n13888, Z => n21291);
   U39 : NAND2_X1 port map( A1 => n7039, A2 => n9494, ZN => n21213);
   U46 : INV_X1 port map( I => n20965, ZN => n1072);
   U71 : NOR2_X1 port map( A1 => n26146, A2 => n24929, ZN => n15313);
   U73 : AOI21_X1 port map( A1 => n23323, A2 => n20598, B => n28017, ZN => 
                           n20408);
   U86 : NOR2_X1 port map( A1 => n22484, A2 => n22483, ZN => n7645);
   U96 : NAND2_X1 port map( A1 => n11120, A2 => n10532, ZN => n25202);
   U101 : NAND2_X1 port map( A1 => n7772, A2 => n15103, ZN => n24924);
   U109 : NAND3_X1 port map( A1 => n4548, A2 => n950, A3 => n20881, ZN => 
                           n20884);
   U111 : INV_X1 port map( I => n4548, ZN => n25009);
   U114 : AND2_X1 port map( A1 => n9131, A2 => n14914, Z => n10809);
   U118 : INV_X1 port map( I => n21691, ZN => n11076);
   U129 : NAND2_X1 port map( A1 => n12309, A2 => n21099, ZN => n23371);
   U135 : CLKBUF_X2 port map( I => n20180, Z => n26156);
   U136 : AND2_X1 port map( A1 => n7807, A2 => n7518, Z => n24619);
   U142 : INV_X2 port map( I => n14334, ZN => n21664);
   U145 : NAND2_X1 port map( A1 => n24539, A2 => n5753, ZN => n8327);
   U152 : NAND2_X1 port map( A1 => n14281, A2 => n21395, ZN => n25277);
   U156 : NAND2_X1 port map( A1 => n13461, A2 => n10730, ZN => n26521);
   U168 : OR2_X1 port map( A1 => n23454, A2 => n20367, Z => n21579);
   U176 : BUF_X2 port map( I => n24331, Z => n12287);
   U179 : NOR2_X1 port map( A1 => n22227, A2 => n25239, ZN => n26477);
   U209 : INV_X1 port map( I => n21388, ZN => n24817);
   U214 : BUF_X2 port map( I => n22919, Z => n20881);
   U255 : NOR2_X1 port map( A1 => n11543, A2 => n11544, ZN => n26537);
   U258 : AND2_X1 port map( A1 => n8898, A2 => n20224, Z => n24676);
   U276 : NAND2_X1 port map( A1 => n23676, A2 => n13837, ZN => n24744);
   U288 : NAND3_X1 port map( A1 => n25012, A2 => n1106, A3 => n25011, ZN => 
                           n9560);
   U320 : NOR2_X1 port map( A1 => n4537, A2 => n21892, ZN => n680);
   U348 : NOR2_X1 port map( A1 => n20138, A2 => n3958, ZN => n26301);
   U349 : NAND2_X1 port map( A1 => n6264, A2 => n26252, ZN => n20040);
   U352 : AND2_X1 port map( A1 => n13719, A2 => n20043, Z => n10686);
   U365 : NAND3_X1 port map( A1 => n23065, A2 => n19962, A3 => n8300, ZN => 
                           n5029);
   U383 : INV_X1 port map( I => n12986, ZN => n23401);
   U391 : NAND2_X1 port map( A1 => n11048, A2 => n2525, ZN => n20187);
   U400 : NOR2_X1 port map( A1 => n27435, A2 => n10764, ZN => n15584);
   U404 : NOR2_X1 port map( A1 => n24998, A2 => n25934, ZN => n25076);
   U425 : OR2_X1 port map( A1 => n12895, A2 => n12893, Z => n25390);
   U435 : INV_X2 port map( I => n20131, ZN => n20318);
   U441 : NOR2_X1 port map( A1 => n25035, A2 => n9732, ZN => n224);
   U446 : OR2_X1 port map( A1 => n19677, A2 => n19846, Z => n10024);
   U471 : NAND2_X1 port map( A1 => n1348, A2 => n19097, ZN => n25035);
   U477 : AOI21_X1 port map( A1 => n26162, A2 => n19831, B => n14319, ZN => 
                           n9176);
   U490 : NAND2_X1 port map( A1 => n7376, A2 => n19603, ZN => n26162);
   U539 : NAND2_X1 port map( A1 => n15048, A2 => n25899, ZN => n25114);
   U553 : NOR2_X1 port map( A1 => n22140, A2 => n25279, ZN => n3431);
   U555 : NAND3_X1 port map( A1 => n19671, A2 => n24184, A3 => n329, ZN => 
                           n9156);
   U558 : OAI21_X1 port map( A1 => n11369, A2 => n19862, B => n4810, ZN => 
                           n25110);
   U565 : OAI21_X1 port map( A1 => n10272, A2 => n10557, B => n19766, ZN => 
                           n9814);
   U573 : AOI21_X1 port map( A1 => n19671, A2 => n24184, B => n10196, ZN => 
                           n9157);
   U580 : INV_X1 port map( I => n13194, ZN => n25279);
   U581 : AND2_X1 port map( A1 => n21788, A2 => n26354, Z => n11130);
   U611 : AND2_X1 port map( A1 => n10937, A2 => n3563, Z => n670);
   U615 : NAND2_X1 port map( A1 => n26535, A2 => n22744, ZN => n23380);
   U620 : NAND2_X1 port map( A1 => n19767, A2 => n19766, ZN => n12265);
   U632 : NAND2_X1 port map( A1 => n19889, A2 => n2223, ZN => n26527);
   U641 : OAI21_X1 port map( A1 => n19928, A2 => n26625, B => n9612, ZN => 
                           n26099);
   U647 : INV_X1 port map( I => n19890, ZN => n26528);
   U672 : NAND2_X1 port map( A1 => n19466, A2 => n19468, ZN => n26022);
   U709 : BUF_X2 port map( I => n22365, Z => n26447);
   U736 : CLKBUF_X2 port map( I => n12697, Z => n23572);
   U738 : INV_X1 port map( I => n12909, ZN => n26172);
   U740 : INV_X1 port map( I => n19521, ZN => n19563);
   U802 : NAND3_X1 port map( A1 => n23618, A2 => n11696, A3 => n18914, ZN => 
                           n18915);
   U816 : OR2_X1 port map( A1 => n23546, A2 => n11580, Z => n7567);
   U828 : OR2_X1 port map( A1 => n26641, A2 => n1164, Z => n24309);
   U841 : INV_X1 port map( I => n28547, ZN => n26607);
   U849 : CLKBUF_X2 port map( I => n8554, Z => n22260);
   U858 : AND2_X1 port map( A1 => n19057, A2 => n12571, Z => n1923);
   U863 : NAND2_X1 port map( A1 => n18876, A2 => n180, ZN => n12981);
   U866 : NOR2_X1 port map( A1 => n1163, A2 => n19191, ZN => n25201);
   U868 : NAND2_X1 port map( A1 => n24524, A2 => n28299, ZN => n26300);
   U869 : NAND2_X1 port map( A1 => n2247, A2 => n2245, ZN => n25381);
   U873 : INV_X2 port map( I => n13349, ZN => n15246);
   U881 : NOR2_X1 port map( A1 => n7030, A2 => n14098, ZN => n9554);
   U890 : NAND2_X1 port map( A1 => n19124, A2 => n2617, ZN => n2616);
   U898 : OR2_X1 port map( A1 => n4265, A2 => n14580, Z => n4264);
   U903 : AND2_X1 port map( A1 => n18376, A2 => n18375, Z => n25367);
   U912 : CLKBUF_X2 port map( I => n18947, Z => n26345);
   U970 : OAI22_X1 port map( A1 => n24608, A2 => n6512, B1 => n12724, B2 => 
                           n18475, ZN => n22290);
   U982 : NAND3_X1 port map( A1 => n22977, A2 => n18749, A3 => n18643, ZN => 
                           n10479);
   U987 : NAND2_X1 port map( A1 => n18387, A2 => n12979, ZN => n18388);
   U1013 : AOI21_X1 port map( A1 => n10642, A2 => n277, B => n23666, ZN => 
                           n24712);
   U1020 : NAND2_X1 port map( A1 => n24870, A2 => n18487, ZN => n18389);
   U1022 : NOR2_X1 port map( A1 => n18682, A2 => n18685, ZN => n26423);
   U1030 : AND2_X1 port map( A1 => n1015, A2 => n27241, Z => n24634);
   U1032 : BUF_X2 port map( I => n10564, Z => n7078);
   U1036 : NOR2_X1 port map( A1 => n18534, A2 => n1180, ZN => n6075);
   U1038 : NOR2_X1 port map( A1 => n18749, A2 => n18639, ZN => n24700);
   U1054 : INV_X1 port map( I => n18757, ZN => n26282);
   U1058 : NAND2_X1 port map( A1 => n12820, A2 => n18124, ZN => n24818);
   U1069 : OR2_X1 port map( A1 => n18557, A2 => n6014, Z => n8702);
   U1070 : NAND3_X1 port map( A1 => n18664, A2 => n18662, A3 => n24207, ZN => 
                           n3887);
   U1073 : NAND2_X1 port map( A1 => n737, A2 => n2912, ZN => n5457);
   U1079 : INV_X1 port map( I => n18534, ZN => n9784);
   U1094 : AOI21_X1 port map( A1 => n13192, A2 => n13191, B => n15660, ZN => 
                           n25705);
   U1114 : NAND2_X1 port map( A1 => n14376, A2 => n18639, ZN => n18745);
   U1120 : CLKBUF_X1 port map( I => n649, Z => n457);
   U1133 : NAND2_X1 port map( A1 => n18646, A2 => n27871, ZN => n9869);
   U1166 : CLKBUF_X2 port map( I => n2437, Z => n25651);
   U1174 : NAND2_X1 port map( A1 => n9328, A2 => n12371, ZN => n1371);
   U1188 : OR2_X1 port map( A1 => n12913, A2 => n12590, Z => n24624);
   U1240 : AND2_X1 port map( A1 => n7599, A2 => n1349, Z => n1771);
   U1242 : NAND2_X1 port map( A1 => n24969, A2 => n12087, ZN => n24946);
   U1272 : OAI21_X1 port map( A1 => n8365, A2 => n1780, B => n5584, ZN => n5583
                           );
   U1276 : AND2_X1 port map( A1 => n17867, A2 => n17868, Z => n13988);
   U1292 : AND2_X1 port map( A1 => n17607, A2 => n9485, Z => n11834);
   U1309 : BUF_X2 port map( I => n25679, Z => n25515);
   U1312 : INV_X2 port map( I => n1780, ZN => n12850);
   U1314 : OR2_X1 port map( A1 => n5402, A2 => n10673, Z => n14189);
   U1315 : NOR2_X1 port map( A1 => n12027, A2 => n763, ZN => n25200);
   U1321 : OAI21_X1 port map( A1 => n26437, A2 => n25724, B => n1213, ZN => 
                           n25885);
   U1322 : BUF_X2 port map( I => n17726, Z => n26610);
   U1331 : NAND2_X1 port map( A1 => n21768, A2 => n14278, ZN => n11770);
   U1341 : OAI21_X1 port map( A1 => n23563, A2 => n1966, B => n5096, ZN => 
                           n1965);
   U1347 : NAND2_X1 port map( A1 => n3620, A2 => n24613, ZN => n25466);
   U1354 : NOR2_X1 port map( A1 => n17472, A2 => n17244, ZN => n17151);
   U1356 : AOI22_X1 port map( A1 => n23449, A2 => n24612, B1 => n8661, B2 => 
                           n23777, ZN => n22704);
   U1357 : AOI21_X1 port map( A1 => n17187, A2 => n14532, B => n24214, ZN => 
                           n24775);
   U1360 : NAND2_X1 port map( A1 => n17192, A2 => n17175, ZN => n24686);
   U1363 : AOI21_X1 port map( A1 => n13358, A2 => n17335, B => n17565, ZN => 
                           n17184);
   U1384 : INV_X1 port map( I => n9481, ZN => n24688);
   U1393 : AND2_X1 port map( A1 => n14528, A2 => n12438, Z => n17280);
   U1395 : NAND2_X1 port map( A1 => n24517, A2 => n24406, ZN => n26191);
   U1403 : NOR2_X1 port map( A1 => n26226, A2 => n23105, ZN => n22979);
   U1410 : NAND2_X1 port map( A1 => n12455, A2 => n13568, ZN => n26500);
   U1413 : NAND2_X1 port map( A1 => n24517, A2 => n17381, ZN => n26362);
   U1415 : AND2_X1 port map( A1 => n9535, A2 => n7371, Z => n17248);
   U1424 : CLKBUF_X2 port map( I => n17532, Z => n12438);
   U1427 : NAND2_X1 port map( A1 => n23102, A2 => n17468, ZN => n195);
   U1432 : NAND2_X1 port map( A1 => n17515, A2 => n26616, ZN => n10298);
   U1445 : NAND2_X1 port map( A1 => n7912, A2 => n12225, ZN => n25057);
   U1446 : NOR2_X1 port map( A1 => n17381, A2 => n24335, ZN => n26361);
   U1465 : INV_X1 port map( I => n6707, ZN => n336);
   U1479 : NOR2_X1 port map( A1 => n145, A2 => n23236, ZN => n25723);
   U1481 : NOR2_X1 port map( A1 => n25670, A2 => n25554, ZN => n24856);
   U1487 : NAND2_X1 port map( A1 => n26114, A2 => n26113, ZN => n26112);
   U1490 : BUF_X2 port map( I => n16604, Z => n2131);
   U1492 : NAND2_X1 port map( A1 => n14656, A2 => n26244, ZN => n10514);
   U1499 : NOR2_X1 port map( A1 => n16533, A2 => n9830, ZN => n26593);
   U1510 : NOR2_X1 port map( A1 => n1257, A2 => n12117, ZN => n14820);
   U1512 : NOR2_X1 port map( A1 => n16530, A2 => n13964, ZN => n26293);
   U1516 : NOR2_X1 port map( A1 => n24952, A2 => n25415, ZN => n26489);
   U1517 : NAND3_X1 port map( A1 => n26108, A2 => n12949, A3 => n26107, ZN => 
                           n26111);
   U1519 : NOR2_X1 port map( A1 => n24648, A2 => n26298, ZN => n4449);
   U1524 : NAND2_X1 port map( A1 => n16585, A2 => n26244, ZN => n7114);
   U1527 : NOR2_X1 port map( A1 => n16598, A2 => n4555, ZN => n25010);
   U1530 : AOI21_X1 port map( A1 => n26853, A2 => n16438, B => n21809, ZN => 
                           n23780);
   U1532 : NAND2_X1 port map( A1 => n28083, A2 => n7265, ZN => n22715);
   U1536 : INV_X1 port map( I => n905, ZN => n26108);
   U1547 : INV_X1 port map( I => n25940, ZN => n26145);
   U1565 : NAND2_X1 port map( A1 => n15159, A2 => n16691, ZN => n5556);
   U1575 : NOR2_X1 port map( A1 => n905, A2 => n12726, ZN => n26113);
   U1590 : AND2_X1 port map( A1 => n12647, A2 => n16604, Z => n24644);
   U1602 : BUF_X2 port map( I => n14451, Z => n2390);
   U1608 : NAND2_X1 port map( A1 => n11503, A2 => n906, ZN => n26318);
   U1614 : NAND2_X1 port map( A1 => n4589, A2 => n23367, ZN => n10767);
   U1622 : NOR2_X1 port map( A1 => n22862, A2 => n16295, ZN => n25701);
   U1627 : NAND3_X1 port map( A1 => n16132, A2 => n15831, A3 => n25471, ZN => 
                           n15772);
   U1639 : NOR3_X1 port map( A1 => n26692, A2 => n14559, A3 => n16324, ZN => 
                           n25757);
   U1649 : OAI21_X1 port map( A1 => n4763, A2 => n16324, B => n16326, ZN => 
                           n25300);
   U1650 : NAND2_X1 port map( A1 => n2543, A2 => n9706, ZN => n9705);
   U1653 : AOI21_X1 port map( A1 => n799, A2 => n4532, B => n14415, ZN => n4378
                           );
   U1655 : OAI21_X1 port map( A1 => n9393, A2 => n21786, B => n24879, ZN => 
                           n9394);
   U1657 : NAND2_X1 port map( A1 => n7311, A2 => n16318, ZN => n13583);
   U1672 : NOR2_X1 port map( A1 => n4751, A2 => n10707, ZN => n25444);
   U1676 : AND2_X1 port map( A1 => n1721, A2 => n16063, Z => n24603);
   U1677 : NOR2_X1 port map( A1 => n16326, A2 => n15331, ZN => n25825);
   U1681 : NOR2_X1 port map( A1 => n1260, A2 => n12678, ZN => n22862);
   U1683 : INV_X1 port map( I => n16010, ZN => n16008);
   U1688 : NAND2_X1 port map( A1 => n9393, A2 => n10001, ZN => n24879);
   U1689 : NAND2_X1 port map( A1 => n7282, A2 => n16027, ZN => n24696);
   U1694 : NOR2_X1 port map( A1 => n14559, A2 => n10707, ZN => n25826);
   U1699 : AOI21_X1 port map( A1 => n795, A2 => n1263, B => n16106, ZN => 
                           n26134);
   U1703 : NAND2_X1 port map( A1 => n28032, A2 => n12678, ZN => n25917);
   U1705 : NAND2_X1 port map( A1 => n15947, A2 => n16320, ZN => n25464);
   U1708 : OAI21_X1 port map( A1 => n16130, A2 => n14386, B => n7235, ZN => 
                           n14910);
   U1709 : NAND2_X1 port map( A1 => n9223, A2 => n16107, ZN => n16059);
   U1713 : INV_X1 port map( I => n15989, ZN => n25599);
   U1722 : NAND2_X1 port map( A1 => n25764, A2 => n25763, ZN => n7472);
   U1730 : INV_X1 port map( I => n16258, ZN => n25764);
   U1753 : NAND2_X2 port map( A1 => n8534, A2 => n22838, ZN => n24839);
   U1769 : NAND2_X2 port map( A1 => n27359, A2 => n24175, ZN => n17720);
   U1771 : BUF_X2 port map( I => n11816, Z => n26051);
   U1779 : INV_X4 port map( I => n6998, ZN => n20129);
   U1788 : INV_X1 port map( I => n2506, ZN => n868);
   U1801 : NOR3_X2 port map( A1 => n15706, A2 => n1515, A3 => n21664, ZN => 
                           n25821);
   U1816 : OR2_X1 port map( A1 => n26647, A2 => n21734, Z => n9836);
   U1817 : NAND2_X2 port map( A1 => n22319, A2 => n7868, ZN => n11755);
   U1819 : BUF_X2 port map( I => n16306, Z => n13545);
   U1821 : INV_X2 port map( I => n17160, ZN => n17317);
   U1842 : NOR2_X1 port map( A1 => n13607, A2 => n17560, ZN => n10232);
   U1862 : NAND3_X1 port map( A1 => n20728, A2 => n20730, A3 => n24930, ZN => 
                           n3132);
   U1868 : OAI21_X1 port map( A1 => n27822, A2 => n12559, B => n20998, ZN => 
                           n1824);
   U1909 : INV_X1 port map( I => n10347, ZN => n73);
   U1926 : OAI22_X1 port map( A1 => n204, A2 => n14459, B1 => n4810, B2 => 
                           n12941, ZN => n6875);
   U1931 : INV_X1 port map( I => n26626, ZN => n361);
   U1942 : NOR3_X1 port map( A1 => n9378, A2 => n20180, A3 => n3559, ZN => 
                           n2213);
   U1943 : OAI21_X1 port map( A1 => n15471, A2 => n28095, B => n28134, ZN => 
                           n143);
   U1950 : INV_X1 port map( I => n21898, ZN => n24195);
   U1954 : NAND2_X1 port map( A1 => n21222, A2 => n21220, ZN => n24973);
   U1967 : AND2_X1 port map( A1 => n13056, A2 => n11318, Z => n12407);
   U1973 : NOR3_X1 port map( A1 => n28305, A2 => n1091, A3 => n4122, ZN => 
                           n8510);
   U1974 : NAND2_X1 port map( A1 => n3430, A2 => n23956, ZN => n6904);
   U1979 : CLKBUF_X2 port map( I => n7454, Z => n26462);
   U1980 : NAND2_X1 port map( A1 => n22218, A2 => n22668, ZN => n26133);
   U1993 : INV_X1 port map( I => n21087, ZN => n21081);
   U2005 : AND2_X1 port map( A1 => n5797, A2 => n15021, Z => n24626);
   U2014 : INV_X1 port map( I => n6508, ZN => n6794);
   U2026 : CLKBUF_X4 port map( I => n20365, Z => n21622);
   U2032 : AOI21_X1 port map( A1 => n3643, A2 => n21165, B => n3641, ZN => 
                           n3231);
   U2038 : OAI21_X1 port map( A1 => n12191, A2 => n21172, B => n4307, ZN => 
                           n3643);
   U2039 : INV_X2 port map( I => n17914, ZN => n17783);
   U2040 : BUF_X2 port map( I => n17914, Z => n13061);
   U2046 : NOR3_X1 port map( A1 => n1172, A2 => n7165, A3 => n7168, ZN => n7684
                           );
   U2056 : NAND3_X1 port map( A1 => n4984, A2 => n5005, A3 => n21409, ZN => 
                           n22574);
   U2064 : NAND3_X1 port map( A1 => n19700, A2 => n20137, A3 => n14235, ZN => 
                           n5854);
   U2065 : NAND2_X1 port map( A1 => n20137, A2 => n27129, ZN => n12563);
   U2072 : OR2_X1 port map( A1 => n13979, A2 => n21586, Z => n24224);
   U2085 : NOR2_X1 port map( A1 => n968, A2 => n14193, ZN => n14430);
   U2114 : NAND2_X1 port map( A1 => n8447, A2 => n20749, ZN => n8446);
   U2115 : OAI21_X1 port map( A1 => n12002, A2 => n23978, B => n27820, ZN => 
                           n13340);
   U2125 : NOR2_X1 port map( A1 => n12821, A2 => n24818, ZN => n12704);
   U2138 : NOR2_X1 port map( A1 => n4364, A2 => n19697, ZN => n26314);
   U2139 : NAND2_X1 port map( A1 => n9697, A2 => n10771, ZN => n1798);
   U2163 : OR2_X1 port map( A1 => n8982, A2 => n13642, Z => n1764);
   U2166 : INV_X1 port map( I => n13925, ZN => n19992);
   U2170 : INV_X1 port map( I => n22191, ZN => n25824);
   U2176 : NAND3_X1 port map( A1 => n1073, A2 => n20457, A3 => n20462, ZN => 
                           n26303);
   U2184 : NOR2_X1 port map( A1 => n3824, A2 => n2254, ZN => n20655);
   U2186 : NAND2_X1 port map( A1 => n25237, A2 => n25298, ZN => n24961);
   U2191 : NAND2_X1 port map( A1 => n16526, A2 => n16525, ZN => n8249);
   U2200 : BUF_X2 port map( I => n16526, Z => n14579);
   U2201 : INV_X1 port map( I => n16526, ZN => n6911);
   U2206 : OR2_X1 port map( A1 => n11044, A2 => n28121, Z => n10167);
   U2209 : NAND2_X1 port map( A1 => n21565, A2 => n7085, ZN => n12795);
   U2267 : NAND2_X1 port map( A1 => n9131, A2 => n11089, ZN => n25739);
   U2272 : NAND2_X1 port map( A1 => n27924, A2 => n20639, ZN => n24929);
   U2279 : INV_X1 port map( I => n9042, ZN => n8300);
   U2287 : AOI21_X1 port map( A1 => n26970, A2 => n11961, B => n5934, ZN => 
                           n3508);
   U2298 : NAND2_X1 port map( A1 => n13269, A2 => n3644, ZN => n4151);
   U2303 : NOR2_X1 port map( A1 => n22548, A2 => n22547, ZN => n22546);
   U2328 : OAI21_X1 port map( A1 => n24470, A2 => n7904, B => n21066, ZN => 
                           n25264);
   U2332 : OAI22_X1 port map( A1 => n8052, A2 => n8645, B1 => n8054, B2 => 
                           n24332, ZN => n2506);
   U2347 : INV_X1 port map( I => n18443, ZN => n18784);
   U2372 : BUF_X2 port map( I => n24568, Z => n23399);
   U2384 : AOI21_X1 port map( A1 => n12234, A2 => n14037, B => n2516, ZN => 
                           n19023);
   U2414 : NOR2_X1 port map( A1 => n24019, A2 => n875, ZN => n3178);
   U2422 : NOR2_X1 port map( A1 => n3801, A2 => n875, ZN => n26546);
   U2430 : CLKBUF_X2 port map( I => n23128, Z => n22296);
   U2432 : NOR2_X1 port map( A1 => n26226, A2 => n14917, ZN => n8380);
   U2446 : INV_X2 port map( I => n14578, ZN => n1234);
   U2449 : NOR2_X1 port map( A1 => n14578, A2 => n6870, ZN => n2502);
   U2451 : NOR2_X1 port map( A1 => n14578, A2 => n9879, ZN => n6196);
   U2466 : NAND2_X1 port map( A1 => n21061, A2 => n14341, ZN => n26221);
   U2468 : OAI21_X1 port map( A1 => n27734, A2 => n16694, B => n14676, ZN => 
                           n8632);
   U2484 : INV_X1 port map( I => n21695, ZN => n1091);
   U2491 : NAND2_X1 port map( A1 => n24646, A2 => n16619, ZN => n5122);
   U2503 : AND2_X1 port map( A1 => n16274, A2 => n11813, Z => n14764);
   U2533 : NAND2_X1 port map( A1 => n14900, A2 => n4472, ZN => n17374);
   U2536 : INV_X1 port map( I => n1975, ZN => n4304);
   U2537 : CLKBUF_X4 port map( I => n7281, Z => n23749);
   U2541 : NAND2_X1 port map( A1 => n9661, A2 => n8165, ZN => n17269);
   U2571 : AOI21_X1 port map( A1 => n17403, A2 => n14762, B => n10580, ZN => 
                           n17169);
   U2574 : NOR2_X1 port map( A1 => n14356, A2 => n5008, ZN => n9553);
   U2578 : INV_X1 port map( I => n19741, ZN => n14356);
   U2589 : AND2_X1 port map( A1 => n13049, A2 => n14795, Z => n14860);
   U2593 : AND2_X1 port map( A1 => n6763, A2 => n13794, Z => n12526);
   U2595 : INV_X1 port map( I => n13794, ZN => n16676);
   U2596 : BUF_X2 port map( I => n13351, Z => n6996);
   U2600 : CLKBUF_X2 port map( I => n25328, Z => n6652);
   U2604 : CLKBUF_X2 port map( I => n2179, Z => n458);
   U2615 : NAND2_X1 port map( A1 => n17605, A2 => n4719, ZN => n6644);
   U2622 : INV_X2 port map( I => n25922, ZN => n830);
   U2625 : NAND2_X1 port map( A1 => n25922, A2 => n4536, ZN => n17224);
   U2629 : AND2_X1 port map( A1 => n21644, A2 => n24381, Z => n15658);
   U2635 : NOR2_X1 port map( A1 => n10801, A2 => n10474, ZN => n23970);
   U2644 : OR3_X1 port map( A1 => n13794, A2 => n15652, A3 => n13548, Z => 
                           n6935);
   U2652 : INV_X1 port map( I => n18574, ZN => n18759);
   U2670 : INV_X2 port map( I => n17116, ZN => n17068);
   U2673 : AND2_X1 port map( A1 => n23236, A2 => n14562, Z => n24540);
   U2675 : INV_X2 port map( I => n17173, ZN => n2377);
   U2676 : AND2_X1 port map( A1 => n13530, A2 => n18003, Z => n24541);
   U2689 : INV_X2 port map( I => n15284, ZN => n280);
   U2691 : INV_X2 port map( I => n17532, ZN => n17478);
   U2692 : XNOR2_X1 port map( A1 => n18069, A2 => n18088, ZN => n24542);
   U2694 : AOI21_X2 port map( A1 => n6372, A2 => n13350, B => n6171, ZN => 
                           n25312);
   U2697 : CLKBUF_X4 port map( I => n18418, Z => n18750);
   U2698 : INV_X4 port map( I => n18750, ZN => n25828);
   U2699 : CLKBUF_X4 port map( I => n17891, Z => n18749);
   U2711 : INV_X1 port map( I => n22105, ZN => n19138);
   U2720 : AND2_X2 port map( A1 => n19913, A2 => n22842, Z => n24545);
   U2727 : INV_X2 port map( I => n10602, ZN => n20415);
   U2735 : NOR2_X2 port map( A1 => n6756, A2 => n10217, ZN => n25307);
   U2738 : NAND2_X2 port map( A1 => n21015, A2 => n21014, ZN => n25352);
   U2739 : NAND2_X2 port map( A1 => n21015, A2 => n21014, ZN => n9422);
   U2751 : OR2_X1 port map( A1 => n21345, A2 => n25753, Z => n24549);
   U2753 : NOR2_X2 port map( A1 => n14583, A2 => n13395, ZN => n25003);
   U2766 : NOR2_X1 port map( A1 => n3090, A2 => n15592, ZN => n26033);
   U2771 : NOR3_X2 port map( A1 => n10872, A2 => n27871, A3 => n21790, ZN => 
                           n25567);
   U2775 : AND3_X2 port map( A1 => n14284, A2 => n22307, A3 => n17869, Z => 
                           n22112);
   U2778 : NAND2_X1 port map( A1 => n4311, A2 => n20030, ZN => n20031);
   U2781 : AOI21_X2 port map( A1 => n21099, A2 => n12309, B => n1078, ZN => 
                           n12308);
   U2787 : INV_X2 port map( I => n9828, ZN => n9830);
   U2788 : BUF_X2 port map( I => n9828, Z => n8901);
   U2797 : AND2_X2 port map( A1 => n24458, A2 => n6853, Z => n10563);
   U2798 : NOR2_X1 port map( A1 => n26097, A2 => n10164, ZN => n26096);
   U2804 : INV_X1 port map( I => n21161, ZN => n21022);
   U2805 : NAND3_X1 port map( A1 => n13545, A2 => n15916, A3 => n1270, ZN => 
                           n3767);
   U2809 : INV_X1 port map( I => n2131, ZN => n4060);
   U2820 : OR2_X2 port map( A1 => n7940, A2 => n27467, Z => n21462);
   U2823 : INV_X1 port map( I => n14369, ZN => n11783);
   U2830 : OAI21_X1 port map( A1 => n13472, A2 => n21118, B => n11837, ZN => 
                           n11011);
   U2855 : OR2_X2 port map( A1 => n21667, A2 => n21668, Z => n12353);
   U2871 : NAND3_X1 port map( A1 => n27456, A2 => n22370, A3 => n797, ZN => 
                           n26142);
   U2881 : NAND2_X1 port map( A1 => n7910, A2 => n14893, ZN => n2331);
   U2882 : INV_X2 port map( I => n15662, ZN => n4020);
   U2884 : OAI22_X1 port map( A1 => n5923, A2 => n17867, B1 => n1028, B2 => 
                           n17770, ZN => n5922);
   U2893 : INV_X1 port map( I => n17867, ZN => n17770);
   U2904 : AND2_X2 port map( A1 => n14757, A2 => n7182, Z => n22710);
   U2916 : AOI22_X2 port map( A1 => n13376, A2 => n1004, B1 => n25051, B2 => 
                           n8792, ZN => n13375);
   U2921 : NOR2_X1 port map( A1 => n997, A2 => n27464, ZN => n18670);
   U2926 : INV_X1 port map( I => n22919, ZN => n20933);
   U2945 : CLKBUF_X12 port map( I => n13421, Z => n26243);
   U2949 : CLKBUF_X4 port map( I => n15884, Z => n16298);
   U2953 : INV_X1 port map( I => n19349, ZN => n26403);
   U2955 : BUF_X2 port map( I => n12708, Z => n5218);
   U2979 : NOR2_X1 port map( A1 => n17678, A2 => n25679, ZN => n4917);
   U2989 : INV_X2 port map( I => n1483, ZN => n14552);
   U3015 : NOR2_X1 port map( A1 => n18370, A2 => n18455, ZN => n18383);
   U3029 : OAI21_X1 port map( A1 => n21850, A2 => n9553, B => n24184, ZN => 
                           n22875);
   U3031 : NOR2_X1 port map( A1 => n2049, A2 => n12218, ZN => n2491);
   U3033 : AOI21_X1 port map( A1 => n845, A2 => n9460, B => n6802, ZN => n1693)
                           ;
   U3035 : OAI21_X1 port map( A1 => n188, A2 => n6802, B => n13718, ZN => n7998
                           );
   U3062 : AOI22_X1 port map( A1 => n1992, A2 => n4644, B1 => n15351, B2 => 
                           n1048, ZN => n1991);
   U3078 : OR2_X2 port map( A1 => n21754, A2 => n4888, Z => n17429);
   U3081 : NOR3_X1 port map( A1 => n16813, A2 => n12224, A3 => n4518, ZN => 
                           n23809);
   U3104 : NOR2_X1 port map( A1 => n4812, A2 => n17926, ZN => n3233);
   U3121 : INV_X1 port map( I => n17751, ZN => n17987);
   U3128 : CLKBUF_X12 port map( I => n14321, Z => n13968);
   U3139 : INV_X1 port map( I => n10241, ZN => n19877);
   U3147 : OAI22_X1 port map( A1 => n1646, A2 => n3297, B1 => n6683, B2 => 
                           n12039, ZN => n1645);
   U3152 : CLKBUF_X4 port map( I => n20469, Z => n21699);
   U3170 : NOR2_X1 port map( A1 => n8223, A2 => n905, ZN => n7648);
   U3175 : OAI21_X2 port map( A1 => n3693, A2 => n4118, B => n18956, ZN => 
                           n3150);
   U3179 : NOR2_X1 port map( A1 => n5310, A2 => n16224, ZN => n15351);
   U3192 : BUF_X4 port map( I => n6215, Z => n24998);
   U3201 : OAI22_X1 port map( A1 => n16603, A2 => n2131, B1 => n132, B2 => 
                           n7539, ZN => n16607);
   U3219 : AOI21_X1 port map( A1 => n19077, A2 => n19078, B => n12521, ZN => 
                           n6026);
   U3221 : AND2_X2 port map( A1 => n10574, A2 => n25346, Z => n7041);
   U3231 : NAND2_X1 port map( A1 => n18124, A2 => n1191, ZN => n14371);
   U3265 : NAND2_X1 port map( A1 => n13502, A2 => n11874, ZN => n8989);
   U3267 : NOR2_X2 port map( A1 => n9602, A2 => n9603, ZN => n22383);
   U3273 : NAND3_X1 port map( A1 => n11603, A2 => n1111, A3 => n10938, ZN => 
                           n6420);
   U3279 : OR2_X2 port map( A1 => n19850, A2 => n7240, Z => n5739);
   U3304 : NOR2_X2 port map( A1 => n9974, A2 => n15411, ZN => n9973);
   U3307 : CLKBUF_X12 port map( I => n14426, Z => n1629);
   U3312 : BUF_X2 port map( I => n965, Z => n24558);
   U3315 : INV_X1 port map( I => n16959, ZN => n24069);
   U3334 : AOI21_X2 port map( A1 => n10225, A2 => n1108, B => n23599, ZN => 
                           n10222);
   U3341 : NAND3_X1 port map( A1 => n24961, A2 => n3593, A3 => n9378, ZN => 
                           n14443);
   U3357 : INV_X1 port map( I => n21004, ZN => n21007);
   U3365 : INV_X1 port map( I => n17094, ZN => n25414);
   U3370 : NAND2_X1 port map( A1 => n15282, A2 => n10629, ZN => n16038);
   U3377 : INV_X1 port map( I => n13752, ZN => n19344);
   U3378 : NOR2_X1 port map( A1 => n22325, A2 => n18715, ZN => n8746);
   U3390 : NAND2_X1 port map( A1 => n6945, A2 => n18414, ZN => n5561);
   U3401 : OR2_X1 port map( A1 => n18947, A2 => n25339, Z => n14441);
   U3425 : OR2_X2 port map( A1 => n10542, A2 => n24329, Z => n8333);
   U3444 : NAND2_X1 port map( A1 => n11471, A2 => n968, ZN => n11470);
   U3445 : OAI21_X1 port map( A1 => n19544, A2 => n11471, B => n28134, ZN => 
                           n6429);
   U3446 : INV_X1 port map( I => n25439, ZN => n14950);
   U3448 : INV_X1 port map( I => n17869, ZN => n886);
   U3450 : OR2_X1 port map( A1 => n7321, A2 => n17869, Z => n5923);
   U3451 : NAND3_X1 port map( A1 => n1028, A2 => n17867, A3 => n17869, ZN => 
                           n24807);
   U3452 : OR2_X2 port map( A1 => n14748, A2 => n11628, Z => n4346);
   U3455 : AND2_X2 port map( A1 => n14748, A2 => n11628, Z => n16089);
   U3456 : BUF_X4 port map( I => n14748, Z => n22319);
   U3464 : NOR2_X1 port map( A1 => n26145, A2 => n479, ZN => n3949);
   U3465 : INV_X1 port map( I => n479, ZN => n1252);
   U3470 : NOR2_X1 port map( A1 => n479, A2 => n25940, ZN => n16423);
   U3492 : NAND2_X1 port map( A1 => n21111, A2 => n13009, ZN => n21107);
   U3494 : NOR2_X1 port map( A1 => n1035, A2 => n14528, ZN => n24980);
   U3510 : INV_X2 port map( I => n16685, ZN => n16687);
   U3511 : NAND2_X1 port map( A1 => n16685, A2 => n3792, ZN => n26032);
   U3537 : NAND2_X1 port map( A1 => n11223, A2 => n16335, ZN => n1546);
   U3547 : AOI22_X1 port map( A1 => n817, A2 => n5990, B1 => n27432, B2 => 
                           n27044, ZN => n5288);
   U3553 : BUF_X4 port map( I => n16629, Z => n25670);
   U3556 : NAND2_X1 port map( A1 => n23744, A2 => n16629, ZN => n14339);
   U3588 : AND3_X2 port map( A1 => n14759, A2 => n13772, A3 => n21395, Z => 
                           n21447);
   U3591 : OR2_X2 port map( A1 => n19913, A2 => n24558, Z => n1685);
   U3609 : OR2_X2 port map( A1 => n5391, A2 => n8793, Z => n8154);
   U3616 : INV_X2 port map( I => n12571, ZN => n26395);
   U3623 : NAND2_X1 port map( A1 => n16565, A2 => n10543, ZN => n10502);
   U3636 : NOR2_X1 port map( A1 => n16524, A2 => n16525, ZN => n16527);
   U3650 : NAND2_X1 port map( A1 => n28288, A2 => n1024, ZN => n8889);
   U3651 : INV_X1 port map( I => n3834, ZN => n18039);
   U3669 : OAI21_X1 port map( A1 => n7009, A2 => n696, B => n27390, ZN => 
                           n21645);
   U3670 : NOR2_X1 port map( A1 => n7009, A2 => n27390, ZN => n9850);
   U3675 : OR2_X1 port map( A1 => n6843, A2 => n6838, Z => n571);
   U3680 : NAND2_X1 port map( A1 => n6838, A2 => n10393, ZN => n5973);
   U3697 : NOR2_X1 port map( A1 => n21096, A2 => n20559, ZN => n15451);
   U3714 : AND2_X2 port map( A1 => n15892, A2 => n15891, Z => n16351);
   U3726 : INV_X1 port map( I => n10971, ZN => n3903);
   U3762 : CLKBUF_X4 port map( I => n561, Z => n7282);
   U3816 : NAND2_X1 port map( A1 => n21455, A2 => n27431, ZN => n13973);
   U3831 : AND3_X2 port map( A1 => n18741, A2 => n27737, A3 => n18739, Z => 
                           n18742);
   U3833 : INV_X1 port map( I => n21538, ZN => n21530);
   U3852 : CLKBUF_X12 port map( I => n17173, Z => n17347);
   U3860 : INV_X2 port map( I => n8181, ZN => n16563);
   U3861 : NOR2_X1 port map( A1 => n26578, A2 => n8181, ZN => n22378);
   U3871 : NOR2_X1 port map( A1 => n20917, A2 => n20911, ZN => n2838);
   U3873 : AND2_X2 port map( A1 => n8373, A2 => n14906, Z => n21891);
   U3911 : AOI21_X1 port map( A1 => n26234, A2 => n23488, B => n5363, ZN => 
                           n6836);
   U3931 : NAND2_X1 port map( A1 => n17869, A2 => n22202, ZN => n22305);
   U3933 : INV_X1 port map( I => n22738, ZN => n25963);
   U3937 : NAND2_X1 port map( A1 => n13188, A2 => n24575, ZN => n25750);
   U3938 : BUF_X2 port map( I => n20787, Z => n24575);
   U3943 : NOR2_X1 port map( A1 => n857, A2 => n7942, ZN => n20024);
   U3959 : AOI21_X1 port map( A1 => n15286, A2 => n26948, B => n26447, ZN => 
                           n24985);
   U3960 : AND2_X1 port map( A1 => n13110, A2 => n19872, Z => n24601);
   U3961 : NAND2_X1 port map( A1 => n19955, A2 => n19953, ZN => n25936);
   U3964 : NOR2_X1 port map( A1 => n19842, A2 => n3584, ZN => n24866);
   U3968 : BUF_X2 port map( I => n14595, Z => n26120);
   U3979 : NAND2_X1 port map( A1 => n18895, A2 => n18917, ZN => n2541);
   U3984 : INV_X2 port map( I => n2617, ZN => n19062);
   U4015 : INV_X4 port map( I => n2820, ZN => n24572);
   U4016 : CLKBUF_X1 port map( I => n2869, Z => n24019);
   U4027 : INV_X1 port map( I => n25705, ZN => n5586);
   U4030 : OAI21_X1 port map( A1 => n22832, A2 => n18662, B => n18722, ZN => 
                           n26215);
   U4040 : AOI21_X1 port map( A1 => n22482, A2 => n14375, B => n18748, ZN => 
                           n26064);
   U4056 : NAND2_X1 port map( A1 => n18747, A2 => n24701, ZN => n25082);
   U4063 : CLKBUF_X2 port map( I => n18569, Z => n14376);
   U4071 : INV_X1 port map( I => n1197, ZN => n13676);
   U4085 : NAND2_X1 port map( A1 => n26437, A2 => n17948, ZN => n25883);
   U4086 : OR2_X1 port map( A1 => n17795, A2 => n8882, Z => n24665);
   U4090 : NAND2_X1 port map( A1 => n7495, A2 => n14610, ZN => n25394);
   U4093 : NOR2_X1 port map( A1 => n7834, A2 => n12600, ZN => n25734);
   U4099 : NAND2_X1 port map( A1 => n6662, A2 => n6672, ZN => n26128);
   U4106 : AND2_X1 port map( A1 => n23797, A2 => n14990, Z => n15222);
   U4110 : NOR2_X1 port map( A1 => n13623, A2 => n791, ZN => n25871);
   U4113 : BUF_X4 port map( I => n15317, Z => n4536);
   U4117 : CLKBUF_X1 port map( I => n10431, Z => n25983);
   U4126 : INV_X1 port map( I => n16918, ZN => n24968);
   U4136 : BUF_X4 port map( I => n10337, Z => n25772);
   U4138 : BUF_X2 port map( I => n16497, Z => n22660);
   U4143 : AND2_X1 port map( A1 => n15787, A2 => n25373, Z => n4763);
   U4146 : AOI21_X1 port map( A1 => n3298, A2 => n7022, B => n25171, ZN => 
                           n25170);
   U4151 : BUF_X2 port map( I => n16021, Z => n26350);
   U4155 : INV_X2 port map( I => n14224, ZN => n25135);
   U4162 : NAND2_X1 port map( A1 => n25134, A2 => n5847, ZN => n21294);
   U4168 : NOR2_X1 port map( A1 => n11820, A2 => n6051, ZN => n6054);
   U4179 : NAND2_X1 port map( A1 => n21293, A2 => n21292, ZN => n25134);
   U4182 : NAND2_X1 port map( A1 => n8559, A2 => n4767, ZN => n8558);
   U4190 : NAND2_X1 port map( A1 => n929, A2 => n21107, ZN => n5221);
   U4194 : INV_X1 port map( I => n9563, ZN => n24853);
   U4199 : NOR2_X1 port map( A1 => n1338, A2 => n13476, ZN => n25953);
   U4200 : NAND2_X1 port map( A1 => n21348, A2 => n21340, ZN => n2452);
   U4201 : INV_X2 port map( I => n21340, ZN => n21344);
   U4212 : NOR2_X1 port map( A1 => n21659, A2 => n6181, ZN => n21656);
   U4219 : OR2_X1 port map( A1 => n6727, A2 => n6728, Z => n25378);
   U4222 : CLKBUF_X2 port map( I => n21083, Z => n26157);
   U4225 : NAND2_X1 port map( A1 => n26220, A2 => n21096, ZN => n26219);
   U4227 : NAND2_X1 port map( A1 => n12098, A2 => n12097, ZN => n25460);
   U4229 : NAND2_X1 port map( A1 => n21069, A2 => n25264, ZN => n15479);
   U4231 : INV_X4 port map( I => n24225, ZN => n24574);
   U4274 : INV_X2 port map( I => n21389, ZN => n26554);
   U4289 : CLKBUF_X2 port map( I => n24680, Z => n8751);
   U4290 : BUF_X2 port map( I => n3895, Z => n22737);
   U4291 : BUF_X4 port map( I => n20935, Z => n950);
   U4292 : OR2_X1 port map( A1 => n7706, A2 => n3462, Z => n5071);
   U4319 : INV_X2 port map( I => n20581, ZN => n24577);
   U4368 : NAND2_X1 port map( A1 => n13255, A2 => n24590, ZN => n25695);
   U4409 : NAND2_X1 port map( A1 => n807, A2 => n24989, ZN => n24988);
   U4420 : OAI21_X1 port map( A1 => n7122, A2 => n8898, B => n20226, ZN => 
                           n24833);
   U4442 : AND2_X1 port map( A1 => n25455, A2 => n9167, Z => n514);
   U4448 : INV_X1 port map( I => n10356, ZN => n26270);
   U4450 : INV_X2 port map( I => n19999, ZN => n20219);
   U4461 : INV_X1 port map( I => n4021, ZN => n25056);
   U4467 : INV_X2 port map( I => n11947, ZN => n25710);
   U4470 : CLKBUF_X2 port map( I => n14221, Z => n24394);
   U4474 : INV_X1 port map( I => n10344, ZN => n26201);
   U4479 : INV_X1 port map( I => n24985, ZN => n24984);
   U4486 : NAND2_X1 port map( A1 => n19467, A2 => n26021, ZN => n26020);
   U4488 : NAND2_X1 port map( A1 => n19738, A2 => n19876, ZN => n26130);
   U4492 : NAND2_X1 port map( A1 => n26099, A2 => n9813, ZN => n15049);
   U4493 : NAND2_X1 port map( A1 => n19604, A2 => n27730, ZN => n26543);
   U4504 : INV_X1 port map( I => n19620, ZN => n26126);
   U4526 : INV_X2 port map( I => n1460, ZN => n19800);
   U4538 : AOI21_X1 port map( A1 => n15575, A2 => n19877, B => n14307, ZN => 
                           n15521);
   U4540 : NAND2_X1 port map( A1 => n24866, A2 => n14307, ZN => n26399);
   U4549 : INV_X1 port map( I => n19922, ZN => n24820);
   U4550 : CLKBUF_X2 port map( I => n19899, Z => n25230);
   U4551 : NAND2_X1 port map( A1 => n4364, A2 => n19697, ZN => n26023);
   U4558 : BUF_X1 port map( I => n10601, Z => n26061);
   U4564 : INV_X4 port map( I => n11805, ZN => n24579);
   U4591 : INV_X1 port map( I => n25545, ZN => n25544);
   U4593 : NAND2_X1 port map( A1 => n21756, A2 => n14719, ZN => n24883);
   U4610 : NAND2_X1 port map( A1 => n22115, A2 => n24489, ZN => n252);
   U4616 : NOR2_X1 port map( A1 => n22566, A2 => n11117, ZN => n25090);
   U4617 : NOR2_X1 port map( A1 => n8248, A2 => n4224, ZN => n25732);
   U4640 : NOR2_X1 port map( A1 => n994, A2 => n25201, ZN => n5459);
   U4648 : NAND2_X1 port map( A1 => n19038, A2 => n19037, ZN => n7657);
   U4678 : CLKBUF_X2 port map( I => n14162, Z => n24188);
   U4681 : INV_X2 port map( I => n22626, ZN => n24937);
   U4687 : INV_X1 port map( I => n19155, ZN => n22882);
   U4688 : NAND2_X1 port map( A1 => n19163, A2 => n8611, ZN => n5247);
   U4703 : INV_X1 port map( I => n26215, ZN => n26214);
   U4709 : NAND2_X1 port map( A1 => n26283, A2 => n26282, ZN => n26281);
   U4719 : INV_X1 port map( I => n18756, ZN => n26283);
   U4720 : INV_X1 port map( I => n26064, ZN => n13940);
   U4743 : NOR2_X1 port map( A1 => n18714, A2 => n6800, ZN => n6767);
   U4744 : OR2_X1 port map( A1 => n12569, A2 => n15623, Z => n24608);
   U4745 : INV_X1 port map( I => n18783, ZN => n26072);
   U4790 : INV_X1 port map( I => n18745, ZN => n12998);
   U4815 : BUF_X2 port map( I => n18578, Z => n12573);
   U4818 : AND2_X1 port map( A1 => n8855, A2 => n25349, Z => n3416);
   U4824 : NOR2_X1 port map( A1 => n14362, A2 => n18570, ZN => n24699);
   U4834 : BUF_X2 port map( I => n18579, Z => n23062);
   U4837 : INV_X2 port map( I => n6549, ZN => n18455);
   U4838 : CLKBUF_X2 port map( I => n18642, Z => n24701);
   U4899 : BUF_X2 port map( I => n2704, Z => n2873);
   U4907 : INV_X1 port map( I => n23950, ZN => n25677);
   U4910 : CLKBUF_X4 port map( I => n4559, Z => n26486);
   U4916 : NAND2_X1 port map( A1 => n25884, A2 => n25883, ZN => n17698);
   U4919 : NOR2_X1 port map( A1 => n25395, A2 => n25394, ZN => n25393);
   U4938 : INV_X1 port map( I => n25885, ZN => n25884);
   U4944 : INV_X1 port map( I => n7497, ZN => n25395);
   U4954 : OAI21_X1 port map( A1 => n15390, A2 => n25734, B => n17648, ZN => 
                           n9211);
   U4955 : NOR2_X1 port map( A1 => n25578, A2 => n17797, ZN => n17201);
   U4957 : NAND2_X1 port map( A1 => n6965, A2 => n6964, ZN => n17961);
   U4958 : OR2_X1 port map( A1 => n23064, A2 => n7358, Z => n15534);
   U4960 : OR2_X1 port map( A1 => n4319, A2 => n23064, Z => n12731);
   U4964 : CLKBUF_X2 port map( I => n23231, Z => n26387);
   U4966 : NAND2_X1 port map( A1 => n827, A2 => n6709, ZN => n25578);
   U4985 : CLKBUF_X2 port map( I => n17653, Z => n24003);
   U4998 : INV_X1 port map( I => n25214, ZN => n25492);
   U5000 : NAND2_X1 port map( A1 => n17968, A2 => n11112, ZN => n6590);
   U5003 : NAND2_X1 port map( A1 => n5844, A2 => n26195, ZN => n17551);
   U5007 : INV_X2 port map( I => n4110, ZN => n25926);
   U5027 : NOR2_X1 port map( A1 => n22498, A2 => n24688, ZN => n24687);
   U5030 : NOR2_X1 port map( A1 => n24878, A2 => n24017, ZN => n24705);
   U5033 : NAND2_X1 port map( A1 => n10461, A2 => n25672, ZN => n8749);
   U5040 : OAI21_X1 port map( A1 => n26260, A2 => n26259, B => n13623, ZN => 
                           n14688);
   U5049 : NOR2_X1 port map( A1 => n23777, A2 => n25605, ZN => n11296);
   U5053 : NAND2_X1 port map( A1 => n7155, A2 => n11284, ZN => n25180);
   U5061 : NAND3_X1 port map( A1 => n17443, A2 => n10183, A3 => n17268, ZN => 
                           n23600);
   U5062 : AND2_X1 port map( A1 => n17546, A2 => n24234, Z => n12455);
   U5067 : OAI21_X1 port map( A1 => n17565, A2 => n13230, B => n16972, ZN => 
                           n25928);
   U5069 : INV_X1 port map( I => n11270, ZN => n17511);
   U5108 : AND2_X1 port map( A1 => n10539, A2 => n13358, Z => n24620);
   U5109 : BUF_X2 port map( I => n14533, Z => n23956);
   U5116 : BUF_X2 port map( I => n3300, Z => n24335);
   U5126 : INV_X1 port map( I => n16785, ZN => n25410);
   U5136 : CLKBUF_X2 port map( I => n16895, Z => n25582);
   U5144 : CLKBUF_X2 port map( I => n26576, Z => n24740);
   U5160 : INV_X1 port map( I => n14866, ZN => n23918);
   U5162 : NOR2_X1 port map( A1 => n3144, A2 => n7047, ZN => n25740);
   U5165 : INV_X1 port map( I => n1564, ZN => n26368);
   U5188 : NAND2_X1 port map( A1 => n2754, A2 => n24215, ZN => n24868);
   U5191 : NAND2_X1 port map( A1 => n162, A2 => n4630, ZN => n25441);
   U5197 : NAND2_X1 port map( A1 => n22587, A2 => n15420, ZN => n25938);
   U5200 : NOR2_X1 port map( A1 => n9605, A2 => n7758, ZN => n26307);
   U5203 : AND2_X1 port map( A1 => n16507, A2 => n1793, Z => n24657);
   U5205 : INV_X1 port map( I => n2038, ZN => n26124);
   U5208 : NAND2_X1 port map( A1 => n15421, A2 => n16467, ZN => n25939);
   U5218 : BUF_X2 port map( I => n6843, Z => n24334);
   U5220 : INV_X4 port map( I => n16654, ZN => n24580);
   U5223 : BUF_X4 port map( I => n2788, Z => n24089);
   U5224 : INV_X1 port map( I => n13039, ZN => n11122);
   U5227 : INV_X2 port map( I => n12839, ZN => n25834);
   U5228 : INV_X1 port map( I => n13815, ZN => n16175);
   U5238 : NAND2_X1 port map( A1 => n23946, A2 => n379, ZN => n25451);
   U5243 : NAND2_X1 port map( A1 => n25479, A2 => n25478, ZN => n25477);
   U5244 : NAND2_X1 port map( A1 => n16299, A2 => n25170, ZN => n12761);
   U5245 : NAND2_X1 port map( A1 => n26134, A2 => n2495, ZN => n2496);
   U5247 : INV_X1 port map( I => n7472, ZN => n16233);
   U5248 : AOI21_X1 port map( A1 => n16299, A2 => n11568, B => n23525, ZN => 
                           n26373);
   U5249 : NOR2_X1 port map( A1 => n21822, A2 => n24247, ZN => n26075);
   U5250 : NAND2_X1 port map( A1 => n14384, A2 => n10270, ZN => n26116);
   U5258 : NAND2_X1 port map( A1 => n15134, A2 => n15135, ZN => n26115);
   U5264 : OR2_X1 port map( A1 => n16039, A2 => n7152, Z => n10652);
   U5266 : INV_X1 port map( I => n5464, ZN => n15955);
   U5272 : INV_X1 port map( I => n16301, ZN => n25171);
   U5273 : OR2_X1 port map( A1 => n10970, A2 => n15889, Z => n24591);
   U5276 : CLKBUF_X2 port map( I => n21876, Z => n25570);
   U5277 : CLKBUF_X2 port map( I => n16068, Z => n24872);
   U5298 : INV_X2 port map( I => n16123, ZN => n6237);
   U5300 : NOR2_X1 port map( A1 => n6647, A2 => n1987, ZN => n5312);
   U5301 : NAND2_X1 port map( A1 => n16189, A2 => n16301, ZN => n14831);
   U5304 : CLKBUF_X2 port map( I => n16088, Z => n24702);
   U5305 : CLKBUF_X1 port map( I => n8648, Z => n8647);
   U5307 : NOR2_X1 port map( A1 => n13123, A2 => n16063, ZN => n1720);
   U5309 : OR2_X1 port map( A1 => n16203, A2 => n25365, Z => n10882);
   U5314 : CLKBUF_X2 port map( I => n12529, Z => n25224);
   U5315 : AOI21_X1 port map( A1 => n7282, A2 => n24581, B => n8647, ZN => 
                           n16200);
   U5319 : OAI21_X1 port map( A1 => n15994, A2 => n6236, B => n13731, ZN => 
                           n6235);
   U5328 : NOR2_X1 port map( A1 => n15895, A2 => n16339, ZN => n25660);
   U5331 : NAND2_X1 port map( A1 => n23457, A2 => n799, ZN => n23456);
   U5332 : CLKBUF_X2 port map( I => n4485, Z => n26371);
   U5341 : CLKBUF_X4 port map( I => n22991, Z => n16106);
   U5347 : NAND3_X1 port map( A1 => n16041, A2 => n16292, A3 => n12678, ZN => 
                           n16043);
   U5350 : BUF_X2 port map( I => n15881, Z => n16193);
   U5352 : AOI21_X1 port map( A1 => n798, A2 => n769, B => n14385, ZN => n22150
                           );
   U5353 : NAND3_X1 port map( A1 => n16106, A2 => n1259, A3 => n250, ZN => 
                           n7818);
   U5365 : INV_X2 port map( I => n13964, ZN => n1042);
   U5370 : AOI22_X1 port map( A1 => n2283, A2 => n730, B1 => n13877, B2 => 
                           n16196, ZN => n2282);
   U5371 : NOR2_X1 port map( A1 => n14942, A2 => n16241, ZN => n10504);
   U5377 : NOR2_X1 port map( A1 => n9763, A2 => n7631, ZN => n7650);
   U5380 : INV_X1 port map( I => n16704, ZN => n834);
   U5391 : OAI22_X1 port map( A1 => n6898, A2 => n23107, B1 => n6763, B2 => 
                           n15652, ZN => n4756);
   U5395 : NAND2_X1 port map( A1 => n14682, A2 => n16171, ZN => n16172);
   U5412 : NAND2_X1 port map( A1 => n7688, A2 => n24952, ZN => n13047);
   U5418 : NAND2_X1 port map( A1 => n15701, A2 => n16728, ZN => n8340);
   U5421 : OR2_X1 port map( A1 => n3399, A2 => n16679, Z => n24604);
   U5422 : CLKBUF_X2 port map( I => n12482, Z => n25287);
   U5440 : CLKBUF_X2 port map( I => n5861, Z => n25973);
   U5447 : NAND4_X1 port map( A1 => n10192, A2 => n10193, A3 => n11599, A4 => 
                           n11600, ZN => n9533);
   U5455 : NAND2_X1 port map( A1 => n22436, A2 => n16598, ZN => n12876);
   U5458 : INV_X2 port map( I => n16746, ZN => n17098);
   U5459 : AOI22_X1 port map( A1 => n2658, A2 => n13211, B1 => n16490, B2 => 
                           n27381, ZN => n15972);
   U5461 : CLKBUF_X2 port map( I => n16823, Z => n24077);
   U5467 : OAI21_X1 port map( A1 => n3218, A2 => n16405, B => n16638, ZN => 
                           n16032);
   U5471 : CLKBUF_X4 port map( I => n5379, Z => n23750);
   U5474 : NOR2_X1 port map( A1 => n17363, A2 => n25922, ZN => n3838);
   U5486 : NOR2_X1 port map( A1 => n4832, A2 => n25506, ZN => n23604);
   U5510 : NAND2_X1 port map( A1 => n21942, A2 => n12438, ZN => n26195);
   U5524 : AOI21_X1 port map( A1 => n17507, A2 => n17508, B => n17509, ZN => 
                           n7451);
   U5526 : NOR2_X1 port map( A1 => n17525, A2 => n791, ZN => n26260);
   U5557 : NAND3_X1 port map( A1 => n6022, A2 => n898, A3 => n1227, ZN => n327)
                           ;
   U5568 : NAND2_X1 port map( A1 => n17004, A2 => n17005, ZN => n22092);
   U5581 : OAI21_X1 port map( A1 => n892, A2 => n6021, B => n8094, ZN => n8175)
                           ;
   U5608 : NAND3_X1 port map( A1 => n2403, A2 => n826, A3 => n17842, ZN => 
                           n1906);
   U5612 : NAND2_X1 port map( A1 => n25215, A2 => n6681, ZN => n22289);
   U5636 : AND2_X1 port map( A1 => n5920, A2 => n4100, Z => n24661);
   U5638 : NAND2_X1 port map( A1 => n7492, A2 => n25393, ZN => n10890);
   U5649 : INV_X1 port map( I => n18310, ZN => n25143);
   U5656 : INV_X1 port map( I => n18319, ZN => n9144);
   U5681 : OAI21_X1 port map( A1 => n11783, A2 => n482, B => n1191, ZN => 
                           n18515);
   U5682 : INV_X1 port map( I => n18685, ZN => n25680);
   U5684 : NAND2_X1 port map( A1 => n23004, A2 => n15448, ZN => n15449);
   U5688 : NAND2_X1 port map( A1 => n11617, A2 => n18728, ZN => n10215);
   U5699 : NAND2_X1 port map( A1 => n27453, A2 => n18728, ZN => n2948);
   U5701 : INV_X2 port map( I => n5835, ZN => n14649);
   U5703 : NOR2_X1 port map( A1 => n22547, A2 => n18532, ZN => n15460);
   U5707 : NOR2_X1 port map( A1 => n7769, A2 => n6968, ZN => n15131);
   U5711 : NAND2_X1 port map( A1 => n18515, A2 => n18516, ZN => n1380);
   U5722 : OAI21_X1 port map( A1 => n14510, A2 => n1018, B => n14427, ZN => 
                           n22073);
   U5734 : INV_X1 port map( I => n14065, ZN => n18610);
   U5737 : NAND2_X1 port map( A1 => n12048, A2 => n15693, ZN => n7730);
   U5738 : OAI21_X1 port map( A1 => n15137, A2 => n4639, B => n18585, ZN => 
                           n13796);
   U5759 : INV_X2 port map( I => n6598, ZN => n10083);
   U5766 : NAND3_X1 port map( A1 => n26395, A2 => n18396, A3 => n19057, ZN => 
                           n18398);
   U5780 : NAND3_X1 port map( A1 => n3009, A2 => n5877, A3 => n6145, ZN => 
                           n19048);
   U5786 : INV_X1 port map( I => n5877, ZN => n13629);
   U5795 : NAND2_X1 port map( A1 => n10801, A2 => n2398, ZN => n24730);
   U5810 : AOI21_X1 port map( A1 => n23161, A2 => n19160, B => n9922, ZN => 
                           n2816);
   U5816 : NOR2_X1 port map( A1 => n26327, A2 => n19121, ZN => n14181);
   U5847 : NAND2_X1 port map( A1 => n18852, A2 => n25411, ZN => n25543);
   U5848 : OAI21_X1 port map( A1 => n22649, A2 => n26720, B => n22648, ZN => 
                           n18478);
   U5852 : NAND2_X1 port map( A1 => n2701, A2 => n18904, ZN => n25621);
   U5856 : AOI22_X1 port map( A1 => n11981, A2 => n27279, B1 => n3275, B2 => 
                           n22338, ZN => n11613);
   U5863 : INV_X2 port map( I => n19290, ZN => n982);
   U5876 : INV_X1 port map( I => n19314, ZN => n24925);
   U5881 : NOR2_X1 port map( A1 => n19672, A2 => n2941, ZN => n19580);
   U5905 : NAND2_X1 port map( A1 => n19922, A2 => n669, ZN => n26208);
   U5909 : INV_X1 port map( I => n19882, ZN => n975);
   U5925 : OAI21_X1 port map( A1 => n19888, A2 => n19681, B => n19890, ZN => 
                           n2214);
   U5926 : NOR2_X1 port map( A1 => n15265, A2 => n19907, ZN => n23887);
   U5929 : NOR2_X1 port map( A1 => n1118, A2 => n19801, ZN => n3654);
   U5931 : INV_X1 port map( I => n11205, ZN => n12690);
   U5940 : NOR2_X1 port map( A1 => n865, A2 => n5008, ZN => n19885);
   U5946 : NAND2_X1 port map( A1 => n11369, A2 => n4810, ZN => n11329);
   U5948 : OR2_X1 port map( A1 => n19575, A2 => n19914, Z => n11303);
   U5965 : CLKBUF_X4 port map( I => n6219, Z => n3317);
   U5975 : NAND3_X1 port map( A1 => n19903, A2 => n24109, A3 => n26654, ZN => 
                           n19911);
   U5980 : INV_X1 port map( I => n20029, ZN => n22622);
   U5981 : INV_X1 port map( I => n19692, ZN => n19948);
   U5987 : NOR2_X1 port map( A1 => n9042, A2 => n11215, ZN => n1756);
   U5988 : NOR2_X1 port map( A1 => n12757, A2 => n13925, ZN => n12755);
   U5989 : NAND3_X1 port map( A1 => n23229, A2 => n25340, A3 => n23906, ZN => 
                           n10898);
   U6014 : INV_X1 port map( I => n21104, ZN => n25980);
   U6020 : NAND2_X1 port map( A1 => n24989, A2 => n20165, ZN => n19934);
   U6026 : OAI21_X1 port map( A1 => n19992, A2 => n20430, B => n20089, ZN => 
                           n26556);
   U6030 : AOI21_X1 port map( A1 => n19992, A2 => n1580, B => n26556, ZN => 
                           n26555);
   U6052 : INV_X1 port map( I => n13680, ZN => n20579);
   U6056 : NAND2_X1 port map( A1 => n26651, A2 => n6547, ZN => n11689);
   U6059 : INV_X1 port map( I => n13505, ZN => n24930);
   U6068 : INV_X1 port map( I => n21324, ZN => n23251);
   U6074 : NAND2_X1 port map( A1 => n690, A2 => n10314, ZN => n5781);
   U6085 : NAND2_X1 port map( A1 => n13050, A2 => n23036, ZN => n11902);
   U6087 : OAI21_X1 port map( A1 => n14914, A2 => n24978, B => n21278, ZN => 
                           n12098);
   U6094 : NOR2_X1 port map( A1 => n22823, A2 => n6547, ZN => n21360);
   U6097 : NAND2_X1 port map( A1 => n26156, A2 => n26290, ZN => n2415);
   U6098 : INV_X1 port map( I => n21668, ZN => n21571);
   U6102 : INV_X1 port map( I => n13291, ZN => n25064);
   U6111 : NOR2_X1 port map( A1 => n1547, A2 => n844, ZN => n11440);
   U6115 : AOI21_X1 port map( A1 => n5673, A2 => n21666, B => n21571, ZN => 
                           n26586);
   U6117 : NOR2_X1 port map( A1 => n26462, A2 => n11522, ZN => n15125);
   U6122 : INV_X1 port map( I => n6181, ZN => n10173);
   U6123 : NAND2_X1 port map( A1 => n15125, A2 => n24763, ZN => n15124);
   U6127 : INV_X1 port map( I => n21174, ZN => n21165);
   U6139 : INV_X1 port map( I => n14609, ZN => n1292);
   U6142 : BUF_X2 port map( I => Key(173), Z => n21454);
   U6146 : AND2_X2 port map( A1 => n11374, A2 => n16515, Z => n24583);
   U6148 : XNOR2_X1 port map( A1 => n4877, A2 => n14589, ZN => n24584);
   U6149 : XNOR2_X1 port map( A1 => n575, A2 => n16955, ZN => n24585);
   U6151 : INV_X1 port map( I => n5353, ZN => n24507);
   U6153 : AND2_X1 port map( A1 => n16140, A2 => n15686, Z => n24588);
   U6155 : NAND3_X1 port map( A1 => n19697, A2 => n1121, A3 => n19782, ZN => 
                           n24589);
   U6158 : XNOR2_X1 port map( A1 => n12094, A2 => n21453, ZN => n24592);
   U6159 : XNOR2_X1 port map( A1 => n16747, A2 => n13738, ZN => n24593);
   U6162 : XNOR2_X1 port map( A1 => n21311, A2 => n13285, ZN => n24595);
   U6166 : AND2_X2 port map( A1 => n2622, A2 => n22522, Z => n24597);
   U6167 : OR2_X1 port map( A1 => n1990, A2 => n11694, Z => n24598);
   U6176 : OR2_X1 port map( A1 => n20049, A2 => n2023, Z => n24606);
   U6179 : AND3_X1 port map( A1 => n18785, A2 => n15227, A3 => n7087, Z => 
                           n24610);
   U6187 : NOR2_X1 port map( A1 => n14997, A2 => n27826, ZN => n24612);
   U6195 : AND3_X2 port map( A1 => n3857, A2 => n3856, A3 => n16468, Z => 
                           n24614);
   U6196 : AND2_X1 port map( A1 => n4914, A2 => n17713, Z => n24615);
   U6198 : OR2_X1 port map( A1 => n13673, A2 => n27161, Z => n24616);
   U6199 : AND2_X1 port map( A1 => n6522, A2 => n852, Z => n24617);
   U6203 : XNOR2_X1 port map( A1 => n23750, A2 => n14535, ZN => n24618);
   U6204 : AND2_X1 port map( A1 => n5009, A2 => n14679, Z => n24621);
   U6205 : BUF_X4 port map( I => n25854, Z => n25697);
   U6214 : AND2_X1 port map( A1 => n13572, A2 => n23842, Z => n24627);
   U6216 : NOR2_X1 port map( A1 => n12125, A2 => n15887, ZN => n24628);
   U6217 : CLKBUF_X4 port map( I => n11947, Z => n25254);
   U6219 : OR2_X2 port map( A1 => n19156, A2 => n5393, Z => n24630);
   U6221 : CLKBUF_X4 port map( I => n15934, Z => n1269);
   U6224 : AND2_X1 port map( A1 => n19759, A2 => n14279, Z => n24632);
   U6225 : AND2_X1 port map( A1 => n11331, A2 => n19015, Z => n24633);
   U6226 : AND3_X1 port map( A1 => n10385, A2 => n22732, A3 => n24574, Z => 
                           n24635);
   U6230 : INV_X1 port map( I => n1637, ZN => n1881);
   U6236 : INV_X1 port map( I => n3850, ZN => n15610);
   U6243 : AND2_X1 port map( A1 => n25843, A2 => n14221, Z => n24642);
   U6244 : INV_X1 port map( I => n16707, ZN => n26107);
   U6260 : INV_X2 port map( I => n27454, ZN => n745);
   U6262 : OR2_X2 port map( A1 => n15804, A2 => n15805, Z => n24646);
   U6264 : AND2_X2 port map( A1 => n13548, A2 => n13794, Z => n24648);
   U6265 : XOR2_X1 port map( A1 => n10049, A2 => n10047, Z => n24649);
   U6269 : XNOR2_X1 port map( A1 => n16924, A2 => n21288, ZN => n24651);
   U6273 : XNOR2_X1 port map( A1 => n28013, A2 => n14593, ZN => n24652);
   U6274 : AND3_X1 port map( A1 => n17922, A2 => n14397, A3 => n17921, Z => 
                           n24653);
   U6275 : XNOR2_X1 port map( A1 => n5481, A2 => n13450, ZN => n24654);
   U6286 : INV_X1 port map( I => n18579, ZN => n759);
   U6290 : XOR2_X1 port map( A1 => n18182, A2 => n21106, Z => n24658);
   U6302 : CLKBUF_X4 port map( I => n645, Z => n1177);
   U6312 : INV_X1 port map( I => n6870, ZN => n17313);
   U6313 : XNOR2_X1 port map( A1 => n18236, A2 => n11687, ZN => n24662);
   U6318 : XNOR2_X1 port map( A1 => n6123, A2 => n14473, ZN => n24663);
   U6329 : XNOR2_X1 port map( A1 => n19305, A2 => n20208, ZN => n24667);
   U6340 : CLKBUF_X4 port map( I => n16942, Z => n17513);
   U6343 : NOR2_X1 port map( A1 => n8838, A2 => n22845, ZN => n24670);
   U6353 : XNOR2_X1 port map( A1 => n5024, A2 => n5020, ZN => n24672);
   U6354 : CLKBUF_X4 port map( I => n19916, Z => n14459);
   U6356 : XNOR2_X1 port map( A1 => n19194, A2 => n1316, ZN => n24673);
   U6367 : INV_X1 port map( I => n24743, ZN => n3057);
   U6369 : NOR2_X1 port map( A1 => n6047, A2 => n25536, ZN => n24679);
   U6372 : XOR2_X1 port map( A1 => n25925, A2 => n21430, Z => n24680);
   U6378 : INV_X1 port map( I => n6860, ZN => n9377);
   U6379 : CLKBUF_X2 port map( I => n6860, Z => n3559);
   U6386 : XOR2_X1 port map( A1 => n18245, A2 => n24681, Z => n25296);
   U6388 : XOR2_X1 port map( A1 => n25865, A2 => n24682, Z => n24681);
   U6390 : INV_X1 port map( I => n21384, ZN => n24682);
   U6392 : NAND4_X1 port map( A1 => n9579, A2 => n19724, A3 => n20155, A4 => 
                           n19723, ZN => n1643);
   U6393 : NOR2_X2 port map( A1 => n2561, A2 => n24684, ZN => n15777);
   U6394 : NOR2_X1 port map( A1 => n2560, A2 => n16335, ZN => n24684);
   U6395 : NAND2_X1 port map( A1 => n15653, A2 => n15657, ZN => n7059);
   U6401 : AOI21_X2 port map( A1 => n6050, A2 => n15107, B => n6049, ZN => 
                           n17133);
   U6408 : XOR2_X1 port map( A1 => n18144, A2 => n4559, Z => n25105);
   U6409 : NAND2_X2 port map( A1 => n8182, A2 => n8185, ZN => n18144);
   U6418 : XOR2_X1 port map( A1 => n2902, A2 => n2903, Z => n2711);
   U6419 : XOR2_X1 port map( A1 => n1192, A2 => n3777, Z => n25813);
   U6427 : OAI21_X1 port map( A1 => n18566, A2 => n18495, B => n18653, ZN => 
                           n9273);
   U6437 : AND2_X1 port map( A1 => n18953, A2 => n736, Z => n9237);
   U6440 : NOR3_X1 port map( A1 => n647, A2 => n7212, A3 => n23399, ZN => 
                           n18422);
   U6441 : NOR2_X2 port map( A1 => n24691, A2 => n13652, ZN => n5537);
   U6444 : OAI21_X2 port map( A1 => n25621, A2 => n9346, B => n18905, ZN => 
                           n19285);
   U6451 : XOR2_X1 port map( A1 => n13906, A2 => n21712, Z => n6158);
   U6454 : NAND3_X2 port map( A1 => n3316, A2 => n3315, A3 => n18451, ZN => 
                           n13906);
   U6466 : BUF_X2 port map( I => n25176, Z => n24693);
   U6470 : NAND2_X2 port map( A1 => n24350, A2 => n10895, ZN => n22774);
   U6471 : AOI22_X2 port map( A1 => n8974, A2 => n23696, B1 => n12104, B2 => 
                           n26356, ZN => n24350);
   U6478 : NAND2_X1 port map( A1 => n3212, A2 => n13522, ZN => n22779);
   U6487 : AOI22_X1 port map( A1 => n12115, A2 => n16127, B1 => n12116, B2 => 
                           n263, ZN => n15870);
   U6491 : XOR2_X1 port map( A1 => n20361, A2 => n8072, Z => n2554);
   U6506 : NAND2_X1 port map( A1 => n15920, A2 => n8834, ZN => n24697);
   U6519 : OAI22_X2 port map( A1 => n13076, A2 => n20105, B1 => n25063, B2 => 
                           n13864, ZN => n21374);
   U6535 : NOR2_X2 port map( A1 => n24700, A2 => n24699, ZN => n26309);
   U6538 : XOR2_X1 port map( A1 => n4659, A2 => n11844, Z => n11843);
   U6547 : XOR2_X1 port map( A1 => n26246, A2 => n16817, Z => n4659);
   U6548 : XOR2_X1 port map( A1 => n24703, A2 => n23463, Z => n24954);
   U6554 : XOR2_X1 port map( A1 => n21237, A2 => n24955, Z => n24703);
   U6555 : NOR2_X1 port map( A1 => n8834, A2 => n25804, ZN => n16030);
   U6564 : XOR2_X1 port map( A1 => n16981, A2 => n26084, Z => n24193);
   U6574 : NOR2_X2 port map( A1 => n24705, A2 => n23151, ZN => n341);
   U6599 : NOR2_X2 port map( A1 => n1029, A2 => n17326, ZN => n24706);
   U6617 : OR2_X1 port map( A1 => n17495, A2 => n24308, Z => n22650);
   U6623 : NAND2_X2 port map( A1 => n8846, A2 => n8845, ZN => n16943);
   U6624 : NAND2_X1 port map( A1 => n25049, A2 => n5713, ZN => n24710);
   U6630 : XOR2_X1 port map( A1 => n18270, A2 => n24711, Z => n21911);
   U6635 : INV_X1 port map( I => n14575, ZN => n24711);
   U6645 : AOI21_X2 port map( A1 => n18651, A2 => n785, B => n24712, ZN => 
                           n19091);
   U6646 : NAND2_X1 port map( A1 => n65, A2 => n67, ZN => n25074);
   U6648 : OAI21_X2 port map( A1 => n12997, A2 => n12998, B => n18749, ZN => 
                           n25563);
   U6659 : NAND2_X2 port map( A1 => n23957, A2 => n24414, ZN => n16915);
   U6671 : NOR2_X1 port map( A1 => n20800, A2 => n10050, ZN => n24714);
   U6699 : NAND2_X2 port map( A1 => n15331, A2 => n14326, ZN => n15943);
   U6700 : XOR2_X1 port map( A1 => n18299, A2 => n17811, Z => n13850);
   U6704 : OAI22_X2 port map( A1 => n17773, A2 => n17584, B1 => n17928, B2 => 
                           n17742, ZN => n25496);
   U6705 : NAND2_X2 port map( A1 => n4813, A2 => n17924, ZN => n17742);
   U6706 : OR2_X2 port map( A1 => n25266, A2 => n10573, Z => n15975);
   U6710 : XOR2_X1 port map( A1 => n1198, A2 => n18221, Z => n18208);
   U6717 : XOR2_X1 port map( A1 => n19276, A2 => n19172, Z => n1944);
   U6721 : AOI22_X2 port map( A1 => n22977, A2 => n18497, B1 => n14362, B2 => 
                           n28090, ZN => n13939);
   U6726 : NAND2_X2 port map( A1 => n21845, A2 => n2906, ZN => n19201);
   U6732 : XOR2_X1 port map( A1 => n25747, A2 => n6291, Z => n10605);
   U6733 : NOR2_X1 port map( A1 => n20165, A2 => n24862, ZN => n23993);
   U6746 : XOR2_X1 port map( A1 => n25950, A2 => n24718, Z => n23420);
   U6748 : XOR2_X1 port map( A1 => n22846, A2 => n24673, Z => n24718);
   U6765 : AND2_X1 port map( A1 => n19110, A2 => n1156, Z => n19112);
   U6810 : BUF_X4 port map( I => n11077, Z => n24720);
   U6844 : NAND3_X2 port map( A1 => n24725, A2 => n17465, A3 => n17466, ZN => 
                           n21898);
   U6858 : NAND3_X1 port map( A1 => n17461, A2 => n17462, A3 => n14357, ZN => 
                           n24725);
   U6879 : INV_X2 port map( I => n11733, ZN => n24727);
   U6884 : NOR2_X2 port map( A1 => n3029, A2 => n16001, ZN => n3553);
   U6886 : INV_X2 port map( I => n24728, ZN => n6185);
   U6890 : XOR2_X1 port map( A1 => n24729, A2 => n18293, Z => n25038);
   U6891 : XOR2_X1 port map( A1 => n10917, A2 => n22879, Z => n24729);
   U6900 : NOR2_X2 port map( A1 => n9021, A2 => n17506, ZN => n9722);
   U6910 : NAND3_X2 port map( A1 => n10449, A2 => n9457, A3 => n14776, ZN => 
                           n9021);
   U6914 : AND2_X1 port map( A1 => n16159, A2 => n14425, Z => n16112);
   U6924 : XOR2_X1 port map( A1 => n2850, A2 => n6104, Z => n16922);
   U6925 : NAND2_X2 port map( A1 => n15296, A2 => n26590, ZN => n6104);
   U6928 : AOI22_X1 port map( A1 => n11751, A2 => n102, B1 => n8544, B2 => 
                           n4277, ZN => n8543);
   U6929 : OAI22_X2 port map( A1 => n120, A2 => n2061, B1 => n25670, B2 => n729
                           , ZN => n16988);
   U6937 : XOR2_X1 port map( A1 => n24732, A2 => n8649, Z => n22446);
   U6940 : XOR2_X1 port map( A1 => n28541, A2 => n18230, Z => n24732);
   U6954 : NOR3_X1 port map( A1 => n18445, A2 => n25585, A3 => n5407, ZN => 
                           n5211);
   U6958 : XNOR2_X1 port map( A1 => n20514, A2 => n19818, ZN => n25075);
   U6960 : INV_X2 port map( I => n24735, ZN => n7169);
   U6968 : XOR2_X1 port map( A1 => n17045, A2 => n10387, Z => n9841);
   U6970 : XOR2_X1 port map( A1 => n16823, A2 => n12626, Z => n17045);
   U6985 : AOI21_X2 port map( A1 => n2161, A2 => n21729, B => n11076, ZN => 
                           n2160);
   U6999 : NAND2_X2 port map( A1 => n13994, A2 => n24738, ZN => n21644);
   U7018 : XOR2_X1 port map( A1 => n16747, A2 => n24739, Z => n16510);
   U7020 : INV_X2 port map( I => n17147, ZN => n24739);
   U7027 : AOI21_X2 port map( A1 => n5730, A2 => n11495, B => n16408, ZN => 
                           n16747);
   U7028 : NAND2_X1 port map( A1 => n22681, A2 => n22799, ZN => n2136);
   U7034 : INV_X2 port map( I => n9117, ZN => n25914);
   U7035 : OR2_X1 port map( A1 => n4486, A2 => n23391, Z => n17834);
   U7045 : XOR2_X1 port map( A1 => n21151, A2 => n22340, Z => n24741);
   U7047 : INV_X2 port map( I => n24742, ZN => n10209);
   U7050 : XNOR2_X1 port map( A1 => n2124, A2 => n2123, ZN => n24742);
   U7057 : XOR2_X1 port map( A1 => n22159, A2 => n22158, Z => n17369);
   U7061 : NAND4_X2 port map( A1 => n3405, A2 => n7406, A3 => n14012, A4 => 
                           n7407, ZN => n11775);
   U7073 : XOR2_X1 port map( A1 => n18190, A2 => n24592, Z => n26037);
   U7079 : XOR2_X1 port map( A1 => n20250, A2 => n20423, Z => n23014);
   U7082 : NAND3_X2 port map( A1 => n25712, A2 => n1012, A3 => n737, ZN => 
                           n2245);
   U7093 : XOR2_X1 port map( A1 => n13351, A2 => n7399, Z => n2771);
   U7096 : NAND2_X2 port map( A1 => n24797, A2 => n3534, ZN => n13351);
   U7097 : AOI21_X2 port map( A1 => n6542, A2 => n9728, B => n24747, ZN => 
                           n6543);
   U7098 : AOI21_X2 port map( A1 => n6243, A2 => n9648, B => n1081, ZN => 
                           n24747);
   U7104 : XOR2_X1 port map( A1 => n3613, A2 => n9722, Z => n18278);
   U7111 : XOR2_X1 port map( A1 => n14551, A2 => n24108, Z => n8486);
   U7123 : NAND2_X2 port map( A1 => n13769, A2 => n10844, ZN => n12784);
   U7141 : NOR2_X1 port map( A1 => n21004, A2 => n3725, ZN => n3723);
   U7142 : NAND2_X1 port map( A1 => n3921, A2 => n740, ZN => n8528);
   U7143 : NAND2_X1 port map( A1 => n24750, A2 => n5133, ZN => n3852);
   U7144 : NAND2_X1 port map( A1 => n22680, A2 => n22681, ZN => n24750);
   U7147 : NOR2_X2 port map( A1 => n17179, A2 => n24752, ZN => n17470);
   U7159 : XOR2_X1 port map( A1 => n5420, A2 => n11552, Z => n22196);
   U7160 : NOR2_X2 port map( A1 => n24865, A2 => n6026, ZN => n5420);
   U7162 : XOR2_X1 port map( A1 => n24754, A2 => n1296, Z => Ciphertext(122));
   U7165 : OAI22_X1 port map( A1 => n26412, A2 => n14080, B1 => n14078, B2 => 
                           n14079, ZN => n24754);
   U7173 : OR2_X1 port map( A1 => n15985, A2 => n15984, Z => n24772);
   U7178 : AOI21_X2 port map( A1 => n3524, A2 => n10894, B => n24756, ZN => 
                           n4028);
   U7211 : XOR2_X1 port map( A1 => n24761, A2 => n3219, Z => n3746);
   U7212 : XOR2_X1 port map( A1 => n15456, A2 => n3748, Z => n24761);
   U7222 : OR2_X1 port map( A1 => n21111, A2 => n13009, Z => n24763);
   U7256 : NAND2_X1 port map( A1 => n24798, A2 => n26898, ZN => n24797);
   U7261 : NAND2_X1 port map( A1 => n23213, A2 => n1074, ZN => n25424);
   U7275 : NAND2_X1 port map( A1 => n14639, A2 => n17173, ZN => n6370);
   U7281 : NOR2_X2 port map( A1 => n24771, A2 => n15521, ZN => n20288);
   U7291 : NAND2_X2 port map( A1 => n24773, A2 => n24772, ZN => n13815);
   U7293 : AOI22_X1 port map( A1 => n21109, A2 => n11751, B1 => n13013, B2 => 
                           n102, ZN => n13012);
   U7295 : NOR2_X2 port map( A1 => n12699, A2 => n25363, ZN => n18476);
   U7307 : NOR2_X2 port map( A1 => n24791, A2 => n24775, ZN => n23245);
   U7341 : NOR2_X2 port map( A1 => n24883, A2 => n24602, ZN => n19194);
   U7346 : NAND2_X2 port map( A1 => n5126, A2 => n5125, ZN => n4970);
   U7347 : AND3_X1 port map( A1 => n4486, A2 => n4414, A3 => n23391, Z => 
                           n14706);
   U7348 : XOR2_X1 port map( A1 => n23359, A2 => n13008, Z => n13007);
   U7351 : OAI21_X2 port map( A1 => n4690, A2 => n9730, B => n5746, ZN => 
                           n10840);
   U7359 : INV_X2 port map( I => n3470, ZN => n3979);
   U7392 : NAND2_X2 port map( A1 => n12317, A2 => n10295, ZN => n10294);
   U7397 : NAND3_X2 port map( A1 => n6693, A2 => n6692, A3 => n26970, ZN => 
                           n5609);
   U7415 : AND2_X1 port map( A1 => n13267, A2 => n20135, Z => n22783);
   U7418 : OAI21_X2 port map( A1 => n3610, A2 => n656, B => n14188, ZN => n3609
                           );
   U7429 : NAND2_X2 port map( A1 => n16218, A2 => n11325, ZN => n24783);
   U7432 : XOR2_X1 port map( A1 => n16899, A2 => n16510, Z => n22711);
   U7434 : INV_X2 port map( I => n9508, ZN => n25712);
   U7437 : XOR2_X1 port map( A1 => n20577, A2 => n20576, Z => n2273);
   U7441 : XOR2_X1 port map( A1 => n2292, A2 => n9049, Z => n20576);
   U7443 : XOR2_X1 port map( A1 => n17073, A2 => n17074, Z => n17075);
   U7450 : INV_X2 port map( I => n9381, ZN => n20314);
   U7451 : NAND3_X2 port map( A1 => n9382, A2 => n25511, A3 => n7196, ZN => 
                           n9381);
   U7460 : OR2_X1 port map( A1 => n7602, A2 => n7601, Z => n3414);
   U7464 : NOR2_X1 port map( A1 => n19606, A2 => n11421, ZN => n11420);
   U7469 : NOR2_X2 port map( A1 => n11300, A2 => n5115, ZN => n12736);
   U7473 : NAND2_X2 port map( A1 => n1729, A2 => n1727, ZN => n7562);
   U7481 : INV_X2 port map( I => n20146, ZN => n856);
   U7487 : NOR2_X2 port map( A1 => n24785, A2 => n12621, ZN => n17759);
   U7488 : INV_X4 port map( I => n6185, ZN => n3533);
   U7490 : XOR2_X1 port map( A1 => n19347, A2 => n19348, Z => n11247);
   U7492 : NAND2_X2 port map( A1 => n22913, A2 => n1834, ZN => n19347);
   U7494 : NAND2_X2 port map( A1 => n5999, A2 => n24786, ZN => n7257);
   U7503 : XOR2_X1 port map( A1 => n452, A2 => n17028, Z => n4051);
   U7506 : NAND2_X2 port map( A1 => n24787, A2 => n23098, ZN => n7388);
   U7508 : INV_X2 port map( I => n24788, ZN => n11114);
   U7510 : XOR2_X1 port map( A1 => n16909, A2 => n21890, Z => n11002);
   U7527 : XOR2_X1 port map( A1 => n24166, A2 => n17090, Z => n16909);
   U7528 : XOR2_X1 port map( A1 => n19374, A2 => n19219, Z => n3007);
   U7537 : OAI21_X2 port map( A1 => n13202, A2 => n15673, B => n22127, ZN => 
                           n1772);
   U7539 : XOR2_X1 port map( A1 => n6959, A2 => n19180, Z => n3437);
   U7548 : XOR2_X1 port map( A1 => n15661, A2 => n19353, Z => n24111);
   U7549 : XOR2_X1 port map( A1 => n23117, A2 => n8322, Z => n19353);
   U7550 : INV_X4 port map( I => n1163, ZN => n25894);
   U7551 : NAND3_X1 port map( A1 => n11459, A2 => n11456, A3 => n11457, ZN => 
                           n437);
   U7552 : NAND2_X2 port map( A1 => n1104, A2 => n4274, ZN => n7942);
   U7560 : NOR2_X2 port map( A1 => n7330, A2 => n7518, ZN => n12140);
   U7576 : NAND2_X2 port map( A1 => n24867, A2 => n23741, ZN => n24790);
   U7589 : NAND3_X2 port map( A1 => n21133, A2 => n25947, A3 => n21131, ZN => 
                           n21174);
   U7590 : XOR2_X1 port map( A1 => n19248, A2 => n24793, Z => n23608);
   U7591 : XOR2_X1 port map( A1 => n19507, A2 => n24794, Z => n24793);
   U7592 : XOR2_X1 port map( A1 => n6554, A2 => n18125, Z => n18086);
   U7599 : NOR2_X1 port map( A1 => n26384, A2 => n24795, ZN => n6007);
   U7611 : NAND3_X2 port map( A1 => n9644, A2 => n19809, A3 => n25081, ZN => 
                           n24800);
   U7613 : BUF_X2 port map( I => n4034, Z => n24801);
   U7614 : AOI21_X2 port map( A1 => n26686, A2 => n8735, B => n24802, ZN => 
                           n9692);
   U7618 : NOR2_X2 port map( A1 => n21579, A2 => n8735, ZN => n24802);
   U7645 : AOI22_X2 port map( A1 => n12217, A2 => n23145, B1 => n975, B2 => 
                           n966, ZN => n2170);
   U7647 : OAI21_X1 port map( A1 => n10845, A2 => n23245, B => n1214, ZN => 
                           n17350);
   U7651 : XOR2_X1 port map( A1 => n17067, A2 => n24593, Z => n24805);
   U7652 : NOR2_X1 port map( A1 => n21716, A2 => n6046, ZN => n21717);
   U7659 : XOR2_X1 port map( A1 => n7653, A2 => n7654, Z => n9702);
   U7668 : INV_X2 port map( I => n8102, ZN => n24806);
   U7680 : XOR2_X1 port map( A1 => n13918, A2 => n658, Z => n19404);
   U7682 : NOR2_X2 port map( A1 => n252, A2 => n251, ZN => n658);
   U7689 : XOR2_X1 port map( A1 => n17109, A2 => n16965, Z => n16987);
   U7694 : NOR3_X2 port map( A1 => n19087, A2 => n19086, A3 => n25770, ZN => 
                           n8121);
   U7701 : NAND2_X2 port map( A1 => n10868, A2 => n3443, ZN => n16467);
   U7709 : INV_X2 port map( I => n24810, ZN => n14886);
   U7713 : XOR2_X1 port map( A1 => Plaintext(90), A2 => Key(90), Z => n24810);
   U7714 : INV_X4 port map( I => n24811, ZN => n11982);
   U7720 : NOR3_X1 port map( A1 => n10205, A2 => n18828, A3 => n25102, ZN => 
                           n24813);
   U7727 : XOR2_X1 port map( A1 => n521, A2 => n7130, Z => n24814);
   U7729 : NAND2_X2 port map( A1 => n1749, A2 => n24815, ZN => n16883);
   U7731 : NOR2_X1 port map( A1 => n1746, A2 => n1748, ZN => n24815);
   U7741 : XOR2_X1 port map( A1 => n21431, A2 => n25943, Z => n25948);
   U7743 : OAI21_X1 port map( A1 => n10197, A2 => n28428, B => n21332, ZN => 
                           n1739);
   U7747 : OAI21_X2 port map( A1 => n2642, A2 => n2641, B => n16392, ZN => 
                           n17035);
   U7759 : OR2_X1 port map( A1 => n632, A2 => n6779, Z => n10025);
   U7768 : OAI22_X1 port map( A1 => n17417, A2 => n3091, B1 => n17418, B2 => 
                           n3090, ZN => n3095);
   U7769 : INV_X2 port map( I => n3389, ZN => n3090);
   U7776 : NAND2_X2 port map( A1 => n15345, A2 => n13986, ZN => n21451);
   U7808 : AND2_X1 port map( A1 => n16005, A2 => n16006, Z => n14198);
   U7830 : BUF_X2 port map( I => n2788, Z => n24829);
   U7837 : NOR2_X2 port map( A1 => n16579, A2 => n3564, ZN => n22050);
   U7840 : OAI21_X2 port map( A1 => n20746, A2 => n953, B => n24830, ZN => 
                           n6589);
   U7845 : NAND2_X1 port map( A1 => n12890, A2 => n18971, ZN => n12889);
   U7847 : NAND2_X2 port map( A1 => n24831, A2 => n24835, ZN => n21087);
   U7849 : XOR2_X1 port map( A1 => n24832, A2 => n8316, Z => n23284);
   U7850 : XOR2_X1 port map( A1 => n9214, A2 => n26550, Z => n24832);
   U7852 : XOR2_X1 port map( A1 => n23834, A2 => n12522, Z => n13475);
   U7855 : OAI21_X1 port map( A1 => n24676, A2 => n20226, B => n24833, ZN => 
                           n20231);
   U7856 : NOR2_X1 port map( A1 => n7834, A2 => n7298, ZN => n1570);
   U7857 : NOR2_X1 port map( A1 => n20181, A2 => n13719, ZN => n20182);
   U7868 : NOR2_X2 port map( A1 => n2639, A2 => n23191, ZN => n5351);
   U7873 : NOR2_X2 port map( A1 => n25336, A2 => n16630, ZN => n2038);
   U7881 : NAND2_X2 port map( A1 => n2591, A2 => n2590, ZN => n25336);
   U7892 : NAND2_X2 port map( A1 => n11761, A2 => n10942, ZN => n17482);
   U7895 : NAND2_X2 port map( A1 => n24834, A2 => n23477, ZN => n19804);
   U7897 : OAI21_X2 port map( A1 => n27881, A2 => n11936, B => n1459, ZN => 
                           n24834);
   U7899 : NOR2_X1 port map( A1 => n13424, A2 => n22616, ZN => n12296);
   U7911 : AND2_X1 port map( A1 => n756, A2 => n19899, Z => n23296);
   U7917 : INV_X1 port map( I => n13043, ZN => n25106);
   U7923 : XOR2_X1 port map( A1 => n12909, A2 => n12910, Z => n12908);
   U7940 : XOR2_X1 port map( A1 => n22774, A2 => n24840, Z => n25093);
   U7945 : INV_X1 port map( I => n21602, ZN => n24840);
   U7949 : NAND4_X2 port map( A1 => n24842, A2 => n16356, A3 => n16358, A4 => 
                           n24841, ZN => n18002);
   U7953 : NAND2_X1 port map( A1 => n12496, A2 => n1232, ZN => n24842);
   U7957 : XOR2_X1 port map( A1 => n19288, A2 => n19287, Z => n24843);
   U7961 : INV_X2 port map( I => n16699, ZN => n24844);
   U7966 : AOI21_X2 port map( A1 => n14863, A2 => n2814, B => n10355, ZN => 
                           n17617);
   U7973 : INV_X1 port map( I => n13181, ZN => n24846);
   U7987 : OAI21_X2 port map( A1 => n10809, A2 => n10621, B => n21328, ZN => 
                           n24849);
   U8009 : NAND2_X1 port map( A1 => n8388, A2 => n9563, ZN => n24851);
   U8010 : AOI21_X1 port map( A1 => n24853, A2 => n934, B => n27429, ZN => 
                           n24852);
   U8018 : OAI21_X1 port map( A1 => n2307, A2 => n14583, B => n1068, ZN => 
                           n20583);
   U8023 : AOI21_X2 port map( A1 => n6073, A2 => n6074, B => n18372, ZN => 
                           n25514);
   U8029 : NOR2_X2 port map( A1 => n28378, A2 => n19683, ZN => n25910);
   U8031 : NAND3_X1 port map( A1 => n480, A2 => n3759, A3 => n20693, ZN => 
                           n2937);
   U8039 : XOR2_X1 port map( A1 => n3005, A2 => n23279, Z => n3003);
   U8040 : OAI21_X2 port map( A1 => n24868, A2 => n24856, B => n6611, ZN => 
                           n2265);
   U8058 : XOR2_X1 port map( A1 => n24858, A2 => n21104, Z => Ciphertext(90));
   U8067 : OAI21_X2 port map( A1 => n6064, A2 => n15812, B => n24859, ZN => 
                           n6858);
   U8071 : NAND3_X2 port map( A1 => n5050, A2 => n15812, A3 => n25225, ZN => 
                           n24859);
   U8074 : OR2_X1 port map( A1 => n21538, A2 => n12625, Z => n9577);
   U8079 : MUX2_X1 port map( I0 => n14352, I1 => n6052, S => n20751, Z => 
                           n20745);
   U8082 : NAND2_X2 port map( A1 => n10086, A2 => n10087, ZN => n20751);
   U8091 : INV_X2 port map( I => n23687, ZN => n9056);
   U8104 : OAI21_X2 port map( A1 => n628, A2 => n1905, B => n24863, ZN => n7951
                           );
   U8115 : OAI22_X2 port map( A1 => n19074, A2 => n987, B1 => n19075, B2 => 
                           n14791, ZN => n24865);
   U8123 : NAND2_X1 port map( A1 => n12465, A2 => n20979, ZN => n25692);
   U8128 : XOR2_X1 port map( A1 => n18276, A2 => n18275, Z => n9552);
   U8135 : XOR2_X1 port map( A1 => n18211, A2 => n18135, Z => n18275);
   U8152 : NAND2_X2 port map( A1 => n21496, A2 => n21495, ZN => n24867);
   U8198 : INV_X2 port map( I => n21342, ZN => n24874);
   U8208 : NAND2_X2 port map( A1 => n1738, A2 => n1737, ZN => n21340);
   U8218 : NOR2_X1 port map( A1 => n2238, A2 => n25903, ZN => n17682);
   U8219 : OAI21_X1 port map( A1 => n16279, A2 => n12507, B => n24875, ZN => 
                           n26574);
   U8221 : OR2_X1 port map( A1 => n22799, A2 => n14424, Z => n2133);
   U8229 : NOR2_X1 port map( A1 => n24977, A2 => n4925, ZN => n24877);
   U8232 : NAND2_X2 port map( A1 => n24880, A2 => n25549, ZN => n24225);
   U8248 : NAND2_X2 port map( A1 => n16046, A2 => n16047, ZN => n23107);
   U8266 : XOR2_X1 port map( A1 => n24886, A2 => n27423, Z => n26192);
   U8279 : NAND3_X2 port map( A1 => n13208, A2 => n23706, A3 => n11967, ZN => 
                           n14765);
   U8331 : NAND3_X1 port map( A1 => n16517, A2 => n27239, A3 => n24552, ZN => 
                           n16245);
   U8333 : NOR2_X2 port map( A1 => n11876, A2 => n11875, ZN => n12500);
   U8353 : XOR2_X1 port map( A1 => n19264, A2 => n6419, Z => n6416);
   U8375 : NAND2_X2 port map( A1 => n5941, A2 => n5943, ZN => n19264);
   U8404 : XOR2_X1 port map( A1 => n18239, A2 => n18013, Z => n25068);
   U8407 : NAND2_X2 port map( A1 => n17596, A2 => n17595, ZN => n18013);
   U8421 : AOI21_X2 port map( A1 => n24117, A2 => n6440, B => n6439, ZN => 
                           n12493);
   U8426 : OAI22_X2 port map( A1 => n14862, A2 => n14861, B1 => n17188, B2 => 
                           n2713, ZN => n10355);
   U8437 : AOI21_X2 port map( A1 => n8174, A2 => n8175, B => n17449, ZN => 
                           n2910);
   U8438 : XOR2_X1 port map( A1 => n18128, A2 => n3556, Z => n25416);
   U8441 : NAND3_X2 port map( A1 => n20734, A2 => n13506, A3 => n20733, ZN => 
                           n8311);
   U8444 : OR2_X1 port map( A1 => n19878, A2 => n15575, Z => n25638);
   U8451 : NOR2_X2 port map( A1 => n26228, A2 => n26051, ZN => n12419);
   U8467 : NOR2_X2 port map( A1 => n2632, A2 => n23968, ZN => n19627);
   U8473 : XOR2_X1 port map( A1 => n6540, A2 => n13382, Z => n25767);
   U8474 : NAND2_X2 port map( A1 => n6502, A2 => n24596, ZN => n6540);
   U8475 : XOR2_X1 port map( A1 => n5783, A2 => n5782, Z => n24199);
   U8503 : XOR2_X1 port map( A1 => n18282, A2 => n24894, Z => n11015);
   U8507 : XOR2_X1 port map( A1 => n18012, A2 => n14322, Z => n24894);
   U8508 : NAND3_X2 port map( A1 => n18696, A2 => n18613, A3 => n18697, ZN => 
                           n24895);
   U8530 : OAI21_X2 port map( A1 => n23093, A2 => n17432, B => n9434, ZN => 
                           n24897);
   U8542 : NAND2_X2 port map( A1 => n9366, A2 => n3198, ZN => n9365);
   U8544 : NAND3_X2 port map( A1 => n833, A2 => n10422, A3 => n16433, ZN => 
                           n24899);
   U8545 : NAND3_X1 port map( A1 => n12369, A2 => n12331, A3 => n12368, ZN => 
                           n24900);
   U8546 : NOR2_X1 port map( A1 => n1109, A2 => n12946, ZN => n9026);
   U8548 : NOR2_X2 port map( A1 => n20151, A2 => n7057, ZN => n11403);
   U8552 : XOR2_X1 port map( A1 => n24901, A2 => n26833, Z => n15546);
   U8554 : XOR2_X1 port map( A1 => n25006, A2 => n13382, Z => n24901);
   U8573 : XOR2_X1 port map( A1 => n18311, A2 => n2157, Z => n2156);
   U8576 : XOR2_X1 port map( A1 => n18137, A2 => n18125, Z => n18311);
   U8578 : AOI22_X1 port map( A1 => n20066, A2 => n25795, B1 => n19972, B2 => 
                           n4782, ZN => n19973);
   U8579 : NOR2_X2 port map( A1 => n4782, A2 => n4537, ZN => n20066);
   U8580 : NAND2_X2 port map( A1 => n20570, A2 => n734, ZN => n25527);
   U8589 : XOR2_X1 port map( A1 => n5624, A2 => n25647, Z => n24903);
   U8595 : INV_X2 port map( I => n16422, ZN => n11952);
   U8597 : OR2_X1 port map( A1 => n22763, A2 => n5578, Z => n6924);
   U8603 : XOR2_X1 port map( A1 => n28510, A2 => n16826, Z => n23940);
   U8606 : NOR2_X2 port map( A1 => n4493, A2 => n26307, ZN => n25439);
   U8608 : XOR2_X1 port map( A1 => n24906, A2 => n24905, Z => n22478);
   U8610 : XOR2_X1 port map( A1 => n24623, A2 => n20551, Z => n24905);
   U8622 : XOR2_X1 port map( A1 => n24910, A2 => n15201, Z => n1696);
   U8635 : NAND2_X2 port map( A1 => n3726, A2 => n3727, ZN => n19999);
   U8652 : NAND2_X2 port map( A1 => n6159, A2 => n25163, ZN => n5682);
   U8655 : AOI21_X2 port map( A1 => n24914, A2 => n26695, B => n111, ZN => 
                           n2247);
   U8659 : XOR2_X1 port map( A1 => n6416, A2 => n25767, Z => n25762);
   U8660 : XOR2_X1 port map( A1 => n8438, A2 => n21281, Z => n8396);
   U8661 : NAND2_X2 port map( A1 => n10240, A2 => n10238, ZN => n8438);
   U8671 : NAND2_X1 port map( A1 => n17288, A2 => n1030, ZN => n25694);
   U8682 : OAI22_X2 port map( A1 => n25420, A2 => n253, B1 => n8245, B2 => n956
                           , ZN => n24917);
   U8696 : BUF_X2 port map( I => n7971, Z => n24922);
   U8697 : OAI21_X2 port map( A1 => n24576, A2 => n27406, B => n4085, ZN => 
                           n8449);
   U8700 : NAND2_X2 port map( A1 => n24924, A2 => n11806, ZN => n7971);
   U8703 : XOR2_X1 port map( A1 => n24926, A2 => n24925, Z => n25536);
   U8707 : NOR2_X1 port map( A1 => n21658, A2 => n27411, ZN => n24927);
   U8711 : NOR2_X2 port map( A1 => n24541, A2 => n2403, ZN => n13051);
   U8714 : NAND2_X1 port map( A1 => n17574, A2 => n12999, ZN => n25123);
   U8719 : NAND2_X2 port map( A1 => n8393, A2 => n24932, ZN => n13793);
   U8724 : AOI21_X2 port map( A1 => n4653, A2 => n21944, B => n24934, ZN => 
                           n21148);
   U8735 : NAND2_X1 port map( A1 => n28507, A2 => n13028, ZN => n24935);
   U8737 : NAND2_X1 port map( A1 => n13371, A2 => n24937, ZN => n24936);
   U8739 : NOR2_X1 port map( A1 => n484, A2 => n808, ZN => n25575);
   U8757 : NAND2_X1 port map( A1 => n15468, A2 => n15474, ZN => n21601);
   U8771 : XOR2_X1 port map( A1 => n19552, A2 => n11918, Z => n25853);
   U8778 : OR2_X1 port map( A1 => n26633, A2 => n25614, Z => n19590);
   U8781 : OR2_X1 port map( A1 => n17637, A2 => n23110, Z => n10850);
   U8784 : NOR2_X2 port map( A1 => n18555, A2 => n18554, ZN => n25104);
   U8798 : AOI22_X1 port map( A1 => n21225, A2 => n26333, B1 => n26059, B2 => 
                           n21226, ZN => n26337);
   U8803 : NAND2_X2 port map( A1 => n24941, A2 => n8416, ZN => n5751);
   U8806 : NAND2_X2 port map( A1 => n25894, A2 => n994, ZN => n24941);
   U8818 : BUF_X4 port map( I => n15077, Z => n25786);
   U8820 : NAND2_X2 port map( A1 => n4191, A2 => n9525, ZN => n11789);
   U8829 : AND2_X1 port map( A1 => n6725, A2 => n19033, Z => n8828);
   U8833 : XOR2_X1 port map( A1 => n10921, A2 => n10966, Z => n13491);
   U8839 : XOR2_X1 port map( A1 => n25533, A2 => n8959, Z => n24944);
   U8845 : NOR2_X1 port map( A1 => n25575, A2 => n10932, ZN => n23617);
   U8852 : NOR2_X2 port map( A1 => n4774, A2 => n4775, ZN => n25874);
   U8853 : INV_X2 port map( I => n25795, ZN => n859);
   U8865 : AOI21_X2 port map( A1 => n17634, A2 => n14230, B => n17633, ZN => 
                           n18048);
   U8871 : NOR2_X2 port map( A1 => n15331, A2 => n14326, ZN => n16324);
   U8905 : AOI21_X2 port map( A1 => n15648, A2 => n9762, B => n24950, ZN => 
                           n7211);
   U8907 : INV_X2 port map( I => n21118, ZN => n23976);
   U8913 : NAND2_X2 port map( A1 => n25778, A2 => n11904, ZN => n21118);
   U8926 : NOR2_X2 port map( A1 => n12934, A2 => n12935, ZN => n18103);
   U8929 : INV_X2 port map( I => n16336, ZN => n24952);
   U8936 : OAI21_X1 port map( A1 => n21690, A2 => n27403, B => n21691, ZN => 
                           n21584);
   U8937 : NAND3_X2 port map( A1 => n24953, A2 => n22558, A3 => n17922, ZN => 
                           n15284);
   U8939 : NAND3_X1 port map( A1 => n10691, A2 => n22765, A3 => n15096, ZN => 
                           n24953);
   U8940 : XOR2_X1 port map( A1 => n23582, A2 => n24954, Z => n7940);
   U8942 : INV_X2 port map( I => n13253, ZN => n24955);
   U8946 : NAND2_X2 port map( A1 => n15879, A2 => n15880, ZN => n16823);
   U8947 : XOR2_X1 port map( A1 => n24957, A2 => n21649, Z => Ciphertext(167));
   U8949 : NAND3_X2 port map( A1 => n15427, A2 => n15428, A3 => n15426, ZN => 
                           n24957);
   U8950 : NAND2_X1 port map( A1 => n21007, A2 => n14583, ZN => n21002);
   U8952 : OR2_X1 port map( A1 => n17795, A2 => n25688, Z => n26609);
   U8956 : INV_X4 port map( I => n16712, ZN => n12039);
   U8958 : NOR2_X2 port map( A1 => n7720, A2 => n10305, ZN => n16712);
   U8971 : XOR2_X1 port map( A1 => n18119, A2 => n28541, Z => n7717);
   U8979 : NAND2_X1 port map( A1 => n4857, A2 => n25018, ZN => n24185);
   U8990 : NAND2_X2 port map( A1 => n763, A2 => n24564, ZN => n17739);
   U8997 : XOR2_X1 port map( A1 => n19340, A2 => n19339, Z => n6344);
   U9002 : NAND3_X2 port map( A1 => n2981, A2 => n658, A3 => n6242, ZN => n2465
                           );
   U9004 : AND2_X2 port map( A1 => n10548, A2 => n10542, Z => n18543);
   U9015 : INV_X4 port map( I => n10548, ZN => n5554);
   U9019 : AOI21_X2 port map( A1 => n1685, A2 => n1491, B => n724, ZN => n1683)
                           ;
   U9021 : NAND2_X2 port map( A1 => n25707, A2 => n4035, ZN => n4034);
   U9023 : XOR2_X1 port map( A1 => n24960, A2 => n553, Z => n10252);
   U9027 : XOR2_X1 port map( A1 => n9802, A2 => n25946, Z => n24960);
   U9028 : XOR2_X1 port map( A1 => n3614, A2 => n3616, Z => n4263);
   U9030 : XOR2_X1 port map( A1 => n25969, A2 => n24962, Z => n25970);
   U9031 : XOR2_X1 port map( A1 => n17140, A2 => n23659, Z => n24962);
   U9043 : XOR2_X1 port map( A1 => n13793, A2 => n1290, Z => n24963);
   U9053 : NAND2_X1 port map( A1 => n7919, A2 => n14502, ZN => n12096);
   U9058 : XOR2_X1 port map( A1 => n24111, A2 => n24964, Z => n19784);
   U9061 : XOR2_X1 port map( A1 => n19407, A2 => n21838, Z => n24964);
   U9075 : NAND2_X2 port map( A1 => n17549, A2 => n17550, ZN => n14269);
   U9080 : XOR2_X1 port map( A1 => n19325, A2 => n4697, Z => n4696);
   U9100 : NAND3_X2 port map( A1 => n22257, A2 => n6665, A3 => n6666, ZN => 
                           n12644);
   U9104 : NAND2_X2 port map( A1 => n17230, A2 => n17554, ZN => n24966);
   U9105 : XOR2_X1 port map( A1 => n24967, A2 => n3036, Z => n21877);
   U9107 : XOR2_X1 port map( A1 => n14294, A2 => n24968, Z => n24967);
   U9109 : OAI21_X2 port map( A1 => n14635, A2 => n21867, B => n838, ZN => 
                           n14068);
   U9111 : INV_X4 port map( I => n25161, ZN => n23161);
   U9115 : OAI21_X2 port map( A1 => n24970, A2 => n2533, B => n22386, ZN => 
                           n24114);
   U9124 : NOR2_X1 port map( A1 => n1848, A2 => n15187, ZN => n24971);
   U9128 : NAND2_X2 port map( A1 => n17243, A2 => n17242, ZN => n17924);
   U9129 : AND2_X1 port map( A1 => n814, A2 => n10601, Z => n10469);
   U9131 : NAND2_X2 port map( A1 => n24974, A2 => n10804, ZN => n4224);
   U9132 : OAI21_X2 port map( A1 => n15459, A2 => n15460, B => n23062, ZN => 
                           n24974);
   U9136 : XOR2_X1 port map( A1 => n4478, A2 => n20536, Z => n3970);
   U9139 : XOR2_X1 port map( A1 => n12382, A2 => n20450, Z => n20536);
   U9140 : AOI21_X1 port map( A1 => n14458, A2 => n21003, B => n25003, ZN => 
                           n25288);
   U9145 : NAND3_X2 port map( A1 => n24975, A2 => n10228, A3 => n11422, ZN => 
                           n10190);
   U9152 : OAI22_X1 port map( A1 => n2308, A2 => n15678, B1 => n2307, B2 => 
                           n13961, ZN => n23614);
   U9161 : NAND3_X2 port map( A1 => n692, A2 => n2095, A3 => n21004, ZN => 
                           n21006);
   U9168 : XOR2_X1 port map( A1 => n9985, A2 => n19300, Z => n3941);
   U9169 : XOR2_X1 port map( A1 => n22577, A2 => n3372, Z => n19300);
   U9197 : OAI22_X2 port map( A1 => n2469, A2 => n6372, B1 => n17662, B2 => 
                           n12599, ZN => n22207);
   U9205 : AOI22_X2 port map( A1 => n25786, A2 => n17488, B1 => n17561, B2 => 
                           n13997, ZN => n24986);
   U9216 : INV_X2 port map( I => n24990, ZN => n14914);
   U9219 : XNOR2_X1 port map( A1 => n7391, A2 => n11090, ZN => n24990);
   U9222 : XOR2_X1 port map( A1 => n18328, A2 => n24991, Z => n24116);
   U9223 : XOR2_X1 port map( A1 => n18221, A2 => n18290, Z => n24991);
   U9224 : NOR2_X2 port map( A1 => n19582, A2 => n23444, ZN => n22776);
   U9226 : NAND2_X2 port map( A1 => n25639, A2 => n25638, ZN => n19582);
   U9227 : XOR2_X1 port map( A1 => n10208, A2 => n24992, Z => n3586);
   U9230 : XOR2_X1 port map( A1 => n24275, A2 => n19478, Z => n24992);
   U9233 : INV_X1 port map( I => n22879, ZN => n12572);
   U9241 : NAND2_X1 port map( A1 => n6237, A2 => n14584, ZN => n527);
   U9242 : INV_X2 port map( I => n24995, ZN => n9464);
   U9244 : XNOR2_X1 port map( A1 => n26600, A2 => n3760, ZN => n24995);
   U9245 : BUF_X2 port map( I => n15490, Z => n24996);
   U9260 : XOR2_X1 port map( A1 => n9742, A2 => n9739, Z => n304);
   U9269 : INV_X2 port map( I => n14338, ZN => n14912);
   U9271 : NAND2_X2 port map( A1 => n10147, A2 => n12938, ZN => n14338);
   U9282 : AND2_X1 port map( A1 => n15104, A2 => n13417, Z => n14310);
   U9284 : XOR2_X1 port map( A1 => n19518, A2 => n14686, Z => n14151);
   U9287 : NAND2_X2 port map( A1 => n25004, A2 => n23443, ZN => n21237);
   U9288 : NAND2_X1 port map( A1 => n7931, A2 => n7930, ZN => n25004);
   U9289 : XOR2_X1 port map( A1 => n9585, A2 => n25005, Z => n26501);
   U9292 : NAND2_X1 port map( A1 => n9584, A2 => n7186, ZN => n11205);
   U9298 : XOR2_X1 port map( A1 => n25007, A2 => n14614, Z => Ciphertext(57));
   U9303 : NAND2_X1 port map( A1 => n4520, A2 => n4521, ZN => n4519);
   U9304 : OAI21_X2 port map( A1 => n969, A2 => n11936, B => n25635, ZN => 
                           n15250);
   U9309 : AOI21_X2 port map( A1 => n24187, A2 => n19748, B => n15667, ZN => 
                           n25008);
   U9311 : XOR2_X1 port map( A1 => n1876, A2 => n1875, Z => n26257);
   U9314 : OAI21_X2 port map( A1 => n10780, A2 => n25010, B => n16404, ZN => 
                           n22692);
   U9316 : NAND2_X2 port map( A1 => n8468, A2 => n20817, ZN => n9567);
   U9321 : NAND2_X1 port map( A1 => n20255, A2 => n26652, ZN => n25011);
   U9322 : NAND2_X1 port map( A1 => n20021, A2 => n9579, ZN => n25012);
   U9326 : OAI21_X2 port map( A1 => n12518, A2 => n7178, B => n17986, ZN => 
                           n15681);
   U9327 : XOR2_X1 port map( A1 => n3211, A2 => n27461, Z => n6640);
   U9328 : NAND3_X1 port map( A1 => n17401, A2 => n10209, A3 => n11113, ZN => 
                           n22415);
   U9332 : NAND2_X2 port map( A1 => n5081, A2 => n9773, ZN => n16732);
   U9343 : INV_X4 port map( I => n13205, ZN => n25724);
   U9345 : NAND2_X2 port map( A1 => n6007, A2 => n13637, ZN => n13205);
   U9346 : XOR2_X1 port map( A1 => n2352, A2 => n25328, Z => n21142);
   U9366 : NOR2_X2 port map( A1 => n16191, A2 => n14108, ZN => n12151);
   U9368 : NAND2_X2 port map( A1 => n25016, A2 => n25015, ZN => n16191);
   U9371 : INV_X1 port map( I => n15881, ZN => n25015);
   U9375 : INV_X2 port map( I => n15025, ZN => n25016);
   U9378 : BUF_X2 port map( I => n16167, Z => n25017);
   U9379 : OR2_X1 port map( A1 => n25045, A2 => n20165, Z => n25018);
   U9386 : XOR2_X1 port map( A1 => n19173, A2 => n19177, Z => n3845);
   U9408 : OR2_X1 port map( A1 => n21989, A2 => n20339, Z => n22409);
   U9410 : INV_X1 port map( I => n22813, ZN => n25934);
   U9433 : NOR2_X1 port map( A1 => n1431, A2 => n21005, ZN => n3739);
   U9434 : AND2_X1 port map( A1 => n3326, A2 => n23023, Z => n1342);
   U9437 : XOR2_X1 port map( A1 => n8112, A2 => n97, Z => n8109);
   U9441 : OAI21_X2 port map( A1 => n2154, A2 => n2155, B => n15568, ZN => 
                           n25024);
   U9447 : XOR2_X1 port map( A1 => n16859, A2 => n17014, Z => n10169);
   U9449 : OAI22_X2 port map( A1 => n13067, A2 => n9903, B1 => n9902, B2 => 
                           n16858, ZN => n17014);
   U9459 : XOR2_X1 port map( A1 => n2889, A2 => n2888, Z => n8890);
   U9464 : NOR2_X2 port map( A1 => n24440, A2 => n12453, ZN => n25798);
   U9466 : NOR2_X1 port map( A1 => n2857, A2 => n12039, ZN => n16714);
   U9481 : OAI22_X1 port map( A1 => n7054, A2 => n27367, B1 => n16578, B2 => 
                           n8223, ZN => n3564);
   U9491 : XOR2_X1 port map( A1 => n26962, A2 => n15126, Z => n19331);
   U9492 : NAND2_X2 port map( A1 => n9326, A2 => n9327, ZN => n15126);
   U9495 : XOR2_X1 port map( A1 => n16992, A2 => n25028, Z => n5522);
   U9502 : XOR2_X1 port map( A1 => n14294, A2 => n25029, Z => n25028);
   U9509 : OAI22_X2 port map( A1 => n25665, A2 => n1872, B1 => n8270, B2 => 
                           n8269, ZN => n11376);
   U9513 : NOR2_X1 port map( A1 => n3644, A2 => n14256, ZN => n4712);
   U9516 : NAND2_X2 port map( A1 => n4182, A2 => n4180, ZN => n14256);
   U9517 : OAI21_X2 port map( A1 => n5073, A2 => n5074, B => n838, ZN => n5072)
                           ;
   U9519 : INV_X4 port map( I => n6216, ZN => n13788);
   U9528 : OAI21_X2 port map( A1 => n25924, A2 => n4063, B => n25030, ZN => 
                           n18234);
   U9536 : OAI21_X2 port map( A1 => n15550, A2 => n28540, B => n4063, ZN => 
                           n25030);
   U9539 : XOR2_X1 port map( A1 => n16841, A2 => n16840, Z => n16842);
   U9553 : AOI22_X2 port map( A1 => n3040, A2 => n20110, B1 => n4136, B2 => 
                           n2891, ZN => n25687);
   U9555 : XOR2_X1 port map( A1 => n2508, A2 => n25372, Z => n19171);
   U9558 : AOI21_X2 port map( A1 => n3033, A2 => n9226, B => n3031, ZN => n2508
                           );
   U9573 : NAND2_X2 port map( A1 => n20193, A2 => n955, ZN => n14855);
   U9584 : NAND2_X2 port map( A1 => n25768, A2 => n12166, ZN => n12718);
   U9595 : INV_X2 port map( I => n25034, ZN => n8031);
   U9602 : XOR2_X1 port map( A1 => Plaintext(121), A2 => Key(121), Z => n25034)
                           ;
   U9606 : XOR2_X1 port map( A1 => n28370, A2 => n22135, Z => n15108);
   U9608 : XOR2_X1 port map( A1 => n16899, A2 => n25036, Z => n5610);
   U9616 : XOR2_X1 port map( A1 => n25037, A2 => n21227, Z => Ciphertext(112));
   U9617 : NAND2_X1 port map( A1 => n14755, A2 => n26337, ZN => n25037);
   U9620 : XOR2_X1 port map( A1 => n25038, A2 => n24662, Z => n25113);
   U9631 : AND2_X2 port map( A1 => n19189, A2 => n7030, Z => n21757);
   U9632 : BUF_X2 port map( I => n15917, Z => n14456);
   U9638 : XOR2_X1 port map( A1 => n4273, A2 => n4272, Z => n10246);
   U9639 : NAND2_X2 port map( A1 => n7182, A2 => n21788, ZN => n19839);
   U9640 : NAND2_X1 port map( A1 => n765, A2 => n24509, ZN => n4861);
   U9649 : XOR2_X1 port map( A1 => n4302, A2 => n4301, Z => n15632);
   U9650 : NAND2_X1 port map( A1 => n993, A2 => n2356, ZN => n7597);
   U9651 : NOR2_X2 port map( A1 => n2358, A2 => n2357, ZN => n14836);
   U9656 : XOR2_X1 port map( A1 => n7751, A2 => n7763, Z => n25039);
   U9660 : XOR2_X1 port map( A1 => n20008, A2 => n8138, Z => n14961);
   U9667 : NOR2_X1 port map( A1 => n12637, A2 => n16426, ZN => n11194);
   U9676 : NOR2_X1 port map( A1 => n5715, A2 => n21682, ZN => n25049);
   U9682 : AOI21_X2 port map( A1 => n26073, A2 => n27258, B => n26822, ZN => 
                           n25042);
   U9686 : NAND2_X2 port map( A1 => n25043, A2 => n11744, ZN => n11983);
   U9687 : NAND2_X2 port map( A1 => n9675, A2 => n10133, ZN => n26042);
   U9689 : XOR2_X1 port map( A1 => n2439, A2 => n18324, Z => n18313);
   U9690 : AOI22_X2 port map( A1 => n15664, A2 => n1217, B1 => n15663, B2 => 
                           n23927, ZN => n2439);
   U9691 : NAND2_X1 port map( A1 => n18875, A2 => n26395, ZN => n26335);
   U9692 : NAND2_X2 port map( A1 => n19803, A2 => n11936, ZN => n19629);
   U9709 : AOI21_X2 port map( A1 => n19785, A2 => n27443, B => n27730, ZN => 
                           n14522);
   U9720 : XOR2_X1 port map( A1 => n4987, A2 => n4986, Z => n4985);
   U9728 : NAND2_X2 port map( A1 => n19688, A2 => n3152, ZN => n20226);
   U9731 : NAND2_X2 port map( A1 => n5421, A2 => n14565, ZN => n19794);
   U9742 : NAND2_X2 port map( A1 => n10210, A2 => n27380, ZN => n6651);
   U9750 : NOR2_X2 port map( A1 => n17317, A2 => n12040, ZN => n17400);
   U9770 : NOR2_X2 port map( A1 => n26894, A2 => n7212, ZN => n18566);
   U9781 : NAND3_X2 port map( A1 => n21139, A2 => n15463, A3 => n21140, ZN => 
                           n25052);
   U9784 : INV_X1 port map( I => n25102, ZN => n3383);
   U9786 : NAND2_X1 port map( A1 => n25054, A2 => n12235, ZN => n20678);
   U9791 : AND2_X1 port map( A1 => n4705, A2 => n4702, Z => n8321);
   U9792 : NOR2_X1 port map( A1 => n815, A2 => n19836, ZN => n19840);
   U9797 : NOR2_X2 port map( A1 => n24323, A2 => n5353, ZN => n8770);
   U9810 : AND2_X1 port map( A1 => n25322, A2 => n2631, Z => n19626);
   U9834 : OAI22_X2 port map( A1 => n1685, A2 => n27204, B1 => n7794, B2 => 
                           n22174, ZN => n1684);
   U9840 : NAND3_X2 port map( A1 => n25979, A2 => n19834, A3 => n19892, ZN => 
                           n11033);
   U9845 : AND2_X1 port map( A1 => n8193, A2 => n25380, Z => n4885);
   U9871 : NAND2_X2 port map( A1 => n2339, A2 => n23955, ZN => n4559);
   U9878 : INV_X2 port map( I => n1970, ZN => n2604);
   U9880 : NAND2_X2 port map( A1 => n17609, A2 => n13618, ZN => n1970);
   U9886 : BUF_X4 port map( I => n10548, Z => n25935);
   U9889 : XOR2_X1 port map( A1 => n22169, A2 => n24312, Z => n9256);
   U9890 : XOR2_X1 port map( A1 => n9904, A2 => n9670, Z => n7644);
   U9894 : OAI22_X2 port map( A1 => n25069, A2 => n14672, B1 => n6682, B2 => 
                           n26522, ZN => n6215);
   U9896 : NOR2_X2 port map( A1 => n19753, A2 => n10690, ZN => n25069);
   U9900 : INV_X1 port map( I => n19160, ZN => n25070);
   U9901 : NAND2_X2 port map( A1 => n16122, A2 => n3651, ZN => n25071);
   U9917 : NAND2_X2 port map( A1 => n1455, A2 => n25074, ZN => n10268);
   U9930 : INV_X2 port map( I => n25547, ZN => n26627);
   U9948 : XOR2_X1 port map( A1 => n23047, A2 => n11322, Z => n13363);
   U9950 : NOR2_X1 port map( A1 => n7565, A2 => n22391, ZN => n6090);
   U9954 : INV_X2 port map( I => n22718, ZN => n24539);
   U9957 : OR2_X1 port map( A1 => n21220, A2 => n26059, Z => n13526);
   U9964 : XOR2_X1 port map( A1 => n12090, A2 => n25188, Z => n17555);
   U9974 : XOR2_X1 port map( A1 => n20359, A2 => n26453, Z => n23454);
   U9976 : NOR2_X2 port map( A1 => n25670, A2 => n729, ZN => n5709);
   U9979 : XOR2_X1 port map( A1 => n7861, A2 => n23636, Z => n26583);
   U9983 : OAI21_X1 port map( A1 => n18747, A2 => n18643, B => n25082, ZN => 
                           n17893);
   U9987 : NAND2_X2 port map( A1 => n20730, A2 => n8594, ZN => n6243);
   U9997 : AOI21_X2 port map( A1 => n2603, A2 => n10655, B => n2602, ZN => 
                           n25099);
   U10006 : XOR2_X1 port map( A1 => n19311, A2 => n4026, Z => n1712);
   U10012 : OAI21_X2 port map( A1 => n6880, A2 => n6683, B => n25086, ZN => 
                           n6878);
   U10018 : NAND2_X2 port map( A1 => n1893, A2 => n10779, ZN => n12494);
   U10033 : NAND2_X2 port map( A1 => n5708, A2 => n5710, ZN => n5718);
   U10039 : XOR2_X1 port map( A1 => n4811, A2 => n13524, Z => n17037);
   U10043 : NOR2_X2 port map( A1 => n16727, A2 => n3159, ZN => n4811);
   U10062 : XOR2_X1 port map( A1 => n25946, A2 => n10056, Z => n4723);
   U10073 : NAND2_X2 port map( A1 => n25090, A2 => n11118, ZN => n19334);
   U10074 : NAND2_X1 port map( A1 => n25237, A2 => n3645, ZN => n2062);
   U10090 : XOR2_X1 port map( A1 => n17718, A2 => n25093, Z => n25092);
   U10097 : XOR2_X1 port map( A1 => n26066, A2 => n14642, Z => n15228);
   U10099 : XOR2_X1 port map( A1 => n21142, A2 => n19701, Z => n12081);
   U10102 : NAND2_X2 port map( A1 => n11018, A2 => n25094, ZN => n6473);
   U10104 : NAND2_X1 port map( A1 => n14508, A2 => n11017, ZN => n25094);
   U10111 : NAND2_X2 port map( A1 => n6729, A2 => n6730, ZN => n25095);
   U10119 : INV_X2 port map( I => n18120, ZN => n18263);
   U10126 : XOR2_X1 port map( A1 => n13510, A2 => n13511, Z => n24223);
   U10130 : AOI22_X2 port map( A1 => n16387, A2 => n7180, B1 => n15120, B2 => 
                           n5558, ZN => n25097);
   U10132 : NOR2_X1 port map( A1 => n28468, A2 => n2023, ZN => n14090);
   U10138 : XOR2_X1 port map( A1 => n633, A2 => n7723, Z => n1389);
   U10139 : XOR2_X1 port map( A1 => n2467, A2 => n14187, Z => n12909);
   U10140 : NOR2_X2 port map( A1 => n4543, A2 => n4546, ZN => n14187);
   U10141 : OR2_X1 port map( A1 => n25173, A2 => n25547, Z => n3974);
   U10142 : XOR2_X1 port map( A1 => n2611, A2 => n26409, Z => n19932);
   U10143 : XOR2_X1 port map( A1 => n2378, A2 => n26037, Z => n23415);
   U10145 : AOI21_X2 port map( A1 => n17328, A2 => n17269, B => n17507, ZN => 
                           n1485);
   U10149 : OAI21_X2 port map( A1 => n13567, A2 => n13566, B => n14552, ZN => 
                           n13565);
   U10153 : BUF_X2 port map( I => n6419, Z => n25098);
   U10169 : AOI21_X2 port map( A1 => n3710, A2 => n22785, B => n22555, ZN => 
                           n13395);
   U10172 : XOR2_X1 port map( A1 => n16817, A2 => n16883, Z => n16992);
   U10176 : NOR2_X2 port map( A1 => n1760, A2 => n1759, ZN => n16817);
   U10187 : NOR2_X2 port map( A1 => n15979, A2 => n16136, ZN => n14150);
   U10192 : NAND2_X1 port map( A1 => n23674, A2 => n20316, ZN => n19969);
   U10195 : XOR2_X1 port map( A1 => n25488, A2 => n17037, Z => n23528);
   U10202 : NAND2_X2 port map( A1 => n23951, A2 => n3783, ZN => n23391);
   U10212 : OR2_X1 port map( A1 => n25106, A2 => n23391, Z => n5892);
   U10222 : BUF_X4 port map( I => n18646, Z => n11299);
   U10235 : AOI22_X2 port map( A1 => n17902, A2 => n23115, B1 => n17900, B2 => 
                           n28247, ZN => n18171);
   U10256 : NAND2_X2 port map( A1 => n28444, A2 => n27432, ZN => n25109);
   U10257 : NAND2_X2 port map( A1 => n6874, A2 => n25110, ZN => n13248);
   U10260 : INV_X2 port map( I => n25111, ZN => n14815);
   U10261 : XOR2_X1 port map( A1 => Plaintext(119), A2 => Key(119), Z => n25111
                           );
   U10262 : OAI22_X2 port map( A1 => n6197, A2 => n6198, B1 => n6195, B2 => 
                           n6196, ZN => n14397);
   U10283 : OAI21_X2 port map( A1 => n12375, A2 => n14648, B => n5801, ZN => 
                           n23332);
   U10284 : BUF_X4 port map( I => n19861, Z => n4810);
   U10285 : NAND2_X2 port map( A1 => n23669, A2 => n1929, ZN => n5874);
   U10290 : INV_X2 port map( I => n25113, ZN => n18527);
   U10294 : NAND2_X2 port map( A1 => n2591, A2 => n2590, ZN => n24236);
   U10299 : NAND2_X2 port map( A1 => n24114, A2 => n2530, ZN => n10494);
   U10300 : NAND3_X2 port map( A1 => n9689, A2 => n9687, A3 => n25114, ZN => 
                           n25421);
   U10306 : OAI21_X1 port map( A1 => n26206, A2 => n4021, B => n25115, ZN => 
                           n4108);
   U10312 : OAI22_X1 port map( A1 => n17962, A2 => n13981, B1 => n23023, B2 => 
                           n13235, ZN => n13428);
   U10329 : NAND2_X1 port map( A1 => n22378, A2 => n22453, ZN => n22280);
   U10346 : OR2_X1 port map( A1 => n28088, A2 => n6315, Z => n6840);
   U10349 : XOR2_X1 port map( A1 => n1833, A2 => n1831, Z => n8598);
   U10354 : NAND2_X1 port map( A1 => n21352, A2 => n21353, ZN => n21354);
   U10367 : NOR2_X1 port map( A1 => n25316, A2 => n21160, ZN => n13525);
   U10376 : NAND2_X2 port map( A1 => n8864, A2 => n12314, ZN => n13099);
   U10384 : NAND2_X2 port map( A1 => n28378, A2 => n19683, ZN => n23424);
   U10397 : XOR2_X1 port map( A1 => n25120, A2 => n8238, Z => n6853);
   U10413 : OAI22_X2 port map( A1 => n14648, A2 => n27887, B1 => n28542, B2 => 
                           n9464, ZN => n9323);
   U10450 : NAND2_X2 port map( A1 => n25123, A2 => n2740, ZN => n18003);
   U10465 : NOR2_X1 port map( A1 => n27456, A2 => n840, ZN => n15952);
   U10466 : INV_X2 port map( I => n2404, ZN => n238);
   U10473 : XOR2_X1 port map( A1 => n25125, A2 => n21262, Z => Ciphertext(16));
   U10484 : AOI22_X2 port map( A1 => n11468, A2 => n22747, B1 => n1765, B2 => 
                           n9737, ZN => n21641);
   U10494 : NAND2_X2 port map( A1 => n23313, A2 => n1764, ZN => n11468);
   U10525 : INV_X2 port map( I => n25128, ZN => n19759);
   U10527 : XNOR2_X1 port map( A1 => n7471, A2 => n672, ZN => n25128);
   U10533 : XOR2_X1 port map( A1 => n8710, A2 => n25129, Z => n26620);
   U10542 : XOR2_X1 port map( A1 => n13157, A2 => n9197, Z => n25129);
   U10556 : XOR2_X1 port map( A1 => n7598, A2 => n8608, Z => n18300);
   U10563 : INV_X2 port map( I => n9773, ZN => n25130);
   U10589 : INV_X2 port map( I => n20153, ZN => n20151);
   U10605 : XOR2_X1 port map( A1 => n7976, A2 => n5359, Z => n8545);
   U10618 : XOR2_X1 port map( A1 => n20376, A2 => n21085, Z => n517);
   U10620 : INV_X2 port map( I => n25133, ZN => n18646);
   U10667 : NAND2_X2 port map( A1 => n25136, A2 => n8635, ZN => n11319);
   U10717 : XOR2_X1 port map( A1 => n8776, A2 => n1709, Z => n7727);
   U10719 : NAND2_X2 port map( A1 => n25137, A2 => n17181, ZN => n26308);
   U10720 : OAI21_X2 port map( A1 => n17565, A2 => n13358, B => n7361, ZN => 
                           n25137);
   U10721 : OR2_X1 port map( A1 => n11089, A2 => n9131, Z => n12254);
   U10727 : NAND2_X2 port map( A1 => n6491, A2 => n6494, ZN => n6490);
   U10729 : NAND2_X1 port map( A1 => n1886, A2 => n665, ZN => n15575);
   U10730 : XOR2_X1 port map( A1 => n25531, A2 => n12031, Z => n1886);
   U10743 : XOR2_X1 port map( A1 => n18194, A2 => n18193, Z => n25138);
   U10753 : INV_X2 port map( I => n22598, ZN => n25141);
   U10769 : XOR2_X1 port map( A1 => n1680, A2 => n25143, Z => n10313);
   U10783 : OAI21_X1 port map( A1 => n8576, A2 => n7791, B => n5098, ZN => 
                           n4035);
   U10789 : OR2_X1 port map( A1 => n1045, A2 => n6373, Z => n5603);
   U10792 : NAND2_X2 port map( A1 => n25144, A2 => n4110, ZN => n6628);
   U10794 : BUF_X2 port map( I => n20730, Z => n25145);
   U10798 : INV_X2 port map( I => n23546, ZN => n7568);
   U10811 : NOR2_X2 port map( A1 => n23488, A2 => n998, ZN => n2894);
   U10812 : NAND3_X2 port map( A1 => n873, A2 => n26570, A3 => n8554, ZN => 
                           n1813);
   U10814 : AND2_X1 port map( A1 => n9446, A2 => n23642, Z => n21808);
   U10817 : XNOR2_X1 port map( A1 => n9035, A2 => n9037, ZN => n19792);
   U10818 : OR2_X1 port map( A1 => n14815, A2 => n14814, Z => n16050);
   U10830 : INV_X2 port map( I => n14033, ZN => n23542);
   U10831 : INV_X4 port map( I => n6006, ZN => n9450);
   U10851 : NAND2_X2 port map( A1 => n1977, A2 => n1980, ZN => n17053);
   U10859 : NOR2_X2 port map( A1 => n13573, A2 => n12111, ZN => n18970);
   U10862 : XOR2_X1 port map( A1 => n27661, A2 => n16883, Z => n1725);
   U10867 : NAND3_X2 port map( A1 => n8148, A2 => n2249, A3 => n11633, ZN => 
                           n12674);
   U10871 : NAND2_X2 port map( A1 => n21775, A2 => n13432, ZN => n25150);
   U10873 : NAND2_X2 port map( A1 => n25151, A2 => n23401, ZN => n4491);
   U10877 : XOR2_X1 port map( A1 => n25152, A2 => n5792, Z => n24344);
   U10878 : XOR2_X1 port map( A1 => n5772, A2 => n28550, Z => n25152);
   U10888 : XOR2_X1 port map( A1 => n20411, A2 => n25156, Z => n4064);
   U10890 : XOR2_X1 port map( A1 => n11021, A2 => n21868, Z => n25156);
   U10910 : NAND3_X2 port map( A1 => n22238, A2 => n26284, A3 => n18425, ZN => 
                           n25162);
   U10916 : XOR2_X1 port map( A1 => n3665, A2 => n25165, Z => n6291);
   U10917 : XOR2_X1 port map( A1 => n3419, A2 => n20344, Z => n3665);
   U10921 : NAND2_X1 port map( A1 => n6162, A2 => n11629, ZN => n25163);
   U10931 : INV_X1 port map( I => n25166, ZN => n2459);
   U10933 : XOR2_X1 port map( A1 => n27360, A2 => n20872, Z => n25165);
   U10937 : NAND2_X2 port map( A1 => n15725, A2 => n18382, ZN => n4212);
   U10955 : NAND2_X1 port map( A1 => n25168, A2 => n20658, ZN => n20659);
   U10956 : INV_X1 port map( I => n3824, ZN => n25168);
   U10957 : NAND2_X2 port map( A1 => n3828, A2 => n25243, ZN => n3824);
   U10958 : XOR2_X1 port map( A1 => n16862, A2 => n16937, Z => n10705);
   U10959 : NAND2_X2 port map( A1 => n15336, A2 => n15337, ZN => n16862);
   U10968 : XOR2_X1 port map( A1 => n20449, A2 => n9055, Z => n9982);
   U10980 : XOR2_X1 port map( A1 => n4707, A2 => n14733, Z => n4159);
   U10981 : XOR2_X1 port map( A1 => n172, A2 => n25439, Z => n14733);
   U10996 : XOR2_X1 port map( A1 => n25174, A2 => n21917, Z => n3236);
   U11000 : NAND2_X1 port map( A1 => n21124, A2 => n21118, ZN => n21122);
   U11002 : NAND2_X2 port map( A1 => n17436, A2 => n17508, ZN => n17328);
   U11010 : NAND2_X1 port map( A1 => n21166, A2 => n11107, ZN => n2228);
   U11012 : OAI21_X2 port map( A1 => n15606, A2 => n849, B => n24422, ZN => 
                           n21166);
   U11022 : XOR2_X1 port map( A1 => n18189, A2 => n25178, Z => n23116);
   U11023 : XOR2_X1 port map( A1 => n3834, A2 => n25651, Z => n25178);
   U11039 : XOR2_X1 port map( A1 => n1098, A2 => n25362, Z => n2193);
   U11041 : NAND3_X2 port map( A1 => n25180, A2 => n10165, A3 => n25179, ZN => 
                           n9734);
   U11043 : NOR2_X1 port map( A1 => n25359, A2 => n16676, ZN => n16049);
   U11055 : NAND3_X2 port map( A1 => n5225, A2 => n7253, A3 => n7254, ZN => 
                           n13794);
   U11056 : XOR2_X1 port map( A1 => n25181, A2 => n17122, Z => n7242);
   U11063 : XOR2_X1 port map( A1 => n22597, A2 => n16991, Z => n25183);
   U11064 : NAND2_X2 port map( A1 => n20261, A2 => n19956, ZN => n19957);
   U11066 : XOR2_X1 port map( A1 => n18084, A2 => n2796, Z => n23319);
   U11070 : INV_X2 port map( I => n25184, ZN => n7824);
   U11086 : XOR2_X1 port map( A1 => n16839, A2 => n25185, Z => n1473);
   U11088 : XOR2_X1 port map( A1 => n16838, A2 => n24651, Z => n25185);
   U11094 : NAND2_X2 port map( A1 => n21397, A2 => n23802, ZN => n24422);
   U11107 : OAI21_X2 port map( A1 => n11123, A2 => n20253, B => n25186, ZN => 
                           n14876);
   U11112 : XOR2_X1 port map( A1 => n4095, A2 => n23829, Z => n23269);
   U11117 : NAND2_X2 port map( A1 => n1813, A2 => n22075, ZN => n1811);
   U11118 : NAND3_X1 port map( A1 => n24563, A2 => n4898, A3 => n17580, ZN => 
                           n25720);
   U11122 : XOR2_X1 port map( A1 => n11678, A2 => n24625, Z => n25507);
   U11123 : XOR2_X1 port map( A1 => n16989, A2 => n11679, Z => n11678);
   U11132 : XOR2_X1 port map( A1 => n19313, A2 => n14600, Z => n6135);
   U11134 : NOR2_X2 port map( A1 => n24339, A2 => n1624, ZN => n19313);
   U11145 : NAND2_X2 port map( A1 => n8290, A2 => n22727, ZN => n23422);
   U11146 : XOR2_X1 port map( A1 => n12089, A2 => n17103, Z => n25188);
   U11148 : XOR2_X1 port map( A1 => n17153, A2 => n17152, Z => n17156);
   U11151 : XOR2_X1 port map( A1 => n21237, A2 => n12995, Z => n20577);
   U11158 : OAI21_X2 port map( A1 => n4449, A2 => n4002, B => n25191, ZN => 
                           n24343);
   U11166 : NAND2_X2 port map( A1 => n10345, A2 => n2730, ZN => n2832);
   U11169 : OR2_X1 port map( A1 => n15003, A2 => n20852, Z => n7955);
   U11170 : XOR2_X1 port map( A1 => n25372, A2 => n2508, Z => n2504);
   U11171 : OAI22_X2 port map( A1 => n8054, A2 => n24332, B1 => n8052, B2 => 
                           n8645, ZN => n25372);
   U11182 : NOR2_X1 port map( A1 => n21872, A2 => n480, ZN => n26568);
   U11184 : OAI21_X2 port map( A1 => n26585, A2 => n26586, B => n21576, ZN => 
                           n21608);
   U11189 : INV_X2 port map( I => n2434, ZN => n9854);
   U11201 : NOR2_X2 port map( A1 => n15187, A2 => n9538, ZN => n2394);
   U11205 : INV_X4 port map( I => n4224, ZN => n15187);
   U11208 : NAND2_X2 port map( A1 => n6476, A2 => n25196, ZN => n5442);
   U11210 : NAND3_X2 port map( A1 => n6479, A2 => n16300, A3 => n14732, ZN => 
                           n25196);
   U11211 : INV_X2 port map( I => n25197, ZN => n16544);
   U11218 : OAI21_X2 port map( A1 => n24050, A2 => n24049, B => n18702, ZN => 
                           n25198);
   U11224 : XOR2_X1 port map( A1 => n3603, A2 => n3602, Z => n3601);
   U11225 : XOR2_X1 port map( A1 => n19465, A2 => n19463, Z => n3086);
   U11226 : XOR2_X1 port map( A1 => n2462, A2 => n868, Z => n19463);
   U11230 : NAND2_X1 port map( A1 => n21349, A2 => n11156, ZN => n25203);
   U11232 : BUF_X2 port map( I => n21970, Z => n25199);
   U11237 : NOR2_X2 port map( A1 => n10629, A2 => n14385, ZN => n15104);
   U11248 : XOR2_X1 port map( A1 => n24343, A2 => n23352, Z => n1526);
   U11250 : OAI22_X2 port map( A1 => n1504, A2 => n14254, B1 => n1503, B2 => 
                           n13964, ZN => n23352);
   U11258 : OR2_X1 port map( A1 => n19661, A2 => n598, Z => n24474);
   U11261 : XOR2_X1 port map( A1 => n19356, A2 => n25208, Z => n13425);
   U11265 : XOR2_X1 port map( A1 => n299, A2 => n19355, Z => n25208);
   U11271 : INV_X4 port map( I => n12521, ZN => n14791);
   U11282 : AOI22_X1 port map( A1 => n21226, A2 => n7039, B1 => n10217, B2 => 
                           n14901, ZN => n12394);
   U11288 : OAI21_X2 port map( A1 => n8025, A2 => n14332, B => n18726, ZN => 
                           n15379);
   U11293 : NOR3_X1 port map( A1 => n25755, A2 => n734, A3 => n25756, ZN => 
                           n22071);
   U11305 : OR2_X1 port map( A1 => n19011, A2 => n22626, Z => n4734);
   U11314 : NAND2_X1 port map( A1 => n25216, A2 => n3389, ZN => n1470);
   U11316 : NOR2_X2 port map( A1 => n17802, A2 => n17588, ZN => n25789);
   U11328 : NAND3_X1 port map( A1 => n14409, A2 => n21064, A3 => n9377, ZN => 
                           n6851);
   U11329 : NOR2_X2 port map( A1 => n13819, A2 => n17976, ZN => n26264);
   U11330 : NAND2_X2 port map( A1 => n25684, A2 => n4463, ZN => n13819);
   U11333 : NAND2_X1 port map( A1 => n25218, A2 => n25217, ZN => n17579);
   U11335 : NAND2_X1 port map( A1 => n2895, A2 => n17578, ZN => n25217);
   U11337 : NAND2_X1 port map( A1 => n17787, A2 => n6076, ZN => n25218);
   U11340 : NAND2_X2 port map( A1 => n14320, A2 => n13415, ZN => n8999);
   U11347 : XOR2_X1 port map( A1 => n11328, A2 => n19220, Z => n9339);
   U11348 : NAND2_X2 port map( A1 => n18855, A2 => n18854, ZN => n19220);
   U11349 : XOR2_X1 port map( A1 => n9832, A2 => n9357, Z => n8244);
   U11356 : XOR2_X1 port map( A1 => n18077, A2 => n18029, Z => n9357);
   U11357 : NAND2_X1 port map( A1 => n25949, A2 => n21087, ZN => n10622);
   U11360 : BUF_X2 port map( I => n16288, Z => n6427);
   U11362 : NAND2_X2 port map( A1 => n17355, A2 => n26614, ZN => n17480);
   U11387 : NAND2_X2 port map( A1 => n17253, A2 => n17252, ZN => n17927);
   U11388 : NOR2_X2 port map( A1 => n20430, A2 => n14611, ZN => n20287);
   U11399 : AOI22_X2 port map( A1 => n25907, A2 => n27713, B1 => n2418, B2 => 
                           n3937, ZN => n9117);
   U11401 : BUF_X2 port map( I => n15964, Z => n25225);
   U11410 : OAI21_X2 port map( A1 => n19185, A2 => n24674, B => n19799, ZN => 
                           n26445);
   U11412 : AOI22_X2 port map( A1 => n8192, A2 => n19796, B1 => n23968, B2 => 
                           n19633, ZN => n19799);
   U11422 : NAND2_X2 port map( A1 => n23187, A2 => n8013, ZN => n25445);
   U11443 : XOR2_X1 port map( A1 => n20534, A2 => n20485, Z => n8808);
   U11444 : AOI21_X1 port map( A1 => n12434, A2 => n26578, B => n2391, ZN => 
                           n16512);
   U11451 : NAND2_X2 port map( A1 => n10989, A2 => n10990, ZN => n13443);
   U11460 : NOR2_X2 port map( A1 => n17220, A2 => n21824, ZN => n11217);
   U11461 : XOR2_X1 port map( A1 => Plaintext(190), A2 => Key(190), Z => n15964
                           );
   U11471 : NAND2_X2 port map( A1 => n16673, A2 => n5973, ZN => n25671);
   U11473 : AOI21_X2 port map( A1 => n7840, A2 => n15429, B => n987, ZN => 
                           n10348);
   U11476 : NOR2_X1 port map( A1 => n16220, A2 => n6063, ZN => n25235);
   U11480 : XOR2_X1 port map( A1 => n24582, A2 => n5474, Z => n25648);
   U11481 : XOR2_X1 port map( A1 => n26962, A2 => n7659, Z => n7204);
   U11482 : NAND2_X2 port map( A1 => n7657, A2 => n6601, ZN => n7659);
   U11490 : NOR2_X2 port map( A1 => n25236, A2 => n12863, ZN => n2653);
   U11497 : INV_X2 port map( I => n20856, ZN => n25628);
   U11500 : NAND2_X2 port map( A1 => n25629, A2 => n25630, ZN => n20856);
   U11505 : XOR2_X1 port map( A1 => n19533, A2 => n592, Z => n2673);
   U11513 : XOR2_X1 port map( A1 => Plaintext(12), A2 => Key(12), Z => n22623);
   U11517 : XOR2_X1 port map( A1 => n21260, A2 => n6616, Z => n11026);
   U11531 : NAND2_X2 port map( A1 => n15078, A2 => n25242, ZN => n14920);
   U11532 : NAND2_X1 port map( A1 => n7452, A2 => n7453, ZN => n13034);
   U11536 : XOR2_X1 port map( A1 => n27466, A2 => n13077, Z => n2071);
   U11537 : NOR2_X2 port map( A1 => n21843, A2 => n22388, ZN => n25243);
   U11552 : AND2_X1 port map( A1 => n18863, A2 => n25339, Z => n10720);
   U11558 : NAND2_X1 port map( A1 => n19605, A2 => n19785, ZN => n5606);
   U11560 : NOR2_X2 port map( A1 => n12617, A2 => n1711, ZN => n19605);
   U11564 : OAI21_X2 port map( A1 => n8473, A2 => n8435, B => n17291, ZN => 
                           n25246);
   U11569 : XOR2_X1 port map( A1 => n17121, A2 => n25247, Z => n10524);
   U11570 : XOR2_X1 port map( A1 => n25744, A2 => n16875, Z => n25247);
   U11579 : XOR2_X1 port map( A1 => n3368, A2 => n24711, Z => n18790);
   U11580 : AOI21_X2 port map( A1 => n3906, A2 => n3905, B => n18789, ZN => 
                           n3368);
   U11581 : AOI21_X2 port map( A1 => n1049, A2 => n13758, B => n4162, ZN => 
                           n25249);
   U11584 : XOR2_X1 port map( A1 => n16774, A2 => n16751, Z => n5435);
   U11585 : NAND2_X1 port map( A1 => n2749, A2 => n10992, ZN => n21710);
   U11588 : NAND2_X2 port map( A1 => n22924, A2 => n2160, ZN => n2749);
   U11596 : XOR2_X1 port map( A1 => n18136, A2 => n10754, Z => n12855);
   U11603 : OAI21_X1 port map( A1 => n23399, A2 => n27867, B => n8357, ZN => 
                           n25252);
   U11612 : XNOR2_X1 port map( A1 => Key(164), A2 => Plaintext(164), ZN => 
                           n25253);
   U11620 : BUF_X2 port map( I => n25693, Z => n25255);
   U11623 : XOR2_X1 port map( A1 => n25257, A2 => n13859, Z => Ciphertext(121))
                           ;
   U11631 : AOI22_X1 port map( A1 => n21339, A2 => n21338, B1 => n21356, B2 => 
                           n21343, ZN => n25257);
   U11645 : XOR2_X1 port map( A1 => n16951, A2 => n14145, Z => n17074);
   U11661 : NAND2_X2 port map( A1 => n9912, A2 => n13357, ZN => n3398);
   U11668 : NOR2_X2 port map( A1 => n17442, A2 => n24509, ZN => n6425);
   U11673 : OR2_X1 port map( A1 => n26461, A2 => n11947, Z => n11792);
   U11678 : INV_X2 port map( I => n4832, ZN => n7275);
   U11684 : AOI22_X1 port map( A1 => n13602, A2 => n12918, B1 => n15104, B2 => 
                           n16332, ZN => n13601);
   U11694 : INV_X2 port map( I => n19975, ZN => n961);
   U11695 : NAND2_X2 port map( A1 => n13002, A2 => n7236, ZN => n19975);
   U11697 : NOR2_X1 port map( A1 => n16360, A2 => n25693, ZN => n11547);
   U11698 : NOR2_X2 port map( A1 => n14657, A2 => n16075, ZN => n25693);
   U11701 : XOR2_X1 port map( A1 => n24004, A2 => n14715, Z => n14712);
   U11718 : NAND2_X2 port map( A1 => n13434, A2 => n22875, ZN => n11947);
   U11722 : NAND2_X1 port map( A1 => n16403, A2 => n4556, ZN => n25550);
   U11729 : NAND3_X2 port map( A1 => n24391, A2 => n24330, A3 => n6642, ZN => 
                           n17716);
   U11730 : AOI21_X1 port map( A1 => n17386, A2 => n17385, B => n10183, ZN => 
                           n4805);
   U11731 : INV_X2 port map( I => n24234, ZN => n10183);
   U11736 : XOR2_X1 port map( A1 => n8016, A2 => n8017, Z => n24234);
   U11744 : NAND2_X2 port map( A1 => n11870, A2 => n22835, ZN => n20260);
   U11763 : OAI21_X1 port map( A1 => n20950, A2 => n23662, B => n477, ZN => 
                           n14466);
   U11764 : NOR2_X2 port map( A1 => n12235, A2 => n10534, ZN => n20670);
   U11769 : NOR2_X2 port map( A1 => n25263, A2 => n24142, ZN => n627);
   U11780 : XOR2_X1 port map( A1 => n11672, A2 => n20549, Z => n25541);
   U11794 : INV_X1 port map( I => n16784, ZN => n147);
   U11797 : XNOR2_X1 port map( A1 => n26823, A2 => n4811, ZN => n17149);
   U11801 : XOR2_X1 port map( A1 => n2439, A2 => n1777, Z => n18189);
   U11808 : NAND2_X2 port map( A1 => n14446, A2 => n17927, ZN => n17773);
   U11810 : NOR2_X2 port map( A1 => n6426, A2 => n878, ZN => n1500);
   U11811 : NAND2_X2 port map( A1 => n11185, A2 => n11184, ZN => n15725);
   U11812 : BUF_X2 port map( I => n15872, Z => n25266);
   U11823 : NAND2_X2 port map( A1 => n16462, A2 => n25267, ZN => n94);
   U11833 : OAI22_X2 port map( A1 => n12383, A2 => n13758, B1 => n3981, B2 => 
                           n12384, ZN => n25267);
   U11847 : AND2_X1 port map( A1 => n26292, A2 => n18427, Z => n3886);
   U11855 : NOR2_X2 port map( A1 => n23018, A2 => n21761, ZN => n8726);
   U11860 : XOR2_X1 port map( A1 => n19411, A2 => n24669, Z => n25271);
   U11861 : XOR2_X1 port map( A1 => n3538, A2 => n3540, Z => n8012);
   U11862 : INV_X2 port map( I => n2231, ZN => n3060);
   U11867 : NAND2_X1 port map( A1 => n21123, A2 => n21122, ZN => n21127);
   U11879 : OR2_X1 port map( A1 => n16651, A2 => n9116, Z => n10891);
   U11880 : NAND2_X2 port map( A1 => n24151, A2 => n22672, ZN => n24481);
   U11897 : NAND2_X1 port map( A1 => n13518, A2 => n6193, ZN => n26481);
   U11899 : XOR2_X1 port map( A1 => n16958, A2 => n16897, Z => n16537);
   U11901 : NAND3_X2 port map( A1 => n7241, A2 => n15370, A3 => n16056, ZN => 
                           n16958);
   U11905 : XNOR2_X1 port map( A1 => n26216, A2 => n15609, ZN => n16940);
   U11906 : NAND2_X2 port map( A1 => n25619, A2 => n1596, ZN => n15609);
   U11919 : NAND2_X2 port map( A1 => n10820, A2 => n10819, ZN => n3729);
   U11925 : NOR2_X2 port map( A1 => n25484, A2 => n3467, ZN => n10820);
   U11928 : OAI22_X2 port map( A1 => n17994, A2 => n24391, B1 => n14342, B2 => 
                           n17845, ZN => n6430);
   U11931 : XOR2_X1 port map( A1 => n19331, A2 => n10671, Z => n13156);
   U11940 : NAND2_X2 port map( A1 => n8411, A2 => n20139, ZN => n20249);
   U11944 : NAND2_X2 port map( A1 => n696, A2 => n21641, ZN => n13908);
   U11960 : XOR2_X1 port map( A1 => n5858, A2 => n18916, Z => n2609);
   U11964 : INV_X2 port map( I => n19411, ZN => n5858);
   U11970 : OAI21_X2 port map( A1 => n26349, A2 => n25280, B => n15737, ZN => 
                           n5298);
   U11976 : NAND2_X2 port map( A1 => n20110, A2 => n978, ZN => n19726);
   U11982 : NOR2_X2 port map( A1 => n18749, A2 => n14376, ZN => n18497);
   U11994 : XOR2_X1 port map( A1 => n19276, A2 => n24035, Z => n24034);
   U12011 : XOR2_X1 port map( A1 => n18016, A2 => n18351, Z => n14979);
   U12015 : NAND2_X2 port map( A1 => n6518, A2 => n25282, ZN => n10359);
   U12023 : XOR2_X1 port map( A1 => n13514, A2 => n14000, Z => n1710);
   U12024 : XOR2_X1 port map( A1 => n28517, A2 => n11124, Z => n13514);
   U12027 : XOR2_X1 port map( A1 => n25284, A2 => n21010, Z => Ciphertext(76));
   U12028 : AND2_X1 port map( A1 => n18581, A2 => n22547, Z => n15459);
   U12029 : NOR2_X2 port map( A1 => n28378, A2 => n3317, ZN => n13911);
   U12031 : NAND2_X2 port map( A1 => n15903, A2 => n22984, ZN => n5861);
   U12038 : OR2_X1 port map( A1 => n11992, A2 => n17003, Z => n16969);
   U12043 : NOR2_X2 port map( A1 => n7096, A2 => n13062, ZN => n5938);
   U12046 : INV_X1 port map( I => n26104, ZN => n21866);
   U12058 : XOR2_X1 port map( A1 => n24079, A2 => n13464, Z => n9559);
   U12059 : OAI21_X2 port map( A1 => n10728, A2 => n14252, B => n1267, ZN => 
                           n6846);
   U12062 : XOR2_X1 port map( A1 => n25288, A2 => n1299, Z => Ciphertext(72));
   U12065 : XOR2_X1 port map( A1 => n23329, A2 => n4286, Z => n12315);
   U12067 : AND2_X2 port map( A1 => n18370, A2 => n2989, Z => n18381);
   U12076 : NAND2_X2 port map( A1 => n17200, A2 => n25290, ZN => n26076);
   U12077 : NOR2_X2 port map( A1 => n254, A2 => n12607, ZN => n26576);
   U12080 : XOR2_X1 port map( A1 => n25292, A2 => n18186, Z => n15177);
   U12084 : XOR2_X1 port map( A1 => n18360, A2 => n9076, Z => n18186);
   U12086 : XOR2_X1 port map( A1 => n1192, A2 => n27459, Z => n25292);
   U12089 : INV_X2 port map( I => n25293, ZN => n21890);
   U12099 : NOR2_X2 port map( A1 => n17463, A2 => n9459, ZN => n17458);
   U12105 : NAND2_X2 port map( A1 => n7964, A2 => n8512, ZN => n16391);
   U12106 : NAND2_X1 port map( A1 => n14858, A2 => n14174, ZN => n5464);
   U12129 : OAI21_X2 port map( A1 => n3088, A2 => n16346, B => n3089, ZN => 
                           n3297);
   U12134 : XOR2_X1 port map( A1 => n19533, A2 => n27388, Z => n1540);
   U12137 : AND2_X1 port map( A1 => n13009, A2 => n7454, Z => n13013);
   U12139 : INV_X1 port map( I => n8642, ZN => n20256);
   U12143 : NAND2_X1 port map( A1 => n22830, A2 => n20155, ZN => n8642);
   U12153 : INV_X2 port map( I => n18575, ZN => n11262);
   U12168 : AOI22_X2 port map( A1 => n24639, A2 => n815, B1 => n11130, B2 => 
                           n19836, ZN => n5249);
   U12186 : NOR2_X2 port map( A1 => n18101, A2 => n22396, ZN => n4014);
   U12189 : NOR2_X2 port map( A1 => n25477, A2 => n16030, ZN => n16640);
   U12192 : NAND3_X1 port map( A1 => n18446, A2 => n18534, A3 => n18533, ZN => 
                           n25662);
   U12193 : NAND2_X2 port map( A1 => n1180, A2 => n5407, ZN => n18446);
   U12194 : AOI21_X2 port map( A1 => n16169, A2 => n15787, B => n25303, ZN => 
                           n16483);
   U12200 : NAND2_X2 port map( A1 => n25426, A2 => n14328, ZN => n25303);
   U12201 : INV_X4 port map( I => n23437, ZN => n3347);
   U12204 : XOR2_X1 port map( A1 => n9455, A2 => n17077, Z => n11041);
   U12212 : INV_X2 port map( I => n18793, ZN => n18873);
   U12222 : NAND2_X2 port map( A1 => n6999, A2 => n9050, ZN => n18944);
   U12232 : AND2_X1 port map( A1 => n25318, A2 => n4822, Z => n4820);
   U12242 : NOR2_X1 port map( A1 => n22767, A2 => n20894, ZN => n12129);
   U12261 : BUF_X2 port map( I => n24344, Z => n25304);
   U12271 : INV_X1 port map( I => n24344, ZN => n690);
   U12273 : NAND2_X1 port map( A1 => n13398, A2 => n22925, ZN => n22924);
   U12284 : AOI21_X1 port map( A1 => n24316, A2 => n11937, B => n22734, ZN => 
                           n24461);
   U12285 : NAND2_X1 port map( A1 => n20171, A2 => n859, ZN => n6160);
   U12297 : NAND3_X1 port map( A1 => n132, A2 => n2131, A3 => n703, ZN => 
                           n16056);
   U12301 : INV_X1 port map( I => n16284, ZN => n14452);
   U12318 : NAND2_X1 port map( A1 => n7908, A2 => n14663, ZN => n7925);
   U12344 : INV_X2 port map( I => n6589, ZN => n11820);
   U12347 : INV_X1 port map( I => n12195, ZN => n11558);
   U12350 : CLKBUF_X4 port map( I => n5118, Z => n26169);
   U12356 : NOR2_X1 port map( A1 => n9446, A2 => n23642, ZN => n20126);
   U12376 : AND2_X2 port map( A1 => n5367, A2 => n14666, Z => n14665);
   U12377 : NOR2_X1 port map( A1 => n5367, A2 => n20868, ZN => n13037);
   U12380 : CLKBUF_X4 port map( I => n19584, Z => n978);
   U12389 : NAND2_X1 port map( A1 => n10133, A2 => n237, ZN => n17710);
   U12392 : NAND2_X1 port map( A1 => n10133, A2 => n10136, ZN => n10132);
   U12414 : XOR2_X1 port map( A1 => n8652, A2 => n25991, Z => n25308);
   U12425 : OR2_X1 port map( A1 => n13490, A2 => n27432, Z => n21845);
   U12434 : NAND2_X1 port map( A1 => n25692, A2 => n7354, ZN => n20779);
   U12456 : NAND2_X1 port map( A1 => n10194, A2 => n17032, ZN => n5076);
   U12457 : OAI22_X1 port map( A1 => n2537, A2 => n17501, B1 => n17345, B2 => 
                           n1233, ZN => n26166);
   U12471 : NOR2_X1 port map( A1 => n13799, A2 => n23578, ZN => n13950);
   U12473 : NAND2_X1 port map( A1 => n13979, A2 => n21616, ZN => n13992);
   U12481 : XOR2_X1 port map( A1 => n20538, A2 => n11885, Z => n25310);
   U12488 : INV_X1 port map( I => n20917, ZN => n22728);
   U12489 : OAI21_X1 port map( A1 => n1071, A2 => n20917, B => n26006, ZN => 
                           n7906);
   U12495 : NAND4_X1 port map( A1 => n17552, A2 => n17551, A3 => n17549, A4 => 
                           n17550, ZN => n17542);
   U12505 : NAND2_X1 port map( A1 => n19961, A2 => n7364, ZN => n5031);
   U12511 : AND2_X1 port map( A1 => n22385, A2 => n26764, Z => n8130);
   U12523 : OR2_X2 port map( A1 => n9083, A2 => n10026, Z => n25313);
   U12527 : NAND2_X1 port map( A1 => n25750, A2 => n20781, ZN => n22040);
   U12536 : INV_X2 port map( I => n6543, ZN => n14750);
   U12537 : NOR2_X1 port map( A1 => n28295, A2 => n25679, ZN => n2955);
   U12539 : OR2_X1 port map( A1 => n10593, A2 => n27409, Z => n9135);
   U12543 : NOR2_X1 port map( A1 => n14584, A2 => n5095, ZN => n15868);
   U12552 : AND2_X1 port map( A1 => n26317, A2 => n13372, Z => n2155);
   U12565 : INV_X2 port map( I => n20030, ZN => n1105);
   U12567 : INV_X1 port map( I => n20030, ZN => n25999);
   U12573 : NAND2_X1 port map( A1 => n19064, A2 => n4669, ZN => n4668);
   U12574 : XNOR2_X1 port map( A1 => n17754, A2 => n13122, ZN => n2621);
   U12592 : NAND2_X1 port map( A1 => n7525, A2 => n796, ZN => n16142);
   U12596 : OAI21_X1 port map( A1 => n19869, A2 => n11474, B => n19650, ZN => 
                           n11473);
   U12599 : NOR3_X1 port map( A1 => n20915, A2 => n846, A3 => n20911, ZN => 
                           n7440);
   U12600 : AOI22_X1 port map( A1 => n20152, A2 => n7618, B1 => n20338, B2 => 
                           n7057, ZN => n7634);
   U12613 : AND2_X1 port map( A1 => n10810, A2 => n20277, Z => n4649);
   U12616 : NAND3_X1 port map( A1 => n27924, A2 => n1081, A3 => n13505, ZN => 
                           n13506);
   U12630 : NAND2_X1 port map( A1 => n17458, A2 => n28035, ZN => n17466);
   U12637 : AOI21_X1 port map( A1 => n26435, A2 => n13291, B => n21620, ZN => 
                           n13993);
   U12645 : CLKBUF_X4 port map( I => n8246, Z => n7807);
   U12649 : AND2_X1 port map( A1 => n23753, A2 => n20803, Z => n8990);
   U12657 : AOI22_X1 port map( A1 => n26574, A2 => n13533, B1 => n16282, B2 => 
                           n14346, ZN => n14728);
   U12658 : NOR2_X1 port map( A1 => n15897, A2 => n8191, ZN => n25659);
   U12685 : INV_X1 port map( I => n20588, ZN => n15316);
   U12693 : INV_X1 port map( I => n13131, ZN => n25488);
   U12700 : INV_X1 port map( I => n852, ZN => n25509);
   U12701 : NAND2_X1 port map( A1 => n2215, A2 => n11856, ZN => n25321);
   U12709 : NAND2_X2 port map( A1 => n5196, A2 => n21028, ZN => n9653);
   U12717 : BUF_X2 port map( I => n20436, Z => n7130);
   U12718 : OAI21_X1 port map( A1 => n6865, A2 => n7682, B => n19893, ZN => 
                           n12425);
   U12719 : CLKBUF_X12 port map( I => n19891, Z => n26158);
   U12720 : XOR2_X1 port map( A1 => n13561, A2 => n13560, Z => n25322);
   U12737 : NAND2_X1 port map( A1 => n26306, A2 => n14954, ZN => n26286);
   U12742 : NOR2_X1 port map( A1 => n20868, A2 => n10578, ZN => n12887);
   U12747 : INV_X1 port map( I => n10588, ZN => n10512);
   U12752 : AOI21_X1 port map( A1 => n4440, A2 => n15375, B => n6055, ZN => 
                           n3491);
   U12754 : NAND2_X1 port map( A1 => n21274, A2 => n3530, ZN => n21133);
   U12755 : OAI21_X2 port map( A1 => n20033, A2 => n13091, B => n806, ZN => 
                           n13090);
   U12756 : INV_X1 port map( I => n7319, ZN => n927);
   U12767 : NAND2_X1 port map( A1 => n21584, A2 => n27379, ZN => n15270);
   U12768 : OAI21_X1 port map( A1 => n800, A2 => n20803, B => n20801, ZN => 
                           n20800);
   U12773 : NAND2_X2 port map( A1 => n9074, A2 => n15713, ZN => n25324);
   U12784 : INV_X1 port map( I => n19045, ZN => n18930);
   U12785 : NAND2_X1 port map( A1 => n13788, A2 => n19045, ZN => n11494);
   U12788 : AOI21_X1 port map( A1 => n25809, A2 => n13234, B => n20685, ZN => 
                           n20668);
   U12800 : INV_X2 port map( I => n20938, ZN => n25326);
   U12812 : NAND3_X1 port map( A1 => n6498, A2 => n4537, A3 => n15412, ZN => 
                           n12897);
   U12816 : NOR2_X1 port map( A1 => n20732, A2 => n20730, ZN => n26146);
   U12823 : NOR2_X2 port map( A1 => n24443, A2 => n27411, ZN => n10124);
   U12842 : NOR2_X1 port map( A1 => n5415, A2 => n20316, ZN => n13835);
   U12845 : NOR2_X1 port map( A1 => n24209, A2 => n722, ZN => n5994);
   U12854 : INV_X1 port map( I => n16521, ZN => n2585);
   U12856 : INV_X1 port map( I => n23973, ZN => n19303);
   U12861 : INV_X1 port map( I => n26264, ZN => n5117);
   U12876 : NAND2_X1 port map( A1 => n20647, A2 => n4121, ZN => n7671);
   U12878 : NAND2_X1 port map( A1 => n20647, A2 => n8449, ZN => n4084);
   U12879 : NOR2_X1 port map( A1 => n20647, A2 => n20591, ZN => n5461);
   U12883 : AOI21_X1 port map( A1 => n18933, A2 => n19019, B => n24170, ZN => 
                           n18767);
   U12887 : XOR2_X1 port map( A1 => n3419, A2 => n20344, Z => n25330);
   U12894 : CLKBUF_X12 port map( I => n11809, Z => n25331);
   U12901 : NAND2_X1 port map( A1 => n6838, A2 => n10393, ZN => n24119);
   U12907 : INV_X2 port map( I => n25841, ZN => n731);
   U12913 : INV_X2 port map( I => n18661, ZN => n15423);
   U12918 : NAND3_X2 port map( A1 => n25637, A2 => n9495, A3 => n10300, ZN => 
                           n25333);
   U12921 : NAND3_X1 port map( A1 => n13187, A2 => n22812, A3 => n28234, ZN => 
                           n11633);
   U12927 : NOR2_X1 port map( A1 => n19833, A2 => n26447, ZN => n1598);
   U12928 : NOR2_X1 port map( A1 => n3559, A2 => n3593, ZN => n26290);
   U12947 : OAI22_X1 port map( A1 => n21416, A2 => n21415, B1 => n21414, B2 => 
                           n13741, ZN => n22607);
   U12949 : INV_X1 port map( I => n11820, ZN => n25334);
   U12950 : NAND2_X1 port map( A1 => n15724, A2 => n20852, ZN => n20853);
   U12955 : NOR2_X1 port map( A1 => n13050, A2 => n21160, ZN => n11134);
   U12973 : INV_X2 port map( I => n25305, ZN => n866);
   U12974 : OAI21_X2 port map( A1 => n24215, A2 => n2038, B => n5685, ZN => 
                           n5684);
   U12975 : NAND2_X1 port map( A1 => n3165, A2 => n25367, ZN => n3164);
   U12976 : NOR2_X1 port map( A1 => n826, A2 => n2403, ZN => n22285);
   U12985 : AND2_X2 port map( A1 => n13964, A2 => n14228, Z => n22418);
   U13000 : INV_X1 port map( I => n21290, ZN => n26010);
   U13005 : NAND2_X1 port map( A1 => n4110, A2 => n25854, ZN => n17968);
   U13018 : NAND2_X1 port map( A1 => n9722, A2 => n6718, ZN => n7873);
   U13031 : INV_X2 port map( I => n5317, ZN => n17664);
   U13032 : NOR2_X1 port map( A1 => n20598, A2 => n10666, ZN => n9977);
   U13036 : AOI21_X1 port map( A1 => n9376, A2 => n25914, B => n18914, ZN => 
                           n9409);
   U13046 : OAI21_X2 port map( A1 => n12419, A2 => n10789, B => n22054, ZN => 
                           n25339);
   U13050 : CLKBUF_X8 port map( I => n11553, Z => n25592);
   U13054 : NAND2_X1 port map( A1 => n6323, A2 => n13095, ZN => n20798);
   U13065 : OAI22_X2 port map( A1 => n11013, A2 => n216, B1 => n22209, B2 => 
                           n22208, ZN => n25342);
   U13069 : OAI22_X1 port map( A1 => n10263, A2 => n4131, B1 => n18580, B2 => 
                           n18581, ZN => n25907);
   U13070 : AOI22_X1 port map( A1 => n10263, A2 => n4131, B1 => n18580, B2 => 
                           n18581, ZN => n6074);
   U13076 : INV_X2 port map( I => n2689, ZN => n19623);
   U13079 : INV_X1 port map( I => n24312, ZN => n9709);
   U13084 : XOR2_X1 port map( A1 => n7079, A2 => n10033, Z => n25346);
   U13089 : AND2_X1 port map( A1 => n11619, A2 => n25346, Z => n10428);
   U13092 : XOR2_X1 port map( A1 => n15637, A2 => n1237, Z => n25347);
   U13095 : INV_X2 port map( I => n12610, ZN => n17986);
   U13110 : XOR2_X1 port map( A1 => n5142, A2 => n5144, Z => n25348);
   U13111 : XOR2_X1 port map( A1 => n10379, A2 => n22330, Z => n25349);
   U13115 : INV_X1 port map( I => n26646, ZN => n2703);
   U13135 : OAI22_X1 port map( A1 => n2469, A2 => n6372, B1 => n17662, B2 => 
                           n12599, ZN => n25351);
   U13143 : INV_X1 port map( I => n18048, ZN => n5602);
   U13147 : XOR2_X1 port map( A1 => n2507, A2 => n2389, Z => n25353);
   U13151 : OAI21_X1 port map( A1 => n17349, A2 => n7961, B => n7110, ZN => 
                           n11782);
   U13152 : AND2_X1 port map( A1 => n21228, A2 => n10268, Z => n7038);
   U13158 : NAND3_X1 port map( A1 => n10924, A2 => n6725, A3 => n874, ZN => 
                           n18339);
   U13163 : AOI21_X1 port map( A1 => n6725, A2 => n8290, B => n3960, ZN => 
                           n18340);
   U13164 : INV_X1 port map( I => n6725, ZN => n18942);
   U13172 : OAI21_X1 port map( A1 => n23823, A2 => n23824, B => n10268, ZN => 
                           n14755);
   U13179 : XOR2_X1 port map( A1 => n24176, A2 => n9034, Z => n25357);
   U13184 : INV_X1 port map( I => n20482, ZN => n26550);
   U13185 : NOR2_X1 port map( A1 => n4934, A2 => n20654, ZN => n20656);
   U13190 : INV_X2 port map( I => n15010, ZN => n18454);
   U13193 : AOI21_X1 port map( A1 => n14291, A2 => n820, B => n18546, ZN => 
                           n25665);
   U13194 : NAND2_X1 port map( A1 => n235, A2 => n18628, ZN => n7581);
   U13195 : NOR2_X2 port map( A1 => n12942, A2 => n12537, ZN => n25358);
   U13208 : NAND2_X1 port map( A1 => n7185, A2 => n10652, ZN => n25359);
   U13219 : NAND2_X2 port map( A1 => n23872, A2 => n11307, ZN => n25360);
   U13227 : NAND2_X1 port map( A1 => n5974, A2 => n6779, ZN => n12078);
   U13233 : INV_X2 port map( I => n25412, ZN => n18971);
   U13238 : OAI21_X1 port map( A1 => n12117, A2 => n9759, B => n16731, ZN => 
                           n9758);
   U13240 : INV_X1 port map( I => n26084, ZN => n8178);
   U13266 : OAI21_X1 port map( A1 => n1460, A2 => n14302, B => n1458, ZN => 
                           n23477);
   U13271 : XOR2_X1 port map( A1 => n9745, A2 => n9746, Z => n25363);
   U13276 : NAND2_X1 port map( A1 => n9051, A2 => n17855, ZN => n17856);
   U13286 : NAND2_X1 port map( A1 => n6056, A2 => n11891, ZN => n4440);
   U13288 : XNOR2_X1 port map( A1 => n15182, A2 => n5921, ZN => n12681);
   U13291 : INV_X1 port map( I => n15182, ZN => n1194);
   U13297 : NAND2_X1 port map( A1 => n17912, A2 => n17783, ZN => n13805);
   U13298 : XOR2_X1 port map( A1 => Plaintext(87), A2 => Key(87), Z => n25365);
   U13304 : NAND2_X1 port map( A1 => n14975, A2 => n23817, ZN => n4520);
   U13307 : NAND2_X1 port map( A1 => n7018, A2 => n19101, ZN => n13270);
   U13318 : NAND2_X1 port map( A1 => n7018, A2 => n18799, ZN => n5667);
   U13322 : NAND2_X1 port map( A1 => n7018, A2 => n27704, ZN => n18802);
   U13323 : NOR2_X1 port map( A1 => n12542, A2 => n7018, ZN => n14288);
   U13326 : INV_X1 port map( I => n19405, ZN => n4530);
   U13328 : OR2_X2 port map( A1 => n20078, A2 => n9365, Z => n20054);
   U13334 : INV_X1 port map( I => n12528, ZN => n15913);
   U13338 : AOI21_X1 port map( A1 => n799, A2 => n7460, B => n12528, ZN => 
                           n23367);
   U13342 : NOR3_X1 port map( A1 => n799, A2 => n7460, A3 => n12528, ZN => 
                           n3467);
   U13345 : XOR2_X1 port map( A1 => n4823, A2 => n4825, Z => n25366);
   U13356 : NOR2_X1 port map( A1 => n19106, A2 => n6778, ZN => n19108);
   U13357 : NAND2_X1 port map( A1 => n7319, A2 => n6543, ZN => n9166);
   U13366 : INV_X1 port map( I => n18168, ZN => n18307);
   U13368 : NOR2_X1 port map( A1 => n2869, A2 => n18879, ZN => n18417);
   U13370 : OAI22_X1 port map( A1 => n17770, A2 => n28322, B1 => n14284, B2 => 
                           n22307, ZN => n17238);
   U13371 : NOR2_X1 port map( A1 => n16597, A2 => n16639, ZN => n22703);
   U13375 : OAI21_X1 port map( A1 => n15180, A2 => n6321, B => n6318, ZN => 
                           n25369);
   U13404 : AOI21_X1 port map( A1 => n20915, A2 => n12486, B => n26006, ZN => 
                           n20916);
   U13407 : INV_X2 port map( I => n19110, ZN => n19117);
   U13408 : AOI22_X2 port map( A1 => n15664, A2 => n1217, B1 => n23927, B2 => 
                           n15663, ZN => n25371);
   U13417 : NAND2_X1 port map( A1 => n3178, A2 => n28019, ZN => n23264);
   U13438 : AND2_X1 port map( A1 => n24190, A2 => n25368, Z => n15622);
   U13441 : AOI21_X1 port map( A1 => n21608, A2 => n9611, B => n21609, ZN => 
                           n13829);
   U13445 : XOR2_X1 port map( A1 => Plaintext(130), A2 => Key(130), Z => n25373
                           );
   U13447 : XOR2_X1 port map( A1 => n22855, A2 => n11336, Z => n25374);
   U13451 : INV_X1 port map( I => n18748, ZN => n25375);
   U13453 : AOI21_X2 port map( A1 => n22155, A2 => n22154, B => n18962, ZN => 
                           n25376);
   U13464 : INV_X4 port map( I => n20263, ZN => n946);
   U13466 : INV_X2 port map( I => n3707, ZN => n12344);
   U13475 : NAND2_X1 port map( A1 => n26814, A2 => n16429, ZN => n10777);
   U13476 : AND3_X1 port map( A1 => n13768, A2 => n15524, A3 => n13052, Z => 
                           n25377);
   U13486 : AOI21_X2 port map( A1 => n7881, A2 => n20757, B => n7880, ZN => 
                           n6728);
   U13489 : INV_X2 port map( I => n28353, ZN => n11581);
   U13493 : NAND2_X1 port map( A1 => n25378, A2 => n11319, ZN => n20833);
   U13497 : INV_X2 port map( I => n15502, ZN => n18927);
   U13501 : AND2_X2 port map( A1 => n9779, A2 => n26323, Z => n25899);
   U13505 : CLKBUF_X12 port map( I => n21406, Z => n7199);
   U13511 : OAI22_X1 port map( A1 => n21416, A2 => n21407, B1 => n21403, B2 => 
                           n21402, ZN => n21404);
   U13513 : INV_X1 port map( I => n16526, ZN => n26518);
   U13515 : AOI21_X1 port map( A1 => n4479, A2 => n8250, B => n3171, ZN => 
                           n25386);
   U13517 : AOI21_X1 port map( A1 => n4479, A2 => n8250, B => n3171, ZN => 
                           n23344);
   U13534 : NAND2_X1 port map( A1 => n21000, A2 => n12186, ZN => n26492);
   U13535 : NAND2_X1 port map( A1 => n13467, A2 => n18686, ZN => n652);
   U13548 : XOR2_X1 port map( A1 => Plaintext(129), A2 => Key(129), Z => n25384
                           );
   U13555 : XOR2_X1 port map( A1 => n6706, A2 => n626, Z => n25385);
   U13562 : AOI21_X2 port map( A1 => n4479, A2 => n8250, B => n3171, ZN => 
                           n25387);
   U13568 : AND2_X2 port map( A1 => n5264, A2 => n6185, Z => n17232);
   U13573 : INV_X2 port map( I => n26465, ZN => n18924);
   U13576 : NOR2_X1 port map( A1 => n25390, A2 => n11854, ZN => n26421);
   U13577 : OAI21_X1 port map( A1 => n6145, A2 => n5877, B => n3014, ZN => 
                           n3013);
   U13578 : XOR2_X1 port map( A1 => n14248, A2 => n13359, Z => n25388);
   U13584 : NOR2_X1 port map( A1 => n18891, A2 => n26764, ZN => n5053);
   U13585 : NAND2_X1 port map( A1 => n7382, A2 => n15881, ZN => n11940);
   U13598 : INV_X1 port map( I => n24236, ZN => n14165);
   U13600 : OAI21_X2 port map( A1 => n9452, A2 => n24026, B => n9453, ZN => 
                           n25389);
   U13606 : INV_X2 port map( I => n7612, ZN => n19903);
   U13612 : NAND2_X1 port map( A1 => n11837, A2 => n21120, ZN => n21123);
   U13615 : XOR2_X1 port map( A1 => n4618, A2 => n3701, Z => n25391);
   U13618 : NOR2_X1 port map( A1 => n17522, A2 => n25385, ZN => n4887);
   U13624 : NAND4_X2 port map( A1 => n7510, A2 => n1883, A3 => n24273, A4 => 
                           n25392, ZN => n2460);
   U13638 : NAND2_X2 port map( A1 => n7897, A2 => n7898, ZN => n2179);
   U13639 : XOR2_X1 port map( A1 => n25396, A2 => n14589, Z => Ciphertext(105))
                           ;
   U13641 : NAND2_X1 port map( A1 => n25800, A2 => n7059, ZN => n25396);
   U13646 : NAND2_X2 port map( A1 => n22692, A2 => n4215, ZN => n22926);
   U13652 : XOR2_X1 port map( A1 => n25399, A2 => n6452, Z => n7004);
   U13653 : XOR2_X1 port map( A1 => n7309, A2 => n2528, Z => n25399);
   U13658 : AND2_X1 port map( A1 => n6522, A2 => n21545, Z => n25538);
   U13662 : NAND2_X2 port map( A1 => n6019, A2 => n327, ZN => n6018);
   U13666 : AOI21_X2 port map( A1 => n1771, A2 => n1023, B => n25930, ZN => 
                           n25400);
   U13675 : NAND2_X2 port map( A1 => n1475, A2 => n1914, ZN => n21314);
   U13676 : XOR2_X1 port map( A1 => n9102, A2 => n4525, Z => n4524);
   U13679 : XOR2_X1 port map( A1 => n5129, A2 => n5127, Z => n11719);
   U13685 : NAND2_X2 port map( A1 => n26158, A2 => n21769, ZN => n19835);
   U13686 : XOR2_X1 port map( A1 => n13661, A2 => n25401, Z => n1548);
   U13687 : XOR2_X1 port map( A1 => n17028, A2 => n12523, Z => n25401);
   U13693 : NAND2_X1 port map( A1 => n25403, A2 => n9867, ZN => n6883);
   U13700 : NAND2_X1 port map( A1 => n21084, A2 => n25952, ZN => n25403);
   U13714 : OAI21_X2 port map( A1 => n25405, A2 => n1938, B => n10742, ZN => 
                           n5047);
   U13719 : XOR2_X1 port map( A1 => n25407, A2 => n8440, Z => n8439);
   U13722 : XOR2_X1 port map( A1 => n3437, A2 => n3368, Z => n25520);
   U13723 : XOR2_X1 port map( A1 => n19501, A2 => n587, Z => n25408);
   U13724 : XOR2_X1 port map( A1 => n19231, A2 => n19382, Z => n19509);
   U13727 : NAND2_X2 port map( A1 => n25940, A2 => n16380, ZN => n16422);
   U13728 : INV_X4 port map( I => n15159, ZN => n15186);
   U13737 : NAND2_X2 port map( A1 => n25658, A2 => n15898, ZN => n15159);
   U13740 : NAND2_X2 port map( A1 => n9713, A2 => n9712, ZN => n25586);
   U13743 : XOR2_X1 port map( A1 => n18306, A2 => n25409, Z => n3501);
   U13748 : XOR2_X1 port map( A1 => n28292, A2 => n7256, Z => n25409);
   U13756 : XOR2_X1 port map( A1 => n17149, A2 => n25410, Z => n22877);
   U13763 : XOR2_X1 port map( A1 => n17039, A2 => n16924, Z => n16785);
   U13775 : XOR2_X1 port map( A1 => n2964, A2 => n2965, Z => n14426);
   U13783 : XOR2_X1 port map( A1 => n25414, A2 => n24885, Z => n538);
   U13786 : XOR2_X1 port map( A1 => n27430, A2 => n9876, Z => n4358);
   U13791 : NAND2_X2 port map( A1 => n4353, A2 => n4354, ZN => n9876);
   U13800 : AOI21_X1 port map( A1 => n8593, A2 => n13230, B => n25928, ZN => 
                           n22998);
   U13801 : NAND3_X2 port map( A1 => n6846, A2 => n6845, A3 => n6844, ZN => 
                           n6843);
   U13802 : XOR2_X1 port map( A1 => n25416, A2 => n3558, Z => n15010);
   U13805 : NAND2_X1 port map( A1 => n25500, A2 => n18454, ZN => n8527);
   U13807 : NAND2_X1 port map( A1 => n25366, A2 => n25357, ZN => n8464);
   U13827 : INV_X4 port map( I => n12117, ZN => n15701);
   U13828 : NAND2_X2 port map( A1 => n8286, A2 => n25451, ZN => n12117);
   U13829 : INV_X2 port map( I => n17139, ZN => n26449);
   U13832 : NAND2_X2 port map( A1 => n16252, A2 => n8796, ZN => n17139);
   U13842 : INV_X2 port map( I => n25419, ZN => n10730);
   U13848 : XOR2_X1 port map( A1 => n14972, A2 => n15318, Z => n25419);
   U13849 : AOI22_X2 port map( A1 => n15415, A2 => n26700, B1 => n10043, B2 => 
                           n7799, ZN => n18879);
   U13851 : XOR2_X1 port map( A1 => n13855, A2 => n6764, Z => n20420);
   U13859 : NAND2_X1 port map( A1 => n12586, A2 => n21542, ZN => n25422);
   U13862 : XOR2_X1 port map( A1 => n14796, A2 => n25423, Z => n11966);
   U13864 : XOR2_X1 port map( A1 => n16545, A2 => n11312, Z => n25423);
   U13873 : NOR2_X1 port map( A1 => n875, A2 => n18879, ZN => n26013);
   U13876 : XOR2_X1 port map( A1 => n11097, A2 => n25427, Z => n23973);
   U13877 : NAND2_X2 port map( A1 => n25332, A2 => n1137, ZN => n12433);
   U13881 : XOR2_X1 port map( A1 => n25428, A2 => n16852, Z => n24012);
   U13887 : NOR2_X1 port map( A1 => n7395, A2 => n16524, ZN => n25429);
   U13890 : INV_X1 port map( I => n7416, ZN => n25430);
   U13894 : AOI22_X2 port map( A1 => n18872, A2 => n15187, B1 => n19141, B2 => 
                           n10323, ZN => n25432);
   U13896 : XOR2_X1 port map( A1 => n6024, A2 => n823, Z => n18309);
   U13900 : OAI21_X2 port map( A1 => n11939, A2 => n11938, B => n1437, ZN => 
                           n6024);
   U13902 : NAND2_X2 port map( A1 => n2995, A2 => n17480, ZN => n5176);
   U13914 : XOR2_X1 port map( A1 => n985, A2 => n19405, Z => n12910);
   U13916 : NAND2_X2 port map( A1 => n25436, A2 => n25464, ZN => n15949);
   U13917 : NAND2_X2 port map( A1 => n25462, A2 => n27162, ZN => n25436);
   U13921 : INV_X2 port map( I => n7181, ZN => n10593);
   U13924 : INV_X4 port map( I => n19115, ZN => n997);
   U13926 : AOI22_X2 port map( A1 => n22430, A2 => n28184, B1 => n783, B2 => 
                           n7607, ZN => n19115);
   U13927 : NOR2_X2 port map( A1 => n27862, A2 => n5218, ZN => n17980);
   U13931 : XOR2_X1 port map( A1 => n2873, A2 => n18301, Z => n2690);
   U13974 : INV_X2 port map( I => n25497, ZN => n17047);
   U13982 : NOR2_X1 port map( A1 => n26068, A2 => n25596, ZN => n4114);
   U13987 : NOR2_X1 port map( A1 => n19899, A2 => n19901, ZN => n8562);
   U13991 : NAND2_X1 port map( A1 => n17541, A2 => n17472, ZN => n13280);
   U13993 : INV_X1 port map( I => n13887, ZN => n25726);
   U13994 : NAND3_X1 port map( A1 => n11494, A2 => n3014, A3 => n25726, ZN => 
                           n22576);
   U14000 : NAND2_X2 port map( A1 => n20231, A2 => n25440, ZN => n20452);
   U14002 : AOI21_X1 port map( A1 => n21799, A2 => n25441, B => n15203, ZN => 
                           n3429);
   U14005 : XOR2_X1 port map( A1 => n22504, A2 => n22541, Z => n25442);
   U14008 : NAND2_X2 port map( A1 => n10767, A2 => n26659, ZN => n7265);
   U14011 : XOR2_X1 port map( A1 => n12580, A2 => n7268, Z => n19691);
   U14031 : NAND2_X2 port map( A1 => n3793, A2 => n25448, ZN => n3792);
   U14032 : NOR2_X1 port map( A1 => n2706, A2 => n25455, ZN => n26189);
   U14038 : AOI22_X2 port map( A1 => n17151, A2 => n764, B1 => n17216, B2 => 
                           n17472, ZN => n25449);
   U14040 : INV_X2 port map( I => n25450, ZN => n13900);
   U14046 : OR2_X1 port map( A1 => n18646, A2 => n5115, Z => n13160);
   U14048 : XOR2_X1 port map( A1 => n15242, A2 => n22755, Z => n22340);
   U14049 : NAND2_X2 port map( A1 => n3047, A2 => n20001, ZN => n22755);
   U14059 : NOR2_X2 port map( A1 => n12257, A2 => n5425, ZN => n12621);
   U14063 : AOI21_X2 port map( A1 => n4800, A2 => n4799, B => n23188, ZN => 
                           n12257);
   U14066 : OAI21_X2 port map( A1 => n25453, A2 => n17980, B => n25688, ZN => 
                           n26248);
   U14068 : NOR2_X2 port map( A1 => n17881, A2 => n25, ZN => n25453);
   U14069 : NAND2_X2 port map( A1 => n24162, A2 => n17358, ZN => n15121);
   U14072 : NAND2_X2 port map( A1 => n11541, A2 => n11542, ZN => n12533);
   U14084 : XOR2_X1 port map( A1 => n21142, A2 => n11279, Z => n22719);
   U14088 : XOR2_X1 port map( A1 => n17136, A2 => n22631, Z => n25485);
   U14090 : OAI21_X2 port map( A1 => n19678, A2 => n671, B => n19587, ZN => 
                           n15009);
   U14097 : NAND3_X2 port map( A1 => n26679, A2 => n21095, A3 => n15721, ZN => 
                           n12057);
   U14098 : INV_X1 port map( I => n25458, ZN => n25457);
   U14099 : NOR2_X1 port map( A1 => n15787, A2 => n25373, ZN => n25458);
   U14100 : NAND2_X2 port map( A1 => n25459, A2 => n13574, ZN => n20875);
   U14103 : NAND2_X2 port map( A1 => n25460, A2 => n22990, ZN => n7039);
   U14109 : NAND2_X2 port map( A1 => n25461, A2 => n15645, ZN => n16700);
   U14113 : AND2_X1 port map( A1 => n15643, A2 => n15847, Z => n25461);
   U14115 : NOR2_X2 port map( A1 => n7921, A2 => n16710, ZN => n11684);
   U14128 : INV_X2 port map( I => n25465, ZN => n26154);
   U14132 : NAND2_X2 port map( A1 => n6743, A2 => n25466, ZN => n14792);
   U14134 : OR2_X1 port map( A1 => n7180, A2 => n22614, Z => n16430);
   U14154 : INV_X2 port map( I => n6030, ZN => n18782);
   U14155 : XOR2_X1 port map( A1 => n22940, A2 => n18131, Z => n6030);
   U14157 : AND2_X1 port map( A1 => n25717, A2 => n25254, Z => n25779);
   U14158 : XOR2_X1 port map( A1 => n8957, A2 => n1319, Z => n25781);
   U14160 : XOR2_X1 port map( A1 => n18172, A2 => n13996, Z => n18230);
   U14164 : INV_X2 port map( I => n75, ZN => n25468);
   U14176 : AND2_X1 port map( A1 => n9285, A2 => n632, Z => n13486);
   U14178 : XOR2_X1 port map( A1 => n25469, A2 => n14848, Z => n21443);
   U14180 : XOR2_X1 port map( A1 => n21370, A2 => n14850, Z => n25469);
   U14183 : NAND2_X2 port map( A1 => n25470, A2 => n15091, ZN => n19462);
   U14185 : NAND2_X1 port map( A1 => n18655, A2 => n9354, ZN => n25470);
   U14192 : XOR2_X1 port map( A1 => n18099, A2 => n20908, Z => n5872);
   U14208 : XOR2_X1 port map( A1 => n25474, A2 => n11965, Z => n13610);
   U14214 : AOI21_X2 port map( A1 => n14532, A2 => n13245, B => n23507, ZN => 
                           n25904);
   U14217 : OAI21_X2 port map( A1 => n5603, A2 => n1647, B => n1644, ZN => 
                           n2025);
   U14220 : AND2_X1 port map( A1 => n25896, A2 => n9133, Z => n9469);
   U14239 : AOI22_X2 port map( A1 => n25542, A2 => n14826, B1 => n4192, B2 => 
                           n28104, ZN => n4972);
   U14242 : NAND2_X1 port map( A1 => n16028, A2 => n7282, ZN => n25478);
   U14243 : NAND2_X1 port map( A1 => n10575, A2 => n1059, ZN => n25479);
   U14254 : XOR2_X1 port map( A1 => n20436, A2 => n20873, Z => n8579);
   U14275 : XOR2_X1 port map( A1 => n25481, A2 => n14340, Z => Ciphertext(93));
   U14281 : AOI21_X2 port map( A1 => n19022, A2 => n19021, B => n18929, ZN => 
                           n11239);
   U14288 : AND2_X1 port map( A1 => n4380, A2 => n799, Z => n25484);
   U14289 : XOR2_X1 port map( A1 => n2065, A2 => n25485, Z => n3296);
   U14304 : BUF_X2 port map( I => n10868, Z => n25487);
   U14309 : XOR2_X1 port map( A1 => n11513, A2 => n11511, Z => n22845);
   U14313 : XOR2_X1 port map( A1 => n11512, A2 => n10852, Z => n11511);
   U14320 : NAND2_X2 port map( A1 => n16994, A2 => n16995, ZN => n17580);
   U14323 : NAND2_X1 port map( A1 => n10366, A2 => n6247, ZN => n6246);
   U14341 : NAND2_X2 port map( A1 => n8035, A2 => n25491, ZN => n8032);
   U14342 : XOR2_X1 port map( A1 => n12411, A2 => n22761, Z => n2620);
   U14345 : NAND2_X2 port map( A1 => n3873, A2 => n3872, ZN => n22761);
   U14350 : INV_X1 port map( I => n26626, ZN => n25799);
   U14356 : XOR2_X1 port map( A1 => n4159, A2 => n6276, Z => n5391);
   U14359 : AND2_X1 port map( A1 => n3850, A2 => n16201, Z => n8834);
   U14377 : AOI22_X2 port map( A1 => n5759, A2 => n18465, B1 => n5642, B2 => 
                           n23199, ZN => n23302);
   U14380 : AND2_X1 port map( A1 => n7181, A2 => n19864, Z => n19642);
   U14381 : BUF_X2 port map( I => n1243, Z => n25498);
   U14387 : INV_X1 port map( I => n18510, ZN => n18511);
   U14388 : NAND2_X2 port map( A1 => n25769, A2 => n23062, ZN => n18510);
   U14393 : NAND2_X2 port map( A1 => n7618, A2 => n20339, ZN => n20099);
   U14396 : AOI21_X2 port map( A1 => n1961, A2 => n1960, B => n23899, ZN => 
                           n22757);
   U14404 : NOR2_X2 port map( A1 => n1959, A2 => n24306, ZN => n23899);
   U14412 : OAI21_X2 port map( A1 => n18371, A2 => n18381, B => n4198, ZN => 
                           n7939);
   U14418 : INV_X2 port map( I => n2989, ZN => n25500);
   U14419 : NAND2_X1 port map( A1 => n21628, A2 => n21627, ZN => n6567);
   U14425 : NOR2_X2 port map( A1 => n14406, A2 => n13426, ZN => n21628);
   U14440 : XOR2_X1 port map( A1 => n2140, A2 => n25333, Z => n26584);
   U14450 : INV_X2 port map( I => n25503, ZN => n19775);
   U14469 : INV_X2 port map( I => n25506, ZN => n26081);
   U14482 : XNOR2_X1 port map( A1 => n16948, A2 => n13403, ZN => n25506);
   U14485 : BUF_X2 port map( I => n11391, Z => n25508);
   U14495 : NAND3_X1 port map( A1 => n24026, A2 => n27889, A3 => n19800, ZN => 
                           n25511);
   U14512 : XOR2_X1 port map( A1 => n5914, A2 => n14572, Z => n20410);
   U14517 : NAND2_X1 port map( A1 => n17794, A2 => n25688, ZN => n25524);
   U14521 : INV_X4 port map( I => n8512, ZN => n26262);
   U14526 : XOR2_X1 port map( A1 => n25520, A2 => n19179, Z => n15740);
   U14529 : XOR2_X1 port map( A1 => n5026, A2 => n21375, Z => n5013);
   U14530 : XOR2_X1 port map( A1 => n24577, A2 => n6535, Z => n21375);
   U14538 : XOR2_X1 port map( A1 => n22829, A2 => n4310, Z => n12646);
   U14539 : AOI21_X1 port map( A1 => n9578, A2 => n21527, B => n25523, ZN => 
                           n9576);
   U14540 : OAI22_X1 port map( A1 => n9577, A2 => n21526, B1 => n770, B2 => 
                           n21525, ZN => n25523);
   U14545 : NAND2_X1 port map( A1 => n13489, A2 => n19081, ZN => n25526);
   U14551 : NOR2_X1 port map( A1 => n15352, A2 => n21690, ZN => n2161);
   U14561 : NAND2_X2 port map( A1 => n128, A2 => n22576, ZN => n3372);
   U14570 : INV_X4 port map( I => n7132, ZN => n905);
   U14571 : NAND2_X2 port map( A1 => n2497, A2 => n2496, ZN => n7132);
   U14585 : XOR2_X1 port map( A1 => n25528, A2 => n3601, Z => n9916);
   U14597 : NOR2_X1 port map( A1 => n935, A2 => n6323, ZN => n20802);
   U14599 : NAND2_X2 port map( A1 => n24112, A2 => n25846, ZN => n6323);
   U14601 : NAND2_X1 port map( A1 => n21943, A2 => n17783, ZN => n15532);
   U14603 : NAND2_X1 port map( A1 => n1431, A2 => n21006, ZN => n2427);
   U14605 : XOR2_X1 port map( A1 => n25343, A2 => n20941, Z => n15329);
   U14606 : NAND3_X1 port map( A1 => n16557, A2 => n26396, A3 => n13786, ZN => 
                           n1984);
   U14608 : XOR2_X1 port map( A1 => n8149, A2 => n10460, Z => n8386);
   U14613 : XOR2_X1 port map( A1 => n26922, A2 => n27969, Z => n25533);
   U14617 : NAND2_X2 port map( A1 => n25534, A2 => n16542, ZN => n16938);
   U14618 : OAI21_X2 port map( A1 => n24540, A2 => n25723, B => n25498, ZN => 
                           n25534);
   U14621 : XOR2_X1 port map( A1 => n25535, A2 => n5653, Z => n7592);
   U14625 : NAND2_X1 port map( A1 => n7595, A2 => n7594, ZN => n25535);
   U14626 : INV_X2 port map( I => n25536, ZN => n11805);
   U14629 : NAND3_X2 port map( A1 => n9668, A2 => n9667, A3 => n4068, ZN => 
                           n14753);
   U14638 : XNOR2_X1 port map( A1 => n25371, A2 => n20584, ZN => n25601);
   U14652 : INV_X2 port map( I => n26257, ZN => n19923);
   U14655 : NAND2_X1 port map( A1 => n19645, A2 => n26257, ZN => n19922);
   U14656 : XOR2_X1 port map( A1 => n4896, A2 => n25540, Z => n4893);
   U14658 : XOR2_X1 port map( A1 => n4895, A2 => n15537, Z => n25540);
   U14659 : XOR2_X1 port map( A1 => n25541, A2 => n10458, Z => n3895);
   U14663 : NAND2_X2 port map( A1 => n23466, A2 => n13499, ZN => n25966);
   U14665 : XNOR2_X1 port map( A1 => n12691, A2 => n11655, ZN => n25998);
   U14671 : OAI21_X2 port map( A1 => n2542, A2 => n12058, B => n2540, ZN => 
                           n19480);
   U14677 : XOR2_X1 port map( A1 => n9339, A2 => n25632, Z => n14129);
   U14684 : AOI21_X2 port map( A1 => n11577, A2 => n18895, B => n25411, ZN => 
                           n25545);
   U14713 : OR2_X2 port map( A1 => n25644, A2 => n26323, Z => n19766);
   U14720 : NAND2_X2 port map( A1 => n18692, A2 => n25548, ZN => n18798);
   U14735 : XOR2_X1 port map( A1 => n20521, A2 => n1536, Z => n1535);
   U14740 : XOR2_X1 port map( A1 => n27410, A2 => n25551, Z => n10887);
   U14742 : NAND2_X1 port map( A1 => n10890, A2 => n10889, ZN => n25551);
   U14759 : XOR2_X1 port map( A1 => n4893, A2 => n4897, Z => n20777);
   U14772 : NAND2_X2 port map( A1 => n10181, A2 => n10182, ZN => n11373);
   U14782 : NAND2_X2 port map( A1 => n12754, A2 => n25552, ZN => n12759);
   U14786 : NAND2_X2 port map( A1 => n25553, A2 => n16626, ZN => n16930);
   U14790 : NAND2_X2 port map( A1 => n15864, A2 => n25599, ZN => n16010);
   U14796 : NAND2_X1 port map( A1 => n12391, A2 => n24617, ZN => n12463);
   U14813 : NOR2_X2 port map( A1 => n764, A2 => n6977, ZN => n25560);
   U14822 : NAND2_X2 port map( A1 => n25563, A2 => n12996, ZN => n2516);
   U14826 : XOR2_X1 port map( A1 => n25564, A2 => n20344, Z => n21309);
   U14834 : NAND3_X2 port map( A1 => n10073, A2 => n10074, A3 => n17767, ZN => 
                           n18072);
   U14836 : XOR2_X1 port map( A1 => n20771, A2 => n20773, Z => n21370);
   U14838 : XOR2_X1 port map( A1 => n28510, A2 => n21281, Z => n7726);
   U14839 : NOR2_X2 port map( A1 => n21409, A2 => n13741, ZN => n21407);
   U14844 : XOR2_X1 port map( A1 => n18269, A2 => n633, Z => n8039);
   U14861 : OAI21_X2 port map( A1 => n9157, A2 => n9162, B => n9156, ZN => 
                           n23120);
   U14865 : NAND2_X2 port map( A1 => n18640, A2 => n18748, ZN => n8126);
   U14866 : OAI21_X1 port map( A1 => n9934, A2 => n24574, B => n25566, ZN => 
                           n21556);
   U14874 : NAND3_X2 port map( A1 => n25571, A2 => n2074, A3 => n3509, ZN => 
                           n3506);
   U14883 : XOR2_X1 port map( A1 => n12258, A2 => n25572, Z => n12221);
   U14888 : XOR2_X1 port map( A1 => n18283, A2 => n5314, Z => n25572);
   U14897 : BUF_X2 port map( I => n26076, Z => n25576);
   U14898 : XOR2_X1 port map( A1 => n17033, A2 => n25577, Z => n12341);
   U14900 : XOR2_X1 port map( A1 => n26082, A2 => n14782, Z => n25577);
   U14901 : INV_X2 port map( I => n25579, ZN => n8937);
   U14902 : XOR2_X1 port map( A1 => n8938, A2 => n13784, Z => n25579);
   U14906 : OAI21_X2 port map( A1 => n25874, A2 => n23380, B => n4771, ZN => 
                           n25795);
   U14907 : INV_X2 port map( I => n23107, ZN => n26298);
   U14912 : NAND2_X2 port map( A1 => n5678, A2 => n5676, ZN => n25679);
   U14913 : NAND2_X2 port map( A1 => n25584, A2 => n15300, ZN => n19565);
   U14915 : INV_X2 port map( I => n25585, ZN => n18776);
   U14916 : XOR2_X1 port map( A1 => n12853, A2 => n12855, Z => n25585);
   U14917 : XOR2_X1 port map( A1 => n511, A2 => n19289, Z => n26066);
   U14919 : XOR2_X1 port map( A1 => n22120, A2 => n19480, Z => n19289);
   U14920 : XOR2_X1 port map( A1 => n4777, A2 => n18076, Z => n7902);
   U14921 : AOI21_X2 port map( A1 => n2248, A2 => n6050, B => n15338, ZN => 
                           n12532);
   U14937 : NAND2_X1 port map( A1 => n12879, A2 => n16599, ZN => n25590);
   U14940 : NAND2_X1 port map( A1 => n23454, A2 => n20374, ZN => n26078);
   U14949 : NOR2_X2 port map( A1 => n2726, A2 => n22894, ZN => n25591);
   U14957 : XOR2_X1 port map( A1 => n24115, A2 => n11667, Z => n6777);
   U14968 : XOR2_X1 port map( A1 => n7885, A2 => n7882, Z => n22819);
   U14974 : XOR2_X1 port map( A1 => n7884, A2 => n7883, Z => n7882);
   U14982 : NAND2_X2 port map( A1 => n22425, A2 => n11431, ZN => n237);
   U14983 : XOR2_X1 port map( A1 => n13803, A2 => n13802, Z => n26342);
   U14985 : NAND2_X2 port map( A1 => n7012, A2 => n25595, ZN => n9161);
   U14986 : AOI22_X1 port map( A1 => n9026, A2 => n13422, B1 => n1108, B2 => 
                           n3016, ZN => n25595);
   U14987 : OAI21_X2 port map( A1 => n19737, A2 => n2792, B => n2791, ZN => 
                           n12986);
   U14988 : XOR2_X1 port map( A1 => n1776, A2 => n18189, Z => n26416);
   U14989 : INV_X2 port map( I => n25596, ZN => n15822);
   U14991 : XNOR2_X1 port map( A1 => Key(83), A2 => Plaintext(83), ZN => n25596
                           );
   U14992 : XOR2_X1 port map( A1 => n19357, A2 => n19469, Z => n8800);
   U14997 : AOI21_X2 port map( A1 => n25597, A2 => n15790, B => n23135, ZN => 
                           n16707);
   U15006 : NAND2_X2 port map( A1 => n20237, A2 => n20043, ZN => n25598);
   U15007 : OR2_X1 port map( A1 => n11763, A2 => n28490, Z => n11572);
   U15009 : OAI22_X2 port map( A1 => n1911, A2 => n15921, B1 => n21814, B2 => 
                           n1908, ZN => n8722);
   U15011 : XOR2_X1 port map( A1 => n1676, A2 => n25600, Z => n26176);
   U15012 : XOR2_X1 port map( A1 => n18164, A2 => n25601, Z => n25600);
   U15029 : XOR2_X1 port map( A1 => n18152, A2 => n25604, Z => n10077);
   U15031 : XOR2_X1 port map( A1 => n24357, A2 => n27410, Z => n25604);
   U15037 : NAND2_X1 port map( A1 => n28538, A2 => n613, ZN => n25605);
   U15045 : INV_X2 port map( I => n25606, ZN => n26624);
   U15061 : AOI21_X2 port map( A1 => n1459, A2 => n26624, B => n19801, ZN => 
                           n25635);
   U15062 : INV_X2 port map( I => n17475, ZN => n25608);
   U15067 : INV_X2 port map( I => n25611, ZN => n17123);
   U15074 : XOR2_X1 port map( A1 => n17035, A2 => n16929, Z => n25611);
   U15079 : NAND2_X2 port map( A1 => n15425, A2 => n24373, ZN => n13070);
   U15090 : NAND3_X1 port map( A1 => n18080, A2 => n10263, A3 => n22547, ZN => 
                           n13617);
   U15105 : XOR2_X1 port map( A1 => n25948, A2 => n25616, Z => n15670);
   U15112 : XOR2_X1 port map( A1 => n25617, A2 => n19235, Z => n4582);
   U15113 : XOR2_X1 port map( A1 => n25618, A2 => n26358, Z => n11785);
   U15126 : NOR2_X2 port map( A1 => n17889, A2 => n17888, ZN => n25946);
   U15128 : OR2_X1 port map( A1 => n26293, A2 => n24025, Z => n308);
   U15135 : XOR2_X1 port map( A1 => n25622, A2 => n17105, Z => n5862);
   U15142 : NAND2_X2 port map( A1 => n22977, A2 => n18640, ZN => n18746);
   U15155 : NAND2_X2 port map( A1 => n25455, A2 => n10007, ZN => n22672);
   U15156 : AOI21_X2 port map( A1 => n3545, A2 => n25624, B => n1029, ZN => 
                           n24345);
   U15158 : NAND2_X2 port map( A1 => n125, A2 => n123, ZN => n25626);
   U15162 : OAI21_X1 port map( A1 => n20876, A2 => n27468, B => n13553, ZN => 
                           n11640);
   U15173 : NAND2_X2 port map( A1 => n11869, A2 => n20875, ZN => n13553);
   U15188 : XOR2_X1 port map( A1 => n25166, A2 => n19500, Z => n25627);
   U15221 : NAND2_X1 port map( A1 => n20665, A2 => n4934, ZN => n20657);
   U15225 : NAND2_X2 port map( A1 => n23546, A2 => n7569, ZN => n8226);
   U15243 : NOR2_X2 port map( A1 => n3853, A2 => n3854, ZN => n7281);
   U15252 : NAND2_X2 port map( A1 => n5779, A2 => n5780, ZN => n6718);
   U15258 : XOR2_X1 port map( A1 => n13825, A2 => n19233, Z => n25632);
   U15271 : INV_X4 port map( I => n24482, ZN => n4705);
   U15272 : NAND2_X2 port map( A1 => n4704, A2 => n24483, ZN => n24482);
   U15276 : XOR2_X1 port map( A1 => n25000, A2 => n9722, Z => n25633);
   U15289 : XOR2_X1 port map( A1 => n28233, A2 => n25333, Z => n25634);
   U15291 : XOR2_X1 port map( A1 => n20763, A2 => n25636, Z => n21180);
   U15293 : XOR2_X1 port map( A1 => n8736, A2 => n5174, Z => n3083);
   U15295 : XOR2_X1 port map( A1 => n12410, A2 => n10773, Z => n17062);
   U15297 : NAND3_X1 port map( A1 => n18749, A2 => n18640, A3 => n14362, ZN => 
                           n18501);
   U15308 : NAND3_X2 port map( A1 => n13880, A2 => n5298, A3 => n17218, ZN => 
                           n11497);
   U15315 : AOI22_X2 port map( A1 => n4885, A2 => n26532, B1 => n4252, B2 => 
                           n17522, ZN => n22603);
   U15318 : NOR2_X2 port map( A1 => n5612, A2 => n900, ZN => n4252);
   U15321 : OAI22_X1 port map( A1 => n4245, A2 => n1219, B1 => n890, B2 => 
                           n8849, ZN => n26504);
   U15323 : NAND2_X1 port map( A1 => n17337, A2 => n16972, ZN => n5222);
   U15325 : XOR2_X1 port map( A1 => n22969, A2 => n23998, Z => n17337);
   U15351 : NAND2_X1 port map( A1 => n4499, A2 => n19878, ZN => n25639);
   U15358 : NOR2_X2 port map( A1 => n17803, A2 => n27458, ZN => n25640);
   U15360 : NAND2_X2 port map( A1 => n25641, A2 => n17819, ZN => n24126);
   U15367 : XOR2_X1 port map( A1 => n13514, A2 => n16911, Z => n23735);
   U15368 : XOR2_X1 port map( A1 => n12147, A2 => n4179, Z => n16911);
   U15370 : XOR2_X1 port map( A1 => n7896, A2 => n20577, Z => n7391);
   U15377 : NAND2_X2 port map( A1 => n15093, A2 => n18838, ZN => n19412);
   U15379 : OAI22_X2 port map( A1 => n9474, A2 => n13159, B1 => n25355, B2 => 
                           n18764, ZN => n5511);
   U15385 : XNOR2_X1 port map( A1 => n220, A2 => n25762, ZN => n25644);
   U15389 : NAND2_X1 port map( A1 => n21741, A2 => n27471, ZN => n25645);
   U15393 : NAND2_X2 port map( A1 => n18684, A2 => n18685, ZN => n8619);
   U15395 : OAI21_X1 port map( A1 => n14306, A2 => n14415, B => n12125, ZN => 
                           n3794);
   U15398 : NAND2_X1 port map( A1 => n21087, A2 => n22796, ZN => n9863);
   U15399 : NOR2_X1 port map( A1 => n20655, A2 => n4766, ZN => n25646);
   U15402 : OAI21_X2 port map( A1 => n23223, A2 => n23222, B => n10631, ZN => 
                           n20459);
   U15405 : XOR2_X1 port map( A1 => n4956, A2 => n5625, Z => n25647);
   U15406 : NAND2_X2 port map( A1 => n4122, A2 => n15103, ZN => n20647);
   U15407 : OAI21_X1 port map( A1 => n844, A2 => n20663, B => n3824, ZN => 
                           n8481);
   U15414 : INV_X2 port map( I => n8937, ZN => n25650);
   U15418 : XOR2_X1 port map( A1 => n19374, A2 => n19372, Z => n8938);
   U15443 : XOR2_X1 port map( A1 => n25652, A2 => n1302, Z => Ciphertext(188));
   U15455 : OAI22_X1 port map( A1 => n7384, A2 => n26647, B1 => n10975, B2 => 
                           n21738, ZN => n25652);
   U15461 : OAI21_X1 port map( A1 => n19930, A2 => n11354, B => n27452, ZN => 
                           n11093);
   U15468 : INV_X2 port map( I => n19397, ZN => n19930);
   U15473 : XOR2_X1 port map( A1 => n13132, A2 => n13130, Z => n24289);
   U15475 : INV_X1 port map( I => n22365, ZN => n7611);
   U15479 : INV_X2 port map( I => n5722, ZN => n10797);
   U15482 : NAND2_X1 port map( A1 => n25799, A2 => n5722, ZN => n21691);
   U15483 : NAND2_X2 port map( A1 => n22170, A2 => n6048, ZN => n6050);
   U15487 : NAND2_X2 port map( A1 => n25653, A2 => n9786, ZN => n16651);
   U15489 : OAI21_X2 port map( A1 => n15830, A2 => n15829, B => n15926, ZN => 
                           n25653);
   U15492 : XOR2_X1 port map( A1 => n16521, A2 => n16520, Z => n26386);
   U15498 : XOR2_X1 port map( A1 => n26449, A2 => n16801, Z => n16521);
   U15504 : XOR2_X1 port map( A1 => n25654, A2 => n15400, Z => n17419);
   U15505 : XOR2_X1 port map( A1 => n6137, A2 => n16854, Z => n25654);
   U15511 : NAND3_X1 port map( A1 => n25753, A2 => n24874, A3 => n21355, ZN => 
                           n23800);
   U15512 : NOR3_X1 port map( A1 => n17906, A2 => n17665, A3 => n24127, ZN => 
                           n12169);
   U15513 : AOI21_X2 port map( A1 => n17406, A2 => n17405, B => n17404, ZN => 
                           n17906);
   U15520 : XOR2_X1 port map( A1 => n21182, A2 => n20475, Z => n20477);
   U15527 : XOR2_X1 port map( A1 => n20479, A2 => n20478, Z => n20631);
   U15541 : XOR2_X1 port map( A1 => n23022, A2 => n10382, Z => n22330);
   U15548 : NAND2_X2 port map( A1 => n26043, A2 => n4495, ZN => n172);
   U15550 : NAND2_X2 port map( A1 => n25671, A2 => n8373, ZN => n22273);
   U15557 : XOR2_X1 port map( A1 => n10669, A2 => n336, Z => n25674);
   U15575 : XOR2_X1 port map( A1 => n17045, A2 => n3945, Z => n58);
   U15593 : XOR2_X1 port map( A1 => n25677, A2 => n25676, Z => n21907);
   U15594 : XOR2_X1 port map( A1 => n18106, A2 => n22802, Z => n25676);
   U15600 : NAND2_X2 port map( A1 => n2420, A2 => n9470, ZN => n2820);
   U15618 : XOR2_X1 port map( A1 => n26443, A2 => n18360, Z => n25681);
   U15625 : NAND2_X2 port map( A1 => n21958, A2 => n21957, ZN => n23474);
   U15631 : NOR2_X1 port map( A1 => n22727, A2 => n8290, ZN => n21841);
   U15647 : XOR2_X1 port map( A1 => n4029, A2 => n4031, Z => n16998);
   U15660 : NAND2_X2 port map( A1 => n25713, A2 => n9400, ZN => n11756);
   U15672 : OAI21_X2 port map( A1 => n26672, A2 => n23501, B => n25687, ZN => 
                           n12946);
   U15683 : AOI21_X2 port map( A1 => n12162, A2 => n23126, B => n25689, ZN => 
                           n26392);
   U15684 : NOR2_X2 port map( A1 => n18974, A2 => n11331, ZN => n25689);
   U15693 : NAND2_X2 port map( A1 => n18810, A2 => n14338, ZN => n18974);
   U15698 : NOR2_X2 port map( A1 => n19582, A2 => n23444, ZN => n26461);
   U15705 : NAND2_X2 port map( A1 => n26399, A2 => n23445, ZN => n23444);
   U15719 : NAND2_X2 port map( A1 => n25694, A2 => n17290, ZN => n17761);
   U15720 : XOR2_X1 port map( A1 => n13891, A2 => n18234, Z => n18214);
   U15721 : AOI22_X1 port map( A1 => n21407, A2 => n21408, B1 => n11466, B2 => 
                           n21409, ZN => n25977);
   U15728 : OAI21_X1 port map( A1 => n10371, A2 => n10372, B => n25977, ZN => 
                           n10370);
   U15734 : NAND2_X1 port map( A1 => n26638, A2 => n7611, ZN => n15265);
   U15741 : INV_X2 port map( I => n16612, ZN => n25698);
   U15748 : XOR2_X1 port map( A1 => n25699, A2 => n24384, Z => n6530);
   U15751 : XOR2_X1 port map( A1 => n8132, A2 => n12114, Z => n25699);
   U15762 : OAI21_X2 port map( A1 => n25498, A2 => n6131, B => n4217, ZN => 
                           n4877);
   U15769 : AND2_X1 port map( A1 => n26620, A2 => n26624, Z => n11516);
   U15787 : XOR2_X1 port map( A1 => n4533, A2 => n22313, Z => n5506);
   U15788 : AND2_X1 port map( A1 => n7176, A2 => n19605, Z => n19606);
   U15792 : INV_X2 port map( I => n20376, ZN => n5520);
   U15795 : XOR2_X1 port map( A1 => n9802, A2 => n18112, Z => n18212);
   U15796 : NAND2_X2 port map( A1 => n14904, A2 => n14903, ZN => n18112);
   U15799 : XOR2_X1 port map( A1 => n16739, A2 => n16740, Z => n16741);
   U15819 : NAND2_X1 port map( A1 => n14339, A2 => n24215, ZN => n5685);
   U15828 : AOI21_X2 port map( A1 => n23623, A2 => n21777, B => n4038, ZN => 
                           n25707);
   U15829 : NAND2_X2 port map( A1 => n21499, A2 => n14525, ZN => n21496);
   U15850 : AND3_X1 port map( A1 => n4191, A2 => n25710, A3 => n9525, Z => 
                           n25790);
   U15860 : AOI22_X2 port map( A1 => n20928, A2 => n28197, B1 => n10350, B2 => 
                           n7956, ZN => n25727);
   U15861 : NOR2_X2 port map( A1 => n28198, A2 => n26001, ZN => n20928);
   U15868 : XOR2_X1 port map( A1 => n13895, A2 => n13894, Z => n13896);
   U15883 : INV_X2 port map( I => n26461, ZN => n21932);
   U15889 : NAND2_X1 port map( A1 => n26461, A2 => n22398, ZN => n25717);
   U15894 : NAND2_X1 port map( A1 => n5459, A2 => n12428, ZN => n25811);
   U15895 : OAI21_X2 port map( A1 => n23743, A2 => n14308, B => n8254, ZN => 
                           n25718);
   U15904 : NOR2_X1 port map( A1 => n21622, A2 => n21624, ZN => n25721);
   U15914 : NOR2_X2 port map( A1 => n22737, A2 => n25841, ZN => n4581);
   U15923 : XOR2_X1 port map( A1 => n19482, A2 => n22381, Z => n11174);
   U15926 : NAND2_X2 port map( A1 => n12750, A2 => n12751, ZN => n19482);
   U15945 : AOI21_X1 port map( A1 => n15513, A2 => n15374, B => n1699, ZN => 
                           n12172);
   U15958 : AOI22_X2 port map( A1 => n8772, A2 => n19956, B1 => n19634, B2 => 
                           n20150, ZN => n21249);
   U15964 : XOR2_X1 port map( A1 => n7745, A2 => n18179, Z => n7744);
   U15968 : NAND2_X2 port map( A1 => n10462, A2 => n17625, ZN => n18179);
   U15971 : XOR2_X1 port map( A1 => n12908, A2 => n12907, Z => n5445);
   U15973 : OAI21_X2 port map( A1 => n10351, A2 => n20887, B => n25727, ZN => 
                           n2588);
   U15974 : NAND2_X2 port map( A1 => n9705, A2 => n25728, ZN => n16585);
   U15975 : OAI21_X2 port map( A1 => n4810, A2 => n12614, B => n25729, ZN => 
                           n14896);
   U15977 : NAND2_X2 port map( A1 => n1115, A2 => n4810, ZN => n25729);
   U15978 : INV_X2 port map( I => n25730, ZN => n5140);
   U15980 : XOR2_X1 port map( A1 => Plaintext(144), A2 => Key(144), Z => n25730
                           );
   U15988 : OAI21_X2 port map( A1 => n2512, A2 => n12339, B => n20050, ZN => 
                           n2511);
   U15997 : XOR2_X1 port map( A1 => n16822, A2 => n17090, Z => n16754);
   U15999 : NAND2_X2 port map( A1 => n2722, A2 => n26123, ZN => n17090);
   U16003 : XOR2_X1 port map( A1 => n17125, A2 => n21313, Z => n9536);
   U16005 : AOI21_X1 port map( A1 => n25745, A2 => n4726, B => n1071, ZN => 
                           n4725);
   U16007 : XOR2_X1 port map( A1 => n13115, A2 => n13113, Z => n13628);
   U16021 : XOR2_X1 port map( A1 => n18097, A2 => n25865, Z => n18267);
   U16030 : NOR2_X2 port map( A1 => n25740, A2 => n7356, ZN => n16875);
   U16037 : XOR2_X1 port map( A1 => n2664, A2 => n2665, Z => n25741);
   U16041 : XOR2_X1 port map( A1 => n17015, A2 => n14650, Z => n25744);
   U16042 : XOR2_X1 port map( A1 => n6996, A2 => n1638, Z => n21433);
   U16047 : AOI21_X2 port map( A1 => n9174, A2 => n8093, B => n2036, ZN => 
                           n25856);
   U16050 : OR2_X1 port map( A1 => n20910, A2 => n22803, Z => n25745);
   U16052 : INV_X2 port map( I => n6018, ZN => n11514);
   U16053 : XOR2_X1 port map( A1 => n19311, A2 => n19284, Z => n2176);
   U16062 : NAND2_X1 port map( A1 => n7782, A2 => n7783, ZN => n7781);
   U16063 : XOR2_X1 port map( A1 => n9982, A2 => n23799, Z => n25747);
   U16065 : XOR2_X1 port map( A1 => n22091, A2 => n8371, Z => n8370);
   U16067 : XOR2_X1 port map( A1 => n20409, A2 => n22761, Z => n25748);
   U16084 : NAND2_X2 port map( A1 => n26513, A2 => n8306, ZN => n11261);
   U16088 : XOR2_X1 port map( A1 => n28541, A2 => n24134, Z => n22686);
   U16090 : NOR2_X2 port map( A1 => n27372, A2 => n1681, ZN => n16481);
   U16091 : OAI22_X2 port map( A1 => n1543, A2 => n1544, B1 => n7053, B2 => 
                           n2543, ZN => n1681);
   U16094 : NOR2_X2 port map( A1 => n26430, A2 => n2293, ZN => n25751);
   U16095 : OR2_X1 port map( A1 => n5140, A2 => n8407, Z => n13123);
   U16105 : AOI22_X2 port map( A1 => n5883, A2 => n15067, B1 => n19890, B2 => 
                           n3986, ZN => n22011);
   U16109 : AOI22_X2 port map( A1 => n17691, A2 => n727, B1 => n3346, B2 => 
                           n17692, ZN => n25752);
   U16111 : NAND3_X1 port map( A1 => n929, A2 => n13009, A3 => n21113, ZN => 
                           n21102);
   U16125 : NAND2_X2 port map( A1 => n6315, A2 => n16266, ZN => n9970);
   U16148 : NOR2_X1 port map( A1 => n260, A2 => n4393, ZN => n25756);
   U16156 : NOR2_X2 port map( A1 => n25758, A2 => n25757, ZN => n16336);
   U16164 : OR2_X1 port map( A1 => n23875, A2 => n16323, Z => n25758);
   U16172 : XOR2_X1 port map( A1 => n10529, A2 => n13840, Z => n5971);
   U16173 : OAI21_X2 port map( A1 => n25760, A2 => n807, B => n25759, ZN => 
                           n23141);
   U16174 : INV_X2 port map( I => n25045, ZN => n25759);
   U16178 : XOR2_X1 port map( A1 => n981, A2 => n19477, Z => n7279);
   U16183 : XOR2_X1 port map( A1 => n8500, A2 => n12147, Z => n17106);
   U16184 : NAND2_X2 port map( A1 => n25761, A2 => n4561, ZN => n4558);
   U16193 : OR2_X2 port map( A1 => n8314, A2 => n17745, Z => n4508);
   U16196 : NAND2_X2 port map( A1 => n4225, A2 => n19967, ZN => n20011);
   U16205 : NAND2_X2 port map( A1 => n16003, A2 => n16002, ZN => n16957);
   U16226 : AND2_X1 port map( A1 => n14997, A2 => n613, Z => n5677);
   U16228 : OAI21_X2 port map( A1 => n24666, A2 => n11035, B => n15623, ZN => 
                           n4256);
   U16232 : AOI22_X2 port map( A1 => n13723, A2 => n17925, B1 => n17743, B2 => 
                           n17928, ZN => n25768);
   U16233 : BUF_X2 port map( I => n26494, Z => n25769);
   U16247 : OAI21_X1 port map( A1 => n16289, A2 => n6428, B => n13274, ZN => 
                           n25774);
   U16250 : AOI22_X2 port map( A1 => n21753, A2 => n23811, B1 => n4730, B2 => 
                           n1021, ZN => n10125);
   U16254 : INV_X2 port map( I => n10136, ZN => n4730);
   U16265 : XOR2_X1 port map( A1 => n18230, A2 => n18352, Z => n9558);
   U16276 : NAND2_X1 port map( A1 => n12292, A2 => n16604, ZN => n12092);
   U16277 : NAND2_X2 port map( A1 => n4113, A2 => n4116, ZN => n12292);
   U16283 : XOR2_X1 port map( A1 => n24012, A2 => n9054, Z => n9053);
   U16286 : XOR2_X1 port map( A1 => n1946, A2 => n1041, Z => n9054);
   U16293 : INV_X2 port map( I => n26323, ZN => n26625);
   U16299 : XOR2_X1 port map( A1 => n25780, A2 => n3941, Z => n3940);
   U16306 : XOR2_X1 port map( A1 => n9673, A2 => n25781, Z => n25780);
   U16308 : XOR2_X1 port map( A1 => n26085, A2 => n24654, Z => n25988);
   U16312 : XOR2_X1 port map( A1 => n20540, A2 => n21197, Z => n4866);
   U16313 : NAND2_X2 port map( A1 => n19980, A2 => n19979, ZN => n20540);
   U16329 : OR2_X1 port map( A1 => n5047, A2 => n675, Z => n19813);
   U16332 : OAI22_X2 port map( A1 => n1608, A2 => n1609, B1 => n1610, B2 => n45
                           , ZN => n5573);
   U16339 : NAND2_X2 port map( A1 => n21901, A2 => n17887, ZN => n17803);
   U16341 : OAI22_X1 port map( A1 => n25784, A2 => n22751, B1 => n21169, B2 => 
                           n25377, ZN => n500);
   U16347 : OAI21_X2 port map( A1 => n24426, A2 => n25902, B => n6978, ZN => 
                           n11680);
   U16360 : XOR2_X1 port map( A1 => n18356, A2 => n11682, Z => n11681);
   U16366 : NOR2_X1 port map( A1 => n6247, A2 => n9166, ZN => n8934);
   U16373 : NAND2_X2 port map( A1 => n23134, A2 => n7487, ZN => n16472);
   U16376 : NAND2_X2 port map( A1 => n9163, A2 => n24297, ZN => n2110);
   U16379 : OAI22_X2 port map( A1 => n18666, A2 => n18665, B1 => n18667, B2 => 
                           n1018, ZN => n9163);
   U16388 : NOR2_X2 port map( A1 => n12658, A2 => n25790, ZN => n12656);
   U16394 : NAND3_X1 port map( A1 => n20835, A2 => n20836, A3 => n20850, ZN => 
                           n25791);
   U16395 : XOR2_X1 port map( A1 => n25792, A2 => n14404, Z => n7707);
   U16396 : NAND3_X1 port map( A1 => n4596, A2 => n4595, A3 => n4597, ZN => 
                           n25793);
   U16404 : OAI22_X2 port map( A1 => n864, A2 => n26625, B1 => n9612, B2 => 
                           n19744, ZN => n19764);
   U16405 : XOR2_X1 port map( A1 => n25797, A2 => n23737, Z => n14844);
   U16414 : AND2_X1 port map( A1 => n17388, A2 => n26614, Z => n22275);
   U16438 : XOR2_X1 port map( A1 => n21377, A2 => n20568, Z => n14972);
   U16444 : XOR2_X1 port map( A1 => n11371, A2 => n20575, Z => n21377);
   U16445 : NOR2_X1 port map( A1 => n15655, A2 => n15656, ZN => n25800);
   U16448 : NAND2_X2 port map( A1 => n25801, A2 => n16371, ZN => n16801);
   U16464 : INV_X1 port map( I => n4265, ZN => n22019);
   U16470 : NAND2_X1 port map( A1 => n26640, A2 => n14580, ZN => n24497);
   U16475 : OR2_X1 port map( A1 => n16029, A2 => n24581, Z => n25804);
   U16493 : XOR2_X1 port map( A1 => n27400, A2 => n25807, Z => n24377);
   U16495 : XOR2_X1 port map( A1 => n19220, A2 => n25808, Z => n25807);
   U16499 : INV_X1 port map( I => n14630, ZN => n25808);
   U16527 : NAND2_X1 port map( A1 => n16231, A2 => n21904, ZN => n175);
   U16535 : NAND2_X2 port map( A1 => n25812, A2 => n18877, ZN => n19365);
   U16542 : NOR2_X2 port map( A1 => n26169, A2 => n1793, ZN => n13305);
   U16558 : NAND2_X2 port map( A1 => n13697, A2 => n20987, ZN => n21000);
   U16561 : NAND2_X2 port map( A1 => n12180, A2 => n26660, ZN => n13697);
   U16582 : OR2_X1 port map( A1 => n7612, A2 => n15228, Z => n1601);
   U16613 : NAND2_X2 port map( A1 => n3617, A2 => n3618, ZN => n19445);
   U16617 : XOR2_X1 port map( A1 => n24034, A2 => n23343, Z => n19615);
   U16620 : NAND2_X2 port map( A1 => n25818, A2 => n2927, ZN => n4147);
   U16626 : XOR2_X1 port map( A1 => n2554, A2 => n25819, Z => n24097);
   U16628 : XOR2_X1 port map( A1 => n4314, A2 => n28549, Z => n25819);
   U16631 : AOI21_X2 port map( A1 => n2163, A2 => n13174, B => n25821, ZN => 
                           n12581);
   U16638 : INV_X2 port map( I => n25822, ZN => n10707);
   U16640 : XOR2_X1 port map( A1 => Key(127), A2 => Plaintext(127), Z => n25822
                           );
   U16641 : NAND2_X2 port map( A1 => n25823, A2 => n18882, ZN => n19349);
   U16649 : NAND4_X2 port map( A1 => n12852, A2 => n13697, A3 => n20987, A4 => 
                           n12851, ZN => n12179);
   U16650 : NAND2_X2 port map( A1 => n20974, A2 => n731, ZN => n12852);
   U16651 : XOR2_X1 port map( A1 => n26486, A2 => n25824, Z => n15001);
   U16661 : OR2_X1 port map( A1 => n16413, A2 => n16712, Z => n9819);
   U16665 : AND2_X1 port map( A1 => n20041, A2 => n8100, Z => n25831);
   U16674 : OAI22_X1 port map( A1 => n16216, A2 => n16511, B1 => n16563, B2 => 
                           n16394, ZN => n16223);
   U16680 : INV_X1 port map( I => n11339, ZN => n26100);
   U16703 : NAND2_X2 port map( A1 => n9426, A2 => n3303, ZN => n10635);
   U16705 : AND2_X1 port map( A1 => n16704, A2 => n25834, Z => n22587);
   U16707 : AOI21_X1 port map( A1 => n25835, A2 => n12075, B => n9425, ZN => 
                           n12074);
   U16708 : NAND2_X1 port map( A1 => n21041, A2 => n27392, ZN => n25835);
   U16709 : NOR2_X1 port map( A1 => n17036, A2 => n14250, ZN => n17287);
   U16710 : XOR2_X1 port map( A1 => n17029, A2 => n14000, Z => n10826);
   U16711 : OAI21_X2 port map( A1 => n12419, A2 => n10789, B => n22054, ZN => 
                           n19004);
   U16716 : XOR2_X1 port map( A1 => n27623, A2 => n10529, Z => n17876);
   U16719 : OAI21_X2 port map( A1 => n7153, A2 => n11129, B => n11126, ZN => 
                           n10529);
   U16720 : XNOR2_X1 port map( A1 => n17028, A2 => n4877, ZN => n17127);
   U16726 : XOR2_X1 port map( A1 => n8441, A2 => n25838, Z => n22960);
   U16731 : XOR2_X1 port map( A1 => n3291, A2 => n7752, Z => n25838);
   U16733 : NAND3_X2 port map( A1 => n15479, A2 => n21071, A3 => n10687, ZN => 
                           n21082);
   U16734 : NAND2_X1 port map( A1 => n25504, A2 => n8125, ZN => n3335);
   U16748 : INV_X1 port map( I => n14503, ZN => n25840);
   U16749 : INV_X2 port map( I => n9671, ZN => n25841);
   U16753 : NAND2_X2 port map( A1 => n5512, A2 => n5513, ZN => n22253);
   U16765 : XOR2_X1 port map( A1 => n7437, A2 => n7435, Z => n17198);
   U16791 : NAND2_X2 port map( A1 => n12493, A2 => n18388, ZN => n7919);
   U16808 : XOR2_X1 port map( A1 => n19437, A2 => n19436, Z => n5398);
   U16817 : NAND3_X1 port map( A1 => n11132, A2 => n7682, A3 => n11078, ZN => 
                           n22376);
   U16824 : NAND3_X2 port map( A1 => n13047, A2 => n28400, A3 => n16660, ZN => 
                           n25845);
   U16826 : XOR2_X1 port map( A1 => n16895, A2 => n21341, Z => n7509);
   U16827 : NAND3_X2 port map( A1 => n24029, A2 => n300, A3 => n301, ZN => 
                           n16895);
   U16829 : NAND2_X1 port map( A1 => n20760, A2 => n27380, ZN => n25846);
   U16860 : NOR2_X2 port map( A1 => n17188, A2 => n1232, ZN => n14724);
   U16861 : INV_X2 port map( I => n22620, ZN => n17188);
   U16870 : XOR2_X1 port map( A1 => n19389, A2 => n19348, Z => n3734);
   U16871 : XOR2_X1 port map( A1 => n6309, A2 => n22768, Z => n19348);
   U16880 : NAND2_X2 port map( A1 => n2693, A2 => n1246, ZN => n3415);
   U16881 : XOR2_X1 port map( A1 => n18316, A2 => n18315, Z => n18321);
   U16887 : NAND3_X2 port map( A1 => n24606, A2 => n24230, A3 => n24605, ZN => 
                           n20052);
   U16888 : NOR2_X2 port map( A1 => n9939, A2 => n25852, ZN => n10627);
   U16892 : AOI22_X2 port map( A1 => n5631, A2 => n17722, B1 => n5630, B2 => 
                           n6794, ZN => n18077);
   U16896 : XOR2_X1 port map( A1 => n25855, A2 => n15195, Z => Ciphertext(172))
                           ;
   U16901 : XOR2_X1 port map( A1 => n9130, A2 => n9129, Z => n10971);
   U16902 : INV_X4 port map( I => n25857, ZN => n24524);
   U16906 : NOR2_X2 port map( A1 => n2946, A2 => n2944, ZN => n25857);
   U16912 : OAI21_X2 port map( A1 => n26544, A2 => n24599, B => n24479, ZN => 
                           n9430);
   U16915 : XOR2_X1 port map( A1 => n6308, A2 => n25859, Z => n24415);
   U16916 : XOR2_X1 port map( A1 => n2467, A2 => n22349, Z => n25859);
   U16920 : AOI21_X2 port map( A1 => n5818, A2 => n4735, B => n25861, ZN => 
                           n5817);
   U16935 : NAND3_X2 port map( A1 => n6928, A2 => n6927, A3 => n6931, ZN => 
                           n9414);
   U16936 : AOI22_X1 port map( A1 => n15766, A2 => n15998, B1 => n15767, B2 => 
                           n15995, ZN => n9405);
   U16937 : NAND3_X2 port map( A1 => n15701, A2 => n9759, A3 => n16731, ZN => 
                           n25862);
   U16944 : BUF_X2 port map( I => n25914, Z => n25864);
   U16963 : NAND3_X2 port map( A1 => n14008, A2 => n7113, A3 => n16671, ZN => 
                           n2708);
   U16964 : INV_X2 port map( I => n24531, ZN => n968);
   U16977 : XOR2_X1 port map( A1 => n6344, A2 => n15589, Z => n24531);
   U16978 : XOR2_X1 port map( A1 => n16990, A2 => n25866, Z => n1438);
   U16989 : XOR2_X1 port map( A1 => n26132, A2 => n20851, Z => n25866);
   U17010 : XOR2_X1 port map( A1 => n451, A2 => n21210, Z => n25867);
   U17014 : NOR3_X2 port map( A1 => n25868, A2 => n5375, A3 => n5376, ZN => 
                           n6019);
   U17018 : NOR3_X2 port map( A1 => n892, A2 => n898, A3 => n8093, ZN => n25868
                           );
   U17021 : AOI22_X2 port map( A1 => n25869, A2 => n309, B1 => n16548, B2 => 
                           n3741, ZN => n17843);
   U17028 : OAI21_X2 port map( A1 => n25871, A2 => n11171, B => n11170, ZN => 
                           n17745);
   U17031 : NAND2_X1 port map( A1 => n14318, A2 => n14317, ZN => n13618);
   U17045 : XOR2_X1 port map( A1 => n22126, A2 => n6108, Z => n2748);
   U17049 : XOR2_X1 port map( A1 => n11430, A2 => n3946, Z => n26067);
   U17057 : XOR2_X1 port map( A1 => n25877, A2 => n14335, Z => n7507);
   U17063 : XOR2_X1 port map( A1 => n7509, A2 => n25683, Z => n25877);
   U17073 : NOR2_X2 port map( A1 => n3839, A2 => n3836, ZN => n22602);
   U17085 : NAND2_X1 port map( A1 => n11983, A2 => n28237, ZN => n8377);
   U17086 : OAI21_X2 port map( A1 => n7274, A2 => n7518, B => n25881, ZN => 
                           n20746);
   U17092 : NAND3_X2 port map( A1 => n11642, A2 => n9265, A3 => n9266, ZN => 
                           n14586);
   U17101 : NOR2_X2 port map( A1 => n17315, A2 => n14250, ZN => n10913);
   U17107 : OR2_X1 port map( A1 => n2346, A2 => n26570, Z => n4544);
   U17124 : OAI21_X2 port map( A1 => n13765, A2 => n10908, B => n23745, ZN => 
                           n22194);
   U17135 : OAI22_X1 port map( A1 => n21632, A2 => n21647, B1 => n13908, B2 => 
                           n27390, ZN => n15217);
   U17136 : XOR2_X1 port map( A1 => n25889, A2 => n24266, Z => n14287);
   U17141 : XOR2_X1 port map( A1 => n18275, A2 => n1194, Z => n25889);
   U17142 : XNOR2_X1 port map( A1 => n18114, A2 => n23888, ZN => n25912);
   U17147 : INV_X4 port map( I => n6293, ZN => n9459);
   U17149 : XOR2_X1 port map( A1 => n5597, A2 => n12205, Z => n26180);
   U17153 : NAND2_X2 port map( A1 => n22206, A2 => n10125, ZN => n12205);
   U17154 : XOR2_X1 port map( A1 => n16889, A2 => n16890, Z => n11656);
   U17159 : XOR2_X1 port map( A1 => n7917, A2 => n12709, Z => n16890);
   U17163 : NAND2_X1 port map( A1 => n3013, A2 => n26048, ZN => n3012);
   U17177 : OAI21_X2 port map( A1 => n3272, A2 => n680, B => n11746, ZN => n103
                           );
   U17186 : XOR2_X1 port map( A1 => n18097, A2 => n25333, Z => n9228);
   U17187 : XOR2_X1 port map( A1 => n4055, A2 => n4053, Z => n4826);
   U17192 : OAI22_X2 port map( A1 => n24579, A2 => n22140, B1 => n3226, B2 => 
                           n9401, ZN => n19709);
   U17193 : NAND3_X1 port map( A1 => n13674, A2 => n17204, A3 => n17415, ZN => 
                           n25896);
   U17195 : NAND2_X2 port map( A1 => n9469, A2 => n9468, ZN => n25903);
   U17197 : OAI21_X2 port map( A1 => n15269, A2 => n16085, B => n9203, ZN => 
                           n9773);
   U17208 : NOR2_X2 port map( A1 => n22936, A2 => n22935, ZN => n25898);
   U17214 : XOR2_X1 port map( A1 => n17142, A2 => n9614, Z => n26274);
   U17216 : XOR2_X1 port map( A1 => n25900, A2 => n11427, Z => n2458);
   U17224 : OAI22_X2 port map( A1 => n6022, A2 => n13509, B1 => n892, B2 => 
                           n26255, ZN => n9174);
   U17227 : INV_X4 port map( I => n25904, ZN => n11112);
   U17234 : XOR2_X1 port map( A1 => n27391, A2 => n14505, Z => n10798);
   U17251 : OR2_X2 port map( A1 => n22905, A2 => n14287, Z => n10708);
   U17252 : XOR2_X1 port map( A1 => n8039, A2 => n25906, Z => n17850);
   U17253 : XOR2_X1 port map( A1 => n13000, A2 => n8037, Z => n25906);
   U17269 : XOR2_X1 port map( A1 => n4126, A2 => n7659, Z => n15661);
   U17278 : AOI22_X2 port map( A1 => n6600, A2 => n6599, B1 => n24572, B2 => 
                           n4125, ZN => n4126);
   U17279 : NOR2_X2 port map( A1 => n7535, A2 => n5796, ZN => n6588);
   U17280 : NAND2_X2 port map( A1 => n26299, A2 => n13838, ZN => n9759);
   U17302 : NAND2_X1 port map( A1 => n16130, A2 => n15828, ZN => n15776);
   U17310 : NAND2_X2 port map( A1 => n25911, A2 => n15842, ZN => n16468);
   U17320 : XOR2_X1 port map( A1 => n8848, A2 => n12405, Z => n4106);
   U17321 : XOR2_X1 port map( A1 => n4107, A2 => n14077, Z => n8848);
   U17323 : INV_X1 port map( I => n1172, ZN => n7841);
   U17329 : XOR2_X1 port map( A1 => n7843, A2 => n25912, Z => n1172);
   U17336 : NAND2_X1 port map( A1 => n27402, A2 => n19645, ZN => n26535);
   U17337 : AOI22_X2 port map( A1 => n15821, A2 => n15820, B1 => n3780, B2 => 
                           n9443, ZN => n9790);
   U17349 : NAND2_X1 port map( A1 => n14907, A2 => n14911, ZN => n26299);
   U17350 : INV_X4 port map( I => n24638, ZN => n4537);
   U17358 : AOI21_X1 port map( A1 => n24572, A2 => n25914, B => n10083, ZN => 
                           n2298);
   U17370 : NAND2_X2 port map( A1 => n22893, A2 => n1717, ZN => n6110);
   U17375 : NOR2_X1 port map( A1 => n15268, A2 => n11175, ZN => n7167);
   U17399 : XOR2_X1 port map( A1 => n27863, A2 => n21650, Z => n21854);
   U17404 : OR2_X1 port map( A1 => n17362, A2 => n25922, Z => n10620);
   U17406 : NAND2_X2 port map( A1 => n6612, A2 => n24236, ZN => n3017);
   U17411 : INV_X2 port map( I => n25923, ZN => n4667);
   U17412 : XOR2_X1 port map( A1 => n3970, A2 => n3968, Z => n25923);
   U17416 : XOR2_X1 port map( A1 => n2064, A2 => n21429, Z => n25925);
   U17419 : AOI22_X2 port map( A1 => n11952, A2 => n16687, B1 => n3948, B2 => 
                           n16423, ZN => n11951);
   U17427 : NAND2_X2 port map( A1 => n16642, A2 => n16643, ZN => n17028);
   U17430 : NOR2_X2 port map( A1 => n17809, A2 => n14180, ZN => n25930);
   U17439 : NAND2_X2 port map( A1 => n27658, A2 => n11391, ZN => n17809);
   U17447 : AND2_X1 port map( A1 => n3874, A2 => n15610, Z => n3853);
   U17451 : OR2_X1 port map( A1 => n4883, A2 => n4198, Z => n7938);
   U17475 : BUF_X2 port map( I => n16836, Z => n25933);
   U17506 : AND2_X1 port map( A1 => n8723, A2 => n25934, Z => n13454);
   U17509 : NAND2_X1 port map( A1 => n28537, A2 => n17388, ZN => n10821);
   U17510 : XOR2_X1 port map( A1 => n17075, A2 => n17076, Z => n17388);
   U17517 : NAND2_X2 port map( A1 => n24104, A2 => n24105, ZN => n6999);
   U17520 : NAND2_X2 port map( A1 => n13502, A2 => n4199, ZN => n26152);
   U17524 : NAND2_X2 port map( A1 => n5827, A2 => n23363, ZN => n4199);
   U17527 : NOR2_X1 port map( A1 => n13854, A2 => n19866, ZN => n19577);
   U17533 : INV_X2 port map( I => n13363, ZN => n13854);
   U17560 : XOR2_X1 port map( A1 => n16863, A2 => n337, Z => n6707);
   U17565 : NAND2_X2 port map( A1 => n25939, A2 => n25938, ZN => n337);
   U17573 : OAI21_X2 port map( A1 => n15189, A2 => n17490, B => n17489, ZN => 
                           n7151);
   U17578 : NAND2_X2 port map( A1 => n25942, A2 => n6235, ZN => n2788);
   U17596 : NAND2_X2 port map( A1 => n8731, A2 => n13090, ZN => n20379);
   U17609 : XOR2_X1 port map( A1 => n25356, A2 => n25944, Z => n25943);
   U17618 : INV_X1 port map( I => n14360, ZN => n25944);
   U17620 : XOR2_X1 port map( A1 => n25945, A2 => n1310, Z => Ciphertext(103));
   U17621 : NAND3_X1 port map( A1 => n21129, A2 => n23786, A3 => n13448, ZN => 
                           n25947);
   U17625 : XOR2_X1 port map( A1 => n20535, A2 => n14421, Z => n26389);
   U17626 : NAND2_X2 port map( A1 => n9342, A2 => n9340, ZN => n14421);
   U17629 : INV_X1 port map( I => n21080, ZN => n25949);
   U17631 : XOR2_X1 port map( A1 => n15819, A2 => Key(73), Z => n16007);
   U17636 : NOR2_X1 port map( A1 => n11891, A2 => n15375, ZN => n3518);
   U17639 : NAND2_X2 port map( A1 => n749, A2 => n21279, ZN => n11891);
   U17642 : XOR2_X1 port map( A1 => n5858, A2 => n2702, Z => n25950);
   U17644 : OAI21_X2 port map( A1 => n1442, A2 => n1446, B => n1441, ZN => 
                           n22760);
   U17662 : OAI21_X1 port map( A1 => n21666, A2 => n5675, B => n23999, ZN => 
                           n201);
   U17702 : NOR2_X1 port map( A1 => n6976, A2 => n25308, ZN => n9629);
   U17704 : NAND2_X1 port map( A1 => n22738, A2 => n20964, ZN => n25961);
   U17706 : XOR2_X1 port map( A1 => n3569, A2 => n3566, Z => n5535);
   U17725 : NAND3_X2 port map( A1 => n5203, A2 => n13301, A3 => n5202, ZN => 
                           n25965);
   U17730 : XOR2_X1 port map( A1 => n16754, A2 => n4030, Z => n4029);
   U17742 : OAI21_X2 port map( A1 => n24607, A2 => n11716, B => n17370, ZN => 
                           n26476);
   U17753 : XOR2_X1 port map( A1 => n9982, A2 => n24595, Z => n26606);
   U17757 : INV_X2 port map( I => n25968, ZN => n8113);
   U17758 : XOR2_X1 port map( A1 => n8114, A2 => n18289, Z => n25968);
   U17766 : INV_X1 port map( I => n11200, ZN => n26079);
   U17769 : XOR2_X1 port map( A1 => n13293, A2 => n24618, Z => n25969);
   U17784 : INV_X2 port map( I => n25970, ZN => n17244);
   U17791 : OAI22_X2 port map( A1 => n8134, A2 => n9268, B1 => n3619, B2 => 
                           n8226, ZN => n8122);
   U17797 : OR2_X1 port map( A1 => n13741, A2 => n21408, Z => n5005);
   U17798 : XOR2_X1 port map( A1 => n14753, A2 => n16755, Z => n4067);
   U17804 : XOR2_X1 port map( A1 => n22010, A2 => n9723, Z => n10332);
   U17810 : XOR2_X1 port map( A1 => n26246, A2 => n25980, Z => n548);
   U17825 : NAND2_X2 port map( A1 => n15870, A2 => n15871, ZN => n479);
   U17827 : NOR2_X1 port map( A1 => n705, A2 => n21880, ZN => n20950);
   U17828 : NAND3_X2 port map( A1 => n25986, A2 => n5981, A3 => n10271, ZN => 
                           n19562);
   U17835 : NAND2_X1 port map( A1 => n14461, A2 => n18416, ZN => n25986);
   U17845 : XOR2_X1 port map( A1 => n15256, A2 => n24107, Z => n5212);
   U17854 : INV_X2 port map( I => n25988, ZN => n24523);
   U17865 : NAND2_X2 port map( A1 => n2981, A2 => n6242, ZN => n2462);
   U17873 : NAND2_X2 port map( A1 => n9374, A2 => n7213, ZN => n2981);
   U17874 : XOR2_X1 port map( A1 => n8652, A2 => n25991, Z => n12695);
   U17878 : XOR2_X1 port map( A1 => n10208, A2 => n19390, Z => n25991);
   U17884 : NAND2_X2 port map( A1 => n17854, A2 => n15311, ZN => n18225);
   U17886 : INV_X1 port map( I => n16685, ZN => n25994);
   U17890 : XOR2_X1 port map( A1 => n11656, A2 => n25998, Z => n24416);
   U17891 : XOR2_X1 port map( A1 => n2029, A2 => n21907, Z => n18498);
   U17917 : INV_X2 port map( I => n9550, ZN => n26001);
   U17920 : XOR2_X1 port map( A1 => n5089, A2 => n18242, Z => n22637);
   U17921 : XOR2_X1 port map( A1 => n5921, A2 => n18123, Z => n18242);
   U17941 : OAI21_X2 port map( A1 => n26062, A2 => n26063, B => n17158, ZN => 
                           n7553);
   U17945 : AOI22_X2 port map( A1 => n15866, A2 => n12010, B1 => n15865, B2 => 
                           n9443, ZN => n26388);
   U17947 : XOR2_X1 port map( A1 => n1096, A2 => n8582, Z => n8581);
   U17954 : NAND2_X2 port map( A1 => n2035, A2 => n26005, ZN => n20153);
   U17973 : AOI22_X2 port map( A1 => n23514, A2 => n5483, B1 => n23499, B2 => 
                           n15463, ZN => n13267);
   U17976 : NOR2_X1 port map( A1 => n25307, A2 => n7039, ZN => n6833);
   U17979 : OAI22_X2 port map( A1 => n16276, A2 => n16277, B1 => n7868, B2 => 
                           n13562, ZN => n11614);
   U17982 : NOR2_X2 port map( A1 => n7868, A2 => n22319, ZN => n16276);
   U17986 : NAND2_X2 port map( A1 => n13758, A2 => n14177, ZN => n16370);
   U17999 : NOR2_X1 port map( A1 => n8541, A2 => n8542, ZN => n26015);
   U18041 : NOR2_X2 port map( A1 => n7298, A2 => n12600, ZN => n12599);
   U18045 : NAND2_X2 port map( A1 => n26027, A2 => n26028, ZN => n10681);
   U18062 : NAND2_X2 port map( A1 => n2728, A2 => n5120, ZN => n6600);
   U18063 : AOI21_X2 port map( A1 => n6937, A2 => n16676, B => n26024, ZN => 
                           n4002);
   U18067 : XOR2_X1 port map( A1 => n4876, A2 => n4877, Z => n9900);
   U18068 : AOI21_X2 port map( A1 => n4871, A2 => n7805, B => n4870, ZN => 
                           n4876);
   U18078 : OAI22_X2 port map( A1 => n13389, A2 => n17986, B1 => n7023, B2 => 
                           n23002, ZN => n17649);
   U18089 : OAI21_X2 port map( A1 => n14069, A2 => n25940, B => n26032, ZN => 
                           n5997);
   U18091 : XOR2_X1 port map( A1 => n19441, A2 => n19440, Z => n11709);
   U18092 : OAI22_X2 port map( A1 => n11241, A2 => n783, B1 => n11240, B2 => 
                           n1189, ZN => n15677);
   U18097 : XNOR2_X1 port map( A1 => n3834, A2 => n13746, ZN => n26168);
   U18105 : OAI21_X1 port map( A1 => n16336, A2 => n6110, B => n25415, ZN => 
                           n7092);
   U18111 : INV_X2 port map( I => n26034, ZN => n21873);
   U18113 : XOR2_X1 port map( A1 => n9861, A2 => Plaintext(0), Z => n26034);
   U18120 : OR2_X1 port map( A1 => n15890, A2 => n16350, Z => n26074);
   U18130 : NAND2_X1 port map( A1 => n22799, A2 => n26036, ZN => n26035);
   U18136 : INV_X2 port map( I => n10702, ZN => n26036);
   U18138 : XOR2_X1 port map( A1 => n8705, A2 => n7303, Z => n9143);
   U18169 : INV_X2 port map( I => n8605, ZN => n26038);
   U18180 : AND2_X1 port map( A1 => n25843, A2 => n20174, Z => n26439);
   U18182 : NAND3_X2 port map( A1 => n945, A2 => n21720, A3 => n21719, ZN => 
                           n26091);
   U18193 : OAI21_X2 port map( A1 => n9675, A2 => n27101, B => n26042, ZN => 
                           n15663);
   U18194 : XOR2_X1 port map( A1 => n19322, A2 => n10944, Z => n10945);
   U18210 : NAND3_X2 port map( A1 => n9560, A2 => n677, A3 => n7359, ZN => 
                           n14653);
   U18226 : XOR2_X1 port map( A1 => n12230, A2 => n26046, Z => n638);
   U18232 : INV_X1 port map( I => n14597, ZN => n26046);
   U18236 : NAND2_X2 port map( A1 => n14932, A2 => n14933, ZN => n12230);
   U18241 : XNOR2_X1 port map( A1 => n25337, A2 => n10294, ZN => n26480);
   U18243 : NAND2_X2 port map( A1 => n13147, A2 => n20087, ZN => n20049);
   U18245 : OR2_X1 port map( A1 => n6217, A2 => n3014, Z => n26048);
   U18248 : NOR2_X1 port map( A1 => n1014, A2 => n26317, ZN => n22326);
   U18257 : XOR2_X1 port map( A1 => n10055, A2 => n10052, Z => n10097);
   U18258 : INV_X2 port map( I => n26049, ZN => n10875);
   U18265 : OAI22_X2 port map( A1 => n6684, A2 => n2857, B1 => n6685, B2 => 
                           n10304, ZN => n26050);
   U18267 : OAI21_X2 port map( A1 => n26489, A2 => n1750, B => n25772, ZN => 
                           n1749);
   U18270 : NAND2_X1 port map( A1 => n12113, A2 => n14037, ZN => n12112);
   U18281 : XOR2_X1 port map( A1 => n12909, A2 => n25353, Z => n3753);
   U18284 : XOR2_X1 port map( A1 => n2507, A2 => n2389, Z => n2505);
   U18287 : XOR2_X1 port map( A1 => n16836, A2 => n26053, Z => n17115);
   U18288 : INV_X2 port map( I => n10123, ZN => n26053);
   U18292 : NOR2_X2 port map( A1 => n16470, A2 => n3133, ZN => n10123);
   U18297 : XOR2_X1 port map( A1 => Plaintext(158), A2 => Key(158), Z => n26106
                           );
   U18301 : NAND2_X2 port map( A1 => n23884, A2 => n10008, ZN => n2398);
   U18307 : OR2_X1 port map( A1 => n5299, A2 => n22790, Z => n26054);
   U18314 : XOR2_X1 port map( A1 => n19507, A2 => n27422, Z => n26056);
   U18320 : NAND2_X2 port map( A1 => n14687, A2 => n14688, ZN => n17847);
   U18321 : XOR2_X1 port map( A1 => n22806, A2 => n9161, Z => n12604);
   U18334 : NOR2_X2 port map( A1 => n3694, A2 => n6413, ZN => n26058);
   U18337 : NAND2_X2 port map( A1 => n19892, A2 => n19834, ZN => n14734);
   U18338 : NOR2_X1 port map( A1 => n20161, A2 => n9440, ZN => n8057);
   U18339 : NAND2_X2 port map( A1 => n26060, A2 => n23395, ZN => n12477);
   U18348 : NOR2_X2 port map( A1 => n22560, A2 => n8180, ZN => n26063);
   U18373 : XOR2_X1 port map( A1 => n26067, A2 => n58, Z => n8985);
   U18382 : NAND2_X2 port map( A1 => n3278, A2 => n23379, ZN => n26084);
   U18383 : NAND2_X1 port map( A1 => n4762, A2 => n25373, ZN => n4752);
   U18384 : XOR2_X1 port map( A1 => Plaintext(130), A2 => Key(130), Z => n4522)
                           ;
   U18386 : XOR2_X1 port map( A1 => Plaintext(80), A2 => Key(80), Z => n26068);
   U18398 : XOR2_X1 port map( A1 => n26071, A2 => n12709, Z => n2363);
   U18404 : XOR2_X1 port map( A1 => n10004, A2 => n23312, Z => n19882);
   U18405 : NAND2_X2 port map( A1 => n26075, A2 => n26074, ZN => n16691);
   U18442 : XOR2_X1 port map( A1 => n14285, A2 => n10678, Z => n11816);
   U18446 : XOR2_X1 port map( A1 => n10333, A2 => n26386, Z => n17157);
   U18451 : NAND2_X2 port map( A1 => n26079, A2 => n26078, ZN => n6181);
   U18453 : INV_X2 port map( I => n26080, ZN => n10629);
   U18455 : XNOR2_X1 port map( A1 => Plaintext(140), A2 => Key(140), ZN => 
                           n26080);
   U18468 : OAI21_X2 port map( A1 => n26102, A2 => n1175, B => n23960, ZN => 
                           n12571);
   U18490 : INV_X1 port map( I => n3943, ZN => n26087);
   U18492 : NAND2_X1 port map( A1 => n12913, A2 => n12611, ZN => n26088);
   U18495 : XOR2_X1 port map( A1 => n4067, A2 => n26093, Z => n4095);
   U18501 : NAND2_X2 port map( A1 => n5667, A2 => n781, ZN => n19206);
   U18515 : AOI21_X2 port map( A1 => n26423, A2 => n18467, B => n26159, ZN => 
                           n3329);
   U18528 : XOR2_X1 port map( A1 => n2266, A2 => n10279, Z => n12620);
   U18537 : NOR2_X2 port map( A1 => n24304, A2 => n5305, ZN => n17586);
   U18538 : OAI21_X2 port map( A1 => n51, A2 => n25222, B => n12025, ZN => 
                           n11927);
   U18544 : NAND2_X2 port map( A1 => n13613, A2 => n8173, ZN => n12025);
   U18549 : AOI22_X2 port map( A1 => n17938, A2 => n17937, B1 => n17939, B2 => 
                           n17940, ZN => n9748);
   U18578 : NAND2_X2 port map( A1 => n12272, A2 => n15989, ZN => n26104);
   U18584 : BUF_X2 port map( I => n12292, Z => n26105);
   U18585 : XNOR2_X1 port map( A1 => n9534, A2 => n16755, ZN => n17126);
   U18601 : OAI22_X2 port map( A1 => n15439, A2 => n14778, B1 => n15438, B2 => 
                           n15436, ZN => n16755);
   U18603 : INV_X2 port map( I => n26106, ZN => n22991);
   U18605 : XOR2_X1 port map( A1 => n20512, A2 => n20522, Z => n4631);
   U18618 : XOR2_X1 port map( A1 => n18214, A2 => n4901, Z => n18216);
   U18619 : AND2_X1 port map( A1 => n10875, A2 => n17250, Z => n26153);
   U18620 : NAND3_X1 port map( A1 => n7698, A2 => n20685, A3 => n25324, ZN => 
                           n20682);
   U18623 : NAND2_X1 port map( A1 => n13546, A2 => n14894, ZN => n26109);
   U18635 : NAND2_X2 port map( A1 => n26111, A2 => n26112, ZN => n12942);
   U18641 : NAND2_X2 port map( A1 => n22043, A2 => n8234, ZN => n12181);
   U18644 : NAND2_X2 port map( A1 => n26116, A2 => n26115, ZN => n13039);
   U18647 : NAND2_X1 port map( A1 => n26117, A2 => n2765, ZN => n24414);
   U18652 : INV_X1 port map( I => n13305, ZN => n26117);
   U18658 : XOR2_X1 port map( A1 => n7264, A2 => n1710, Z => n2671);
   U18661 : XOR2_X1 port map( A1 => n26118, A2 => n7375, Z => n315);
   U18671 : XOR2_X1 port map( A1 => n20498, A2 => n23898, Z => n26119);
   U18675 : XOR2_X1 port map( A1 => n6631, A2 => n6633, Z => n18549);
   U18700 : AOI21_X2 port map( A1 => n8453, A2 => n27494, B => n8452, ZN => 
                           n24445);
   U18717 : NOR2_X1 port map( A1 => n21079, A2 => n21072, ZN => n21074);
   U18719 : XOR2_X1 port map( A1 => n9357, A2 => n18218, Z => n7885);
   U18729 : AND2_X1 port map( A1 => n10830, A2 => n15834, Z => n23457);
   U18738 : NAND2_X2 port map( A1 => n20173, A2 => n24554, ZN => n26438);
   U18749 : NAND3_X1 port map( A1 => n26124, A2 => n3017, A3 => n24215, ZN => 
                           n26123);
   U18750 : OR2_X1 port map( A1 => n17724, A2 => n26144, Z => n17591);
   U18763 : NAND2_X2 port map( A1 => n26128, A2 => n26448, ZN => n4531);
   U18769 : OAI21_X1 port map( A1 => n6488, A2 => n19028, B => n19154, ZN => 
                           n8043);
   U18770 : NOR2_X2 port map( A1 => n9065, A2 => n3325, ZN => n9063);
   U18772 : AOI21_X2 port map( A1 => n18952, A2 => n9642, B => n28147, ZN => 
                           n9065);
   U18773 : NOR3_X2 port map( A1 => n16106, A2 => n22801, A3 => n8867, ZN => 
                           n26488);
   U18781 : XOR2_X1 port map( A1 => n6891, A2 => n27745, Z => n17105);
   U18806 : XOR2_X1 port map( A1 => n16909, A2 => n8115, Z => n7859);
   U18811 : NAND3_X2 port map( A1 => n7818, A2 => n16110, A3 => n7227, ZN => 
                           n10282);
   U18826 : OAI21_X2 port map( A1 => n26133, A2 => n4450, B => n8433, ZN => 
                           n2869);
   U18828 : XOR2_X1 port map( A1 => n21300, A2 => n26135, Z => n6698);
   U18829 : XOR2_X1 port map( A1 => n4259, A2 => n4258, Z => n26135);
   U18833 : INV_X2 port map( I => n17142, ZN => n1041);
   U18834 : OAI21_X2 port map( A1 => n6934, A2 => n6933, B => n24604, ZN => 
                           n17142);
   U18840 : NAND2_X2 port map( A1 => n26136, A2 => n6284, ZN => n9055);
   U18854 : NOR2_X2 port map( A1 => n8473, A2 => n748, ZN => n13282);
   U18862 : XOR2_X1 port map( A1 => n19496, A2 => n23917, Z => n19389);
   U18886 : XOR2_X1 port map( A1 => n17150, A2 => n26143, Z => n575);
   U18887 : OR2_X1 port map( A1 => n18497, A2 => n22977, Z => n14204);
   U18888 : AND2_X1 port map( A1 => n631, A2 => n26081, Z => n15322);
   U18895 : INV_X4 port map( I => n26144, ZN => n3929);
   U18896 : XOR2_X1 port map( A1 => n23703, A2 => n6379, Z => n15698);
   U18900 : NAND2_X1 port map( A1 => n846, A2 => n22803, ZN => n4726);
   U18907 : NAND2_X1 port map( A1 => n5458, A2 => n447, ZN => n22279);
   U18913 : AOI21_X2 port map( A1 => n26381, A2 => n5274, B => n24431, ZN => 
                           n24430);
   U18930 : BUF_X2 port map( I => n15930, Z => n26147);
   U18938 : XOR2_X1 port map( A1 => n26149, A2 => n20919, Z => Ciphertext(59));
   U18943 : OAI22_X1 port map( A1 => n20918, A2 => n22729, B1 => n20916, B2 => 
                           n2587, ZN => n26149);
   U18956 : XOR2_X1 port map( A1 => n19507, A2 => n19487, Z => n19501);
   U18968 : OAI21_X2 port map( A1 => n7963, A2 => n22061, B => n26150, ZN => 
                           n7200);
   U18975 : OAI21_X2 port map( A1 => n24141, A2 => n16696, B => n22061, ZN => 
                           n26150);
   U18989 : BUF_X2 port map( I => n10613, Z => n26155);
   U18990 : AOI22_X2 port map( A1 => n26651, A2 => n21544, B1 => n15697, B2 => 
                           n6547, ZN => n21512);
   U18992 : XOR2_X1 port map( A1 => n11671, A2 => n8378, Z => n9456);
   U19003 : XOR2_X1 port map( A1 => n7948, A2 => n24652, Z => n8077);
   U19007 : OR2_X1 port map( A1 => n3062, A2 => n22856, Z => n26160);
   U19021 : XOR2_X1 port map( A1 => n18217, A2 => n24357, Z => n7884);
   U19025 : OAI21_X2 port map( A1 => n4581, A2 => n21021, B => n1090, ZN => 
                           n3045);
   U19032 : XOR2_X1 port map( A1 => n9339, A2 => n19515, Z => n15161);
   U19040 : OR2_X1 port map( A1 => n6281, A2 => n6339, Z => n21740);
   U19052 : NOR3_X2 port map( A1 => n8896, A2 => n24278, A3 => n10598, ZN => 
                           n6281);
   U19056 : OR2_X1 port map( A1 => n19244, A2 => n9762, Z => n19246);
   U19078 : NAND2_X1 port map( A1 => n26166, A2 => n17502, ZN => n26165);
   U19079 : NAND3_X2 port map( A1 => n1085, A2 => n20986, A3 => n7535, ZN => 
                           n20987);
   U19080 : INV_X4 port map( I => n5324, ZN => n3948);
   U19082 : NAND2_X2 port map( A1 => n21964, A2 => n15877, ZN => n5324);
   U19090 : XOR2_X1 port map( A1 => n13747, A2 => n26168, Z => n23347);
   U19123 : XOR2_X1 port map( A1 => n19234, A2 => n4076, Z => n6912);
   U19138 : XOR2_X1 port map( A1 => n26172, A2 => n26173, Z => n5929);
   U19139 : XOR2_X1 port map( A1 => n26545, A2 => n21367, Z => n26173);
   U19154 : AOI22_X2 port map( A1 => n4101, A2 => n1203, B1 => n2736, B2 => 
                           n6076, ZN => n5920);
   U19159 : NAND2_X1 port map( A1 => n14320, A2 => n13721, ZN => n16498);
   U19167 : NAND2_X2 port map( A1 => n8239, A2 => n3440, ZN => n14320);
   U19173 : INV_X2 port map( I => n26176, ZN => n7817);
   U19181 : XOR2_X1 port map( A1 => n4618, A2 => n3701, Z => n6946);
   U19182 : XOR2_X1 port map( A1 => n26177, A2 => n19564, Z => n4658);
   U19196 : NOR2_X2 port map( A1 => n18824, A2 => n18823, ZN => n26178);
   U19204 : NAND2_X2 port map( A1 => n26179, A2 => n6362, ZN => n5368);
   U19208 : OAI21_X2 port map( A1 => n1566, A2 => n6183, B => n894, ZN => 
                           n26179);
   U19210 : INV_X2 port map( I => n26180, ZN => n21893);
   U19216 : XOR2_X1 port map( A1 => n26181, A2 => n19547, Z => n3211);
   U19219 : XOR2_X1 port map( A1 => n19546, A2 => n27397, Z => n26181);
   U19220 : XOR2_X1 port map( A1 => n5964, A2 => n5962, Z => n9362);
   U19222 : XOR2_X1 port map( A1 => n23568, A2 => n26182, Z => n5835);
   U19224 : XOR2_X1 port map( A1 => n18086, A2 => n15057, Z => n26182);
   U19227 : XOR2_X1 port map( A1 => n27421, A2 => n1136, Z => n6200);
   U19234 : INV_X2 port map( I => n26183, ZN => n617);
   U19239 : NOR2_X1 port map( A1 => n19937, A2 => n704, ZN => n21987);
   U19244 : INV_X1 port map( I => n20379, ZN => n20453);
   U19253 : XNOR2_X1 port map( A1 => n20452, A2 => n20379, ZN => n20517);
   U19294 : BUF_X2 port map( I => n16202, Z => n26186);
   U19301 : OR2_X1 port map( A1 => n26187, A2 => n7964, Z => n12891);
   U19317 : OAI22_X2 port map( A1 => n26483, A2 => n7603, B1 => n17791, B2 => 
                           n17630, ZN => n13944);
   U19327 : NAND2_X2 port map( A1 => n2083, A2 => n2082, ZN => n2068);
   U19332 : XOR2_X1 port map( A1 => n18203, A2 => n24658, Z => n13816);
   U19336 : XOR2_X1 port map( A1 => n26193, A2 => n20375, Z => n15374);
   U19354 : XOR2_X1 port map( A1 => n20443, A2 => n10950, Z => n8319);
   U19355 : XOR2_X1 port map( A1 => n21318, A2 => n22777, Z => n20443);
   U19360 : INV_X2 port map( I => n26196, ZN => n5853);
   U19361 : XOR2_X1 port map( A1 => Plaintext(174), A2 => Key(174), Z => n26196
                           );
   U19363 : INV_X1 port map( I => n9527, ZN => n26198);
   U19364 : AOI21_X2 port map( A1 => n72, A2 => n73, B => n26201, ZN => n11593)
                           ;
   U19367 : NAND2_X2 port map( A1 => n9659, A2 => n969, ZN => n10344);
   U19373 : OAI22_X1 port map( A1 => n18757, A2 => n3502, B1 => n22856, B2 => 
                           n18424, ZN => n26202);
   U19385 : NAND2_X2 port map( A1 => n1023, A2 => n14180, ZN => n14777);
   U19388 : NOR2_X2 port map( A1 => n16015, A2 => n26205, ZN => n16639);
   U19393 : NAND2_X2 port map( A1 => n25360, A2 => n8760, ZN => n20843);
   U19397 : XOR2_X1 port map( A1 => n5435, A2 => n26210, Z => n14723);
   U19398 : XOR2_X1 port map( A1 => n11102, A2 => n12862, Z => n26210);
   U19405 : NOR2_X1 port map( A1 => n10794, A2 => n4710, ZN => n26212);
   U19406 : NAND2_X2 port map( A1 => n12773, A2 => n26214, ZN => n19134);
   U19411 : XNOR2_X1 port map( A1 => n18209, A2 => n21367, ZN => n22988);
   U19421 : OAI21_X1 port map( A1 => n1211, A2 => n4192, B => n24570, ZN => 
                           n4974);
   U19423 : XOR2_X1 port map( A1 => n19314, A2 => n3155, Z => n10255);
   U19425 : XOR2_X1 port map( A1 => n12204, A2 => n16930, Z => n16829);
   U19445 : XOR2_X1 port map( A1 => n18155, A2 => n18169, Z => n18053);
   U19497 : INV_X2 port map( I => n18366, ZN => n26277);
   U19500 : NAND2_X2 port map( A1 => n11079, A2 => n6865, ZN => n26231);
   U19507 : NAND2_X1 port map( A1 => n20203, A2 => n709, ZN => n8774);
   U19518 : OR2_X1 port map( A1 => n20064, A2 => n26461, Z => n11955);
   U19538 : NOR2_X2 port map( A1 => n12470, A2 => n26233, ZN => n19016);
   U19573 : NAND2_X1 port map( A1 => n18786, A2 => n24243, ZN => n26235);
   U19577 : AND2_X1 port map( A1 => n19048, A2 => n26237, Z => n159);
   U19583 : NAND3_X1 port map( A1 => n19046, A2 => n5877, A3 => n19045, ZN => 
                           n26237);
   U19594 : XOR2_X1 port map( A1 => n491, A2 => n22759, Z => n26238);
   U19603 : XOR2_X1 port map( A1 => n4684, A2 => n4686, Z => n12598);
   U19633 : OAI21_X2 port map( A1 => n15941, A2 => n21787, B => n7144, ZN => 
                           n16224);
   U19634 : NOR2_X1 port map( A1 => n7390, A2 => n25319, ZN => n22346);
   U19649 : NAND3_X2 port map( A1 => n11824, A2 => n17657, A3 => n14994, ZN => 
                           n15237);
   U19651 : XOR2_X1 port map( A1 => n8957, A2 => n11275, Z => n10071);
   U19689 : AOI21_X1 port map( A1 => n10461, A2 => n15055, B => n9827, ZN => 
                           n8106);
   U19697 : NOR2_X2 port map( A1 => n10790, A2 => n10791, ZN => n16704);
   U19700 : OAI22_X2 port map( A1 => n4287, A2 => n15913, B1 => n4231, B2 => 
                           n799, ZN => n10790);
   U19733 : OAI22_X2 port map( A1 => n15956, A2 => n16206, B1 => n5668, B2 => 
                           n1058, ZN => n26254);
   U19735 : NAND2_X2 port map( A1 => n12185, A2 => n12184, ZN => n2656);
   U19743 : AOI21_X2 port map( A1 => n12058, A2 => n10812, B => n26256, ZN => 
                           n11575);
   U19755 : NAND2_X2 port map( A1 => n6958, A2 => n18958, ZN => n11417);
   U19756 : NAND2_X2 port map( A1 => n26258, A2 => n22570, ZN => n7543);
   U19768 : XOR2_X1 port map( A1 => n16860, A2 => n8900, Z => n3323);
   U19785 : NOR2_X2 port map( A1 => n23616, A2 => n6643, ZN => n15443);
   U19791 : NOR2_X1 port map( A1 => n17390, A2 => n12692, ZN => n26259);
   U19792 : XOR2_X1 port map( A1 => n7744, A2 => n26261, Z => n11698);
   U19799 : XOR2_X1 port map( A1 => n18044, A2 => n23375, Z => n26261);
   U19805 : XOR2_X1 port map( A1 => n20436, A2 => n14587, Z => n20437);
   U19811 : XOR2_X1 port map( A1 => n4558, A2 => n15431, Z => n18283);
   U19838 : NAND2_X2 port map( A1 => n26262, A2 => n26187, ZN => n14866);
   U19845 : XOR2_X1 port map( A1 => n26263, A2 => n5334, Z => n14416);
   U19847 : XOR2_X1 port map( A1 => n22540, A2 => n20438, Z => n26263);
   U19854 : XOR2_X1 port map( A1 => n17051, A2 => n21940, Z => n26391);
   U19864 : NOR3_X2 port map( A1 => n26267, A2 => n12449, A3 => n26266, ZN => 
                           n17806);
   U19867 : XOR2_X1 port map( A1 => n6062, A2 => n3489, Z => n26494);
   U19872 : NAND2_X2 port map( A1 => n22701, A2 => n26268, ZN => n11100);
   U19880 : XOR2_X1 port map( A1 => n25332, A2 => n26273, Z => n10683);
   U19884 : INV_X1 port map( I => n21631, ZN => n26273);
   U19908 : NAND2_X1 port map( A1 => n9461, A2 => n9462, ZN => n20340);
   U19917 : OAI22_X1 port map( A1 => n2114, A2 => n934, B1 => n2115, B2 => 
                           n2916, ZN => n22055);
   U19921 : XOR2_X1 port map( A1 => n26274, A2 => n16783, Z => n4922);
   U19924 : NOR2_X1 port map( A1 => n21768, A2 => n25214, ZN => n17278);
   U19932 : XOR2_X1 port map( A1 => n14694, A2 => n9638, Z => n9637);
   U19950 : AOI21_X2 port map( A1 => n9040, A2 => n17895, B => n22812, ZN => 
                           n2317);
   U19959 : NOR2_X1 port map( A1 => n12241, A2 => n26276, ZN => n12239);
   U19961 : NOR2_X1 port map( A1 => n10964, A2 => n25390, ZN => n26276);
   U19964 : NAND2_X2 port map( A1 => n24847, A2 => n26277, ZN => n1387);
   U19969 : XOR2_X1 port map( A1 => n2026, A2 => n9507, Z => n26278);
   U19970 : XOR2_X1 port map( A1 => n19366, A2 => n19290, Z => n26279);
   U19984 : XOR2_X1 port map( A1 => n26286, A2 => n20396, Z => Ciphertext(82));
   U19985 : OAI21_X2 port map( A1 => n1940, A2 => n6551, B => n17227, ZN => 
                           n26288);
   U19989 : NOR2_X1 port map( A1 => n20492, A2 => n20493, ZN => n20494);
   U19994 : XOR2_X1 port map( A1 => n16957, A2 => n26289, Z => n12664);
   U20015 : NAND2_X2 port map( A1 => n21980, A2 => n26156, ZN => n23158);
   U20026 : NAND2_X2 port map( A1 => n23288, A2 => n23475, ZN => n13891);
   U20027 : NOR2_X1 port map( A1 => n15509, A2 => n23115, ZN => n13734);
   U20028 : XOR2_X1 port map( A1 => n12484, A2 => n14085, Z => n23713);
   U20029 : NOR2_X1 port map( A1 => n7119, A2 => n24178, ZN => n22008);
   U20030 : XOR2_X1 port map( A1 => n13966, A2 => n26294, Z => n19403);
   U20034 : XOR2_X1 port map( A1 => n3291, A2 => n22890, Z => n26294);
   U20040 : XOR2_X1 port map( A1 => n18244, A2 => n18270, Z => n23202);
   U20047 : AOI21_X2 port map( A1 => n26295, A2 => n14634, B => n13321, ZN => 
                           n13295);
   U20049 : INV_X4 port map( I => n19161, ZN => n22338);
   U20059 : INV_X2 port map( I => n24251, ZN => n26296);
   U20061 : AOI21_X2 port map( A1 => n20080, A2 => n6470, B => n26301, ZN => 
                           n14889);
   U20066 : NAND2_X1 port map( A1 => n9618, A2 => n9619, ZN => n5510);
   U20084 : XOR2_X1 port map( A1 => n12532, A2 => n16988, Z => n8673);
   U20086 : XNOR2_X1 port map( A1 => n7885, A2 => n7882, ZN => n26302);
   U20088 : INV_X1 port map( I => n5950, ZN => n21614);
   U20100 : AOI22_X2 port map( A1 => n3629, A2 => n25834, B1 => n16434, B2 => 
                           n16701, ZN => n1664);
   U20102 : AOI21_X2 port map( A1 => n12839, A2 => n16468, B => n3443, ZN => 
                           n16434);
   U20106 : AND2_X1 port map( A1 => n10956, A2 => n674, Z => n10864);
   U20114 : NOR2_X2 port map( A1 => n21699, A2 => n21724, ZN => n21722);
   U20122 : XOR2_X1 port map( A1 => n26305, A2 => n15719, Z => n15081);
   U20141 : XOR2_X1 port map( A1 => n19383, A2 => n24667, Z => n8628);
   U20144 : OAI21_X2 port map( A1 => n26310, A2 => n24614, B => n22510, ZN => 
                           n1425);
   U20148 : NOR2_X2 port map( A1 => n26330, A2 => n11913, ZN => n8704);
   U20149 : BUF_X2 port map( I => n22057, Z => n26311);
   U20153 : OR2_X1 port map( A1 => n413, A2 => n17694, Z => n17645);
   U20159 : INV_X4 port map( I => n26312, ZN => n21842);
   U20174 : XOR2_X1 port map( A1 => n4993, A2 => n4992, Z => n8903);
   U20184 : NOR2_X2 port map( A1 => n4475, A2 => n17676, ZN => n26316);
   U20193 : OAI21_X2 port map( A1 => n23651, A2 => n23652, B => n18744, ZN => 
                           n14037);
   U20198 : OAI22_X2 port map( A1 => n1400, A2 => n9961, B1 => n22409, B2 => 
                           n7618, ZN => n1355);
   U20218 : AOI22_X2 port map( A1 => n26319, A2 => n2168, B1 => n27558, B2 => 
                           n19003, ZN => n2164);
   U20222 : NAND2_X2 port map( A1 => n675, A2 => n20142, ZN => n12362);
   U20252 : XOR2_X1 port map( A1 => n4317, A2 => n5168, Z => n26323);
   U20254 : XOR2_X1 port map( A1 => n26324, A2 => n10383, Z => n21619);
   U20264 : XOR2_X1 port map( A1 => n2193, A2 => n13589, Z => n26324);
   U20274 : AOI22_X2 port map( A1 => n11443, A2 => n5266, B1 => n3949, B2 => 
                           n3948, ZN => n26325);
   U20277 : XOR2_X1 port map( A1 => n1355, A2 => n14544, Z => n1354);
   U20298 : OAI21_X2 port map( A1 => n28544, A2 => n8697, B => n15674, ZN => 
                           n26331);
   U20323 : INV_X1 port map( I => n15081, ZN => n26405);
   U20337 : NAND2_X2 port map( A1 => n3283, A2 => n22907, ZN => n5373);
   U20350 : NOR2_X2 port map( A1 => n11382, A2 => n18613, ZN => n8697);
   U20351 : INV_X2 port map( I => n8727, ZN => n11382);
   U20363 : XOR2_X1 port map( A1 => n26334, A2 => n9383, Z => n10057);
   U20369 : OAI21_X2 port map( A1 => n24580, A2 => n2390, B => n12026, ZN => 
                           n26338);
   U20390 : NOR2_X1 port map( A1 => n4861, A2 => n17268, ZN => n13567);
   U20403 : AOI22_X2 port map( A1 => n19003, A2 => n14502, B1 => n15622, B2 => 
                           n26631, ZN => n11154);
   U20436 : XOR2_X1 port map( A1 => n26344, A2 => n14999, Z => n14082);
   U20443 : XOR2_X1 port map( A1 => n24166, A2 => n27394, Z => n26344);
   U20444 : XOR2_X1 port map( A1 => n19498, A2 => n12354, Z => n4823);
   U20476 : NOR2_X1 port map( A1 => n9269, A2 => n1214, ZN => n26347);
   U20480 : XOR2_X1 port map( A1 => n26348, A2 => n12714, Z => n22429);
   U20516 : NOR2_X1 port map( A1 => n27881, A2 => n26624, ZN => n14241);
   U20531 : XOR2_X1 port map( A1 => n8678, A2 => n19408, Z => n8677);
   U20536 : NOR2_X2 port map( A1 => n9252, A2 => n12692, ZN => n26349);
   U20541 : OR2_X1 port map( A1 => n16731, A2 => n5502, Z => n16151);
   U20548 : NOR2_X1 port map( A1 => n17363, A2 => n6672, ZN => n26351);
   U20568 : XOR2_X1 port map( A1 => n1392, A2 => n26353, Z => n24308);
   U20570 : XOR2_X1 port map( A1 => n16753, A2 => n16464, Z => n26353);
   U20590 : NAND2_X2 port map( A1 => n5198, A2 => n8898, ZN => n11603);
   U20591 : NOR2_X2 port map( A1 => n12895, A2 => n12893, ZN => n8898);
   U20595 : OR2_X1 port map( A1 => n16468, A2 => n12839, Z => n3361);
   U20610 : NOR2_X1 port map( A1 => n14906, A2 => n10393, ZN => n16361);
   U20634 : INV_X2 port map( I => n26354, ZN => n26621);
   U20644 : AOI21_X2 port map( A1 => n23718, A2 => n16670, B => n908, ZN => 
                           n9523);
   U20652 : XOR2_X1 port map( A1 => n23764, A2 => n19448, Z => n26358);
   U20665 : NAND2_X1 port map( A1 => n15482, A2 => n15483, ZN => n10486);
   U20704 : XOR2_X1 port map( A1 => n17661, A2 => n17660, Z => n18661);
   U20732 : BUF_X2 port map( I => n20156, Z => n26365);
   U20740 : INV_X2 port map( I => n26367, ZN => n2266);
   U20746 : NAND3_X2 port map( A1 => n26368, A2 => n1562, A3 => n1563, ZN => 
                           n26367);
   U20759 : NOR2_X1 port map( A1 => n13430, A2 => n15885, ZN => n11565);
   U20777 : NOR2_X1 port map( A1 => n16021, A2 => n15982, ZN => n16145);
   U20779 : XOR2_X1 port map( A1 => n14744, A2 => n17085, Z => n2699);
   U20786 : NAND2_X2 port map( A1 => n16636, A2 => n16635, ZN => n17085);
   U20790 : NAND2_X1 port map( A1 => n23062, A2 => n18581, ZN => n3937);
   U20796 : NOR2_X2 port map( A1 => n16172, A2 => n26373, ZN => n16525);
   U20804 : XOR2_X1 port map( A1 => n2440, A2 => n2441, Z => n18579);
   U20816 : OR2_X2 port map( A1 => n7608, A2 => n10204, Z => n3651);
   U20817 : NOR2_X1 port map( A1 => n10602, A2 => n7289, ZN => n11402);
   U20824 : OR2_X1 port map( A1 => n9140, A2 => n2800, Z => n23726);
   U20826 : INV_X2 port map( I => n26374, ZN => n21798);
   U20829 : XOR2_X1 port map( A1 => n16742, A2 => n16741, Z => n26374);
   U20831 : OAI22_X2 port map( A1 => n16118, A2 => n4926, B1 => n26375, B2 => 
                           n13256, ZN => n9831);
   U20832 : INV_X2 port map( I => n16150, ZN => n26375);
   U20846 : NOR2_X2 port map( A1 => n1269, A2 => n16119, ZN => n16150);
   U20856 : NAND2_X2 port map( A1 => n8009, A2 => n21792, ZN => n17666);
   U20857 : INV_X2 port map( I => n23753, ZN => n800);
   U20892 : XOR2_X1 port map( A1 => n17709, A2 => n22392, Z => n12023);
   U20914 : XOR2_X1 port map( A1 => n9780, A2 => n22432, Z => n1618);
   U20916 : NOR2_X2 port map( A1 => n26377, A2 => n9565, ZN => n9563);
   U20927 : NOR2_X2 port map( A1 => n24619, A2 => n8247, ZN => n26377);
   U20933 : XOR2_X1 port map( A1 => n12596, A2 => n9504, Z => n12595);
   U20935 : NOR2_X2 port map( A1 => n26378, A2 => n19810, ZN => n20771);
   U20940 : OAI22_X2 port map( A1 => n15281, A2 => n733, B1 => n27984, B2 => 
                           n15280, ZN => n26378);
   U20965 : NAND2_X2 port map( A1 => n15975, A2 => n15358, ZN => n15874);
   U20966 : INV_X1 port map( I => n16678, ZN => n23880);
   U20976 : NAND2_X2 port map( A1 => n7255, A2 => n14214, ZN => n16678);
   U20985 : OAI21_X1 port map( A1 => n26380, A2 => n14148, B => n24443, ZN => 
                           n22203);
   U20998 : NOR2_X1 port map( A1 => n1067, A2 => n22848, ZN => n26380);
   U21010 : AOI21_X1 port map( A1 => n6654, A2 => n6653, B => n23556, ZN => 
                           n26384);
   U21011 : NAND2_X2 port map( A1 => n1927, A2 => n4645, ZN => n4644);
   U21020 : XOR2_X1 port map( A1 => n137, A2 => n11821, Z => n19693);
   U21034 : XOR2_X1 port map( A1 => n21309, A2 => n26389, Z => n22254);
   U21038 : NAND2_X2 port map( A1 => n13651, A2 => n13650, ZN => n2544);
   U21060 : XOR2_X1 port map( A1 => n18130, A2 => n1306, Z => n6129);
   U21064 : AOI22_X2 port map( A1 => n23386, A2 => n22628, B1 => n17852, B2 => 
                           n23064, ZN => n18130);
   U21102 : XOR2_X1 port map( A1 => n26391, A2 => n23373, Z => n23684);
   U21178 : XOR2_X1 port map( A1 => n16822, A2 => n22926, Z => n26398);
   U21179 : NAND2_X2 port map( A1 => n9851, A2 => n21057, ZN => n21086);
   U21191 : NAND2_X2 port map( A1 => n1255, A2 => n3729, ZN => n26400);
   U21204 : NAND2_X2 port map( A1 => n26401, A2 => n6895, ZN => n20138);
   U21205 : XOR2_X1 port map( A1 => n20770, A2 => n20769, Z => n24281);
   U21208 : XOR2_X1 port map( A1 => n26402, A2 => n6071, Z => n24530);
   U21211 : XOR2_X1 port map( A1 => n16754, A2 => n4173, Z => n2903);
   U21223 : XOR2_X1 port map( A1 => n7874, A2 => n15057, Z => n26406);
   U21230 : XOR2_X1 port map( A1 => n11261, A2 => n7751, Z => n3640);
   U21236 : NOR2_X2 port map( A1 => n22689, A2 => n7239, ZN => n7751);
   U21246 : OR2_X1 port map( A1 => n21086, A2 => n6485, Z => n21079);
   U21265 : NOR2_X1 port map( A1 => n21109, A2 => n21110, ZN => n21112);
   U21270 : NOR2_X1 port map( A1 => n7291, A2 => n25753, ZN => n26412);
   U21290 : XOR2_X1 port map( A1 => n26414, A2 => n641, Z => n2013);
   U21300 : NOR2_X2 port map( A1 => n24829, A2 => n25875, ZN => n16668);
   U21302 : OAI22_X2 port map( A1 => n11344, A2 => n1152, B1 => n24572, B2 => 
                           n5120, ZN => n10389);
   U21329 : NAND2_X2 port map( A1 => n10695, A2 => n22533, ZN => n21435);
   U21339 : XOR2_X1 port map( A1 => n27459, A2 => n12230, Z => n9750);
   U21362 : XOR2_X1 port map( A1 => n9745, A2 => n9746, Z => n13303);
   U21368 : XOR2_X1 port map( A1 => n19388, A2 => n3368, Z => n6753);
   U21385 : OAI21_X2 port map( A1 => n26421, A2 => n26420, B => n20225, ZN => 
                           n9115);
   U21387 : NOR2_X1 port map( A1 => n8898, A2 => n20224, ZN => n26420);
   U21411 : NAND3_X2 port map( A1 => n1334, A2 => n1330, A3 => n1328, ZN => 
                           n19507);
   U21416 : OAI21_X2 port map( A1 => n5150, A2 => n5152, B => n26425, ZN => 
                           n18110);
   U21417 : OAI21_X1 port map( A1 => n5149, A2 => n15539, B => n11497, ZN => 
                           n26425);
   U21418 : NAND2_X2 port map( A1 => n26426, A2 => n22891, ZN => n23907);
   U21438 : NAND2_X2 port map( A1 => n16058, A2 => n16106, ZN => n26426);
   U21439 : XOR2_X1 port map( A1 => n26012, A2 => n27446, Z => n6155);
   U21457 : XOR2_X1 port map( A1 => n26427, A2 => n2274, Z => n2277);
   U21459 : XOR2_X1 port map( A1 => n16767, A2 => n2276, Z => n26427);
   U21503 : XOR2_X1 port map( A1 => n18133, A2 => n24542, Z => n26429);
   U21505 : XOR2_X1 port map( A1 => n24094, A2 => n20535, Z => n20518);
   U21520 : INV_X1 port map( I => n9115, ZN => n26432);
   U21541 : OAI21_X2 port map( A1 => n24554, A2 => n26439, B => n26438, ZN => 
                           n3873);
   U21551 : XOR2_X1 port map( A1 => n26440, A2 => n10495, Z => n15564);
   U21552 : XOR2_X1 port map( A1 => n2795, A2 => n6087, Z => n26440);
   U21555 : NAND2_X2 port map( A1 => n12143, A2 => n27129, ZN => n19700);
   U21558 : OAI21_X2 port map( A1 => n10347, A2 => n3655, B => n10344, ZN => 
                           n11487);
   U21572 : NOR2_X1 port map( A1 => n1258, A2 => n11024, ZN => n11528);
   U21579 : XOR2_X1 port map( A1 => n5870, A2 => n18011, Z => n22940);
   U21584 : XOR2_X1 port map( A1 => n27470, A2 => n11707, Z => n6664);
   U21586 : NAND2_X2 port map( A1 => n26445, A2 => n19186, ZN => n20142);
   U21594 : NAND2_X2 port map( A1 => n14500, A2 => n22559, ZN => n13349);
   U21599 : NAND3_X1 port map( A1 => n12831, A2 => n2576, A3 => n2490, ZN => 
                           n2488);
   U21600 : NAND2_X2 port map( A1 => n23780, A2 => n2353, ZN => n12831);
   U21611 : NOR2_X2 port map( A1 => n334, A2 => n24383, ZN => n26451);
   U21613 : NOR2_X1 port map( A1 => n16275, A2 => n16088, ZN => n7536);
   U21614 : XOR2_X1 port map( A1 => n26479, A2 => n8422, Z => n21941);
   U21617 : XOR2_X1 port map( A1 => n9598, A2 => n20358, Z => n26453);
   U21618 : INV_X2 port map( I => n26455, ZN => n9979);
   U21622 : XOR2_X1 port map( A1 => n9980, A2 => n9983, Z => n26455);
   U21623 : XOR2_X1 port map( A1 => n5613, A2 => n4412, Z => n7918);
   U21645 : NAND2_X2 port map( A1 => n19611, A2 => n19610, ZN => n20131);
   U21651 : XOR2_X1 port map( A1 => n21198, A2 => n11815, Z => n20546);
   U21653 : NOR2_X2 port map( A1 => n9519, A2 => n9518, ZN => n21198);
   U21654 : OAI21_X1 port map( A1 => n28537, A2 => n26614, B => n17479, ZN => 
                           n4465);
   U21655 : XNOR2_X1 port map( A1 => n2188, A2 => n24477, ZN => n26614);
   U21658 : INV_X2 port map( I => n8982, ZN => n21692);
   U21664 : XOR2_X1 port map( A1 => n24096, A2 => n8984, Z => n8982);
   U21668 : NOR2_X1 port map( A1 => n18516, A2 => n12672, ZN => n21795);
   U21677 : NAND2_X1 port map( A1 => n26464, A2 => n26463, ZN => n23628);
   U21679 : NAND2_X1 port map( A1 => n15239, A2 => n11733, ZN => n26464);
   U21682 : XOR2_X1 port map( A1 => n9982, A2 => n9981, Z => n9980);
   U21684 : XOR2_X1 port map( A1 => n21311, A2 => n8629, Z => n9981);
   U21685 : XOR2_X1 port map( A1 => n14940, A2 => n8628, Z => n8627);
   U21689 : XOR2_X1 port map( A1 => n15708, A2 => n26141, Z => n13856);
   U21690 : XOR2_X1 port map( A1 => n8490, A2 => n5283, Z => n20395);
   U21706 : OAI21_X2 port map( A1 => n3082, A2 => n27447, B => n3080, ZN => 
                           n3107);
   U21711 : XOR2_X1 port map( A1 => n26471, A2 => n4747, Z => n4743);
   U21712 : XOR2_X1 port map( A1 => n16826, A2 => n28058, Z => n26471);
   U21713 : OAI21_X2 port map( A1 => n26472, A2 => n17478, B => n8986, ZN => 
                           n17061);
   U21717 : INV_X2 port map( I => n6780, ZN => n19873);
   U21725 : INV_X1 port map( I => n21712, ZN => n26473);
   U21733 : XOR2_X1 port map( A1 => n6251, A2 => n22725, Z => n3562);
   U21748 : XOR2_X1 port map( A1 => n19428, A2 => n8399, Z => n13157);
   U21751 : XOR2_X1 port map( A1 => n8424, A2 => n26480, Z => n26479);
   U21760 : NAND2_X2 port map( A1 => n26481, A2 => n4062, ZN => n16604);
   U21765 : NAND2_X1 port map( A1 => n6585, A2 => n6586, ZN => n6584);
   U21767 : XOR2_X1 port map( A1 => n17129, A2 => n12778, Z => n2962);
   U21770 : XOR2_X1 port map( A1 => n26575, A2 => n16863, Z => n17129);
   U21772 : AND2_X1 port map( A1 => n9042, A2 => n26485, Z => n23073);
   U21779 : NAND2_X2 port map( A1 => n6141, A2 => n11473, ZN => n22000);
   U21783 : XOR2_X1 port map( A1 => n13519, A2 => n26493, Z => n21774);
   U21787 : XOR2_X1 port map( A1 => n17066, A2 => n15466, Z => n26493);
   U21789 : NAND2_X2 port map( A1 => n8826, A2 => n8827, ZN => n22529);
   U21798 : NAND2_X2 port map( A1 => n22011, A2 => n3277, ZN => n3644);
   U21800 : NAND2_X1 port map( A1 => n7118, A2 => n7117, ZN => n22891);
   U21801 : XOR2_X1 port map( A1 => n7431, A2 => n26053, Z => n11337);
   U21809 : NAND2_X2 port map( A1 => n5326, A2 => n7428, ZN => n7431);
   U21810 : BUF_X2 port map( I => n1436, Z => n26496);
   U21812 : OAI22_X1 port map( A1 => n21637, A2 => n438, B1 => n13908, B2 => 
                           n932, ZN => n26497);
   U21815 : INV_X2 port map( I => n28546, ZN => n6593);
   U21821 : INV_X2 port map( I => n14041, ZN => n19003);
   U21822 : NAND2_X2 port map( A1 => n7919, A2 => n25368, ZN => n14041);
   U21823 : NAND2_X1 port map( A1 => n26498, A2 => n22256, ZN => n11601);
   U21828 : OAI21_X1 port map( A1 => n11587, A2 => n21112, B => n21111, ZN => 
                           n26498);
   U21830 : XOR2_X1 port map( A1 => n26499, A2 => n17105, Z => n9454);
   U21838 : XOR2_X1 port map( A1 => n8040, A2 => n9456, Z => n26499);
   U21843 : NOR3_X1 port map( A1 => n12784, A2 => n27431, A3 => n13987, ZN => 
                           n11765);
   U21846 : NAND3_X1 port map( A1 => n19962, A2 => n12712, A3 => n1731, ZN => 
                           n5030);
   U21847 : INV_X2 port map( I => n26501, ZN => n9584);
   U21848 : INV_X2 port map( I => n7454, ZN => n21110);
   U21849 : NAND2_X2 port map( A1 => n3788, A2 => n3789, ZN => n7454);
   U21865 : BUF_X2 port map( I => n14529, Z => n26505);
   U21874 : XOR2_X1 port map( A1 => Plaintext(173), A2 => Key(173), Z => n14748
                           );
   U21877 : XOR2_X1 port map( A1 => n1527, A2 => n23518, Z => n1565);
   U21878 : XOR2_X1 port map( A1 => n26507, A2 => n21607, Z => Ciphertext(160))
                           ;
   U21880 : NOR2_X1 port map( A1 => n16630, A2 => n21970, ZN => n4967);
   U21881 : INV_X2 port map( I => n26510, ZN => n612);
   U21894 : OAI22_X1 port map( A1 => n21579, A2 => n21624, B1 => n11286, B2 => 
                           n21627, ZN => n82);
   U21895 : NOR3_X1 port map( A1 => n16686, A2 => n8344, A3 => n5324, ZN => 
                           n24051);
   U21900 : INV_X2 port map( I => n26515, ZN => n26616);
   U21901 : XOR2_X1 port map( A1 => n1438, A2 => n8143, Z => n26515);
   U21902 : INV_X4 port map( I => n4455, ZN => n14255);
   U21903 : OAI21_X2 port map( A1 => n7785, A2 => n372, B => n13687, ZN => 
                           n4455);
   U21905 : NAND2_X2 port map( A1 => n20052, A2 => n20051, ZN => n21158);
   U21909 : XOR2_X1 port map( A1 => n4222, A2 => n22686, Z => n11809);
   U21910 : NOR2_X2 port map( A1 => n3387, A2 => n3388, ZN => n11478);
   U21911 : XOR2_X1 port map( A1 => n18438, A2 => n18437, Z => n19864);
   U21912 : NAND2_X2 port map( A1 => n20240, A2 => n20183, ZN => n1475);
   U21913 : OAI22_X2 port map( A1 => n20181, A2 => n20044, B1 => n20016, B2 => 
                           n20237, ZN => n20240);
   U21916 : NAND2_X2 port map( A1 => n5000, A2 => n4999, ZN => n7395);
   U21919 : XOR2_X1 port map( A1 => n12925, A2 => n21144, Z => n15710);
   U21920 : OAI21_X2 port map( A1 => n23055, A2 => n18369, B => n26520, ZN => 
                           n2582);
   U21922 : NAND3_X1 port map( A1 => n2842, A2 => n2844, A3 => n846, ZN => 
                           n2841);
   U21925 : NOR2_X2 port map( A1 => n3046, A2 => n13352, ZN => n3042);
   U21928 : BUF_X2 port map( I => n7464, Z => n26522);
   U21929 : AOI21_X1 port map( A1 => n26523, A2 => n9848, B => n9847, ZN => 
                           n9846);
   U21930 : OAI21_X1 port map( A1 => n9850, A2 => n15658, B => n932, ZN => 
                           n26523);
   U21932 : OAI21_X2 port map( A1 => n2471, A2 => n20240, B => n2470, ZN => 
                           n21302);
   U21935 : INV_X2 port map( I => n26531, ZN => n24517);
   U21936 : XOR2_X1 port map( A1 => n7859, A2 => n7856, Z => n26531);
   U21938 : OAI21_X2 port map( A1 => n13075, A2 => n19957, B => n13074, ZN => 
                           n20344);
   U21940 : XOR2_X1 port map( A1 => n7644, A2 => n26536, Z => n23203);
   U21941 : NAND2_X2 port map( A1 => n9079, A2 => n9077, ZN => n9076);
   U21942 : NAND2_X1 port map( A1 => n26540, A2 => n26538, ZN => n17699);
   U21943 : INV_X1 port map( I => n26539, ZN => n26538);
   U21945 : NAND2_X1 port map( A1 => n17695, A2 => n728, ZN => n26540);
   U21947 : XOR2_X1 port map( A1 => n16778, A2 => n10535, Z => n17132);
   U21948 : AND2_X1 port map( A1 => n26541, A2 => n1974, Z => n6073);
   U21949 : NAND2_X2 port map( A1 => n12295, A2 => n26542, ZN => n13987);
   U21950 : OR2_X1 port map( A1 => n12294, A2 => n1703, Z => n26542);
   U21953 : NOR2_X2 port map( A1 => n9522, A2 => n9523, ZN => n17013);
   U21954 : NOR2_X1 port map( A1 => n9569, A2 => n26989, ZN => n2139);
   U21955 : NAND2_X2 port map( A1 => n11420, A2 => n26543, ZN => n3803);
   U21956 : XOR2_X1 port map( A1 => n20539, A2 => n22108, Z => n3806);
   U21957 : XOR2_X1 port map( A1 => n21254, A2 => n22099, Z => n20539);
   U21958 : NAND2_X2 port map( A1 => n2247, A2 => n2245, ZN => n26570);
   U21959 : XOR2_X1 port map( A1 => n20283, A2 => n21154, Z => n20284);
   U21960 : XOR2_X1 port map( A1 => n27371, A2 => n20773, Z => n21154);
   U21962 : BUF_X2 port map( I => n985, Z => n26545);
   U21963 : INV_X1 port map( I => n19064, ZN => n26547);
   U21965 : XOR2_X1 port map( A1 => n18228, A2 => n22802, Z => n26548);
   U21966 : XOR2_X1 port map( A1 => n26549, A2 => n14491, Z => Ciphertext(123))
                           ;
   U21968 : OAI21_X1 port map( A1 => n21275, A2 => n4143, B => n21389, ZN => 
                           n26552);
   U21969 : NOR2_X2 port map( A1 => n26555, A2 => n19855, ZN => n20404);
   U21973 : XOR2_X1 port map( A1 => n19351, A2 => n23539, Z => n26559);
   U21976 : INV_X2 port map( I => n26561, ZN => n4410);
   U21977 : XOR2_X1 port map( A1 => n10077, A2 => n4411, Z => n26561);
   U21978 : INV_X2 port map( I => n26562, ZN => n5139);
   U21979 : XNOR2_X1 port map( A1 => Plaintext(180), A2 => Key(180), ZN => 
                           n26562);
   U21982 : INV_X2 port map( I => n24083, ZN => n20132);
   U21984 : NAND2_X1 port map( A1 => n20564, A2 => n26566, ZN => n4908);
   U21987 : NAND2_X2 port map( A1 => n19073, A2 => n22643, ZN => n7840);
   U21992 : XOR2_X1 port map( A1 => n21150, A2 => n9640, Z => n26569);
   U21994 : XOR2_X1 port map( A1 => n6445, A2 => n4768, Z => n19345);
   U21998 : XOR2_X1 port map( A1 => n14047, A2 => n14048, Z => n14046);
   U22006 : NOR2_X1 port map( A1 => n14611, A2 => n20200, ZN => n26577);
   U22008 : XOR2_X1 port map( A1 => Plaintext(188), A2 => Key(188), Z => n6063)
                           ;
   U22010 : NAND3_X2 port map( A1 => n17768, A2 => n3141, A3 => n17872, ZN => 
                           n12164);
   U22013 : XOR2_X1 port map( A1 => n26579, A2 => n7187, Z => n7701);
   U22019 : XOR2_X1 port map( A1 => n26583, A2 => n23409, Z => n19280);
   U22022 : NAND2_X1 port map( A1 => n13719, A2 => n20043, ZN => n7345);
   U22023 : XOR2_X1 port map( A1 => n26584, A2 => n10053, Z => n10052);
   U22029 : XOR2_X1 port map( A1 => n26589, A2 => n8991, Z => n3600);
   U22031 : NAND2_X2 port map( A1 => n6190, A2 => n6188, ZN => n2525);
   U22032 : XOR2_X1 port map( A1 => n5537, A2 => n21143, Z => n13361);
   U22033 : NOR3_X1 port map( A1 => n3835, A2 => n19759, A3 => n7464, ZN => 
                           n6811);
   U22034 : NOR2_X2 port map( A1 => n22281, A2 => n13069, ZN => n26590);
   U22037 : NAND3_X2 port map( A1 => n24598, A2 => n2562, A3 => n18043, ZN => 
                           n18173);
   U22038 : XOR2_X1 port map( A1 => n26592, A2 => n14550, Z => Ciphertext(66));
   U22040 : NAND2_X1 port map( A1 => n722, A2 => n1699, ZN => n15562);
   U22043 : NOR2_X1 port map( A1 => n11835, A2 => n14858, ZN => n10230);
   U22045 : XOR2_X1 port map( A1 => n20513, A2 => n20515, Z => n12474);
   U22051 : NAND2_X2 port map( A1 => n26599, A2 => n5649, ZN => n23018);
   U22053 : XOR2_X1 port map( A1 => n6946, A2 => n18082, Z => n26600);
   U22056 : OR2_X1 port map( A1 => n20986, A2 => n24078, Z => n22407);
   U22057 : NAND2_X2 port map( A1 => n1839, A2 => n26603, ZN => n23744);
   U22059 : XOR2_X1 port map( A1 => n26604, A2 => n1300, Z => Ciphertext(133));
   U22060 : XOR2_X1 port map( A1 => n24536, A2 => n26606, Z => n126);
   U22061 : NOR2_X1 port map( A1 => n2447, A2 => n21342, ZN => n4829);
   U22063 : NOR2_X2 port map( A1 => n26611, A2 => n1598, ZN => n15638);
   U22066 : NAND2_X1 port map( A1 => n22365, A2 => n26638, ZN => n19587);
   U22067 : OR2_X1 port map( A1 => n16730, A2 => n16728, Z => n23162);
   U22068 : XOR2_X1 port map( A1 => n10676, A2 => n26612, Z => n12489);
   U22069 : XOR2_X1 port map( A1 => n12285, A2 => n13852, Z => n26612);
   U22070 : XOR2_X1 port map( A1 => n3529, A2 => n24500, Z => n24499);
   U22073 : XOR2_X1 port map( A1 => n19485, A2 => n19286, Z => n26613);
   U22074 : NAND3_X2 port map( A1 => n16623, A2 => n14102, A3 => n16624, ZN => 
                           n12204);
   U22075 : INV_X2 port map( I => n17548, ZN => n1224);
   U22077 : INV_X2 port map( I => n17983, ZN => n18673);
   U22078 : INV_X2 port map( I => n10499, ZN => n10601);
   U22079 : INV_X2 port map( I => n19707, ZN => n14726);
   U22081 : XOR2_X1 port map( A1 => n2522, A2 => n2618, Z => n26626);
   U22082 : INV_X2 port map( I => n14712, ZN => n22767);
   U3271 : NAND2_X2 port map( A1 => n10392, A2 => n415, ZN => n12686);
   U5714 : NOR2_X2 port map( A1 => n14128, A2 => n14649, ZN => n5230);
   U8861 : INV_X2 port map( I => n12933, ZN => n3113);
   U5992 : NOR2_X2 port map( A1 => n9446, A2 => n9264, ZN => n8236);
   U3232 : NOR2_X2 port map( A1 => n3960, A2 => n8290, ZN => n5458);
   U8167 : OAI22_X2 port map( A1 => n15761, A2 => n11693, B1 => n16219, B2 => 
                           n24132, ZN => n15507);
   U2083 : INV_X2 port map( I => n16630, ZN => n907);
   U4622 : NAND2_X2 port map( A1 => n26675, A2 => n9569, ZN => n10181);
   U2145 : OAI21_X2 port map( A1 => n13809, A2 => n15560, B => n19945, ZN => 
                           n11642);
   U2393 : INV_X2 port map( I => n8636, ZN => n9912);
   U765 : INV_X4 port map( I => n1189, ZN => n1014);
   U21697 : INV_X2 port map( I => n14364, ZN => n5502);
   U700 : INV_X2 port map( I => n18256, ZN => n23199);
   U4008 : BUF_X4 port map( I => n13757, Z => n23126);
   U5501 : BUF_X2 port map( I => n17217, Z => n26343);
   U4776 : INV_X2 port map( I => n11382, ZN => n1185);
   U1037 : INV_X4 port map( I => n8986, ZN => n1035);
   U3560 : INV_X2 port map( I => n14991, ZN => n25063);
   U8583 : BUF_X4 port map( I => n12195, Z => n11577);
   U64 : NAND2_X2 port map( A1 => n22821, A2 => n9047, ZN => n12809);
   U1467 : INV_X2 port map( I => n7431, ZN => n17114);
   U5211 : NAND2_X2 port map( A1 => n9323, A2 => n13390, ZN => n6115);
   U544 : INV_X2 port map( I => n18612, ZN => n18613);
   U1202 : NAND2_X2 port map( A1 => n16713, A2 => n12050, ZN => n9820);
   U242 : INV_X2 port map( I => n7562, ZN => n20565);
   U9557 : AOI21_X2 port map( A1 => n13160, A2 => n12870, B => n27871, ZN => 
                           n13159);
   U2351 : INV_X2 port map( I => n24646, ZN => n7487);
   U4022 : BUF_X4 port map( I => n15339, Z => n24258);
   U15054 : NOR2_X2 port map( A1 => n7449, A2 => n27341, ZN => n23987);
   U4506 : BUF_X2 port map( I => n19931, Z => n25103);
   U17767 : NOR3_X2 port map( A1 => n18628, A2 => n820, A3 => n18546, ZN => 
                           n22457);
   U13073 : AOI21_X2 port map( A1 => n17440, A2 => n17384, B => n12340, ZN => 
                           n4803);
   U3657 : NOR2_X2 port map( A1 => n19360, A2 => n8048, ZN => n19640);
   U13335 : NOR2_X2 port map( A1 => n12528, A2 => n14306, ZN => n3797);
   U1675 : NAND2_X2 port map( A1 => n24267, A2 => n24270, ZN => n15877);
   U201 : INV_X2 port map( I => n20894, ZN => n25630);
   U7339 : INV_X2 port map( I => n9674, ZN => n981);
   U3459 : NAND2_X2 port map( A1 => n16687, A2 => n479, ZN => n25731);
   U18083 : BUF_X4 port map( I => n14243, Z => n26029);
   U3092 : OR2_X2 port map( A1 => n10246, A2 => n7950, Z => n17493);
   U1578 : NOR2_X2 port map( A1 => n6763, A2 => n23107, ZN => n16418);
   U1618 : OAI21_X2 port map( A1 => n25826, A2 => n25825, B => n25657, ZN => 
                           n16046);
   U20762 : OAI21_X2 port map( A1 => n25796, A2 => n14367, B => n748, ZN => 
                           n17294);
   U22005 : NOR2_X2 port map( A1 => n4308, A2 => n21445, ZN => n5626);
   U58 : NAND2_X2 port map( A1 => n1090, A2 => n9677, ZN => n10687);
   U15350 : OR2_X2 port map( A1 => n3932, A2 => n12195, Z => n1412);
   U2162 : AND2_X2 port map( A1 => n1458, A2 => n14302, Z => n19652);
   U1031 : NOR2_X2 port map( A1 => n309, A2 => n3741, ZN => n22560);
   U3200 : BUF_X4 port map( I => n16602, Z => n132);
   U8174 : INV_X2 port map( I => n21342, ZN => n21348);
   U20717 : OAI21_X2 port map( A1 => n26147, A2 => n16138, B => n7332, ZN => 
                           n7331);
   U6208 : INV_X2 port map( I => n19651, ZN => n1133);
   U4410 : INV_X4 port map( I => n14520, ZN => n11423);
   U3944 : BUF_X2 port map( I => n19967, Z => n25294);
   U842 : NOR2_X2 port map( A1 => n1882, A2 => n829, ZN => n17813);
   U8048 : INV_X4 port map( I => n13211, ZN => n9379);
   U19771 : INV_X4 port map( I => n15443, ZN => n14026);
   U12001 : NAND2_X2 port map( A1 => n8418, A2 => n10207, ZN => n23079);
   U2546 : NAND2_X2 port map( A1 => n14059, A2 => n24862, ZN => n20166);
   U21785 : NAND2_X2 port map( A1 => n17600, A2 => n17599, ZN => n15339);
   U3611 : NAND2_X2 port map( A1 => n12571, A2 => n12781, ZN => n12980);
   U495 : AOI21_X2 port map( A1 => n11936, A2 => n26624, B => n10562, ZN => 
                           n9452);
   U1376 : INV_X2 port map( I => n17181, ZN => n23171);
   U14171 : NOR2_X2 port map( A1 => n12702, A2 => n12704, ZN => n19056);
   U252 : INV_X2 port map( I => n103, ZN => n1611);
   U19148 : OAI21_X2 port map( A1 => n13979, A2 => n21586, B => n27023, ZN => 
                           n12012);
   U8045 : AOI22_X2 port map( A1 => n16662, A2 => n9500, B1 => n16661, B2 => 
                           n16663, ZN => n4495);
   U1541 : NOR2_X2 port map( A1 => n390, A2 => n14177, ZN => n16662);
   U5150 : BUF_X2 port map( I => n172, Z => n25159);
   U4340 : INV_X2 port map( I => n16167, ZN => n719);
   U1299 : INV_X2 port map( I => n19056, ZN => n12781);
   U6215 : BUF_X2 port map( I => n10338, Z => n9768);
   U220 : NOR2_X2 port map( A1 => n22987, A2 => n21963, ZN => n25383);
   U1131 : INV_X2 port map( I => n22803, ZN => n20915);
   U12224 : INV_X4 port map( I => n20064, ZN => n1110);
   U5097 : INV_X2 port map( I => n3971, ZN => n802);
   U20481 : INV_X2 port map( I => n14306, ZN => n15887);
   U3109 : NAND2_X2 port map( A1 => n7539, A2 => n16419, ZN => n1413);
   U3237 : NAND2_X2 port map( A1 => n4070, A2 => n2897, ZN => n17864);
   U10800 : INV_X2 port map( I => n1398, ZN => n15282);
   U942 : NAND2_X2 port map( A1 => n13573, A2 => n14037, ZN => n19021);
   U2294 : NAND2_X2 port map( A1 => n3927, A2 => n28402, ZN => n4859);
   U8742 : INV_X2 port map( I => n10445, ZN => n1094);
   U1171 : OAI21_X2 port map( A1 => n13690, A2 => n793, B => n13572, ZN => 
                           n24025);
   U914 : NAND2_X2 port map( A1 => n16333, A2 => n16332, ZN => n13265);
   U4288 : INV_X4 port map( I => n4070, ZN => n713);
   U8450 : AOI21_X1 port map( A1 => n27407, A2 => n9894, B => n9893, ZN => 
                           n7384);
   U5047 : INV_X2 port map( I => n10868, ZN => n16701);
   U11445 : INV_X4 port map( I => n11114, ZN => n19748);
   U3882 : AOI21_X2 port map( A1 => n26640, A2 => n14358, B => n19091, ZN => 
                           n1959);
   U5394 : INV_X2 port map( I => n16380, ZN => n16176);
   U15068 : INV_X4 port map( I => n1458, ZN => n1459);
   U239 : INV_X4 port map( I => n10151, ZN => n20186);
   U4982 : NOR2_X2 port map( A1 => n1023, A2 => n8009, ZN => n9331);
   U13564 : NAND2_X2 port map( A1 => n13104, A2 => n25340, ZN => n20192);
   U481 : INV_X2 port map( I => n11874, ZN => n18807);
   U2973 : INV_X2 port map( I => n20194, ZN => n20147);
   U13009 : INV_X2 port map( I => n27858, ZN => n8629);
   U2686 : NAND2_X2 port map( A1 => n25542, A2 => n24570, ZN => n17998);
   U5615 : INV_X2 port map( I => n20277, ZN => n21944);
   U595 : INV_X2 port map( I => n18130, ZN => n8432);
   U3718 : INV_X2 port map( I => n19090, ZN => n11839);
   U3648 : OAI21_X2 port map( A1 => n23216, A2 => n19790, B => n23215, ZN => 
                           n19670);
   U10619 : BUF_X2 port map( I => n14542, Z => n6316);
   U5599 : NAND2_X2 port map( A1 => n18380, A2 => n878, ZN => n11184);
   U1978 : NAND2_X2 port map( A1 => n2587, A2 => n20911, ZN => n12034);
   U1300 : INV_X2 port map( I => n2068, ZN => n17791);
   U17888 : NAND2_X2 port map( A1 => n17529, A2 => n14324, ZN => n13902);
   U1471 : INV_X2 port map( I => n27661, ZN => n23502);
   U1338 : NAND2_X2 port map( A1 => n26165, A2 => n1350, ZN => n17824);
   U12738 : INV_X2 port map( I => n5130, ZN => n10930);
   U6024 : INV_X2 port map( I => n4679, ZN => n12672);
   U17816 : NOR2_X2 port map( A1 => n18424, A2 => n26121, ZN => n11058);
   U1229 : NAND2_X2 port map( A1 => n22117, A2 => n836, ZN => n15945);
   U9853 : INV_X2 port map( I => n16858, ZN => n13067);
   U13229 : INV_X2 port map( I => n18755, ZN => n10594);
   U438 : NAND2_X2 port map( A1 => n23936, A2 => n23937, ZN => n18836);
   U12601 : NAND2_X2 port map( A1 => n20336, A2 => n7057, ZN => n7704);
   U9568 : INV_X2 port map( I => n4706, ZN => n18379);
   U178 : NAND2_X2 port map( A1 => n20644, A2 => n9979, ZN => n20643);
   U15127 : INV_X4 port map( I => n9472, ZN => n12617);
   U7970 : NAND2_X2 port map( A1 => n1802, A2 => n6347, ZN => n2303);
   U417 : NAND2_X2 port map( A1 => n12143, A2 => n27010, ZN => n26456);
   U1587 : INV_X2 port map( I => n5861, ZN => n6347);
   U17263 : NOR2_X2 port map( A1 => n17447, A2 => n1036, ZN => n10634);
   U992 : AND2_X2 port map( A1 => n12699, A2 => n13303, Z => n24666);
   U13502 : NAND2_X2 port map( A1 => n10862, A2 => n4246, ZN => n23552);
   U1574 : NAND2_X2 port map( A1 => n16508, A2 => n16605, ZN => n25482);
   U17709 : INV_X2 port map( I => n19267, ZN => n19330);
   U4242 : INV_X2 port map( I => n20234, ZN => n20235);
   U20944 : NAND2_X2 port map( A1 => n18873, A2 => n180, ZN => n18399);
   U5916 : OAI21_X2 port map( A1 => n19805, A2 => n510, B => n11778, ZN => 
                           n22460);
   U4900 : INV_X2 port map( I => n19806, ZN => n11778);
   U3890 : NOR2_X2 port map( A1 => n28552, A2 => n20709, ZN => n13879);
   U3230 : NOR2_X2 port map( A1 => n18742, A2 => n8781, ZN => n24157);
   U18577 : INV_X2 port map( I => n17419, ZN => n17421);
   U20245 : NAND2_X2 port map( A1 => n15147, A2 => n15145, ZN => n20713);
   U172 : BUF_X4 port map( I => n20709, Z => n20899);
   U534 : NOR2_X2 port map( A1 => n9367, A2 => n19712, ZN => n9366);
   U1850 : NOR2_X2 port map( A1 => n3830, A2 => n9873, ZN => n6740);
   U21834 : NAND2_X2 port map( A1 => n9309, A2 => n9308, ZN => n24480);
   U17274 : AOI21_X2 port map( A1 => n4701, A2 => n881, B => n23594, ZN => 
                           n24483);
   U1871 : NAND2_X2 port map( A1 => n16337, A2 => n16339, ZN => n7142);
   U12811 : OAI21_X2 port map( A1 => n18747, A2 => n14362, B => n12931, ZN => 
                           n12996);
   U11592 : INV_X2 port map( I => n28552, ZN => n14806);
   U4074 : INV_X2 port map( I => n12910, ZN => n19287);
   U13228 : INV_X2 port map( I => n3502, ZN => n18755);
   U7646 : OAI21_X2 port map( A1 => n3289, A2 => n3288, B => n17987, ZN => 
                           n15136);
   U13386 : NOR2_X2 port map( A1 => n1271, A2 => n15864, ZN => n3780);
   U7214 : OAI22_X2 port map( A1 => n13226, A2 => n6981, B1 => n19869, B2 => 
                           n1130, ZN => n5301);
   U557 : INV_X2 port map( I => n10537, ZN => n18532);
   U812 : NAND2_X2 port map( A1 => n19167, A2 => n5990, ZN => n13490);
   U3440 : NOR2_X2 port map( A1 => n27640, A2 => n4192, ZN => n23692);
   U3220 : AOI22_X2 port map( A1 => n10239, A2 => n12521, B1 => n14791, B2 => 
                           n15429, ZN => n10238);
   U20605 : NOR2_X2 port map( A1 => n10304, A2 => n1053, ZN => n16432);
   U4302 : BUF_X4 port map( I => n619, Z => n17415);
   U3932 : NAND2_X2 port map( A1 => n21487, A2 => n10878, ZN => n15458);
   U950 : INV_X2 port map( I => n16209, ZN => n9308);
   U5368 : INV_X4 port map( I => n11962, ZN => n6688);
   U304 : NAND2_X2 port map( A1 => n7849, A2 => n19705, ZN => n7667);
   U21626 : OR2_X2 port map( A1 => n7817, A2 => n643, Z => n8425);
   U1390 : INV_X4 port map( I => n10533, ZN => n892);
   U2358 : NOR2_X2 port map( A1 => n6522, A2 => n852, ZN => n10547);
   U4454 : INV_X2 port map( I => n7138, ZN => n15674);
   U1864 : INV_X2 port map( I => n19201, ZN => n23117);
   U5924 : NAND2_X2 port map( A1 => n19747, A2 => n15667, ZN => n13148);
   U5667 : NAND3_X2 port map( A1 => n28457, A2 => n1207, A3 => n13350, ZN => 
                           n1706);
   U6638 : INV_X2 port map( I => n16998, ZN => n17175);
   U13231 : NAND2_X2 port map( A1 => n20336, A2 => n20153, ZN => n20337);
   U3551 : AND2_X1 port map( A1 => n25336, A2 => n16629, Z => n2607);
   U411 : OAI22_X2 port map( A1 => n21846, A2 => n209, B1 => n18866, B2 => 
                           n2218, ZN => n15207);
   U3578 : NAND3_X2 port map( A1 => n5718, A2 => n11143, A3 => n27072, ZN => 
                           n2596);
   U7497 : AOI21_X2 port map( A1 => n26701, A2 => n28160, B => n11280, ZN => 
                           n12950);
   U5784 : NOR2_X2 port map( A1 => n25984, A2 => n2798, ZN => n25850);
   U4226 : INV_X2 port map( I => n10435, ZN => n8976);
   U2525 : NAND3_X2 port map( A1 => n15186, A2 => n16690, A3 => n26734, ZN => 
                           n11360);
   U7202 : AOI21_X2 port map( A1 => n4088, A2 => n19941, B => n1120, ZN => 
                           n3497);
   U3880 : NAND2_X2 port map( A1 => n1164, A2 => n26640, ZN => n11840);
   U18688 : BUF_X4 port map( I => n18673, Z => n26121);
   U6161 : INV_X2 port map( I => n28237, ZN => n5055);
   U240 : NOR2_X2 port map( A1 => n19794, A2 => n8952, ZN => n5471);
   U15449 : NOR2_X2 port map( A1 => n23548, A2 => n10433, ZN => n3071);
   U475 : AOI21_X2 port map( A1 => n26631, A2 => n14502, B => n14382, ZN => 
                           n23774);
   U4742 : BUF_X2 port map( I => n5985, Z => n450);
   U4605 : OAI21_X2 port map( A1 => n25704, A2 => n15246, B => n3074, ZN => 
                           n3073);
   U9646 : INV_X2 port map( I => n18773, ZN => n18620);
   U3227 : OR2_X1 port map( A1 => n17435, A2 => n17198, Z => n7510);
   U910 : NOR2_X2 port map( A1 => n13502, A2 => n4199, ZN => n10205);
   U2648 : INV_X4 port map( I => n13548, ZN => n16679);
   U7965 : NAND2_X2 port map( A1 => n6936, A2 => n6935, ZN => n6934);
   U8257 : INV_X4 port map( I => n16332, ZN => n13990);
   U776 : INV_X2 port map( I => n823, ZN => n23041);
   U974 : INV_X2 port map( I => n8314, ZN => n4319);
   U8740 : AOI22_X2 port map( A1 => n12828, A2 => n26898, B1 => n20149, B2 => 
                           n6819, ZN => n12827);
   U264 : NOR2_X2 port map( A1 => n19974, A2 => n3439, ZN => n12828);
   U1081 : BUF_X4 port map( I => n8855, Z => n18588);
   U865 : NAND2_X2 port map( A1 => n2578, A2 => n2579, ZN => n2576);
   U154 : NOR2_X2 port map( A1 => n26436, A2 => n21616, ZN => n21589);
   U5096 : INV_X2 port map( I => n12251, ZN => n21286);
   U303 : NAND2_X2 port map( A1 => n6998, A2 => n5415, ZN => n24083);
   U13081 : NAND2_X2 port map( A1 => n18995, A2 => n19107, ZN => n18994);
   U18665 : INV_X2 port map( I => n11580, ZN => n18995);
   U12952 : NOR2_X2 port map( A1 => n6098, A2 => n3292, ZN => n7985);
   U20173 : INV_X4 port map( I => n15025, ZN => n16005);
   U10430 : NAND2_X2 port map( A1 => n443, A2 => n13389, ZN => n22494);
   U644 : NAND2_X2 port map( A1 => n28481, A2 => n1387, ZN => n8090);
   U22009 : AOI22_X2 port map( A1 => n5910, A2 => n11403, B1 => n20337, B2 => 
                           n20338, ZN => n1400);
   U13726 : NOR2_X2 port map( A1 => n1152, A2 => n22894, ZN => n4125);
   U4936 : AOI22_X2 port map( A1 => n23462, A2 => n10041, B1 => n19751, B2 => 
                           n23869, ZN => n9719);
   U488 : NAND2_X2 port map( A1 => n24579, A2 => n6987, ZN => n19598);
   U538 : NAND2_X2 port map( A1 => n15009, A2 => n15265, ZN => n25951);
   U8112 : NAND2_X1 port map( A1 => n8409, A2 => n16062, ZN => n2482);
   U4647 : INV_X2 port map( I => n5118, ZN => n16694);
   U6777 : OAI21_X2 port map( A1 => n21904, A2 => n15607, B => n25816, ZN => 
                           n3203);
   U244 : BUF_X4 port map( I => n6006, Z => n23642);
   U5855 : INV_X2 port map( I => n3830, ZN => n7752);
   U653 : INV_X2 port map( I => n12218, ZN => n865);
   U5303 : AND2_X2 port map( A1 => n7168, A2 => n1172, Z => n21825);
   U18352 : OAI21_X2 port map( A1 => n21757, A2 => n22981, B => n25894, ZN => 
                           n11996);
   U9624 : BUF_X2 port map( I => n9761, Z => n7190);
   U546 : INV_X2 port map( I => n649, ZN => n1001);
   U8251 : NOR2_X2 port map( A1 => n24882, A2 => n17367, ZN => n23118);
   U2255 : BUF_X2 port map( I => n18740, Z => n7212);
   U14719 : INV_X1 port map( I => n13660, ZN => n9813);
   U8148 : NAND2_X2 port map( A1 => n24081, A2 => n460, ZN => n8315);
   U18479 : NAND3_X2 port map( A1 => n24624, A2 => n26088, A3 => n26087, ZN => 
                           n8187);
   U6551 : AOI22_X2 port map( A1 => n4010, A2 => n24881, B1 => n5478, B2 => 
                           n24403, ZN => n22052);
   U648 : NAND2_X2 port map( A1 => n14255, A2 => n17981, ZN => n6592);
   U963 : INV_X2 port map( I => n19134, ZN => n13028);
   U2395 : NAND2_X2 port map( A1 => n22081, A2 => n8636, ZN => n4824);
   U5616 : NOR2_X2 port map( A1 => n632, A2 => n1022, ZN => n11264);
   U7185 : NAND2_X2 port map( A1 => n11079, A2 => n21769, ZN => n3678);
   U12281 : NAND2_X2 port map( A1 => n9105, A2 => n11937, ZN => n11910);
   U2844 : NAND2_X2 port map( A1 => n11580, A2 => n6778, ZN => n19105);
   U61 : AOI21_X2 port map( A1 => n708, A2 => n4742, B => n1087, ZN => n8060);
   U2810 : AOI21_X2 port map( A1 => n23645, A2 => n17683, B => n9480, ZN => 
                           n17620);
   U485 : AOI22_X2 port map( A1 => n9310, A2 => n24579, B1 => n24679, B2 => 
                           n6394, ZN => n25713);
   U5201 : INV_X2 port map( I => n8554, ZN => n18977);
   U314 : NOR2_X2 port map( A1 => n19917, A2 => n25236, ZN => n24364);
   U1540 : AOI21_X2 port map( A1 => n24442, A2 => n2177, B => n13171, ZN => 
                           n2178);
   U1298 : NAND2_X2 port map( A1 => n1786, A2 => n9149, ZN => n1785);
   U13171 : OAI21_X2 port map( A1 => n16653, A2 => n10597, B => n24552, ZN => 
                           n16566);
   U12502 : OAI21_X2 port map( A1 => n22703, A2 => n15751, B => n26008, ZN => 
                           n16643);
   U1085 : INV_X2 port map( I => n16972, ZN => n17563);
   U3936 : BUF_X2 port map( I => n8594, Z => n24327);
   U3613 : BUF_X2 port map( I => n24531, Z => n510);
   U1461 : BUF_X2 port map( I => n360, Z => n24774);
   U1234 : NAND2_X2 port map( A1 => n2910, A2 => n9691, ZN => n17637);
   U640 : AOI21_X2 port map( A1 => n19733, A2 => n13854, B => n2653, ZN => 
                           n2413);
   U9866 : NAND2_X2 port map( A1 => n17959, A2 => n23542, ZN => n15406);
   U3694 : NAND3_X2 port map( A1 => n13915, A2 => n13914, A3 => n1419, ZN => 
                           n7899);
   U13358 : INV_X2 port map( I => n15545, ZN => n21100);
   U12316 : INV_X4 port map( I => n20338, ZN => n5910);
   U3003 : AOI22_X2 port map( A1 => n9108, A2 => n14737, B1 => n9107, B2 => 
                           n11514, ZN => n22657);
   U218 : INV_X1 port map( I => n12533, ZN => n2998);
   U11496 : NOR2_X2 port map( A1 => n22164, A2 => n9573, ZN => n9571);
   U8846 : NAND2_X2 port map( A1 => n14284, A2 => n27029, ZN => n3910);
   U7382 : NOR2_X2 port map( A1 => n2394, A2 => n1331, ZN => n1330);
   U4372 : AOI21_X2 port map( A1 => n2716, A2 => n24496, B => n26710, ZN => 
                           n25860);
   U1480 : OAI21_X2 port map( A1 => n21791, A2 => n14342, B => n17847, ZN => 
                           n14351);
   U5496 : INV_X2 port map( I => n15255, ZN => n23571);
   U2356 : NOR2_X2 port map( A1 => n4385, A2 => n852, ZN => n6701);
   U4338 : BUF_X2 port map( I => n15916, Z => n1419);
   U2086 : INV_X2 port map( I => n574, ZN => n15760);
   U4156 : NOR2_X2 port map( A1 => n22399, A2 => n9989, ZN => n22506);
   U1537 : NOR2_X2 port map( A1 => n16433, A2 => n12331, ZN => n16503);
   U1220 : AOI22_X2 port map( A1 => n11264, A2 => n25903, B1 => n13486, B2 => 
                           n25966, ZN => n24932);
   U586 : INV_X2 port map( I => n19046, ZN => n24062);
   U40 : INV_X2 port map( I => n7039, ZN => n26059);
   U1920 : INV_X2 port map( I => n25322, ZN => n19633);
   U2919 : NAND2_X2 port map( A1 => n997, A2 => n27464, ZN => n19085);
   U5665 : INV_X2 port map( I => n13819, ZN => n17629);
   U7643 : OAI21_X2 port map( A1 => n17700, A2 => n1990, B => n18043, ZN => 
                           n14027);
   U2076 : NAND2_X2 port map( A1 => n18927, A2 => n22345, ZN => n13066);
   U4881 : INV_X2 port map( I => n9055, ZN => n13342);
   U734 : NAND2_X2 port map( A1 => n22856, A2 => n18424, ZN => n18425);
   U3125 : NOR2_X2 port map( A1 => n23000, A2 => n23001, ZN => n22195);
   U5878 : NAND2_X2 port map( A1 => n19819, A2 => n814, ZN => n19711);
   U5589 : INV_X4 port map( I => n2238, ZN => n23645);
   U6573 : OR2_X2 port map( A1 => n542, A2 => n24509, Z => n17440);
   U9068 : AOI21_X2 port map( A1 => n6279, A2 => n5571, B => n10690, ZN => 
                           n5570);
   U8096 : OAI21_X2 port map( A1 => n25287, A2 => n5062, B => n16632, ZN => 
                           n5061);
   U1200 : NAND2_X2 port map( A1 => n26681, A2 => n17952, ZN => n3304);
   U3733 : NOR2_X2 port map( A1 => n852, A2 => n21544, ZN => n6520);
   U1903 : NOR2_X2 port map( A1 => n19785, A2 => n28168, ZN => n19786);
   U2834 : NAND2_X2 port map( A1 => n9660, A2 => n27889, ZN => n24056);
   U470 : INV_X2 port map( I => n19088, ZN => n18920);
   U12824 : NAND2_X2 port map( A1 => n13009, A2 => n102, ZN => n21114);
   U7974 : INV_X4 port map( I => n1177, ZN => n24847);
   U2154 : INV_X2 port map( I => n13505, ZN => n20639);
   U729 : NOR2_X2 port map( A1 => n1177, A2 => n7168, ZN => n22873);
   U9532 : NOR2_X2 port map( A1 => n6312, A2 => n25828, ZN => n6311);
   U763 : OR2_X2 port map( A1 => n25381, A2 => n15326, Z => n1809);
   U2743 : INV_X2 port map( I => n22345, ZN => n18866);
   U9231 : NAND3_X2 port map( A1 => n22353, A2 => n9630, A3 => n25926, ZN => 
                           n23955);
   U6589 : INV_X2 port map( I => n8125, ZN => n1031);
   U3973 : BUF_X4 port map( I => n10494, Z => n26495);
   U6643 : INV_X1 port map( I => n9527, ZN => n901);
   U1115 : NAND2_X2 port map( A1 => n6430, A2 => n17605, ZN => n12619);
   U6328 : BUF_X2 port map( I => n704, Z => n22775);
   U1101 : NAND2_X2 port map( A1 => n1004, A2 => n18487, ZN => n18700);
   U6001 : OAI21_X2 port map( A1 => n11372, A2 => n25870, B => n20166, ZN => 
                           n22216);
   U1307 : NAND4_X2 port map( A1 => n13517, A2 => n20599, A3 => n20601, A4 => 
                           n20600, ZN => n24231);
   U12628 : INV_X2 port map( I => n25370, ZN => n21412);
   U8520 : NAND2_X2 port map( A1 => n18407, A2 => n233, ZN => n20);
   U2426 : OAI21_X2 port map( A1 => n20, A2 => n28019, B => n875, ZN => n5363);
   U4939 : BUF_X4 port map( I => n8467, Z => n4735);
   U12534 : NAND2_X2 port map( A1 => n4847, A2 => n4846, ZN => n7811);
   U1183 : INV_X2 port map( I => n26396, ZN => n16559);
   U3106 : NOR2_X2 port map( A1 => n10224, A2 => n10221, ZN => n23599);
   U13360 : INV_X2 port map( I => n11215, ZN => n26485);
   U3309 : OR2_X1 port map( A1 => n17302, A2 => n1629, Z => n3110);
   U4208 : INV_X4 port map( I => n7421, ZN => n708);
   U3326 : NOR3_X2 port map( A1 => n13925, A2 => n15717, A3 => n20430, ZN => 
                           n6801);
   U11257 : INV_X1 port map( I => n18665, ZN => n26031);
   U861 : OAI21_X2 port map( A1 => n25850, A2 => n15202, B => n778, ZN => n7372
                           );
   U783 : AOI21_X2 port map( A1 => n25732, A2 => n24730, B => n24971, ZN => 
                           n1846);
   U4669 : AOI21_X2 port map( A1 => n6834, A2 => n24573, B => n998, ZN => n1581
                           );
   U1260 : NOR2_X2 port map( A1 => n12590, A2 => n23002, ZN => n25532);
   U2634 : INV_X2 port map( I => n10474, ZN => n10323);
   U3229 : OAI21_X2 port map( A1 => n9917, A2 => n24167, B => n25583, ZN => 
                           n10119);
   U8664 : INV_X2 port map( I => n20502, ZN => n20728);
   U7904 : NAND2_X1 port map( A1 => n4715, A2 => n28389, ZN => n7449);
   U1884 : BUF_X4 port map( I => n13685, Z => n11372);
   U7350 : AND2_X2 port map( A1 => n23002, A2 => n7553, Z => n3943);
   U744 : BUF_X4 port map( I => n18527, Z => n11685);
   U1991 : NAND2_X2 port map( A1 => n23578, A2 => n27431, ZN => n13934);
   U2851 : NAND3_X2 port map( A1 => n21630, A2 => n28433, A3 => n21668, ZN => 
                           n15500);
   U13736 : OAI21_X2 port map( A1 => n19624, A2 => n12444, B => n866, ZN => 
                           n22901);
   U12580 : OAI21_X2 port map( A1 => n23966, A2 => n11299, B => n9869, ZN => 
                           n11300);
   U3171 : NAND3_X2 port map( A1 => n12949, A2 => n12726, A3 => n8223, ZN => 
                           n7756);
   U817 : AOI21_X2 port map( A1 => n10748, A2 => n5502, B => n9059, ZN => 
                           n11042);
   U9318 : NAND2_X2 port map( A1 => n14441, A2 => n19005, ZN => n19007);
   U15725 : NAND2_X2 port map( A1 => n23682, A2 => n21860, ZN => n19793);
   U3408 : NAND2_X2 port map( A1 => n15187, A2 => n19140, ZN => n18871);
   U9904 : NAND2_X2 port map( A1 => n5568, A2 => n27201, ZN => n5566);
   U3163 : AOI22_X2 port map( A1 => n7648, A2 => n26114, B1 => n7647, B2 => 
                           n8223, ZN => n24168);
   U1271 : NOR2_X2 port map( A1 => n12850, A2 => n12676, ZN => n13657);
   U8526 : NOR2_X1 port map( A1 => n10482, A2 => n20780, ZN => n5302);
   U293 : INV_X2 port map( I => n3497, ZN => n1607);
   U2228 : NAND2_X2 port map( A1 => n10267, A2 => n10708, ZN => n15142);
   U1583 : NOR2_X2 port map( A1 => n9829, A2 => n13964, ZN => n26240);
   U2310 : INV_X4 port map( I => n756, ZN => n3861);
   U3617 : NOR2_X2 port map( A1 => n19055, A2 => n12571, ZN => n18796);
   U5747 : NOR2_X2 port map( A1 => n7759, A2 => n913, ZN => n11894);
   U1088 : NOR2_X2 port map( A1 => n18723, A2 => n14332, ZN => n25067);
   U12479 : OR2_X2 port map( A1 => n24234, A2 => n3527, Z => n17384);
   U13103 : NOR2_X2 port map( A1 => n756, A2 => n26621, ZN => n15118);
   U4405 : OAI21_X2 port map( A1 => n1116, A2 => n19848, B => n14726, ZN => 
                           n7325);
   U9823 : INV_X2 port map( I => n17844, ZN => n1870);
   U18714 : NOR2_X2 port map( A1 => n10993, A2 => n27497, ZN => n14924);
   U4380 : NAND2_X2 port map( A1 => n25155, A2 => n25154, ZN => n24919);
   U5887 : INV_X4 port map( I => n11936, ZN => n1118);
   U3382 : AOI22_X2 port map( A1 => n4290, A2 => n28184, B1 => n1189, B2 => 
                           n8604, ZN => n22449);
   U12435 : OAI21_X2 port map( A1 => n13019, A2 => n13018, B => n21100, ZN => 
                           n22451);
   U427 : INV_X4 port map( I => n25421, ZN => n675);
   U8882 : NAND2_X2 port map( A1 => n808, A2 => n19664, ZN => n5307);
   U15253 : INV_X2 port map( I => n5816, ZN => n21686);
   U4180 : NAND2_X2 port map( A1 => n2777, A2 => n12061, ZN => n5816);
   U458 : AOI21_X2 port map( A1 => n14735, A2 => n14734, B => n4929, ZN => 
                           n20200);
   U2874 : INV_X4 port map( I => n238, ZN => n914);
   U2872 : AOI21_X2 port map( A1 => n238, A2 => n24216, B => n797, ZN => n2687)
                           ;
   U1429 : INV_X2 port map( I => n4797, ZN => n24981);
   U20145 : NAND2_X2 port map( A1 => n13788, A2 => n5877, ZN => n18931);
   U5877 : INV_X2 port map( I => n10593, ZN => n19919);
   U2607 : INV_X4 port map( I => n27043, ZN => n2798);
   U19119 : NOR2_X2 port map( A1 => n23887, A2 => n23886, ZN => n1114);
   U108 : INV_X2 port map( I => n10558, ZN => n2093);
   U2638 : BUF_X4 port map( I => n15234, Z => n13979);
   U1236 : NAND2_X2 port map( A1 => n17701, A2 => n9040, ZN => n1990);
   U547 : NAND2_X2 port map( A1 => n14883, A2 => n18757, ZN => n18490);
   U792 : INV_X2 port map( I => n18173, ZN => n18044);
   U20130 : NOR2_X2 port map( A1 => n24056, A2 => n3654, ZN => n10347);
   U275 : AOI22_X2 port map( A1 => n856, A2 => n22807, B1 => n7731, B2 => n733,
                           ZN => n1573);
   U1951 : NAND2_X2 port map( A1 => n21898, A2 => n4610, ZN => n17812);
   U1751 : NOR2_X2 port map( A1 => n7062, A2 => n7063, ZN => n4912);
   U1726 : INV_X2 port map( I => n24643, ZN => n22370);
   U4458 : INV_X4 port map( I => n632, ZN => n2238);
   U19866 : INV_X2 port map( I => n5683, ZN => n21511);
   U2910 : BUF_X4 port map( I => n12500, Z => n24552);
   U2906 : BUF_X2 port map( I => n12500, Z => n24550);
   U4864 : OAI21_X2 port map( A1 => n18233, A2 => n23138, B => n18808, ZN => 
                           n23430);
   U496 : NAND2_X2 port map( A1 => n10243, A2 => n10242, ZN => n488);
   U21507 : NOR2_X2 port map( A1 => n26432, A2 => n26431, ZN => n26430);
   U21514 : NAND2_X2 port map( A1 => n15679, A2 => n923, ZN => n26431);
   U12408 : NOR2_X2 port map( A1 => n1383, A2 => n14334, ZN => n15411);
   U957 : OAI21_X2 port map( A1 => n23534, A2 => n18693, B => n25802, ZN => 
                           n26465);
   U3383 : AOI21_X2 port map( A1 => n22326, A2 => n22325, B => n8604, ZN => 
                           n2150);
   U11475 : NOR2_X2 port map( A1 => n15812, A2 => n25225, ZN => n25234);
   U7041 : INV_X2 port map( I => n13432, ZN => n1080);
   U186 : NOR2_X2 port map( A1 => n24554, A2 => n806, ZN => n683);
   U5652 : NAND2_X2 port map( A1 => n24142, A2 => n787, ZN => n21827);
   U5354 : CLKBUF_X4 port map( I => n6687, Z => n2045);
   U12889 : INV_X2 port map( I => n22421, ZN => n3530);
   U3222 : INV_X2 port map( I => n12434, ZN => n16511);
   U6035 : INV_X2 port map( I => n3706, ZN => n12279);
   U8101 : AOI21_X1 port map( A1 => n22889, A2 => n18605, B => n22217, ZN => 
                           n12967);
   U66 : OAI21_X2 port map( A1 => n3938, A2 => n3826, B => n24327, ZN => n3825)
                           ;
   U13412 : NAND2_X2 port map( A1 => n24573, A2 => n28019, ZN => n19064);
   U3735 : NAND2_X2 port map( A1 => n22823, A2 => n21544, ZN => n4385);
   U2948 : INV_X2 port map( I => n11124, ZN => n21995);
   U5968 : NOR2_X2 port map( A1 => n11213, A2 => n754, ZN => n19763);
   U123 : NAND2_X2 port map( A1 => n20642, A2 => n21715, ZN => n20645);
   U5090 : BUF_X2 port map( I => n616, Z => n25971);
   U4325 : INV_X1 port map( I => n16314, ZN => n15075);
   U4638 : INV_X2 port map( I => n17198, ZN => n17508);
   U2656 : NAND2_X2 port map( A1 => n18424, A2 => n18574, ZN => n18675);
   U1328 : BUF_X2 port map( I => n14552, Z => n25493);
   U6152 : INV_X2 port map( I => n19883, ZN => n19742);
   U7055 : OAI21_X2 port map( A1 => n8471, A2 => n4624, B => n18821, ZN => 
                           n18824);
   U2669 : INV_X2 port map( I => n17522, ZN => n4888);
   U202 : AND2_X2 port map( A1 => n7561, A2 => n23687, Z => n21671);
   U1336 : INV_X2 port map( I => n28295, ZN => n1512);
   U9794 : INV_X4 port map( I => n4812, ZN => n4063);
   U3068 : BUF_X4 port map( I => n6447, Z => n2726);
   U3874 : OAI21_X2 port map( A1 => n9379, A2 => n24119, B => n16673, ZN => 
                           n16675);
   U233 : INV_X4 port map( I => n24720, ZN => n19974);
   U3477 : INV_X2 port map( I => n679, ZN => n10520);
   U1813 : INV_X2 port map( I => n11488, ZN => n17954);
   U15790 : NOR2_X2 port map( A1 => n22396, A2 => n6770, ZN => n8221);
   U7380 : INV_X2 port map( I => n26920, ZN => n10164);
   U1451 : BUF_X4 port map( I => n14859, Z => n3091);
   U5824 : NAND2_X2 port map( A1 => n18994, A2 => n8133, ZN => n19094);
   U3906 : INV_X4 port map( I => n778, ZN => n23597);
   U3270 : INV_X2 port map( I => n22487, ZN => n9524);
   U21131 : NAND2_X2 port map( A1 => n19726, A2 => n19858, ZN => n19585);
   U530 : INV_X1 port map( I => n15623, ZN => n1188);
   U11295 : INV_X2 port map( I => n13571, ZN => n19842);
   U3891 : NOR2_X2 port map( A1 => n9167, A2 => n24283, ZN => n8459);
   U3530 : BUF_X4 port map( I => n20471, Z => n21724);
   U18536 : INV_X2 port map( I => n18410, ZN => n18693);
   U8003 : NOR2_X2 port map( A1 => n1042, A2 => n13927, ZN => n9616);
   U2043 : NAND2_X2 port map( A1 => n7165, A2 => n7168, ZN => n18409);
   U401 : NOR2_X2 port map( A1 => n1156, A2 => n997, ZN => n19087);
   U4018 : INV_X2 port map( I => n18309, ZN => n22556);
   U12620 : OAI21_X2 port map( A1 => n8491, A2 => n8492, B => n27924, ZN => 
                           n8493);
   U3728 : AOI21_X2 port map( A1 => n6522, A2 => n21544, B => n22823, ZN => 
                           n21440);
   U1396 : NAND2_X2 port map( A1 => n17490, A2 => n15189, ZN => n25140);
   U10435 : NAND2_X2 port map( A1 => n7142, A2 => n15965, ZN => n9309);
   U12614 : NOR2_X2 port map( A1 => n27924, A2 => n13505, ZN => n3938);
   U1318 : BUF_X4 port map( I => n5402, Z => n22312);
   U5322 : CLKBUF_X4 port map( I => n13242, Z => n6345);
   U2477 : NOR2_X2 port map( A1 => n28166, A2 => n1062, ZN => n15921);
   U1610 : INV_X2 port map( I => n9978, ZN => n912);
   U5562 : NOR2_X2 port map( A1 => n21767, A2 => n27043, ZN => n3524);
   U13561 : NOR2_X2 port map( A1 => n404, A2 => n703, ZN => n15438);
   U5226 : BUF_X2 port map( I => n9261, Z => n390);
   U13028 : NOR2_X2 port map( A1 => n8221, A2 => n100, ZN => n8220);
   U16973 : NAND2_X2 port map( A1 => n7282, A2 => n8648, ZN => n13783);
   U3402 : OAI21_X2 port map( A1 => n16409, A2 => n9116, B => n23439, ZN => 
                           n14173);
   U918 : INV_X2 port map( I => n14580, ZN => n19089);
   U7182 : AOI21_X2 port map( A1 => n10733, A2 => n27984, B => n14973, ZN => 
                           n20199);
   U6829 : NAND2_X2 port map( A1 => n8926, A2 => n16120, ZN => n16118);
   U11980 : OAI21_X2 port map( A1 => n9502, A2 => n9503, B => n16822, ZN => 
                           n2980);
   U4644 : OAI21_X2 port map( A1 => n26013, A2 => n26014, B => n998, ZN => 
                           n25823);
   U12561 : AOI22_X2 port map( A1 => n8236, A2 => n25431, B1 => n9264, B2 => 
                           n8235, ZN => n22043);
   U10373 : AOI21_X2 port map( A1 => n16019, A2 => n16018, B => n16146, ZN => 
                           n16023);
   U3257 : INV_X1 port map( I => n15227, ZN => n21783);
   U12635 : OAI21_X2 port map( A1 => n24261, A2 => n15249, B => n26435, ZN => 
                           n22691);
   U194 : INV_X2 port map( I => n24680, ZN => n26435);
   U20994 : OAI21_X2 port map( A1 => n18709, A2 => n14207, B => n12711, ZN => 
                           n18702);
   U5415 : INV_X2 port map( I => n5197, ZN => n16488);
   U3424 : BUF_X4 port map( I => n18694, Z => n18697);
   U15624 : INV_X2 port map( I => n23474, ZN => n25685);
   U1472 : OAI21_X2 port map( A1 => n23531, A2 => n14177, B => n16370, ZN => 
                           n25801);
   U12158 : NAND2_X2 port map( A1 => n19117, A2 => n7609, ZN => n4079);
   U3443 : INV_X2 port map( I => n8311, ZN => n8447);
   U11457 : NAND2_X2 port map( A1 => n797, A2 => n1266, ZN => n16355);
   U577 : INV_X2 port map( I => n25099, ZN => n23268);
   U5642 : NAND2_X2 port map( A1 => n17874, A2 => n17894, ZN => n18043);
   U5462 : OAI21_X2 port map( A1 => n22342, A2 => n26065, B => n14090, ZN => 
                           n8698);
   U5742 : BUF_X2 port map( I => n2013, Z => n26321);
   U584 : INV_X2 port map( I => n9994, ZN => n19821);
   U12563 : OAI21_X2 port map( A1 => n8236, A2 => n23913, B => n8265, ZN => 
                           n8234);
   U12475 : AOI21_X2 port map( A1 => n27023, A2 => n13979, B => n21620, ZN => 
                           n23990);
   U5705 : NOR2_X2 port map( A1 => n18583, A2 => n1013, ZN => n23390);
   U6606 : INV_X2 port map( I => n12225, ZN => n17323);
   U18940 : INV_X1 port map( I => n16193, ZN => n14197);
   U1924 : OAI21_X2 port map( A1 => n20338, A2 => n19985, B => n20336, ZN => 
                           n7396);
   U16466 : INV_X2 port map( I => n18142, ZN => n18290);
   U1715 : INV_X4 port map( I => n7053, ZN => n836);
   U4893 : NOR2_X2 port map( A1 => n12441, A2 => n19945, ZN => n9995);
   U5296 : NOR2_X2 port map( A1 => n12116, A2 => n16127, ZN => n15996);
   U2141 : NOR2_X2 port map( A1 => n10293, A2 => n15560, ZN => n12441);
   U1475 : NOR2_X2 port map( A1 => n26593, A2 => n13953, ZN => n23301);
   U11565 : NAND2_X2 port map( A1 => n22912, A2 => n15068, ZN => n6245);
   U20504 : NOR2_X1 port map( A1 => n15918, A2 => n14197, ZN => n15857);
   U380 : BUF_X4 port map( I => n24553, Z => n24554);
   U15598 : NOR2_X2 port map( A1 => n18588, A2 => n820, ZN => n18547);
   U2423 : AOI21_X2 port map( A1 => n6835, A2 => n6834, B => n875, ZN => n3170)
                           ;
   U1667 : OAI21_X2 port map( A1 => n12690, A2 => n10121, B => n813, ZN => 
                           n12689);
   U2580 : NOR2_X2 port map( A1 => n11294, A2 => n11292, ZN => n4999);
   U743 : OAI21_X2 port map( A1 => n19026, A2 => n19154, B => n22860, ZN => 
                           n9674);
   U47 : BUF_X4 port map( I => n21563, Z => n10385);
   U3679 : INV_X2 port map( I => n19669, ZN => n23216);
   U4988 : NAND2_X2 port map( A1 => n22901, A2 => n28425, ZN => n13650);
   U17817 : INV_X2 port map( I => n19133, ZN => n18929);
   U13498 : AOI22_X2 port map( A1 => n13758, A2 => n14177, B1 => n2976, B2 => 
                           n16466, ZN => n2975);
   U14360 : OAI21_X2 port map( A1 => n15434, A2 => n12521, B => n13, ZN => 
                           n25494);
   U14894 : NAND2_X1 port map( A1 => n17870, A2 => n14284, ZN => n23288);
   U25 : INV_X2 port map( I => n9611, ZN => n940);
   U1763 : INV_X2 port map( I => n17345, ZN => n17227);
   U6031 : OAI21_X2 port map( A1 => n19665, A2 => n808, B => n5307, ZN => 
                           n10288);
   U2300 : AOI22_X2 port map( A1 => n10931, A2 => n751, B1 => n25959, B2 => 
                           n287, ZN => n19665);
   U21841 : INV_X2 port map( I => n24487, ZN => n613);
   U1546 : NOR2_X2 port map( A1 => n14177, A2 => n16461, ZN => n26175);
   U8160 : NOR2_X2 port map( A1 => n15878, A2 => n10452, ZN => n10451);
   U4070 : INV_X4 port map( I => n10810, ZN => n751);
   U213 : INV_X4 port map( I => n13301, ZN => n12659);
   U10386 : NOR2_X2 port map( A1 => n8347, A2 => n9792, ZN => n8346);
   U1883 : INV_X4 port map( I => n11319, ZN => n20842);
   U2583 : NOR2_X2 port map( A1 => n16134, A2 => n16132, ZN => n9792);
   U6909 : INV_X2 port map( I => n21343, ZN => n2450);
   U5213 : NAND3_X1 port map( A1 => n21848, A2 => n14539, A3 => n14017, ZN => 
                           n23805);
   U4067 : INV_X2 port map( I => n26302, ZN => n18256);
   U5782 : NAND2_X2 port map( A1 => n16321, A2 => n9095, ZN => n16157);
   U2565 : NOR2_X2 port map( A1 => n7970, A2 => n27465, ZN => n3156);
   U5527 : NAND2_X2 port map( A1 => n12236, A2 => n1037, ZN => n17234);
   U6245 : AOI21_X2 port map( A1 => n23126, A2 => n444, B => n18933, ZN => 
                           n8729);
   U1831 : NAND2_X2 port map( A1 => n11778, A2 => n968, ZN => n19770);
   U13068 : INV_X4 port map( I => n15812, ZN => n16083);
   U5382 : AOI22_X2 port map( A1 => n15812, A2 => n5050, B1 => n16254, B2 => 
                           n16255, ZN => n5051);
   U5128 : INV_X2 port map( I => n7228, ZN => n24470);
   U3076 : BUF_X2 port map( I => n15119, Z => n24197);
   U1798 : NAND4_X1 port map( A1 => n8759, A2 => n8758, A3 => n20999, A4 => 
                           n13272, ZN => n26592);
   U13543 : BUF_X2 port map( I => n5505, Z => n25382);
   U271 : INV_X2 port map( I => n11225, ZN => n12512);
   U6099 : NAND2_X2 port map( A1 => n28552, A2 => n20901, ZN => n20757);
   U1621 : BUF_X4 port map( I => n16567, Z => n434);
   U2473 : INV_X4 port map( I => n814, ZN => n12666);
   U12619 : OAI21_X2 port map( A1 => n27924, A2 => n20639, B => n28553, ZN => 
                           n6542);
   U2510 : INV_X2 port map( I => n25559, ZN => n19165);
   U3186 : INV_X2 port map( I => n12477, ZN => n23913);
   U10509 : INV_X2 port map( I => n16267, ZN => n6317);
   U683 : NOR2_X2 port map( A1 => n19726, A2 => n10613, ZN => n8837);
   U6382 : INV_X2 port map( I => n14649, ZN => n1174);
   U5858 : NOR2_X2 port map( A1 => n990, A2 => n13371, ZN => n26222);
   U20018 : BUF_X4 port map( I => n15796, Z => n16271);
   U3294 : INV_X2 port map( I => n13662, ZN => n1169);
   U210 : NOR2_X2 port map( A1 => n15697, A2 => n6547, ZN => n10795);
   U8849 : NAND2_X2 port map( A1 => n24946, A2 => n17623, ZN => n7090);
   U8750 : NAND2_X2 port map( A1 => n20413, A2 => n14262, ZN => n6716);
   U3644 : NOR2_X2 port map( A1 => n16524, A2 => n3537, ZN => n13608);
   U7409 : NAND2_X1 port map( A1 => n25550, A2 => n22299, ZN => n24781);
   U3700 : OAI22_X1 port map( A1 => n21801, A2 => n15667, B1 => n19168, B2 => 
                           n24187, ZN => n22612);
   U6485 : OAI22_X2 port map( A1 => n24337, A2 => n27856, B1 => n22775, B2 => 
                           n12617, ZN => n5836);
   U2617 : CLKBUF_X4 port map( I => n4719, Z => n24330);
   U321 : INV_X2 port map( I => n19700, ZN => n26459);
   U13603 : INV_X2 port map( I => n10554, ZN => n21025);
   U1878 : NAND2_X2 port map( A1 => n10554, A2 => n21024, ZN => n12160);
   U10291 : NOR2_X2 port map( A1 => n16401, A2 => n16644, ZN => n14965);
   U1585 : BUF_X4 port map( I => n16612, Z => n14562);
   U3822 : INV_X2 port map( I => n21534, ZN => n21528);
   U4051 : NOR2_X2 port map( A1 => n9078, A2 => n12169, ZN => n9077);
   U10031 : NOR2_X1 port map( A1 => n14658, A2 => n9018, ZN => n17219);
   U9335 : OAI21_X2 port map( A1 => n10563, A2 => n17407, B => n8237, ZN => 
                           n9686);
   U11587 : OR2_X1 port map( A1 => n16639, A2 => n2179, Z => n4597);
   U21750 : NOR2_X2 port map( A1 => n9642, A2 => n19009, ZN => n24424);
   U8842 : INV_X4 port map( I => n22202, ZN => n22307);
   U15663 : OAI21_X2 port map( A1 => n1216, A2 => n8314, B => n17542, ZN => 
                           n17852);
   U3067 : AND2_X1 port map( A1 => n6447, A2 => n14210, Z => n26336);
   U15638 : INV_X2 port map( I => n23307, ZN => n4657);
   U897 : INV_X2 port map( I => n24089, ZN => n1247);
   U19724 : INV_X2 port map( I => n26254, ZN => n8534);
   U2460 : BUF_X4 port map( I => n3109, Z => n21767);
   U578 : BUF_X2 port map( I => n3109, Z => n21765);
   U6919 : NAND2_X2 port map( A1 => n22087, A2 => n2782, ZN => n3109);
   U13205 : AOI22_X2 port map( A1 => n3217, A2 => n24421, B1 => n253, B2 => 
                           n27385, ZN => n8506);
   U4013 : BUF_X4 port map( I => n10027, Z => n699);
   U5416 : NOR2_X2 port map( A1 => n13758, A2 => n4162, ZN => n23530);
   U1180 : INV_X2 port map( I => n27344, ZN => n11702);
   U13016 : NAND2_X2 port map( A1 => n23064, A2 => n4318, ZN => n23042);
   U13510 : INV_X2 port map( I => n3843, ZN => n6293);
   U12531 : NAND2_X2 port map( A1 => n20124, A2 => n8265, ZN => n3138);
   U3189 : NAND2_X2 port map( A1 => n3803, A2 => n12477, ZN => n20122);
   U15343 : INV_X1 port map( I => n5969, ZN => n13811);
   U5567 : AOI21_X2 port map( A1 => n2835, A2 => n17460, B => n897, ZN => 
                           n15305);
   U3070 : OAI22_X2 port map( A1 => n8447, A2 => n26914, B1 => n20749, B2 => 
                           n6589, ZN => n20754);
   U7172 : INV_X4 port map( I => n14683, ZN => n1012);
   U727 : INV_X2 port map( I => n25767, ZN => n6539);
   U6990 : AOI21_X2 port map( A1 => n15316, A2 => n20403, B => n15315, ZN => 
                           n15314);
   U4356 : BUF_X2 port map( I => n23825, Z => n25023);
   U3001 : OR2_X1 port map( A1 => n6219, A2 => n15619, Z => n15618);
   U14631 : INV_X2 port map( I => n14162, ZN => n18959);
   U1104 : INV_X2 port map( I => n15352, ZN => n21689);
   U8528 : INV_X1 port map( I => n20680, ZN => n7698);
   U576 : AND2_X2 port map( A1 => n19899, A2 => n21788, Z => n24639);
   U15761 : NAND2_X2 port map( A1 => n18379, A2 => n24133, ZN => n6731);
   U2730 : INV_X4 port map( I => n9464, ZN => n24092);
   U1848 : NAND2_X2 port map( A1 => n8180, A2 => n3741, ZN => n17360);
   U2495 : BUF_X2 port map( I => n10175, Z => n95);
   U6090 : NAND2_X2 port map( A1 => n2085, A2 => n5057, ZN => n21989);
   U12625 : AOI21_X2 port map( A1 => n9672, A2 => n20645, B => n3995, ZN => 
                           n3994);
   U5499 : BUF_X4 port map( I => n8314, Z => n4318);
   U12331 : AOI21_X2 port map( A1 => n17528, A2 => n17527, B => n10015, ZN => 
                           n4320);
   U3634 : INV_X2 port map( I => n16524, ZN => n16725);
   U20056 : INV_X1 port map( I => n10045, ZN => n11812);
   U1729 : INV_X2 port map( I => n15565, ZN => n25763);
   U5078 : INV_X1 port map( I => n15565, ZN => n16230);
   U16353 : INV_X2 port map( I => n23448, ZN => n17036);
   U11711 : AOI21_X2 port map( A1 => n15534, A2 => n15533, B => n4319, ZN => 
                           n22689);
   U1330 : NOR2_X2 port map( A1 => n12197, A2 => n20890, ZN => n5196);
   U1072 : NOR2_X2 port map( A1 => n9370, A2 => n14859, ZN => n23797);
   U650 : INV_X2 port map( I => n25644, ZN => n19928);
   U4854 : OR2_X2 port map( A1 => n11719, A2 => n9619, Z => n18479);
   U463 : INV_X2 port map( I => n20, ZN => n998);
   U1219 : NAND2_X2 port map( A1 => n22485, A2 => n17681, ZN => n2287);
   U19044 : INV_X2 port map( I => n18549, ZN => n18728);
   U8574 : NAND2_X1 port map( A1 => n7671, A2 => n20591, ZN => n7192);
   U20428 : OAI22_X1 port map( A1 => n17612, A2 => n237, B1 => n17614, B2 => 
                           n1217, ZN => n17613);
   U7829 : OAI21_X2 port map( A1 => n15037, A2 => n5353, B => n17518, ZN => 
                           n5092);
   U1881 : NOR3_X2 port map( A1 => n10554, A2 => n21024, A3 => n708, ZN => 
                           n12197);
   U5751 : AOI22_X2 port map( A1 => n12573, A2 => n27739, B1 => n3902, B2 => 
                           n1175, ZN => n1874);
   U2516 : INV_X4 port map( I => n10015, ZN => n17529);
   U7889 : NOR2_X2 port map( A1 => n7901, A2 => n4417, ZN => n4416);
   U3953 : NAND2_X2 port map( A1 => n464, A2 => n24601, ZN => n23846);
   U6025 : NAND2_X2 port map( A1 => n9760, A2 => n11462, ZN => n21298);
   U12840 : NAND2_X1 port map( A1 => n16527, A2 => n4998, ZN => n9373);
   U6848 : INV_X2 port map( I => n14174, ZN => n15930);
   U8857 : NAND2_X1 port map( A1 => n7734, A2 => n7732, ZN => n1572);
   U3793 : INV_X2 port map( I => n11658, ZN => n835);
   U14783 : NAND3_X2 port map( A1 => n26705, A2 => n10701, A3 => n1580, ZN => 
                           n25552);
   U366 : INV_X2 port map( I => n8399, ZN => n10447);
   U4756 : NOR2_X2 port map( A1 => n12245, A2 => n5250, ZN => n7788);
   U227 : NAND2_X2 port map( A1 => n2199, A2 => n25830, ZN => n25362);
   U1016 : NOR2_X2 port map( A1 => n23199, A2 => n18465, ZN => n26159);
   U11535 : AOI21_X2 port map( A1 => n13184, A2 => n10958, B => n18505, ZN => 
                           n15085);
   U1632 : NOR2_X2 port map( A1 => n15988, A2 => n22932, ZN => n24773);
   U9635 : INV_X2 port map( I => n9699, ZN => n1175);
   U7324 : INV_X2 port map( I => n19516, ZN => n10331);
   U10049 : NAND2_X2 port map( A1 => n8770, A2 => n3545, ZN => n1799);
   U12578 : NOR2_X1 port map( A1 => n5294, A2 => n11299, ZN => n26044);
   U10458 : NOR2_X2 port map( A1 => n14948, A2 => n15878, ZN => n8347);
   U5583 : OAI21_X2 port map( A1 => n24502, A2 => n10725, B => n25796, ZN => 
                           n13957);
   U4351 : INV_X2 port map( I => n2710, ZN => n25636);
   U11954 : NOR2_X2 port map( A1 => n18929, A2 => n2516, ZN => n13105);
   U18001 : NAND2_X2 port map( A1 => n24664, A2 => n994, ZN => n23732);
   U9936 : OAI21_X2 port map( A1 => n17344, A2 => n23787, B => n12506, ZN => 
                           n13055);
   U9103 : OAI21_X1 port map( A1 => n6861, A2 => n19730, B => n8208, ZN => 
                           n19596);
   U9799 : NAND3_X2 port map( A1 => n17834, A2 => n4590, A3 => n17833, ZN => 
                           n17835);
   U2674 : BUF_X4 port map( I => n17261, Z => n17519);
   U6822 : NAND2_X2 port map( A1 => n16134, A2 => n15926, ZN => n9892);
   U3176 : OAI21_X2 port map( A1 => n22472, A2 => n22471, B => n23405, ZN => 
                           n6443);
   U6171 : INV_X2 port map( I => n24351, ZN => n5227);
   U15215 : AOI21_X2 port map( A1 => n28081, A2 => n835, B => n13481, ZN => 
                           n5757);
   U12558 : INV_X4 port map( I => n6339, ZN => n21734);
   U1006 : AOI21_X2 port map( A1 => n24047, A2 => n23743, B => n25718, ZN => 
                           n24045);
   U5661 : NAND2_X2 port map( A1 => n11327, A2 => n7451, ZN => n7450);
   U5938 : INV_X2 port map( I => n8326, ZN => n10611);
   U290 : INV_X2 port map( I => n19849, ZN => n1116);
   U1012 : BUF_X2 port map( I => n27780, Z => n14634);
   U13469 : NOR2_X2 port map( A1 => n1256, A2 => n24552, ZN => n16564);
   U4931 : NAND2_X1 port map( A1 => n11236, A2 => n19768, ZN => n11235);
   U4724 : AOI21_X2 port map( A1 => n22329, A2 => n12989, B => n18613, ZN => 
                           n26233);
   U7306 : INV_X2 port map( I => n13387, ZN => n971);
   U968 : NAND2_X2 port map( A1 => n18615, A2 => n24895, ZN => n18616);
   U6008 : INV_X4 port map( I => n9175, ZN => n14179);
   U2785 : OR2_X1 port map( A1 => n16534, A2 => n6766, Z => n25289);
   U12339 : NOR2_X2 port map( A1 => n5141, A2 => n21136, ZN => n12944);
   U2640 : AND2_X2 port map( A1 => n21456, A2 => n15234, Z => n552);
   U4738 : NAND2_X2 port map( A1 => n25891, A2 => n11817, ZN => n25233);
   U5633 : BUF_X2 port map( I => n6144, Z => n3106);
   U3239 : OR2_X1 port map( A1 => n4070, A2 => n2897, Z => n17787);
   U642 : NAND3_X1 port map( A1 => n9923, A2 => n7581, A3 => n18588, ZN => 
                           n5936);
   U10037 : INV_X2 port map( I => n21754, ZN => n17426);
   U2371 : OR2_X2 port map( A1 => n6575, A2 => n17324, Z => n21754);
   U2189 : NAND2_X2 port map( A1 => n14153, A2 => n675, ZN => n20108);
   U8139 : OAI21_X2 port map( A1 => n12535, A2 => n12536, B => n1259, ZN => 
                           n2497);
   U5902 : BUF_X2 port map( I => n19757, Z => n8192);
   U4174 : BUF_X4 port map( I => n15255, Z => n9358);
   U15182 : NAND2_X1 port map( A1 => n11121, A2 => n5683, ZN => n11120);
   U6675 : INV_X2 port map( I => n12973, ZN => n22066);
   U964 : NAND2_X2 port map( A1 => n26598, A2 => n24092, ZN => n7787);
   U13954 : NOR3_X1 port map( A1 => n4403, A2 => n6681, A3 => n14062, ZN => 
                           n4402);
   U18550 : INV_X2 port map( I => n11816, ZN => n11817);
   U9967 : AOI21_X2 port map( A1 => n20570, A2 => n7060, B => n24421, ZN => 
                           n22438);
   U7092 : NAND2_X2 port map( A1 => n26637, A2 => n3460, ZN => n4911);
   U20870 : AOI21_X2 port map( A1 => n17999, A2 => n1020, B => n4976, ZN => 
                           n18000);
   U4273 : BUF_X2 port map( I => n10519, Z => n25829);
   U3190 : BUF_X4 port map( I => n12477, Z => n26355);
   U14179 : AOI22_X2 port map( A1 => n10118, A2 => n27734, B1 => n14676, B2 => 
                           n9917, ZN => n10117);
   U13467 : BUF_X2 port map( I => n14554, Z => n9087);
   U206 : INV_X2 port map( I => n20155, ZN => n958);
   U12968 : OR2_X1 port map( A1 => n1892, A2 => n14658, Z => n3935);
   U5263 : INV_X2 port map( I => n25508, ZN => n17826);
   U1327 : INV_X4 port map( I => n7481, ZN => n1211);
   U3184 : AOI22_X2 port map( A1 => n20125, A2 => n9264, B1 => n26355, B2 => 
                           n8265, ZN => n19971);
   U3740 : INV_X2 port map( I => n10578, ZN => n20866);
   U21250 : BUF_X4 port map( I => n7379, Z => n26410);
   U895 : INV_X2 port map( I => n3537, ZN => n7517);
   U8791 : NAND2_X2 port map( A1 => n21932, A2 => n25254, ZN => n5202);
   U4708 : INV_X4 port map( I => n19004, ZN => n13563);
   U7565 : OAI21_X2 port map( A1 => n5704, A2 => n14683, B => n9508, ZN => 
                           n3373);
   U5333 : OAI22_X2 port map( A1 => n16186, A2 => n13533, B1 => n13142, B2 => 
                           n16185, ZN => n8970);
   U4917 : INV_X2 port map( I => n19630, ZN => n1122);
   U18121 : NOR2_X1 port map( A1 => n26035, A2 => n10930, ZN => n21826);
   U15002 : INV_X2 port map( I => n14961, ZN => n21160);
   U18254 : INV_X2 port map( I => n10097, ZN => n26317);
   U7612 : INV_X2 port map( I => n5704, ZN => n5749);
   U5251 : OAI21_X2 port map( A1 => n6481, A2 => n9690, B => n17822, ZN => 
                           n13586);
   U10365 : NOR2_X2 port map( A1 => n703, A2 => n132, ZN => n14778);
   U3094 : NAND2_X2 port map( A1 => n19731, A2 => n19846, ZN => n26272);
   U12019 : INV_X2 port map( I => n19919, ZN => n23821);
   U2216 : INV_X4 port map( I => n15453, ZN => n20263);
   U1051 : INV_X4 port map( I => n17515, ZN => n24323);
   U2758 : NAND2_X2 port map( A1 => n11514, A2 => n27146, ZN => n3235);
   U70 : NOR2_X2 port map( A1 => n3362, A2 => n21135, ZN => n110);
   U8779 : OAI21_X2 port map( A1 => n15178, A2 => n4342, B => n20144, ZN => 
                           n4341);
   U3113 : NOR2_X2 port map( A1 => n20071, A2 => n22735, ZN => n4342);
   U3393 : BUF_X4 port map( I => n16184, Z => n21787);
   U13024 : NAND2_X1 port map( A1 => n1125, A2 => n27905, ZN => n19168);
   U11326 : INV_X2 port map( I => n6063, ZN => n15812);
   U3545 : INV_X4 port map( I => n11223, ZN => n1055);
   U2355 : INV_X2 port map( I => n8459, ZN => n24151);
   U4137 : BUF_X4 port map( I => n16419, Z => n703);
   U4928 : NAND2_X2 port map( A1 => n4735, A2 => n19138, ZN => n19135);
   U1952 : OAI21_X2 port map( A1 => n19599, A2 => n777, B => n775, ZN => n9441)
                           ;
   U5329 : NOR2_X2 port map( A1 => n16240, A2 => n16239, ZN => n9769);
   U6792 : INV_X1 port map( I => n15831, ZN => n15770);
   U7277 : NAND2_X2 port map( A1 => n1154, A2 => n994, ZN => n14959);
   U14995 : NAND3_X2 port map( A1 => n994, A2 => n4471, A3 => n27813, ZN => 
                           n12817);
   U263 : NAND2_X2 port map( A1 => n6646, A2 => n23558, ZN => n25048);
   U4509 : INV_X2 port map( I => n10064, ZN => n14557);
   U8012 : OAI21_X2 port map( A1 => n24614, A2 => n16701, B => n16469, ZN => 
                           n4426);
   U9338 : NAND3_X2 port map( A1 => n728, A2 => n25724, A3 => n27550, ZN => 
                           n3119);
   U13403 : OAI21_X2 port map( A1 => n14519, A2 => n1271, B => n12010, ZN => 
                           n15991);
   U610 : NOR2_X2 port map( A1 => n9628, A2 => n9627, ZN => n25491);
   U2020 : BUF_X2 port map( I => n18452, Z => n7165);
   U1824 : BUF_X4 port map( I => n11100, Z => n6523);
   U1449 : NAND3_X2 port map( A1 => n12937, A2 => n22172, A3 => n22171, ZN => 
                           n23553);
   U4130 : INV_X2 port map( I => n26298, ZN => n26024);
   U4833 : NAND2_X2 port map( A1 => n14569, A2 => n14883, ZN => n22239);
   U16775 : INV_X4 port map( I => n7553, ZN => n17984);
   U8359 : BUF_X2 port map( I => Key(119), Z => n21422);
   U15532 : CLKBUF_X4 port map( I => n14326, Z => n25657);
   U143 : INV_X2 port map( I => n12055, ZN => n3481);
   U10728 : OR2_X1 port map( A1 => n6859, A2 => n14632, Z => n16401);
   U13992 : INV_X2 port map( I => n9642, ZN => n13905);
   U9661 : BUF_X2 port map( I => n18549, Z => n14594);
   U598 : NAND3_X2 port map( A1 => n13806, A2 => n13805, A3 => n7358, ZN => 
                           n6847);
   U16867 : INV_X2 port map( I => n8408, ZN => n16063);
   U4422 : NAND2_X2 port map( A1 => n18731, A2 => n24937, ZN => n18732);
   U4415 : NOR2_X2 port map( A1 => n204, A2 => n6529, ZN => n10357);
   U1002 : NAND2_X1 port map( A1 => n23338, A2 => n17558, ZN => n3034);
   U7447 : NOR2_X1 port map( A1 => n816, A2 => n21767, ZN => n6351);
   U15662 : BUF_X2 port map( I => n13274, Z => n23309);
   U469 : INV_X4 port map( I => n7030, ZN => n994);
   U12766 : INV_X2 port map( I => n20102, ZN => n10808);
   U6258 : NOR2_X2 port map( A1 => n8007, A2 => n27704, ZN => n19104);
   U5387 : INV_X2 port map( I => n15686, ZN => n1262);
   U1538 : NAND2_X2 port map( A1 => n3981, A2 => n16663, ZN => n16665);
   U5173 : INV_X2 port map( I => n172, ZN => n26071);
   U1484 : NOR2_X2 port map( A1 => n431, A2 => n3330, ZN => n24792);
   U16027 : INV_X2 port map( I => n5305, ZN => n25738);
   U5849 : AOI21_X2 port map( A1 => n18526, A2 => n12980, B => n7084, ZN => 
                           n14019);
   U2119 : NAND3_X2 port map( A1 => n14835, A2 => n6699, A3 => n14833, ZN => 
                           n12432);
   U6083 : OAI21_X2 port map( A1 => n4742, A2 => n21024, B => n708, ZN => 
                           n11140);
   U4230 : NAND2_X1 port map( A1 => n23630, A2 => n23628, ZN => n16003);
   U1988 : NOR2_X2 port map( A1 => n19968, A2 => n3223, ZN => n6501);
   U8656 : AOI21_X2 port map( A1 => n5704, A2 => n14683, B => n737, ZN => 
                           n24914);
   U341 : INV_X4 port map( I => n26624, ZN => n19802);
   U1843 : INV_X2 port map( I => n17559, ZN => n13607);
   U3483 : CLKBUF_X8 port map( I => n679, Z => n2891);
   U5408 : INV_X4 port map( I => n7486, ZN => n797);
   U13471 : OR2_X1 port map( A1 => n18661, A2 => n14745, Z => n18662);
   U12287 : NOR2_X2 port map( A1 => n2670, A2 => n4738, ZN => n25517);
   U17295 : INV_X2 port map( I => n9370, ZN => n17418);
   U900 : NOR2_X2 port map( A1 => n14777, A2 => n22197, ZN => n17506);
   U687 : NAND2_X2 port map( A1 => n8330, A2 => n12393, ZN => n22903);
   U9352 : INV_X4 port map( I => n797, ZN => n22371);
   U4711 : INV_X2 port map( I => n20316, ZN => n744);
   U15191 : NAND3_X1 port map( A1 => n23226, A2 => n21392, A3 => n23225, ZN => 
                           n21393);
   U13128 : BUF_X4 port map( I => n3932, Z => n1558);
   U15927 : INV_X2 port map( I => n14981, ZN => n18355);
   U4238 : NOR2_X1 port map( A1 => n1994, A2 => n22908, ZN => n23349);
   U7763 : INV_X4 port map( I => n17957, ZN => n17785);
   U4949 : OAI21_X1 port map( A1 => n12955, A2 => n18583, B => n12953, ZN => 
                           n12579);
   U9250 : NOR2_X2 port map( A1 => n18796, A2 => n18795, ZN => n3386);
   U1803 : NAND3_X2 port map( A1 => n12175, A2 => n9910, A3 => n13169, ZN => 
                           n22036);
   U879 : INV_X2 port map( I => n6763, ZN => n6898);
   U3295 : NAND2_X2 port map( A1 => n14804, A2 => n9304, ZN => n23953);
   U3945 : OR2_X1 port map( A1 => n1325, A2 => n12189, Z => n24105);
   U1508 : NAND2_X2 port map( A1 => n16665, A2 => n25249, ZN => n26043);
   U1062 : NAND2_X2 port map( A1 => n18585, A2 => n18586, ZN => n18584);
   U18096 : NOR2_X2 port map( A1 => n1001, A2 => n23624, ZN => n11414);
   U21013 : NAND2_X2 port map( A1 => n778, A2 => n28240, ZN => n18860);
   U6021 : OAI21_X2 port map( A1 => n20182, A2 => n20239, B => n13995, ZN => 
                           n11210);
   U1026 : INV_X4 port map( I => n1882, ZN => n14804);
   U13159 : BUF_X4 port map( I => n3982, Z => n3981);
   U17266 : NAND2_X2 port map( A1 => n23592, A2 => n8032, ZN => n23591);
   U13223 : INV_X2 port map( I => n20852, ZN => n7956);
   U12830 : NAND2_X2 port map( A1 => n797, A2 => n24643, ZN => n16213);
   U2965 : OAI22_X2 port map( A1 => n4108, A2 => n857, B1 => n3870, B2 => n7942
                           , ZN => n1358);
   U2118 : OAI22_X2 port map( A1 => n3110, A2 => n17303, B1 => n17307, B2 => 
                           n2963, ZN => n23815);
   U13248 : NOR2_X2 port map( A1 => n1882, A2 => n27177, ZN => n9804);
   U9643 : BUF_X2 port map( I => n15362, Z => n7769);
   U18303 : NAND2_X2 port map( A1 => n11959, A2 => n9040, ZN => n11958);
   U12884 : OAI22_X2 port map( A1 => n2952, A2 => n28295, B1 => n22519, B2 => 
                           n25679, ZN => n2388);
   U2657 : NAND2_X2 port map( A1 => n9691, A2 => n11968, ZN => n17638);
   U18631 : NAND2_X2 port map( A1 => n10823, A2 => n17957, ZN => n17376);
   U4045 : NAND2_X2 port map( A1 => n23953, A2 => n23952, ZN => n22897);
   U13250 : AOI21_X2 port map( A1 => n12964, A2 => n27177, B => n21778, ZN => 
                           n23952);
   U21585 : NOR2_X2 port map( A1 => n11447, A2 => n15751, ZN => n24447);
   U2386 : INV_X2 port map( I => n7354, ZN => n15724);
   U1647 : OAI21_X2 port map( A1 => n9629, A2 => n8033, B => n26061, ZN => 
                           n8035);
   U16702 : NAND2_X2 port map( A1 => n18949, A2 => n27569, ZN => n8095);
   U14264 : INV_X1 port map( I => n2284, ZN => n24443);
   U13923 : OAI22_X2 port map( A1 => n18587, A2 => n18586, B1 => n14494, B2 => 
                           n1013, ZN => n7171);
   U1663 : NOR2_X2 port map( A1 => n19951, A2 => n19952, ZN => n422);
   U9093 : AOI22_X2 port map( A1 => n19717, A2 => n19716, B1 => n19827, B2 => 
                           n19715, ZN => n19718);
   U6363 : INV_X1 port map( I => n19684, ZN => n19955);
   U256 : NOR3_X2 port map( A1 => n23676, A2 => n20318, A3 => n14104, ZN => 
                           n8478);
   U2382 : NOR2_X2 port map( A1 => n10963, A2 => n7122, ZN => n12250);
   U418 : NAND3_X2 port map( A1 => n5189, A2 => n19005, A3 => n18956, ZN => 
                           n11028);
   U17826 : NAND2_X2 port map( A1 => n8326, A2 => n19689, ZN => n10957);
   U3117 : OAI21_X2 port map( A1 => n2316, A2 => n2315, B => n10498, ZN => 
                           n2314);
   U1624 : INV_X4 port map( I => n5402, ZN => n17959);
   U3479 : CLKBUF_X4 port map( I => n18146, Z => n18583);
   U1544 : BUF_X4 port map( I => n14260, Z => n216);
   U5794 : INV_X2 port map( I => n19073, ZN => n15434);
   U5930 : NOR3_X1 port map( A1 => n3959, A2 => n950, A3 => n20931, ZN => n4081
                           );
   U4722 : OAI21_X2 port map( A1 => n10746, A2 => n11704, B => n11703, ZN => 
                           n25043);
   U7812 : OAI21_X2 port map( A1 => n1952, A2 => n1951, B => n1950, ZN => n1949
                           );
   U2428 : AOI21_X2 port map( A1 => n1158, A2 => n447, B => n2733, ZN => n8711)
                           ;
   U1078 : NOR2_X2 port map( A1 => n18785, A2 => n18629, ZN => n12324);
   U13621 : NAND3_X2 port map( A1 => n12732, A2 => n5192, A3 => n25051, ZN => 
                           n11907);
   U9969 : OAI21_X2 port map( A1 => n3175, A2 => n17022, B => n17021, ZN => 
                           n13956);
   U11534 : NOR2_X1 port map( A1 => n24610, A2 => n18630, ZN => n7789);
   U17090 : INV_X2 port map( I => n17318, ZN => n23556);
   U6715 : INV_X4 port map( I => n8882, ZN => n25688);
   U19946 : NOR2_X2 port map( A1 => n24442, A2 => n14271, ZN => n19225);
   U3672 : INV_X4 port map( I => n21024, ZN => n1087);
   U3211 : OAI21_X2 port map( A1 => n744, A2 => n13754, B => n14104, ZN => 
                           n8480);
   U10570 : INV_X2 port map( I => n6428, ZN => n3572);
   U3991 : INV_X1 port map( I => n13467, ZN => n18608);
   U2440 : NAND2_X2 port map( A1 => n17785, A2 => n5449, ZN => n15407);
   U18666 : INV_X4 port map( I => n10875, ZN => n14900);
   U20752 : OAI21_X2 port map( A1 => n23915, A2 => n1212, B => n27852, ZN => 
                           n17257);
   U14256 : NAND2_X2 port map( A1 => n4536, A2 => n25971, ZN => n6258);
   U1603 : NAND2_X2 port map( A1 => n16610, A2 => n9978, ZN => n16507);
   U14558 : NAND2_X2 port map( A1 => n23857, A2 => n7895, ZN => n7894);
   U748 : INV_X2 port map( I => n10923, ZN => n17569);
   U8146 : NAND2_X1 port map( A1 => n1930, A2 => n12918, ZN => n1929);
   U593 : OAI21_X2 port map( A1 => n27756, A2 => n17974, B => n116, ZN => n5236
                           );
   U3098 : BUF_X2 port map( I => n10638, Z => n14883);
   U7301 : NOR2_X2 port map( A1 => n19952, A2 => n14651, ZN => n19715);
   U14876 : NOR2_X2 port map( A1 => n3229, A2 => n5574, ZN => n25571);
   U11100 : INV_X2 port map( I => n12648, ZN => n13354);
   U1301 : NAND2_X2 port map( A1 => n1200, A2 => n4318, ZN => n13806);
   U419 : NAND2_X2 port map( A1 => n8515, A2 => n8514, ZN => n14239);
   U1543 : NAND2_X2 port map( A1 => n216, A2 => n21933, ZN => n22209);
   U9050 : INV_X1 port map( I => n18645, ZN => n25355);
   U12926 : OAI22_X2 port map( A1 => n19833, A2 => n28207, B1 => n19832, B2 => 
                           n19906, ZN => n13649);
   U17117 : INV_X2 port map( I => n12595, ZN => n8986);
   U3233 : NOR2_X1 port map( A1 => n22459, A2 => n1014, ZN => n22458);
   U6778 : INV_X2 port map( I => n16069, ZN => n16275);
   U14337 : INV_X4 port map( I => n26654, ZN => n19906);
   U10379 : NOR2_X2 port map( A1 => n13220, A2 => n9793, ZN => n13838);
   U1605 : NOR2_X2 port map( A1 => n1256, A2 => n10597, ZN => n12318);
   U273 : INV_X2 port map( I => n19798, ZN => n19754);
   U9472 : NOR2_X2 port map( A1 => n4961, A2 => n4960, ZN => n2257);
   U7777 : NOR2_X2 port map( A1 => n11591, A2 => n11590, ZN => n11589);
   U9804 : NOR2_X1 port map( A1 => n2751, A2 => n17766, ZN => n2318);
   U8992 : AOI21_X2 port map( A1 => n17620, A2 => n17621, B => n17619, ZN => 
                           n25476);
   U415 : INV_X2 port map( I => n12980, ZN => n18525);
   U7687 : AOI22_X2 port map( A1 => n17616, A2 => n17618, B1 => n17615, B2 => 
                           n7614, ZN => n8708);
   U17496 : INV_X2 port map( I => n9916, ZN => n21324);
   U8561 : OAI22_X2 port map( A1 => n11980, A2 => n11978, B1 => n11977, B2 => 
                           n23225, ZN => n11976);
   U5645 : OAI21_X2 port map( A1 => n13421, A2 => n17898, B => n7120, ZN => 
                           n17902);
   U4484 : INV_X4 port map( I => n15425, ZN => n17381);
   U14860 : NAND2_X2 port map( A1 => n11257, A2 => n24027, ZN => n6776);
   U197 : INV_X2 port map( I => n20291, ZN => n20196);
   U4187 : BUF_X4 port map( I => n15425, Z => n24406);
   U18178 : OAI21_X2 port map( A1 => n20881, A2 => n950, B => n20931, ZN => 
                           n13584);
   U19328 : NAND2_X2 port map( A1 => n26191, A2 => n13070, ZN => n7774);
   U2263 : OAI21_X1 port map( A1 => n12583, A2 => n10617, B => n13401, ZN => 
                           n18890);
   U6046 : INV_X1 port map( I => n21428, ZN => n23799);
   U2261 : NOR2_X2 port map( A1 => n7820, A2 => n7293, ZN => n7819);
   U4393 : OAI21_X2 port map( A1 => n24642, A2 => n25960, B => n20270, ZN => 
                           n9957);
   U15518 : INV_X2 port map( I => n17457, ZN => n6294);
   U591 : NAND2_X2 port map( A1 => n17862, A2 => n727, ZN => n14716);
   U12958 : NOR2_X2 port map( A1 => n15434, A2 => n15429, ZN => n23752);
   U16440 : INV_X4 port map( I => n7561, ZN => n9057);
   U2364 : NOR2_X2 port map( A1 => n17529, A2 => n9358, ZN => n9696);
   U980 : OAI22_X2 port map( A1 => n25147, A2 => n14498, B1 => n7212, B2 => 
                           n9041, ZN => n3495);
   U8418 : NOR2_X2 port map( A1 => n26272, A2 => n26271, ZN => n24972);
   U13142 : BUF_X4 port map( I => n12947, Z => n10221);
   U716 : INV_X4 port map( I => n15560, ZN => n964);
   U3640 : OR2_X1 port map( A1 => n16524, A2 => n16525, Z => n2692);
   U219 : INV_X4 port map( I => n5415, ZN => n20317);
   U7835 : NAND3_X2 port map( A1 => n10897, A2 => n17408, A3 => n897, ZN => 
                           n3675);
   U2610 : INV_X2 port map( I => n8031, ZN => n16329);
   U1744 : CLKBUF_X4 port map( I => n20057, Z => n19);
   U18467 : NAND3_X1 port map( A1 => n27822, A2 => n12082, A3 => n12179, ZN => 
                           n20994);
   U4813 : INV_X2 port map( I => n19124, ZN => n986);
   U9937 : NAND2_X2 port map( A1 => n10416, A2 => n790, ZN => n10415);
   U10056 : NAND2_X2 port map( A1 => n26335, A2 => n4675, ZN => n25812);
   U4984 : NOR2_X1 port map( A1 => n9329, A2 => n1411, ZN => n3814);
   U6655 : BUF_X4 port map( I => n16699, Z => n22061);
   U131 : INV_X4 port map( I => n6375, ZN => n10610);
   U4883 : NAND2_X1 port map( A1 => n22266, A2 => n15220, ZN => n10775);
   U6233 : AOI22_X2 port map( A1 => n23268, A2 => n13183, B1 => n18956, B2 => 
                           n757, ZN => n9326);
   U9435 : INV_X2 port map( I => n6908, ZN => n6907);
   U4779 : OAI21_X2 port map( A1 => n10039, A2 => n5645, B => n18685, ZN => 
                           n25956);
   U5254 : OAI21_X2 port map( A1 => n26704, A2 => n8784, B => n24391, ZN => 
                           n8013);
   U12848 : AND3_X2 port map( A1 => n7940, A2 => n21495, A3 => n21500, Z => 
                           n13321);
   U10419 : INV_X2 port map( I => n1545, ZN => n1544);
   U2708 : OAI21_X2 port map( A1 => n836, A2 => n11223, B => n16063, ZN => 
                           n1545);
   U2553 : AOI22_X2 port map( A1 => n14819, A2 => n13532, B1 => n3106, B2 => 
                           n1997, ZN => n1996);
   U17016 : INV_X2 port map( I => n8724, ZN => n17460);
   U1740 : INV_X1 port map( I => n9598, ZN => n26122);
   U754 : INV_X4 port map( I => n17534, ZN => n764);
   U9208 : NOR2_X2 port map( A1 => n9351, A2 => n9353, ZN => n9350);
   U14932 : INV_X4 port map( I => n17301, ZN => n9481);
   U15356 : AOI21_X2 port map( A1 => n11808, A2 => n17803, B => n25640, ZN => 
                           n15563);
   U13920 : INV_X2 port map( I => n4344, ZN => n6681);
   U3100 : INV_X4 port map( I => n17926, ZN => n17928);
   U10702 : BUF_X2 port map( I => Key(149), Z => n21607);
   U1103 : CLKBUF_X4 port map( I => n10904, Z => n26228);
   U20118 : INV_X2 port map( I => n14673, ZN => n17497);
   U4539 : INV_X2 port map( I => n20817, ZN => n732);
   U4532 : NAND3_X2 port map( A1 => n10554, A2 => n708, A3 => n27689, ZN => 
                           n21028);
   U2475 : NOR2_X2 port map( A1 => n2481, A2 => n9917, ZN => n10118);
   U5515 : NAND2_X2 port map( A1 => n19800, A2 => n19801, ZN => n9660);
   U8150 : OAI21_X1 port map( A1 => n13942, A2 => n12338, B => n757, ZN => 
                           n23059);
   U2392 : INV_X4 port map( I => n10556, ZN => n14128);
   U2002 : NOR3_X2 port map( A1 => n21540, A2 => n21669, A3 => n21666, ZN => 
                           n15175);
   U2415 : INV_X4 port map( I => n11627, ZN => n22732);
   U2486 : INV_X2 port map( I => n16063, ZN => n22798);
   U9590 : OAI21_X1 port map( A1 => n9248, A2 => n15674, B => n18611, ZN => 
                           n18615);
   U6962 : NOR2_X2 port map( A1 => n27689, A2 => n7421, ZN => n20541);
   U2557 : BUF_X4 port map( I => n12974, Z => n12647);
   U15633 : NAND2_X1 port map( A1 => n23306, A2 => n20314, ZN => n7636);
   U16971 : NAND2_X2 port map( A1 => n8645, A2 => n13812, ZN => n18965);
   U1562 : INV_X2 port map( I => n14501, ZN => n18629);
   U6365 : INV_X2 port map( I => n24092, ZN => n1006);
   U6816 : INV_X4 port map( I => n24581, ZN => n16027);
   U14108 : INV_X4 port map( I => n16700, ZN => n16469);
   U4620 : INV_X4 port map( I => n21842, ZN => n739);
   U4671 : BUF_X2 port map( I => n7533, Z => n25664);
   U5853 : NOR2_X1 port map( A1 => n1604, A2 => n1603, ZN => n1602);
   U3622 : BUF_X4 port map( I => n10543, Z => n1256);
   U7496 : NOR2_X1 port map( A1 => n27653, A2 => n9429, ZN => n24786);
   U1217 : OAI21_X2 port map( A1 => n7617, A2 => n17680, B => n27100, ZN => 
                           n7616);
   U9182 : NOR2_X2 port map( A1 => n27699, A2 => n7614, ZN => n7617);
   U14420 : INV_X4 port map( I => n20129, ZN => n23676);
   U10278 : NOR2_X2 port map( A1 => n21830, A2 => n11547, ZN => n11546);
   U1995 : OAI22_X2 port map( A1 => n10761, A2 => n7251, B1 => n27557, B2 => 
                           n19821, ZN => n5100);
   U4433 : INV_X2 port map( I => n16610, ZN => n1792);
   U2983 : INV_X2 port map( I => n25679, ZN => n17618);
   U556 : INV_X1 port map( I => n25769, ZN => n18531);
   U7806 : NAND2_X2 port map( A1 => n5679, A2 => n24214, ZN => n5678);
   U4164 : NAND2_X2 port map( A1 => n24613, A2 => n17342, ZN => n5679);
   U3946 : NOR2_X2 port map( A1 => n22119, A2 => n22118, ZN => n22185);
   U780 : INV_X1 port map( I => n13411, ZN => n15592);
   U1152 : NOR2_X2 port map( A1 => n16695, A2 => n24167, ZN => n5850);
   U10023 : OR2_X1 port map( A1 => n26264, A2 => n2068, Z => n26483);
   U3428 : AND2_X2 port map( A1 => n12062, A2 => n12064, Z => n22821);
   U7479 : NOR2_X2 port map( A1 => n15599, A2 => n1169, ZN => n15598);
   U4855 : OR2_X2 port map( A1 => n6489, A2 => n19154, Z => n8485);
   U2313 : BUF_X4 port map( I => n9887, Z => n26129);
   U311 : NAND2_X2 port map( A1 => n21759, A2 => n27414, ZN => n20248);
   U5593 : NOR2_X2 port map( A1 => n47, A2 => n23197, ZN => n4101);
   U3410 : NOR2_X2 port map( A1 => n9538, A2 => n19140, ZN => n13171);
   U8653 : NAND2_X2 port map( A1 => n3067, A2 => n26338, ZN => n22309);
   U4261 : BUF_X2 port map( I => n21545, Z => n10532);
   U4329 : NAND2_X2 port map( A1 => n14442, A2 => n22801, ZN => n8696);
   U3901 : OAI22_X2 port map( A1 => n13659, A2 => n25984, B1 => n14222, B2 => 
                           n25514, ZN => n4171);
   U7511 : NAND2_X2 port map( A1 => n1168, A2 => n8022, ZN => n4392);
   U11975 : NAND2_X2 port map( A1 => n23926, A2 => n17480, ZN => n13355);
   U4348 : INV_X2 port map( I => n21292, ZN => n15375);
   U20314 : NOR2_X2 port map( A1 => n11196, A2 => n15416, ZN => n15415);
   U8238 : NAND3_X1 port map( A1 => n23104, A2 => n10440, A3 => n9393, ZN => 
                           n10439);
   U1682 : NAND3_X2 port map( A1 => n10665, A2 => n14222, A3 => n21765, ZN => 
                           n15300);
   U17834 : INV_X2 port map( I => n21376, ZN => n15130);
   U2552 : NOR2_X2 port map( A1 => n13532, A2 => n13184, ZN => n18406);
   U2786 : OAI21_X2 port map( A1 => n23870, A2 => n5806, B => n20637, ZN => 
                           n2624);
   U7183 : NOR2_X2 port map( A1 => n27043, A2 => n25514, ZN => n24756);
   U4699 : AOI22_X2 port map( A1 => n23064, A2 => n23063, B1 => n13264, B2 => 
                           n17783, ZN => n6848);
   U3660 : OAI21_X2 port map( A1 => n24632, A2 => n15489, B => n22748, ZN => 
                           n6855);
   U5054 : OR3_X2 port map( A1 => n17418, A2 => n14990, A3 => n3091, Z => 
                           n11569);
   U16010 : NAND2_X2 port map( A1 => n20213, A2 => n12946, ZN => n10224);
   U20624 : NAND2_X2 port map( A1 => n476, A2 => n8442, ZN => n24123);
   U6996 : OAI21_X2 port map( A1 => n21097, A2 => n21096, B => n28139, ZN => 
                           n7263);
   U13777 : NAND2_X2 port map( A1 => n10415, A2 => n13355, ZN => n22907);
   U10881 : INV_X2 port map( I => n26705, ZN => n25155);
   U7007 : BUF_X2 port map( I => n631, Z => n5489);
   U1724 : INV_X4 port map( I => n4705, ZN => n989);
   U13949 : NOR2_X1 port map( A1 => n9181, A2 => n23287, ZN => n7261);
   U1549 : NAND2_X2 port map( A1 => n24644, A2 => n404, ZN => n21833);
   U1665 : INV_X1 port map( I => n2264, ZN => n1402);
   U4993 : NOR2_X2 port map( A1 => n28295, A2 => n4914, ZN => n7615);
   U4560 : NAND3_X2 port map( A1 => n13771, A2 => n10293, A3 => n27557, ZN => 
                           n9265);
   U21188 : INV_X2 port map( I => n24219, ZN => n19937);
   U19143 : BUF_X2 port map( I => n24127, Z => n26437);
   U17732 : NAND2_X2 port map( A1 => n28091, A2 => n1108, ZN => n20307);
   U15284 : INV_X2 port map( I => n5862, ZN => n8237);
   U10208 : NAND3_X1 port map( A1 => n7114, A2 => n16587, A3 => n7112, ZN => 
                           n11548);
   U5214 : BUF_X2 port map( I => n14766, Z => n26244);
   U8008 : OAI21_X2 port map( A1 => n13261, A2 => n4630, B => n12881, ZN => 
                           n12328);
   U2357 : INV_X4 port map( I => n16813, ZN => n15029);
   U929 : INV_X4 port map( I => n16283, ZN => n13533);
   U4305 : BUF_X4 port map( I => n12694, Z => n24215);
   U11586 : NOR2_X2 port map( A1 => n4597, A2 => n16597, ZN => n11447);
   U2445 : NAND2_X2 port map( A1 => n6904, A2 => n14578, ZN => n2101);
   U2812 : INV_X2 port map( I => n14724, ZN => n24841);
   U5114 : BUF_X4 port map( I => n6853, Z => n25013);
   U1989 : NOR2_X2 port map( A1 => n21097, A2 => n14341, ZN => n8278);
   U248 : NOR2_X2 port map( A1 => n4438, A2 => n4437, ZN => n4436);
   U10935 : OR2_X2 port map( A1 => n25357, A2 => n8439, Z => n8004);
   U3952 : BUF_X2 port map( I => n7057, Z => n1366);
   U13837 : INV_X2 port map( I => n14117, ZN => n17495);
   U22047 : NAND2_X2 port map( A1 => n12244, A2 => n18624, ZN => n26598);
   U7161 : INV_X2 port map( I => n16602, ZN => n1054);
   U5911 : NOR2_X2 port map( A1 => n3317, A2 => n14304, ZN => n21837);
   U8411 : NAND2_X2 port map( A1 => n6150, A2 => n6149, ZN => n5412);
   U17053 : NAND2_X1 port map( A1 => n6584, A2 => n15028, ZN => n25908);
   U2582 : NOR2_X1 port map( A1 => n18383, A2 => n11186, ZN => n11185);
   U1136 : NOR2_X2 port map( A1 => n145, A2 => n25698, ZN => n16412);
   U16482 : INV_X2 port map( I => n25806, ZN => n18487);
   U8867 : NOR2_X2 port map( A1 => n28419, A2 => n15544, ZN => n9010);
   U10000 : AOI21_X2 port map( A1 => n6525, A2 => n20030, B => n25084, ZN => 
                           n22701);
   U19653 : OAI21_X2 port map( A1 => n826, A2 => n14885, B => n22594, ZN => 
                           n8974);
   U1956 : NAND2_X1 port map( A1 => n24904, A2 => n12625, ZN => n21514);
   U8362 : BUF_X2 port map( I => Key(7), Z => n14560);
   U19137 : NAND2_X2 port map( A1 => n3276, A2 => n11982, ZN => n13919);
   U1175 : INV_X4 port map( I => n18432, ZN => n18666);
   U3836 : BUF_X2 port map( I => n19238, Z => n23691);
   U522 : AOI22_X2 port map( A1 => n10080, A2 => n864, B1 => n26625, B2 => 
                           n19746, ZN => n23167);
   U10239 : AOI22_X2 port map( A1 => n552, A2 => n26435, B1 => n21589, B2 => 
                           n8751, ZN => n25549);
   U16402 : BUF_X4 port map( I => n766, Z => n25796);
   U6974 : OAI22_X2 port map( A1 => n20643, A2 => n10512, B1 => n21714, B2 => 
                           n20644, ZN => n10515);
   U2846 : OAI21_X2 port map( A1 => n19647, A2 => n10739, B => n27204, ZN => 
                           n22671);
   U5922 : BUF_X4 port map( I => n19913, Z => n23857);
   U6450 : OAI21_X1 port map( A1 => n24633, A2 => n19017, B => n24745, ZN => 
                           n18975);
   U6231 : BUF_X4 port map( I => n3914, Z => n404);
   U8022 : AOI21_X2 port map( A1 => n9139, A2 => n26039, B => n23439, ZN => 
                           n7877);
   U5963 : AOI21_X2 port map( A1 => n8621, A2 => n23857, B => n24545, ZN => 
                           n15231);
   U760 : NOR2_X2 port map( A1 => n2356, A2 => n1658, ZN => n25245);
   U21167 : NOR3_X2 port map( A1 => n7919, A2 => n25368, A3 => n24190, ZN => 
                           n1816);
   U2977 : NOR2_X2 port map( A1 => n4914, A2 => n25679, ZN => n17680);
   U11969 : OAI21_X2 port map( A1 => n2790, A2 => n5677, B => n2527, ZN => 
                           n5676);
   U5893 : NAND2_X2 port map( A1 => n19748, A2 => n669, ZN => n2034);
   U7216 : NAND2_X2 port map( A1 => n6593, A2 => n10941, ZN => n13341);
   U510 : OAI21_X2 port map( A1 => n10654, A2 => n14516, B => n19847, ZN => 
                           n3212);
   U4856 : BUF_X2 port map( I => n18575, Z => n14510);
   U2396 : INV_X2 port map( I => n21029, ZN => n20890);
   U13353 : INV_X2 port map( I => n8290, ZN => n8716);
   U721 : OR2_X2 port map( A1 => n10255, A2 => n19593, Z => n19849);
   U8855 : NOR2_X2 port map( A1 => n20223, A2 => n13294, ZN => n15744);
   U18634 : OAI22_X1 port map( A1 => n3431, A2 => n13962, B1 => n5634, B2 => 
                           n24579, ZN => n26401);
   U4991 : INV_X2 port map( I => n6211, ZN => n8621);
   U2899 : BUF_X2 port map( I => n19649, Z => n19915);
   U2863 : OR2_X1 port map( A1 => n10251, A2 => n649, Z => n14096);
   U1498 : NAND2_X2 port map( A1 => n24900, A2 => n24899, ZN => n4493);
   U9172 : BUF_X2 port map( I => n19651, Z => n11988);
   U5494 : OR2_X2 port map( A1 => n6018, A2 => n17855, Z => n21905);
   U11091 : OR2_X2 port map( A1 => n6575, A2 => n25385, Z => n12748);
   U1734 : INV_X4 port map( I => n26434, ZN => n12678);
   U9044 : OAI21_X2 port map( A1 => n14241, A2 => n11901, B => n19801, ZN => 
                           n7196);
   U18563 : NOR2_X1 port map( A1 => n16514, A2 => n23749, ZN => n26103);
   U1342 : OAI21_X2 port map( A1 => n14724, A2 => n2815, B => n3018, ZN => 
                           n23497);
   U1765 : NOR2_X2 port map( A1 => n24076, A2 => n24825, ZN => n17596);
   U1222 : NOR3_X2 port map( A1 => n17727, A2 => n14230, A3 => n23245, ZN => 
                           n24825);
   U4132 : INV_X4 port map( I => n17989, ZN => n21791);
   U3120 : BUF_X4 port map( I => n15806, Z => n6315);
   U3913 : BUF_X4 port map( I => n23871, Z => n427);
   U939 : INV_X2 port map( I => n24524, ZN => n26097);
   U3026 : NAND2_X2 port map( A1 => n6820, A2 => n15461, ZN => n12014);
   U7428 : NOR2_X2 port map( A1 => n10632, A2 => n24783, ZN => n11082);
   U15056 : NAND3_X2 port map( A1 => n9139, A2 => n16249, A3 => n16455, ZN => 
                           n16252);
   U13458 : NAND3_X2 port map( A1 => n745, A2 => n26252, A3 => n27679, ZN => 
                           n5173);
   U9996 : OAI21_X2 port map( A1 => n10694, A2 => n10954, B => n1032, ZN => 
                           n10953);
   U17479 : AOI21_X2 port map( A1 => n5055, A2 => n11983, B => n26822, ZN => 
                           n13489);
   U3063 : INV_X2 port map( I => n4644, ZN => n1046);
   U1502 : NOR2_X2 port map( A1 => n19758, A2 => n19752, ZN => n6279);
   U11025 : NOR2_X2 port map( A1 => n9645, A2 => n8073, ZN => n22563);
   U6505 : INV_X1 port map( I => n17927, ZN => n1212);
   U4377 : NAND2_X1 port map( A1 => n20116, A2 => n25518, ZN => n20118);
   U229 : AND2_X2 port map( A1 => n8098, A2 => n8099, Z => n955);
   U21325 : INV_X2 port map( I => n20783, ZN => n20633);
   U5021 : NAND2_X2 port map( A1 => n28539, A2 => n14762, ZN => n17467);
   U3355 : NOR2_X1 port map( A1 => n11095, A2 => n4939, ZN => n6496);
   U2976 : OAI21_X2 port map( A1 => n23772, A2 => n5990, B => n27044, ZN => 
                           n18899);
   U8821 : NAND2_X1 port map( A1 => n20295, A2 => n15279, ZN => n11542);
   U20959 : NAND2_X2 port map( A1 => n13584, A2 => n20938, ZN => n24186);
   U2247 : NOR2_X2 port map( A1 => n20852, A2 => n15724, ZN => n20887);
   U17344 : NAND2_X2 port map( A1 => n17174, A2 => n12236, ZN => n24006);
   U8175 : NAND2_X2 port map( A1 => n11330, A2 => n11693, ZN => n3089);
   U769 : INV_X1 port map( I => n17520, ZN => n13035);
   U18361 : INV_X2 port map( I => n19412, ZN => n11234);
   U1090 : INV_X4 port map( I => n26627, ZN => n21097);
   U1664 : INV_X1 port map( I => n21062, ZN => n20561);
   U7139 : NAND3_X2 port map( A1 => n1108, A2 => n20213, A3 => n26009, ZN => 
                           n20214);
   U6636 : INV_X2 port map( I => n7972, ZN => n14990);
   U4169 : INV_X2 port map( I => n17941, ZN => n1217);
   U10180 : NOR2_X2 port map( A1 => n17315, A2 => n1030, ZN => n7194);
   U652 : INV_X1 port map( I => n6770, ZN => n7247);
   U12579 : BUF_X4 port map( I => n7183, Z => n4710);
   U5506 : INV_X1 port map( I => n25380, ZN => n17322);
   U6650 : AOI21_X1 port map( A1 => n1693, A2 => n1692, B => n22060, ZN => 
                           n1690);
   U12233 : INV_X2 port map( I => n26129, ZN => n966);
   U159 : INV_X2 port map( I => n20180, ZN => n25237);
   U3883 : AND2_X1 port map( A1 => n13613, A2 => n15894, Z => n7721);
   U6846 : INV_X2 port map( I => n2671, ZN => n15514);
   U4468 : INV_X2 port map( I => n17942, ZN => n10816);
   U923 : NAND2_X2 port map( A1 => n19159, A2 => n15502, ZN => n6113);
   U18170 : INV_X2 port map( I => n665, ZN => n23748);
   U753 : INV_X4 port map( I => n5612, ZN => n17427);
   U5392 : INV_X4 port map( I => n16244, ZN => n795);
   U689 : OAI21_X2 port map( A1 => n18483, A2 => n18484, B => n880, ZN => 
                           n22561);
   U13551 : NOR2_X2 port map( A1 => n17771, A2 => n886, ZN => n24156);
   U1969 : BUF_X4 port map( I => n13473, Z => n4057);
   U249 : BUF_X2 port map( I => n12995, Z => n25642);
   U766 : NOR2_X2 port map( A1 => n22634, A2 => n19154, ZN => n26446);
   U5826 : INV_X2 port map( I => n10894, ZN => n14222);
   U9496 : INV_X2 port map( I => n3612, ZN => n15523);
   U6331 : NAND2_X2 port map( A1 => n18720, A2 => n14420, ZN => n3612);
   U2222 : NAND2_X1 port map( A1 => n149, A2 => n148, ZN => n9809);
   U12338 : NAND2_X1 port map( A1 => n23196, A2 => n9135, ZN => n22871);
   U18013 : OAI21_X2 port map( A1 => n13877, A2 => n16197, B => n1056, ZN => 
                           n13876);
   U9461 : NAND2_X1 port map( A1 => n23583, A2 => n25798, ZN => n25297);
   U1433 : INV_X2 port map( I => n14450, ZN => n21498);
   U1770 : NAND3_X2 port map( A1 => n24710, A2 => n6035, A3 => n6034, ZN => 
                           n5712);
   U12141 : INV_X2 port map( I => n5529, ZN => n18301);
   U9049 : OR2_X1 port map( A1 => n14997, A2 => n24487, Z => n17187);
   U12940 : NAND3_X2 port map( A1 => n18737, A2 => n18736, A3 => n760, ZN => 
                           n24262);
   U2277 : BUF_X2 port map( I => n9042, Z => n7364);
   U2218 : CLKBUF_X4 port map( I => n16678, Z => n3399);
   U8376 : BUF_X2 port map( I => Key(187), Z => n14598);
   U6170 : OAI21_X2 port map( A1 => n24196, A2 => n971, B => n19947, ZN => 
                           n9178);
   U4122 : INV_X1 port map( I => n9095, ZN => n6122);
   U8134 : NAND3_X2 port map( A1 => n6118, A2 => n6121, A3 => n915, ZN => n6117
                           );
   U1539 : NAND2_X2 port map( A1 => n16224, A2 => n5310, ZN => n16378);
   U12260 : INV_X1 port map( I => n19171, ZN => n2510);
   U1754 : INV_X2 port map( I => n20255, ZN => n20021);
   U2713 : INV_X2 port map( I => n19468, ZN => n26021);
   U10606 : INV_X4 port map( I => n9173, ZN => n14442);
   U12750 : INV_X2 port map( I => n12208, ZN => n1011);
   U12548 : NOR2_X1 port map( A1 => n11295, A2 => n11296, ZN => n6743);
   U8240 : NAND2_X2 port map( A1 => n11693, A2 => n16348, ZN => n13705);
   U20813 : OAI21_X2 port map( A1 => n27456, A2 => n27240, B => n2687, ZN => 
                           n2686);
   U10892 : NAND3_X2 port map( A1 => n6471, A2 => n20054, A3 => n20053, ZN => 
                           n9371);
   U1358 : NOR3_X2 port map( A1 => n8093, A2 => n10533, A3 => n13509, ZN => 
                           n5376);
   U12989 : BUF_X4 port map( I => n14228, Z => n9829);
   U7049 : NOR2_X2 port map( A1 => n6022, A2 => n7798, ZN => n5078);
   U4092 : BUF_X4 port map( I => n5955, Z => n25192);
   U844 : NOR2_X2 port map( A1 => n17915, A2 => n4319, ZN => n13264);
   U17255 : AOI22_X2 port map( A1 => n7615, A2 => n25515, B1 => n2952, B2 => 
                           n17618, ZN => n3877);
   U13411 : INV_X1 port map( I => n28019, ZN => n4452);
   U19047 : NOR2_X1 port map( A1 => n21826, A2 => n8283, ZN => n23878);
   U7150 : INV_X2 port map( I => n8723, ZN => n12973);
   U3236 : BUF_X4 port map( I => n18782, Z => n6031);
   U2199 : NAND2_X2 port map( A1 => n16303, A2 => n16329, ZN => n9364);
   U3262 : AOI21_X2 port map( A1 => n1626, A2 => n5247, B => n19164, ZN => 
                           n1624);
   U5691 : INV_X2 port map( I => n18552, ZN => n18720);
   U10203 : NAND2_X2 port map( A1 => n26920, A2 => n2647, ZN => n9945);
   U7505 : NAND2_X2 port map( A1 => n783, A2 => n22325, ZN => n18716);
   U15021 : INV_X2 port map( I => n20308, ZN => n25603);
   U2319 : INV_X2 port map( I => n237, ZN => n1021);
   U10186 : NOR2_X1 port map( A1 => n6493, A2 => n6492, ZN => n6491);
   U8129 : OR2_X2 port map( A1 => n16109, A2 => n16108, Z => n16110);
   U6917 : NOR2_X1 port map( A1 => n13423, A2 => n22086, ZN => n17859);
   U17881 : NAND2_X1 port map( A1 => n15382, A2 => n16456, ZN => n15381);
   U5198 : NAND3_X1 port map( A1 => n18434, A2 => n736, A3 => n19147, ZN => 
                           n18435);
   U7717 : BUF_X2 port map( I => n13138, Z => n24812);
   U4764 : OAI22_X2 port map( A1 => n5879, A2 => n18781, B1 => n5545, B2 => 
                           n1174, ZN => n3473);
   U18786 : INV_X1 port map( I => n22237, ZN => n9922);
   U12274 : INV_X4 port map( I => n17664, ZN => n13350);
   U1 : OAI21_X2 port map( A1 => n26712, A2 => n20998, B => n26492, ZN => 
                           n21001);
   U664 : OAI21_X2 port map( A1 => n6223, A2 => n2337, B => n18752, ZN => 
                           n23291);
   U9367 : NAND2_X2 port map( A1 => n27558, A2 => n26631, ZN => n2167);
   U751 : OAI21_X2 port map( A1 => n26167, A2 => n3670, B => n11580, ZN => 
                           n3647);
   U422 : INV_X2 port map( I => n4021, ZN => n13255);
   U14685 : NAND3_X2 port map( A1 => n166, A2 => n18779, A3 => n14649, ZN => 
                           n6649);
   U116 : INV_X1 port map( I => n7807, ZN => n7274);
   U20513 : NAND2_X2 port map( A1 => n13, A2 => n12521, ZN => n3181);
   U7453 : BUF_X4 port map( I => n3960, Z => n1158);
   U12111 : INV_X1 port map( I => n19873, ZN => n1131);
   U1256 : NAND2_X1 port map( A1 => n5729, A2 => n16245, ZN => n431);
   U3215 : BUF_X2 port map( I => n14391, Z => n4136);
   U6314 : NAND2_X2 port map( A1 => n9041, A2 => n5306, ZN => n7288);
   U12632 : OAI22_X2 port map( A1 => n13096, A2 => n8735, B1 => n21546, B2 => 
                           n21624, ZN => n9939);
   U5650 : INV_X4 port map( I => n391, ZN => n23564);
   U3148 : INV_X2 port map( I => n23026, ZN => n11363);
   U4598 : INV_X4 port map( I => n879, ZN => n18512);
   U12832 : INV_X4 port map( I => n9911, ZN => n14683);
   U4250 : INV_X2 port map( I => n19870, ZN => n19650);
   U3405 : BUF_X2 port map( I => n18710, Z => n448);
   U21731 : NAND3_X2 port map( A1 => n2938, A2 => n2936, A3 => n2937, ZN => 
                           n24399);
   U1425 : BUF_X2 port map( I => n7371, Z => n401);
   U21681 : NOR2_X2 port map( A1 => n16563, A2 => n16511, ZN => n12668);
   U6323 : NAND2_X2 port map( A1 => n18781, A2 => n1174, ZN => n18504);
   U3780 : NAND2_X2 port map( A1 => n20168, A2 => n7388, ZN => n8610);
   U11227 : OR2_X2 port map( A1 => n9696, A2 => n9698, Z => n1797);
   U7644 : NOR2_X2 port map( A1 => n25655, A2 => n4136, ZN => n24804);
   U3360 : BUF_X2 port map( I => Key(129), Z => n20674);
   U6863 : BUF_X2 port map( I => Key(189), Z => n20908);
   U5121 : NAND2_X2 port map( A1 => n21098, A2 => n12067, ZN => n24260);
   U9774 : BUF_X2 port map( I => n9583, Z => n113);
   U6387 : INV_X2 port map( I => n5985, ZN => n6438);
   U1957 : NAND3_X2 port map( A1 => n6516, A2 => n11689, A3 => n852, ZN => 
                           n6518);
   U2359 : INV_X2 port map( I => n15513, ZN => n15706);
   U4552 : OR2_X2 port map( A1 => n7681, A2 => n25366, Z => n19893);
   U3174 : BUF_X2 port map( I => n19565, Z => n22169);
   U10331 : INV_X2 port map( I => n5243, ZN => n4940);
   U9739 : INV_X2 port map( I => n17666, ZN => n17938);
   U7884 : INV_X1 port map( I => n5541, ZN => n7996);
   U12726 : INV_X2 port map( I => n20189, ZN => n23771);
   U22004 : BUF_X4 port map( I => n23641, Z => n26575);
   U6406 : OR2_X1 port map( A1 => n21740, A2 => n21739, Z => n11168);
   U4674 : AOI21_X2 port map( A1 => n25304, A2 => n14718, B => n773, ZN => 
                           n9823);
   U627 : INV_X4 port map( I => n12885, ZN => n19033);
   U10028 : INV_X2 port map( I => n10559, ZN => n17372);
   U1264 : INV_X2 port map( I => n16338, ZN => n23609);
   U932 : INV_X2 port map( I => n25135, ZN => n915);
   U13537 : INV_X2 port map( I => n21052, ZN => n9425);
   U14923 : OAI21_X2 port map( A1 => n10709, A2 => n15641, B => n13629, ZN => 
                           n13224);
   U18015 : NAND3_X2 port map( A1 => n16350, A2 => n21873, A3 => n7374, ZN => 
                           n11424);
   U2041 : NAND2_X2 port map( A1 => n25795, A2 => n4790, ZN => n10356);
   U5187 : BUF_X2 port map( I => n10190, Z => n62);
   U3711 : OAI21_X2 port map( A1 => n4719, A2 => n6642, B => n10509, ZN => 
                           n9386);
   U7950 : CLKBUF_X4 port map( I => n15609, Z => n1593);
   U15553 : INV_X2 port map( I => n14759, ZN => n21445);
   U7156 : NAND2_X2 port map( A1 => n1108, A2 => n26365, ZN => n5280);
   U7366 : NOR2_X1 port map( A1 => n24424, A2 => n24425, ZN => n4448);
   U14518 : AOI21_X2 port map( A1 => n25517, A2 => n27435, B => n22906, ZN => 
                           n3505);
   U702 : INV_X1 port map( I => n14304, ZN => n19898);
   U21571 : OAI21_X2 port map( A1 => n23864, A2 => n23322, B => n19623, ZN => 
                           n12443);
   U4873 : INV_X2 port map( I => n21063, ZN => n21091);
   U17011 : INV_X2 port map( I => n3960, ZN => n8714);
   U16452 : INV_X4 port map( I => n7586, ZN => n20938);
   U4083 : INV_X2 port map( I => n4508, ZN => n23063);
   U2075 : INV_X2 port map( I => n13066, ZN => n2533);
   U671 : INV_X1 port map( I => n23245, ZN => n11872);
   U1343 : BUF_X4 port map( I => n1483, Z => n21768);
   U7452 : NAND2_X1 port map( A1 => n18697, A2 => n18698, ZN => n18699);
   U4963 : OAI22_X2 port map( A1 => n13565, A2 => n12983, B1 => n11770, B2 => 
                           n28247, ZN => n12789);
   U9307 : AOI21_X2 port map( A1 => n4844, A2 => n22981, B => n8049, ZN => 
                           n18950);
   U10275 : NAND2_X2 port map( A1 => n16725, A2 => n3537, ZN => n16723);
   U8337 : BUF_X2 port map( I => Key(25), Z => n20941);
   U15549 : OR3_X2 port map( A1 => n16559, A2 => n16558, A3 => n12637, Z => 
                           n11726);
   U6186 : AND3_X1 port map( A1 => n1175, A2 => n23761, A3 => n18578, Z => 
                           n24611);
   U14124 : NAND2_X2 port map( A1 => n25135, A2 => n16318, ZN => n25462);
   U2628 : OR2_X2 port map( A1 => n11842, A2 => n25349, Z => n14821);
   U2334 : NOR2_X2 port map( A1 => n5310, A2 => n27019, ZN => n1982);
   U9680 : NAND2_X1 port map( A1 => n7801, A2 => n7800, ZN => n7804);
   U15849 : NAND3_X2 port map( A1 => n25709, A2 => n8113, A3 => n25708, ZN => 
                           n3742);
   U13586 : OAI21_X2 port map( A1 => n6910, A2 => n2068, B => n5117, ZN => 
                           n4459);
   U65 : NAND2_X1 port map( A1 => n20063, A2 => n13448, ZN => n13445);
   U2928 : OR2_X2 port map( A1 => n21388, A2 => n15209, Z => n21273);
   U20368 : NOR2_X2 port map( A1 => n26336, A2 => n18914, ZN => n2727);
   U10320 : INV_X1 port map( I => n1711, ZN => n9950);
   U1791 : NOR2_X2 port map( A1 => n3343, A2 => n3342, ZN => n25684);
   U1629 : INV_X2 port map( I => n8786, ZN => n19689);
   U17202 : INV_X4 port map( I => n9116, ZN => n9139);
   U245 : NAND2_X2 port map( A1 => n19797, A2 => n26120, ZN => n4632);
   U11228 : INV_X4 port map( I => n9143, ZN => n5353);
   U12410 : INV_X4 port map( I => n4531, ZN => n10133);
   U3043 : NAND2_X2 port map( A1 => n24260, A2 => n24259, ZN => n20925);
   U663 : INV_X4 port map( I => n864, ZN => n10272);
   U4973 : NAND2_X1 port map( A1 => n7412, A2 => n7411, ZN => n18059);
   U16688 : INV_X2 port map( I => n977, ZN => n15376);
   U6407 : NOR2_X2 port map( A1 => n8843, A2 => n1119, ZN => n22109);
   U5866 : NAND2_X2 port map( A1 => n978, A2 => n10520, ZN => n8843);
   U4808 : OAI21_X2 port map( A1 => n18685, A2 => n18466, B => n18256, ZN => 
                           n7888);
   U1523 : OAI21_X2 port map( A1 => n15701, A2 => n16435, B => n25862, ZN => 
                           n9275);
   U4700 : BUF_X4 port map( I => n819, Z => n24454);
   U2662 : NAND2_X1 port map( A1 => n4981, A2 => n13963, ZN => n270);
   U12967 : NOR4_X2 port map( A1 => n7289, A2 => n2544, A3 => n5837, A4 => 
                           n5836, ZN => n22906);
   U15224 : INV_X1 port map( I => n16534, ZN => n13496);
   U4775 : INV_X2 port map( I => n15362, ZN => n18458);
   U16409 : NOR2_X2 port map( A1 => n7395, A2 => n26760, ZN => n16484);
   U6529 : NOR3_X2 port map( A1 => n3545, A2 => n27959, A3 => n5353, ZN => 
                           n2499);
   U2244 : AOI21_X2 port map( A1 => n11803, A2 => n21022, B => n11801, ZN => 
                           n11800);
   U10991 : AOI22_X1 port map( A1 => n15720, A2 => n9421, B1 => n21045, B2 => 
                           n25352, ZN => n26306);
   U9832 : AOI22_X1 port map( A1 => n17793, A2 => n27424, B1 => n23806, B2 => 
                           n5218, ZN => n17796);
   U5014 : INV_X4 port map( I => n3347, ZN => n17727);
   U16781 : INV_X1 port map( I => n8032, ZN => n25843);
   U5966 : NAND2_X2 port map( A1 => n19714, A2 => n19468, ZN => n19950);
   U5186 : NAND2_X2 port map( A1 => n12495, A2 => n15246, ZN => n3074);
   U11304 : OAI21_X2 port map( A1 => n12104, A2 => n1893, B => n12494, ZN => 
                           n4390);
   U5822 : INV_X2 port map( I => n9509, ZN => n4618);
   U5348 : INV_X2 port map( I => n15916, ZN => n730);
   U6500 : NAND3_X2 port map( A1 => n13920, A2 => n27492, A3 => n13919, ZN => 
                           n13917);
   U21590 : AOI21_X2 port map( A1 => n20590, A2 => n5042, B => n24285, ZN => 
                           n7672);
   U8230 : NAND2_X2 port map( A1 => n16303, A2 => n720, ZN => n9363);
   U2975 : INV_X2 port map( I => n18221, ZN => n9727);
   U4520 : NAND2_X2 port map( A1 => n3401, A2 => n8735, ZN => n8742);
   U18389 : BUF_X4 port map( I => n20523, Z => n13808);
   U614 : NAND2_X1 port map( A1 => n25096, A2 => n19646, ZN => n2021);
   U2559 : NAND2_X1 port map( A1 => n11243, A2 => n8245, ZN => n243);
   U10427 : AOI21_X2 port map( A1 => n15837, A2 => n15836, B => n11429, ZN => 
                           n12837);
   U21663 : OAI21_X2 port map( A1 => n524, A2 => n16340, B => n15615, ZN => 
                           n14571);
   U9286 : OAI21_X1 port map( A1 => n8313, A2 => n28547, B => n8312, ZN => 
                           n10807);
   U16809 : INV_X4 port map( I => n8423, ZN => n10580);
   U12514 : AOI21_X2 port map( A1 => n25315, A2 => n22764, B => n842, ZN => 
                           n6923);
   U3667 : BUF_X4 port map( I => n1062, Z => n524);
   U4279 : BUF_X4 port map( I => n5197, Z => n2789);
   U11273 : INV_X4 port map( I => n1062, ZN => n16113);
   U12209 : NAND2_X2 port map( A1 => n18496, A2 => n18750, ZN => n15266);
   U14544 : NAND2_X2 port map( A1 => n13488, A2 => n26822, ZN => n25525);
   U589 : BUF_X4 port map( I => n14210, Z => n22894);
   U11018 : NAND2_X2 port map( A1 => n10520, A2 => n19728, ZN => n25655);
   U8673 : INV_X2 port map( I => n3880, ZN => n26052);
   U4443 : NAND3_X2 port map( A1 => n18727, A2 => n18728, A3 => n10930, ZN => 
                           n5131);
   U394 : NOR2_X1 port map( A1 => n2652, A2 => n5263, ZN => n12185);
   U17964 : NAND2_X2 port map( A1 => n7263, A2 => n20561, ZN => n23728);
   U20137 : INV_X1 port map( I => n17956, ZN => n8117);
   U7791 : NAND3_X1 port map( A1 => n11029, A2 => n22578, A3 => n11030, ZN => 
                           n2752);
   U13604 : NAND2_X2 port map( A1 => n21529, A2 => n12625, ZN => n21535);
   U10453 : AOI22_X2 port map( A1 => n1856, A2 => n8530, B1 => n22496, B2 => 
                           n27160, ZN => n1854);
   U21313 : INV_X2 port map( I => n21153, ZN => n20475);
   U806 : OAI22_X2 port map( A1 => n26327, A2 => n2091, B1 => n19044, B2 => 
                           n23575, ZN => n251);
   U20650 : NAND2_X2 port map( A1 => n23828, A2 => n703, ZN => n26357);
   U13052 : INV_X1 port map( I => n18245, ZN => n22363);
   U2889 : CLKBUF_X4 port map( I => n6698, Z => n852);
   U117 : INV_X4 port map( I => n26882, ZN => n951);
   U9475 : NAND2_X1 port map( A1 => n18439, A2 => n2594, ZN => n2603);
   U5538 : INV_X2 port map( I => n19949, ZN => n19828);
   U397 : NAND2_X2 port map( A1 => n18825, A2 => n10323, ZN => n1845);
   U19110 : NOR2_X1 port map( A1 => n7107, A2 => n26157, ZN => n26170);
   U12993 : NAND2_X1 port map( A1 => n6852, A2 => n6851, ZN => n6850);
   U1265 : AOI21_X2 port map( A1 => n16196, A2 => n16307, B => n14886, ZN => 
                           n12840);
   U14962 : NAND2_X2 port map( A1 => n19742, A2 => n26129, ZN => n13345);
   U20615 : NAND2_X2 port map( A1 => n28369, A2 => n14579, ZN => n16476);
   U1099 : AOI22_X2 port map( A1 => n16386, A2 => n24183, B1 => n5558, B2 => 
                           n15571, ZN => n23113);
   U5419 : NOR2_X2 port map( A1 => n15186, A2 => n22614, ZN => n16386);
   U10154 : NOR2_X1 port map( A1 => n25660, A2 => n25659, ZN => n25658);
   U5964 : NOR2_X2 port map( A1 => n12512, A2 => n14423, ZN => n19600);
   U2808 : BUF_X4 port map( I => n26646, Z => n16303);
   U16685 : NAND2_X1 port map( A1 => n26137, A2 => n6282, ZN => n26136);
   U10723 : BUF_X4 port map( I => n14586, Z => n9264);
   U11878 : AND2_X2 port map( A1 => n6777, A2 => n7169, Z => n9348);
   U7278 : NOR2_X1 port map( A1 => n13722, A2 => n5253, ZN => n8525);
   U12953 : AOI21_X1 port map( A1 => n11994, A2 => n759, B => n18582, ZN => 
                           n10804);
   U21232 : INV_X2 port map( I => n665, ZN => n13571);
   U7120 : NOR2_X2 port map( A1 => n745, A2 => n22224, ZN => n5248);
   U4522 : NAND2_X1 port map( A1 => n11464, A2 => n25936, ZN => n26413);
   U16437 : INV_X1 port map( I => n20680, ZN => n25809);
   U7335 : AOI21_X1 port map( A1 => n19061, A2 => n13596, B => n13595, ZN => 
                           n13594);
   U4299 : BUF_X1 port map( I => n17457, Z => n3752);
   U2339 : NAND2_X1 port map( A1 => n11113, A2 => n22840, ZN => n6653);
   U7421 : INV_X2 port map( I => n19101, ZN => n18800);
   U18596 : NAND2_X2 port map( A1 => n23984, A2 => n12573, ZN => n11890);
   U19550 : NAND2_X2 port map( A1 => n18537, A2 => n1010, ZN => n23984);
   U5921 : OR2_X2 port map( A1 => n19693, A2 => n19778, Z => n19597);
   U426 : INV_X2 port map( I => n114, ZN => n19082);
   U9938 : NAND3_X2 port map( A1 => n5503, A2 => n8146, A3 => n8144, ZN => 
                           n6894);
   U14722 : NAND2_X2 port map( A1 => n12911, A2 => n12912, ZN => n25548);
   U12835 : BUF_X4 port map( I => n114, Z => n24265);
   U5683 : INV_X4 port map( I => n15037, ZN => n3545);
   U7017 : INV_X2 port map( I => n773, ZN => n15208);
   U1893 : NAND2_X2 port map( A1 => n5055, A2 => n18837, ZN => n26070);
   U2767 : NAND2_X1 port map( A1 => n12402, A2 => n22045, ZN => n15153);
   U5134 : NAND2_X1 port map( A1 => n23537, A2 => n26109, ZN => n26057);
   U5819 : NOR2_X1 port map( A1 => n8128, A2 => n8127, ZN => n8131);
   U16803 : NAND2_X2 port map( A1 => n11023, A2 => n460, ZN => n12153);
   U7588 : INV_X4 port map( I => n20269, ZN => n23592);
   U10167 : NAND2_X2 port map( A1 => n26457, A2 => n18830, ZN => n25818);
   U6981 : NAND3_X2 port map( A1 => n26676, A2 => n13172, A3 => n13432, ZN => 
                           n9805);
   U11124 : NAND3_X2 port map( A1 => n7888, A2 => n18467, A3 => n26209, ZN => 
                           n8171);
   U12449 : INV_X1 port map( I => n25829, ZN => n10604);
   U7454 : INV_X2 port map( I => n26644, ZN => n7980);
   U3514 : AND2_X2 port map( A1 => n15557, A2 => n14567, Z => n21669);
   U10942 : NAND2_X1 port map( A1 => n3164, A2 => n3166, ZN => n18657);
   U5972 : NAND2_X2 port map( A1 => n11372, A2 => n24862, ZN => n11370);
   U14365 : NAND2_X2 port map( A1 => n4953, A2 => n26644, ZN => n18946);
   U509 : NAND2_X1 port map( A1 => n23822, A2 => n23821, ZN => n12459);
   U7608 : NOR2_X1 port map( A1 => n24796, A2 => n26504, ZN => n17731);
   U447 : NAND2_X1 port map( A1 => n23059, A2 => n23057, ZN => n18911);
   U9296 : NAND2_X2 port map( A1 => n10323, A2 => n1329, ZN => n1328);
   U15616 : INV_X1 port map( I => n25104, ZN => n9946);
   U4477 : BUF_X4 port map( I => n20234, Z => n26252);
   U8372 : BUF_X2 port map( I => Key(117), Z => n21419);
   U5635 : CLKBUF_X4 port map( I => n18772, Z => n14648);
   U10668 : CLKBUF_X2 port map( I => Key(126), Z => n14479);
   U5056 : NAND2_X2 port map( A1 => n3966, A2 => n3965, ZN => n11748);
   U1872 : NOR2_X2 port map( A1 => n16337, A2 => n9308, ZN => n7722);
   U504 : NAND2_X1 port map( A1 => n26208, A2 => n26207, ZN => n23098);
   U4839 : INV_X2 port map( I => n18891, ZN => n19079);
   U9362 : AOI21_X2 port map( A1 => n18802, A2 => n18801, B => n18800, ZN => 
                           n18803);
   U3571 : OAI21_X1 port map( A1 => n11370, A2 => n4858, B => n11255, ZN => 
                           n22199);
   U19824 : INV_X2 port map( I => n14852, ZN => n14679);
   U2990 : NOR2_X2 port map( A1 => n2761, A2 => n23958, ZN => n23957);
   U13055 : NOR2_X2 port map( A1 => n1202, A2 => n9344, ZN => n11663);
   U9565 : AND3_X2 port map( A1 => n877, A2 => n25500, A3 => n18455, Z => n1499
                           );
   U12760 : NAND2_X2 port map( A1 => n15315, A2 => n20588, ZN => n15288);
   U2378 : INV_X2 port map( I => n477, ZN => n23088);
   U1053 : BUF_X2 port map( I => n10971, Z => n3902);
   U2907 : INV_X2 port map( I => n11982, ZN => n21776);
   U5493 : INV_X4 port map( I => n11992, ZN => n7498);
   U2746 : NAND2_X1 port map( A1 => n294, A2 => n293, ZN => n8815);
   U7334 : AOI21_X2 port map( A1 => n10709, A2 => n28173, B => n15641, ZN => 
                           n12751);
   U7283 : NOR2_X2 port map( A1 => n19714, A2 => n19828, ZN => n19467);
   U1660 : OAI21_X2 port map( A1 => n1658, A2 => n7567, B => n19105, ZN => 
                           n7174);
   U17776 : NAND3_X2 port map( A1 => n27557, A2 => n9994, A3 => n11110, ZN => 
                           n19713);
   U7546 : NAND3_X2 port map( A1 => n14417, A2 => n5457, A3 => n25712, ZN => 
                           n5750);
   U6633 : INV_X1 port map( I => n2960, ZN => n17303);
   U12360 : INV_X2 port map( I => n18479, ZN => n2949);
   U6581 : INV_X2 port map( I => n26110, ZN => n21901);
   U4021 : NAND2_X2 port map( A1 => n22113, A2 => n14980, ZN => n7412);
   U18586 : INV_X1 port map( I => Key(164), ZN => n13859);
   U8355 : CLKBUF_X2 port map( I => Key(3), Z => n20605);
   U4344 : BUF_X2 port map( I => Key(24), Z => n21436);
   U5230 : CLKBUF_X2 port map( I => Key(132), Z => n21090);
   U8379 : BUF_X2 port map( I => Key(160), Z => n14340);
   U4399 : BUF_X2 port map( I => Key(84), Z => n14588);
   U8365 : BUF_X2 port map( I => Key(0), Z => n21357);
   U8374 : BUF_X2 port map( I => Key(131), Z => n21411);
   U8391 : BUF_X2 port map( I => Key(124), Z => n14473);
   U10679 : BUF_X2 port map( I => Key(154), Z => n14506);
   U10711 : BUF_X2 port map( I => Key(4), Z => n14558);
   U8328 : BUF_X2 port map( I => Key(142), Z => n20952);
   U6874 : BUF_X2 port map( I => Key(177), Z => n10544);
   U5086 : CLKBUF_X2 port map( I => Key(123), Z => n20369);
   U10644 : BUF_X2 port map( I => Key(37), Z => n7355);
   U10707 : BUF_X2 port map( I => Key(34), Z => n14404);
   U8282 : INV_X1 port map( I => n13418, ZN => n16077);
   U10615 : BUF_X2 port map( I => n16006, Z => n14108);
   U13177 : CLKBUF_X4 port map( I => n16228, Z => n10001);
   U5401 : CLKBUF_X1 port map( I => n16158, Z => n7311);
   U11582 : OR2_X1 port map( A1 => n5448, A2 => n22590, Z => n15831);
   U10633 : INV_X1 port map( I => n14537, ZN => n13787);
   U11608 : INV_X2 port map( I => n25253, ZN => n21904);
   U10649 : INV_X1 port map( I => n20674, ZN => n1277);
   U10587 : BUF_X2 port map( I => n12271, Z => n5362);
   U8291 : INV_X1 port map( I => n14543, ZN => n1298);
   U3517 : CLKBUF_X4 port map( I => n11813, Z => n7868);
   U10622 : INV_X1 port map( I => n20961, ZN => n15731);
   U2645 : CLKBUF_X4 port map( I => n21874, Z => n21773);
   U5396 : CLKBUF_X1 port map( I => n15491, Z => n7351);
   U4153 : CLKBUF_X2 port map( I => n16128, Z => n263);
   U5285 : CLKBUF_X4 port map( I => n15832, Z => n24581);
   U4656 : CLKBUF_X2 port map( I => n16342, Z => n14293);
   U15530 : NOR2_X1 port map( A1 => n6314, A2 => n7374, ZN => n13438);
   U10638 : BUF_X2 port map( I => n14843, Z => n7152);
   U4846 : INV_X2 port map( I => n16196, ZN => n2111);
   U1727 : CLKBUF_X4 port map( I => n10629, Z => n12918);
   U11932 : CLKBUF_X4 port map( I => n841, Z => n250);
   U13294 : CLKBUF_X2 port map( I => n27469, Z => n24198);
   U2084 : CLKBUF_X4 port map( I => n15886, Z => n121);
   U8258 : INV_X2 port map( I => n14557, ZN => n16239);
   U16245 : NAND2_X1 port map( A1 => n12678, A2 => n25774, ZN => n25773);
   U1693 : NAND2_X1 port map( A1 => n12507, A2 => n11291, ZN => n24875);
   U1845 : OAI21_X1 port map( A1 => n24588, A2 => n15955, B => n11830, ZN => 
                           n11829);
   U14841 : AOI21_X1 port map( A1 => n4751, A2 => n15788, B => n6647, ZN => 
                           n23135);
   U14026 : AOI21_X1 port map( A1 => n25457, A2 => n4751, B => n25444, ZN => 
                           n25597);
   U1084 : CLKBUF_X4 port map( I => n11775, Z => n9725);
   U1706 : NAND2_X1 port map( A1 => n7125, A2 => n7123, ZN => n10321);
   U3366 : CLKBUF_X1 port map( I => n16466, Z => n23529);
   U5212 : CLKBUF_X2 port map( I => n23744, Z => n25554);
   U5046 : CLKBUF_X2 port map( I => n16585, Z => n7115);
   U2285 : INV_X2 port map( I => n6373, ZN => n16713);
   U1189 : CLKBUF_X4 port map( I => n124, Z => n23439);
   U2472 : INV_X2 port map( I => n27734, ZN => n16695);
   U22041 : CLKBUF_X2 port map( I => n28400, Z => n26594);
   U4313 : CLKBUF_X4 port map( I => n7395, Z => n4998);
   U10282 : INV_X1 port map( I => n16540, ZN => n2118);
   U15998 : NAND2_X1 port map( A1 => n15528, A2 => n15527, ZN => n15337);
   U1711 : NAND2_X1 port map( A1 => n1792, A2 => n7308, ZN => n16693);
   U983 : NAND2_X1 port map( A1 => n10260, A2 => n10259, ZN => n16424);
   U5192 : NAND2_X1 port map( A1 => n16663, A2 => n26174, ZN => n16371);
   U3461 : CLKBUF_X2 port map( I => n14618, Z => n465);
   U7163 : OAI21_X1 port map( A1 => n16500, A2 => n22110, B => n1761, ZN => 
                           n1760);
   U18820 : CLKBUF_X2 port map( I => n23053, Z => n26132);
   U18043 : INV_X1 port map( I => n15256, ZN => n17065);
   U8264 : CLKBUF_X4 port map( I => n26084, Z => n24885);
   U3593 : CLKBUF_X4 port map( I => n10443, Z => n1709);
   U18461 : CLKBUF_X4 port map( I => n16915, Z => n26082);
   U5472 : INV_X1 port map( I => n13856, ZN => n7209);
   U6931 : CLKBUF_X4 port map( I => n14723, Z => n1232);
   U3840 : BUF_X2 port map( I => n17369, Z => n24567);
   U10096 : CLKBUF_X2 port map( I => n17414, Z => n5500);
   U17291 : INV_X2 port map( I => n3296, ZN => n17541);
   U694 : INV_X1 port map( I => n12040, ZN => n17286);
   U10121 : BUF_X2 port map( I => n17003, Z => n17452);
   U7942 : INV_X2 port map( I => n26081, ZN => n1040);
   U5104 : BUF_X2 port map( I => n21774, Z => n26418);
   U789 : INV_X2 port map( I => n899, ZN => n1233);
   U5101 : CLKBUF_X4 port map( I => n17160, Z => n11113);
   U749 : INV_X2 port map( I => n21798, ZN => n14061);
   U13071 : NAND2_X1 port map( A1 => n12340, A2 => n17543, ZN => n15031);
   U2122 : NAND2_X1 port map( A1 => n17307, A2 => n17303, ZN => n17304);
   U20306 : NOR2_X1 port map( A1 => n5845, A2 => n26332, ZN => n5844);
   U14697 : OR2_X1 port map( A1 => n10912, A2 => n10913, Z => n5282);
   U8644 : OAI21_X1 port map( A1 => n22275, A2 => n23926, B => n22274, ZN => 
                           n17243);
   U11802 : INV_X1 port map( I => n6183, ZN => n25265);
   U2514 : NAND2_X1 port map( A1 => n231, A2 => n229, ZN => n17001);
   U5697 : NAND2_X1 port map( A1 => n21952, A2 => n1231, ZN => n16828);
   U9934 : NAND2_X1 port map( A1 => n9610, A2 => n10160, ZN => n9607);
   U20686 : NAND3_X1 port map( A1 => n16878, A2 => n1224, A3 => n10546, ZN => 
                           n16879);
   U3601 : NAND2_X1 port map( A1 => n17393, A2 => n17472, ZN => n508);
   U13649 : NAND2_X1 port map( A1 => n23025, A2 => n25568, ZN => n23151);
   U9939 : NOR2_X1 port map( A1 => n17383, A2 => n13374, ZN => n14615);
   U4123 : CLKBUF_X2 port map( I => n413, Z => n23441);
   U4283 : CLKBUF_X4 port map( I => n2460, Z => n1882);
   U5018 : CLKBUF_X2 port map( I => n14397, Z => n24881);
   U5023 : INV_X2 port map( I => n14397, ZN => n11419);
   U4124 : CLKBUF_X2 port map( I => n17665, Z => n7140);
   U7785 : BUF_X4 port map( I => n17992, Z => n6642);
   U1755 : CLKBUF_X4 port map( I => n391, Z => n47);
   U4096 : CLKBUF_X4 port map( I => n17578, Z => n23197);
   U1308 : CLKBUF_X4 port map( I => n17926, Z => n25929);
   U4980 : INV_X2 port map( I => n5368, ZN => n1026);
   U3328 : CLKBUF_X2 port map( I => n3292, Z => n23963);
   U2693 : INV_X2 port map( I => n17962, ZN => n787);
   U4972 : INV_X1 port map( I => n17656, ZN => n25787);
   U1259 : NAND2_X1 port map( A1 => n8884, A2 => n27424, ZN => n26608);
   U4965 : AOI21_X1 port map( A1 => n5892, A2 => n13216, B => n4590, ZN => 
                           n24796);
   U5600 : NOR2_X1 port map( A1 => n10059, A2 => n17847, ZN => n17848);
   U1294 : INV_X1 port map( I => n17739, ZN => n24958);
   U14548 : NOR2_X1 port map( A1 => n13848, A2 => n13849, ZN => n9210);
   U16712 : INV_X1 port map( I => n25837, ZN => n22176);
   U5597 : OAI21_X1 port map( A1 => n9905, A2 => n1025, B => n4503, ZN => n4502
                           );
   U3216 : NAND2_X1 port map( A1 => n14111, A2 => n14112, ZN => n17600);
   U791 : BUF_X2 port map( I => n4970, Z => n24255);
   U4029 : NAND2_X1 port map( A1 => n4502, A2 => n4504, ZN => n23283);
   U1463 : NAND2_X1 port map( A1 => n3172, A2 => n3173, ZN => n24065);
   U12713 : CLKBUF_X4 port map( I => n12205, Z => n24357);
   U4602 : INV_X2 port map( I => n21923, ZN => n820);
   U10897 : INV_X2 port map( I => n6777, ZN => n10437);
   U2350 : CLKBUF_X4 port map( I => n18443, Z => n18785);
   U9653 : CLKBUF_X2 port map( I => n18725, Z => n14427);
   U10123 : INV_X2 port map( I => n22799, ZN => n7591);
   U732 : INV_X2 port map( I => n10437, ZN => n8269);
   U1646 : NAND2_X1 port map( A1 => n2325, A2 => n18780, ZN => n2120);
   U5723 : INV_X1 port map( I => n3215, ZN => n18568);
   U6398 : NOR2_X1 port map( A1 => n1013, A2 => n18507, ZN => n12954);
   U3527 : INV_X2 port map( I => n1018, ZN => n2081);
   U13027 : INV_X2 port map( I => n18442, ZN => n18774);
   U17807 : NAND2_X1 port map( A1 => n18706, A2 => n28306, ZN => n15397);
   U17805 : NOR2_X1 port map( A1 => n5561, A2 => n25261, ZN => n111);
   U7605 : INV_X2 port map( I => n18445, ZN => n1180);
   U9476 : NAND2_X1 port map( A1 => n3699, A2 => n8113, ZN => n3698);
   U4716 : NAND2_X1 port map( A1 => n11058, A2 => n18755, ZN => n26284);
   U3967 : NOR2_X1 port map( A1 => n23006, A2 => n23005, ZN => n1378);
   U7486 : NOR2_X1 port map( A1 => n18707, A2 => n25708, ZN => n15599);
   U14489 : NAND2_X1 port map( A1 => n18700, A2 => n24870, ZN => n23037);
   U7600 : OR2_X1 port map( A1 => n24054, A2 => n5691, Z => n5690);
   U430 : INV_X2 port map( I => n18933, ZN => n19017);
   U1470 : INV_X1 port map( I => n8611, ZN => n1153);
   U1947 : INV_X2 port map( I => n19126, ZN => n12583);
   U902 : INV_X2 port map( I => n18921, ZN => n873);
   U956 : CLKBUF_X4 port map( I => n10894, Z => n25984);
   U933 : CLKBUF_X4 port map( I => n2617, Z => n26327);
   U2274 : CLKBUF_X4 port map( I => n11906, Z => n447);
   U4614 : NAND2_X1 port map( A1 => n3671, A2 => n7597, ZN => n3646);
   U1464 : INV_X1 port map( I => n19373, ZN => n24189);
   U3827 : CLKBUF_X2 port map( I => n7126, Z => n22939);
   U12178 : NAND2_X1 port map( A1 => n23434, A2 => n23432, ZN => n18855);
   U3818 : INV_X1 port map( I => n19565, ZN => n22120);
   U11786 : NAND2_X1 port map( A1 => n27441, A2 => n25006, ZN => n12546);
   U3785 : CLKBUF_X4 port map( I => n10105, Z => n10041);
   U9179 : INV_X1 port map( I => n19410, ZN => n2702);
   U6364 : CLKBUF_X4 port map( I => n19778, Z => n13194);
   U4556 : CLKBUF_X4 port map( I => n19684, Z => n19951);
   U1345 : BUF_X2 port map( I => n664, Z => n6976);
   U9151 : CLKBUF_X4 port map( I => n19614, Z => n12393);
   U4580 : CLKBUF_X4 port map( I => n7681, Z => n21769);
   U4735 : CLKBUF_X4 port map( I => n13909, Z => n8754);
   U10447 : CLKBUF_X4 port map( I => n22978, Z => n10498);
   U3140 : INV_X1 port map( I => n19791, ZN => n14531);
   U21306 : INV_X4 port map( I => n26415, ZN => n14304);
   U21758 : INV_X2 port map( I => n2057, ZN => n24431);
   U3708 : CLKBUF_X2 port map( I => n19741, Z => n329);
   U7302 : CLKBUF_X2 port map( I => n11619, Z => n10293);
   U3134 : CLKBUF_X4 port map( I => n26621, Z => n22422);
   U21273 : BUF_X1 port map( I => n9612, Z => n24235);
   U2575 : BUF_X2 port map( I => n14356, Z => n23145);
   U594 : INV_X1 port map( I => n19766, ZN => n10080);
   U3722 : NAND2_X1 port map( A1 => n13660, A2 => n4132, ZN => n13666);
   U646 : CLKBUF_X4 port map( I => n12218, Z => n24184);
   U11747 : NAND2_X1 port map( A1 => n22883, A2 => n11063, ZN => n11061);
   U6147 : NAND2_X1 port map( A1 => n19938, A2 => n27730, ZN => n15367);
   U9130 : INV_X1 port map( I => n8048, ZN => n13760);
   U6104 : OAI21_X1 port map( A1 => n19283, A2 => n10196, B => n329, ZN => 
                           n2171);
   U8985 : NAND2_X1 port map( A1 => n4480, A2 => n3424, ZN => n3727);
   U17301 : OR2_X1 port map( A1 => n19629, A2 => n10562, Z => n9382);
   U3635 : CLKBUF_X2 port map( I => n5934, Z => n23558);
   U1736 : CLKBUF_X4 port map( I => n20059, Z => n7122);
   U1854 : INV_X1 port map( I => n8135, ZN => n20143);
   U12612 : CLKBUF_X4 port map( I => n8135, Z => n5049);
   U266 : CLKBUF_X2 port map( I => n14213, Z => n24315);
   U8938 : INV_X2 port map( I => n11871, ZN => n11870);
   U2146 : CLKBUF_X2 port map( I => n5231, Z => n135);
   U4459 : CLKBUF_X1 port map( I => n20168, Z => n25175);
   U1284 : NOR2_X1 port map( A1 => n12746, A2 => n20290, ZN => n13076);
   U8802 : INV_X1 port map( I => n6313, ZN => n20185);
   U20195 : NAND2_X1 port map( A1 => n8610, A2 => n11372, ZN => n3302);
   U4390 : INV_X1 port map( I => n20287, ZN => n25154);
   U6033 : OR2_X1 port map( A1 => n20039, A2 => n5967, Z => n2199);
   U6017 : AOI21_X1 port map( A1 => n20114, A2 => n20192, B => n955, ZN => 
                           n5014);
   U12667 : NOR2_X1 port map( A1 => n809, A2 => n22745, ZN => n9960);
   U2159 : CLKBUF_X4 port map( I => n21148, Z => n136);
   U4218 : CLKBUF_X4 port map( I => n21369, Z => n9678);
   U15201 : NAND2_X1 port map( A1 => n3081, A2 => n15391, ZN => n3080);
   U12064 : INV_X2 port map( I => n12315, ZN => n12309);
   U4872 : BUF_X2 port map( I => n21547, Z => n14406);
   U12415 : CLKBUF_X1 port map( I => n3592, Z => n25309);
   U6070 : INV_X2 port map( I => n21507, ZN => n21592);
   U15248 : INV_X2 port map( I => n5807, ZN => n13505);
   U6376 : BUF_X2 port map( I => n21271, Z => n14409);
   U5961 : AND2_X1 port map( A1 => n20972, A2 => n25388, Z => n21094);
   U8675 : BUF_X1 port map( I => n20593, Z => n3299);
   U3324 : OR2_X1 port map( A1 => n9702, A2 => n13642, Z => n8215);
   U21158 : INV_X1 port map( I => n21140, ZN => n21138);
   U6998 : INV_X1 port map( I => n20860, ZN => n20861);
   U4232 : CLKBUF_X4 port map( I => n20817, Z => n7330);
   U9133 : OR3_X1 port map( A1 => n21549, A2 => n12900, A3 => n14679, Z => 
                           n10883);
   U7900 : OAI21_X1 port map( A1 => n10623, A2 => n216, B => n13388, ZN => 
                           n24835);
   U10978 : NAND2_X1 port map( A1 => n13088, A2 => n8327, ZN => n22555);
   U5425 : NAND2_X1 port map( A1 => n13847, A2 => n14460, ZN => n13845);
   U4673 : NAND2_X1 port map( A1 => n11468, A2 => n4879, ZN => n9976);
   U10240 : INV_X2 port map( I => n24381, ZN => n696);
   U1908 : BUF_X4 port map( I => n4890, Z => n24562);
   U28 : CLKBUF_X2 port map( I => n21538, Z => n9575);
   U12792 : OAI21_X1 port map( A1 => n20997, A2 => n12188, B => n12186, ZN => 
                           n12187);
   U3411 : NAND2_X1 port map( A1 => n6406, A2 => n20748, ZN => n24071);
   U16096 : NOR2_X2 port map( A1 => n15980, A2 => n15981, ZN => n16135);
   U5660 : INV_X4 port map( I => n11364, ZN => n13996);
   U8932 : INV_X2 port map( I => n9956, ZN => n1102);
   U541 : OAI21_X2 port map( A1 => n5883, A2 => n15067, B => n24365, ZN => 
                           n19853);
   U3153 : OAI21_X2 port map( A1 => n12393, A2 => n8330, B => n15067, ZN => 
                           n24365);
   U1306 : NAND4_X2 port map( A1 => n1349, A2 => n21792, A3 => n17504, A4 => 
                           n17505, ZN => n14776);
   U3842 : BUF_X2 port map( I => n13825, Z => n22123);
   U7656 : BUF_X2 port map( I => n17806, Z => n22165);
   U18385 : INV_X1 port map( I => n26068, ZN => n10830);
   U6825 : INV_X2 port map( I => n16273, ZN => n1263);
   U5080 : INV_X1 port map( I => n16274, ZN => n13562);
   U3584 : INV_X1 port map( I => n10035, ZN => n16269);
   U12834 : NAND2_X1 port map( A1 => n24216, A2 => n24643, ZN => n2405);
   U3512 : INV_X1 port map( I => n11813, ZN => n16226);
   U1635 : BUF_X2 port map( I => n333, Z => n11);
   U3368 : INV_X1 port map( I => n10629, ZN => n769);
   U5406 : INV_X1 port map( I => n16143, ZN => n15983);
   U4508 : INV_X1 port map( I => n14843, ZN => n16334);
   U5821 : INV_X1 port map( I => n16107, ZN => n8867);
   U1267 : INV_X1 port map( I => n15491, ZN => n23104);
   U4367 : NOR2_X1 port map( A1 => n11940, A2 => n15918, ZN => n12152);
   U21863 : INV_X1 port map( I => n28284, ZN => n16076);
   U4353 : NOR2_X1 port map( A1 => n8696, A2 => n795, ZN => n22935);
   U4436 : BUF_X2 port map( I => n7910, Z => n460);
   U3430 : INV_X2 port map( I => n16220, ZN => n16254);
   U16594 : CLKBUF_X2 port map( I => n16231, Z => n25816);
   U3272 : INV_X2 port map( I => n6315, ZN => n1264);
   U3585 : BUF_X2 port map( I => n10035, Z => n9393);
   U1266 : NOR2_X1 port map( A1 => n9223, A2 => n841, ZN => n12536);
   U13186 : CLKBUF_X2 port map( I => n15859, Z => n16292);
   U935 : INV_X1 port map( I => n16021, ZN => n13717);
   U5800 : INV_X1 port map( I => n577, ZN => n16041);
   U4333 : INV_X2 port map( I => n16111, ZN => n16320);
   U20356 : INV_X1 port map( I => n16258, ZN => n15607);
   U15312 : INV_X1 port map( I => n16335, ZN => n13307);
   U15108 : INV_X2 port map( I => n5580, ZN => n16132);
   U15827 : INV_X1 port map( I => n10707, ZN => n16326);
   U2502 : INV_X1 port map( I => n16131, ZN => n14636);
   U4335 : INV_X1 port map( I => n16227, ZN => n16080);
   U6812 : INV_X2 port map( I => n1269, ZN => n16148);
   U11129 : INV_X1 port map( I => n22590, ZN => n15980);
   U8272 : NOR2_X1 port map( A1 => n9095, A2 => n16321, ZN => n7007);
   U5812 : NAND2_X1 port map( A1 => n16266, A2 => n28088, ZN => n6256);
   U14499 : OAI21_X1 port map( A1 => n9967, A2 => n15970, B => n5139, ZN => 
                           n9966);
   U20220 : OAI21_X1 port map( A1 => n1264, A2 => n22910, B => n6316, ZN => 
                           n16081);
   U14010 : NAND2_X1 port map( A1 => n13677, A2 => n1269, ZN => n15935);
   U8252 : NOR2_X1 port map( A1 => n10001, A2 => n16271, ZN => n7124);
   U1707 : OAI21_X1 port map( A1 => n3797, A2 => n4114, B => n14171, ZN => 
                           n25448);
   U3124 : NAND2_X1 port map( A1 => n12116, A2 => n15998, ZN => n379);
   U6857 : INV_X1 port map( I => n10303, ZN => n16206);
   U3689 : INV_X1 port map( I => n16080, ZN => n5884);
   U21390 : NAND2_X1 port map( A1 => n15930, A2 => n1262, ZN => n7014);
   U21561 : INV_X1 port map( I => n15984, ZN => n16146);
   U5815 : INV_X1 port map( I => n21787, ZN => n16185);
   U2367 : INV_X1 port map( I => n7910, ZN => n2195);
   U1762 : NOR3_X1 port map( A1 => n12918, A2 => n798, A3 => n7266, ZN => n5381
                           );
   U3626 : BUF_X2 port map( I => n15936, Z => n516);
   U9594 : NOR2_X1 port map( A1 => n8031, A2 => n14303, ZN => n9595);
   U15692 : NOR2_X1 port map( A1 => n16220, A2 => n16253, ZN => n6605);
   U5384 : INV_X2 port map( I => n16132, ZN => n10453);
   U5787 : NOR2_X1 port map( A1 => n524, A2 => n25570, ZN => n6240);
   U16325 : NAND2_X1 port map( A1 => n16231, A2 => n16072, ZN => n15676);
   U8275 : INV_X1 port map( I => n5139, ZN => n6837);
   U8170 : NOR2_X1 port map( A1 => n16299, A2 => n16189, ZN => n6192);
   U19270 : NAND2_X1 port map( A1 => n795, A2 => n14442, ZN => n23908);
   U20847 : NAND2_X1 port map( A1 => n16063, A2 => n16062, ZN => n2543);
   U1662 : AOI22_X1 port map( A1 => n3232, A2 => n16267, B1 => n5884, B2 => 
                           n5744, ZN => n26280);
   U6773 : NAND2_X1 port map( A1 => n1264, A2 => n6256, ZN => n6255);
   U14188 : NAND2_X1 port map( A1 => n15925, A2 => n16136, ZN => n25471);
   U924 : NOR2_X1 port map( A1 => n15676, A2 => n21904, ZN => n16092);
   U10522 : AOI21_X1 port map( A1 => n15928, A2 => n15980, B => n10453, ZN => 
                           n8085);
   U18009 : NAND2_X1 port map( A1 => n16299, A2 => n13430, ZN => n14732);
   U8190 : NAND2_X1 port map( A1 => n6315, A2 => n16267, ZN => n6257);
   U10449 : NAND2_X1 port map( A1 => n24198, A2 => n24485, ZN => n6729);
   U16400 : NAND2_X1 port map( A1 => n7868, A2 => n16069, ZN => n14012);
   U5767 : NOR2_X1 port map( A1 => n1268, A2 => n914, ZN => n2629);
   U10451 : INV_X1 port map( I => n16122, ZN => n2147);
   U14867 : NOR2_X1 port map( A1 => n14830, A2 => n6304, ZN => n6303);
   U1687 : NAND2_X1 port map( A1 => n1271, A2 => n14178, ZN => n10870);
   U6791 : NAND2_X1 port map( A1 => n9393, A2 => n5853, ZN => n10037);
   U19629 : NAND2_X1 port map( A1 => n15874, A2 => n21764, ZN => n14067);
   U13872 : NAND2_X1 port map( A1 => n5312, A2 => n25657, ZN => n25426);
   U1239 : NAND2_X1 port map( A1 => n16086, A2 => n21873, ZN => n22975);
   U20492 : NOR2_X1 port map( A1 => n838, A2 => n14636, ZN => n15841);
   U10406 : INV_X1 port map( I => n16016, ZN => n16019);
   U3057 : OAI21_X1 port map( A1 => n16147, A2 => n11429, B => n16146, ZN => 
                           n15511);
   U2489 : AOI22_X1 port map( A1 => n9704, A2 => n16063, B1 => n22798, B2 => 
                           n7053, ZN => n25728);
   U5066 : NOR2_X1 port map( A1 => n25225, A2 => n5050, ZN => n5052);
   U5367 : OAI22_X1 port map( A1 => n15971, A2 => n6317, B1 => n16080, B2 => 
                           n6316, ZN => n22984);
   U2067 : AOI21_X1 port map( A1 => n16022, A2 => n16144, B => n26350, ZN => 
                           n14881);
   U5765 : AOI22_X1 port map( A1 => n2629, A2 => n797, B1 => n15953, B2 => 
                           n1268, ZN => n2627);
   U1019 : OAI21_X1 port map( A1 => n16298, A2 => n6480, B => n6477, ZN => 
                           n6476);
   U6779 : NAND2_X1 port map( A1 => n4942, A2 => n12678, ZN => n8498);
   U17319 : OAI21_X1 port map( A1 => n15840, A2 => n15841, B => n8303, ZN => 
                           n25911);
   U5231 : BUF_X4 port map( I => n3792, Z => n25940);
   U21819 : NAND3_X1 port map( A1 => n16303, A2 => n25017, A3 => n14107, ZN => 
                           n10609);
   U1147 : BUF_X2 port map( I => n7308, Z => n1793);
   U9607 : BUF_X2 port map( I => n16610, Z => n24167);
   U14147 : OR2_X1 port map( A1 => n15942, A2 => n25657, Z => n4645);
   U2245 : INV_X2 port map( I => n12637, ZN => n8199);
   U6708 : INV_X1 port map( I => n16525, ZN => n1246);
   U18040 : NAND2_X1 port map( A1 => n434, A2 => n27239, ZN => n13298);
   U880 : CLKBUF_X2 port map( I => n13415, Z => n7378);
   U12149 : INV_X1 port map( I => n5874, ZN => n2149);
   U2555 : INV_X2 port map( I => n3914, ZN => n16605);
   U16459 : INV_X1 port map( I => n10337, ZN => n7688);
   U19618 : NOR2_X1 port map( A1 => n16530, A2 => n23842, ZN => n26241);
   U3486 : INV_X1 port map( I => n16597, ZN => n16638);
   U14177 : NOR2_X1 port map( A1 => n16694, A2 => n27734, ZN => n5438);
   U5052 : NOR2_X1 port map( A1 => n5197, A2 => n24829, ZN => n14626);
   U11915 : AOI21_X1 port map( A1 => n912, A2 => n26169, B => n2481, ZN => 
                           n2765);
   U3508 : NAND2_X1 port map( A1 => n16422, A2 => n16685, ZN => n25995);
   U10234 : INV_X1 port map( I => n16551, ZN => n11144);
   U16737 : INV_X1 port map( I => n124, ZN => n8021);
   U8037 : INV_X1 port map( I => n7395, ZN => n16523);
   U11050 : INV_X2 port map( I => n22572, ZN => n10597);
   U1553 : OAI21_X1 port map( A1 => n2607, A2 => n11721, B => n25199, ZN => 
                           n5710);
   U19299 : INV_X1 port map( I => n8722, ZN => n26187);
   U10732 : INV_X2 port map( I => n23907, ZN => n7113);
   U19765 : NAND2_X1 port map( A1 => n13298, A2 => n16519, ZN => n26258);
   U1185 : NAND2_X1 port map( A1 => n7668, A2 => n16497, ZN => n16573);
   U4297 : CLKBUF_X2 port map( I => n9773, Z => n9202);
   U1588 : NAND2_X1 port map( A1 => n9759, A2 => n12117, ZN => n14908);
   U2439 : NOR2_X1 port map( A1 => n10282, A2 => n14632, ZN => n25736);
   U13629 : INV_X2 port map( I => n2179, ZN => n4556);
   U17133 : INV_X1 port map( I => n16644, ZN => n16736);
   U4267 : BUF_X2 port map( I => n9978, Z => n9917);
   U10276 : NOR2_X1 port map( A1 => n1054, A2 => n12647, ZN => n15613);
   U1963 : INV_X1 port map( I => n12292, ZN => n7539);
   U21185 : NAND2_X1 port map( A1 => n4644, A2 => n5874, ZN => n6538);
   U13943 : INV_X1 port map( I => n14228, ZN => n13572);
   U2129 : INV_X1 port map( I => n6843, ZN => n741);
   U4649 : INV_X1 port map( I => n25940, ZN => n10261);
   U855 : INV_X1 port map( I => n13739, ZN => n1251);
   U1570 : NAND2_X1 port map( A1 => n7964, A2 => n8722, ZN => n7531);
   U13955 : NOR2_X1 port map( A1 => n703, A2 => n1054, ZN => n16057);
   U8068 : NAND2_X1 port map( A1 => n16647, A2 => n5244, ZN => n3551);
   U2499 : OAI22_X1 port map( A1 => n13211, A2 => n27381, B1 => n741, B2 => 
                           n6838, ZN => n9315);
   U1593 : AOI21_X1 port map( A1 => n3017, A2 => n24341, B => n25670, ZN => 
                           n25197);
   U10297 : NAND2_X1 port map( A1 => n16700, A2 => n3443, ZN => n4296);
   U10279 : NAND2_X1 port map( A1 => n907, A2 => n25199, ZN => n2060);
   U8097 : NAND2_X1 port map( A1 => n14401, A2 => n16644, ZN => n6048);
   U5043 : NAND2_X1 port map( A1 => n14676, A2 => n16507, ZN => n8916);
   U2992 : OAI21_X1 port map( A1 => n16609, A2 => n23935, B => n1048, ZN => 
                           n1981);
   U8024 : NAND2_X1 port map( A1 => n16679, A2 => n15652, ZN => n14309);
   U7995 : NAND3_X1 port map( A1 => n14579, A2 => n14264, A3 => n16523, ZN => 
                           n9372);
   U9147 : OAI21_X1 port map( A1 => n26240, A2 => n26241, B => n13927, ZN => 
                           n24975);
   U8122 : NOR2_X1 port map( A1 => n132, A2 => n26105, ZN => n10567);
   U15744 : NOR2_X1 port map( A1 => n25698, A2 => n5442, ZN => n21809);
   U10266 : NAND2_X1 port map( A1 => n2045, A2 => n12039, ZN => n6879);
   U4826 : INV_X1 port map( I => n16400, ZN => n7957);
   U21678 : INV_X2 port map( I => n4281, ZN => n26463);
   U5417 : INV_X2 port map( I => n12949, ZN => n26114);
   U8085 : NOR2_X1 port map( A1 => n6347, A2 => n7180, ZN => n15120);
   U5750 : NOR2_X1 port map( A1 => n24845, A2 => n22061, ZN => n10142);
   U15985 : NAND2_X1 port map( A1 => n25995, A2 => n25731, ZN => n15880);
   U5388 : NOR2_X1 port map( A1 => n26169, A2 => n27734, ZN => n25583);
   U18173 : BUF_X2 port map( I => n16649, Z => n26039);
   U17254 : NAND2_X1 port map( A1 => n28141, A2 => n23474, ZN => n16667);
   U20645 : NAND2_X1 port map( A1 => n24089, A2 => n5197, ZN => n16670);
   U8066 : OAI21_X1 port map( A1 => n15536, A2 => n28231, B => n16681, ZN => 
                           n3552);
   U5362 : INV_X2 port map( I => n16530, ZN => n793);
   U4498 : INV_X1 port map( I => n16640, ZN => n16598);
   U5042 : INV_X1 port map( I => n16391, ZN => n16408);
   U891 : INV_X2 port map( I => n8534, ZN => n8530);
   U1191 : NAND2_X1 port map( A1 => n14177, A2 => n3479, ZN => n24484);
   U7031 : OR2_X1 port map( A1 => n5442, A2 => n16612, Z => n16614);
   U6267 : AND2_X1 port map( A1 => n24236, A2 => n16630, Z => n24650);
   U1138 : INV_X1 port map( I => n24727, ZN => n24374);
   U8081 : NOR2_X1 port map( A1 => n6688, A2 => n2045, ZN => n1647);
   U19462 : INV_X2 port map( I => n16471, ZN => n16555);
   U12933 : AOI22_X1 port map( A1 => n9830, A2 => n13572, B1 => n13964, B2 => 
                           n13927, ZN => n1504);
   U1478 : NOR3_X1 port map( A1 => n25772, A2 => n1251, A3 => n16336, ZN => 
                           n25902);
   U15092 : OAI22_X1 port map( A1 => n16556, A2 => n4940, B1 => n16554, B2 => 
                           n16555, ZN => n14270);
   U9698 : NAND2_X1 port map( A1 => n16611, A2 => n14562, ZN => n15418);
   U6692 : AOI21_X1 port map( A1 => n16732, A2 => n13496, B => n9484, ZN => 
                           n9483);
   U12777 : NAND2_X1 port map( A1 => n16647, A2 => n24727, ZN => n14802);
   U5762 : OAI21_X1 port map( A1 => n14165, A2 => n25670, B => n14339, ZN => 
                           n2723);
   U5725 : AOI21_X1 port map( A1 => n14254, A2 => n9830, B => n793, ZN => n1503
                           );
   U1082 : OAI21_X1 port map( A1 => n7957, A2 => n16399, B => n9830, ZN => 
                           n11599);
   U10304 : NAND2_X1 port map( A1 => n16476, A2 => n13608, ZN => n16478);
   U11192 : NOR2_X1 port map( A1 => n23719, A2 => n22542, ZN => n1750);
   U7204 : NAND2_X1 port map( A1 => n12949, A2 => n16707, ZN => n16708);
   U8109 : NAND2_X1 port map( A1 => n2045, A2 => n10304, ZN => n6684);
   U19978 : AOI21_X1 port map( A1 => n9907, A2 => n8530, B => n2789, ZN => 
                           n9522);
   U1806 : NOR2_X1 port map( A1 => n1247, A2 => n2789, ZN => n16363);
   U10267 : INV_X1 port map( I => n16481, ZN => n2248);
   U17882 : AOI21_X1 port map( A1 => n16409, A2 => n26039, B => n14173, ZN => 
                           n14172);
   U6684 : AOI21_X1 port map( A1 => n3196, A2 => n16467, B => n16700, ZN => 
                           n16470);
   U20698 : NOR2_X1 port map( A1 => n24845, A2 => n8097, ZN => n24141);
   U11933 : NAND2_X1 port map( A1 => n22715, A2 => n23439, ZN => n123);
   U13365 : INV_X1 port map( I => n25670, ZN => n904);
   U10268 : NAND2_X1 port map( A1 => n3552, A2 => n3551, ZN => n9870);
   U1515 : OAI21_X1 port map( A1 => n8511, A2 => n16696, B => n7963, ZN => 
                           n8295);
   U12905 : NOR2_X1 port map( A1 => n16669, A2 => n8534, ZN => n15538);
   U15118 : NOR2_X1 port map( A1 => n1595, A2 => n23809, ZN => n25619);
   U2079 : NAND2_X1 port map( A1 => n2060, A2 => n3017, ZN => n120);
   U1737 : INV_X2 port map( I => n5718, ZN => n902);
   U14427 : NAND2_X1 port map( A1 => n25501, A2 => n16660, ZN => n24426);
   U17877 : NOR2_X1 port map( A1 => n28231, A2 => n15239, ZN => n13214);
   U15114 : NOR2_X1 port map( A1 => n4281, A2 => n5244, ZN => n13215);
   U11200 : NOR2_X1 port map( A1 => n1048, A2 => n5874, ZN => n25195);
   U823 : OAI22_X1 port map( A1 => n16614, A2 => n16615, B1 => n6147, B2 => 
                           n1243, ZN => n254);
   U19103 : INV_X1 port map( I => n16853, ZN => n22358);
   U7976 : OAI22_X1 port map( A1 => n10514, A2 => n1242, B1 => n16421, B2 => 
                           n23758, ZN => n7356);
   U7944 : OAI21_X1 port map( A1 => n13309, A2 => n7323, B => n3751, ZN => 
                           n1919);
   U10162 : INV_X1 port map( I => n11143, ZN => n10189);
   U9989 : AOI21_X1 port map( A1 => n16611, A2 => n23236, B => n910, ZN => 
                           n6131);
   U10151 : NAND2_X1 port map( A1 => n5240, A2 => n16812, ZN => n3428);
   U10259 : NAND2_X1 port map( A1 => n2723, A2 => n729, ZN => n2722);
   U7992 : OAI21_X1 port map( A1 => n6812, A2 => n16418, B => n25359, ZN => 
                           n6400);
   U10131 : NAND2_X1 port map( A1 => n24347, A2 => n17117, ZN => n1920);
   U1096 : OAI21_X1 port map( A1 => n6402, A2 => n6403, B => n16679, ZN => 
                           n22252);
   U14788 : AOI22_X1 port map( A1 => n8363, A2 => n904, B1 => n24650, B2 => 
                           n24215, ZN => n25553);
   U20216 : AOI21_X1 port map( A1 => n26318, A2 => n10425, B => n24770, ZN => 
                           n10423);
   U13869 : NAND2_X1 port map( A1 => n7877, A2 => n7466, ZN => n25425);
   U18864 : NAND3_X1 port map( A1 => n13496, A2 => n835, A3 => n28126, ZN => 
                           n13495);
   U12298 : NAND3_X1 port map( A1 => n16669, A2 => n16667, A3 => n2789, ZN => 
                           n23896);
   U13061 : NOR2_X1 port map( A1 => n16569, A2 => n16568, ZN => n16845);
   U4515 : OAI21_X1 port map( A1 => n24583, A2 => n465, B => n16760, ZN => 
                           n15637);
   U1483 : NAND2_X1 port map( A1 => n5684, A2 => n16544, ZN => n25337);
   U4534 : CLKBUF_X2 port map( I => n12626, Z => n452);
   U20074 : OAI21_X1 port map( A1 => n15061, A2 => n16681, B => n4281, ZN => 
                           n24066);
   U2668 : INV_X1 port map( I => n26246, ZN => n22597);
   U5141 : INV_X1 port map( I => n17032, ZN => n25029);
   U2185 : INV_X1 port map( I => n17133, ZN => n6101);
   U18402 : NAND2_X1 port map( A1 => n5684, A2 => n16544, ZN => n12709);
   U4382 : INV_X1 port map( I => n7362, ZN => n22673);
   U6840 : INV_X1 port map( I => n14574, ZN => n1273);
   U13831 : NAND2_X1 port map( A1 => n1920, A2 => n1919, ZN => n16932);
   U2985 : CLKBUF_X2 port map( I => n7786, Z => n24000);
   U3454 : INV_X1 port map( I => n7257, ZN => n11794);
   U811 : INV_X1 port map( I => n9027, ZN => n8880);
   U6140 : INV_X1 port map( I => n20519, ZN => n21281);
   U5146 : INV_X1 port map( I => n13443, ZN => n25785);
   U18198 : INV_X1 port map( I => n7973, ZN => n17044);
   U7947 : INV_X1 port map( I => n2265, ZN => n17069);
   U15254 : INV_X1 port map( I => n10999, ZN => n14999);
   U6137 : BUF_X2 port map( I => Key(101), Z => n21262);
   U5124 : INV_X1 port map( I => n16981, ZN => n24956);
   U7943 : INV_X1 port map( I => n16820, ZN => n16916);
   U4378 : INV_X1 port map( I => n20652, ZN => n22512);
   U16761 : INV_X1 port map( I => n9399, ZN => n17033);
   U4542 : INV_X1 port map( I => n12691, ZN => n7988);
   U20262 : INV_X2 port map( I => n15190, ZN => n17489);
   U3475 : INV_X1 port map( I => n360, ZN => n9018);
   U772 : INV_X1 port map( I => n17157, ZN => n1892);
   U3794 : BUF_X2 port map( I => n1565, Z => n24566);
   U16548 : INV_X1 port map( I => n26615, ZN => n17526);
   U12459 : NOR2_X1 port map( A1 => n17501, A2 => n17346, ZN => n23723);
   U9283 : NOR2_X1 port map( A1 => n6185, A2 => n24566, ZN => n25206);
   U12458 : NOR2_X1 port map( A1 => n17501, A2 => n899, ZN => n1940);
   U5106 : BUF_X2 port map( I => n17463, Z => n14357);
   U2765 : INV_X2 port map( I => n3090, ZN => n17166);
   U19318 : BUF_X2 port map( I => n28537, Z => n23926);
   U2363 : NAND2_X1 port map( A1 => n9358, A2 => n14324, ZN => n22399);
   U10750 : INV_X2 port map( I => n10209, ZN => n8692);
   U5479 : INV_X1 port map( I => n542, ZN => n17543);
   U5317 : INV_X2 port map( I => n6637, ZN => n791);
   U17122 : INV_X1 port map( I => n8995, ZN => n8996);
   U20738 : INV_X1 port map( I => n17302, ZN => n17192);
   U15885 : INV_X1 port map( I => n17446, ZN => n17547);
   U5718 : INV_X2 port map( I => n17230, ZN => n17558);
   U1442 : NOR2_X1 port map( A1 => n17244, A2 => n13693, ZN => n17213);
   U1435 : INV_X2 port map( I => n17519, ZN => n26226);
   U16372 : NOR3_X1 port map( A1 => n17381, A2 => n21785, A3 => n17548, ZN => 
                           n7433);
   U18460 : INV_X2 port map( I => n23269, ZN => n17561);
   U19413 : OAI21_X1 port map( A1 => n17415, A2 => n5500, B => n1030, ZN => 
                           n26217);
   U12104 : INV_X1 port map( I => n10183, ZN => n14697);
   U3702 : INV_X2 port map( I => n9898, ZN => n897);
   U13669 : NOR2_X1 port map( A1 => n15189, A2 => n6672, ZN => n6663);
   U9992 : OAI21_X1 port map( A1 => n830, A2 => n4536, B => n26655, ZN => n6662
                           );
   U17231 : INV_X1 port map( I => n9224, ZN => n10568);
   U19714 : NOR2_X1 port map( A1 => n24018, A2 => n1040, ZN => n24017);
   U3488 : NAND2_X1 port map( A1 => n14963, A2 => n17166, ZN => n476);
   U11974 : NOR2_X1 port map( A1 => n11761, A2 => n10942, ZN => n25280);
   U1450 : INV_X2 port map( I => n12692, ZN => n15504);
   U16745 : NAND2_X1 port map( A1 => n17219, A2 => n8180, ZN => n15122);
   U5685 : NOR2_X1 port map( A1 => n17335, A2 => n7361, ZN => n7620);
   U2570 : INV_X2 port map( I => n17403, ZN => n8473);
   U3361 : CLKBUF_X1 port map( I => n9224, Z => n461);
   U5536 : BUF_X2 port map( I => n5541, Z => n26213);
   U1742 : NOR2_X1 port map( A1 => n23723, A2 => n23724, ZN => n26287);
   U4633 : INV_X2 port map( I => n17492, ZN => n9569);
   U4635 : INV_X1 port map( I => n900, ZN => n1231);
   U2217 : INV_X1 port map( I => n12340, ZN => n13568);
   U720 : INV_X2 port map( I => n10150, ZN => n17370);
   U12568 : NOR2_X1 port map( A1 => n24560, A2 => n14944, ZN => n25672);
   U1935 : NAND2_X1 port map( A1 => n17522, A2 => n900, ZN => n2934);
   U745 : INV_X2 port map( I => n23926, ZN => n790);
   U5692 : INV_X2 port map( I => n791, ZN => n15737);
   U16138 : OR2_X1 port map( A1 => n6637, A2 => n15344, Z => n17483);
   U1059 : AND2_X1 port map( A1 => n15273, A2 => n5506, Z => n14504);
   U750 : INV_X1 port map( I => n28538, ZN => n12882);
   U5507 : INV_X1 port map( I => n10942, ZN => n17390);
   U19010 : CLKBUF_X2 port map( I => n7269, Z => n26161);
   U2481 : BUF_X2 port map( I => n11610, Z => n8093);
   U1448 : INV_X1 port map( I => n766, ZN => n8435);
   U6619 : INV_X1 port map( I => n17343, ZN => n2527);
   U6188 : OR2_X1 port map( A1 => n14997, A2 => n540, Z => n24613);
   U10035 : NAND2_X1 port map( A1 => n2934, A2 => n12748, ZN => n6342);
   U5572 : NAND3_X1 port map( A1 => n17177, A2 => n16999, A3 => n17175, ZN => 
                           n17000);
   U17763 : NOR2_X1 port map( A1 => n4797, A2 => n14592, ZN => n12641);
   U7877 : NAND2_X1 port map( A1 => n13509, A2 => n8093, ZN => n5416);
   U11219 : NAND2_X1 port map( A1 => n17510, A2 => n24585, ZN => n23040);
   U13588 : NAND3_X1 port map( A1 => n23275, A2 => n17478, A3 => n25608, ZN => 
                           n13356);
   U1003 : NAND3_X1 port map( A1 => n17518, A2 => n7996, A3 => n24323, ZN => 
                           n630);
   U6592 : AOI21_X1 port map( A1 => n17524, A2 => n11761, B => n791, ZN => 
                           n5254);
   U15496 : NAND2_X1 port map( A1 => n17400, A2 => n23556, ZN => n13637);
   U1400 : NAND2_X1 port map( A1 => n4415, A2 => n14453, ZN => n25215);
   U3843 : INV_X2 port map( I => n10603, ZN => n894);
   U6552 : OAI21_X1 port map( A1 => n1030, A2 => n9132, B => n27132, ZN => 
                           n1950);
   U4585 : NAND2_X1 port map( A1 => n26852, A2 => n17514, ZN => n17203);
   U7355 : NOR2_X1 port map( A1 => n17460, A2 => n17408, ZN => n24779);
   U4592 : NOR2_X1 port map( A1 => n17436, A2 => n9661, ZN => n17437);
   U14814 : NOR2_X1 port map( A1 => n17472, A2 => n17541, ZN => n25561);
   U16420 : NOR2_X1 port map( A1 => n17534, A2 => n17541, ZN => n23471);
   U18058 : NOR2_X1 port map( A1 => n831, A2 => n26161, ZN => n12496);
   U5032 : INV_X1 port map( I => n26349, ZN => n12485);
   U1218 : INV_X1 port map( I => n17402, ZN => n10972);
   U4142 : NAND2_X1 port map( A1 => n13535, A2 => n24159, ZN => n24103);
   U10744 : NAND3_X1 port map( A1 => n6258, A2 => n25140, A3 => n17362, ZN => 
                           n6966);
   U4478 : INV_X1 port map( I => n7370, ZN => n17527);
   U5019 : NAND3_X1 port map( A1 => n790, A2 => n26418, A3 => n13740, ZN => 
                           n4463);
   U14447 : NOR2_X1 port map( A1 => n6022, A2 => n1227, ZN => n7797);
   U15077 : NOR2_X1 port map( A1 => n1036, A2 => n13070, ZN => n7096);
   U15937 : INV_X1 port map( I => n17163, ZN => n17162);
   U5436 : BUF_X2 port map( I => n17230, Z => n17496);
   U5313 : INV_X1 port map( I => n10081, ZN => n1229);
   U21630 : NOR3_X1 port map( A1 => n8094, A2 => n10046, A3 => n1227, ZN => 
                           n5375);
   U13507 : NAND3_X1 port map( A1 => n7357, A2 => n791, A3 => n17525, ZN => 
                           n13880);
   U4480 : NAND3_X1 port map( A1 => n25504, A2 => n17492, A3 => n8125, ZN => 
                           n10182);
   U20793 : NOR2_X1 port map( A1 => n14592, A2 => n27073, ZN => n17476);
   U6569 : NAND2_X1 port map( A1 => n4254, A2 => n4888, ZN => n4253);
   U17751 : NOR2_X1 port map( A1 => n8996, A2 => n10875, ZN => n11716);
   U13013 : NOR2_X1 port map( A1 => n17306, A2 => n17301, ZN => n11674);
   U9102 : NOR2_X1 port map( A1 => n6293, A2 => n17463, ZN => n8335);
   U739 : INV_X1 port map( I => n11763, ZN => n17417);
   U1375 : NOR2_X1 port map( A1 => n3980, A2 => n6977, ZN => n17216);
   U6575 : INV_X2 port map( I => n17569, ZN => n1032);
   U1288 : INV_X1 port map( I => n9879, ZN => n17314);
   U10075 : INV_X1 port map( I => n17570, ZN => n1566);
   U16040 : OR2_X1 port map( A1 => n15514, A2 => n8430, Z => n9651);
   U5514 : INV_X1 port map( I => n2037, ZN => n372);
   U18454 : NOR2_X1 port map( A1 => n17486, A2 => n17561, ZN => n17488);
   U21671 : NOR2_X1 port map( A1 => n17230, A2 => n17556, ZN => n17223);
   U21722 : INV_X2 port map( I => n15077, ZN => n24387);
   U10085 : AOI21_X1 port map( A1 => n17317, A2 => n27288, B => n8692, ZN => 
                           n5016);
   U1825 : OAI21_X1 port map( A1 => n17227, A2 => n899, B => n17577, ZN => 
                           n17228);
   U4629 : NAND3_X1 port map( A1 => n17166, A2 => n24159, A3 => n17418, ZN => 
                           n3092);
   U1040 : NAND2_X1 port map( A1 => n17510, A2 => n7275, ZN => n7033);
   U1362 : AOI21_X1 port map( A1 => n17370, A2 => n10577, B => n17372, ZN => 
                           n23852);
   U2123 : AOI21_X1 port map( A1 => n17175, A2 => n2963, B => n17307, ZN => 
                           n17308);
   U1452 : OAI21_X1 port map( A1 => n15737, A2 => n15504, B => n17525, ZN => 
                           n11171);
   U17899 : NAND2_X1 port map( A1 => n27648, A2 => n17452, ZN => n12707);
   U7860 : NOR2_X1 port map( A1 => n6672, A2 => n17489, ZN => n13268);
   U9471 : NAND2_X1 port map( A1 => n17347, A2 => n24091, ZN => n3786);
   U10040 : NOR2_X1 port map( A1 => n4415, A2 => n17496, ZN => n9089);
   U8256 : AOI21_X1 port map( A1 => n17365, A2 => n17364, B => n25786, ZN => 
                           n24882);
   U1353 : AOI21_X1 port map( A1 => n17192, A2 => n24688, B => n17177, ZN => 
                           n24752);
   U9942 : AOI21_X1 port map( A1 => n16743, A2 => n9593, B => n15063, ZN => 
                           n11532);
   U4630 : NAND2_X1 port map( A1 => n17437, A2 => n4715, ZN => n1883);
   U9973 : NAND2_X1 port map( A1 => n6342, A2 => n17427, ZN => n15722);
   U2375 : OAI21_X1 port map( A1 => n1030, A2 => n5500, B => n17415, ZN => n184
                           );
   U7783 : NAND3_X1 port map( A1 => n17433, A2 => n24513, A3 => n17436, ZN => 
                           n24273);
   U9888 : OAI21_X1 port map( A1 => n7797, A2 => n9556, B => n896, ZN => n5958)
                           ;
   U9982 : AOI21_X1 port map( A1 => n17265, A2 => n5612, B => n17426, ZN => 
                           n2753);
   U6788 : NOR2_X1 port map( A1 => n12641, A2 => n17280, ZN => n25107);
   U9883 : AOI21_X1 port map( A1 => n9555, A2 => n6022, B => n5078, ZN => n5959
                           );
   U1033 : CLKBUF_X2 port map( I => n17185, Z => n23787);
   U19979 : NOR2_X1 port map( A1 => n24059, A2 => n5563, ZN => n5562);
   U14206 : NAND2_X1 port map( A1 => n4715, A2 => n27341, ZN => n11327);
   U15462 : AOI21_X1 port map( A1 => n27946, A2 => n27530, B => n764, ZN => 
                           n13281);
   U1364 : INV_X1 port map( I => n17337, ZN => n17735);
   U6567 : NOR2_X1 port map( A1 => n832, A2 => n8692, ZN => n5257);
   U6522 : AOI21_X1 port map( A1 => n1036, A2 => n24406, B => n16872, ZN => 
                           n16880);
   U2531 : AOI22_X1 port map( A1 => n9609, A2 => n14900, B1 => n4472, B2 => 
                           n11284, ZN => n9608);
   U7859 : OAI21_X1 port map( A1 => n27161, A2 => n1234, B => n25013, ZN => 
                           n6197);
   U13803 : NAND2_X1 port map( A1 => n5016, A2 => n832, ZN => n5015);
   U20792 : NAND2_X1 port map( A1 => n17464, A2 => n9898, ZN => n17465);
   U5629 : OAI21_X1 port map( A1 => n27580, A2 => n2963, B => n17308, ZN => 
                           n17309);
   U13589 : NAND2_X1 port map( A1 => n8986, A2 => n25608, ZN => n4799);
   U13717 : NOR2_X1 port map( A1 => n17464, A2 => n9898, ZN => n25406);
   U2374 : OAI21_X1 port map( A1 => n17287, A2 => n17415, B => n184, ZN => 
                           n17290);
   U9955 : NAND2_X1 port map( A1 => n23327, A2 => n17558, ZN => n25077);
   U7866 : OAI21_X1 port map( A1 => n8692, A2 => n17318, B => n17401, ZN => 
                           n17022);
   U989 : NAND3_X1 port map( A1 => n12707, A2 => n12706, A3 => n11992, ZN => 
                           n6484);
   U7234 : INV_X2 port map( I => n15462, ZN => n22519);
   U14542 : NAND3_X1 port map( A1 => n5187, A2 => n13779, A3 => n28535, ZN => 
                           n10566);
   U1634 : NAND2_X1 port map( A1 => n25796, A2 => n13282, ZN => n13499);
   U975 : NOR2_X1 port map( A1 => n11216, A2 => n11217, ZN => n22817);
   U5591 : INV_X1 port map( I => n17976, ZN => n15539);
   U5010 : INV_X1 port map( I => n17617, ZN => n17678);
   U16714 : OAI21_X1 port map( A1 => n23979, A2 => n17962, B => n11182, ZN => 
                           n25837);
   U16192 : INV_X2 port map( I => n17665, ZN => n728);
   U9851 : NAND2_X1 port map( A1 => n17607, A2 => n18005, ZN => n11818);
   U12403 : NAND2_X1 port map( A1 => n10133, A2 => n17942, ZN => n12312);
   U3395 : INV_X1 port map( I => n17953, ZN => n25530);
   U629 : INV_X1 port map( I => n5955, ZN => n5957);
   U9722 : NOR2_X1 port map( A1 => n14552, A2 => n17872, ZN => n12791);
   U11983 : INV_X2 port map( I => n7321, ZN => n14284);
   U674 : INV_X2 port map( I => n283, ZN => n17845);
   U3316 : BUF_X2 port map( I => n6018, Z => n24316);
   U4087 : CLKBUF_X2 port map( I => n14269, Z => n21943);
   U675 : INV_X2 port map( I => n6910, ZN => n4475);
   U5509 : INV_X2 port map( I => n11182, ZN => n9905);
   U17806 : BUF_X2 port map( I => n10779, Z => n23696);
   U860 : INV_X1 port map( I => n17935, ZN => n24397);
   U668 : INV_X2 port map( I => n13530, ZN => n826);
   U937 : INV_X2 port map( I => n23118, ZN => n10673);
   U977 : INV_X1 port map( I => n10779, ZN => n22153);
   U12791 : INV_X1 port map( I => n8155, ZN => n14986);
   U5376 : INV_X2 port map( I => n11112, ZN => n6629);
   U11385 : NAND2_X1 port map( A1 => n17927, A2 => n4813, ZN => n12429);
   U17417 : INV_X1 port map( I => n9691, ZN => n13329);
   U12708 : NAND2_X1 port map( A1 => n5584, A2 => n17607, ZN => n17608);
   U16397 : NOR2_X1 port map( A1 => n24304, A2 => n17881, ZN => n7496);
   U5268 : NAND2_X1 port map( A1 => n11182, A2 => n17761, ZN => n17764);
   U1316 : NAND2_X1 port map( A1 => n17687, A2 => n22646, ZN => n15098);
   U20810 : INV_X1 port map( I => n18002, ZN => n17842);
   U1949 : NAND2_X1 port map( A1 => n21898, A2 => n23110, ZN => n13208);
   U4981 : INV_X2 port map( I => n9285, ZN => n1022);
   U13265 : INV_X2 port map( I => n14446, ZN => n17925);
   U4295 : INV_X1 port map( I => n17580, ZN => n17920);
   U3321 : BUF_X2 port map( I => n17919, Z => n22244);
   U12559 : NOR2_X1 port map( A1 => n7823, A2 => n6709, ZN => n7822);
   U5627 : NOR2_X1 port map( A1 => n7023, A2 => n9606, ZN => n7178);
   U2970 : NAND2_X1 port map( A1 => n22812, A2 => n22253, ZN => n23469);
   U656 : INV_X1 port map( I => n17722, ZN => n789);
   U3052 : INV_X2 port map( I => n891, ZN => n17830);
   U666 : INV_X2 port map( I => n11579, ZN => n8365);
   U877 : NOR2_X1 port map( A1 => n8070, A2 => n6709, ZN => n8071);
   U11303 : NAND2_X1 port map( A1 => n26356, A2 => n1893, ZN => n13547);
   U19368 : NOR2_X1 port map( A1 => n23963, A2 => n14255, ZN => n7821);
   U2658 : BUF_X2 port map( I => n11968, Z => n23706);
   U5659 : INV_X2 port map( I => n1211, ZN => n1020);
   U18612 : INV_X1 port map( I => n17943, ZN => n23811);
   U2968 : BUF_X2 port map( I => n283, Z => n24391);
   U18293 : NAND2_X1 port map( A1 => n12312, A2 => n24916, ZN => n12311);
   U1319 : BUF_X2 port map( I => n17953, Z => n24175);
   U4094 : INV_X2 port map( I => n23110, ZN => n885);
   U4471 : INV_X1 port map( I => n9734, ZN => n10030);
   U3437 : NAND2_X1 port map( A1 => n28105, A2 => n27640, ZN => n25002);
   U11773 : INV_X2 port map( I => n25856, ZN => n9040);
   U1805 : INV_X2 port map( I => n25697, ZN => n25144);
   U1223 : AND2_X1 port map( A1 => n17935, A2 => n17824, Z => n24586);
   U4457 : INV_X2 port map( I => n11937, ZN => n4828);
   U6764 : NAND3_X1 port map( A1 => n891, A2 => n18101, A3 => n22396, ZN => 
                           n5956);
   U634 : INV_X1 port map( I => n17868, ZN => n716);
   U11772 : NAND2_X1 port map( A1 => n9905, A2 => n17761, ZN => n25263);
   U4464 : INV_X1 port map( I => n17470, ZN => n17713);
   U13029 : OAI21_X1 port map( A1 => n17830, A2 => n7247, B => n8220, ZN => 
                           n8219);
   U5607 : INV_X1 port map( I => n10673, ZN => n17958);
   U11035 : OAI21_X1 port map( A1 => n789, A2 => n11112, B => n1617, ZN => 
                           n2221);
   U7723 : NOR2_X1 port map( A1 => n28118, A2 => n12964, ZN => n12086);
   U4658 : NAND2_X1 port map( A1 => n13237, A2 => n21792, ZN => n8502);
   U18761 : NOR2_X1 port map( A1 => n17963, A2 => n24142, ZN => n11129);
   U624 : INV_X1 port map( I => n12670, ZN => n17874);
   U7766 : NOR2_X1 port map( A1 => n4976, A2 => n27640, ZN => n4973);
   U4799 : NAND2_X1 port map( A1 => n17964, A2 => n9905, ZN => n7153);
   U20753 : NOR2_X1 port map( A1 => n17924, A2 => n4812, ZN => n17256);
   U19353 : NOR2_X1 port map( A1 => n1200, A2 => n13061, ZN => n26194);
   U7671 : AOI21_X1 port map( A1 => n887, A2 => n9105, B => n11937, ZN => 
                           n11938);
   U3119 : NAND2_X1 port map( A1 => n7023, A2 => n17751, ZN => n17159);
   U6453 : NAND2_X1 port map( A1 => n17812, A2 => n23110, ZN => n6482);
   U836 : BUF_X2 port map( I => n17941, Z => n23927);
   U6423 : NAND2_X1 port map( A1 => n21905, A2 => n9105, ZN => n9109);
   U12272 : NOR2_X1 port map( A1 => n17349, A2 => n890, ZN => n2206);
   U15364 : OAI21_X1 port map( A1 => n10178, A2 => n17816, B => n21778, ZN => 
                           n25641);
   U1269 : NOR2_X1 port map( A1 => n1219, A2 => n23391, ZN => n4591);
   U6469 : NOR2_X1 port map( A1 => n12611, A2 => n17986, ZN => n3288);
   U7666 : INV_X1 port map( I => n17742, ZN => n17743);
   U2966 : INV_X1 port map( I => n27359, ZN => n762);
   U4696 : INV_X1 port map( I => n17803, ZN => n17802);
   U1263 : NAND2_X1 port map( A1 => n25002, A2 => n28104, ZN => n24766);
   U832 : OAI21_X1 port map( A1 => n11579, A2 => n22896, B => n22895, ZN => 
                           n13656);
   U5663 : INV_X1 port map( I => n17640, ZN => n15550);
   U7681 : NAND2_X1 port map( A1 => n17956, A2 => n10823, ZN => n6964);
   U4659 : NAND2_X1 port map( A1 => n1217, A2 => n17942, ZN => n8994);
   U622 : AOI21_X1 port map( A1 => n23197, A2 => n23564, B => n1203, ZN => 
                           n2900);
   U8981 : OAI21_X1 port map( A1 => n24958, A2 => n25200, B => n11419, ZN => 
                           n4006);
   U20868 : NOR2_X1 port map( A1 => n27820, A2 => n24175, ZN => n17955);
   U21601 : NOR2_X1 port map( A1 => n1203, A2 => n24292, ZN => n4103);
   U1305 : BUF_X2 port map( I => n17924, Z => n23915);
   U2599 : INV_X2 port map( I => n3929, ZN => n17729);
   U17903 : INV_X1 port map( I => n14255, ZN => n17797);
   U6431 : NAND2_X1 port map( A1 => n4461, A2 => n25192, ZN => n8218);
   U18610 : NAND2_X1 port map( A1 => n28022, A2 => n9675, ZN => n23810);
   U13961 : NAND2_X1 port map( A1 => n4976, A2 => n27640, ZN => n17997);
   U4713 : AOI21_X1 port map( A1 => n7825, A2 => n7247, B => n17830, ZN => 
                           n17831);
   U21906 : NAND2_X1 port map( A1 => n17791, A2 => n10030, ZN => n9733);
   U5648 : AOI22_X1 port map( A1 => n25929, A2 => n26533, B1 => n23915, B2 => 
                           n17928, ZN => n25924);
   U17911 : NAND2_X1 port map( A1 => n17656, A2 => n17729, ZN => n14994);
   U9775 : NAND2_X1 port map( A1 => n21778, A2 => n21779, ZN => n1863);
   U1204 : NAND3_X1 port map( A1 => n28105, A2 => n28104, A3 => n14826, ZN => 
                           n25078);
   U1184 : NAND3_X1 port map( A1 => n25493, A2 => n23115, A3 => n28247, ZN => 
                           n3207);
   U8564 : NOR2_X1 port map( A1 => n10823, A2 => n17959, ZN => n14816);
   U4611 : NOR2_X1 port map( A1 => n24586, A2 => n21792, ZN => n17939);
   U7718 : NAND2_X1 port map( A1 => n17651, A2 => n6629, ZN => n9165);
   U9745 : OAI21_X1 port map( A1 => n17985, A2 => n17984, B => n443, ZN => 
                           n17988);
   U1195 : INV_X1 port map( I => n17649, ZN => n5926);
   U3135 : OAI21_X1 port map( A1 => n17955, A2 => n12621, B => n17954, ZN => 
                           n7530);
   U9783 : NAND2_X1 port map( A1 => n15408, A2 => n24003, ZN => n6719);
   U4607 : NOR2_X1 port map( A1 => n17679, A2 => n17680, ZN => n2099);
   U15117 : NAND2_X1 port map( A1 => n12676, A2 => n5584, ZN => n10982);
   U7679 : AOI21_X1 port map( A1 => n15531, A2 => n15532, B => n4318, ZN => 
                           n7239);
   U1190 : OAI21_X1 port map( A1 => n4591, A2 => n2206, B => n4486, ZN => n2538
                           );
   U7703 : OAI21_X1 port map( A1 => n14230, A2 => n3929, B => n24808, ZN => 
                           n11824);
   U4983 : AOI21_X1 port map( A1 => n13730, A2 => n17972, B => n13217, ZN => 
                           n2328);
   U7638 : NOR2_X1 port map( A1 => n8184, A2 => n8183, ZN => n8182);
   U1198 : NAND2_X1 port map( A1 => n25719, A2 => n25720, ZN => n25212);
   U1317 : NAND3_X1 port map( A1 => n8917, A2 => n9675, A3 => n10816, ZN => 
                           n7322);
   U3300 : AOI21_X1 port map( A1 => n21859, A2 => n4306, B => n25192, ZN => 
                           n13275);
   U4987 : OAI21_X1 port map( A1 => n28540, A2 => n12516, B => n17928, ZN => 
                           n4561);
   U4996 : NOR2_X1 port map( A1 => n10058, A2 => n17989, ZN => n10509);
   U5609 : INV_X1 port map( I => n6718, ZN => n15056);
   U16168 : INV_X1 port map( I => n6867, ZN => n18105);
   U5260 : NAND2_X1 port map( A1 => n6642, A2 => n24391, ZN => n10508);
   U5641 : NAND2_X1 port map( A1 => n15056, A2 => n5300, ZN => n10163);
   U14050 : INV_X1 port map( I => n12276, ZN => n25631);
   U7695 : INV_X1 port map( I => n18125, ZN => n1777);
   U4880 : NAND2_X1 port map( A1 => n7413, A2 => n26473, ZN => n7801);
   U6414 : NAND3_X1 port map( A1 => n9854, A2 => n7002, A3 => n21436, ZN => 
                           n4238);
   U7667 : INV_X1 port map( I => n17731, ZN => n3613);
   U1402 : NOR2_X1 port map( A1 => n4072, A2 => n4288, ZN => n4071);
   U9582 : INV_X1 port map( I => n12718, ZN => n23681);
   U1164 : CLKBUF_X2 port map( I => n14139, Z => n25901);
   U5242 : CLKBUF_X2 port map( I => n7103, Z => n4310);
   U7398 : CLKBUF_X2 port map( I => n18359, Z => n22135);
   U6239 : INV_X1 port map( I => n18021, ZN => n1019);
   U554 : INV_X1 port map( I => n18649, ZN => n18444);
   U2530 : CLKBUF_X2 port map( I => n21923, Z => n235);
   U2306 : INV_X2 port map( I => n4131, ZN => n22547);
   U3392 : CLKBUF_X2 port map( I => n18427, Z => n22832);
   U511 : INV_X2 port map( I => n18455, ZN => n4198);
   U4774 : INV_X2 port map( I => n13184, ZN => n18778);
   U499 : INV_X2 port map( I => n18715, ZN => n783);
   U13452 : INV_X1 port map( I => n18498, ZN => n18748);
   U542 : INV_X1 port map( I => n7383, ZN => n1013);
   U16560 : INV_X1 port map( I => n18601, ZN => n7770);
   U18804 : NOR2_X1 port map( A1 => n11262, A2 => n18667, ZN => n18668);
   U2548 : NAND2_X1 port map( A1 => n18778, A2 => n13532, ZN => n14141);
   U1097 : INV_X2 port map( I => n18581, ZN => n10263);
   U7617 : INV_X1 port map( I => n18487, ZN => n18709);
   U3384 : BUF_X2 port map( I => n18414, Z => n5746);
   U2914 : CLKBUF_X2 port map( I => n14369, Z => n24133);
   U2703 : INV_X2 port map( I => n8113, ZN => n18705);
   U1108 : INV_X2 port map( I => n13619, ZN => n1179);
   U3988 : INV_X2 port map( I => n18687, ZN => n11453);
   U4969 : BUF_X2 port map( I => n18341, Z => n18585);
   U7616 : INV_X1 port map( I => n28542, ZN => n1187);
   U2080 : INV_X2 port map( I => n5986, ZN => n15623);
   U8768 : INV_X1 port map( I => n10564, ZN => n12569);
   U2568 : NAND2_X1 port map( A1 => n15448, A2 => n13969, ZN => n12732);
   U11037 : INV_X1 port map( I => n1618, ZN => n6800);
   U2018 : INV_X1 port map( I => n14287, ZN => n1003);
   U21734 : INV_X1 port map( I => n25609, ZN => n877);
   U519 : INV_X1 port map( I => n18642, ZN => n14362);
   U18145 : INV_X1 port map( I => n23415, ZN => n6041);
   U757 : OAI21_X1 port map( A1 => n18785, A2 => n2072, B => n18444, ZN => 
                           n12325);
   U20915 : NAND2_X1 port map( A1 => n26277, A2 => n4661, ZN => n22031);
   U2137 : INV_X2 port map( I => n18527, ZN => n18590);
   U3805 : INV_X2 port map( I => n18646, ZN => n18763);
   U6303 : INV_X1 port map( I => n6800, ZN => n25708);
   U1369 : NAND2_X1 port map( A1 => n18590, A2 => n1011, ZN => n10011);
   U5694 : NAND2_X1 port map( A1 => n18628, A2 => n18588, ZN => n12843);
   U713 : NOR2_X1 port map( A1 => n357, A2 => n7446, ZN => n7499);
   U9611 : INV_X1 port map( I => n14424, ZN => n10116);
   U9618 : NAND2_X1 port map( A1 => n4639, A2 => n18585, ZN => n18587);
   U15100 : OAI21_X1 port map( A1 => n758, A2 => n5554, B => n6593, ZN => 
                           n18064);
   U1077 : OAI21_X1 port map( A1 => n18706, A2 => n8113, B => n27895, ZN => 
                           n3744);
   U12762 : INV_X1 port map( I => n18424, ZN => n18489);
   U4017 : BUF_X2 port map( I => n18344, Z => n482);
   U17937 : AOI21_X1 port map( A1 => n18747, A2 => n25375, B => n18749, ZN => 
                           n12931);
   U6344 : NOR2_X1 port map( A1 => n11783, A2 => n4158, ZN => n4701);
   U14557 : OAI22_X1 port map( A1 => n1012, A2 => n11425, B1 => n5704, B2 => 
                           n14683, ZN => n23055);
   U4811 : NAND2_X1 port map( A1 => n14883, A2 => n18755, ZN => n4300);
   U9604 : NOR2_X1 port map( A1 => n8025, A2 => n1018, ZN => n18669);
   U6321 : NAND2_X1 port map( A1 => n18546, A2 => n820, ZN => n2783);
   U17942 : OAI21_X1 port map( A1 => n18705, A2 => n28306, B => n18706, ZN => 
                           n15405);
   U4732 : INV_X1 port map( I => n18700, ZN => n18703);
   U19120 : NOR2_X1 port map( A1 => n24523, A2 => n25382, ZN => n12200);
   U9438 : NOR2_X1 port map( A1 => n18439, A2 => n18769, ZN => n5246);
   U528 : INV_X2 port map( I => n24286, ZN => n2253);
   U5678 : NAND2_X1 port map( A1 => n3106, A2 => n13184, ZN => n25993);
   U9633 : BUF_X2 port map( I => n18683, Z => n11911);
   U9460 : INV_X1 port map( I => n14821, ZN => n7867);
   U4807 : NOR2_X1 port map( A1 => n2478, A2 => n25680, ZN => n12403);
   U12503 : NAND2_X1 port map( A1 => n1387, A2 => n13963, ZN => n14154);
   U9547 : NAND2_X1 port map( A1 => n18447, A2 => n18512, ZN => n13508);
   U9512 : NOR2_X1 port map( A1 => n18425, A2 => n26121, ZN => n9603);
   U7585 : INV_X1 port map( I => n18746, ZN => n12997);
   U19937 : INV_X2 port map( I => n14097, ZN => n18463);
   U1064 : NAND2_X1 port map( A1 => n22518, A2 => n820, ZN => n22955);
   U503 : NOR2_X1 port map( A1 => n18784, A2 => n18444, ZN => n18630);
   U9576 : NAND2_X1 port map( A1 => n11711, A2 => n9348, ZN => n2787);
   U20279 : NOR2_X1 port map( A1 => n11685, A2 => n1011, ZN => n18529);
   U513 : INV_X1 port map( I => n6041, ZN => n18751);
   U3251 : INV_X1 port map( I => n12672, ZN => n1722);
   U15435 : NOR2_X1 port map( A1 => n28481, A2 => n7841, ZN => n23876);
   U1566 : NOR2_X1 port map( A1 => n18785, A2 => n24243, ZN => n3387);
   U18098 : NOR2_X1 port map( A1 => n2072, A2 => n18444, ZN => n18786);
   U9586 : INV_X1 port map( I => n6438, ZN => n6512);
   U4594 : NOR2_X1 port map( A1 => n12699, A2 => n18475, ZN => n11035);
   U16364 : NAND2_X1 port map( A1 => n12375, A2 => n18623, ZN => n23453);
   U5622 : NOR2_X1 port map( A1 => n23743, A2 => n8254, ZN => n7500);
   U1039 : INV_X1 port map( I => n27026, ZN => n25709);
   U11527 : OR2_X1 port map( A1 => n26561, A2 => n25585, Z => n18534);
   U533 : INV_X2 port map( I => n18605, ZN => n15416);
   U5632 : INV_X1 port map( I => n18588, ZN => n8877);
   U16656 : NAND2_X1 port map( A1 => n6042, A2 => n25828, ZN => n2385);
   U15946 : NAND2_X1 port map( A1 => n18590, A2 => n1440, ZN => n10012);
   U4451 : INV_X2 port map( I => n18782, ZN => n18779);
   U2391 : NAND2_X1 port map( A1 => n10556, A2 => n18780, ZN => n18783);
   U725 : AOI21_X1 port map( A1 => n10437, A2 => n235, B => n18546, ZN => 
                           n15068);
   U14963 : OAI21_X1 port map( A1 => n13532, A2 => n11817, B => n1179, ZN => 
                           n10789);
   U5614 : INV_X1 port map( I => n1184, ZN => n880);
   U20988 : NAND2_X1 port map( A1 => n18747, A2 => n18749, ZN => n18641);
   U11067 : NAND3_X1 port map( A1 => n5746, A2 => n9508, A3 => n25261, ZN => 
                           n323);
   U984 : AOI22_X1 port map( A1 => n23761, A2 => n3902, B1 => n18537, B2 => 
                           n1326, ZN => n26102);
   U10355 : OAI22_X1 port map( A1 => n26721, A2 => n25935, B1 => n8333, B2 => 
                           n758, ZN => n25118);
   U711 : NOR2_X1 port map( A1 => n18145, A2 => n18585, ZN => n22993);
   U6327 : AOI21_X1 port map( A1 => n10872, A2 => n18763, B => n27830, ZN => 
                           n9474);
   U5606 : NOR2_X1 port map( A1 => n14022, A2 => n18763, ZN => n5116);
   U5704 : NOR2_X1 port map( A1 => n1722, A2 => n4959, ZN => n4961);
   U19506 : NAND3_X1 port map( A1 => n18684, A2 => n18682, A3 => n10596, ZN => 
                           n12886);
   U2323 : AOI21_X1 port map( A1 => n18586, A2 => n18507, B => n23540, ZN => 
                           n5439);
   U9487 : OAI21_X1 port map( A1 => n12375, A2 => n27888, B => n3310, ZN => 
                           n8436);
   U18979 : NAND2_X1 port map( A1 => n18703, A2 => n27497, ZN => n13984);
   U16456 : INV_X1 port map( I => n18463, ZN => n25803);
   U14036 : INV_X1 port map( I => n25500, ZN => n18509);
   U994 : NOR2_X1 port map( A1 => n15677, A2 => n11242, ZN => n22105);
   U1021 : OAI21_X1 port map( A1 => n2478, A2 => n18685, B => n8619, ZN => 
                           n4450);
   U17847 : NOR2_X1 port map( A1 => n5749, A2 => n11425, ZN => n25987);
   U3963 : NOR2_X1 port map( A1 => n18563, A2 => n11299, ZN => n22119);
   U16598 : NOR2_X1 port map( A1 => n5246, A2 => n5245, ZN => n10491);
   U7517 : OAI21_X1 port map( A1 => n3435, A2 => n3434, B => n1188, ZN => n4255
                           );
   U6334 : NOR3_X1 port map( A1 => n14569, A2 => n18489, A3 => n26282, ZN => 
                           n5037);
   U5588 : NAND2_X1 port map( A1 => n1010, A2 => n26657, ZN => n18539);
   U9597 : NOR2_X1 port map( A1 => n15693, A2 => n9248, ZN => n18468);
   U16270 : OAI21_X1 port map( A1 => n12711, A2 => n14207, B => n13969, ZN => 
                           n18488);
   U2198 : INV_X1 port map( I => n21790, ZN => n1000);
   U2225 : NOR2_X1 port map( A1 => n15144, A2 => n10708, ZN => n15143);
   U4814 : INV_X1 port map( I => n26209, ZN => n10039);
   U9175 : OAI21_X1 port map( A1 => n26744, A2 => n10152, B => n10930, ZN => 
                           n10929);
   U18127 : AOI21_X1 port map( A1 => n28090, A2 => n18748, B => n24701, ZN => 
                           n11636);
   U11662 : NOR2_X1 port map( A1 => n2253, A2 => n18458, ZN => n7677);
   U13113 : NAND2_X1 port map( A1 => n18488, A2 => n1004, ZN => n9712);
   U4002 : INV_X2 port map( I => n4549, ZN => n23392);
   U2821 : OR2_X1 port map( A1 => n14649, A2 => n18779, Z => n5879);
   U9477 : NAND2_X1 port map( A1 => n10908, A2 => n8123, ZN => n10919);
   U9523 : NOR2_X1 port map( A1 => n18468, A2 => n11382, ZN => n15673);
   U4749 : NAND2_X1 port map( A1 => n18511, A2 => n10537, ZN => n23791);
   U11737 : NAND2_X1 port map( A1 => n23332, A2 => n1006, ZN => n25262);
   U12359 : NAND2_X1 port map( A1 => n2949, A2 => n2948, ZN => n2947);
   U20055 : OAI21_X1 port map( A1 => n12385, A2 => n5645, B => n11911, ZN => 
                           n23428);
   U677 : NOR2_X1 port map( A1 => n23966, A2 => n1000, ZN => n22272);
   U4272 : OR2_X1 port map( A1 => n18693, A2 => n26700, Z => n10668);
   U7534 : OAI21_X1 port map( A1 => n880, A2 => n2982, B => n4091, ZN => n4090)
                           ;
   U19291 : NAND2_X1 port map( A1 => n23392, A2 => n7468, ZN => n15223);
   U2837 : INV_X1 port map( I => n6778, ZN => n993);
   U9540 : NAND2_X1 port map( A1 => n7677, A2 => n18472, ZN => n7676);
   U6293 : INV_X1 port map( I => n19189, ZN => n1154);
   U3907 : INV_X1 port map( I => n25514, ZN => n816);
   U12590 : NAND2_X1 port map( A1 => n5112, A2 => n5113, ZN => n25319);
   U5531 : INV_X2 port map( I => n22391, ZN => n736);
   U3061 : INV_X2 port map( I => n19091, ZN => n1164);
   U941 : AND2_X1 port map( A1 => n25563, A2 => n12996, Z => n25327);
   U4264 : INV_X2 port map( I => n1159, ZN => n990);
   U607 : INV_X1 port map( I => n18999, ZN => n1156);
   U2745 : NAND2_X1 port map( A1 => n19159, A2 => n22345, ZN => n8514);
   U10774 : INV_X2 port map( I => n8049, ZN => n18949);
   U11398 : NAND2_X1 port map( A1 => n9117, A2 => n6598, ZN => n5120);
   U12979 : NOR2_X1 port map( A1 => n23844, A2 => n19155, ZN => n6488);
   U3922 : BUF_X2 port map( I => n1716, Z => n24294);
   U4926 : NOR2_X1 port map( A1 => n987, A2 => n12521, ZN => n2993);
   U7519 : INV_X1 port map( I => n18939, ZN => n1166);
   U7426 : INV_X1 port map( I => n13028, ZN => n8471);
   U4940 : INV_X1 port map( I => n18953, ZN => n780);
   U3992 : CLKBUF_X2 port map( I => n14237, Z => n5393);
   U4698 : CLKBUF_X2 port map( I => n14338, Z => n444);
   U4588 : INV_X1 port map( I => n18794, ZN => n19055);
   U12133 : INV_X2 port map( I => n15429, ZN => n15040);
   U1117 : INV_X2 port map( I => n4702, ZN => n4703);
   U11147 : NOR2_X1 port map( A1 => n18920, A2 => n19091, ZN => n18996);
   U915 : INV_X1 port map( I => n1772, ZN => n12978);
   U6322 : OR2_X1 port map( A1 => n19191, A2 => n9216, Z => n24664);
   U901 : INV_X1 port map( I => n4034, ZN => n24061);
   U3282 : INV_X1 port map( I => n14382, ZN => n19152);
   U5741 : INV_X1 port map( I => n12584, ZN => n19122);
   U5195 : INV_X2 port map( I => n19143, ZN => n778);
   U5571 : NAND2_X1 port map( A1 => n1716, A2 => n23905, ZN => n18917);
   U20023 : NOR2_X1 port map( A1 => n24061, A2 => n23017, ZN => n5114);
   U5779 : NAND2_X1 port map( A1 => n26762, A2 => n19062, ZN => n19060);
   U21026 : OAI21_X1 port map( A1 => n23431, A2 => n19015, B => n14912, ZN => 
                           n19018);
   U8649 : INV_X1 port map( I => n3833, ZN => n24912);
   U14004 : NAND2_X1 port map( A1 => n873, A2 => n26570, ZN => n4545);
   U11520 : NAND2_X1 port map( A1 => n986, A2 => n26327, ZN => n10617);
   U795 : NOR2_X1 port map( A1 => n2177, A2 => n10801, ZN => n18872);
   U6248 : NOR2_X1 port map( A1 => n15041, A2 => n13812, ZN => n15518);
   U19839 : NOR2_X1 port map( A1 => n5393, A2 => n6487, ZN => n8695);
   U388 : INV_X1 port map( I => n19014, ZN => n12162);
   U12259 : NOR2_X1 port map( A1 => n24572, A2 => n1152, ZN => n9407);
   U19525 : OAI21_X1 port map( A1 => n18525, A2 => n180, B => n12981, ZN => 
                           n18877);
   U9395 : NOR2_X1 port map( A1 => n4705, A2 => n4702, ZN => n1396);
   U2936 : NAND2_X1 port map( A1 => n1494, A2 => n874, ZN => n1493);
   U4581 : INV_X1 port map( I => n9322, ZN => n13550);
   U2895 : NOR2_X1 port map( A1 => n9376, A2 => n9117, ZN => n24200);
   U6242 : NOR2_X1 port map( A1 => n818, A2 => n15041, ZN => n5944);
   U3899 : BUF_X2 port map( I => n3030, Z => n3009);
   U3905 : NOR2_X1 port map( A1 => n25514, A2 => n10894, ZN => n13229);
   U4685 : NOR2_X1 port map( A1 => n24265, A2 => n19079, ZN => n13488);
   U6268 : INV_X1 port map( I => n4212, ZN => n18945);
   U3548 : NOR2_X1 port map( A1 => n12978, A2 => n5990, ZN => n18898);
   U6438 : OR2_X1 port map( A1 => n22105, A2 => n19134, Z => n18968);
   U16278 : INV_X1 port map( I => n25592, ZN => n19103);
   U820 : INV_X1 port map( I => n19163, ZN => n18980);
   U9721 : INV_X2 port map( I => n27492, ZN => n19068);
   U412 : NOR2_X1 port map( A1 => n19145, A2 => n21767, ZN => n1897);
   U9342 : NOR2_X1 port map( A1 => n15224, A2 => n23392, ZN => n1814);
   U6220 : OAI21_X1 port map( A1 => n6602, A2 => n27868, B => n19036, ZN => 
                           n6601);
   U532 : NOR2_X1 port map( A1 => n1658, A2 => n7568, ZN => n19109);
   U17155 : NAND3_X1 port map( A1 => n23835, A2 => n1165, A3 => n28147, ZN => 
                           n18858);
   U17950 : NAND3_X1 port map( A1 => n14441, A2 => n14440, A3 => n23268, ZN => 
                           n14438);
   U21951 : NAND2_X1 port map( A1 => n23844, A2 => n19155, ZN => n23663);
   U779 : NAND2_X1 port map( A1 => n19073, A2 => n15435, ZN => n19075);
   U13011 : NAND2_X1 port map( A1 => n18990, A2 => n27813, ZN => n7994);
   U9323 : NAND2_X1 port map( A1 => n18974, A2 => n11331, ZN => n18253);
   U13681 : NAND3_X1 port map( A1 => n22949, A2 => n28548, A3 => n27787, ZN => 
                           n6768);
   U16699 : INV_X1 port map( I => n18945, ZN => n8082);
   U4835 : OAI21_X1 port map( A1 => n1396, A2 => n13812, B => n818, ZN => n3832
                           );
   U18351 : NAND2_X1 port map( A1 => n19131, A2 => n19132, ZN => n12627);
   U15326 : NAND3_X1 port map( A1 => n1150, A2 => n818, A3 => n5942, ZN => 
                           n5941);
   U4432 : NAND3_X1 port map( A1 => n23161, A2 => n14119, A3 => n18866, ZN => 
                           n2530);
   U551 : NOR2_X1 port map( A1 => n427, A2 => n782, ZN => n22551);
   U453 : OAI21_X1 port map( A1 => n18953, A2 => n19148, B => n22391, ZN => 
                           n22240);
   U12524 : NAND2_X1 port map( A1 => n987, A2 => n15040, ZN => n19077);
   U3194 : OAI21_X1 port map( A1 => n24201, A2 => n24200, B => n10083, ZN => 
                           n7213);
   U8080 : NAND2_X1 port map( A1 => n12542, A2 => n27704, ZN => n12698);
   U797 : NOR2_X1 port map( A1 => n23835, A2 => n19009, ZN => n9234);
   U5564 : INV_X1 port map( I => n19013, ZN => n13338);
   U5563 : INV_X1 port map( I => n18936, ZN => n8730);
   U396 : NAND2_X1 port map( A1 => n869, A2 => n11576, ZN => n12196);
   U13569 : NAND2_X1 port map( A1 => n14925, A2 => n26465, ZN => n19151);
   U14914 : AOI21_X1 port map( A1 => n15299, A2 => n778, B => n24466, ZN => 
                           n25584);
   U7404 : NAND2_X1 port map( A1 => n9032, A2 => n23161, ZN => n7503);
   U6957 : OAI21_X1 port map( A1 => n4736, A2 => n1159, B => n4734, ZN => n4731
                           );
   U1835 : NAND3_X1 port map( A1 => n14791, A2 => n13, A3 => n15434, ZN => 
                           n23665);
   U9214 : NOR2_X1 port map( A1 => n18399, A2 => n18796, ZN => n2908);
   U9844 : NAND3_X1 port map( A1 => n10735, A2 => n13587, A3 => n28444, ZN => 
                           n22605);
   U4104 : AOI21_X1 port map( A1 => n1818, A2 => n1817, B => n1816, ZN => n1815
                           );
   U12986 : AOI21_X1 port map( A1 => n4545, A2 => n4544, B => n22260, ZN => 
                           n4543);
   U3167 : NAND2_X1 port map( A1 => n95, A2 => n27647, ZN => n19120);
   U1964 : NAND3_X1 port map( A1 => n9881, A2 => n24055, A3 => n22634, ZN => 
                           n9880);
   U2609 : NOR2_X1 port map( A1 => n5138, A2 => n27043, ZN => n1976);
   U516 : NAND2_X1 port map( A1 => n1558, A2 => n24294, ZN => n18851);
   U11283 : AND2_X1 port map( A1 => n18847, A2 => n18827, Z => n3905);
   U2883 : INV_X1 port map( I => n9971, ZN => n8829);
   U3902 : AND2_X1 port map( A1 => n10894, A2 => n25514, Z => n3076);
   U18362 : NOR2_X1 port map( A1 => n18920, A2 => n9354, ZN => n15181);
   U3900 : OAI21_X1 port map( A1 => n26997, A2 => n21767, B => n2798, ZN => 
                           n3077);
   U13310 : AOI21_X1 port map( A1 => n11558, A2 => n23905, B => n11576, ZN => 
                           n18839);
   U2011 : INV_X1 port map( I => n19489, ZN => n2675);
   U11231 : OAI21_X1 port map( A1 => n1811, A2 => n1814, B => n1809, ZN => 
                           n19265);
   U13459 : NAND2_X1 port map( A1 => n23405, A2 => n14041, ZN => n22154);
   U12858 : INV_X1 port map( I => n1436, ZN => n25427);
   U6238 : NAND3_X1 port map( A1 => n25984, A2 => n21767, A3 => n27043, ZN => 
                           n1898);
   U12798 : INV_X1 port map( I => n19536, ZN => n1138);
   U20710 : AOI22_X1 port map( A1 => n18934, A2 => n23431, B1 => n13338, B2 => 
                           n18810, ZN => n18811);
   U374 : OAI21_X1 port map( A1 => n13869, A2 => n15181, B => n24306, ZN => 
                           n13868);
   U19457 : NAND2_X1 port map( A1 => n6930, A2 => n27647, ZN => n6927);
   U9358 : INV_X1 port map( I => n28548, ZN => n5984);
   U389 : NOR2_X1 port map( A1 => n1976, A2 => n1897, ZN => n1896);
   U12997 : AOI21_X1 port map( A1 => n22514, A2 => n18994, B => n23183, ZN => 
                           n13883);
   U20161 : NAND3_X1 port map( A1 => n6417, A2 => n6418, A3 => n18915, ZN => 
                           n6419);
   U6610 : NOR2_X1 port map( A1 => n3077, A2 => n3076, ZN => n14582);
   U4260 : NOR2_X1 port map( A1 => n6600, A2 => n24572, ZN => n11445);
   U4587 : BUF_X2 port map( I => n19453, Z => n26469);
   U15995 : INV_X2 port map( I => n21758, ZN => n7050);
   U793 : NAND2_X1 port map( A1 => n23161, A2 => n25070, ZN => n10843);
   U4860 : INV_X1 port map( I => n13357, ZN => n22081);
   U2204 : INV_X1 port map( I => n8374, ZN => n19166);
   U2308 : INV_X1 port map( I => n12527, ZN => n10828);
   U5181 : INV_X1 port map( I => n25270, ZN => n2581);
   U2012 : NAND2_X1 port map( A1 => n19236, A2 => n19489, ZN => n2676);
   U14680 : NAND2_X1 port map( A1 => n25544, A2 => n25543, ZN => n18854);
   U3352 : BUF_X2 port map( I => n19363, Z => n26012);
   U14576 : NAND2_X1 port map( A1 => n12546, A2 => n12545, ZN => n13982);
   U416 : INV_X1 port map( I => n19261, ZN => n984);
   U16294 : INV_X1 port map( I => n19302, ZN => n12202);
   U4737 : INV_X1 port map( I => n22845, ZN => n19728);
   U11278 : INV_X1 port map( I => n12952, ZN => n19645);
   U325 : INV_X2 port map( I => n11354, ZN => n754);
   U17272 : INV_X2 port map( I => n669, ZN => n19921);
   U3662 : INV_X2 port map( I => n1459, ZN => n19803);
   U1279 : NAND2_X1 port map( A1 => n9762, A2 => n10041, ZN => n11092);
   U1922 : BUF_X2 port map( I => n19755, Z => n2632);
   U12542 : INV_X2 port map( I => n4657, ZN => n14393);
   U3717 : INV_X2 port map( I => n9896, ZN => n19658);
   U9137 : INV_X1 port map( I => n19645, ZN => n2492);
   U3731 : INV_X2 port map( I => n14343, ZN => n19892);
   U623 : INV_X2 port map( I => n22140, ZN => n1120);
   U5541 : INV_X2 port map( I => n19808, ZN => n813);
   U4892 : NAND2_X1 port map( A1 => n8192, A2 => n2632, ZN => n8256);
   U6190 : INV_X1 port map( I => n27402, ZN => n1125);
   U14591 : INV_X2 port map( I => n25650, ZN => n19694);
   U4145 : INV_X1 port map( I => n7767, ZN => n19632);
   U645 : INV_X2 port map( I => n14726, ZN => n26271);
   U9807 : NAND2_X1 port map( A1 => n19915, A2 => n19914, ZN => n8887);
   U4736 : INV_X1 port map( I => n13121, ZN => n1130);
   U2549 : INV_X1 port map( I => n21916, ZN => n6394);
   U16681 : NOR2_X1 port map( A1 => n12666, A2 => n19935, ZN => n8033);
   U4054 : INV_X2 port map( I => n15478, ZN => n1491);
   U9277 : INV_X1 port map( I => n19923, ZN => n972);
   U11403 : NAND2_X1 port map( A1 => n10978, A2 => n19499, ZN => n19834);
   U4571 : INV_X1 port map( I => n27588, ZN => n755);
   U272 : INV_X1 port map( I => n24317, ZN => n19624);
   U6202 : INV_X1 port map( I => n26158, ZN => n11078);
   U14552 : INV_X1 port map( I => n10951, ZN => n8418);
   U654 : NAND2_X1 port map( A1 => n2320, A2 => n19623, ZN => n19635);
   U11946 : INV_X1 port map( I => n7326, ZN => n19676);
   U375 : INV_X1 port map( I => n4432, ZN => n22748);
   U1533 : INV_X1 port map( I => n19830, ZN => n15383);
   U2435 : INV_X1 port map( I => n10549, ZN => n211);
   U19997 : NOR2_X1 port map( A1 => n19758, A2 => n14279, ZN => n15489);
   U7819 : NAND2_X1 port map( A1 => n24196, A2 => n13387, ZN => n10862);
   U7258 : NAND2_X1 port map( A1 => n19749, A2 => n23868, ZN => n10042);
   U1759 : NOR2_X1 port map( A1 => n978, A2 => n10613, ZN => n3040);
   U8980 : AOI21_X1 port map( A1 => n19857, A2 => n4136, B => n24670, ZN => 
                           n10698);
   U2205 : AOI21_X1 port map( A1 => n23968, A2 => n19798, B => n2632, ZN => 
                           n5274);
   U2853 : NAND2_X1 port map( A1 => n19890, A2 => n19888, ZN => n23709);
   U10392 : OAI21_X1 port map( A1 => n976, A2 => n13110, B => n22688, ZN => 
                           n22687);
   U9084 : OAI21_X1 port map( A1 => n6393, A2 => n24579, B => n3226, ZN => 
                           n19779);
   U487 : NAND2_X1 port map( A1 => n14304, A2 => n211, ZN => n25014);
   U9026 : NAND2_X1 port map( A1 => n463, A2 => n14789, ZN => n14790);
   U18135 : NOR2_X1 port map( A1 => n19633, A2 => n19754, ZN => n19185);
   U636 : NOR2_X1 port map( A1 => n28268, A2 => n14393, ZN => n14410);
   U1786 : AOI21_X1 port map( A1 => n24861, A2 => n6191, B => n6811, ZN => 
                           n6190);
   U18156 : NAND3_X1 port map( A1 => n14304, A2 => n28378, A3 => n19823, ZN => 
                           n15748);
   U6753 : NAND2_X1 port map( A1 => n19750, A2 => n19930, ZN => n19573);
   U1826 : NOR2_X1 port map( A1 => n11778, A2 => n968, ZN => n14191);
   U4402 : INV_X1 port map( I => n19629, ZN => n9659);
   U10952 : OAI22_X1 port map( A1 => n8119, A2 => n10498, B1 => n863, B2 => 
                           n19936, ZN => n25167);
   U9411 : NAND2_X1 port map( A1 => n10498, A2 => n9561, ZN => n9368);
   U21343 : NOR2_X1 port map( A1 => n13926, A2 => n26415, ZN => n4181);
   U2091 : NAND2_X1 port map( A1 => n19946, A2 => n19947, ZN => n12389);
   U5947 : NOR2_X1 port map( A1 => n13110, A2 => n19650, ZN => n6143);
   U4909 : NOR2_X1 port map( A1 => n4810, A2 => n11369, ZN => n24102);
   U2290 : NOR2_X1 port map( A1 => n755, A2 => n15478, ZN => n7893);
   U600 : INV_X1 port map( I => n13854, ZN => n1117);
   U9035 : INV_X1 port map( I => n19671, ZN => n18862);
   U5960 : INV_X1 port map( I => n12617, ZN => n5839);
   U1438 : NAND2_X1 port map( A1 => n815, A2 => n19899, ZN => n19673);
   U4905 : INV_X2 port map( I => n26621, ZN => n4565);
   U307 : INV_X2 port map( I => n811, ZN => n7849);
   U15503 : INV_X2 port map( I => n11471, ZN => n15471);
   U14306 : NOR2_X1 port map( A1 => n12395, A2 => n1133, ZN => n25489);
   U6209 : INV_X1 port map( I => n11363, ZN => n8145);
   U19761 : INV_X1 port map( I => n19801, ZN => n24026);
   U1505 : AOI21_X1 port map( A1 => n19758, A2 => n19752, B => n3835, ZN => 
                           n6854);
   U2562 : AOI21_X1 port map( A1 => n7251, A2 => n11110, B => n9994, ZN => 
                           n6668);
   U3159 : INV_X1 port map( I => n21788, ZN => n21782);
   U16850 : OAI21_X1 port map( A1 => n15295, A2 => n13110, B => n1131, ZN => 
                           n25847);
   U2054 : OAI21_X1 port map( A1 => n964, A2 => n7251, B => n6668, ZN => n22257
                           );
   U10549 : OAI22_X1 port map( A1 => n967, A2 => n8004, B1 => n8464, B2 => 
                           n6865, ZN => n8463);
   U5149 : AOI21_X1 port map( A1 => n2891, A2 => n11988, B => n12395, ZN => 
                           n2823);
   U7176 : OAI21_X1 port map( A1 => n6561, A2 => n26522, B => n6560, ZN => 
                           n19963);
   U1559 : AOI21_X1 port map( A1 => n10520, A2 => n11988, B => n2925, ZN => 
                           n23501);
   U18188 : OAI21_X1 port map( A1 => n19768, A2 => n23977, B => n15471, ZN => 
                           n26041);
   U4894 : OAI21_X1 port map( A1 => n12441, A2 => n12440, B => n19945, ZN => 
                           n5099);
   U13519 : NAND2_X1 port map( A1 => n19838, A2 => n3861, ZN => n13797);
   U12248 : NOR2_X1 port map( A1 => n7849, A2 => n19893, ZN => n21961);
   U9085 : OAI21_X1 port map( A1 => n24109, A2 => n19903, B => n19706, ZN => 
                           n2121);
   U536 : NOR2_X1 port map( A1 => n7251, A2 => n11175, ZN => n13809);
   U19624 : OAI21_X1 port map( A1 => n26314, A2 => n19782, B => n1121, ZN => 
                           n3726);
   U7081 : NOR2_X1 port map( A1 => n174, A2 => n814, ZN => n11442);
   U5156 : OAI21_X1 port map( A1 => n11454, A2 => n2304, B => n3563, ZN => 
                           n10979);
   U17750 : OAI21_X1 port map( A1 => n18862, A2 => n2491, B => n23145, ZN => 
                           n23680);
   U6185 : NAND2_X1 port map( A1 => n19876, A2 => n3584, ZN => n10242);
   U13787 : OAI21_X1 port map( A1 => n4181, A2 => n211, B => n3317, ZN => n4180
                           );
   U9065 : NAND2_X1 port map( A1 => n6854, A2 => n6451, ZN => n1933);
   U2087 : NAND2_X1 port map( A1 => n15009, A2 => n24109, ZN => n13539);
   U3665 : NAND2_X1 port map( A1 => n10042, A2 => n9418, ZN => n23945);
   U3155 : NAND2_X1 port map( A1 => n27202, A2 => n756, ZN => n8561);
   U3412 : OAI21_X1 port map( A1 => n14411, A2 => n14410, B => n5421, ZN => 
                           n9825);
   U4945 : OR2_X1 port map( A1 => n8525, A2 => n19870, Z => n6057);
   U19646 : OAI21_X1 port map( A1 => n14429, A2 => n14430, B => n11471, ZN => 
                           n13311);
   U8954 : CLKBUF_X2 port map( I => n6821, Z => n3439);
   U7251 : NAND2_X1 port map( A1 => n19750, A2 => n14109, ZN => n19244);
   U5143 : NOR2_X1 port map( A1 => n8359, A2 => n22422, ZN => n15117);
   U21844 : NOR2_X1 port map( A1 => n6976, A2 => n12666, ZN => n24491);
   U4726 : NAND2_X1 port map( A1 => n972, A2 => n19921, ZN => n1687);
   U1948 : AOI22_X1 port map( A1 => n24413, A2 => n23169, B1 => n13345, B2 => 
                           n4241, ZN => n20096);
   U20723 : OAI21_X1 port map( A1 => n19612, A2 => n19952, B => n26021, ZN => 
                           n24144);
   U235 : NAND2_X1 port map( A1 => n11987, A2 => n20111, ZN => n11986);
   U8991 : NOR2_X1 port map( A1 => n2653, A2 => n11822, ZN => n12472);
   U7191 : NAND3_X1 port map( A1 => n19867, A2 => n27916, A3 => n23821, ZN => 
                           n6365);
   U5939 : NAND2_X1 port map( A1 => n6885, A2 => n24579, ZN => n13962);
   U2677 : INV_X1 port map( I => n24553, ZN => n20267);
   U216 : INV_X2 port map( I => n6821, ZN => n15461);
   U4555 : INV_X2 port map( I => n9579, ZN => n5577);
   U2969 : INV_X2 port map( I => n20023, ZN => n857);
   U5483 : INV_X2 port map( I => n25389, ZN => n10931);
   U2399 : INV_X1 port map( I => n3891, ZN => n15076);
   U2237 : INV_X1 port map( I => n12946, ZN => n2599);
   U4388 : INV_X1 port map( I => n20096, ZN => n20149);
   U3629 : CLKBUF_X2 port map( I => n20326, Z => n24383);
   U11961 : BUF_X2 port map( I => n7061, Z => n24421);
   U5022 : INV_X1 port map( I => n4191, ZN => n1113);
   U13060 : NAND2_X1 port map( A1 => n488, A2 => n19880, ZN => n25340);
   U15724 : INV_X2 port map( I => n23120, ZN => n20308);
   U12313 : INV_X1 port map( I => n2890, ZN => n20050);
   U12391 : INV_X1 port map( I => n14213, ZN => n11052);
   U10760 : INV_X1 port map( I => n7057, ZN => n19985);
   U6588 : NAND2_X1 port map( A1 => n2890, A2 => n20087, ZN => n20085);
   U5979 : NAND2_X1 port map( A1 => n956, A2 => n20272, ZN => n5905);
   U2353 : OAI21_X1 port map( A1 => n10721, A2 => n12479, B => n22342, ZN => 
                           n2513);
   U8886 : OAI21_X1 port map( A1 => n24027, A2 => n858, B => n23408, ZN => 
                           n1408);
   U13059 : NAND2_X1 port map( A1 => n12570, A2 => n19793, ZN => n22807);
   U7155 : OAI21_X1 port map( A1 => n21759, A2 => n26741, B => n20245, ZN => 
                           n3965);
   U3572 : NAND2_X1 port map( A1 => n23146, A2 => n3891, ZN => n8411);
   U12163 : NAND2_X1 port map( A1 => n25455, A2 => n2706, ZN => n8453);
   U3602 : INV_X1 port map( I => n7704, ZN => n24085);
   U2033 : INV_X1 port map( I => n6511, ZN => n5575);
   U238 : BUF_X2 port map( I => n8910, Z => n23725);
   U3362 : NOR2_X1 port map( A1 => n10436, A2 => n24534, ZN => n10433);
   U5464 : NAND2_X1 port map( A1 => n6264, A2 => n20235, ZN => n11151);
   U12198 : BUF_X2 port map( I => n12986, Z => n1108);
   U237 : NAND2_X1 port map( A1 => n20018, A2 => n22598, ZN => n20203);
   U3706 : CLKBUF_X1 port map( I => n20294, Z => n13252);
   U7075 : OAI21_X1 port map( A1 => n20259, A2 => n9921, B => n1103, ZN => 
                           n8895);
   U10455 : INV_X2 port map( I => n751, ZN => n23450);
   U1961 : INV_X2 port map( I => n857, ZN => n3870);
   U12744 : INV_X1 port map( I => n25959, ZN => n4660);
   U2231 : NOR2_X1 port map( A1 => n20018, A2 => n22374, ZN => n13315);
   U437 : INV_X1 port map( I => n20168, ZN => n807);
   U6065 : INV_X1 port map( I => n1104, ZN => n3460);
   U3160 : BUF_X2 port map( I => n11756, Z => n9446);
   U4418 : OR2_X1 port map( A1 => n10963, A2 => n8898, Z => n10662);
   U12615 : AND2_X1 port map( A1 => n4859, A2 => n12267, Z => n22758);
   U3521 : INV_X1 port map( I => n22374, ZN => n20290);
   U16145 : NOR2_X1 port map( A1 => n956, A2 => n27091, ZN => n25755);
   U12932 : INV_X1 port map( I => n14221, ZN => n10885);
   U12678 : NOR2_X1 port map( A1 => n12933, A2 => n23725, ZN => n21965);
   U8765 : NOR2_X1 port map( A1 => n22843, A2 => n1366, ZN => n7702);
   U5038 : NOR3_X1 port map( A1 => n20255, A2 => n22830, A3 => n26652, ZN => 
                           n3229);
   U2967 : NOR2_X1 port map( A1 => n20023, A2 => n4274, ZN => n3461);
   U3889 : NAND2_X1 port map( A1 => n751, A2 => n25959, ZN => n22625);
   U2006 : NOR3_X1 port map( A1 => n745, A2 => n20235, A3 => n6264, ZN => n6265
                           );
   U1394 : INV_X1 port map( I => n20136, ZN => n2767);
   U3102 : NOR2_X1 port map( A1 => n20290, A2 => n28277, ZN => n22373);
   U8874 : NOR2_X1 port map( A1 => n5576, A2 => n5575, ZN => n5574);
   U8876 : INV_X1 port map( I => n20099, ZN => n11072);
   U6043 : NAND2_X1 port map( A1 => n20127, A2 => n20166, ZN => n6606);
   U8815 : INV_X1 port map( I => n11398, ZN => n15597);
   U4421 : CLKBUF_X2 port map( I => n3803, Z => n25431);
   U12690 : NOR2_X1 port map( A1 => n13578, A2 => n27347, ZN => n11991);
   U7128 : NOR2_X1 port map( A1 => n21772, A2 => n334, ZN => n1757);
   U6022 : NAND2_X1 port map( A1 => n24720, A2 => n22835, ZN => n2971);
   U5859 : NOR2_X1 port map( A1 => n20213, A2 => n26009, ZN => n10225);
   U18423 : NOR2_X1 port map( A1 => n22295, A2 => n1110, ZN => n11957);
   U12165 : NAND2_X1 port map( A1 => n26410, A2 => n27668, ZN => n9877);
   U1811 : NOR3_X1 port map( A1 => n26189, A2 => n514, A3 => n27345, ZN => 
                           n24282);
   U3025 : INV_X1 port map( I => n12014, ZN => n8852);
   U8900 : INV_X1 port map( I => n14179, ZN => n20309);
   U15164 : NAND2_X1 port map( A1 => n4710, A2 => n24534, ZN => n23209);
   U7066 : INV_X1 port map( I => n8810, ZN => n20205);
   U371 : INV_X2 port map( I => n20317, ZN => n14104);
   U190 : NAND2_X1 port map( A1 => n4739, A2 => n2670, ZN => n14184);
   U170 : NOR2_X1 port map( A1 => n20188, A2 => n26252, ZN => n20041);
   U200 : NAND2_X1 port map( A1 => n4739, A2 => n27484, ZN => n24463);
   U2543 : AOI21_X1 port map( A1 => n15151, A2 => n20089, B => n1580, ZN => 
                           n20432);
   U6618 : NOR2_X1 port map( A1 => n24709, A2 => n22596, ZN => n15391);
   U21145 : NOR2_X1 port map( A1 => n27219, A2 => n22943, ZN => n19634);
   U5009 : NAND2_X1 port map( A1 => n958, A2 => n21863, ZN => n13259);
   U13572 : OAI21_X1 port map( A1 => n4781, A2 => n25999, B => n3933, ZN => 
                           n11544);
   U10366 : NAND2_X1 port map( A1 => n20130, A2 => n20129, ZN => n23481);
   U12604 : NOR2_X1 port map( A1 => n4269, A2 => n27129, ZN => n13396);
   U19963 : OAI21_X1 port map( A1 => n675, A2 => n5047, B => n14152, ZN => 
                           n19814);
   U14328 : NAND2_X1 port map( A1 => n733, A2 => n22807, ZN => n15280);
   U7119 : OAI21_X1 port map( A1 => n19965, A2 => n1110, B => n21932, ZN => 
                           n12247);
   U3949 : NOR2_X1 port map( A1 => n20269, A2 => n24394, ZN => n25960);
   U21602 : NAND3_X1 port map( A1 => n24293, A2 => n14497, A3 => n11920, ZN => 
                           n6422);
   U153 : OAI21_X1 port map( A1 => n26727, A2 => n11957, B => n25710, ZN => 
                           n11956);
   U6016 : NAND2_X1 port map( A1 => n19986, A2 => n955, ZN => n19991);
   U13474 : AOI21_X1 port map( A1 => n25431, A2 => n8265, B => n14179, ZN => 
                           n3802);
   U18237 : AOI21_X1 port map( A1 => n1101, A2 => n20317, B => n23676, ZN => 
                           n26089);
   U12639 : AOI21_X1 port map( A1 => n24083, A2 => n19969, B => n28408, ZN => 
                           n24495);
   U175 : NAND2_X1 port map( A1 => n14992, A2 => n14448, ZN => n14447);
   U1310 : NOR2_X1 port map( A1 => n22625, A2 => n12826, ZN => n23223);
   U183 : OAI22_X1 port map( A1 => n27487, A2 => n20171, B1 => n15413, B2 => 
                           n4783, ZN => n3990);
   U6173 : OR2_X1 port map( A1 => n2890, A2 => n13145, Z => n24605);
   U2811 : NAND2_X1 port map( A1 => n12701, A2 => n9919, ZN => n19579);
   U6686 : NAND3_X1 port map( A1 => n2655, A2 => n5213, A3 => n5609, ZN => 
                           n2518);
   U18397 : NAND2_X1 port map( A1 => n13271, A2 => n20011, ZN => n19578);
   U11044 : NAND2_X1 port map( A1 => n12632, A2 => n22569, ZN => n12629);
   U6517 : INV_X1 port map( I => n21374, ZN => n3419);
   U12734 : NAND2_X1 port map( A1 => n1573, A2 => n1572, ZN => n22771);
   U1714 : CLKBUF_X1 port map( I => n14601, Z => n36);
   U226 : CLKBUF_X2 port map( I => n9789, Z => n3390);
   U236 : INV_X1 port map( I => n23314, ZN => n21144);
   U3573 : NAND2_X1 port map( A1 => n7566, A2 => n11059, ZN => n22791);
   U1640 : INV_X1 port map( I => n20540, ZN => n8655);
   U167 : NOR3_X1 port map( A1 => n8479, A2 => n8478, A3 => n8477, ZN => n22820
                           );
   U215 : INV_X1 port map( I => n7813, ZN => n7812);
   U12311 : INV_X1 port map( I => n23173, ZN => n2888);
   U2591 : BUF_X2 port map( I => n13585, Z => n26329);
   U21635 : NAND2_X1 port map( A1 => n2519, A2 => n2518, ZN => n2520);
   U163 : NAND2_X1 port map( A1 => n3873, A2 => n3872, ZN => n3868);
   U1340 : INV_X1 port map( I => n3506, ZN => n1096);
   U15957 : INV_X1 port map( I => n21249, ZN => n20566);
   U1500 : INV_X2 port map( I => n21699, ZN => n945);
   U16576 : INV_X2 port map( I => n15501, ZN => n8050);
   U5444 : INV_X2 port map( I => n612, ZN => n20931);
   U12254 : INV_X2 port map( I => n25304, ZN => n21775);
   U11685 : BUF_X2 port map( I => n20405, Z => n20644);
   U11504 : INV_X1 port map( I => n8668, ZN => n25239);
   U128 : INV_X1 port map( I => n3462, ZN => n10578);
   U17297 : INV_X1 port map( I => n21270, ZN => n21064);
   U21318 : INV_X1 port map( I => n20631, ZN => n21721);
   U13021 : INV_X1 port map( I => n21723, ZN => n21696);
   U19779 : INV_X1 port map( I => n13642, ZN => n21716);
   U2770 : INV_X2 port map( I => n13979, ZN => n1077);
   U3737 : NAND2_X1 port map( A1 => n852, A2 => n21544, ZN => n11121);
   U127 : INV_X1 port map( I => n21924, ZN => n20920);
   U12429 : INV_X1 port map( I => n21027, ZN => n1082);
   U12448 : INV_X1 port map( I => n10519, ZN => n22747);
   U19667 : NAND2_X1 port map( A1 => n28027, A2 => n21699, ZN => n3923);
   U12159 : NAND2_X1 port map( A1 => n10591, A2 => n20345, ZN => n21572);
   U2602 : INV_X2 port map( I => n8050, ZN => n1083);
   U20120 : INV_X1 port map( I => n5675, ZN => n15616);
   U4374 : INV_X2 port map( I => n21624, ZN => n8735);
   U11888 : INV_X2 port map( I => n13900, ZN => n21395);
   U2212 : BUF_X2 port map( I => n21068, Z => n1090);
   U1554 : NAND2_X1 port map( A1 => n21444, A2 => n3549, ZN => n11743);
   U12196 : INV_X1 port map( I => n21715, ZN => n15315);
   U14123 : INV_X1 port map( I => n10591, ZN => n4623);
   U4278 : INV_X2 port map( I => n21586, ZN => n21618);
   U5446 : INV_X2 port map( I => n20736, ZN => n20781);
   U12486 : OR2_X1 port map( A1 => n10591, A2 => n14677, Z => n21630);
   U5105 : INV_X1 port map( I => n10732, ZN => n11490);
   U112 : INV_X1 port map( I => n26636, ZN => n20516);
   U4690 : INV_X1 port map( I => n9057, ZN => n10636);
   U12305 : INV_X1 port map( I => n2882, ZN => n7299);
   U4211 : INV_X1 port map( I => n21629, ZN => n21539);
   U10913 : OR2_X1 port map( A1 => n15670, A2 => n14348, Z => n21332);
   U177 : INV_X2 port map( I => n6547, ZN => n6522);
   U13472 : OR2_X1 port map( A1 => n27426, A2 => n6860, Z => n3560);
   U12818 : INV_X1 port map( I => n20732, ZN => n1081);
   U1778 : NOR2_X1 port map( A1 => n2569, A2 => n361, ZN => n21615);
   U12020 : AOI22_X1 port map( A1 => n6520, A2 => n6547, B1 => n10795, B2 => 
                           n21545, ZN => n25282);
   U12890 : NOR2_X1 port map( A1 => n21719, A2 => n21721, ZN => n20484);
   U10716 : OAI21_X1 port map( A1 => n24626, A2 => n28015, B => n20920, ZN => 
                           n25136);
   U103 : NOR3_X1 port map( A1 => n21720, A2 => n15307, A3 => n21719, ZN => 
                           n22388);
   U5958 : OAI21_X1 port map( A1 => n7807, A2 => n14113, B => n953, ZN => n8230
                           );
   U7046 : NAND3_X1 port map( A1 => n21507, A2 => n15646, A3 => n27363, ZN => 
                           n21459);
   U12117 : INV_X1 port map( I => n21462, ZN => n21259);
   U4262 : NAND2_X1 port map( A1 => n21205, A2 => n26554, ZN => n26553);
   U138 : AOI21_X1 port map( A1 => n15562, A2 => n15129, B => n11263, ZN => 
                           n23867);
   U12633 : INV_X2 port map( I => n3549, ZN => n849);
   U17593 : INV_X1 port map( I => n21572, ZN => n15570);
   U13242 : INV_X1 port map( I => n21666, ZN => n11759);
   U3460 : INV_X1 port map( I => n15208, ZN => n22046);
   U12906 : NAND2_X1 port map( A1 => n22737, A2 => n25841, ZN => n20556);
   U5971 : NAND2_X1 port map( A1 => n1078, A2 => n21100, ZN => n6676);
   U130 : NAND2_X1 port map( A1 => n731, A2 => n22737, ZN => n14460);
   U2258 : NAND2_X1 port map( A1 => n20938, A2 => n20932, ZN => n13440);
   U6100 : NAND2_X1 port map( A1 => n8198, A2 => n13287, ZN => n8469);
   U3336 : INV_X1 port map( I => n3593, ZN => n943);
   U3742 : OAI21_X1 port map( A1 => n7807, A2 => n10610, B => n732, ZN => n8247
                           );
   U8645 : NOR2_X1 port map( A1 => n13174, A2 => n8757, ZN => n9974);
   U5995 : INV_X2 port map( I => n27356, ZN => n15463);
   U1159 : INV_X1 port map( I => n21275, ZN => n13448);
   U3028 : AND2_X1 port map( A1 => n15353, A2 => n5722, Z => n5950);
   U13746 : INV_X1 port map( I => n4143, ZN => n13447);
   U5438 : NOR2_X1 port map( A1 => n13600, A2 => n21136, ZN => n21012);
   U12213 : OAI21_X1 port map( A1 => n20885, A2 => n20882, B => n10484, ZN => 
                           n6405);
   U5180 : AOI21_X1 port map( A1 => n12128, A2 => n20809, B => n20900, ZN => 
                           n24036);
   U3337 : NAND3_X1 port map( A1 => n25237, A2 => n3593, A3 => n3559, ZN => 
                           n22501);
   U21393 : NOR2_X1 port map( A1 => n9179, A2 => n20818, ZN => n20819);
   U12477 : NOR2_X1 port map( A1 => n13979, A2 => n21618, ZN => n15249);
   U18184 : NAND2_X1 port map( A1 => n21506, A2 => n14679, ZN => n21510);
   U6095 : NAND2_X1 port map( A1 => n8449, A2 => n5042, ZN => n11806);
   U83 : OAI21_X1 port map( A1 => n24548, A2 => n25721, B => n22364, ZN => 
                           n9694);
   U5934 : AOI21_X1 port map( A1 => n23802, A2 => n3549, B => n3195, ZN => 
                           n3661);
   U1932 : NAND3_X1 port map( A1 => n20856, A2 => n20758, A3 => n14806, ZN => 
                           n23334);
   U22016 : NAND2_X1 port map( A1 => n11562, A2 => n23225, ZN => n26580);
   U80 : NAND2_X1 port map( A1 => n25628, A2 => n20858, ZN => n25459);
   U7461 : NAND2_X1 port map( A1 => n11076, A2 => n2569, ZN => n3855);
   U91 : NAND2_X1 port map( A1 => n21328, A2 => n21324, ZN => n24976);
   U15907 : INV_X1 port map( I => n9567, ZN => n20710);
   U5138 : NAND2_X1 port map( A1 => n946, A2 => n13600, ZN => n65);
   U9148 : OAI21_X1 port map( A1 => n23514, A2 => n21328, B => n24976, ZN => 
                           n21331);
   U12692 : AOI22_X1 port map( A1 => n20968, A2 => n12067, B1 => n12066, B2 => 
                           n20969, ZN => n24444);
   U15499 : OAI21_X1 port map( A1 => n20401, A2 => n20639, B => n6243, ZN => 
                           n15312);
   U12783 : NAND2_X1 port map( A1 => n9074, A2 => n15713, ZN => n10534);
   U4862 : AOI21_X1 port map( A1 => n7088, A2 => n21614, B => n1076, ZN => 
                           n1769);
   U14245 : INV_X1 port map( I => n20654, ZN => n4767);
   U29 : NAND2_X1 port map( A1 => n23247, A2 => n8069, ZN => n22738);
   U41 : OR2_X1 port map( A1 => n12160, A2 => n1083, Z => n10658);
   U4183 : INV_X1 port map( I => n20875, ZN => n11868);
   U51 : OAI22_X1 port map( A1 => n11013, A2 => n216, B1 => n22209, B2 => 
                           n22208, ZN => n11837);
   U11949 : INV_X1 port map( I => n12011, ZN => n23578);
   U6949 : AOI21_X1 port map( A1 => n20747, A2 => n6408, B => n6407, ZN => 
                           n20748);
   U1620 : INV_X1 port map( I => n10851, ZN => n13799);
   U14955 : INV_X1 port map( I => n12797, ZN => n21565);
   U2736 : INV_X1 port map( I => n9894, ZN => n14350);
   U36 : INV_X1 port map( I => n13021, ZN => n21109);
   U17717 : INV_X1 port map( I => n20803, ZN => n10477);
   U32 : INV_X1 port map( I => n4413, ZN => n4604);
   U5901 : INV_X1 port map( I => n8271, ZN => n12517);
   U4178 : INV_X1 port map( I => n21606, ZN => n21612);
   U4220 : AND2_X1 port map( A1 => n8069, A2 => n23247, Z => n21880);
   U3966 : INV_X2 port map( I => n6052, ZN => n20749);
   U4853 : INV_X1 port map( I => n15470, ZN => n15475);
   U23 : INV_X1 port map( I => n21609, ZN => n15469);
   U1513 : INV_X1 port map( I => n8672, ZN => n6803);
   U27 : INV_X1 port map( I => n15287, ZN => n20624);
   U18101 : NOR2_X1 port map( A1 => n21734, A2 => n9894, ZN => n9893);
   U5872 : INV_X1 port map( I => n2749, ZN => n9460);
   U20 : INV_X1 port map( I => n13395, ZN => n1068);
   U1915 : NAND2_X1 port map( A1 => n24574, A2 => n11627, ZN => n25566);
   U2262 : INV_X1 port map( I => n934, ZN => n3759);
   U13539 : CLKBUF_X2 port map( I => n21052, Z => n9421);
   U3356 : CLKBUF_X2 port map( I => n21004, Z => n2307);
   U6943 : NAND3_X1 port map( A1 => n13842, A2 => n13841, A3 => n3725, ZN => 
                           n13961);
   U19566 : NOR2_X1 port map( A1 => n10385, A2 => n28308, ZN => n13126);
   U3746 : INV_X1 port map( I => n6517, ZN => n21483);
   U11 : INV_X1 port map( I => n6323, ZN => n10050);
   U14743 : INV_X1 port map( I => n12559, ZN => n10858);
   U9261 : INV_X1 port map( I => n21536, ZN => n770);
   U6 : OR2_X1 port map( A1 => n21663, A2 => n27395, Z => n25314);
   U12872 : OR2_X1 port map( A1 => n26377, A2 => n9565, Z => n25329);
   U12 : INV_X1 port map( I => n21487, ZN => n21473);
   U5095 : INV_X1 port map( I => n20704, ZN => n20695);
   U3 : INV_X1 port map( I => n2254, ZN => n20663);
   U8777 : OAI22_X1 port map( A1 => n7038, A2 => n26059, B1 => n21230, B2 => 
                           n26311, ZN => n11912);
   U2 : NAND3_X1 port map( A1 => n13921, A2 => n22892, A3 => n5486, ZN => 
                           n28114);
   U4 : NAND3_X1 port map( A1 => n9302, A2 => n9301, A3 => n12684, ZN => n27851
                           );
   U5 : AND2_X1 port map( A1 => n15458, A2 => n22844, Z => n26711);
   U8 : NAND2_X1 port map( A1 => n21741, A2 => n26647, ZN => n10975);
   U14 : NAND3_X1 port map( A1 => n11923, A2 => n13476, A3 => n21083, ZN => 
                           n26855);
   U16 : OAI21_X1 port map( A1 => n28347, A2 => n21738, B => n24685, ZN => 
                           n25562);
   U17 : NOR2_X1 port map( A1 => n21647, A2 => n21641, ZN => n21648);
   U18 : INV_X1 port map( I => n10268, ZN => n21222);
   U22 : AND2_X1 port map( A1 => n15470, A2 => n8271, Z => n21599);
   U24 : CLKBUF_X2 port map( I => n20680, Z => n7342);
   U31 : NAND2_X1 port map( A1 => n28055, A2 => n24951, ZN => n26952);
   U34 : INV_X1 port map( I => n21412, ZN => n27317);
   U37 : INV_X1 port map( I => n21711, ZN => n12018);
   U38 : INV_X1 port map( I => n20878, ZN => n1070);
   U42 : NAND2_X1 port map( A1 => n15199, A2 => n21659, ZN => n9319);
   U44 : NAND2_X1 port map( A1 => n21647, A2 => n21641, ZN => n21637);
   U48 : NAND2_X1 port map( A1 => n12046, A2 => n21000, ZN => n2514);
   U50 : AND2_X1 port map( A1 => n7296, A2 => n492, Z => n27439);
   U52 : INV_X1 port map( I => n1065, ZN => n27097);
   U53 : INV_X1 port map( I => n11492, ZN => n23579);
   U59 : INV_X1 port map( I => n3725, ZN => n27859);
   U62 : NAND2_X1 port map( A1 => n28274, A2 => n350, ZN => n27386);
   U69 : CLKBUF_X2 port map( I => n7516, Z => n6051);
   U75 : INV_X1 port map( I => n21086, ZN => n26649);
   U76 : BUF_X2 port map( I => n5578, Z => n5195);
   U78 : CLKBUF_X2 port map( I => n20654, Z => n4766);
   U84 : AND2_X1 port map( A1 => n21729, A2 => n2813, Z => n24278);
   U87 : AOI22_X1 port map( A1 => n552, A2 => n23991, B1 => n8751, B2 => n12476
                           , ZN => n28007);
   U88 : OAI22_X1 port map( A1 => n8278, A2 => n21059, B1 => n20560, B2 => 
                           n20971, ZN => n24765);
   U89 : OR2_X1 port map( A1 => n5071, A2 => n27380, Z => n7043);
   U92 : AOI22_X1 port map( A1 => n25509, A2 => n26651, B1 => n10547, B2 => 
                           n21543, ZN => n27076);
   U93 : NAND3_X1 port map( A1 => n8010, A2 => n8059, A3 => n1083, ZN => n22880
                           );
   U105 : NAND2_X1 port map( A1 => n21581, A2 => n21580, ZN => n22259);
   U110 : AOI21_X1 port map( A1 => n20923, A2 => n20922, B => n21099, ZN => 
                           n20924);
   U113 : NAND3_X1 port map( A1 => n23251, A2 => n24978, A3 => n26650, ZN => 
                           n27738);
   U115 : OAI21_X1 port map( A1 => n9005, A2 => n9004, B => n23054, ZN => 
                           n22937);
   U119 : NAND2_X1 port map( A1 => n21615, A2 => n1076, ZN => n1768);
   U120 : INV_X1 port map( I => n28017, ZN => n27260);
   U122 : NAND2_X1 port map( A1 => n1077, A2 => n23991, ZN => n28340);
   U124 : NOR2_X1 port map( A1 => n20900, A2 => n20899, ZN => n28040);
   U126 : AOI21_X1 port map( A1 => n1726, A2 => n22767, B => n14806, ZN => 
                           n2181);
   U133 : NOR2_X1 port map( A1 => n3096, A2 => n14679, ZN => n25696);
   U137 : AND2_X1 port map( A1 => n20732, A2 => n20728, Z => n20729);
   U140 : AND2_X1 port map( A1 => n25348, A2 => n12653, Z => n21591);
   U141 : NAND2_X1 port map( A1 => n22767, A2 => n20897, ZN => n20895);
   U147 : NOR2_X1 port map( A1 => n11905, A2 => n10031, ZN => n20558);
   U149 : AND2_X1 port map( A1 => n20932, A2 => n612, Z => n10586);
   U155 : NAND2_X1 port map( A1 => n20897, A2 => n20894, ZN => n1726);
   U157 : NOR2_X1 port map( A1 => n13791, A2 => n24538, ZN => n13790);
   U158 : INV_X1 port map( I => n11089, ZN => n26650);
   U161 : AND2_X1 port map( A1 => n14406, A2 => n13426, Z => n26686);
   U162 : INV_X1 port map( I => n9737, ZN => n21781);
   U164 : NAND2_X1 port map( A1 => n7956, A2 => n28197, ZN => n20926);
   U169 : NAND2_X1 port map( A1 => n12180, A2 => n20516, ZN => n8635);
   U173 : NAND2_X1 port map( A1 => n12654, A2 => n21506, ZN => n28020);
   U180 : INV_X1 port map( I => n950, ZN => n28059);
   U181 : NAND2_X1 port map( A1 => n25610, A2 => n20931, ZN => n28200);
   U182 : INV_X1 port map( I => n1515, ZN => n23125);
   U187 : NAND2_X1 port map( A1 => n14634, A2 => n3504, ZN => n21267);
   U188 : NOR2_X1 port map( A1 => n946, A2 => n13600, ZN => n26771);
   U192 : NOR2_X1 port map( A1 => n21775, A2 => n14718, ZN => n28508);
   U193 : NAND2_X1 port map( A1 => n15646, A2 => n14679, ZN => n8721);
   U195 : BUF_X2 port map( I => n21027, Z => n27689);
   U198 : INV_X1 port map( I => n20932, ZN => n25610);
   U199 : CLKBUF_X2 port map( I => n5841, Z => n27455);
   U203 : NAND2_X1 port map( A1 => n22767, A2 => n20894, ZN => n20860);
   U205 : NOR2_X1 port map( A1 => n26774, A2 => n26773, ZN => n26772);
   U207 : INV_X1 port map( I => n21092, ZN => n26773);
   U208 : CLKBUF_X2 port map( I => n21092, Z => n21136);
   U211 : BUF_X2 port map( I => n21101, Z => n13050);
   U212 : CLKBUF_X1 port map( I => n3466, Z => n27450);
   U217 : NAND2_X1 port map( A1 => n2199, A2 => n25830, ZN => n25361);
   U221 : INV_X1 port map( I => n15242, ZN => n11371);
   U225 : CLKBUF_X2 port map( I => n14653, Z => n7284);
   U232 : INV_X1 port map( I => n23849, ZN => n27302);
   U241 : AND2_X1 port map( A1 => n9760, A2 => n11462, Z => n26634);
   U243 : INV_X1 port map( I => n11880, ZN => n27650);
   U250 : INV_X1 port map( I => n12531, ZN => n23770);
   U253 : INV_X1 port map( I => n14243, ZN => n28159);
   U254 : INV_X2 port map( I => n27534, ZN => n5446);
   U257 : AND2_X1 port map( A1 => n24383, A2 => n12712, Z => n10770);
   U259 : OR2_X1 port map( A1 => n20122, A2 => n6006, Z => n21929);
   U260 : AOI21_X1 port map( A1 => n7618, A2 => n11519, B => n7457, ZN => n7635
                           );
   U261 : OAI21_X1 port map( A1 => n24464, A2 => n4739, B => n24463, ZN => 
                           n26909);
   U262 : NAND2_X1 port map( A1 => n27835, A2 => n26729, ZN => n10939);
   U267 : OAI21_X1 port map( A1 => n10582, A2 => n12631, B => n7457, ZN => 
                           n22569);
   U268 : NOR2_X1 port map( A1 => n14514, A2 => n24921, ZN => n27643);
   U269 : NAND2_X1 port map( A1 => n22183, A2 => n20330, ZN => n27158);
   U278 : NOR2_X1 port map( A1 => n8775, A2 => n27197, ZN => n8773);
   U280 : NAND3_X1 port map( A1 => n12362, A2 => n5049, A3 => n12801, ZN => 
                           n10487);
   U284 : AOI22_X1 port map( A1 => n11219, A2 => n26410, B1 => n27345, B2 => 
                           n15752, ZN => n6004);
   U285 : INV_X1 port map( I => n20141, ZN => n13732);
   U286 : NAND2_X1 port map( A1 => n26706, A2 => n14235, ZN => n28316);
   U287 : NOR2_X1 port map( A1 => n15752, A2 => n28098, ZN => n28097);
   U289 : NAND3_X1 port map( A1 => n9219, A2 => n28512, A3 => n4710, ZN => 
                           n23683);
   U292 : NAND3_X1 port map( A1 => n20260, A2 => n11463, A3 => n24720, ZN => 
                           n11462);
   U295 : NOR2_X1 port map( A1 => n959, A2 => n26969, ZN => n27778);
   U296 : NOR2_X1 port map( A1 => n20011, A2 => n20071, ZN => n10847);
   U299 : OAI22_X1 port map( A1 => n13429, A2 => n20318, B1 => n23674, B2 => 
                           n22815, ZN => n27953);
   U300 : NAND2_X1 port map( A1 => n3882, A2 => n7942, ZN => n22157);
   U301 : NAND2_X1 port map( A1 => n10356, A2 => n1105, ZN => n4791);
   U302 : NAND2_X1 port map( A1 => n6470, A2 => n20000, ZN => n26836);
   U306 : AOI22_X1 port map( A1 => n25056, A2 => n19981, B1 => n20254, B2 => 
                           n27846, ZN => n11123);
   U309 : NAND2_X1 port map( A1 => n135, A2 => n4710, ZN => n28511);
   U310 : NAND2_X1 port map( A1 => n1110, A2 => n4191, ZN => n27932);
   U312 : OAI21_X1 port map( A1 => n20232, A2 => n27347, B => n12933, ZN => 
                           n27509);
   U313 : INV_X1 port map( I => n20262, ZN => n27286);
   U315 : NOR2_X1 port map( A1 => n5248, A2 => n22921, ZN => n24380);
   U322 : INV_X1 port map( I => n4311, ZN => n15413);
   U323 : BUF_X2 port map( I => n20131, Z => n28408);
   U328 : NOR2_X1 port map( A1 => n26738, A2 => n9042, ZN => n20493);
   U337 : NAND3_X1 port map( A1 => n20238, A2 => n25598, A3 => n28519, ZN => 
                           n27006);
   U346 : NAND3_X1 port map( A1 => n26252, A2 => n28151, A3 => n20188, ZN => 
                           n27071);
   U350 : NAND3_X1 port map( A1 => n27434, A2 => n20237, A3 => n27674, ZN => 
                           n19169);
   U354 : NAND3_X1 port map( A1 => n27929, A2 => n27930, A3 => n20237, ZN => 
                           n26946);
   U355 : CLKBUF_X2 port map( I => n11487, Z => n25722);
   U356 : NAND2_X1 port map( A1 => n22066, A2 => n25076, ZN => n22291);
   U358 : AND2_X1 port map( A1 => n135, A2 => n13578, Z => n26703);
   U359 : AOI21_X1 port map( A1 => n13551, A2 => n26229, B => n20186, ZN => 
                           n24691);
   U360 : AOI21_X1 port map( A1 => n13682, A2 => n25141, B => n26890, ZN => 
                           n27525);
   U361 : AND2_X1 port map( A1 => n1110, A2 => n22776, Z => n26727);
   U362 : NOR2_X1 port map( A1 => n5664, A2 => n25455, ZN => n11219);
   U368 : INV_X2 port map( I => n26009, ZN => n25602);
   U372 : INV_X1 port map( I => n13864, ZN => n26995);
   U373 : INV_X1 port map( I => n6634, ZN => n1758);
   U376 : NAND3_X1 port map( A1 => n7345, A2 => n27951, A3 => n12177, ZN => 
                           n26947);
   U379 : NAND2_X1 port map( A1 => n858, A2 => n23416, ZN => n7931);
   U381 : NAND2_X1 port map( A1 => n20413, A2 => n27484, ZN => n20330);
   U384 : NAND3_X1 port map( A1 => n4709, A2 => n13578, A3 => n28512, ZN => 
                           n27519);
   U387 : OAI21_X1 port map( A1 => n1580, A2 => n20431, B => n14611, ZN => 
                           n24977);
   U390 : NAND2_X1 port map( A1 => n25418, A2 => n956, ZN => n9092);
   U393 : INV_X1 port map( I => n12644, ZN => n14991);
   U395 : NAND2_X1 port map( A1 => n5049, A2 => n675, ZN => n26825);
   U398 : INV_X1 port map( I => n12643, ZN => n14176);
   U399 : AND2_X1 port map( A1 => n7388, A2 => n12643, Z => n25760);
   U402 : NAND2_X1 port map( A1 => n5577, A2 => n5573, ZN => n5576);
   U403 : INV_X1 port map( I => n24283, ZN => n8452);
   U405 : BUF_X2 port map( I => n20490, Z => n334);
   U406 : CLKBUF_X2 port map( I => n14641, Z => n4709);
   U407 : INV_X1 port map( I => n7618, ZN => n27143);
   U408 : INV_X1 port map( I => n11583, ZN => n12492);
   U409 : NAND2_X1 port map( A1 => n7457, A2 => n5910, ZN => n9461);
   U414 : CLKBUF_X2 port map( I => n20174, Z => n9103);
   U420 : NOR2_X1 port map( A1 => n14059, A2 => n24862, ZN => n9298);
   U424 : NAND2_X1 port map( A1 => n2185, A2 => n4021, ZN => n25115);
   U429 : NAND2_X1 port map( A1 => n9365, A2 => n5080, ZN => n27815);
   U432 : AOI22_X1 port map( A1 => n26270, A2 => n27487, B1 => n25999, B2 => 
                           n4537, ZN => n26268);
   U436 : NOR2_X1 port map( A1 => n15076, A2 => n20139, ZN => n26863);
   U442 : NAND2_X1 port map( A1 => n20183, A2 => n20016, ZN => n27930);
   U445 : NAND2_X1 port map( A1 => n7969, A2 => n20023, ZN => n20022);
   U448 : INV_X1 port map( I => n20273, ZN => n27235);
   U451 : AND2_X1 port map( A1 => n15334, A2 => n1114, Z => n27398);
   U455 : NOR2_X1 port map( A1 => n20267, A2 => n20174, ZN => n20033);
   U459 : INV_X2 port map( I => n27873, ZN => n24534);
   U462 : INV_X1 port map( I => n20044, ZN => n28326);
   U465 : BUF_X2 port map( I => n6511, Z => n26652);
   U468 : CLKBUF_X2 port map( I => n20100, Z => n28525);
   U473 : INV_X2 port map( I => n20490, ZN => n1731);
   U478 : INV_X1 port map( I => n24533, ZN => n5906);
   U480 : NAND2_X1 port map( A1 => n12364, A2 => n11861, ZN => n27838);
   U482 : INV_X1 port map( I => n22374, ZN => n28399);
   U483 : INV_X1 port map( I => n2023, ZN => n13145);
   U486 : AOI21_X1 port map( A1 => n19633, A2 => n24431, B => n28484, ZN => 
                           n28119);
   U491 : NAND3_X1 port map( A1 => n8326, A2 => n27350, A3 => n10937, ZN => 
                           n12594);
   U492 : OAI21_X1 port map( A1 => n19840, A2 => n3861, B => n28441, ZN => 
                           n22707);
   U493 : NOR2_X1 port map( A1 => n24820, A2 => n27905, ZN => n27581);
   U497 : NOR2_X1 port map( A1 => n9732, A2 => n19099, ZN => n11692);
   U500 : NAND2_X1 port map( A1 => n9186, A2 => n27634, ZN => n25879);
   U501 : OAI21_X1 port map( A1 => n19903, A2 => n26948, B => n19906, ZN => 
                           n26933);
   U502 : OAI21_X1 port map( A1 => n28130, A2 => n28207, B => n26654, ZN => 
                           n12033);
   U506 : OAI21_X1 port map( A1 => n19951, A2 => n19952, B => n26021, ZN => 
                           n27786);
   U508 : NAND2_X1 port map( A1 => n19685, A2 => n19952, ZN => n27154);
   U515 : NAND2_X1 port map( A1 => n14240, A2 => n19928, ZN => n27708);
   U520 : NAND2_X1 port map( A1 => n27537, A2 => n8004, ZN => n22916);
   U521 : OAI21_X1 port map( A1 => n27881, A2 => n523, B => n11936, ZN => n9390
                           );
   U523 : NAND2_X1 port map( A1 => n19920, A2 => n1117, ZN => n161);
   U525 : NAND2_X1 port map( A1 => n19764, A2 => n15048, ZN => n28473);
   U527 : NAND3_X1 port map( A1 => n777, A2 => n775, A3 => n19694, ZN => n8146)
                           ;
   U537 : OAI21_X1 port map( A1 => n25230, A2 => n4565, B => n21782, ZN => 
                           n27336);
   U543 : NAND2_X1 port map( A1 => n19764, A2 => n19926, ZN => n12266);
   U548 : NOR2_X1 port map( A1 => n674, A2 => n14929, ZN => n2304);
   U550 : AOI21_X1 port map( A1 => n14651, A2 => n19951, B => n19952, ZN => 
                           n27153);
   U561 : NOR2_X1 port map( A1 => n26129, A2 => n24184, ZN => n12217);
   U562 : NOR2_X1 port map( A1 => n22775, A2 => n19937, ZN => n26994);
   U563 : AND2_X1 port map( A1 => n9701, A2 => n9583, Z => n5400);
   U564 : CLKBUF_X2 port map( I => n19798, Z => n28121);
   U567 : INV_X1 port map( I => n28377, ZN => n12467);
   U568 : NAND2_X1 port map( A1 => n26963, A2 => n14044, ZN => n19944);
   U570 : AND2_X1 port map( A1 => n19889, A2 => n19280, Z => n3916);
   U571 : AND2_X1 port map( A1 => n1121, A2 => n3954, Z => n26661);
   U572 : INV_X1 port map( I => n19892, ZN => n26990);
   U579 : NOR2_X1 port map( A1 => n28199, A2 => n19638, ZN => n27325);
   U583 : BUF_X2 port map( I => n19866, Z => n27916);
   U587 : CLKBUF_X2 port map( I => n14929, Z => n28264);
   U590 : NOR2_X1 port map( A1 => n5008, A2 => n12218, ZN => n10196);
   U596 : NAND2_X1 port map( A1 => n5738, A2 => n5739, ZN => n27037);
   U599 : CLKBUF_X2 port map( I => n19586, Z => n28130);
   U601 : NAND2_X1 port map( A1 => n4931, A2 => n6865, ZN => n26991);
   U602 : OAI21_X1 port map( A1 => n813, A2 => n9645, B => n9644, ZN => n6233);
   U603 : OAI21_X1 port map( A1 => n8417, A2 => n10956, B => n26296, ZN => 
                           n4394);
   U605 : NAND2_X1 port map( A1 => n24135, A2 => n14193, ZN => n26839);
   U608 : INV_X2 port map( I => n11110, ZN => n19945);
   U609 : NOR2_X1 port map( A1 => n1121, A2 => n3954, ZN => n19360);
   U612 : INV_X1 port map( I => n19586, ZN => n19678);
   U613 : INV_X1 port map( I => n4364, ZN => n15027);
   U617 : INV_X2 port map( I => n21769, ZN => n4931);
   U618 : BUF_X2 port map( I => n1127, Z => n28199);
   U625 : CLKBUF_X2 port map( I => n28224, Z => n27730);
   U626 : CLKBUF_X2 port map( I => n1459, Z => n27889);
   U628 : CLKBUF_X2 port map( I => n4364, Z => n27064);
   U635 : BUF_X2 port map( I => n606, Z => n34);
   U637 : NAND2_X1 port map( A1 => n14423, A2 => n26758, ZN => n26840);
   U643 : NAND2_X1 port map( A1 => n19658, A2 => n14393, ZN => n26986);
   U649 : NAND2_X1 port map( A1 => n2223, A2 => n15067, ZN => n5738);
   U651 : NAND2_X1 port map( A1 => n26447, A2 => n7612, ZN => n26828);
   U657 : BUF_X2 port map( I => n24336, Z => n27856);
   U658 : NOR2_X1 port map( A1 => n3954, A2 => n15310, ZN => n4324);
   U660 : INV_X1 port map( I => n24228, ZN => n24317);
   U662 : NOR2_X1 port map( A1 => n19400, A2 => n15573, ZN => n14568);
   U665 : CLKBUF_X2 port map( I => n8627, Z => n25081);
   U667 : CLKBUF_X4 port map( I => n19850, Z => n27823);
   U670 : INV_X2 port map( I => n19827, ZN => n19953);
   U676 : NAND3_X1 port map( A1 => n754, A2 => n19931, A3 => n19750, ZN => 
                           n25087);
   U680 : INV_X2 port map( I => n19400, ZN => n19809);
   U681 : INV_X1 port map( I => n28149, ZN => n14642);
   U684 : NAND2_X1 port map( A1 => n3150, A2 => n5467, ZN => n27422);
   U685 : CLKBUF_X2 port map( I => n12527, Z => n28460);
   U686 : INV_X1 port map( I => n5351, ZN => n28358);
   U688 : INV_X1 port map( I => n19496, ZN => n4626);
   U691 : INV_X1 port map( I => n982, ZN => n28096);
   U696 : BUF_X2 port map( I => n4126, Z => n27624);
   U697 : INV_X1 port map( I => n5698, ZN => n24794);
   U701 : INV_X1 port map( I => n9952, ZN => n5108);
   U705 : INV_X1 port map( I => n13918, ZN => n25794);
   U707 : NAND3_X1 port map( A1 => n994, A2 => n1163, A3 => n4471, ZN => n8063)
                           ;
   U708 : NAND2_X1 port map( A1 => n27626, A2 => n27894, ZN => n28179);
   U715 : NAND2_X1 port map( A1 => n27613, A2 => n19019, ZN => n18812);
   U741 : NOR3_X1 port map( A1 => n26446, A2 => n6040, A3 => n5393, ZN => 
                           n27646);
   U742 : OAI21_X1 port map( A1 => n2256, A2 => n28043, B => n23392, ZN => 
                           n23331);
   U747 : NAND2_X1 port map( A1 => n24630, A2 => n8485, ZN => n27906);
   U756 : NAND2_X1 port map( A1 => n8557, A2 => n25381, ZN => n22635);
   U759 : NAND3_X1 port map( A1 => n7260, A2 => n18807, A3 => n14257, ZN => 
                           n18451);
   U762 : NOR2_X1 port map( A1 => n28444, A2 => n28311, ZN => n7879);
   U764 : INV_X1 port map( I => n15704, ZN => n19053);
   U767 : NOR2_X1 port map( A1 => n13788, A2 => n5877, ZN => n14664);
   U771 : INV_X1 port map( I => n18808, ZN => n27613);
   U775 : OR2_X1 port map( A1 => n19081, A2 => n19082, Z => n15002);
   U778 : NAND2_X1 port map( A1 => n18964, A2 => n989, ZN => n27038);
   U781 : CLKBUF_X2 port map( I => n11376, Z => n7260);
   U784 : NAND2_X1 port map( A1 => n24265, A2 => n28237, ZN => n26903);
   U786 : OR2_X1 port map( A1 => n26764, A2 => n114, Z => n7072);
   U787 : NAND2_X1 port map( A1 => n18806, A2 => n18807, ZN => n27007);
   U788 : INV_X1 port map( I => n27432, ZN => n27277);
   U790 : NOR2_X1 port map( A1 => n11718, A2 => n19033, ZN => n28053);
   U794 : NAND3_X1 port map( A1 => n24442, A2 => n14271, A3 => n25664, ZN => 
                           n2399);
   U796 : NAND2_X1 port map( A1 => n18826, A2 => n19227, ZN => n27114);
   U801 : AOI21_X1 port map( A1 => n6013, A2 => n19167, B => n28444, ZN => 
                           n12566);
   U804 : NOR2_X1 port map( A1 => n26822, A2 => n18837, ZN => n26821);
   U808 : AOI21_X1 port map( A1 => n11839, A2 => n14580, B => n9354, ZN => 
                           n10480);
   U809 : AND2_X1 port map( A1 => n4735, A2 => n1159, Z => n26685);
   U810 : CLKBUF_X2 port map( I => n10362, Z => n25411);
   U814 : NAND2_X1 port map( A1 => n28499, A2 => n25327, ZN => n19131);
   U815 : NOR2_X1 port map( A1 => n95, A2 => n27799, ZN => n26756);
   U818 : BUF_X2 port map( I => n6089, Z => n23835);
   U825 : INV_X1 port map( I => n2701, ZN => n1443);
   U831 : NAND2_X1 port map( A1 => n19017, A2 => n18972, ZN => n24745);
   U834 : NOR2_X1 port map( A1 => n18999, A2 => n28547, ZN => n19086);
   U835 : OAI21_X1 port map( A1 => n4264, A2 => n19091, B => n27817, ZN => 
                           n9351);
   U838 : AOI21_X1 port map( A1 => n27775, A2 => n12542, B => n22809, ZN => 
                           n11913);
   U843 : OAI21_X1 port map( A1 => n1159, A2 => n13371, B => n13946, ZN => 
                           n10128);
   U847 : OAI22_X1 port map( A1 => n27942, A2 => n27941, B1 => n15704, B2 => 
                           n18797, ZN => n9311);
   U848 : INV_X1 port map( I => n28299, ZN => n26918);
   U856 : OR2_X1 port map( A1 => n19161, A2 => n8611, Z => n24340);
   U862 : INV_X1 port map( I => n18798, ZN => n8007);
   U864 : INV_X2 port map( I => n22727, ZN => n11718);
   U872 : CLKBUF_X2 port map( I => n8646, Z => n8645);
   U875 : BUF_X2 port map( I => n14098, Z => n22981);
   U884 : NOR2_X1 port map( A1 => n8988, A2 => n25176, ZN => n25102);
   U885 : INV_X1 port map( I => n18828, ZN => n28381);
   U894 : INV_X1 port map( I => n15224, ZN => n27948);
   U899 : NAND2_X1 port map( A1 => n14502, A2 => n24190, ZN => n18926);
   U904 : INV_X1 port map( I => n28384, ZN => n18932);
   U906 : INV_X2 port map( I => n988, ZN => n23017);
   U907 : BUF_X2 port map( I => n14654, Z => n22537);
   U909 : CLKBUF_X4 port map( I => n8683, Z => n24170);
   U916 : NAND2_X1 port map( A1 => n19057, A2 => n18396, ZN => n18526);
   U917 : NAND2_X1 port map( A1 => n27941, A2 => n24801, ZN => n28255);
   U919 : NOR2_X1 port map( A1 => n19155, A2 => n18939, ZN => n18940);
   U920 : NAND2_X1 port map( A1 => n18921, A2 => n8554, ZN => n18841);
   U922 : INV_X2 port map( I => n18799, ZN => n12542);
   U927 : INV_X2 port map( I => n10175, ZN => n28299);
   U936 : CLKBUF_X1 port map( I => n25099, Z => n27506);
   U947 : NAND2_X1 port map( A1 => n12967, A2 => n18693, ZN => n5070);
   U952 : INV_X1 port map( I => n4034, ZN => n27927);
   U959 : NAND2_X1 port map( A1 => n12991, A2 => n27207, ZN => n12470);
   U960 : NAND2_X1 port map( A1 => n15085, A2 => n15084, ZN => n27016);
   U962 : NAND2_X1 port map( A1 => n22035, A2 => n28515, ZN => n4787);
   U965 : NOR2_X1 port map( A1 => n27768, A2 => n22546, ZN => n11085);
   U966 : OR2_X1 port map( A1 => n10642, A2 => n18784, Z => n10759);
   U969 : NAND2_X1 port map( A1 => n18391, A2 => n11911, ZN => n27600);
   U971 : OAI21_X1 port map( A1 => n4552, A2 => n15131, B => n18602, ZN => 
                           n13244);
   U973 : AOI21_X1 port map( A1 => n881, A2 => n4158, B => n12671, ZN => n3122)
                           ;
   U976 : OAI21_X1 port map( A1 => n7078, A2 => n15623, B => n18476, ZN => 
                           n7678);
   U986 : AND2_X1 port map( A1 => n18585, A2 => n18583, Z => n26677);
   U988 : INV_X1 port map( I => n28437, ZN => n28436);
   U990 : AOI21_X1 port map( A1 => n6031, A2 => n14784, B => n6558, ZN => 
                           n28406);
   U991 : NOR2_X1 port map( A1 => n5341, A2 => n5342, ZN => n23544);
   U993 : NAND2_X1 port map( A1 => n18653, A2 => n7212, ZN => n25147);
   U995 : NAND2_X1 port map( A1 => n25993, A2 => n27050, ZN => n25891);
   U997 : NOR2_X1 port map( A1 => n23876, A2 => n13963, ZN => n28202);
   U999 : NAND3_X1 port map( A1 => n6031, A2 => n14128, A3 => n22973, ZN => 
                           n28379);
   U1000 : OAI22_X1 port map( A1 => n21852, A2 => n7190, B1 => n18584, B2 => 
                           n18583, ZN => n27096);
   U1001 : AOI21_X1 port map( A1 => n15019, A2 => n18580, B => n23062, ZN => 
                           n27768);
   U1004 : NOR3_X1 port map( A1 => n14498, A2 => n647, A3 => n5306, ZN => 
                           n18420);
   U1005 : NOR3_X1 port map( A1 => n13619, A2 => n13532, A3 => n10904, ZN => 
                           n27880);
   U1007 : INV_X1 port map( I => n18580, ZN => n18530);
   U1011 : NAND3_X1 port map( A1 => n2445, A2 => n10437, A3 => n18627, ZN => 
                           n28163);
   U1017 : CLKBUF_X2 port map( I => n22325, Z => n28184);
   U1023 : NOR2_X1 port map( A1 => n23624, A2 => n7791, ZN => n23623);
   U1027 : NOR2_X1 port map( A1 => n23761, A2 => n3902, ZN => n25275);
   U1035 : CLKBUF_X2 port map( I => n23004, Z => n25051);
   U1042 : NAND2_X1 port map( A1 => n4131, A2 => n18581, ZN => n15019);
   U1044 : OR2_X1 port map( A1 => n21790, A2 => n18645, Z => n10874);
   U1046 : OAI21_X1 port map( A1 => n3612, A2 => n1184, B => n2982, ZN => 
                           n18554);
   U1047 : NOR2_X1 port map( A1 => n18750, A2 => n6042, ZN => n6223);
   U1049 : NOR2_X1 port map( A1 => n12569, A2 => n6438, ZN => n3435);
   U1050 : NAND2_X1 port map( A1 => n13619, A2 => n13532, ZN => n27050);
   U1052 : NAND2_X1 port map( A1 => n18580, A2 => n25769, ZN => n22548);
   U1055 : INV_X1 port map( I => n15137, ZN => n14494);
   U1056 : INV_X1 port map( I => n18535, ZN => n1005);
   U1057 : OR2_X1 port map( A1 => n18782, A2 => n7965, Z => n13210);
   U1063 : CLKBUF_X2 port map( I => n14065, Z => n11919);
   U1065 : CLKBUF_X2 port map( I => n27797, Z => n27631);
   U1066 : CLKBUF_X1 port map( I => n23841, Z => n27715);
   U1067 : OAI21_X1 port map( A1 => n12672, A2 => n881, B => n4158, ZN => 
                           n28346);
   U1074 : NOR2_X1 port map( A1 => n14408, A2 => n18602, ZN => n28504);
   U1076 : INV_X2 port map( I => n15343, ZN => n27871);
   U1089 : INV_X1 port map( I => n28362, ZN => n28546);
   U1093 : BUF_X2 port map( I => n6945, Z => n9508);
   U1098 : BUF_X2 port map( I => n7087, Z => n2072);
   U1106 : CLKBUF_X2 port map( I => n18654, Z => n5306);
   U1113 : BUF_X2 port map( I => n11426, Z => n25261);
   U1119 : INV_X1 port map( I => n25985, ZN => n27710);
   U1123 : BUF_X2 port map( I => n18246, Z => n27137);
   U1127 : INV_X1 port map( I => n18058, ZN => n27732);
   U1128 : CLKBUF_X2 port map( I => n12439, Z => n28393);
   U1129 : INV_X1 port map( I => n7951, ZN => n27891);
   U1135 : NOR2_X1 port map( A1 => n27633, A2 => n18092, ZN => n11734);
   U1137 : NAND2_X1 port map( A1 => n14474, A2 => n25158, ZN => n27348);
   U1139 : CLKBUF_X2 port map( I => n24318, Z => n28466);
   U1142 : CLKBUF_X2 port map( I => n7413, Z => n25000);
   U1144 : NAND2_X1 port map( A1 => n28439, A2 => n13826, ZN => n27489);
   U1145 : OAI21_X1 port map( A1 => n27307, A2 => n14816, B => n10673, ZN => 
                           n17379);
   U1146 : INV_X1 port map( I => n18331, ZN => n1199);
   U1148 : BUF_X2 port map( I => n6675, Z => n27564);
   U1149 : NOR2_X1 port map( A1 => n739, A2 => n27766, ZN => n27765);
   U1151 : NAND2_X1 port map( A1 => n22584, A2 => n28003, ZN => n3711);
   U1153 : AOI22_X1 port map( A1 => n14052, A2 => n23696, B1 => n826, B2 => 
                           n14053, ZN => n25158);
   U1154 : NAND2_X1 port map( A1 => n17376, A2 => n23542, ZN => n27116);
   U1155 : OR2_X1 port map( A1 => n17722, A2 => n6629, Z => n17320);
   U1156 : INV_X1 port map( I => n6415, ZN => n17662);
   U1163 : OAI21_X1 port map( A1 => n17629, A2 => n13698, B => n27008, ZN => 
                           n5150);
   U1165 : NOR2_X1 port map( A1 => n27323, A2 => n1203, ZN => n6136);
   U1167 : NAND3_X1 port map( A1 => n17642, A2 => n22765, A3 => n17739, ZN => 
                           n17643);
   U1169 : NAND2_X1 port map( A1 => n24599, A2 => n22812, ZN => n10074);
   U1172 : AOI22_X1 port map( A1 => n11632, A2 => n828, B1 => n17873, B2 => 
                           n9040, ZN => n2249);
   U1173 : NAND2_X1 port map( A1 => n12815, A2 => n17687, ZN => n10871);
   U1178 : NAND2_X1 port map( A1 => n25903, A2 => n1022, ZN => n17681);
   U1187 : NOR2_X1 port map( A1 => n11514, A2 => n9105, ZN => n28037);
   U1192 : AND2_X1 port map( A1 => n11112, A2 => n17722, Z => n5361);
   U1197 : NOR3_X1 port map( A1 => n27458, A2 => n23923, A3 => n12815, ZN => 
                           n13217);
   U1199 : NAND2_X1 port map( A1 => n17918, A2 => n11419, ZN => n25719);
   U1201 : NAND2_X1 port map( A1 => n28005, A2 => n28004, ZN => n28003);
   U1206 : AOI21_X1 port map( A1 => n17933, A2 => n17637, B => n24195, ZN => 
                           n24194);
   U1207 : BUF_X2 port map( I => n1026, Z => n28457);
   U1208 : NOR2_X1 port map( A1 => n21779, A2 => n1882, ZN => n27496);
   U1211 : CLKBUF_X2 port map( I => n17976, Z => n13698);
   U1212 : OR2_X1 port map( A1 => n24570, A2 => n27749, Z => n5480);
   U1215 : AND2_X1 port map( A1 => n26144, A2 => n17728, Z => n26671);
   U1221 : NAND2_X1 port map( A1 => n23245, A2 => n3347, ZN => n27164);
   U1224 : NAND2_X1 port map( A1 => n28234, A2 => n23469, ZN => n2705);
   U1225 : NAND3_X1 port map( A1 => n27521, A2 => n2401, A3 => n22153, ZN => 
                           n25061);
   U1226 : NAND2_X1 port map( A1 => n26387, A2 => n21881, ZN => n14903);
   U1230 : NOR2_X1 port map( A1 => n5238, A2 => n26897, ZN => n27185);
   U1232 : AOI21_X1 port map( A1 => n28194, A2 => n6038, B => n716, ZN => 
                           n27825);
   U1233 : NOR2_X1 port map( A1 => n11182, A2 => n17761, ZN => n14196);
   U1235 : INV_X2 port map( I => n23231, ZN => n21778);
   U1237 : INV_X1 port map( I => n23923, ZN => n27756);
   U1244 : NAND2_X1 port map( A1 => n8626, A2 => n8625, ZN => n27359);
   U1245 : INV_X2 port map( I => n17974, ZN => n12815);
   U1246 : INV_X1 port map( I => n17969, ZN => n17723);
   U1255 : INV_X1 port map( I => n27211, ZN => n24599);
   U1258 : NOR2_X1 port map( A1 => n24570, A2 => n1211, ZN => n6916);
   U1261 : INV_X1 port map( I => n17957, ZN => n27483);
   U1262 : BUF_X2 port map( I => n12600, Z => n28288);
   U1268 : INV_X1 port map( I => n26356, ZN => n26897);
   U1273 : NAND2_X1 port map( A1 => n25787, A2 => n17657, ZN => n17634);
   U1274 : INV_X1 port map( I => n17470, ZN => n27556);
   U1277 : INV_X1 port map( I => n9630, ZN => n4470);
   U1280 : INV_X1 port map( I => n17614, ZN => n28456);
   U1283 : INV_X1 port map( I => n17767, ZN => n26544);
   U1285 : INV_X1 port map( I => n8000, ZN => n27577);
   U1289 : AOI21_X1 port map( A1 => n17636, A2 => n829, B => n23231, ZN => 
                           n27178);
   U1291 : BUF_X2 port map( I => n4610, Z => n28401);
   U1293 : NAND2_X1 port map( A1 => n23064, A2 => n4319, ZN => n23233);
   U1295 : INV_X1 port map( I => n10513, ZN => n17943);
   U1296 : NAND2_X1 port map( A1 => n17766, A2 => n25856, ZN => n17767);
   U1297 : INV_X1 port map( I => n12708, ZN => n17881);
   U1302 : INV_X1 port map( I => n17897, ZN => n17871);
   U1304 : NAND2_X1 port map( A1 => n17941, A2 => n10513, ZN => n10136);
   U1313 : NAND2_X1 port map( A1 => n8658, A2 => n4531, ZN => n17614);
   U1326 : BUF_X2 port map( I => n12610, Z => n12590);
   U1329 : BUF_X2 port map( I => n17617, Z => n4914);
   U1332 : BUF_X4 port map( I => n26218, Z => n24570);
   U1333 : CLKBUF_X2 port map( I => n28302, Z => n27029);
   U1334 : INV_X1 port map( I => n22817, ZN => n27055);
   U1335 : NAND2_X1 port map( A1 => n13281, A2 => n13280, ZN => n27230);
   U1337 : OAI21_X1 port map( A1 => n17314, A2 => n8237, B => n17312, ZN => 
                           n6195);
   U1344 : NOR2_X1 port map( A1 => n17174, A2 => n27561, ZN => n1513);
   U1346 : OAI21_X1 port map( A1 => n17518, A2 => n7996, B => n27959, ZN => 
                           n9142);
   U1348 : NAND3_X1 port map( A1 => n24018, A2 => n5639, A3 => n17514, ZN => 
                           n5887);
   U1352 : NOR3_X1 port map( A1 => n6425, A2 => n26691, A3 => n26782, ZN => 
                           n199);
   U1365 : OAI21_X1 port map( A1 => n26873, A2 => n26872, B => n10903, ZN => 
                           n26930);
   U1366 : OAI21_X1 port map( A1 => n5093, A2 => n17518, B => n5092, ZN => 
                           n28036);
   U1367 : NAND2_X1 port map( A1 => n4687, A2 => n17427, ZN => n27106);
   U1368 : OAI21_X1 port map( A1 => n2610, A2 => n17541, B => n26796, ZN => 
                           n2083);
   U1370 : NAND3_X1 port map( A1 => n17360, A2 => n17359, A3 => n9018, ZN => 
                           n27047);
   U1372 : AOI21_X1 port map( A1 => n5488, A2 => n9898, B => n17460, ZN => 
                           n16934);
   U1373 : AOI21_X1 port map( A1 => n27180, A2 => n5488, B => n8335, ZN => 
                           n3676);
   U1374 : AOI22_X1 port map( A1 => n17575, A2 => n17346, B1 => n17185, B2 => 
                           n17501, ZN => n2740);
   U1377 : INV_X1 port map( I => n6681, ZN => n17554);
   U1378 : NAND2_X1 port map( A1 => n17347, A2 => n17232, ZN => n5408);
   U1379 : NAND2_X1 port map( A1 => n24091, A2 => n2377, ZN => n17573);
   U1382 : NOR2_X1 port map( A1 => n14367, A2 => n28539, ZN => n28244);
   U1383 : OR2_X1 port map( A1 => n14990, A2 => n28490, Z => n13534);
   U1388 : OAI21_X1 port map( A1 => n15322, A2 => n23604, B => n17513, ZN => 
                           n5767);
   U1389 : CLKBUF_X2 port map( I => n17546, Z => n24368);
   U1391 : NAND2_X1 port map( A1 => n4250, A2 => n25057, ZN => n27886);
   U1392 : NOR2_X1 port map( A1 => n24706, A2 => n2499, ZN => n27925);
   U1398 : NOR2_X1 port map( A1 => n8538, A2 => n7498, ZN => n27478);
   U1399 : NAND2_X1 port map( A1 => n13218, A2 => n17328, ZN => n27804);
   U1401 : AOI21_X1 port map( A1 => n24214, A2 => n24419, B => n23449, ZN => 
                           n3620);
   U1404 : AOI21_X1 port map( A1 => n17560, A2 => n17559, B => n17561, ZN => 
                           n24349);
   U1405 : NOR2_X1 port map( A1 => n26628, A2 => n4832, ZN => n26923);
   U1409 : OAI22_X1 port map( A1 => n17326, A2 => n17518, B1 => n17450, B2 => 
                           n26213, ZN => n27963);
   U1417 : INV_X1 port map( I => n17463, ZN => n17409);
   U1419 : INV_X1 port map( I => n17414, ZN => n9132);
   U1420 : NOR2_X1 port map( A1 => n3091, A2 => n193, ZN => n13535);
   U1423 : INV_X1 port map( I => n14990, ZN => n717);
   U1426 : CLKBUF_X2 port map( I => n8165, Z => n28389);
   U1428 : CLKBUF_X2 port map( I => n13247, Z => n7357);
   U1430 : OR2_X1 port map( A1 => n8165, A2 => n5391, Z => n17435);
   U1434 : NAND2_X1 port map( A1 => n25013, A2 => n8237, ZN => n3430);
   U1439 : NAND2_X1 port map( A1 => n11270, A2 => n17510, ZN => n25568);
   U1440 : NOR2_X1 port map( A1 => n17447, A2 => n21785, ZN => n27299);
   U1443 : INV_X1 port map( I => n27088, ZN => n28539);
   U1447 : INV_X2 port map( I => n3980, ZN => n27946);
   U1453 : NOR2_X1 port map( A1 => n2377, A2 => n14639, ZN => n28218);
   U1455 : INV_X1 port map( I => n26616, ZN => n27958);
   U1459 : INV_X1 port map( I => n26616, ZN => n1435);
   U1460 : INV_X1 port map( I => n7399, ZN => n26793);
   U1462 : INV_X1 port map( I => n14492, ZN => n26656);
   U1466 : INV_X1 port map( I => n12192, ZN => n27591);
   U1468 : INV_X1 port map( I => n15609, ZN => n27108);
   U1473 : BUF_X2 port map( I => n6104, Z => n27084);
   U1476 : NAND2_X1 port map( A1 => n16420, A2 => n13211, ZN => n14761);
   U1477 : AOI22_X1 port map( A1 => n25195, A2 => n1046, B1 => n2313, B2 => 
                           n16688, ZN => n6348);
   U1482 : NAND2_X1 port map( A1 => n9829, A2 => n14254, ZN => n16533);
   U1491 : NAND2_X1 port map( A1 => n4518, A2 => n4940, ZN => n10981);
   U1493 : NOR2_X1 port map( A1 => n16692, A2 => n26734, ZN => n12464);
   U1496 : OAI21_X1 port map( A1 => n14562, A2 => n28172, B => n25397, ZN => 
                           n2353);
   U1501 : NOR2_X1 port map( A1 => n13786, A2 => n26396, ZN => n28107);
   U1503 : NAND3_X1 port map( A1 => n2422, A2 => n13137, A3 => n25772, ZN => 
                           n27165);
   U1504 : NOR2_X1 port map( A1 => n24484, A2 => n2976, ZN => n27017);
   U1507 : NAND2_X1 port map( A1 => n27781, A2 => n1984, ZN => n1983);
   U1520 : AND2_X1 port map( A1 => n5324, A2 => n25940, Z => n11443);
   U1521 : OR2_X1 port map( A1 => n6766, A2 => n11413, Z => n6618);
   U1522 : INV_X1 port map( I => n3751, ZN => n24347);
   U1528 : INV_X1 port map( I => n28356, ZN => n23531);
   U1545 : OR2_X1 port map( A1 => n16516, A2 => n12637, Z => n10714);
   U1550 : NAND2_X1 port map( A1 => n27975, A2 => n25482, ZN => n15888);
   U1552 : NAND2_X1 port map( A1 => n3087, A2 => n6688, ZN => n27133);
   U1557 : NAND2_X1 port map( A1 => n28400, A2 => n27543, ZN => n25501);
   U1563 : NAND2_X1 port map( A1 => n16410, A2 => n906, ZN => n7432);
   U1564 : INV_X2 port map( I => n8199, ZN => n28108);
   U1567 : NOR2_X1 port map( A1 => n16471, A2 => n4518, ZN => n6815);
   U1569 : NAND2_X1 port map( A1 => n16507, A2 => n2481, ZN => n27328);
   U1572 : INV_X1 port map( I => n16649, ZN => n28083);
   U1573 : NAND2_X1 port map( A1 => n404, A2 => n132, ZN => n27975);
   U1576 : NAND2_X1 port map( A1 => n7378, A2 => n16513, ZN => n16575);
   U1582 : INV_X1 port map( I => n4518, ZN => n4737);
   U1584 : CLKBUF_X4 port map( I => n12331, Z => n24770);
   U1586 : OAI21_X1 port map( A1 => n25685, A2 => n22838, B => n24839, ZN => 
                           n8533);
   U1594 : NOR2_X1 port map( A1 => n8199, A2 => n26396, ZN => n4339);
   U1596 : INV_X2 port map( I => n13138, ZN => n28400);
   U1598 : AND2_X1 port map( A1 => n5118, A2 => n4683, Z => n26690);
   U1600 : NAND2_X1 port map( A1 => n5081, A2 => n9773, ZN => n3123);
   U1606 : INV_X2 port map( I => n27472, ZN => n6763);
   U1607 : NAND3_X1 port map( A1 => n16355, A2 => n7226, A3 => n2044, ZN => 
                           n27263);
   U1609 : NAND2_X1 port map( A1 => n13265, A2 => n14880, ZN => n27978);
   U1612 : OR2_X1 port map( A1 => n26104, A2 => n121, Z => n10827);
   U1613 : NAND2_X1 port map( A1 => n7219, A2 => n915, ZN => n15950);
   U1615 : NOR2_X1 port map( A1 => n1419, A2 => n1270, ZN => n26895);
   U1617 : NAND2_X1 port map( A1 => n4954, A2 => n6842, ZN => n6841);
   U1626 : AOI22_X1 port map( A1 => n2703, A2 => n719, B1 => n516, B2 => n16329
                           , ZN => n2825);
   U1628 : AOI22_X1 port map( A1 => n6713, A2 => n3262, B1 => n15615, B2 => 
                           n11647, ZN => n26603);
   U1630 : NAND2_X1 port map( A1 => n11223, A2 => n7053, ZN => n2560);
   U1631 : INV_X1 port map( I => n121, ZN => n28012);
   U1638 : NOR3_X1 port map( A1 => n22454, A2 => n13306, A3 => n16086, ZN => 
                           n27508);
   U1641 : INV_X1 port map( I => n16191, ZN => n24081);
   U1642 : NOR2_X1 port map( A1 => n14519, A2 => n5362, ZN => n28011);
   U1643 : NAND2_X1 port map( A1 => n14218, A2 => n16278, ZN => n27666);
   U1644 : NOR2_X1 port map( A1 => n12035, A2 => n15812, ZN => n24388);
   U1645 : NOR2_X1 port map( A1 => n16113, A2 => n25570, ZN => n16114);
   U1648 : INV_X1 port map( I => n27002, ZN => n15984);
   U1651 : INV_X1 port map( I => n4522, ZN => n6647);
   U1656 : INV_X1 port map( I => n12271, ZN => n16011);
   U1658 : AND2_X1 port map( A1 => n561, A2 => n25365, Z => n16202);
   U1666 : BUF_X4 port map( I => n26814, Z => n26734);
   U1673 : NAND2_X2 port map( A1 => n9198, A2 => n11382, ZN => n11596);
   U1674 : INV_X2 port map( I => n17728, ZN => n10845);
   U1685 : BUF_X4 port map( I => n22643, Z => n13);
   U1686 : AOI22_X2 port map( A1 => n21592, A2 => n14679, B1 => n11490, B2 => 
                           n21593, ZN => n21383);
   U1690 : AOI21_X2 port map( A1 => n17632, A2 => n10845, B => n26610, ZN => 
                           n17633);
   U1691 : INV_X4 port map( I => n21792, ZN => n1023);
   U1697 : OAI21_X2 port map( A1 => n28401, A2 => n825, B => n17812, ZN => 
                           n5897);
   U1701 : NAND2_X2 port map( A1 => n5897, A2 => n885, ZN => n5896);
   U1702 : NOR2_X2 port map( A1 => n10474, A2 => n2398, ZN => n8248);
   U1704 : AOI22_X2 port map( A1 => n1701, A2 => n17520, B1 => n8263, B2 => 
                           n23105, ZN => n23739);
   U1710 : NAND2_X2 port map( A1 => n7350, A2 => n10941, ZN => n14872);
   U1719 : INV_X2 port map( I => n562, ZN => n12035);
   U1720 : NAND2_X2 port map( A1 => n11658, A2 => n9484, ZN => n9482);
   U1721 : OAI21_X2 port map( A1 => n16005, A2 => n16193, B => n14108, ZN => 
                           n27669);
   U1723 : AOI21_X2 port map( A1 => n913, A2 => n22529, B => n11503, ZN => 
                           n6268);
   U1731 : BUF_X4 port map( I => n562, Z => n5050);
   U1735 : NAND2_X2 port map( A1 => n6634, A2 => n20323, ZN => n1729);
   U1738 : NAND2_X2 port map( A1 => n15999, A2 => n26998, ZN => n3029);
   U1739 : INV_X2 port map( I => n24562, ZN => n4851);
   U1745 : OAI21_X2 port map( A1 => n882, A2 => n26317, B => n18491, ZN => 
                           n7607);
   U1746 : CLKBUF_X2 port map( I => n20982, Z => n27332);
   U1747 : INV_X1 port map( I => n12982, ZN => n14411);
   U1748 : OAI22_X1 port map( A1 => n19659, A2 => n28268, B1 => n5421, B2 => 
                           n12982, ZN => n19660);
   U1749 : INV_X1 port map( I => n21730, ZN => n851);
   U1752 : NAND2_X1 port map( A1 => n21730, A2 => n1079, ZN => n8897);
   U1756 : NOR2_X1 port map( A1 => n1079, A2 => n21730, ZN => n13416);
   U1757 : OAI22_X1 port map( A1 => n18840, A2 => n18839, B1 => n18896, B2 => 
                           n11577, ZN => n19428);
   U1758 : INV_X1 port map( I => n15004, ZN => n20982);
   U1764 : NOR2_X1 port map( A1 => n19590, A2 => n463, ZN => n9732);
   U1766 : AOI21_X1 port map( A1 => n19590, A2 => n5253, B => n1131, ZN => 
                           n27312);
   U1772 : NAND2_X1 port map( A1 => n20979, A2 => n15003, ZN => n7954);
   U1774 : NAND3_X1 port map( A1 => n2841, A2 => n2837, A3 => n2840, ZN => 
                           n23873);
   U1776 : NAND3_X1 port map( A1 => n9320, A2 => n9317, A3 => n9318, ZN => 
                           n27884);
   U1777 : NOR2_X1 port map( A1 => n21730, A2 => n10797, ZN => n2759);
   U1782 : NOR2_X1 port map( A1 => n1701, A2 => n17520, ZN => n12499);
   U1783 : NOR2_X1 port map( A1 => n950, A2 => n20933, ZN => n11306);
   U1784 : NAND2_X1 port map( A1 => n25238, A2 => n22046, ZN => n25863);
   U1799 : NAND2_X1 port map( A1 => n26974, A2 => n14606, ZN => n14605);
   U1800 : OAI21_X1 port map( A1 => n20848, A2 => n20849, B => n20847, ZN => 
                           n26974);
   U1802 : NAND2_X1 port map( A1 => n5931, A2 => n11048, ZN => n20158);
   U1809 : INV_X1 port map( I => n11048, ZN => n959);
   U1810 : AOI21_X1 port map( A1 => n20311, A2 => n11048, B => n13614, ZN => 
                           n13652);
   U1812 : NOR2_X1 port map( A1 => n10126, A2 => n8757, ZN => n22863);
   U1818 : NAND2_X1 port map( A1 => n20910, A2 => n3042, ZN => n15026);
   U1820 : NOR2_X1 port map( A1 => n20910, A2 => n26006, ZN => n20913);
   U1822 : INV_X2 port map( I => n12486, ZN => n20910);
   U1823 : OAI21_X1 port map( A1 => n7702, A2 => n11403, B => n20338, ZN => 
                           n5069);
   U1834 : NOR2_X1 port map( A1 => n6212, A2 => n28006, ZN => n1934);
   U1837 : NOR2_X1 port map( A1 => n7794, A2 => n755, ZN => n6212);
   U1838 : NOR2_X1 port map( A1 => n848, A2 => n4766, ZN => n4401);
   U1839 : NAND2_X1 port map( A1 => n6517, A2 => n11622, ZN => n21486);
   U1841 : OAI21_X1 port map( A1 => n21477, A2 => n21484, B => n11622, ZN => 
                           n11731);
   U1844 : NAND2_X1 port map( A1 => n20158, A2 => n20311, ZN => n6695);
   U1846 : NOR2_X1 port map( A1 => n19043, A2 => n28299, ZN => n28028);
   U1847 : NAND2_X1 port map( A1 => n10124, A2 => n27386, ZN => n9320);
   U1849 : INV_X1 port map( I => n11174, ZN => n6808);
   U1851 : NAND2_X1 port map( A1 => n2587, A2 => n3042, ZN => n2844);
   U1853 : NAND2_X1 port map( A1 => n20645, A2 => n723, ZN => n27261);
   U1855 : INV_X1 port map( I => n10666, ZN => n723);
   U1858 : NAND3_X1 port map( A1 => n17319, A2 => n17166, A3 => n25216, ZN => 
                           n13536);
   U1863 : NAND2_X1 port map( A1 => n24978, A2 => n21325, ZN => n21139);
   U1865 : CLKBUF_X2 port map( I => n21443, Z => n454);
   U1866 : NAND2_X1 port map( A1 => n2447, A2 => n21340, ZN => n21353);
   U1867 : OR2_X1 port map( A1 => n20099, A2 => n22843, Z => n24622);
   U1869 : OAI21_X1 port map( A1 => n18516, A2 => n13564, B => n22869, ZN => 
                           n2258);
   U1870 : NAND2_X1 port map( A1 => n18980, A2 => n26408, ZN => n18833);
   U1873 : NOR2_X1 port map( A1 => n11982, A2 => n26408, ZN => n11612);
   U1874 : CLKBUF_X1 port map( I => n19161, Z => n26408);
   U1875 : INV_X2 port map( I => n15706, ZN => n21780);
   U1876 : NAND2_X1 port map( A1 => n25240, A2 => n25239, ZN => n25238);
   U1880 : OAI21_X1 port map( A1 => n19731, A2 => n14726, B => n19846, ZN => 
                           n28298);
   U1885 : CLKBUF_X2 port map( I => n11842, Z => n22518);
   U1886 : CLKBUF_X2 port map( I => n26206, Z => n27846);
   U1891 : NAND2_X1 port map( A1 => n18939, A2 => n6889, ZN => n19156);
   U1894 : NAND2_X1 port map( A1 => n22800, A2 => n690, ZN => n25240);
   U1895 : OAI21_X1 port map( A1 => n22046, A2 => n22800, B => n13431, ZN => 
                           n15152);
   U1896 : OAI21_X1 port map( A1 => n21723, A2 => n21719, B => n28027, ZN => 
                           n27122);
   U1897 : NAND2_X1 port map( A1 => n21723, A2 => n21720, ZN => n21700);
   U1899 : OAI21_X1 port map( A1 => n21775, A2 => n10314, B => n773, ZN => 
                           n22045);
   U1900 : AOI21_X1 port map( A1 => n5357, A2 => n19841, B => n19844, ZN => 
                           n24771);
   U1901 : AOI21_X1 port map( A1 => n19737, A2 => n19844, B => n19739, ZN => 
                           n14823);
   U1904 : NOR2_X1 port map( A1 => n27690, A2 => n26738, ZN => n7328);
   U1910 : NAND2_X1 port map( A1 => n8299, A2 => n9042, ZN => n27690);
   U1912 : CLKBUF_X2 port map( I => n751, Z => n28071);
   U1916 : INV_X2 port map( I => n13477, ZN => n19844);
   U1917 : OAI22_X1 port map( A1 => n14307, A2 => n19878, B1 => n13477, B2 => 
                           n19877, ZN => n27962);
   U1919 : NAND2_X1 port map( A1 => n17920, A2 => n22244, ZN => n17921);
   U1927 : OAI21_X1 port map( A1 => n22622, A2 => n9298, B => n20165, ZN => 
                           n2834);
   U1928 : NOR3_X1 port map( A1 => n25870, A2 => n20165, A3 => n14176, ZN => 
                           n11355);
   U1929 : NAND2_X1 port map( A1 => n5367, A2 => n20868, ZN => n5532);
   U1933 : NAND2_X1 port map( A1 => n21564, A2 => n12797, ZN => n21567);
   U1936 : NOR2_X1 port map( A1 => n26422, A2 => n21711, ZN => n21706);
   U1938 : INV_X1 port map( I => n26422, ZN => n27248);
   U1939 : CLKBUF_X4 port map( I => n7971, Z => n26422);
   U1940 : NAND2_X1 port map( A1 => n3186, A2 => n1022, ZN => n8393);
   U1944 : NOR2_X1 port map( A1 => n21279, A2 => n13888, ZN => n3516);
   U1945 : CLKBUF_X2 port map( I => n18040, Z => n23375);
   U1959 : INV_X1 port map( I => n25222, ZN => n14684);
   U1962 : CLKBUF_X2 port map( I => n12181, Z => n28222);
   U1966 : INV_X1 port map( I => n26152, ZN => n24473);
   U1970 : NOR2_X1 port map( A1 => n26152, A2 => n18828, ZN => n18789);
   U1971 : NAND3_X1 port map( A1 => n22343, A2 => n20682, A3 => n20681, ZN => 
                           n26844);
   U1972 : NOR2_X1 port map( A1 => n27460, A2 => n2800, ZN => n9141);
   U1975 : BUF_X1 port map( I => n21641, Z => n23154);
   U1976 : AND2_X1 port map( A1 => n19730, A2 => n1128, Z => n10654);
   U1977 : NAND2_X1 port map( A1 => n6903, A2 => n8237, ZN => n5696);
   U1981 : OAI21_X1 port map( A1 => n6902, A2 => n6903, B => n24022, ZN => 
                           n23337);
   U1982 : NAND2_X1 port map( A1 => n11848, A2 => n7944, ZN => n13780);
   U1983 : NOR2_X1 port map( A1 => n26632, A2 => n27142, ZN => n24602);
   U1984 : NAND2_X1 port map( A1 => n26632, A2 => n27277, ZN => n22746);
   U1986 : NAND2_X1 port map( A1 => n3824, A2 => n2254, ZN => n8559);
   U1990 : NAND3_X1 port map( A1 => n1187, A2 => n5801, A3 => n18774, ZN => 
                           n8574);
   U1992 : OAI21_X1 port map( A1 => n26917, A2 => n26711, B => n21478, ZN => 
                           n11728);
   U1994 : NOR2_X1 port map( A1 => n11731, A2 => n21485, ZN => n26917);
   U1996 : CLKBUF_X4 port map( I => n21424, Z => n28278);
   U1997 : NAND2_X1 port map( A1 => n845, A2 => n13718, ZN => n12176);
   U1998 : INV_X1 port map( I => n20685, ZN => n25054);
   U1999 : NAND2_X1 port map( A1 => n20685, A2 => n12235, ZN => n20684);
   U2000 : NOR2_X1 port map( A1 => n19873, A2 => n5253, ZN => n19869);
   U2003 : INV_X2 port map( I => n20897, ZN => n25629);
   U2008 : OAI21_X1 port map( A1 => n25630, A2 => n20897, B => n20895, ZN => 
                           n20898);
   U2009 : OAI21_X1 port map( A1 => n20897, A2 => n22767, B => n20899, ZN => 
                           n14627);
   U2015 : OAI21_X1 port map( A1 => n21457, A2 => n13791, B => n24538, ZN => 
                           n11166);
   U2016 : NAND2_X1 port map( A1 => n7143, A2 => n13378, ZN => n5028);
   U2017 : NOR2_X1 port map( A1 => n7061, A2 => n14256, ZN => n13269);
   U2019 : INV_X2 port map( I => n14256, ZN => n734);
   U2021 : CLKBUF_X2 port map( I => n14256, Z => n25418);
   U2022 : CLKBUF_X4 port map( I => n21202, Z => n21457);
   U2023 : OAI21_X1 port map( A1 => n5516, A2 => n10209, B => n17401, ZN => 
                           n23557);
   U2024 : NOR2_X1 port map( A1 => n6051, A2 => n6052, ZN => n6406);
   U2025 : NAND2_X1 port map( A1 => n6589, A2 => n6052, ZN => n3650);
   U2027 : NAND3_X1 port map( A1 => n12176, A2 => n21710, A3 => n24922, ZN => 
                           n12175);
   U2029 : CLKBUF_X4 port map( I => n10359, Z => n6517);
   U2030 : OAI22_X1 port map( A1 => n3059, A2 => n14406, B1 => n13097, B2 => 
                           n21622, ZN => n25852);
   U2034 : CLKBUF_X1 port map( I => n10992, Z => n188);
   U2037 : NAND2_X1 port map( A1 => n11622, A2 => n21487, ZN => n8741);
   U2042 : NOR2_X1 port map( A1 => n10984, A2 => n722, ZN => n2163);
   U2047 : INV_X1 port map( I => n722, ZN => n772);
   U2049 : NOR3_X1 port map( A1 => n17401, A2 => n11113, A3 => n8692, ZN => 
                           n24795);
   U2050 : CLKBUF_X4 port map( I => n1715, Z => n491);
   U2051 : CLKBUF_X2 port map( I => n15209, Z => n22942);
   U2052 : NAND2_X1 port map( A1 => n705, A2 => n22738, ZN => n20956);
   U2055 : AOI22_X1 port map( A1 => n23088, A2 => n705, B1 => n20963, B2 => 
                           n4413, ZN => n15023);
   U2058 : CLKBUF_X4 port map( I => n20965, Z => n705);
   U2059 : NAND3_X1 port map( A1 => n27009, A2 => n21399, A3 => n21398, ZN => 
                           n21401);
   U2060 : NAND2_X1 port map( A1 => n15513, A2 => n8757, ZN => n23124);
   U2061 : CLKBUF_X2 port map( I => n21374, Z => n27604);
   U2062 : CLKBUF_X4 port map( I => n21054, Z => n13461);
   U2063 : OAI21_X1 port map( A1 => n27856, A2 => n9950, B => n19786, ZN => 
                           n26315);
   U2066 : NOR3_X1 port map( A1 => n9950, A2 => n27730, A3 => n22269, ZN => 
                           n11421);
   U2070 : NOR2_X1 port map( A1 => n9121, A2 => n9950, ZN => n26763);
   U2071 : CLKBUF_X2 port map( I => n13308, Z => n1515);
   U2073 : NOR2_X1 port map( A1 => n20070, A2 => n855, ZN => n8831);
   U2078 : AOI21_X1 port map( A1 => n17713, A2 => n23056, B => n17678, ZN => 
                           n17679);
   U2081 : INV_X2 port map( I => n23056, ZN => n2952);
   U2082 : BUF_X2 port map( I => n11785, Z => n7251);
   U2088 : NAND2_X1 port map( A1 => n9056, A2 => n7561, ZN => n23313);
   U2089 : OAI21_X1 port map( A1 => n9056, A2 => n10519, B => n9057, ZN => 
                           n21693);
   U2090 : CLKBUF_X1 port map( I => n10978, Z => n25979);
   U2092 : NOR2_X1 port map( A1 => n10978, A2 => n14343, ZN => n14170);
   U2093 : INV_X1 port map( I => n666, ZN => n10881);
   U2094 : INV_X1 port map( I => n20066, ZN => n11616);
   U2095 : AOI21_X1 port map( A1 => n22155, A2 => n22154, B => n18962, ZN => 
                           n19382);
   U2097 : NAND2_X1 port map( A1 => n6588, A2 => n24539, ZN => n27147);
   U2098 : NAND2_X1 port map( A1 => n20927, A2 => n24040, ZN => n9030);
   U2099 : NAND2_X1 port map( A1 => n15005, A2 => n27998, ZN => n20927);
   U2102 : NOR2_X1 port map( A1 => n21725, A2 => n3923, ZN => n6334);
   U2103 : NOR2_X1 port map( A1 => n28027, A2 => n21725, ZN => n28026);
   U2104 : BUF_X2 port map( I => n21638, Z => n438);
   U2105 : BUF_X2 port map( I => n8672, Z => n6802);
   U2106 : NAND2_X1 port map( A1 => n8672, A2 => n26422, ZN => n9943);
   U2107 : NAND2_X1 port map( A1 => n19779, A2 => n13194, ZN => n27011);
   U2109 : AND2_X1 port map( A1 => n19164, A2 => n24811, Z => n23559);
   U2110 : NAND2_X1 port map( A1 => n23577, A2 => n15539, ZN => n26801);
   U2111 : NAND3_X1 port map( A1 => n23577, A2 => n6910, A3 => n13698, ZN => 
                           n28439);
   U2112 : CLKBUF_X2 port map( I => n9734, Z => n23577);
   U2116 : NAND2_X1 port map( A1 => n5028, A2 => n774, ZN => n23071);
   U2117 : NAND3_X1 port map( A1 => n16853, A2 => n13593, A3 => n13592, ZN => 
                           n1790);
   U2124 : CLKBUF_X2 port map( I => n20770, Z => n28483);
   U2126 : INV_X1 port map( I => n5675, ZN => n28432);
   U2127 : CLKBUF_X2 port map( I => n25305, Z => n23864);
   U2128 : CLKBUF_X2 port map( I => n22000, Z => n26065);
   U2130 : INV_X1 port map( I => n21456, ZN => n26436);
   U2132 : CLKBUF_X4 port map( I => n21456, Z => n21620);
   U2133 : OAI21_X1 port map( A1 => n27318, A2 => n27317, B => n22794, ZN => 
                           n27009);
   U2135 : BUF_X2 port map( I => n20312, Z => n23700);
   U2140 : OAI22_X1 port map( A1 => n17905, A2 => n27550, B1 => n413, B2 => 
                           n25724, ZN => n14116);
   U2142 : INV_X1 port map( I => n413, ZN => n1213);
   U2143 : INV_X1 port map( I => n11961, ZN => n1112);
   U2148 : NAND2_X1 port map( A1 => n11961, A2 => n2525, ZN => n20311);
   U2151 : NAND2_X1 port map( A1 => n26970, A2 => n11961, ZN => n26969);
   U2153 : NOR2_X1 port map( A1 => n21564, A2 => n9934, ZN => n27119);
   U2155 : OAI21_X1 port map( A1 => n24574, A2 => n9934, B => n12797, ZN => 
                           n13127);
   U2157 : NOR2_X1 port map( A1 => n19630, A2 => n304, ZN => n19753);
   U2161 : CLKBUF_X1 port map( I => n304, Z => n24997);
   U2165 : INV_X1 port map( I => n7017, ZN => n1210);
   U2168 : AOI21_X1 port map( A1 => n5584, A2 => n7017, B => n1780, ZN => 
                           n28110);
   U2171 : NOR2_X1 port map( A1 => n18469, A2 => n11596, ZN => n13202);
   U2172 : INV_X1 port map( I => n11596, ZN => n15008);
   U2173 : NOR2_X1 port map( A1 => n7080, A2 => n18691, ZN => n18692);
   U2175 : NOR2_X1 port map( A1 => n9188, A2 => n8911, ZN => n4124);
   U2178 : AOI21_X1 port map( A1 => n24044, A2 => n27404, B => n10674, ZN => 
                           n21611);
   U2179 : NAND2_X1 port map( A1 => n11593, A2 => n24998, ZN => n10345);
   U2192 : NAND2_X1 port map( A1 => n11077, A2 => n6821, ZN => n20098);
   U2193 : NOR2_X1 port map( A1 => n9887, A2 => n25354, ZN => n9296);
   U2202 : NAND2_X1 port map( A1 => n26720, A2 => n5990, ZN => n13587);
   U2207 : AOI22_X1 port map( A1 => n375, A2 => n6013, B1 => n7879, B2 => 
                           n26720, ZN => n3480);
   U2211 : AOI21_X1 port map( A1 => n10595, A2 => n21716, B => n21781, ZN => 
                           n22204);
   U2213 : AOI21_X1 port map( A1 => n16585, A2 => n23907, B => n23758, ZN => 
                           n9726);
   U2215 : INV_X1 port map( I => n16585, ZN => n16671);
   U2220 : OR2_X1 port map( A1 => n23269, A2 => n15432, Z => n17226);
   U2223 : NAND4_X1 port map( A1 => n10842, A2 => n10668, A3 => n10840, A4 => 
                           n10841, ZN => n14779);
   U2229 : AOI21_X1 port map( A1 => n24997, A2 => n14671, B => n14279, ZN => 
                           n24861);
   U2233 : NAND2_X1 port map( A1 => n20868, A2 => n10578, ZN => n20462);
   U2235 : NAND2_X1 port map( A1 => n5532, A2 => n10578, ZN => n8495);
   U2236 : INV_X2 port map( I => n19918, ZN => n25236);
   U2238 : NOR3_X1 port map( A1 => n19866, A2 => n14282, A3 => n19918, ZN => 
                           n5263);
   U2242 : OAI21_X1 port map( A1 => n19918, A2 => n13854, B => n19866, ZN => 
                           n27059);
   U2243 : NAND2_X1 port map( A1 => n19917, A2 => n19918, ZN => n22082);
   U2250 : NOR2_X1 port map( A1 => n19918, A2 => n19917, ZN => n19865);
   U2251 : CLKBUF_X1 port map( I => n21118, Z => n28055);
   U2252 : NAND2_X1 port map( A1 => n10444, A2 => n11905, ZN => n11136);
   U2253 : INV_X1 port map( I => n13196, ZN => n25417);
   U2254 : NAND3_X1 port map( A1 => n2974, A2 => n13196, A3 => n3439, ZN => 
                           n2973);
   U2257 : NAND2_X1 port map( A1 => n11846, A2 => n22835, ZN => n13196);
   U2259 : INV_X1 port map( I => n22385, ZN => n18982);
   U2260 : NAND2_X1 port map( A1 => n22385, A2 => n11983, ZN => n26073);
   U2264 : AOI22_X1 port map( A1 => n26070, A2 => n22385, B1 => n5053, B2 => 
                           n24265, ZN => n15093);
   U2265 : CLKBUF_X4 port map( I => n20138, Z => n6470);
   U2266 : NOR2_X1 port map( A1 => n24951, A2 => n13444, ZN => n13638);
   U2270 : AOI22_X1 port map( A1 => n4038, A2 => n8576, B1 => n11414, B2 => 
                           n18633, ZN => n8575);
   U2273 : INV_X1 port map( I => n22050, ZN => n57);
   U2275 : INV_X2 port map( I => n19603, ZN => n974);
   U2276 : NOR2_X1 port map( A1 => n4246, A2 => n19603, ZN => n4247);
   U2278 : OAI21_X1 port map( A1 => n25149, A2 => n18476, B => n1800, ZN => 
                           n10147);
   U2280 : NOR2_X1 port map( A1 => n1800, A2 => n12569, ZN => n6439);
   U2282 : INV_X1 port map( I => n19734, ZN => n19872);
   U2286 : CLKBUF_X2 port map( I => n19734, Z => n14789);
   U2288 : CLKBUF_X2 port map( I => n20222, Z => n23374);
   U2289 : NOR2_X1 port map( A1 => n20222, A2 => n19999, ZN => n20000);
   U2291 : NOR2_X1 port map( A1 => n26456, A2 => n20222, ZN => n27642);
   U2296 : INV_X1 port map( I => n20222, ZN => n13294);
   U2297 : NAND2_X1 port map( A1 => n20219, A2 => n20222, ZN => n3958);
   U2301 : NAND2_X1 port map( A1 => n1159, A2 => n13873, ZN => n27894);
   U2302 : INV_X2 port map( I => n13873, ZN => n13872);
   U2304 : INV_X1 port map( I => n8468, ZN => n20818);
   U2305 : NAND2_X1 port map( A1 => n2450, A2 => n2448, ZN => n2449);
   U2309 : CLKBUF_X2 port map( I => n21355, Z => n2448);
   U2311 : NAND2_X1 port map( A1 => n19676, A2 => n13167, ZN => n26601);
   U2314 : CLKBUF_X2 port map( I => n14194, Z => n23540);
   U2317 : INV_X1 port map( I => n22760, ZN => n11676);
   U2318 : CLKBUF_X1 port map( I => n19150, Z => n28303);
   U2320 : NOR2_X1 port map( A1 => n11080, A2 => n11, ZN => n15966);
   U2321 : OAI21_X1 port map( A1 => n11080, A2 => n16076, B => n10905, ZN => 
                           n15906);
   U2322 : NOR2_X1 port map( A1 => n11080, A2 => n16348, ZN => n16349);
   U2325 : NAND2_X1 port map( A1 => n28468, A2 => n5616, ZN => n20210);
   U2326 : CLKBUF_X2 port map( I => n8468, Z => n25927);
   U2327 : NAND2_X1 port map( A1 => n4782, A2 => n4537, ZN => n11629);
   U2329 : INV_X1 port map( I => n27291, ZN => n17296);
   U2331 : NAND2_X1 port map( A1 => n26400, A2 => n4556, ZN => n10780);
   U2338 : NOR2_X1 port map( A1 => n16640, A2 => n4556, ZN => n16405);
   U2341 : OAI21_X1 port map( A1 => n1255, A2 => n4556, B => n16597, ZN => 
                           n22436);
   U2348 : CLKBUF_X1 port map( I => n14795, Z => n27594);
   U2352 : AOI22_X1 port map( A1 => n21361, A2 => n10541, B1 => n21543, B2 => 
                           n21360, ZN => n24433);
   U2354 : INV_X2 port map( I => n21544, ZN => n10541);
   U2360 : CLKBUF_X2 port map( I => n6364, Z => n5801);
   U2365 : OR2_X1 port map( A1 => n6364, A2 => n23203, Z => n18622);
   U2370 : INV_X1 port map( I => n6364, ZN => n27887);
   U2373 : NAND2_X1 port map( A1 => n8810, A2 => n20107, ZN => n12524);
   U2376 : OR2_X1 port map( A1 => n4664, A2 => n19694, Z => n24600);
   U2383 : NOR2_X1 port map( A1 => n2398, A2 => n7533, ZN => n18825);
   U2387 : NAND2_X1 port map( A1 => n7533, A2 => n2398, ZN => n1335);
   U2389 : OAI22_X1 port map( A1 => n1030, A2 => n17415, B1 => n14250, B2 => 
                           n9865, ZN => n6368);
   U2390 : INV_X1 port map( I => n8963, ZN => n14666);
   U2394 : CLKBUF_X2 port map( I => n8963, Z => n27380);
   U2397 : BUF_X2 port map( I => n15447, Z => n26443);
   U2398 : NOR2_X1 port map( A1 => n26546, A2 => n26547, ZN => n18958);
   U2400 : NOR2_X1 port map( A1 => n27548, A2 => n18474, ZN => n7675);
   U2406 : INV_X1 port map( I => n21536, ZN => n24904);
   U2407 : OAI21_X1 port map( A1 => n21530, A2 => n21536, B => n21531, ZN => 
                           n21521);
   U2408 : NOR2_X1 port map( A1 => n27359, A2 => n4802, ZN => n11157);
   U2412 : INV_X2 port map( I => n5425, ZN => n4802);
   U2416 : INV_X1 port map( I => n3525, ZN => n11846);
   U2418 : OAI21_X1 port map( A1 => n11870, A2 => n20096, B => n3525, ZN => 
                           n3535);
   U2420 : NAND2_X1 port map( A1 => n3525, A2 => n11871, ZN => n20097);
   U2421 : INV_X2 port map( I => n7346, ZN => n13299);
   U2424 : INV_X2 port map( I => n5373, ZN => n7023);
   U2427 : BUF_X2 port map( I => n5373, Z => n443);
   U2429 : CLKBUF_X2 port map( I => n18410, Z => n13646);
   U2431 : NAND2_X1 port map( A1 => n18791, A2 => n12584, ZN => n19061);
   U2441 : NAND3_X1 port map( A1 => n27736, A2 => n18573, A3 => n18791, ZN => 
                           n3239);
   U2442 : INV_X1 port map( I => n18791, ZN => n13597);
   U2443 : NAND2_X1 port map( A1 => n18791, A2 => n23575, ZN => n19123);
   U2447 : CLKBUF_X2 port map( I => n21609, Z => n24044);
   U2450 : NOR2_X1 port map( A1 => n21606, A2 => n21609, ZN => n21603);
   U2452 : INV_X1 port map( I => n17388, ZN => n17355);
   U2456 : CLKBUF_X2 port map( I => n17388, Z => n13766);
   U2457 : NAND2_X1 port map( A1 => n17400, A2 => n17318, ZN => n1902);
   U2458 : NAND2_X1 port map( A1 => n11487, A2 => n24998, ZN => n19956);
   U2459 : AOI22_X1 port map( A1 => n16594, A2 => n741, B1 => n16593, B2 => 
                           n9379, ZN => n16595);
   U2462 : AOI21_X1 port map( A1 => n23663, A2 => n19156, B => n19157, ZN => 
                           n6887);
   U2463 : NAND2_X1 port map( A1 => n19157, A2 => n19154, ZN => n19025);
   U2470 : NOR2_X1 port map( A1 => n19157, A2 => n6487, ZN => n15486);
   U2474 : NOR2_X1 port map( A1 => n19157, A2 => n19154, ZN => n8045);
   U2479 : INV_X2 port map( I => n14237, ZN => n19157);
   U2480 : NOR2_X1 port map( A1 => n8594, A2 => n27416, ZN => n3821);
   U2482 : NOR2_X1 port map( A1 => n27416, A2 => n28553, ZN => n8491);
   U2485 : OR2_X1 port map( A1 => n19845, A2 => n19849, Z => n10023);
   U2487 : INV_X1 port map( I => n20207, ZN => n1955);
   U2488 : NAND2_X1 port map( A1 => n5616, A2 => n2023, ZN => n20084);
   U2490 : NAND2_X1 port map( A1 => n26636, A2 => n5796, ZN => n20986);
   U2494 : NAND3_X1 port map( A1 => n10963, A2 => n20226, A3 => n20225, ZN => 
                           n10940);
   U2497 : AOI21_X1 port map( A1 => n10963, A2 => n20226, B => n20225, ZN => 
                           n27663);
   U2498 : INV_X2 port map( I => n20226, ZN => n20474);
   U2500 : OAI21_X1 port map( A1 => n2767, A2 => n12250, B => n20226, ZN => 
                           n28410);
   U2509 : INV_X1 port map( I => n10627, ZN => n9934);
   U2512 : CLKBUF_X4 port map( I => n10627, Z => n28308);
   U2517 : INV_X1 port map( I => n16485, ZN => n2696);
   U2518 : NAND2_X1 port map( A1 => n6952, A2 => n26710, ZN => n19988);
   U2520 : NOR2_X1 port map( A1 => n6952, A2 => n23906, ZN => n19875);
   U2522 : INV_X1 port map( I => n17850, ZN => n18640);
   U2523 : BUF_X2 port map( I => n17850, Z => n18747);
   U2527 : AND2_X1 port map( A1 => n13349, A2 => n7390, Z => n21919);
   U2528 : INV_X1 port map( I => n7390, ZN => n18797);
   U2529 : NAND2_X1 port map( A1 => n7390, A2 => n25319, ZN => n18522);
   U2532 : AOI21_X1 port map( A1 => n28255, A2 => n19036, B => n7390, ZN => 
                           n9312);
   U2534 : INV_X1 port map( I => n28176, ZN => n26557);
   U2535 : NAND2_X1 port map( A1 => n23450, A2 => n25573, ZN => n10811);
   U2538 : OAI21_X1 port map( A1 => n25573, A2 => n287, B => n10811, ZN => 
                           n20276);
   U2539 : AOI21_X1 port map( A1 => n4660, A2 => n20217, B => n25573, ZN => 
                           n24934);
   U2540 : AOI21_X1 port map( A1 => n4296, A2 => n4295, B => n16704, ZN => 
                           n3133);
   U2542 : NOR2_X1 port map( A1 => n25834, A2 => n16704, ZN => n26310);
   U2544 : NAND3_X1 port map( A1 => n16702, A2 => n4295, A3 => n16704, ZN => 
                           n16153);
   U2545 : NAND2_X1 port map( A1 => n16704, A2 => n12839, ZN => n3196);
   U2547 : NAND2_X1 port map( A1 => n1491, A2 => n22842, ZN => n6210);
   U2550 : INV_X1 port map( I => n6959, ZN => n11328);
   U2558 : NAND2_X1 port map( A1 => n11905, A2 => n13049, ZN => n9003);
   U2560 : NAND2_X1 port map( A1 => n825, A2 => n2910, ZN => n8169);
   U2561 : NAND2_X1 port map( A1 => n22337, A2 => n17920, ZN => n17642);
   U2564 : NOR2_X1 port map( A1 => n10941, A2 => n7350, ZN => n14120);
   U2567 : NAND2_X1 port map( A1 => n18512, A2 => n7350, ZN => n27729);
   U2569 : OAI22_X1 port map( A1 => n10322, A2 => n25935, B1 => n879, B2 => 
                           n7350, ZN => n11088);
   U2573 : OAI21_X1 port map( A1 => n27895, A2 => n18556, B => n27710, ZN => 
                           n3699);
   U2581 : INV_X2 port map( I => n27710, ZN => n18706);
   U2584 : INV_X1 port map( I => n2777, ZN => n21682);
   U2585 : AOI21_X1 port map( A1 => n22244, A2 => n24563, B => n17920, ZN => 
                           n17581);
   U2588 : INV_X2 port map( I => n24563, ZN => n22337);
   U2590 : NAND2_X1 port map( A1 => n24563, A2 => n17580, ZN => n17922);
   U2592 : NAND2_X1 port map( A1 => n17956, A2 => n5402, ZN => n4779);
   U2594 : NOR2_X1 port map( A1 => n10673, A2 => n5402, ZN => n14034);
   U2598 : AND2_X1 port map( A1 => n10764, A2 => n2544, Z => n20416);
   U2601 : NOR2_X1 port map( A1 => n1349, A2 => n7599, ZN => n13237);
   U2605 : BUF_X2 port map( I => n5243, Z => n4938);
   U2606 : BUF_X2 port map( I => n16810, Z => n23505);
   U2608 : NAND2_X1 port map( A1 => n16810, A2 => n12224, ZN => n16554);
   U2611 : NAND2_X1 port map( A1 => n16555, A2 => n16810, ZN => n13261);
   U2612 : NAND2_X1 port map( A1 => n22796, A2 => n6473, ZN => n21080);
   U2613 : CLKBUF_X2 port map( I => n2656, Z => n28468);
   U2614 : CLKBUF_X2 port map( I => n19365, Z => n25941);
   U2621 : NAND2_X1 port map( A1 => n27895, A2 => n27026, ZN => n15398);
   U2624 : AOI22_X1 port map( A1 => n8113, A2 => n15399, B1 => n18704, B2 => 
                           n27026, ZN => n27717);
   U2626 : INV_X1 port map( I => n8912, ZN => n4689);
   U2627 : CLKBUF_X1 port map( I => n5682, Z => n24887);
   U2632 : NAND2_X1 port map( A1 => n694, A2 => n21481, ZN => n24213);
   U2637 : NOR2_X1 port map( A1 => n21481, A2 => n694, ZN => n21485);
   U2639 : INV_X2 port map( I => n11053, ZN => n694);
   U2642 : OAI22_X1 port map( A1 => n9919, A2 => n20145, B1 => n25294, B2 => 
                           n20070, ZN => n15066);
   U2643 : OAI22_X1 port map( A1 => n20145, A2 => n12475, B1 => n26140, B2 => 
                           n20073, ZN => n15065);
   U2646 : NAND2_X1 port map( A1 => n20145, A2 => n4225, ZN => n20075);
   U2649 : INV_X2 port map( I => n19967, ZN => n20145);
   U2653 : CLKBUF_X4 port map( I => n2016, Z => n28263);
   U2654 : INV_X1 port map( I => n5920, ZN => n4357);
   U2660 : NAND2_X1 port map( A1 => n28108, A2 => n16557, ZN => n24124);
   U2661 : NAND2_X1 port map( A1 => n16558, A2 => n16557, ZN => n11604);
   U2663 : INV_X1 port map( I => n2467, ZN => n19298);
   U2672 : BUF_X2 port map( I => n6779, Z => n2285);
   U2678 : INV_X1 port map( I => n6779, ZN => n17683);
   U2679 : INV_X2 port map( I => n22840, ZN => n832);
   U2680 : NOR2_X1 port map( A1 => n18473, A2 => n7770, ZN => n28422);
   U2683 : NAND2_X1 port map( A1 => n7769, A2 => n7770, ZN => n27548);
   U2687 : NOR2_X1 port map( A1 => n24286, A2 => n7770, ZN => n4552);
   U2701 : NAND2_X1 port map( A1 => n8354, A2 => n7770, ZN => n26885);
   U2706 : NOR3_X1 port map( A1 => n24286, A2 => n18602, A3 => n7770, ZN => 
                           n26870);
   U2707 : INV_X1 port map( I => n7364, ZN => n28154);
   U2709 : INV_X1 port map( I => n16288, ZN => n6428);
   U2710 : OAI22_X1 port map( A1 => n5497, A2 => n24881, B1 => n17918, B2 => 
                           n11419, ZN => n17644);
   U2714 : AOI21_X1 port map( A1 => n22536, A2 => n23753, B => n10477, ZN => 
                           n27140);
   U2715 : INV_X2 port map( I => n17495, ZN => n740);
   U2718 : NOR2_X1 port map( A1 => n17556, A2 => n17495, ZN => n4403);
   U2722 : OAI21_X1 port map( A1 => n17554, A2 => n14062, B => n17495, ZN => 
                           n3649);
   U2723 : BUF_X2 port map( I => n27877, Z => n16262);
   U2724 : NOR2_X1 port map( A1 => n15169, A2 => n21702, ZN => n15168);
   U2731 : NAND2_X1 port map( A1 => n21702, A2 => n13432, ZN => n26829);
   U2732 : OAI21_X1 port map( A1 => n11032, A2 => n11031, B => n21702, ZN => 
                           n12588);
   U2733 : NOR2_X1 port map( A1 => n16261, A2 => n16262, ZN => n24898);
   U2734 : NOR2_X1 port map( A1 => n16262, A2 => n16230, ZN => n16232);
   U2737 : NAND2_X1 port map( A1 => n671, A2 => n19586, ZN => n27305);
   U2740 : NOR2_X1 port map( A1 => n6427, A2 => n577, ZN => n13326);
   U2750 : OAI21_X1 port map( A1 => n16293, A2 => n577, B => n16292, ZN => 
                           n16295);
   U2755 : INV_X1 port map( I => n577, ZN => n28033);
   U2756 : CLKBUF_X1 port map( I => n17475, Z => n27073);
   U2761 : INV_X2 port map( I => n15586, ZN => n19768);
   U2762 : OAI21_X1 port map( A1 => n14192, A2 => n14191, B => n15586, ZN => 
                           n28522);
   U2763 : CLKBUF_X2 port map( I => n15586, Z => n28134);
   U2764 : NOR3_X1 port map( A1 => n19808, A2 => n7767, A3 => n28285, ZN => 
                           n6231);
   U2768 : AOI21_X1 port map( A1 => n7767, A2 => n19808, B => n24146, ZN => 
                           n1938);
   U2773 : NAND2_X1 port map( A1 => n19808, A2 => n28111, ZN => n27346);
   U2774 : INV_X1 port map( I => n704, ZN => n7176);
   U2779 : AOI21_X1 port map( A1 => n22609, A2 => n15227, B => n28459, ZN => 
                           n27340);
   U2782 : NAND3_X1 port map( A1 => n20855, A2 => n24040, A3 => n26924, ZN => 
                           n20813);
   U2784 : CLKBUF_X1 port map( I => n20852, Z => n26924);
   U2789 : INV_X1 port map( I => n20596, ZN => n12290);
   U2799 : CLKBUF_X4 port map( I => n20596, Z => n21719);
   U2801 : BUF_X2 port map( I => n17868, Z => n28322);
   U2802 : NAND2_X1 port map( A1 => n22307, A2 => n17868, ZN => n22306);
   U2825 : CLKBUF_X2 port map( I => n15414, Z => n4738);
   U2827 : CLKBUF_X1 port map( I => n4064, Z => n28300);
   U2829 : AOI22_X1 port map( A1 => n1908, A2 => n1881, B1 => n14644, B2 => 
                           n1866, ZN => n1865);
   U2831 : NAND2_X1 port map( A1 => n14571, A2 => n14644, ZN => n26950);
   U2835 : NAND2_X1 port map( A1 => n524, A2 => n14644, ZN => n9438);
   U2836 : CLKBUF_X4 port map( I => n7169, Z => n2445);
   U2838 : INV_X2 port map( I => n7169, ZN => n18628);
   U2839 : NAND2_X1 port map( A1 => n19035, A2 => n209, ZN => n5875);
   U2840 : OAI21_X1 port map( A1 => n15116, A2 => n15114, B => n19675, ZN => 
                           n15113);
   U2842 : OAI22_X1 port map( A1 => n19675, A2 => n19702, B1 => n13797, B2 => 
                           n4565, ZN => n4564);
   U2845 : NAND2_X1 port map( A1 => n60, A2 => n8344, ZN => n15879);
   U2847 : INV_X2 port map( I => n13461, ZN => n1078);
   U2848 : OAI21_X1 port map( A1 => n21056, A2 => n13461, B => n22505, ZN => 
                           n9851);
   U2850 : NAND2_X1 port map( A1 => n12066, A2 => n13461, ZN => n22505);
   U2852 : NOR2_X1 port map( A1 => n13461, A2 => n12309, ZN => n2094);
   U2857 : NOR2_X1 port map( A1 => n13461, A2 => n12067, ZN => n27094);
   U2858 : CLKBUF_X2 port map( I => n24331, Z => n27528);
   U2859 : NAND2_X1 port map( A1 => n19143, A2 => n19144, ZN => n19145);
   U2860 : NAND2_X1 port map( A1 => n8717, A2 => n8968, ZN => n8755);
   U2864 : INV_X2 port map( I => n8717, ZN => n14565);
   U2865 : NAND2_X1 port map( A1 => n28268, A2 => n8717, ZN => n8949);
   U2870 : NOR3_X1 port map( A1 => n19823, A2 => n19720, A3 => n28377, ZN => 
                           n28523);
   U2873 : NOR2_X1 port map( A1 => n13926, A2 => n19720, ZN => n12894);
   U2876 : NOR2_X1 port map( A1 => n18370, A2 => n10206, ZN => n11186);
   U2877 : NAND2_X1 port map( A1 => n18370, A2 => n10206, ZN => n4883);
   U2879 : INV_X2 port map( I => n18370, ZN => n1015);
   U2885 : INV_X1 port map( I => n9880, ZN => n27907);
   U2886 : NAND2_X1 port map( A1 => n2523, A2 => n15953, ZN => n21957);
   U2887 : CLKBUF_X2 port map( I => n9702, Z => n6354);
   U2892 : INV_X1 port map( I => n9702, ZN => n6046);
   U2894 : INV_X1 port map( I => n8472, ZN => n17963);
   U2897 : CLKBUF_X4 port map( I => n8472, Z => n23979);
   U2900 : INV_X1 port map( I => n8985, ZN => n17475);
   U2901 : CLKBUF_X2 port map( I => n8985, Z => n26754);
   U2902 : NAND2_X1 port map( A1 => n14788, A2 => n17845, ZN => n22492);
   U2903 : OAI21_X1 port map( A1 => n17993, A2 => n17994, B => n14788, ZN => 
                           n11283);
   U2905 : OAI22_X1 port map( A1 => n14788, A2 => n17605, B1 => n17845, B2 => 
                           n6644, ZN => n6643);
   U2908 : BUF_X1 port map( I => n24070, Z => n27201);
   U2915 : NAND2_X1 port map( A1 => n24070, A2 => n9224, ZN => n27291);
   U2923 : NAND2_X1 port map( A1 => n17452, A2 => n24070, ZN => n17211);
   U2925 : INV_X2 port map( I => n17843, ZN => n1893);
   U2927 : BUF_X2 port map( I => n17843, Z => n2403);
   U2929 : NAND2_X1 port map( A1 => n28400, A2 => n6110, ZN => n7690);
   U2930 : OR2_X1 port map( A1 => n6110, A2 => n24812, Z => n2422);
   U2932 : INV_X1 port map( I => n19231, ZN => n19355);
   U2937 : NOR2_X1 port map( A1 => n11988, A2 => n14391, ZN => n24854);
   U2940 : INV_X1 port map( I => n21315, ZN => n26958);
   U2941 : NAND2_X1 port map( A1 => n22828, A2 => n27450, ZN => n4121);
   U2944 : OAI21_X1 port map( A1 => n22828, A2 => n24576, B => n6509, ZN => 
                           n7772);
   U2946 : BUF_X2 port map( I => n10104, Z => n22823);
   U2951 : INV_X1 port map( I => n10104, ZN => n15697);
   U2954 : INV_X1 port map( I => n20367, ZN => n21627);
   U2956 : CLKBUF_X2 port map( I => n20367, Z => n21623);
   U2958 : INV_X1 port map( I => n16007, ZN => n15864);
   U2959 : BUF_X2 port map( I => n16007, Z => n14519);
   U2962 : NAND2_X2 port map( A1 => n9116, A2 => n16455, ZN => n7237);
   U2964 : NOR2_X2 port map( A1 => n5353, A2 => n26213, ZN => n3547);
   U2974 : INV_X2 port map( I => n9070, ZN => n10461);
   U2978 : INV_X1 port map( I => n16406, ZN => n1228);
   U2981 : CLKBUF_X4 port map( I => n16406, Z => n17501);
   U2982 : BUF_X2 port map( I => n3963, Z => n3741);
   U2986 : XOR2_X1 port map( A1 => n575, A2 => n16955, Z => n26628);
   U2987 : INV_X2 port map( I => n10856, ZN => n23072);
   U2988 : AND3_X2 port map( A1 => n1031, A2 => n24560, A3 => n9827, Z => 
                           n26629);
   U2991 : INV_X2 port map( I => n12275, ZN => n27854);
   U2997 : NAND2_X2 port map( A1 => n17690, A2 => n17689, ZN => n18226);
   U2998 : NAND2_X2 port map( A1 => n17690, A2 => n17689, ZN => n27459);
   U3000 : AND2_X1 port map( A1 => n13547, A2 => n12494, Z => n26630);
   U3002 : AOI22_X2 port map( A1 => n23418, A2 => n25903, B1 => n17714, B2 => 
                           n17715, ZN => n9802);
   U3005 : AND2_X2 port map( A1 => n12493, A2 => n18388, Z => n26631);
   U3008 : INV_X2 port map( I => n27647, ZN => n27671);
   U3013 : INV_X4 port map( I => n27044, ZN => n28444);
   U3018 : INV_X4 port map( I => n18683, ZN => n18465);
   U3019 : NOR2_X1 port map( A1 => n23772, A2 => n27044, ZN => n26632);
   U3021 : NAND2_X2 port map( A1 => n7673, A2 => n7676, ZN => n27432);
   U3022 : NAND2_X2 port map( A1 => n12433, A2 => n12432, ZN => n27400);
   U3023 : INV_X1 port map( I => n15564, ZN => n19843);
   U3024 : BUF_X2 port map( I => n15564, Z => n14307);
   U3030 : INV_X1 port map( I => n26620, ZN => n10562);
   U3032 : XNOR2_X1 port map( A1 => n19066, A2 => n19067, ZN => n26633);
   U3038 : NOR2_X2 port map( A1 => n7388, A2 => n12643, ZN => n4858);
   U3041 : OR2_X2 port map( A1 => n12364, A2 => n3101, Z => n26635);
   U3042 : INV_X2 port map( I => n687, ZN => n27023);
   U3044 : XNOR2_X1 port map( A1 => n12860, A2 => n12474, ZN => n26636);
   U3047 : AOI21_X2 port map( A1 => n25695, A2 => n26007, B => n20024, ZN => 
                           n6535);
   U3048 : AND2_X2 port map( A1 => n19981, A2 => n2185, Z => n26637);
   U3053 : INV_X4 port map( I => n21091, ZN => n944);
   U3056 : INV_X2 port map( I => n20751, ZN => n26914);
   U3058 : INV_X2 port map( I => n15734, ZN => n11183);
   U3060 : NAND2_X2 port map( A1 => n27643, A2 => n24919, ZN => n27396);
   U3064 : INV_X1 port map( I => n26651, ZN => n12391);
   U3065 : NOR2_X2 port map( A1 => n15314, A2 => n20408, ZN => n27429);
   U3072 : NAND3_X2 port map( A1 => n10040, A2 => n3855, A3 => n10174, ZN => 
                           n6182);
   U3074 : CLKBUF_X4 port map( I => n16012, Z => n12272);
   U3075 : OR2_X2 port map( A1 => n6485, A2 => n21082, Z => n2052);
   U3077 : NAND2_X1 port map( A1 => n25952, A2 => n6485, ZN => n8137);
   U3079 : AOI21_X1 port map( A1 => n12066, A2 => n21100, B => n13461, ZN => 
                           n12307);
   U3080 : NAND2_X1 port map( A1 => n13461, A2 => n21055, ZN => n26984);
   U3083 : NAND2_X1 port map( A1 => n10558, A2 => n13461, ZN => n6962);
   U3084 : NAND2_X1 port map( A1 => n27965, A2 => n9216, ZN => n4844);
   U3085 : NAND2_X1 port map( A1 => n16433, A2 => n12331, ZN => n4553);
   U3087 : CLKBUF_X2 port map( I => n6543, Z => n25315);
   U3088 : NOR2_X1 port map( A1 => n4898, A2 => n22337, ZN => n5497);
   U3091 : OR2_X2 port map( A1 => n17582, A2 => n4898, Z => n6207);
   U3093 : OR2_X2 port map( A1 => n11733, A2 => n4462, Z => n11137);
   U3101 : CLKBUF_X4 port map( I => n15835, Z => n15986);
   U3105 : OAI21_X1 port map( A1 => n8232, A2 => n8233, B => n7518, ZN => 
                           n28398);
   U3107 : OAI21_X1 port map( A1 => n7518, A2 => n20593, B => n12406, ZN => 
                           n20821);
   U3112 : NOR2_X1 port map( A1 => n953, A2 => n7518, ZN => n9134);
   U3116 : NAND2_X1 port map( A1 => n14113, A2 => n7518, ZN => n25881);
   U3127 : NAND2_X1 port map( A1 => n7807, A2 => n7518, ZN => n12406);
   U3129 : INV_X2 port map( I => n7518, ZN => n9179);
   U3131 : AOI21_X1 port map( A1 => n817, A2 => n19167, B => n26720, ZN => n375
                           );
   U3132 : INV_X2 port map( I => n7569, ZN => n19106);
   U3133 : CLKBUF_X4 port map( I => n7569, Z => n1658);
   U3136 : INV_X2 port map( I => n19689, ZN => n10937);
   U3137 : OAI21_X1 port map( A1 => n11454, A2 => n19689, B => n14929, ZN => 
                           n8794);
   U3138 : NOR2_X1 port map( A1 => n19689, A2 => n14929, ZN => n10956);
   U3142 : NAND3_X1 port map( A1 => n19435, A2 => n19211, A3 => n19210, ZN => 
                           n12545);
   U3144 : AOI22_X1 port map( A1 => n3820, A2 => n22811, B1 => n3821, B2 => 
                           n20732, ZN => n23765);
   U3145 : INV_X1 port map( I => n20732, ZN => n27923);
   U3146 : INV_X1 port map( I => n13469, ZN => n11103);
   U3150 : NAND2_X1 port map( A1 => n14320, A2 => n7281, ZN => n16515);
   U3151 : AND2_X2 port map( A1 => n12340, A2 => n24234, Z => n13570);
   U3154 : CLKBUF_X12 port map( I => Key(137), Z => n21010);
   U3156 : NOR2_X1 port map( A1 => n1111, A2 => n11854, ZN => n11786);
   U3157 : NOR2_X1 port map( A1 => n14255, A2 => n9772, ZN => n17598);
   U3158 : INV_X1 port map( I => n16639, ZN => n16599);
   U3162 : AOI21_X1 port map( A1 => n20619, A2 => n22766, B => n26765, ZN => 
                           n10273);
   U3164 : NOR3_X1 port map( A1 => n939, A2 => n22766, A3 => n20623, ZN => 
                           n26765);
   U3165 : INV_X1 port map( I => n18950, ZN => n9215);
   U3166 : CLKBUF_X12 port map( I => n21304, Z => n27169);
   U3169 : NOR2_X1 port map( A1 => n11609, A2 => n15222, ZN => n9631);
   U3172 : INV_X1 port map( I => n8132, ZN => n6273);
   U3180 : INV_X1 port map( I => n12600, ZN => n22544);
   U3183 : CLKBUF_X12 port map( I => n8627, Z => n8073);
   U3185 : BUF_X2 port map( I => n3490, Z => n26638);
   U3191 : NAND2_X1 port map( A1 => n3932, A2 => n10362, ZN => n18896);
   U3193 : NAND3_X1 port map( A1 => n13873, A2 => n13028, A3 => n13371, ZN => 
                           n18821);
   U3197 : NAND2_X1 port map( A1 => n26008, A2 => n3729, ZN => n27896);
   U3199 : NAND2_X1 port map( A1 => n4556, A2 => n26008, ZN => n16026);
   U3203 : INV_X2 port map( I => n26008, ZN => n1255);
   U3207 : INV_X2 port map( I => n11497, ZN => n9330);
   U3208 : NAND2_X1 port map( A1 => n6051, A2 => n6589, ZN => n20711);
   U3210 : AOI21_X1 port map( A1 => n12644, A2 => n12364, B => n23253, ZN => 
                           n7933);
   U3218 : INV_X1 port map( I => n12364, ZN => n11259);
   U3223 : CLKBUF_X12 port map( I => n4762, Z => n4750);
   U3224 : CLKBUF_X4 port map( I => n4826, Z => n26639);
   U3226 : CLKBUF_X4 port map( I => n4265, Z => n26640);
   U3240 : CLKBUF_X12 port map( I => n4265, Z => n26641);
   U3241 : AND2_X2 port map( A1 => n2895, A2 => n2897, Z => n24292);
   U3242 : CLKBUF_X12 port map( I => n2897, Z => n27763);
   U3248 : OR2_X2 port map( A1 => n14224, A2 => n15354, Z => n9098);
   U3249 : INV_X1 port map( I => n18227, ZN => n18241);
   U3252 : INV_X1 port map( I => n18090, ZN => n27633);
   U3253 : OR2_X1 port map( A1 => n19016, A2 => n14338, Z => n21915);
   U3254 : BUF_X2 port map( I => n19016, Z => n23431);
   U3256 : INV_X2 port map( I => n19016, ZN => n11331);
   U3264 : NOR2_X1 port map( A1 => n10543, A2 => n22572, ZN => n27653);
   U3266 : NOR3_X1 port map( A1 => n3090, A2 => n3091, A3 => n14990, ZN => 
                           n11609);
   U3268 : AOI22_X1 port map( A1 => n3090, A2 => n14990, B1 => n9370, B2 => 
                           n15592, ZN => n23756);
   U3269 : NAND2_X1 port map( A1 => n17007, A2 => n14990, ZN => n8442);
   U3276 : AOI22_X1 port map( A1 => n17007, A2 => n717, B1 => n193, B2 => 
                           n14990, ZN => n27125);
   U3277 : NAND2_X1 port map( A1 => n17915, A2 => n17912, ZN => n22628);
   U3280 : NAND2_X1 port map( A1 => n21943, A2 => n17912, ZN => n11651);
   U3281 : AND2_X2 port map( A1 => n7587, A2 => n7870, Z => n3959);
   U3283 : INV_X1 port map( I => n12413, ZN => n14718);
   U3284 : NAND2_X1 port map( A1 => n9051, A2 => n14737, ZN => n24902);
   U3287 : INV_X2 port map( I => n14737, ZN => n887);
   U3290 : INV_X2 port map( I => n19775, ZN => n775);
   U3292 : OAI21_X1 port map( A1 => n23026, A2 => n19775, B => n25650, ZN => 
                           n4665);
   U3298 : NAND2_X1 port map( A1 => n19775, A2 => n11363, ZN => n2102);
   U3301 : NAND3_X1 port map( A1 => n8145, A2 => n12512, A3 => n19775, ZN => 
                           n19656);
   U3302 : OAI21_X1 port map( A1 => n8277, A2 => n8276, B => n19775, ZN => 
                           n19776);
   U3310 : AND2_X2 port map( A1 => n12208, A2 => n1440, Z => n5341);
   U3311 : OAI21_X1 port map( A1 => n6725, A2 => n19033, B => n874, ZN => 
                           n23032);
   U3314 : AND2_X2 port map( A1 => n18686, A2 => n15540, Z => n22217);
   U3317 : INV_X1 port map( I => n12365, ZN => n28334);
   U3318 : CLKBUF_X12 port map( I => n15894, Z => n16337);
   U3325 : INV_X2 port map( I => n8084, ZN => n24845);
   U3327 : NOR2_X1 port map( A1 => n8084, A2 => n16699, ZN => n27590);
   U3329 : NOR2_X1 port map( A1 => n20680, A2 => n28176, ZN => n20667);
   U3330 : NAND2_X1 port map( A1 => n17751, A2 => n12610, ZN => n12930);
   U3331 : OR2_X2 port map( A1 => n22905, A2 => n23415, Z => n3215);
   U3333 : INV_X1 port map( I => n9455, ZN => n8041);
   U3335 : NAND2_X1 port map( A1 => n13422, A2 => n23120, ZN => n20121);
   U3339 : CLKBUF_X12 port map( I => n18041, Z => n26642);
   U3340 : BUF_X4 port map( I => n18041, Z => n26643);
   U3350 : CLKBUF_X12 port map( I => n12413, Z => n22800);
   U3353 : OR2_X2 port map( A1 => n19161, A2 => n24811, Z => n1626);
   U3354 : INV_X1 port map( I => n3297, ZN => n1045);
   U3363 : NAND3_X1 port map( A1 => n955, A2 => n25340, A3 => n20286, ZN => 
                           n25518);
   U3364 : AND2_X2 port map( A1 => n23916, A2 => n20273, Z => n9192);
   U3369 : BUF_X2 port map( I => n23916, Z => n25573);
   U3371 : INV_X1 port map( I => n18244, ZN => n275);
   U3372 : NAND2_X1 port map( A1 => n829, A2 => n13129, ZN => n17635);
   U3374 : INV_X1 port map( I => n13129, ZN => n9304);
   U3375 : CLKBUF_X12 port map( I => n13129, Z => n27177);
   U3388 : INV_X1 port map( I => n1681, ZN => n27173);
   U3396 : INV_X1 port map( I => n1681, ZN => n6058);
   U3397 : NAND2_X1 port map( A1 => n1681, A2 => n14632, ZN => n22170);
   U3398 : NAND3_X1 port map( A1 => n4021, A2 => n20022, A3 => n27846, ZN => 
                           n26007);
   U3403 : OR2_X2 port map( A1 => n4274, A2 => n4021, Z => n4109);
   U3409 : NAND2_X1 port map( A1 => n7496, A2 => n8000, ZN => n7495);
   U3413 : OR2_X2 port map( A1 => n3846, A2 => n8000, Z => n17979);
   U3415 : NAND2_X1 port map( A1 => n3846, A2 => n8000, ZN => n17794);
   U3416 : INV_X1 port map( I => n8000, ZN => n23806);
   U3417 : AND2_X2 port map( A1 => n8000, A2 => n5305, Z => n17793);
   U3418 : CLKBUF_X12 port map( I => n16260, Z => n16264);
   U3419 : AND2_X2 port map( A1 => n16260, A2 => n27877, Z => n14347);
   U3421 : NAND2_X1 port map( A1 => n23645, A2 => n25903, ZN => n24969);
   U3422 : NAND2_X1 port map( A1 => n17694, A2 => n17665, ZN => n17903);
   U3423 : NOR2_X1 port map( A1 => n13112, A2 => n27178, ZN => n14904);
   U3427 : OR3_X2 port map( A1 => n7388, A2 => n11372, A3 => n20168, Z => 
                           n24547);
   U3432 : NAND2_X1 port map( A1 => n14176, A2 => n7388, ZN => n24987);
   U3441 : INV_X1 port map( I => n7388, ZN => n24989);
   U3442 : CLKBUF_X12 port map( I => n7388, Z => n25870);
   U3447 : BUF_X4 port map( I => n6301, Z => n26644);
   U3449 : CLKBUF_X4 port map( I => n6301, Z => n26645);
   U3457 : AOI21_X1 port map( A1 => n24922, A2 => n21711, B => n13718, ZN => 
                           n9930);
   U3458 : INV_X1 port map( I => n13718, ZN => n14283);
   U3463 : NAND2_X1 port map( A1 => n2070, A2 => n25099, ZN => n18910);
   U3466 : CLKBUF_X12 port map( I => n26620, Z => n27881);
   U3474 : OAI22_X1 port map( A1 => n20130, A2 => n20129, B1 => n13429, B2 => 
                           n20316, ZN => n28313);
   U3478 : INV_X1 port map( I => n12644, ZN => n26891);
   U3481 : OAI21_X1 port map( A1 => n23253, A2 => n12644, B => n25141, ZN => 
                           n8775);
   U3482 : NAND2_X1 port map( A1 => n18645, A2 => n27830, ZN => n27829);
   U3485 : CLKBUF_X4 port map( I => n18645, Z => n23966);
   U3487 : CLKBUF_X1 port map( I => n18552, Z => n14140);
   U3489 : NAND2_X1 port map( A1 => n26918, A2 => n8740, ZN => n27672);
   U3491 : NAND2_X1 port map( A1 => n8740, A2 => n27647, ZN => n19043);
   U3496 : NOR2_X1 port map( A1 => n8740, A2 => n27647, ZN => n8814);
   U3500 : NAND2_X1 port map( A1 => n1869, A2 => n18005, ZN => n12899);
   U3501 : NOR3_X1 port map( A1 => n19731, A2 => n19676, A3 => n19730, ZN => 
                           n28180);
   U3502 : NAND2_X1 port map( A1 => n6110, A2 => n10337, ZN => n16658);
   U3503 : NAND2_X1 port map( A1 => n6110, A2 => n13739, ZN => n15298);
   U3504 : NOR3_X1 port map( A1 => n25772, A2 => n28400, A3 => n6110, ZN => 
                           n1748);
   U3506 : NOR2_X1 port map( A1 => n12039, A2 => n3297, ZN => n3087);
   U3507 : NAND2_X1 port map( A1 => n3297, A2 => n1053, ZN => n6685);
   U3513 : AND2_X2 port map( A1 => n14663, A2 => n19968, Z => n13379);
   U3515 : CLKBUF_X12 port map( I => n19968, Z => n24027);
   U3516 : AND2_X2 port map( A1 => n19968, A2 => n3223, Z => n2911);
   U3519 : NAND2_X1 port map( A1 => n19877, A2 => n14307, ZN => n2793);
   U3523 : NOR2_X1 port map( A1 => n19842, A2 => n19877, ZN => n19269);
   U3524 : NAND2_X1 port map( A1 => n3439, A2 => n26898, ZN => n11847);
   U3526 : NOR2_X1 port map( A1 => n3439, A2 => n26898, ZN => n10016);
   U3533 : INV_X1 port map( I => n26898, ZN => n1103);
   U3534 : INV_X1 port map( I => n20538, ZN => n12156);
   U3535 : NAND2_X1 port map( A1 => n11658, A2 => n16534, ZN => n16550);
   U3538 : NAND2_X1 port map( A1 => n22643, A2 => n15040, ZN => n19074);
   U3541 : INV_X1 port map( I => n13235, ZN => n1025);
   U3543 : BUF_X2 port map( I => n13235, Z => n24142);
   U3546 : INV_X2 port map( I => n15514, ZN => n1227);
   U3550 : CLKBUF_X4 port map( I => n15514, Z => n26255);
   U3557 : AND2_X1 port map( A1 => n6021, A2 => n15514, Z => n17449);
   U3558 : OR2_X2 port map( A1 => n7966, A2 => n7965, Z => n2325);
   U3561 : CLKBUF_X4 port map( I => n6216, Z => n6145);
   U3562 : CLKBUF_X12 port map( I => n6959, Z => n24501);
   U3563 : NOR2_X1 port map( A1 => n1998, A2 => n14917, ZN => n23093);
   U3564 : NAND2_X1 port map( A1 => n20323, A2 => n20490, ZN => n14377);
   U3565 : AND2_X2 port map( A1 => n22819, A2 => n23713, Z => n5645);
   U3567 : OR2_X2 port map( A1 => n15717, A2 => n20430, Z => n3799);
   U3568 : BUF_X2 port map( I => n15717, Z => n12503);
   U3569 : INV_X2 port map( I => n15717, ZN => n1580);
   U3574 : INV_X2 port map( I => n11376, ZN => n18828);
   U3575 : NAND2_X1 port map( A1 => n1637, A2 => n3493, ZN => n3193);
   U3577 : AND2_X2 port map( A1 => n14193, A2 => n6259, Z => n14429);
   U3579 : OR2_X2 port map( A1 => n6260, A2 => n6259, Z => n6263);
   U3580 : CLKBUF_X12 port map( I => n15861, Z => n26646);
   U3582 : AOI21_X1 port map( A1 => n17971, A2 => n17887, B => n12815, ZN => 
                           n17888);
   U3586 : AND2_X2 port map( A1 => n17976, A2 => n13819, Z => n17977);
   U3587 : NOR2_X1 port map( A1 => n17976, A2 => n2068, ZN => n5296);
   U3590 : INV_X1 port map( I => n2647, ZN => n28248);
   U3594 : AND2_X2 port map( A1 => n25104, A2 => n2647, Z => n26098);
   U3595 : CLKBUF_X12 port map( I => n2647, Z => n22997);
   U3596 : BUF_X4 port map( I => n24400, Z => n26647);
   U3597 : OAI22_X1 port map( A1 => n19473, A2 => n13463, B1 => n19953, B2 => 
                           n11973, ZN => n19474);
   U3603 : NAND3_X1 port map( A1 => n27786, A2 => n19950, A3 => n11973, ZN => 
                           n3152);
   U3604 : INV_X1 port map( I => n11973, ZN => n1807);
   U3605 : INV_X4 port map( I => n3312, ZN => n818);
   U3610 : OR2_X2 port map( A1 => n15732, A2 => n20286, Z => n20114);
   U3614 : INV_X1 port map( I => n15732, ZN => n6952);
   U3615 : CLKBUF_X12 port map( I => n10220, Z => n17442);
   U3618 : INV_X1 port map( I => n3869, ZN => n7386);
   U3619 : AND2_X1 port map( A1 => n2460, A2 => n829, Z => n17817);
   U3624 : NAND2_X1 port map( A1 => n13129, A2 => n2460, ZN => n17636);
   U3625 : OR2_X1 port map( A1 => n2460, A2 => n7156, Z => n12825);
   U3627 : NAND2_X1 port map( A1 => n19019, A2 => n8683, ZN => n18972);
   U3633 : INV_X2 port map( I => n8683, ZN => n18810);
   U3638 : OR2_X2 port map( A1 => n26638, A2 => n27802, Z => n19833);
   U3639 : NAND2_X1 port map( A1 => n5081, A2 => n11413, ZN => n16733);
   U3642 : NOR2_X1 port map( A1 => n3123, A2 => n11413, ZN => n9517);
   U3645 : INV_X2 port map( I => n11413, ZN => n13481);
   U3646 : INV_X1 port map( I => n10635, ZN => n21041);
   U3647 : NAND2_X1 port map( A1 => n3979, A2 => n12637, ZN => n11605);
   U3649 : NOR2_X1 port map( A1 => n12637, A2 => n26396, ZN => n12679);
   U3652 : OAI21_X1 port map( A1 => n4339, A2 => n14093, B => n3470, ZN => 
                           n28074);
   U3654 : AOI21_X1 port map( A1 => n3470, A2 => n16516, B => n13786, ZN => 
                           n5429);
   U3655 : OR3_X2 port map( A1 => n3470, A2 => n16558, A3 => n1519, Z => n4068)
                           ;
   U3656 : OAI21_X1 port map( A1 => n12679, A2 => n3470, B => n1519, ZN => 
                           n27781);
   U3659 : NAND3_X1 port map( A1 => n16558, A2 => n3470, A3 => n1519, ZN => 
                           n11607);
   U3661 : OAI22_X1 port map( A1 => n7147, A2 => n11147, B1 => n10050, B2 => 
                           n27140, ZN => n5304);
   U3664 : NOR2_X1 port map( A1 => n27376, A2 => n20913, ZN => n20918);
   U3671 : NAND3_X1 port map( A1 => n27876, A2 => n13831, A3 => n13889, ZN => 
                           n26507);
   U3673 : NOR2_X1 port map( A1 => n21451, A2 => n13950, ZN => n27078);
   U3676 : NAND2_X1 port map( A1 => n26827, A2 => n21596, ZN => n27625);
   U3682 : OAI22_X1 port map( A1 => n9424, A2 => n21051, B1 => n9423, B2 => 
                           n21036, ZN => n27193);
   U3695 : NAND2_X1 port map( A1 => n20843, A2 => n28214, ZN => n27750);
   U3696 : NOR3_X1 port map( A1 => n7008, A2 => n3273, A3 => n23154, ZN => 
                           n26789);
   U3698 : OAI21_X1 port map( A1 => n9460, A2 => n188, B => n9943, ZN => n22950
                           );
   U3699 : NAND2_X1 port map( A1 => n27098, A2 => n27097, ZN => n27077);
   U3701 : OAI22_X1 port map( A1 => n4851, A2 => n27853, B1 => n1070, B2 => 
                           n24562, ZN => n27315);
   U3703 : NAND2_X1 port map( A1 => n8137, A2 => n27213, ZN => n26419);
   U3704 : NOR2_X1 port map( A1 => n26682, A2 => n27412, ZN => n14148);
   U3707 : INV_X2 port map( I => n12191, ZN => n21173);
   U3709 : BUF_X1 port map( I => n9894, Z => n24685);
   U3715 : NAND2_X1 port map( A1 => n23274, A2 => n13021, ZN => n7452);
   U3716 : BUF_X2 port map( I => n2800, Z => n2778);
   U3721 : CLKBUF_X4 port map( I => n12011, Z => n7944);
   U3725 : NAND2_X1 port map( A1 => n689, A2 => n15307, ZN => n28470);
   U3727 : AND2_X1 port map( A1 => n26978, A2 => n1083, Z => n20891);
   U3730 : BUF_X2 port map( I => n21501, Z => n23741);
   U3732 : AND2_X1 port map( A1 => n8050, A2 => n21024, Z => n26674);
   U3739 : BUF_X2 port map( I => n26626, Z => n1079);
   U3744 : OR2_X1 port map( A1 => n22421, A2 => n21388, Z => n10197);
   U3745 : BUF_X1 port map( I => n10591, Z => n23999);
   U3753 : BUF_X1 port map( I => n20783, Z => n14647);
   U3756 : CLKBUF_X4 port map( I => n20587, Z => n21714);
   U3761 : OR2_X1 port map( A1 => n15728, A2 => n25388, Z => n21095);
   U3765 : BUF_X1 port map( I => n12315, Z => n26512);
   U3766 : CLKBUF_X4 port map( I => n126, Z => n26651);
   U3769 : INV_X1 port map( I => n2201, ZN => n14882);
   U3771 : BUF_X2 port map( I => n12959, Z => n7248);
   U3776 : CLKBUF_X4 port map( I => n21317, Z => n28502);
   U3778 : CLKBUF_X2 port map( I => n10202, Z => n26848);
   U3783 : INV_X1 port map( I => n27021, ZN => n8731);
   U3784 : NAND2_X1 port map( A1 => n5856, A2 => n6471, ZN => n26837);
   U3788 : INV_X2 port map( I => n7134, ZN => n27630);
   U3792 : INV_X1 port map( I => n20187, ZN => n27214);
   U3800 : OR2_X1 port map( A1 => n14554, A2 => n27091, Z => n8245);
   U3802 : NAND2_X1 port map( A1 => n27602, A2 => n22790, ZN => n12746);
   U3803 : CLKBUF_X2 port map( I => n20196, Z => n27984);
   U3807 : INV_X2 port map( I => n26206, ZN => n19981);
   U3811 : INV_X2 port map( I => n24862, ZN => n25045);
   U3817 : CLKBUF_X2 port map( I => n22374, Z => n27197);
   U3824 : NAND2_X1 port map( A1 => n2173, A2 => n5785, ZN => n5784);
   U3830 : NAND2_X1 port map( A1 => n26804, A2 => n1937, ZN => n25405);
   U3834 : INV_X1 port map( I => n22148, ZN => n27236);
   U3841 : INV_X1 port map( I => n19920, ZN => n19868);
   U3845 : OAI21_X1 port map( A1 => n14043, A2 => n14042, B => n19941, ZN => 
                           n26963);
   U3846 : INV_X1 port map( I => n27059, ZN => n23196);
   U3847 : NAND2_X1 port map( A1 => n27305, A2 => n27304, ZN => n27303);
   U3855 : INV_X1 port map( I => n28485, ZN => n28484);
   U3858 : INV_X1 port map( I => n27001, ZN => n19712);
   U3859 : INV_X1 port map( I => n24337, ZN => n15321);
   U3862 : NAND2_X1 port map( A1 => n27154, A2 => n27152, ZN => n19688);
   U3863 : INV_X1 port map( I => n27153, ZN => n27152);
   U3867 : BUF_X1 port map( I => n14531, Z => n28425);
   U3868 : INV_X1 port map( I => n26803, ZN => n27025);
   U3869 : BUF_X1 port map( I => n19759, Z => n14672);
   U3870 : INV_X1 port map( I => n28298, ZN => n28297);
   U3878 : INV_X2 port map( I => n14568, ZN => n26653);
   U3884 : AND2_X1 port map( A1 => n6861, A2 => n13167, Z => n6392);
   U3885 : BUF_X2 port map( I => n19923, Z => n24187);
   U3886 : NAND2_X1 port map( A1 => n26296, A2 => n27608, ZN => n10045);
   U3888 : CLKBUF_X2 port map( I => n23278, Z => n26948);
   U3893 : CLKBUF_X2 port map( I => n24317, Z => n26767);
   U3894 : INV_X1 port map( I => n19905, ZN => n27802);
   U3895 : CLKBUF_X2 port map( I => n7340, Z => n3226);
   U3898 : CLKBUF_X1 port map( I => n26297, Z => n27608);
   U3908 : BUF_X2 port map( I => n19792, Z => n23322);
   U3909 : BUF_X4 port map( I => n19679, Z => n26654);
   U3912 : NAND2_X1 port map( A1 => n6740, A2 => n1135, ZN => n26811);
   U3914 : NAND2_X1 port map( A1 => n27114, A2 => n27113, ZN => n7523);
   U3916 : INV_X1 port map( I => n19237, ZN => n28514);
   U3923 : INV_X1 port map( I => n12697, ZN => n9544);
   U3924 : NAND2_X1 port map( A1 => n27562, A2 => n10316, ZN => n28124);
   U3928 : OR2_X1 port map( A1 => n5138, A2 => n2798, Z => n24449);
   U3934 : CLKBUF_X4 port map( I => n18959, Z => n28240);
   U3939 : NAND2_X1 port map( A1 => n28170, A2 => n15294, ZN => n18656);
   U3940 : INV_X1 port map( I => n1154, ZN => n27536);
   U3941 : NAND2_X1 port map( A1 => n4453, A2 => n998, ZN => n27231);
   U3942 : INV_X1 port map( I => n6489, ZN => n19028);
   U3947 : NOR2_X1 port map( A1 => n4624, A2 => n24937, ZN => n1604);
   U3950 : INV_X1 port map( I => n10128, ZN => n27626);
   U3951 : INV_X1 port map( I => n18926, ZN => n22472);
   U3958 : NAND2_X1 port map( A1 => n19132, A2 => n25327, ZN => n27553);
   U3969 : BUF_X2 port map( I => n19107, Z => n9268);
   U3970 : BUF_X2 port map( I => n19116, Z => n7970);
   U3972 : CLKBUF_X2 port map( I => n13349, Z => n23931);
   U3975 : CLKBUF_X2 port map( I => n19126, Z => n26762);
   U3976 : CLKBUF_X2 port map( I => n988, Z => n27868);
   U3977 : CLKBUF_X2 port map( I => n28237, Z => n27258);
   U3980 : BUF_X2 port map( I => n19052, Z => n28372);
   U3982 : CLKBUF_X2 port map( I => n2582, Z => n26831);
   U3983 : BUF_X2 port map( I => n1772, Z => n28311);
   U3985 : CLKBUF_X4 port map( I => n25412, Z => n28499);
   U3987 : CLKBUF_X2 port map( I => n19163, Z => n27279);
   U3990 : INV_X2 port map( I => n2582, ZN => n19057);
   U3996 : CLKBUF_X4 port map( I => n8049, Z => n4471);
   U3997 : CLKBUF_X2 port map( I => n22626, Z => n28507);
   U3999 : BUF_X2 port map( I => n19088, Z => n14358);
   U4000 : NAND2_X1 port map( A1 => n6689, A2 => n4348, ZN => n1377);
   U4001 : NAND2_X1 port map( A1 => n6913, A2 => n1800, ZN => n5991);
   U4003 : INV_X1 port map( I => n28346, ZN => n28345);
   U4005 : NAND2_X1 port map( A1 => n27713, A2 => n27712, ZN => n9588);
   U4012 : INV_X1 port map( I => n27664, ZN => n9713);
   U4020 : OAI21_X1 port map( A1 => n10660, A2 => n13360, B => n759, ZN => 
                           n18449);
   U4023 : INV_X1 port map( I => n27150, ZN => n3889);
   U4024 : AND2_X1 port map( A1 => n14022, A2 => n18763, Z => n26697);
   U4025 : OR2_X1 port map( A1 => n14140, A2 => n15660, Z => n26699);
   U4031 : NAND2_X1 port map( A1 => n26745, A2 => n26744, ZN => n2950);
   U4033 : NAND2_X1 port map( A1 => n10537, A2 => n759, ZN => n26541);
   U4034 : NAND2_X1 port map( A1 => n18419, A2 => n23399, ZN => n7100);
   U4035 : CLKBUF_X2 port map( I => n18741, Z => n26894);
   U4036 : CLKBUF_X2 port map( I => n3903, Z => n27739);
   U4038 : CLKBUF_X4 port map( I => n18674, Z => n27281);
   U4039 : BUF_X1 port map( I => n23841, Z => n14498);
   U4041 : INV_X2 port map( I => n18452, ZN => n13963);
   U4042 : INV_X1 port map( I => n27436, ZN => n18294);
   U4044 : BUF_X2 port map( I => n10561, Z => n7791);
   U4046 : INV_X1 port map( I => n3153, ZN => n28073);
   U4047 : CLKBUF_X2 port map( I => n1970, Z => n28315);
   U4050 : NOR2_X1 port map( A1 => n27157, A2 => n3269, ZN => n5764);
   U4064 : NAND2_X1 port map( A1 => n17703, A2 => n17704, ZN => n15430);
   U4068 : INV_X1 port map( I => n24902, ZN => n28038);
   U4069 : AND3_X1 port map( A1 => n4812, A2 => n17926, A3 => n17924, Z => 
                           n26716);
   U4073 : NAND2_X1 port map( A1 => n12001, A2 => n8365, ZN => n28335);
   U4076 : INV_X2 port map( I => n17912, ZN => n1200);
   U4077 : INV_X1 port map( I => n27068, ZN => n27521);
   U4078 : NAND2_X1 port map( A1 => n7986, A2 => n8070, ZN => n24933);
   U4079 : NAND3_X1 port map( A1 => n28239, A2 => n25738, A3 => n8882, ZN => 
                           n27342);
   U4080 : INV_X1 port map( I => n1210, ZN => n28327);
   U4081 : INV_X1 port map( I => n18004, ZN => n27186);
   U4091 : NOR2_X1 port map( A1 => n28057, A2 => n28056, ZN => n9636);
   U4097 : BUF_X2 port map( I => n22834, Z => n27820);
   U4100 : INV_X1 port map( I => n23072, ZN => n28004);
   U4101 : BUF_X1 port map( I => n24304, Z => n28239);
   U4102 : NAND2_X1 port map( A1 => n27619, A2 => n5166, ZN => n5165);
   U4103 : NAND2_X1 port map( A1 => n13767, A2 => n26614, ZN => n17357);
   U4107 : INV_X1 port map( I => n26217, ZN => n26873);
   U4109 : NOR2_X1 port map( A1 => n5579, A2 => n4267, ZN => n26872);
   U4111 : INV_X1 port map( I => n17208, ZN => n17209);
   U4112 : AND2_X1 port map( A1 => n14061, A2 => n17560, Z => n26666);
   U4114 : OAI21_X1 port map( A1 => n26532, A2 => n17323, B => n17322, ZN => 
                           n21952);
   U4115 : INV_X1 port map( I => n17533, ZN => n26332);
   U4118 : INV_X1 port map( I => n15055, ZN => n28535);
   U4119 : CLKBUF_X2 port map( I => n9481, Z => n27580);
   U4125 : OAI21_X1 port map( A1 => n7245, A2 => n26923, B => n1040, ZN => 
                           n28349);
   U4128 : INV_X1 port map( I => n27181, ZN => n27180);
   U4133 : BUF_X1 port map( I => n540, Z => n14532);
   U4135 : BUF_X1 port map( I => n17548, Z => n26363);
   U4139 : INV_X4 port map( I => n17489, ZN => n26655);
   U4140 : CLKBUF_X2 port map( I => n17413, Z => n27132);
   U4150 : AND2_X1 port map( A1 => n26081, A2 => n17513, Z => n10585);
   U4157 : CLKBUF_X2 port map( I => n24585, Z => n28501);
   U4158 : BUF_X2 port map( I => n17412, Z => n14250);
   U4160 : CLKBUF_X2 port map( I => n17469, Z => n28025);
   U4161 : CLKBUF_X2 port map( I => n12040, Z => n27288);
   U4165 : BUF_X2 port map( I => n17343, Z => n24214);
   U4166 : CLKBUF_X2 port map( I => n23352, Z => n27705);
   U4171 : NAND2_X1 port map( A1 => n11606, A2 => n11607, ZN => n1374);
   U4172 : CLKBUF_X2 port map( I => n16858, Z => n27104);
   U4173 : AOI21_X1 port map( A1 => n10988, A2 => n24351, B => n27934, ZN => 
                           n27933);
   U4175 : NAND2_X1 port map( A1 => n27328, A2 => n26169, ZN => n1579);
   U4181 : NAND2_X1 port map( A1 => n9392, A2 => n23261, ZN => n26976);
   U4184 : NAND2_X1 port map( A1 => n9819, A2 => n9820, ZN => n28434);
   U4185 : INV_X1 port map( I => n27653, ZN => n16519);
   U4186 : NAND2_X1 port map( A1 => n23162, A2 => n16435, ZN => n16398);
   U4191 : BUF_X2 port map( I => n25875, Z => n27160);
   U4196 : CLKBUF_X2 port map( I => n28113, Z => n27019);
   U4198 : BUF_X1 port map( I => n16730, Z => n26993);
   U4202 : CLKBUF_X2 port map( I => n16526, Z => n26760);
   U4203 : CLKBUF_X2 port map( I => n10337, Z => n27543);
   U4205 : INV_X2 port map( I => n26578, ZN => n16561);
   U4206 : BUF_X2 port map( I => n16712, Z => n10304);
   U4210 : BUF_X2 port map( I => n11962, Z => n6683);
   U4214 : NOR2_X1 port map( A1 => n15940, A2 => n7152, ZN => n27902);
   U4215 : CLKBUF_X2 port map( I => n15885, Z => n6480);
   U4221 : NAND2_X1 port map( A1 => n14695, A2 => n16335, ZN => n5928);
   U4234 : OR2_X1 port map( A1 => n15936, A2 => n8031, Z => n16304);
   U4236 : INV_X2 port map( I => n9986, ZN => n16229);
   U4239 : CLKBUF_X4 port map( I => n15929, Z => n16140);
   U4241 : CLKBUF_X2 port map( I => n16141, Z => n25873);
   U4243 : CLKBUF_X2 port map( I => n13418, Z => n27878);
   U4245 : CLKBUF_X2 port map( I => n16093, Z => n16072);
   U4246 : INV_X1 port map( I => n14588, ZN => n28342);
   U4249 : BUF_X2 port map( I => n16187, Z => n16188);
   U4251 : CLKBUF_X2 port map( I => Key(114), Z => n20919);
   U4252 : BUF_X2 port map( I => Key(53), Z => n20961);
   U4257 : NOR2_X1 port map( A1 => n12116, A2 => n263, ZN => n23948);
   U4263 : NAND2_X1 port map( A1 => n11, A2 => n24132, ZN => n16218);
   U4266 : NAND2_X1 port map( A1 => n16280, A2 => n12507, ZN => n11293);
   U4268 : CLKBUF_X2 port map( I => n22623, Z => n25222);
   U4269 : OAI21_X1 port map( A1 => n15998, A2 => n14584, B => n263, ZN => 
                           n26018);
   U4270 : NAND2_X1 port map( A1 => n16337, A2 => n9308, ZN => n15895);
   U4271 : AOI21_X1 port map( A1 => n16269, A2 => n15491, B => n5853, ZN => 
                           n10093);
   U4276 : NAND2_X1 port map( A1 => n15936, A2 => n16330, ZN => n16034);
   U4287 : CLKBUF_X2 port map( I => n16227, Z => n28088);
   U4294 : NAND2_X1 port map( A1 => n16264, A2 => n15607, ZN => n16261);
   U4296 : NOR2_X1 port map( A1 => n8873, A2 => n16273, ZN => n16109);
   U4301 : NAND2_X1 port map( A1 => n15986, A2 => n16144, ZN => n24268);
   U4304 : NAND2_X1 port map( A1 => n16304, A2 => n16330, ZN => n15018);
   U4306 : CLKBUF_X2 port map( I => n11407, Z => n26879);
   U4307 : INV_X1 port map( I => n16118, ZN => n15977);
   U4312 : NAND2_X1 port map( A1 => n13457, A2 => n27878, ZN => n10186);
   U4314 : INV_X2 port map( I => n15282, ZN => n16333);
   U4315 : NAND2_X1 port map( A1 => n26018, A2 => n26017, ZN => n25942);
   U4316 : NAND2_X1 port map( A1 => n16140, A2 => n15686, ZN => n7015);
   U4317 : NAND2_X1 port map( A1 => n15760, A2 => n16077, ZN => n16217);
   U4320 : OR2_X1 port map( A1 => n3572, A2 => n23309, Z => n16291);
   U4322 : INV_X1 port map( I => n914, ZN => n27080);
   U4323 : NAND2_X1 port map( A1 => n5637, A2 => n3735, ZN => n25072);
   U4331 : NAND2_X1 port map( A1 => n3771, A2 => n16305, ZN => n13915);
   U4332 : INV_X2 port map( I => n16005, ZN => n1258);
   U4334 : AOI21_X1 port map( A1 => n16265, A2 => n21904, B => n16264, ZN => 
                           n27743);
   U4337 : INV_X1 port map( I => n27669, ZN => n15211);
   U4343 : OAI22_X1 port map( A1 => n3249, A2 => n13677, B1 => n15935, B2 => 
                           n4926, ZN => n3423);
   U4347 : CLKBUF_X2 port map( I => n12529, Z => n7374);
   U4355 : NAND2_X1 port map( A1 => n16215, A2 => n840, ZN => n23166);
   U4357 : NAND2_X1 port map( A1 => n28033, A2 => n28032, ZN => n3573);
   U4360 : INV_X1 port map( I => n15986, ZN => n16020);
   U4363 : NOR2_X1 port map( A1 => n24198, A2 => n5681, ZN => n1842);
   U4364 : INV_X1 port map( I => n3443, ZN => n27572);
   U4366 : INV_X2 port map( I => n1519, ZN => n13786);
   U4369 : INV_X1 port map( I => n16565, ZN => n16518);
   U4371 : NAND2_X1 port map( A1 => n16481, A2 => n1241, ZN => n1562);
   U4373 : NOR2_X1 port map( A1 => n794, A2 => n16730, ZN => n9799);
   U4375 : NOR2_X1 port map( A1 => n1047, A2 => n24215, ZN => n8363);
   U4389 : NOR2_X1 port map( A1 => n10393, A2 => n9314, ZN => n16490);
   U4391 : NOR2_X1 port map( A1 => n14656, A2 => n23907, ZN => n1697);
   U4395 : NOR2_X1 port map( A1 => n8799, A2 => n8797, ZN => n8796);
   U4396 : NOR2_X1 port map( A1 => n390, A2 => n26175, ZN => n26174);
   U4400 : NAND2_X1 port map( A1 => n24028, A2 => n25130, ZN => n10517);
   U4401 : CLKBUF_X4 port map( I => n12884, Z => n4162);
   U4404 : NOR2_X1 port map( A1 => n23749, A2 => n13721, ZN => n22110);
   U4406 : NAND2_X1 port map( A1 => n458, A2 => n27896, ZN => n22299);
   U4413 : OAI21_X1 port map( A1 => n16057, A2 => n10567, B => n404, ZN => 
                           n7241);
   U4419 : AOI21_X1 port map( A1 => n5124, A2 => n24646, B => n173, ZN => 
                           n27728);
   U4431 : NAND3_X1 port map( A1 => n5874, A2 => n16224, A3 => n28113, ZN => 
                           n28475);
   U4434 : OAI21_X1 port map( A1 => n12525, A2 => n12526, B => n6937, ZN => 
                           n23379);
   U4435 : NAND2_X1 port map( A1 => n3948, A2 => n5266, ZN => n10260);
   U4438 : INV_X1 port map( I => n16944, ZN => n17138);
   U4439 : INV_X1 port map( I => n17124, ZN => n2376);
   U4441 : NAND2_X1 port map( A1 => n16692, A2 => n5558, ZN => n6395);
   U4445 : INV_X1 port map( I => n27933, ZN => n17016);
   U4446 : INV_X1 port map( I => n16930, ZN => n26289);
   U4447 : OAI21_X1 port map( A1 => n21809, A2 => n16438, B => n16496, ZN => 
                           n4217);
   U4453 : BUF_X2 port map( I => n12275, Z => n27936);
   U4455 : INV_X1 port map( I => n5624, ZN => n10669);
   U4456 : CLKBUF_X2 port map( I => n16980, Z => n6765);
   U4473 : CLKBUF_X1 port map( I => n17055, Z => n14335);
   U4476 : INV_X1 port map( I => n10516, ZN => n17087);
   U4481 : INV_X1 port map( I => n14016, ZN => n27955);
   U4485 : INV_X1 port map( I => n17102, ZN => n27136);
   U4487 : INV_X1 port map( I => n11780, ZN => n25683);
   U4489 : INV_X1 port map( I => n7701, ZN => n27741);
   U4494 : INV_X2 port map( I => n24070, ZN => n13380);
   U4496 : NAND2_X1 port map( A1 => n1435, A2 => n17518, ZN => n17516);
   U4497 : NAND2_X1 port map( A1 => n5489, A2 => n24018, ZN => n11944);
   U4502 : NOR2_X1 port map( A1 => n17502, A2 => n242, ZN => n6551);
   U4507 : NAND2_X1 port map( A1 => n10985, A2 => n17452, ZN => n16970);
   U4514 : CLKBUF_X2 port map( I => n17419, Z => n17196);
   U4523 : NAND2_X1 port map( A1 => n16996, A2 => n9481, ZN => n231);
   U4528 : CLKBUF_X2 port map( I => n17422, Z => n14324);
   U4529 : NOR2_X1 port map( A1 => n3700, A2 => n13358, ZN => n23170);
   U4530 : NOR2_X1 port map( A1 => n461, A2 => n17454, ZN => n28271);
   U4535 : CLKBUF_X4 port map( I => n24649, Z => n24560);
   U4541 : NAND2_X1 port map( A1 => n23571, A2 => n10015, ZN => n27983);
   U4543 : NAND3_X1 port map( A1 => n5639, A2 => n17513, A3 => n26628, ZN => 
                           n23025);
   U4546 : INV_X1 port map( I => n17543, ZN => n17443);
   U4548 : CLKBUF_X1 port map( I => n17244, Z => n23421);
   U4553 : NAND2_X1 port map( A1 => n17502, A2 => n1228, ZN => n13319);
   U4554 : CLKBUF_X2 port map( I => n17324, Z => n26532);
   U4561 : INV_X2 port map( I => n3533, ZN => n12236);
   U4562 : OAI22_X1 port map( A1 => n17366, A2 => n9593, B1 => n27351, B2 => 
                           n14061, ZN => n17367);
   U4565 : CLKBUF_X1 port map( I => n10183, Z => n26782);
   U4566 : AOI21_X1 port map( A1 => n17372, A2 => n10150, B => n401, ZN => 
                           n9610);
   U4567 : AOI22_X1 port map( A1 => n26655, A2 => n26351, B1 => n14504, B2 => 
                           n25922, ZN => n27960);
   U4570 : NOR2_X1 port map( A1 => n508, A2 => n17471, ZN => n8660);
   U4582 : OR2_X1 port map( A1 => n7651, A2 => n5605, Z => n17295);
   U4583 : INV_X2 port map( I => n14944, ZN => n9827);
   U4586 : OAI21_X1 port map( A1 => n22578, A2 => n17427, B => n17521, ZN => 
                           n12551);
   U4590 : NAND2_X1 port map( A1 => n7151, A2 => n1039, ZN => n7456);
   U4601 : NOR3_X1 port map( A1 => n24406, A2 => n10546, A3 => n21785, ZN => 
                           n16872);
   U4612 : CLKBUF_X2 port map( I => n9070, Z => n25504);
   U4615 : CLKBUF_X2 port map( I => n17137, Z => n17472);
   U4619 : AOI21_X1 port map( A1 => n9767, A2 => n17735, B => n9766, ZN => 
                           n17566);
   U4625 : OAI21_X1 port map( A1 => n6663, A2 => n14504, B => n830, ZN => 
                           n26448);
   U4626 : AOI22_X1 port map( A1 => n17255, A2 => n15189, B1 => n17363, B2 => 
                           n13268, ZN => n27189);
   U4628 : NAND2_X1 port map( A1 => n4486, A2 => n1219, ZN => n7990);
   U4632 : INV_X1 port map( I => n24304, ZN => n2051);
   U4634 : CLKBUF_X2 port map( I => n17917, Z => n24564);
   U4636 : OAI21_X1 port map( A1 => n25013, A2 => n8237, B => n2502, ZN => 
                           n8251);
   U4645 : NAND2_X1 port map( A1 => n787, A2 => n17761, ZN => n5826);
   U4646 : NAND2_X1 port map( A1 => n6709, A2 => n6098, ZN => n17597);
   U4650 : INV_X1 port map( I => n12825, ZN => n10178);
   U4652 : AOI21_X1 port map( A1 => n13061, A2 => n4318, B => n21943, ZN => 
                           n11653);
   U4655 : NAND3_X1 port map( A1 => n15462, A2 => n27699, A3 => n17678, ZN => 
                           n4916);
   U4662 : NAND2_X1 port map( A1 => n27342, A2 => n17794, ZN => n27157);
   U4666 : INV_X1 port map( I => n28302, ZN => n1028);
   U4668 : INV_X1 port map( I => n17818, ZN => n17929);
   U4670 : INV_X2 port map( I => n22519, ZN => n7614);
   U4677 : NAND3_X1 port map( A1 => n14578, A2 => n27161, A3 => n9879, ZN => 
                           n9684);
   U4679 : INV_X1 port map( I => n14278, ZN => n17872);
   U4680 : AOI21_X1 port map( A1 => n28322, A2 => n14284, B => n28194, ZN => 
                           n3041);
   U4683 : NAND2_X1 port map( A1 => n8365, A2 => n12899, ZN => n23031);
   U4686 : NOR2_X1 port map( A1 => n6179, A2 => n17725, ZN => n27772);
   U4689 : NAND3_X1 port map( A1 => n28401, A2 => n11967, A3 => n13329, ZN => 
                           n27339);
   U4693 : NOR2_X1 port map( A1 => n6799, A2 => n789, ZN => n23087);
   U4695 : NAND3_X1 port map( A1 => n17742, A2 => n17925, A3 => n26533, ZN => 
                           n17258);
   U4697 : NAND2_X1 port map( A1 => n23441, A2 => n17903, ZN => n24816);
   U4701 : NAND3_X1 port map( A1 => n12825, A2 => n17636, A3 => n21779, ZN => 
                           n12335);
   U4702 : NAND2_X1 port map( A1 => n12731, A2 => n26194, ZN => n17854);
   U4704 : INV_X1 port map( I => n11858, ZN => n1437);
   U4707 : CLKBUF_X2 port map( I => n14278, Z => n23115);
   U4710 : NAND2_X1 port map( A1 => n24350, A2 => n10895, ZN => n27254);
   U4712 : CLKBUF_X2 port map( I => n25105, Z => n24848);
   U4714 : INV_X1 port map( I => n18267, ZN => n26003);
   U4717 : OAI21_X1 port map( A1 => n2436, A2 => n14980, B => n2433, ZN => 
                           n18082);
   U4718 : INV_X1 port map( I => n25068, ZN => n18348);
   U4725 : NAND2_X1 port map( A1 => n4198, A2 => n10206, ZN => n6426);
   U4727 : NAND2_X1 port map( A1 => n13538, A2 => n22825, ZN => n3984);
   U4739 : INV_X1 port map( I => n18137, ZN => n15719);
   U4741 : INV_X1 port map( I => n18087, ZN => n9914);
   U4750 : NAND2_X1 port map( A1 => n5554, A2 => n348, ZN => n18447);
   U4752 : NOR2_X1 port map( A1 => n14594, A2 => n22799, ZN => n22680);
   U4753 : CLKBUF_X1 port map( I => n18740, Z => n27737);
   U4758 : INV_X1 port map( I => n10555, ZN => n22681);
   U4761 : INV_X2 port map( I => n24032, ZN => n14022);
   U4765 : NOR2_X1 port map( A1 => n10642, A2 => n18785, ZN => n28459);
   U4766 : CLKBUF_X2 port map( I => n18609, Z => n18696);
   U4769 : INV_X1 port map( I => n10708, ZN => n6173);
   U4773 : INV_X2 port map( I => n1015, ZN => n878);
   U4777 : NAND2_X1 port map( A1 => n3062, A2 => n22856, ZN => n18756);
   U4780 : NAND2_X1 port map( A1 => n18445, A2 => n28543, ZN => n18533);
   U4782 : INV_X1 port map( I => n1974, ZN => n11994);
   U4786 : NOR2_X1 port map( A1 => n18778, A2 => n18505, ZN => n14819);
   U4787 : NOR2_X1 port map( A1 => n15448, A2 => n18487, ZN => n8792);
   U4788 : INV_X1 port map( I => n18532, ZN => n27713);
   U4789 : INV_X2 port map( I => n24523, ZN => n18537);
   U4792 : INV_X1 port map( I => n357, ZN => n24047);
   U4795 : INV_X1 port map( I => n7350, ZN => n10322);
   U4798 : NOR2_X1 port map( A1 => n8651, A2 => n18256, ZN => n18391);
   U4800 : NAND2_X1 port map( A1 => n27747, A2 => n1012, ZN => n27746);
   U4801 : OAI22_X1 port map( A1 => n21783, A2 => n2072, B1 => n18784, B2 => 
                           n24243, ZN => n18651);
   U4803 : NOR2_X1 port map( A1 => n23060, A2 => n18947, ZN => n18863);
   U4804 : CLKBUF_X2 port map( I => n18457, Z => n14408);
   U4805 : NAND2_X1 port map( A1 => n24801, A2 => n27175, ZN => n18523);
   U4817 : NAND2_X1 port map( A1 => n18470, A2 => n18697, ZN => n22127);
   U4819 : NAND2_X1 port map( A1 => n19114, A2 => n18999, ZN => n3851);
   U4820 : AOI21_X1 port map( A1 => n1722, A2 => n18516, B => n1191, ZN => 
                           n23479);
   U4822 : OAI21_X1 port map( A1 => n11299, A2 => n21790, B => n27830, ZN => 
                           n13289);
   U4827 : NOR2_X1 port map( A1 => n25586, A2 => n19164, ZN => n18894);
   U4830 : CLKBUF_X1 port map( I => n25514, Z => n26997);
   U4831 : NOR2_X1 port map( A1 => n28303, A2 => n19152, ZN => n14892);
   U4832 : NAND2_X1 port map( A1 => n13573, A2 => n12111, ZN => n12234);
   U4844 : NOR2_X1 port map( A1 => n2726, A2 => n2820, ZN => n19040);
   U4845 : INV_X2 port map( I => n6447, ZN => n9376);
   U4847 : INV_X1 port map( I => n25914, ZN => n23618);
   U4857 : NAND2_X1 port map( A1 => n13015, A2 => n26720, ZN => n22648);
   U4858 : INV_X2 port map( I => n6889, ZN => n23844);
   U4859 : INV_X1 port map( I => n7840, ZN => n10239);
   U4861 : CLKBUF_X2 port map( I => n20, Z => n26234);
   U4863 : INV_X2 port map( I => n18426, ZN => n1165);
   U4865 : NOR3_X1 port map( A1 => n23559, A2 => n18894, A3 => n22338, ZN => 
                           n2108);
   U4866 : OAI21_X1 port map( A1 => n19112, A2 => n19113, B => n25770, ZN => 
                           n10977);
   U4867 : NAND2_X1 port map( A1 => n997, A2 => n7970, ZN => n19001);
   U4868 : NAND2_X1 port map( A1 => n19017, A2 => n24170, ZN => n18254);
   U4869 : NAND2_X1 port map( A1 => n18926, A2 => n18924, ZN => n18393);
   U4870 : OAI21_X1 port map( A1 => n7445, A2 => n14119, B => n9922, ZN => 
                           n6133);
   U4874 : NAND2_X1 port map( A1 => n19102, A2 => n19101, ZN => n9657);
   U4877 : NAND2_X1 port map( A1 => n9407, A2 => n25864, ZN => n6418);
   U4879 : CLKBUF_X4 port map( I => n19056, Z => n23305);
   U4882 : CLKBUF_X4 port map( I => n14836, Z => n2356);
   U4884 : INV_X1 port map( I => n19146, ZN => n28128);
   U4886 : NAND2_X1 port map( A1 => n13270, A2 => n25592, ZN => n14289);
   U4888 : NOR2_X1 port map( A1 => n19192, A2 => n12772, ZN => n12771);
   U4891 : INV_X2 port map( I => n4147, ZN => n19406);
   U4896 : NAND2_X1 port map( A1 => n19375, A2 => n4441, ZN => n4443);
   U4898 : CLKBUF_X4 port map( I => n11575, Z => n24384);
   U4902 : INV_X1 port map( I => n19449, ZN => n23636);
   U4906 : INV_X1 port map( I => n19460, ZN => n24242);
   U4908 : INV_X1 port map( I => n13157, ZN => n5852);
   U4911 : NAND2_X1 port map( A1 => n26654, A2 => n19586, ZN => n15286);
   U4912 : INV_X2 port map( I => n7682, ZN => n11079);
   U4914 : INV_X1 port map( I => n26447, ZN => n27304);
   U4915 : CLKBUF_X2 port map( I => n19693, Z => n6987);
   U4920 : INV_X1 port map( I => n11619, ZN => n19822);
   U4923 : INV_X1 port map( I => n19952, ZN => n13463);
   U4929 : NAND2_X1 port map( A1 => n756, A2 => n815, ZN => n19837);
   U4932 : OAI21_X1 port map( A1 => n22775, A2 => n28168, B => n28225, ZN => 
                           n22148);
   U4933 : INV_X2 port map( I => n10601, ZN => n863);
   U4934 : NAND2_X1 port map( A1 => n19758, A2 => n4432, ZN => n4439);
   U4935 : NAND2_X1 port map( A1 => n10549, A2 => n26623, ZN => n19895);
   U4942 : NOR2_X1 port map( A1 => n9762, A2 => n10041, ZN => n24950);
   U4946 : NAND2_X1 port map( A1 => n19819, A2 => n10601, ZN => n27001);
   U4947 : NOR2_X1 port map( A1 => n9994, A2 => n19822, ZN => n23034);
   U4951 : INV_X1 port map( I => n25899, ZN => n19926);
   U4952 : NOR2_X1 port map( A1 => n19711, A2 => n10498, ZN => n23000);
   U4956 : NOR2_X1 port map( A1 => n19953, A2 => n19952, ZN => n13246);
   U4961 : CLKBUF_X2 port map( I => n7463, Z => n4432);
   U4962 : INV_X1 port map( I => n13665, ZN => n19743);
   U4971 : NOR2_X1 port map( A1 => n864, A2 => n19743, ZN => n19746);
   U4974 : NAND2_X1 port map( A1 => n810, A2 => n19890, ZN => n27913);
   U4975 : NOR2_X1 port map( A1 => n510, A2 => n14193, ZN => n14192);
   U4976 : INV_X1 port map( I => n15457, ZN => n5332);
   U4977 : OAI21_X1 port map( A1 => n21945, A2 => n1655, B => n27001, ZN => 
                           n27000);
   U4978 : NAND2_X1 port map( A1 => n20280, A2 => n14663, ZN => n27276);
   U4989 : INV_X2 port map( I => n19846, ZN => n19847);
   U4992 : INV_X1 port map( I => n27435, ZN => n27195);
   U4997 : INV_X1 port map( I => n19761, ZN => n4775);
   U4999 : NAND2_X1 port map( A1 => n22214, A2 => n22213, ZN => n8299);
   U5001 : INV_X1 port map( I => n19697, ZN => n7129);
   U5006 : OAI21_X1 port map( A1 => n12617, A2 => n19937, B => n7176, ZN => 
                           n19938);
   U5011 : NOR2_X1 port map( A1 => n19936, A2 => n10601, ZN => n9628);
   U5012 : INV_X2 port map( I => n19819, ZN => n9561);
   U5015 : NAND3_X1 port map( A1 => n21782, A2 => n4565, A3 => n815, ZN => 
                           n8563);
   U5016 : AOI21_X1 port map( A1 => n26986, A2 => n26985, B => n8952, ZN => 
                           n27005);
   U5026 : NOR2_X1 port map( A1 => n2891, A2 => n12395, ZN => n24855);
   U5031 : NAND2_X1 port map( A1 => n9583, A2 => n9584, ZN => n1937);
   U5034 : AOI22_X1 port map( A1 => n6142, A2 => n13110, B1 => n976, B2 => 
                           n6143, ZN => n6141);
   U5035 : NAND2_X1 port map( A1 => n7068, A2 => n7069, ZN => n3927);
   U5039 : NAND2_X1 port map( A1 => n15321, A2 => n27856, ZN => n28029);
   U5055 : NOR2_X1 port map( A1 => n11052, A2 => n27195, ZN => n27194);
   U5057 : INV_X1 port map( I => n5934, ZN => n13614);
   U5059 : NOR3_X1 port map( A1 => n25340, A2 => n23906, A3 => n23229, ZN => 
                           n24037);
   U5060 : OAI21_X1 port map( A1 => n4563, A2 => n4564, B => n2231, ZN => n6313
                           );
   U5064 : INV_X2 port map( I => n20072, ZN => n855);
   U5071 : BUF_X2 port map( I => n13853, Z => n28519);
   U5073 : NAND2_X1 port map( A1 => n27434, A2 => n28326, ZN => n27951);
   U5074 : CLKBUF_X2 port map( I => n2890, Z => n22342);
   U5075 : CLKBUF_X4 port map( I => n20189, Z => n1835);
   U5081 : NAND2_X1 port map( A1 => n20107, A2 => n8135, ZN => n1932);
   U5085 : NAND2_X1 port map( A1 => n8099, A2 => n8098, ZN => n22745);
   U5089 : NAND2_X1 port map( A1 => n20085, A2 => n20084, ZN => n1478);
   U5091 : NAND2_X1 port map( A1 => n190, A2 => n11151, ZN => n26137);
   U5094 : INV_X2 port map( I => n11756, ZN => n20125);
   U5098 : NAND2_X1 port map( A1 => n4912, A2 => n4911, ZN => n14868);
   U5099 : INV_X1 port map( I => n2655, ZN => n22129);
   U5102 : NAND3_X1 port map( A1 => n2967, A2 => n1447, A3 => n24677, ZN => 
                           n28405);
   U5107 : NAND2_X1 port map( A1 => n20206, A2 => n20108, ZN => n11211);
   U5111 : NAND2_X1 port map( A1 => n28524, A2 => n20045, ZN => n27649);
   U5112 : INV_X1 port map( I => n5102, ZN => n8072);
   U5113 : INV_X1 port map( I => n21185, ZN => n14077);
   U5119 : CLKBUF_X2 port map( I => n20482, Z => n26884);
   U5127 : INV_X1 port map( I => n20446, ZN => n6105);
   U5131 : NAND2_X1 port map( A1 => n13291, A2 => n21618, ZN => n28131);
   U5132 : NAND2_X1 port map( A1 => n20921, A2 => n21924, ZN => n26211);
   U5135 : NOR2_X1 port map( A1 => n20932, A2 => n950, ZN => n5726);
   U5140 : CLKBUF_X2 port map( I => n21619, Z => n13291);
   U5142 : INV_X1 port map( I => n20735, ZN => n20786);
   U5145 : NOR2_X1 port map( A1 => n3923, A2 => n15307, ZN => n24009);
   U5148 : INV_X1 port map( I => n20921, ZN => n28016);
   U5153 : INV_X2 port map( I => n20728, ZN => n27924);
   U5154 : NAND2_X1 port map( A1 => n1073, A2 => n14183, ZN => n13219);
   U5155 : CLKBUF_X2 port map( I => n21924, Z => n24078);
   U5159 : NAND2_X1 port map( A1 => n6588, A2 => n20516, ZN => n13088);
   U5163 : NAND2_X1 port map( A1 => n3593, A2 => n9377, ZN => n21980);
   U5164 : NOR2_X1 port map( A1 => n3549, A2 => n13900, ZN => n3195);
   U5168 : CLKBUF_X2 port map( I => n21548, Z => n15646);
   U5172 : NOR2_X1 port map( A1 => n21724, A2 => n12290, ZN => n21697);
   U5174 : AOI21_X1 port map( A1 => n21781, A2 => n6046, B => n21693, ZN => 
                           n6805);
   U5177 : CLKBUF_X1 port map( I => n21467, Z => n27885);
   U5182 : AND3_X1 port map( A1 => n21730, A2 => n2569, A3 => n952, Z => n10598
                           );
   U5185 : INV_X2 port map( I => n24538, ZN => n23225);
   U5189 : INV_X1 port map( I => n20885, ZN => n12487);
   U5202 : NAND2_X1 port map( A1 => n6517, A2 => n694, ZN => n12077);
   U5204 : INV_X1 port map( I => n20804, ZN => n6371);
   U5209 : CLKBUF_X2 port map( I => n20816, Z => n14113);
   U5215 : NAND2_X1 port map( A1 => n1085, A2 => n6588, ZN => n25116);
   U5216 : NAND2_X1 port map( A1 => n20927, A2 => n20926, ZN => n20930);
   U5219 : OAI21_X1 port map( A1 => n5753, A2 => n1085, B => n26660, ZN => 
                           n3710);
   U5221 : OAI21_X1 port map( A1 => n13447, A2 => n28428, B => n22511, ZN => 
                           n1737);
   U5222 : OAI21_X1 port map( A1 => n21166, A2 => n27427, B => n21173, ZN => 
                           n4539);
   U5232 : NOR2_X1 port map( A1 => n26942, A2 => n20964, ZN => n4605);
   U5233 : INV_X1 port map( I => n696, ZN => n11380);
   U5234 : INV_X2 port map( I => n694, ZN => n21477);
   U5235 : INV_X2 port map( I => n21166, ZN => n21168);
   U5237 : AOI21_X1 port map( A1 => n21711, A2 => n27248, B => n6802, ZN => 
                           n7348);
   U5239 : OAI21_X1 port map( A1 => n21172, A2 => n21173, B => n11385, ZN => 
                           n2230);
   U5256 : AOI21_X1 port map( A1 => n28308, A2 => n12797, B => n22789, ZN => 
                           n21555);
   U5259 : OAI21_X1 port map( A1 => n803, A2 => n21647, B => n438, ZN => n9848)
                           ;
   U5269 : CLKBUF_X1 port map( I => Key(98), Z => n21476);
   U5270 : CLKBUF_X1 port map( I => Key(27), Z => n21651);
   U5271 : OAI22_X1 port map( A1 => n13073, A2 => n13072, B1 => n20848, B2 => 
                           n20828, ZN => n20829);
   U5279 : INV_X1 port map( I => n14631, ZN => n26566);
   U5281 : INV_X1 port map( I => n21170, ZN => n23021);
   U5282 : CLKBUF_X1 port map( I => Key(69), Z => n20208);
   U5289 : AND2_X2 port map( A1 => n25382, A2 => n24523, Z => n26657);
   U5295 : AND2_X1 port map( A1 => n826, A2 => n23696, Z => n26658);
   U5306 : AND2_X2 port map( A1 => n23456, A2 => n23992, Z => n26659);
   U5308 : OR2_X2 port map( A1 => n5796, A2 => n21924, Z => n26660);
   U5316 : XNOR2_X1 port map( A1 => n11555, A2 => n21044, ZN => n26662);
   U5323 : XNOR2_X1 port map( A1 => n22191, A2 => n25840, ZN => n26663);
   U5324 : XNOR2_X1 port map( A1 => n7052, A2 => n21357, ZN => n26664);
   U5326 : XOR2_X1 port map( A1 => Plaintext(66), A2 => Key(66), Z => n26665);
   U5330 : INV_X1 port map( I => n20294, ZN => n15279);
   U5334 : OR2_X1 port map( A1 => n13167, A2 => n6861, Z => n26667);
   U5339 : OR2_X1 port map( A1 => n26633, A2 => n19870, Z => n26668);
   U5358 : OR2_X1 port map( A1 => n5367, A2 => n20868, Z => n26669);
   U5369 : AND3_X1 port map( A1 => n13389, A2 => n9606, A3 => n17984, Z => 
                           n26670);
   U5373 : AND2_X1 port map( A1 => n2925, A2 => n19727, Z => n26672);
   U5393 : AND2_X2 port map( A1 => n23361, A2 => n10904, Z => n26673);
   U5398 : AND2_X2 port map( A1 => n24567, A2 => n14944, Z => n26675);
   U5405 : OR2_X1 port map( A1 => n14718, A2 => n773, Z => n26676);
   U5424 : NOR2_X1 port map( A1 => n18473, A2 => n24286, ZN => n26678);
   U5426 : OR2_X1 port map( A1 => n14341, A2 => n21058, Z => n26679);
   U5432 : OR2_X1 port map( A1 => n7498, A2 => n10568, Z => n26680);
   U5433 : AND2_X2 port map( A1 => n22834, A2 => n4802, Z => n26681);
   U5434 : AND2_X2 port map( A1 => n28274, A2 => n350, Z => n26682);
   U5441 : OR2_X1 port map( A1 => n27983, A2 => n17526, Z => n26683);
   U5443 : AND2_X1 port map( A1 => n28026, A2 => n945, Z => n26684);
   U5450 : INV_X1 port map( I => n7408, ZN => n11472);
   U5453 : CLKBUF_X4 port map( I => n12885, Z => n10924);
   U5457 : INV_X1 port map( I => n16126, ZN => n15995);
   U5460 : AND2_X1 port map( A1 => n21769, A2 => n14343, Z => n26687);
   U5463 : XNOR2_X1 port map( A1 => n18317, A2 => n27137, ZN => n26688);
   U5466 : AND2_X2 port map( A1 => n13600, A2 => n21136, Z => n26689);
   U5473 : AND2_X1 port map( A1 => n17543, A2 => n24509, Z => n26691);
   U5476 : AND2_X1 port map( A1 => n16326, A2 => n4750, Z => n26692);
   U5478 : AND2_X1 port map( A1 => n19951, A2 => n19827, Z => n26693);
   U5489 : OR2_X1 port map( A1 => n8527, A2 => n11186, Z => n26694);
   U5492 : INV_X1 port map( I => n16618, ZN => n718);
   U5495 : CLKBUF_X2 port map( I => n15182, Z => n7280);
   U5502 : NAND2_X1 port map( A1 => n9911, A2 => n11425, ZN => n26695);
   U5508 : OR2_X1 port map( A1 => n18627, A2 => n7169, Z => n26696);
   U5512 : OR2_X1 port map( A1 => n23977, A2 => n11471, Z => n26698);
   U5518 : OR2_X1 port map( A1 => n14097, A2 => n18687, Z => n26700);
   U5519 : AND2_X1 port map( A1 => n1017, A2 => n5407, Z => n26701);
   U5521 : XNOR2_X1 port map( A1 => Plaintext(91), A2 => Key(91), ZN => n26702)
                           ;
   U5522 : AND2_X1 port map( A1 => n21791, A2 => n10058, Z => n26704);
   U5523 : OR2_X2 port map( A1 => n28525, A2 => n13925, Z => n26705);
   U5529 : AND2_X2 port map( A1 => n20078, A2 => n5080, Z => n26706);
   U5530 : XNOR2_X1 port map( A1 => n1489, A2 => n10051, ZN => n26707);
   U5532 : AND2_X1 port map( A1 => n22153, A2 => n26356, Z => n26708);
   U5537 : INV_X1 port map( I => n28461, ZN => n24641);
   U5545 : AND2_X2 port map( A1 => n28492, A2 => n28384, Z => n26709);
   U5546 : INV_X2 port map( I => n2398, ZN => n14271);
   U5548 : INV_X2 port map( I => n12678, ZN => n16293);
   U5553 : INV_X1 port map( I => n28002, ZN => n20150);
   U5554 : AND2_X2 port map( A1 => n488, A2 => n19880, Z => n26710);
   U5558 : AND2_X2 port map( A1 => n11138, A2 => n10658, Z => n26712);
   U5560 : XNOR2_X1 port map( A1 => n12481, A2 => n7409, ZN => n26713);
   U5576 : CLKBUF_X1 port map( I => n14033, Z => n5449);
   U5577 : OR2_X1 port map( A1 => n13565, A2 => n25492, Z => n26714);
   U5578 : NOR3_X1 port map( A1 => n17751, A2 => n7553, A3 => n5373, ZN => 
                           n26715);
   U5580 : CLKBUF_X1 port map( I => n17522, Z => n22578);
   U5582 : XNOR2_X1 port map( A1 => n18286, A2 => n18008, ZN => n26717);
   U5584 : XNOR2_X1 port map( A1 => n2915, A2 => n27262, ZN => n26718);
   U5587 : CLKBUF_X2 port map( I => n4814, Z => n26533);
   U5603 : XNOR2_X1 port map( A1 => n18048, A2 => n14981, ZN => n26719);
   U5604 : AND2_X2 port map( A1 => n7673, A2 => n7676, Z => n26720);
   U5605 : CLKBUF_X1 port map( I => n18557, Z => n28306);
   U5610 : INV_X2 port map( I => n18557, ZN => n27895);
   U5617 : NAND2_X1 port map( A1 => n5345, A2 => n28362, ZN => n26721);
   U5618 : OR2_X1 port map( A1 => n18871, A2 => n18825, Z => n26722);
   U5619 : INV_X1 port map( I => n19107, ZN => n14545);
   U5620 : XNOR2_X1 port map( A1 => n7744, A2 => n10729, ZN => n26723);
   U5621 : XNOR2_X1 port map( A1 => n19290, A2 => n27444, ZN => n26724);
   U5625 : CLKBUF_X2 port map( I => n5511, Z => n26764);
   U5630 : XNOR2_X1 port map( A1 => n21210, A2 => n22760, ZN => n26725);
   U5646 : XNOR2_X1 port map( A1 => n9002, A2 => n15639, ZN => n26726);
   U5651 : XNOR2_X1 port map( A1 => n19490, A2 => n23917, ZN => n26728);
   U5657 : INV_X1 port map( I => n23278, ZN => n671);
   U5662 : AND2_X1 port map( A1 => n8898, A2 => n20059, Z => n26729);
   U5668 : OR2_X2 port map( A1 => n8910, A2 => n25879, Z => n26730);
   U5669 : OR2_X1 port map( A1 => n4709, A2 => n10794, Z => n26731);
   U5670 : INV_X1 port map( I => n18752, ZN => n27440);
   U5671 : INV_X1 port map( I => n19792, ZN => n12444);
   U5672 : NAND3_X2 port map( A1 => n26732, A2 => n26608, A3 => n26609, ZN => 
                           n9509);
   U5673 : NAND3_X2 port map( A1 => n27172, A2 => n27171, A3 => n17979, ZN => 
                           n26732);
   U5674 : NAND2_X1 port map( A1 => n18624, A2 => n18622, ZN => n28338);
   U5675 : OAI21_X2 port map( A1 => n21772, A2 => n1731, B => n26733, ZN => 
                           n6634);
   U5676 : NAND2_X2 port map( A1 => n11215, A2 => n20326, ZN => n26733);
   U5677 : XOR2_X1 port map( A1 => n9104, A2 => n12604, Z => n25528);
   U5680 : XOR2_X1 port map( A1 => n1097, A2 => n13834, Z => n9104);
   U5686 : XOR2_X1 port map( A1 => n6349, A2 => n28149, Z => n24219);
   U5693 : AOI22_X1 port map( A1 => n7131, A2 => n21208, B1 => n21138, B2 => 
                           n21324, ZN => n27046);
   U5695 : AOI22_X2 port map( A1 => n5944, A2 => n24912, B1 => n14188, B2 => 
                           n13967, ZN => n5943);
   U5698 : NOR2_X2 port map( A1 => n4705, A2 => n13812, ZN => n13967);
   U5700 : NAND3_X2 port map( A1 => n8213, A2 => n8214, A3 => n18166, ZN => 
                           n18816);
   U5710 : INV_X1 port map( I => n2704, ZN => n27700);
   U5715 : OAI22_X2 port map( A1 => n2725, A2 => n2705, B1 => n2318, B2 => 
                           n2317, ZN => n2704);
   U5716 : NAND2_X1 port map( A1 => n19736, A2 => n19735, ZN => n22898);
   U5719 : OAI21_X2 port map( A1 => n14789, A2 => n5253, B => n19570, ZN => 
                           n19736);
   U5720 : XOR2_X1 port map( A1 => n6774, A2 => n6775, Z => n6773);
   U5726 : XOR2_X1 port map( A1 => n19480, A2 => n24312, Z => n6774);
   U5727 : XOR2_X1 port map( A1 => n26737, A2 => n14009, Z => n704);
   U5728 : XOR2_X1 port map( A1 => n5852, A2 => n3812, Z => n26737);
   U5730 : INV_X2 port map( I => n20326, ZN => n26738);
   U5731 : OAI21_X2 port map( A1 => n1024, A2 => n22544, B => n17647, ZN => 
                           n6372);
   U5732 : NAND2_X2 port map( A1 => n14548, A2 => n5368, ZN => n17647);
   U5733 : XOR2_X1 port map( A1 => n19446, A2 => n10494, Z => n7861);
   U5739 : NAND3_X2 port map( A1 => n24630, A2 => n8485, A3 => n9880, ZN => 
                           n19446);
   U5743 : OAI22_X2 port map( A1 => n5051, A2 => n5052, B1 => n5050, B2 => 
                           n16257, ZN => n26814);
   U5745 : NAND2_X1 port map( A1 => n28338, A2 => n1187, ZN => n23201);
   U5746 : AOI22_X2 port map( A1 => n20174, A2 => n24553, B1 => n20269, B2 => 
                           n14221, ZN => n20032);
   U5756 : OAI21_X2 port map( A1 => n9995, A2 => n11111, B => n9992, ZN => 
                           n20174);
   U5760 : XOR2_X1 port map( A1 => n2224, A2 => n20529, Z => n3487);
   U5763 : XOR2_X1 port map( A1 => n8726, A2 => n10445, Z => n2224);
   U5769 : NAND2_X2 port map( A1 => n19014, A2 => n19013, ZN => n26981);
   U5770 : OAI21_X1 port map( A1 => n2952, A2 => n4914, B => n22519, ZN => 
                           n4915);
   U5772 : NAND2_X2 port map( A1 => n2101, A2 => n23337, ZN => n23056);
   U5775 : NAND2_X2 port map( A1 => n26739, A2 => n17687, ZN => n4234);
   U5790 : NAND2_X2 port map( A1 => n17971, A2 => n23365, ZN => n26739);
   U5792 : NOR2_X1 port map( A1 => n2749, A2 => n13718, ZN => n12016);
   U5793 : NAND2_X2 port map( A1 => n26560, A2 => n12588, ZN => n13718);
   U5796 : NAND2_X2 port map( A1 => n26740, A2 => n142, ZN => n27798);
   U5798 : NAND2_X1 port map( A1 => n10215, A2 => n10216, ZN => n26740);
   U5801 : NAND2_X1 port map( A1 => n26022, A2 => n26020, ZN => n27500);
   U5805 : BUF_X2 port map( I => n3891, Z => n26741);
   U5808 : AOI21_X2 port map( A1 => n24340, A2 => n24382, B => n11981, ZN => 
                           n24339);
   U5813 : NOR2_X2 port map( A1 => n22338, A2 => n25586, ZN => n11981);
   U5823 : XOR2_X1 port map( A1 => n5289, A2 => n26742, Z => n27831);
   U5851 : XOR2_X1 port map( A1 => n24848, A2 => n26688, Z => n26742);
   U5854 : OR2_X1 port map( A1 => n2960, A2 => n14426, Z => n17177);
   U5862 : OAI21_X2 port map( A1 => n26222, A2 => n26223, B => n8471, ZN => 
                           n27539);
   U5868 : XOR2_X1 port map( A1 => n9158, A2 => n26743, Z => n4873);
   U5869 : XOR2_X1 port map( A1 => n19093, A2 => n19498, Z => n26743);
   U5874 : NAND2_X2 port map( A1 => n11215, A2 => n9042, ZN => n20491);
   U5879 : OAI22_X1 port map( A1 => n7998, A2 => n7999, B1 => n7348, B2 => 
                           n7347, ZN => n27531);
   U5882 : XOR2_X1 port map( A1 => n24244, A2 => n27343, Z => n19707);
   U5885 : XOR2_X1 port map( A1 => n6220, A2 => n22354, Z => n2076);
   U5890 : NOR3_X1 port map( A1 => n958, A2 => n5573, A3 => n22830, ZN => 
                           n23620);
   U5891 : NOR2_X2 port map( A1 => n26715, A2 => n26670, ZN => n24668);
   U5895 : AOI22_X2 port map( A1 => n26228, A2 => n18405, B1 => n18406, B2 => 
                           n18505, ZN => n22054);
   U5897 : XOR2_X1 port map( A1 => n19479, A2 => n22694, Z => n22693);
   U5904 : XOR2_X1 port map( A1 => n8777, A2 => n19562, Z => n19479);
   U5913 : INV_X1 port map( I => n5510, ZN => n26744);
   U5914 : NAND2_X2 port map( A1 => n18479, A2 => n14594, ZN => n26745);
   U5917 : OR2_X1 port map( A1 => n1806, A2 => n21829, Z => n25119);
   U5918 : XOR2_X1 port map( A1 => n23770, A2 => n8448, Z => n13071);
   U5927 : NAND2_X2 port map( A1 => n23, A2 => n243, ZN => n8448);
   U5928 : XOR2_X1 port map( A1 => n26746, A2 => n20671, Z => Ciphertext(19));
   U5935 : NAND3_X1 port map( A1 => n10410, A2 => n10409, A3 => n10000, ZN => 
                           n26746);
   U5936 : NOR2_X2 port map( A1 => n27498, A2 => n26747, ZN => n6778);
   U5937 : AOI21_X2 port map( A1 => n26696, A2 => n14821, B => n235, ZN => 
                           n26747);
   U5944 : NOR2_X2 port map( A1 => n5908, A2 => n26748, ZN => n5914);
   U5950 : AOI21_X2 port map( A1 => n14134, A2 => n22012, B => n5906, ZN => 
                           n26748);
   U5951 : XOR2_X1 port map( A1 => n26749, A2 => n10544, Z => Ciphertext(164));
   U5955 : NOR2_X1 port map( A1 => n26497, A2 => n26789, ZN => n26749);
   U5962 : NAND3_X2 port map( A1 => n8769, A2 => n224, A3 => n19100, ZN => 
                           n20238);
   U5967 : NAND2_X1 port map( A1 => n28452, A2 => n20660, ZN => n25125);
   U5969 : NAND3_X2 port map( A1 => n26750, A2 => n8390, A3 => n28493, ZN => 
                           n19968);
   U5970 : NAND2_X1 port map( A1 => n19622, A2 => n969, ZN => n26750);
   U5976 : NOR3_X2 port map( A1 => n21812, A2 => n27325, A3 => n27005, ZN => 
                           n15414);
   U5977 : CLKBUF_X4 port map( I => n13437, Z => n3291);
   U5982 : INV_X4 port map( I => n6766, ZN => n9484);
   U5986 : INV_X4 port map( I => n26751, ZN => n5990);
   U5991 : AND2_X2 port map( A1 => n5991, A2 => n7678, Z => n26751);
   U5994 : XOR2_X1 port map( A1 => n21145, A2 => n14551, Z => n20361);
   U5998 : NAND3_X2 port map( A1 => n27158, A2 => n20332, A3 => n10741, ZN => 
                           n21145);
   U5999 : AOI22_X2 port map( A1 => n24922, A2 => n6803, B1 => n13718, B2 => 
                           n2749, ZN => n9267);
   U6000 : NAND2_X2 port map( A1 => n25119, A2 => n26752, ZN => n14513);
   U6002 : AOI22_X2 port map( A1 => n670, A2 => n10611, B1 => n1804, B2 => 
                           n28264, ZN => n26752);
   U6003 : XNOR2_X1 port map( A1 => n2515, A2 => n27848, ZN => n26143);
   U6005 : NOR2_X2 port map( A1 => n27383, A2 => n22438, ZN => n14551);
   U6010 : OAI22_X1 port map( A1 => n6798, A2 => n21531, B1 => n770, B2 => 
                           n26753, ZN => n23634);
   U6011 : OR2_X1 port map( A1 => n21538, A2 => n4827, Z => n26753);
   U6012 : NAND2_X2 port map( A1 => n6913, A2 => n7078, ZN => n7485);
   U6027 : XOR2_X1 port map( A1 => n24498, A2 => n26755, Z => n7189);
   U6028 : XOR2_X1 port map( A1 => n9662, A2 => n28294, Z => n26755);
   U6029 : NAND2_X1 port map( A1 => n27671, A2 => n26756, ZN => n24596);
   U6038 : INV_X1 port map( I => n27175, ZN => n23583);
   U6042 : NAND3_X2 port map( A1 => n6650, A2 => n6649, A3 => n28379, ZN => 
                           n27175);
   U6044 : NAND2_X2 port map( A1 => n17379, A2 => n26757, ZN => n18180);
   U6045 : NAND2_X2 port map( A1 => n27115, A2 => n27116, ZN => n26757);
   U6047 : AOI22_X2 port map( A1 => n26673, A2 => n1179, B1 => n18778, B2 => 
                           n27457, ZN => n22047);
   U6049 : NOR2_X2 port map( A1 => n5845, A2 => n27313, ZN => n8978);
   U6051 : NOR2_X2 port map( A1 => n25608, A2 => n8986, ZN => n5845);
   U6053 : NAND2_X1 port map( A1 => n15984, A2 => n15835, ZN => n15836);
   U6055 : XOR2_X1 port map( A1 => n10029, A2 => n12382, Z => n13458);
   U6060 : NAND2_X2 port map( A1 => n24172, A2 => n11556, ZN => n10029);
   U6061 : INV_X2 port map( I => n20826, ZN => n20848);
   U6063 : NAND2_X2 port map( A1 => n13056, A2 => n8760, ZN => n20826);
   U6064 : BUF_X2 port map( I => n8937, Z => n26758);
   U6067 : XOR2_X1 port map( A1 => Plaintext(70), A2 => Key(70), Z => n27002);
   U6071 : AOI22_X2 port map( A1 => n21134, A2 => n20263, B1 => n12945, B2 => 
                           n12944, ZN => n3627);
   U6072 : INV_X1 port map( I => n12042, ZN => n20434);
   U6077 : AOI21_X2 port map( A1 => n20821, A2 => n27066, B => n20819, ZN => 
                           n8760);
   U6078 : NAND2_X2 port map( A1 => n26315, A2 => n26961, ZN => n11215);
   U6079 : NAND2_X1 port map( A1 => n10555, A2 => n22799, ZN => n11617);
   U6081 : NAND2_X2 port map( A1 => n26451, A2 => n26485, ZN => n21861);
   U6082 : OAI22_X2 port map( A1 => n16724, A2 => n28369, B1 => n8249, B2 => 
                           n16524, ZN => n3171);
   U6091 : NAND2_X2 port map( A1 => n26518, A2 => n7395, ZN => n16724);
   U6092 : OAI22_X2 port map( A1 => n26759, A2 => n26655, B1 => n17224, B2 => 
                           n1039, ZN => n14212);
   U6096 : INV_X2 port map( I => n17255, ZN => n26759);
   U6101 : NOR2_X2 port map( A1 => n17490, A2 => n4536, ZN => n17255);
   U6103 : AND2_X1 port map( A1 => n15834, A2 => n26068, Z => n4380);
   U6105 : INV_X1 port map( I => n19523, ZN => n28009);
   U6106 : AND2_X1 port map( A1 => n9563, A2 => n20704, Z => n28376);
   U6107 : INV_X1 port map( I => n17064, ZN => n28070);
   U6108 : NAND3_X1 port map( A1 => n27217, A2 => n6830, A3 => n13526, ZN => 
                           n27221);
   U6109 : OR2_X1 port map( A1 => n27492, A2 => n11982, Z => n5040);
   U6113 : BUF_X2 port map( I => n7052, Z => n26761);
   U6118 : NOR2_X1 port map( A1 => n27657, A2 => n27656, ZN => n24723);
   U6119 : OAI21_X2 port map( A1 => n15099, A2 => n10875, B => n17372, ZN => 
                           n26197);
   U6120 : AOI22_X1 port map( A1 => n13621, A2 => n17974, B1 => n13620, B2 => 
                           n12815, ZN => n27610);
   U6121 : AOI22_X2 port map( A1 => n26685, A2 => n13872, B1 => n19138, B2 => 
                           n24937, ZN => n22640);
   U6124 : XOR2_X1 port map( A1 => n28358, A2 => n19392, Z => n19486);
   U6125 : XOR2_X1 port map( A1 => n22637, A2 => n11667, Z => n18686);
   U6126 : XOR2_X1 port map( A1 => n24088, A2 => n1192, Z => n11667);
   U6129 : OAI21_X2 port map( A1 => n24570, A2 => n14826, B => n23692, ZN => 
                           n18090);
   U6132 : OAI21_X2 port map( A1 => n27236, A2 => n26763, B => n5606, ZN => 
                           n20189);
   U6133 : NOR2_X2 port map( A1 => n19721, A2 => n19722, ZN => n20255);
   U6134 : AOI22_X2 port map( A1 => n19825, A2 => n25014, B1 => n3190, B2 => 
                           n24392, ZN => n19721);
   U6136 : INV_X2 port map( I => n26766, ZN => n26415);
   U6138 : XOR2_X1 port map( A1 => n19426, A2 => n19425, Z => n26766);
   U6144 : XOR2_X1 port map( A1 => n16627, A2 => n9456, Z => n23637);
   U6145 : XOR2_X1 port map( A1 => n1789, A2 => n27296, Z => n15529);
   U6150 : NAND2_X1 port map( A1 => n24933, A2 => n17878, ZN => n24221);
   U6157 : XOR2_X1 port map( A1 => n6275, A2 => n5653, Z => n19424);
   U6164 : NAND2_X2 port map( A1 => n22420, A2 => n8131, ZN => n6275);
   U6165 : OR2_X2 port map( A1 => n9095, A2 => n14224, Z => n12734);
   U6168 : NAND2_X1 port map( A1 => n26616, A2 => n17325, ZN => n17450);
   U6172 : AOI22_X2 port map( A1 => n26768, A2 => n4715, B1 => n8275, B2 => 
                           n17433, ZN => n23859);
   U6174 : NOR2_X2 port map( A1 => n17433, A2 => n17436, ZN => n26768);
   U6177 : XOR2_X1 port map( A1 => n4211, A2 => n26769, Z => n15545);
   U6178 : XOR2_X1 port map( A1 => n2306, A2 => n2201, Z => n26769);
   U6180 : OAI22_X2 port map( A1 => n10428, A2 => n964, B1 => n15560, B2 => 
                           n9994, ZN => n9186);
   U6189 : XOR2_X1 port map( A1 => n26770, A2 => n8091, Z => Ciphertext(86));
   U6191 : AOI22_X2 port map( A1 => n26170, A2 => n2052, B1 => n26419, B2 => 
                           n26157, ZN => n26770);
   U6193 : OAI21_X2 port map( A1 => n26689, A2 => n26771, B => n21175, ZN => 
                           n24831);
   U6207 : AOI22_X2 port map( A1 => n27265, A2 => n26772, B1 => n5188, B2 => 
                           n21175, ZN => n26847);
   U6210 : INV_X1 port map( I => n15454, ZN => n26774);
   U6213 : OAI21_X2 port map( A1 => n26775, A2 => n5704, B => n9508, ZN => 
                           n10841);
   U6218 : NOR2_X2 port map( A1 => n14683, A2 => n11425, ZN => n26775);
   U6222 : NAND2_X1 port map( A1 => n28271, A2 => n28270, ZN => n28191);
   U6227 : XOR2_X1 port map( A1 => n26776, A2 => n6891, Z => n7218);
   U6228 : XOR2_X1 port map( A1 => n3411, A2 => n16958, Z => n26776);
   U6229 : NAND2_X1 port map( A1 => n26779, A2 => n26777, ZN => n18845);
   U6235 : OAI21_X1 port map( A1 => n18921, A2 => n4549, B => n26778, ZN => 
                           n26777);
   U6237 : INV_X2 port map( I => n2346, ZN => n26778);
   U6240 : NAND2_X1 port map( A1 => n18841, A2 => n2346, ZN => n26779);
   U6241 : AOI22_X1 port map( A1 => n26675, A2 => n25504, B1 => n17247, B2 => 
                           n14944, ZN => n25521);
   U6247 : NOR2_X2 port map( A1 => n24567, A2 => n17492, ZN => n17247);
   U6250 : NAND2_X2 port map( A1 => n26780, A2 => n28500, ZN => n20770);
   U6254 : NOR2_X2 port map( A1 => n9010, A2 => n13399, ZN => n26780);
   U6255 : AOI21_X2 port map( A1 => n14253, A2 => n26781, B => n6627, ZN => 
                           n283);
   U6263 : OAI21_X2 port map( A1 => n27931, A2 => n13570, B => n765, ZN => 
                           n26781);
   U6270 : XOR2_X1 port map( A1 => n26707, A2 => n18216, Z => n28482);
   U6271 : OAI22_X2 port map( A1 => n12403, A2 => n26783, B1 => n5759, B2 => 
                           n18465, ZN => n26163);
   U6272 : NAND2_X2 port map( A1 => n18465, A2 => n18684, ZN => n26783);
   U6276 : XOR2_X1 port map( A1 => n25901, A2 => n8790, Z => n18203);
   U6277 : XOR2_X1 port map( A1 => n21366, A2 => n26784, Z => n5492);
   U6279 : XOR2_X1 port map( A1 => n954, A2 => n10352, Z => n26784);
   U6280 : AOI22_X2 port map( A1 => n26708, A2 => n2403, B1 => n11483, B2 => 
                           n17842, ZN => n26794);
   U6281 : NAND2_X2 port map( A1 => n12643, A2 => n20168, ZN => n20029);
   U6284 : NAND2_X2 port map( A1 => n7211, A2 => n27681, ZN => n12643);
   U6285 : BUF_X4 port map( I => n12360, Z => n27704);
   U6287 : NOR2_X2 port map( A1 => n26886, A2 => n26629, ZN => n27074);
   U6288 : NAND2_X2 port map( A1 => n26785, A2 => n3832, ZN => n3830);
   U6289 : AOI22_X2 port map( A1 => n15518, A2 => n4703, B1 => n3833, B2 => 
                           n3312, ZN => n26785);
   U6291 : NOR2_X2 port map( A1 => n26787, A2 => n26786, ZN => n21135);
   U6295 : INV_X1 port map( I => n15709, ZN => n26786);
   U6296 : INV_X2 port map( I => n15454, ZN => n26787);
   U6297 : NAND2_X2 port map( A1 => n22603, A2 => n26788, ZN => n3292);
   U6300 : OR2_X1 port map( A1 => n4843, A2 => n4887, Z => n26788);
   U6301 : NAND2_X1 port map( A1 => n28087, A2 => n2228, ZN => n3583);
   U6304 : NAND2_X2 port map( A1 => n8049, A2 => n7030, ZN => n7995);
   U6305 : NAND2_X2 port map( A1 => n13244, A2 => n15132, ZN => n8049);
   U6306 : OAI21_X2 port map( A1 => n27270, A2 => n27271, B => n21097, ZN => 
                           n14870);
   U6309 : XOR2_X1 port map( A1 => n27145, A2 => n9748, Z => n18162);
   U6315 : NAND3_X2 port map( A1 => n17945, A2 => n7322, A3 => n26860, ZN => 
                           n27145);
   U6320 : XOR2_X1 port map( A1 => n3977, A2 => n15727, Z => n15728);
   U6332 : NAND2_X2 port map( A1 => n11250, A2 => n11249, ZN => n24381);
   U6336 : NAND2_X2 port map( A1 => n25150, A2 => n9823, ZN => n11250);
   U6337 : OAI21_X2 port map( A1 => n16540, A2 => n14562, B => n26790, ZN => 
                           n15012);
   U6339 : NAND3_X2 port map( A1 => n14562, A2 => n145, A3 => n23048, ZN => 
                           n26790);
   U6342 : NOR2_X2 port map( A1 => n14310, A2 => n26791, ZN => n7185);
   U6346 : OAI22_X2 port map( A1 => n13990, A2 => n16038, B1 => n16334, B2 => 
                           n769, ZN => n26791);
   U6348 : XOR2_X1 port map( A1 => n1041, A2 => n17141, Z => n13293);
   U6349 : NAND2_X1 port map( A1 => n7814, A2 => n19167, ZN => n27142);
   U6355 : BUF_X4 port map( I => n20345, Z => n21666);
   U6357 : AOI22_X1 port map( A1 => n18983, A2 => n22385, B1 => n18984, B2 => 
                           n1149, ZN => n18985);
   U6358 : NAND3_X1 port map( A1 => n19117, A2 => n28547, A3 => n997, ZN => 
                           n10976);
   U6360 : NAND2_X1 port map( A1 => n22744, A2 => n19921, ZN => n26207);
   U6362 : XOR2_X1 port map( A1 => n6475, A2 => n26792, Z => n24938);
   U6366 : XOR2_X1 port map( A1 => n28488, A2 => n26793, Z => n26792);
   U6368 : BUF_X1 port map( I => n7749, Z => n23368);
   U6371 : NAND2_X2 port map( A1 => n11256, A2 => n22199, ZN => n15242);
   U6373 : NOR2_X2 port map( A1 => n15667, A2 => n19925, ZN => n3121);
   U6374 : NAND2_X1 port map( A1 => n201, A2 => n203, ZN => n21576);
   U6375 : NAND2_X2 port map( A1 => n17611, A2 => n26794, ZN => n14139);
   U6381 : NAND2_X1 port map( A1 => n17919, A2 => n17580, ZN => n17582);
   U6391 : NAND3_X2 port map( A1 => n24103, A2 => n13536, A3 => n13534, ZN => 
                           n17919);
   U6397 : XNOR2_X1 port map( A1 => n13131, A2 => n2268, ZN => n27242);
   U6400 : NOR2_X2 port map( A1 => n22128, A2 => n26795, ZN => n27944);
   U6402 : NOR2_X2 port map( A1 => n24361, A2 => n19113, ZN => n26795);
   U6405 : NAND2_X2 port map( A1 => n17214, A2 => n17541, ZN => n26796);
   U6411 : NAND3_X2 port map( A1 => n2021, A2 => n13148, A3 => n22744, ZN => 
                           n2023);
   U6412 : NAND2_X1 port map( A1 => n27696, A2 => n5616, ZN => n50);
   U6416 : AOI21_X2 port map( A1 => n17649, A2 => n12611, B => n26797, ZN => 
                           n18244);
   U6417 : OAI22_X2 port map( A1 => n17750, A2 => n12590, B1 => n12611, B2 => 
                           n12930, ZN => n26797);
   U6421 : OR2_X1 port map( A1 => n26646, A2 => n15937, Z => n4456);
   U6422 : NAND2_X1 port map( A1 => n21604, A2 => n13922, ZN => n22892);
   U6424 : OAI22_X2 port map( A1 => n27811, A2 => n9977, B1 => n21715, B2 => 
                           n8823, ZN => n24400);
   U6425 : AOI22_X2 port map( A1 => n20644, A2 => n20587, B1 => n9979, B2 => 
                           n10666, ZN => n8823);
   U6428 : XOR2_X1 port map( A1 => n26798, A2 => n20605, Z => Ciphertext(2));
   U6429 : NAND2_X1 port map( A1 => n25675, A2 => n27275, ZN => n26798);
   U6430 : AOI21_X2 port map( A1 => n10993, A2 => n15449, B => n18487, ZN => 
                           n27664);
   U6432 : NAND2_X2 port map( A1 => n13969, A2 => n448, ZN => n10993);
   U6433 : NOR2_X2 port map( A1 => n17006, A2 => n22092, ZN => n7481);
   U6435 : XOR2_X1 port map( A1 => n20429, A2 => n2520, Z => n8595);
   U6436 : XOR2_X1 port map( A1 => n2292, A2 => n4383, Z => n20429);
   U6442 : XOR2_X1 port map( A1 => n8879, A2 => n20550, Z => n21238);
   U6446 : NAND2_X2 port map( A1 => n28410, A2 => n8461, ZN => n8879);
   U6448 : AOI21_X2 port map( A1 => n8172, A2 => n7682, B => n19705, ZN => 
                           n27652);
   U6452 : NOR3_X1 port map( A1 => n23719, A2 => n27543, A3 => n24812, ZN => 
                           n1746);
   U6456 : XOR2_X1 port map( A1 => n26799, A2 => n14650, Z => Ciphertext(98));
   U6458 : NAND2_X1 port map( A1 => n5482, A2 => n22585, ZN => n26799);
   U6459 : XOR2_X1 port map( A1 => n26800, A2 => n23021, Z => Ciphertext(106));
   U6460 : NOR2_X1 port map( A1 => n15205, A2 => n500, ZN => n26800);
   U6462 : NAND2_X2 port map( A1 => n4472, A2 => n17370, ZN => n25179);
   U6463 : NAND3_X2 port map( A1 => n26801, A2 => n4474, A3 => n4475, ZN => 
                           n5780);
   U6467 : NAND2_X2 port map( A1 => n26645, A2 => n11485, ZN => n2701);
   U6468 : XOR2_X1 port map( A1 => n1671, A2 => n24377, Z => n27401);
   U6472 : XOR2_X1 port map( A1 => n11675, A2 => n14091, Z => n1671);
   U6473 : XOR2_X1 port map( A1 => n24163, A2 => n26802, Z => n23567);
   U6474 : XOR2_X1 port map( A1 => n902, A2 => n699, Z => n26802);
   U6475 : XOR2_X1 port map( A1 => n20547, A2 => n20536, Z => n20351);
   U6476 : XOR2_X1 port map( A1 => n20580, A2 => n20435, Z => n20547);
   U6477 : NAND2_X1 port map( A1 => n23037, A2 => n27865, ZN => n27546);
   U6479 : INV_X2 port map( I => n22905, ZN => n6042);
   U6480 : XOR2_X1 port map( A1 => n6174, A2 => n27782, Z => n22905);
   U6481 : XOR2_X1 port map( A1 => n23917, A2 => n21607, Z => n19546);
   U6482 : NOR2_X2 port map( A1 => n8711, A2 => n27034, ZN => n23917);
   U6483 : INV_X2 port map( I => n2706, ZN => n5664);
   U6489 : OAI22_X2 port map( A1 => n3391, A2 => n9878, B1 => n6954, B2 => 
                           n10411, ZN => n2706);
   U6490 : AOI21_X1 port map( A1 => n253, A2 => n5292, B => n4393, ZN => n27383
                           );
   U6496 : OAI22_X1 port map( A1 => n16454, A2 => n28083, B1 => n16456, B2 => 
                           n8021, ZN => n16459);
   U6499 : NAND3_X2 port map( A1 => n24135, A2 => n510, A3 => n19768, ZN => 
                           n26803);
   U6501 : BUF_X8 port map( I => n7289, Z => n4739);
   U6504 : NAND2_X1 port map( A1 => n9644, A2 => n25081, ZN => n26804);
   U6509 : NAND2_X2 port map( A1 => n26805, A2 => n8412, ZN => n3891);
   U6511 : NAND2_X1 port map( A1 => n2004, A2 => n15457, ZN => n26805);
   U6512 : INV_X2 port map( I => n26806, ZN => n25305);
   U6515 : XOR2_X1 port map( A1 => n8429, A2 => n8428, Z => n26806);
   U6516 : NOR3_X2 port map( A1 => n25241, A2 => n21561, A3 => n24635, ZN => 
                           n26813);
   U6518 : BUF_X2 port map( I => n27690, Z => n26807);
   U6520 : XOR2_X1 port map( A1 => n19174, A2 => n8224, Z => n1943);
   U6523 : XOR2_X1 port map( A1 => n19388, A2 => n2164, Z => n8224);
   U6526 : NOR2_X2 port map( A1 => n22438, A2 => n22437, ZN => n7848);
   U6527 : AOI22_X2 port map( A1 => n26808, A2 => n20865, B1 => n8495, B2 => 
                           n1073, ZN => n20680);
   U6530 : NAND2_X2 port map( A1 => n6651, A2 => n5071, ZN => n26808);
   U6532 : NOR3_X1 port map( A1 => n23154, A2 => n696, A3 => n843, ZN => n9847)
                           ;
   U6534 : NAND2_X2 port map( A1 => n17539, A2 => n8978, ZN => n17552);
   U6536 : NAND2_X2 port map( A1 => n15266, A2 => n11984, ZN => n114);
   U6537 : NOR2_X1 port map( A1 => n18837, A2 => n1149, ZN => n1704);
   U6542 : NAND3_X2 port map( A1 => n7740, A2 => n7738, A3 => n7742, ZN => 
                           n6301);
   U6543 : XOR2_X1 port map( A1 => n26809, A2 => n549, Z => n5194);
   U6550 : XOR2_X1 port map( A1 => n19166, A2 => n19477, Z => n26809);
   U6553 : XOR2_X1 port map( A1 => n7744, A2 => n26810, Z => n6307);
   U6558 : XOR2_X1 port map( A1 => n18172, A2 => n27702, Z => n26810);
   U6559 : NAND2_X2 port map( A1 => n26811, A2 => n6749, ZN => n6559);
   U6560 : NOR2_X2 port map( A1 => n26812, A2 => n7684, ZN => n22022);
   U6561 : NOR2_X2 port map( A1 => n28031, A2 => n13963, ZN => n26812);
   U6562 : NAND3_X2 port map( A1 => n11924, A2 => n10622, A3 => n26855, ZN => 
                           n28206);
   U6563 : NAND2_X2 port map( A1 => n14227, A2 => n4501, ZN => n3908);
   U6568 : NOR2_X2 port map( A1 => n24917, A2 => n22071, ZN => n4501);
   U6571 : XOR2_X1 port map( A1 => n26813, A2 => n15798, Z => Ciphertext(153));
   U6578 : INV_X2 port map( I => n3846, ZN => n27862);
   U6579 : OAI21_X2 port map( A1 => n24693, A2 => n13502, B => n18827, ZN => 
                           n26457);
   U6580 : XOR2_X1 port map( A1 => n8383, A2 => n26815, Z => n27027);
   U6582 : INV_X2 port map( I => n14754, ZN => n26815);
   U6583 : NAND2_X2 port map( A1 => n8381, A2 => n4469, ZN => n8383);
   U6584 : NAND3_X1 port map( A1 => n8388, A2 => n25329, A3 => n20704, ZN => 
                           n20701);
   U6587 : OR2_X2 port map( A1 => n10571, A2 => n11610, Z => n4446);
   U6590 : INV_X2 port map( I => n26816, ZN => n26623);
   U6594 : XNOR2_X1 port map( A1 => n8863, A2 => n13107, ZN => n26816);
   U6596 : NAND3_X2 port map( A1 => n15034, A2 => n15036, A3 => n20595, ZN => 
                           n6997);
   U6597 : XOR2_X1 port map( A1 => n26817, A2 => n20411, Z => n20787);
   U6602 : XOR2_X1 port map( A1 => n13190, A2 => n13189, Z => n26817);
   U6603 : XOR2_X1 port map( A1 => n22705, A2 => n26818, Z => n14348);
   U6604 : XOR2_X1 port map( A1 => n20012, A2 => n6068, Z => n26818);
   U6607 : NAND2_X2 port map( A1 => n2413, A2 => n22871, ZN => n3525);
   U6611 : NAND2_X2 port map( A1 => n26819, A2 => n9103, ZN => n20176);
   U6612 : NAND2_X2 port map( A1 => n23591, A2 => n23593, ZN => n26819);
   U6614 : NAND2_X2 port map( A1 => n26820, A2 => n11401, ZN => n12411);
   U6615 : NAND3_X2 port map( A1 => n11400, A2 => n15597, A3 => n4739, ZN => 
                           n26820);
   U6616 : XNOR2_X1 port map( A1 => n19510, A2 => n19489, ZN => n19288);
   U6620 : NOR2_X2 port map( A1 => n26943, A2 => n24813, ZN => n19489);
   U6626 : NAND2_X1 port map( A1 => n6833, A2 => n6832, ZN => n27217);
   U6629 : XOR2_X1 port map( A1 => n18111, A2 => n24663, Z => n22592);
   U6634 : XOR2_X1 port map( A1 => n27320, A2 => n761, Z => n18111);
   U6637 : NAND3_X2 port map( A1 => n26829, A2 => n14718, A3 => n25304, ZN => 
                           n12064);
   U6639 : AOI22_X1 port map( A1 => n22216, A2 => n20128, B1 => n26944, B2 => 
                           n11372, ZN => n5224);
   U6644 : NAND2_X2 port map( A1 => n24988, A2 => n24987, ZN => n26944);
   U6649 : AOI21_X2 port map( A1 => n8130, A2 => n11826, B => n26821, ZN => 
                           n22420);
   U6652 : NAND2_X2 port map( A1 => n114, A2 => n18891, ZN => n18837);
   U6656 : INV_X2 port map( I => n1149, ZN => n26822);
   U6658 : BUF_X2 port map( I => n16784, Z => n26823);
   U6660 : XOR2_X1 port map( A1 => n26824, A2 => n20585, Z => Ciphertext(77));
   U6662 : AOI22_X1 port map( A1 => n20583, A2 => n21008, B1 => n15678, B2 => 
                           n24764, ZN => n26824);
   U6663 : NAND3_X2 port map( A1 => n26825, A2 => n14602, A3 => n5048, ZN => 
                           n14951);
   U6666 : BUF_X4 port map( I => n7832, Z => n2140);
   U6668 : OAI22_X2 port map( A1 => n9845, A2 => n24998, B1 => n11593, B2 => 
                           n20261, ZN => n22888);
   U6670 : NAND2_X2 port map( A1 => n24998, A2 => n19978, ZN => n20261);
   U6673 : NAND2_X2 port map( A1 => n26826, A2 => n18501, ZN => n22385);
   U6674 : NAND2_X1 port map( A1 => n14204, A2 => n14206, ZN => n26826);
   U6677 : OR2_X1 port map( A1 => n15642, A2 => n11795, Z => n15169);
   U6680 : INV_X1 port map( I => n26807, ZN => n15146);
   U6681 : XOR2_X1 port map( A1 => n17121, A2 => n17123, Z => n25181);
   U6682 : XOR2_X1 port map( A1 => n26996, A2 => n25582, Z => n17121);
   U6689 : NAND2_X1 port map( A1 => n21595, A2 => n21604, ZN => n26827);
   U6691 : AOI21_X2 port map( A1 => n1601, A2 => n26828, B => n19906, ZN => 
                           n26611);
   U6693 : XOR2_X1 port map( A1 => n9918, A2 => n12959, Z => n7813);
   U6695 : AOI21_X2 port map( A1 => n6449, A2 => n20262, B => n22888, ZN => 
                           n12959);
   U6698 : XOR2_X1 port map( A1 => n26830, A2 => n4208, Z => n4209);
   U6703 : XOR2_X1 port map( A1 => n7812, A2 => n6616, Z => n26830);
   U6709 : INV_X2 port map( I => n21563, ZN => n22789);
   U6713 : NAND2_X2 port map( A1 => n25422, A2 => n25863, ZN => n21563);
   U6714 : AOI21_X1 port map( A1 => n5344, A2 => n13128, B => n13125, ZN => 
                           n26954);
   U6716 : NAND2_X2 port map( A1 => n23746, A2 => n18985, ZN => n19510);
   U6719 : NAND2_X2 port map( A1 => n14210, A2 => n18544, ZN => n18548);
   U6720 : NAND2_X2 port map( A1 => n10278, A2 => n10203, ZN => n14210);
   U6722 : AOI22_X1 port map( A1 => n3583, A2 => n4307, B1 => n11108, B2 => 
                           n12845, ZN => n25945);
   U6723 : OAI21_X1 port map( A1 => n1003, A2 => n6042, B => n23415, ZN => 
                           n18496);
   U6724 : NAND2_X1 port map( A1 => n11923, A2 => n25952, ZN => n6882);
   U6729 : NAND2_X2 port map( A1 => n25521, A2 => n5146, ZN => n14446);
   U6734 : OR2_X1 port map( A1 => n19798, A2 => n13824, Z => n26381);
   U6735 : XOR2_X1 port map( A1 => n14570, A2 => n26832, Z => n15739);
   U6736 : XOR2_X1 port map( A1 => n19435, A2 => n26833, Z => n26832);
   U6739 : INV_X2 port map( I => n19560, ZN => n26833);
   U6741 : XOR2_X1 port map( A1 => n20722, A2 => n20721, Z => n22919);
   U6742 : NAND2_X2 port map( A1 => n5320, A2 => n24429, ZN => n11984);
   U6743 : OAI22_X2 port map( A1 => n6041, A2 => n1003, B1 => n18750, B2 => 
                           n18752, ZN => n5320);
   U6744 : AND2_X1 port map( A1 => n26646, A2 => n8264, Z => n16302);
   U6745 : XOR2_X1 port map( A1 => n9791, A2 => n19487, Z => n19383);
   U6749 : AOI21_X2 port map( A1 => n15100, A2 => n26152, B => n26709, ZN => 
                           n9791);
   U6752 : NAND3_X2 port map( A1 => n19598, A2 => n1120, A3 => n19597, ZN => 
                           n9400);
   U6755 : XOR2_X1 port map( A1 => n18070, A2 => n26058, Z => n18328);
   U6758 : AOI22_X2 port map( A1 => n11282, A2 => n7140, B1 => n6691, B2 => 
                           n11281, ZN => n18070);
   U6759 : NOR2_X1 port map( A1 => n730, A2 => n11407, ZN => n3772);
   U6761 : XOR2_X1 port map( A1 => n21979, A2 => n8879, Z => n20521);
   U6763 : XOR2_X1 port map( A1 => n4188, A2 => n26834, Z => n18710);
   U6767 : XOR2_X1 port map( A1 => n18334, A2 => n590, Z => n26834);
   U6774 : AOI22_X2 port map( A1 => n10983, A2 => n17844, B1 => n10982, B2 => 
                           n16971, ZN => n18161);
   U6776 : NAND2_X2 port map( A1 => n1780, A2 => n9485, ZN => n17844);
   U6782 : NAND2_X2 port map( A1 => n17523, A2 => n6620, ZN => n9250);
   U6789 : OAI21_X2 port map( A1 => n28037, A2 => n28038, B => n27146, ZN => 
                           n17523);
   U6806 : BUF_X4 port map( I => n13467, Z => n11196);
   U6815 : BUF_X4 port map( I => n17497, Z => n24162);
   U6819 : BUF_X4 port map( I => n10422, Z => n26835);
   U6820 : NAND3_X2 port map( A1 => n5854, A2 => n26837, A3 => n26836, ZN => 
                           n25328);
   U6823 : XOR2_X1 port map( A1 => n20767, A2 => n20447, Z => n21303);
   U6824 : NAND2_X2 port map( A1 => n23674, A2 => n22815, ZN => n20130);
   U6828 : NAND3_X1 port map( A1 => n19770, A2 => n26839, A3 => n15471, ZN => 
                           n19771);
   U6830 : NOR2_X1 port map( A1 => n26949, A2 => n22537, ZN => n14921);
   U6832 : NOR2_X2 port map( A1 => n26870, A2 => n9097, ZN => n23029);
   U6833 : AOI21_X2 port map( A1 => n21829, A2 => n10957, B => n10951, ZN => 
                           n3578);
   U6834 : NOR2_X2 port map( A1 => n27606, A2 => n27607, ZN => n21829);
   U6841 : NAND2_X2 port map( A1 => n3870, A2 => n20253, ZN => n15285);
   U6843 : NOR2_X1 port map( A1 => n775, A2 => n26840, ZN => n23934);
   U6855 : XOR2_X1 port map( A1 => n25345, A2 => n19522, Z => n19555);
   U6862 : OAI21_X2 port map( A1 => n1811, A2 => n1814, B => n1809, ZN => 
                           n25345);
   U6887 : OAI22_X2 port map( A1 => n27455, A2 => n28551, B1 => n14281, B2 => 
                           n13900, ZN => n21397);
   U6888 : NOR2_X2 port map( A1 => n8970, A2 => n26841, ZN => n13415);
   U6889 : AOI21_X2 port map( A1 => n26982, A2 => n8972, B => n16283, ZN => 
                           n26841);
   U6898 : XOR2_X1 port map( A1 => n26842, A2 => n19329, Z => n19806);
   U6899 : XOR2_X1 port map( A1 => n4615, A2 => n27470, Z => n26842);
   U6905 : XOR2_X1 port map( A1 => n2615, A2 => n9748, Z => n18087);
   U6906 : OAI21_X2 port map( A1 => n26316, A2 => n4459, B => n4458, ZN => 
                           n2615);
   U6907 : OAI22_X2 port map( A1 => n26843, A2 => n25468, B1 => n19085, B2 => 
                           n7970, ZN => n8120);
   U6908 : NAND2_X1 port map( A1 => n26607, A2 => n19110, ZN => n26843);
   U6911 : OAI21_X1 port map( A1 => n7312, A2 => n26436, B => n21587, ZN => 
                           n10376);
   U6912 : XOR2_X1 port map( A1 => n16757, A2 => n17095, Z => n16440);
   U6915 : XOR2_X1 port map( A1 => n17084, A2 => n16819, Z => n16757);
   U6926 : AOI21_X2 port map( A1 => n26413, A2 => n11465, B => n6552, ZN => 
                           n14221);
   U6927 : INV_X4 port map( I => n27871, ZN => n27830);
   U6935 : AOI22_X2 port map( A1 => n26879, A2 => n730, B1 => n16197, B2 => 
                           n3773, ZN => n8239);
   U6936 : XOR2_X1 port map( A1 => n26844, A2 => n20683, Z => Ciphertext(22));
   U6941 : NAND2_X2 port map( A1 => n26845, A2 => n1029, ZN => n25666);
   U6942 : NAND2_X2 port map( A1 => n12634, A2 => n10298, ZN => n26845);
   U6947 : NOR2_X2 port map( A1 => n27804, A2 => n26846, ZN => n8155);
   U6948 : NOR3_X2 port map( A1 => n8275, A2 => n22865, A3 => n28389, ZN => 
                           n26846);
   U6951 : XOR2_X1 port map( A1 => n22879, A2 => n18155, Z => n18327);
   U6963 : NOR2_X2 port map( A1 => n17267, A2 => n17266, ZN => n18155);
   U6964 : NAND2_X2 port map( A1 => n14401, A2 => n6859, ZN => n16645);
   U6966 : NAND2_X2 port map( A1 => n4361, A2 => n4366, ZN => n9042);
   U6973 : OR2_X1 port map( A1 => n3954, A2 => n19697, Z => n25714);
   U6976 : XOR2_X1 port map( A1 => n8704, A2 => n19238, Z => n19273);
   U6977 : NAND2_X2 port map( A1 => n10807, A2 => n27703, ZN => n19238);
   U6983 : INV_X2 port map( I => n22616, ZN => n24538);
   U6984 : XOR2_X1 port map( A1 => n10927, A2 => n10926, Z => n22616);
   U6986 : XOR2_X1 port map( A1 => n1912, A2 => n25023, Z => n6864);
   U6987 : XOR2_X1 port map( A1 => n25311, A2 => n21376, Z => n21378);
   U6988 : NAND2_X2 port map( A1 => n5761, A2 => n5182, ZN => n25311);
   U6989 : NAND2_X1 port map( A1 => n19805, A2 => n510, ZN => n22883);
   U6991 : NAND2_X2 port map( A1 => n28285, A2 => n8073, ZN => n2868);
   U6992 : NOR2_X1 port map( A1 => n27419, A2 => n25348, ZN => n12900);
   U6997 : XOR2_X1 port map( A1 => n27420, A2 => n21381, Z => n27419);
   U7000 : NAND2_X2 port map( A1 => n20177, A2 => n20176, ZN => n14227);
   U7001 : NAND2_X2 port map( A1 => n27993, A2 => n7418, ZN => n20177);
   U7003 : NAND2_X2 port map( A1 => n18375, A2 => n18376, ZN => n9050);
   U7005 : NAND2_X2 port map( A1 => n26899, A2 => n9738, ZN => n18375);
   U7008 : XOR2_X1 port map( A1 => n21152, A2 => n20424, Z => n21380);
   U7011 : NAND2_X2 port map( A1 => n3047, A2 => n20001, ZN => n21152);
   U7013 : NAND2_X2 port map( A1 => n21268, A2 => n5355, ZN => n21279);
   U7019 : OAI21_X2 port map( A1 => n21259, A2 => n21465, B => n14525, ZN => 
                           n21268);
   U7022 : NAND2_X2 port map( A1 => n27089, A2 => n26847, ZN => n11522);
   U7023 : INV_X2 port map( I => n13333, ZN => n20413);
   U7029 : INV_X2 port map( I => n12701, ZN => n1887);
   U7033 : OAI22_X2 port map( A1 => n4225, A2 => n23212, B1 => n20072, B2 => 
                           n20073, ZN => n12701);
   U7036 : NAND2_X2 port map( A1 => n6429, A2 => n26849, ZN => n25455);
   U7039 : AOI22_X2 port map( A1 => n19545, A2 => n19768, B1 => n28095, B2 => 
                           n19544, ZN => n26849);
   U7043 : NAND2_X1 port map( A1 => n5171, A2 => n27052, ZN => n26295);
   U7044 : NOR2_X1 port map( A1 => n12206, A2 => n27091, ZN => n20573);
   U7051 : NAND3_X2 port map( A1 => n8563, A2 => n5295, A3 => n8561, ZN => 
                           n27091);
   U7052 : XOR2_X1 port map( A1 => n7951, A2 => n8608, Z => n18245);
   U7053 : NAND2_X2 port map( A1 => n3414, A2 => n25400, ZN => n8608);
   U7054 : NAND2_X2 port map( A1 => n22387, A2 => n26850, ZN => n4021);
   U7064 : AOI22_X2 port map( A1 => n3918, A2 => n3916, B1 => n15067, B2 => 
                           n3878, ZN => n26850);
   U7065 : NAND2_X1 port map( A1 => n27784, A2 => n22458, ZN => n27675);
   U7068 : OAI22_X1 port map( A1 => n3738, A2 => n3737, B1 => n3739, B2 => 
                           n3740, ZN => n27126);
   U7070 : NAND3_X2 port map( A1 => n2787, A2 => n2786, A3 => n22955, ZN => 
                           n22087);
   U7071 : AOI22_X2 port map( A1 => n6402, A2 => n25359, B1 => n6763, B2 => 
                           n23107, ZN => n25191);
   U7076 : NOR2_X2 port map( A1 => n28008, A2 => n13794, ZN => n6402);
   U7078 : AOI22_X2 port map( A1 => n10843, A2 => n19034, B1 => n21846, B2 => 
                           n19035, ZN => n26962);
   U7083 : XOR2_X1 port map( A1 => n4627, A2 => n4625, Z => n6260);
   U7086 : OAI21_X2 port map( A1 => n7585, A2 => n19709, B => n7584, ZN => 
                           n27454);
   U7089 : XOR2_X1 port map( A1 => n6108, A2 => n15604, Z => n9904);
   U7102 : NAND2_X2 port map( A1 => n27919, A2 => n27920, ZN => n6108);
   U7108 : OAI21_X2 port map( A1 => n26851, A2 => n13932, B => n17300, ZN => 
                           n17962);
   U7109 : NAND2_X2 port map( A1 => n6199, A2 => n17511, ZN => n26851);
   U7112 : BUF_X2 port map( I => n631, Z => n26852);
   U7114 : NAND2_X2 port map( A1 => n8022, A2 => n738, ZN => n2982);
   U7115 : NAND2_X2 port map( A1 => n20491, A2 => n24383, ZN => n1728);
   U7116 : BUF_X2 port map( I => n25698, Z => n26853);
   U7117 : BUF_X2 port map( I => n15624, Z => n15307);
   U7118 : XOR2_X1 port map( A1 => n26854, A2 => n1540, Z => n6047);
   U7122 : XOR2_X1 port map( A1 => n13537, A2 => n28388, Z => n26854);
   U7125 : XOR2_X1 port map( A1 => n19312, A2 => n1307, Z => n1539);
   U7126 : OAI22_X2 port map( A1 => n9234, A2 => n9232, B1 => n9237, B2 => 
                           n28516, ZN => n19312);
   U7127 : XOR2_X1 port map( A1 => n26100, A2 => n12620, Z => n22855);
   U7129 : NAND2_X1 port map( A1 => n27311, A2 => n6882, ZN => n3319);
   U7131 : XOR2_X1 port map( A1 => n17784, A2 => n25068, Z => n23668);
   U7132 : XOR2_X1 port map( A1 => n18063, A2 => n18081, Z => n17784);
   U7133 : XOR2_X1 port map( A1 => n1713, A2 => n1712, Z => n22554);
   U7134 : NAND3_X2 port map( A1 => n26856, A2 => n22415, A3 => n17164, ZN => 
                           n6779);
   U7135 : NAND3_X2 port map( A1 => n17161, A2 => n17162, A3 => n8692, ZN => 
                           n26856);
   U7136 : XOR2_X1 port map( A1 => n26141, A2 => n920, Z => n3668);
   U7140 : NAND2_X2 port map( A1 => n23113, A2 => n25097, ZN => n26141);
   U7145 : XOR2_X1 port map( A1 => n26857, A2 => n2609, Z => n14039);
   U7149 : XOR2_X1 port map( A1 => n19303, A2 => n19358, Z => n26857);
   U7151 : INV_X2 port map( I => n19159, ZN => n14119);
   U7152 : NAND2_X2 port map( A1 => n18065, A2 => n27733, ZN => n19159);
   U7164 : XOR2_X1 port map( A1 => n26858, A2 => n11525, Z => n26414);
   U7166 : XOR2_X1 port map( A1 => n22191, A2 => n28320, Z => n26858);
   U7169 : NAND3_X1 port map( A1 => n17618, A2 => n22519, A3 => n23056, ZN => 
                           n23184);
   U7171 : NAND3_X2 port map( A1 => n5885, A2 => n22856, A3 => n18675, ZN => 
                           n27282);
   U7177 : NOR2_X2 port map( A1 => n6173, A2 => n26859, ZN => n27507);
   U7184 : NOR2_X1 port map( A1 => n18751, A2 => n6042, ZN => n26859);
   U7186 : NAND2_X2 port map( A1 => n17789, A2 => n17788, ZN => n18330);
   U7188 : NOR2_X2 port map( A1 => n27765, A2 => n6136, ZN => n17789);
   U7193 : NAND2_X2 port map( A1 => n1021, A2 => n23927, ZN => n26860);
   U7195 : AOI22_X2 port map( A1 => n12314, A2 => n20474, B1 => n25390, B2 => 
                           n25321, ZN => n25440);
   U7196 : NOR2_X2 port map( A1 => n7122, A2 => n1111, ZN => n12314);
   U7197 : XNOR2_X1 port map( A1 => n19233, A2 => n11097, ZN => n19515);
   U7198 : NAND3_X2 port map( A1 => n5903, A2 => n23467, A3 => n8694, ZN => 
                           n11097);
   U7200 : NAND2_X1 port map( A1 => n20098, A2 => n20097, ZN => n24798);
   U7201 : AND2_X1 port map( A1 => n18750, A2 => n18753, Z => n2337);
   U7205 : OAI21_X1 port map( A1 => n26568, A2 => n2323, B => n26861, ZN => n89
                           );
   U7206 : NAND2_X1 port map( A1 => n24851, A2 => n24852, ZN => n26861);
   U7207 : INV_X2 port map( I => n17384, ZN => n26862);
   U7209 : NAND2_X2 port map( A1 => n26862, A2 => n17543, ZN => n3459);
   U7210 : AOI21_X2 port map( A1 => n20185, A2 => n21759, B => n26863, ZN => 
                           n11750);
   U7213 : INV_X4 port map( I => n4537, ZN => n27487);
   U7218 : NAND3_X2 port map( A1 => n19002, A2 => n19000, A3 => n19001, ZN => 
                           n19352);
   U7219 : XOR2_X1 port map( A1 => n17970, A2 => n13793, Z => n18310);
   U7221 : NOR2_X2 port map( A1 => n2780, A2 => n2779, ZN => n17970);
   U7223 : INV_X2 port map( I => n26864, ZN => n665);
   U7226 : XOR2_X1 port map( A1 => n3585, A2 => n3586, Z => n26864);
   U7227 : XOR2_X1 port map( A1 => n21317, A2 => n13684, Z => n9597);
   U7228 : NAND2_X2 port map( A1 => n11953, A2 => n11956, ZN => n21317);
   U7229 : XOR2_X1 port map( A1 => n10352, A2 => n13092, Z => n20714);
   U7231 : NAND2_X2 port map( A1 => n27812, A2 => n6070, ZN => n10352);
   U7235 : XOR2_X1 port map( A1 => n26866, A2 => n8448, Z => n7896);
   U7236 : AOI22_X1 port map( A1 => n22216, A2 => n20128, B1 => n26944, B2 => 
                           n11372, ZN => n26866);
   U7237 : NOR3_X2 port map( A1 => n26355, A2 => n23642, A3 => n20310, ZN => 
                           n9440);
   U7240 : NAND2_X2 port map( A1 => n22897, A2 => n26867, ZN => n18147);
   U7241 : AOI22_X2 port map( A1 => n17813, A2 => n12964, B1 => n21778, B2 => 
                           n21881, ZN => n26867);
   U7242 : XOR2_X1 port map( A1 => n26868, A2 => n21075, Z => Ciphertext(85));
   U7244 : NOR3_X1 port map( A1 => n21074, A2 => n21088, A3 => n21073, ZN => 
                           n26868);
   U7245 : NOR3_X2 port map( A1 => n25591, A2 => n22096, A3 => n23618, ZN => 
                           n10388);
   U7248 : XOR2_X1 port map( A1 => n26869, A2 => n20375, Z => n15258);
   U7250 : XOR2_X1 port map( A1 => n27686, A2 => n24715, Z => n26869);
   U7255 : XOR2_X1 port map( A1 => n22191, A2 => n10456, Z => n18351);
   U7257 : NAND2_X2 port map( A1 => n33, A2 => n3711, ZN => n22191);
   U7262 : XOR2_X1 port map( A1 => n15734, A2 => n12531, Z => n3706);
   U7265 : OAI21_X2 port map( A1 => n20289, A2 => n15150, B => n10329, ZN => 
                           n15734);
   U7267 : XOR2_X1 port map( A1 => n2375, A2 => n2374, Z => n10571);
   U7268 : XOR2_X1 port map( A1 => n24848, A2 => n18319, Z => n10379);
   U7269 : NAND3_X2 port map( A1 => n24549, A2 => n25203, A3 => n23800, ZN => 
                           n27280);
   U7273 : XOR2_X1 port map( A1 => n7079, A2 => n10033, Z => n10032);
   U7280 : XOR2_X1 port map( A1 => n28018, A2 => n8441, Z => n7079);
   U7282 : OAI21_X2 port map( A1 => n4976, A2 => n26871, B => n1211, ZN => 
                           n3682);
   U7284 : INV_X2 port map( I => n27640, ZN => n26871);
   U7286 : INV_X2 port map( I => n6145, ZN => n28173);
   U7288 : XOR2_X1 port map( A1 => n18280, A2 => n25312, Z => n22069);
   U7289 : NAND2_X2 port map( A1 => n24668, A2 => n6170, ZN => n18280);
   U7296 : XOR2_X1 port map( A1 => n26874, A2 => n1294, Z => Ciphertext(30));
   U7297 : NOR2_X1 port map( A1 => n7513, A2 => n7514, ZN => n26874);
   U7299 : XOR2_X1 port map( A1 => n19234, A2 => n26469, Z => n25617);
   U7300 : XOR2_X1 port map( A1 => n3900, A2 => n2747, Z => n649);
   U7303 : NAND2_X2 port map( A1 => n26875, A2 => n18948, ZN => n6132);
   U7310 : OAI22_X2 port map( A1 => n27506, A2 => n2070, B1 => n19006, B2 => 
                           n18947, ZN => n26875);
   U7313 : AOI22_X2 port map( A1 => n25417, A2 => n15461, B1 => n20259, B2 => 
                           n26898, ZN => n9760);
   U7314 : NAND2_X2 port map( A1 => n14823, A2 => n26130, ZN => n26898);
   U7318 : NAND2_X1 port map( A1 => n26557, A2 => n13234, ZN => n23883);
   U7319 : NAND3_X2 port map( A1 => n8766, A2 => n8765, A3 => n8764, ZN => 
                           n13234);
   U7320 : XOR2_X1 port map( A1 => n26967, A2 => n11723, Z => n20365);
   U7322 : NAND2_X2 port map( A1 => n7934, A2 => n7932, ZN => n12531);
   U7323 : INV_X4 port map( I => n26876, ZN => n25959);
   U7325 : AND3_X2 port map( A1 => n19656, A2 => n24600, A3 => n9441, Z => 
                           n26876);
   U7327 : INV_X1 port map( I => n8464, ZN => n26877);
   U7328 : NOR2_X1 port map( A1 => n26877, A2 => n19499, ZN => n6655);
   U7330 : NAND2_X1 port map( A1 => n8106, A2 => n3335, ZN => n27540);
   U7331 : NOR2_X2 port map( A1 => n26716, A2 => n27545, ZN => n25761);
   U7332 : XOR2_X1 port map( A1 => n13816, A2 => n13818, Z => n18457);
   U7333 : INV_X1 port map( I => n26878, ZN => n15614);
   U7336 : NAND2_X1 port map( A1 => n16419, A2 => n3914, ZN => n26878);
   U7337 : NAND3_X2 port map( A1 => n2281, A2 => n7483, A3 => n2282, ZN => 
                           n16419);
   U7340 : AOI21_X1 port map( A1 => n999, A2 => n24019, B => n998, ZN => n4669)
                           ;
   U7343 : NOR2_X1 port map( A1 => n24720, A2 => n26898, ZN => n26901);
   U7344 : NAND2_X2 port map( A1 => n5113, A2 => n5112, ZN => n988);
   U7345 : NAND2_X2 port map( A1 => n18761, A2 => n1000, ZN => n5112);
   U7353 : BUF_X2 port map( I => n18609, Z => n26880);
   U7354 : OAI22_X2 port map( A1 => n21383, A2 => n21590, B1 => n25696, B2 => 
                           n24621, ZN => n21406);
   U7356 : NAND2_X2 port map( A1 => n6310, A2 => n26881, ZN => n12584);
   U7358 : NAND3_X2 port map( A1 => n6755, A2 => n25828, A3 => n10708, ZN => 
                           n26881);
   U7360 : NOR2_X2 port map( A1 => n940, A2 => n8271, ZN => n10674);
   U7363 : BUF_X2 port map( I => n21548, Z => n26882);
   U7367 : NAND2_X2 port map( A1 => n2079, A2 => n28339, ZN => n2231);
   U7368 : AOI22_X2 port map( A1 => n3918, A2 => n15067, B1 => n810, B2 => 
                           n3878, ZN => n28339);
   U7369 : NAND2_X2 port map( A1 => n26883, A2 => n19617, ZN => n20316);
   U7371 : NAND2_X1 port map( A1 => n13353, A2 => n27542, ZN => n26883);
   U7374 : XOR2_X1 port map( A1 => n19273, A2 => n19412, Z => n19357);
   U7375 : INV_X1 port map( I => n26984, ZN => n13019);
   U7376 : NAND2_X2 port map( A1 => n10827, A2 => n9790, ZN => n9116);
   U7378 : INV_X4 port map( I => n8330, ZN => n3918);
   U7383 : XOR2_X1 port map( A1 => n6867, A2 => n18205, Z => n13064);
   U7384 : NAND2_X2 port map( A1 => n6847, A2 => n6848, ZN => n6867);
   U7389 : NOR2_X1 port map( A1 => n12186, A2 => n21000, ZN => n11323);
   U7394 : NAND3_X2 port map( A1 => n27977, A2 => n20984, A3 => n24280, ZN => 
                           n12186);
   U7396 : OAI21_X2 port map( A1 => n21919, A2 => n23017, B => n27938, ZN => 
                           n8913);
   U7400 : OAI21_X2 port map( A1 => n26678, A2 => n26885, B => n14244, ZN => 
                           n6967);
   U7402 : AOI22_X1 port map( A1 => n27593, A2 => n27257, B1 => n14319, B2 => 
                           n4247, ZN => n194);
   U7405 : XOR2_X1 port map( A1 => n15174, A2 => n18095, Z => n2129);
   U7406 : NAND2_X1 port map( A1 => n19868, A2 => n27719, ZN => n25209);
   U7408 : NAND2_X2 port map( A1 => n11143, A2 => n27599, ZN => n17026);
   U7410 : NAND2_X2 port map( A1 => n5757, A2 => n11144, ZN => n11143);
   U7411 : INV_X4 port map( I => n27074, ZN => n17956);
   U7412 : NAND2_X2 port map( A1 => n17959, A2 => n27074, ZN => n27806);
   U7413 : NAND2_X2 port map( A1 => n27355, A2 => n8804, ZN => n26886);
   U7417 : INV_X4 port map( I => n23772, ZN => n817);
   U7419 : NOR2_X2 port map( A1 => n13566, A2 => n13567, ZN => n13421);
   U7420 : NAND3_X2 port map( A1 => n26500, A2 => n3459, A3 => n23600, ZN => 
                           n13566);
   U7424 : NOR2_X2 port map( A1 => n27290, A2 => n2097, ZN => n14583);
   U7425 : AOI21_X1 port map( A1 => n26521, A2 => n23371, B => n12066, ZN => 
                           n2097);
   U7427 : NAND2_X2 port map( A1 => n27004, A2 => n23243, ZN => n4827);
   U7430 : NOR2_X2 port map( A1 => n3438, A2 => n26887, ZN => n25854);
   U7435 : NAND2_X2 port map( A1 => n5697, A2 => n5693, ZN => n26887);
   U7446 : AOI22_X2 port map( A1 => n8756, A2 => n28199, B1 => n13775, B2 => 
                           n19774, ZN => n20324);
   U7458 : OAI21_X2 port map( A1 => n8754, A2 => n14393, B => n9896, ZN => 
                           n8756);
   U7462 : XOR2_X1 port map( A1 => n12437, A2 => n7887, Z => n27956);
   U7463 : XOR2_X1 port map( A1 => n24152, A2 => n26888, Z => n7870);
   U7465 : XOR2_X1 port map( A1 => n20724, A2 => n13965, Z => n26888);
   U7467 : XOR2_X1 port map( A1 => n13537, A2 => n19255, Z => n19258);
   U7468 : XOR2_X1 port map( A1 => n10038, A2 => n19462, Z => n13537);
   U7470 : XOR2_X1 port map( A1 => n26889, A2 => n14489, Z => Ciphertext(190));
   U7474 : NAND3_X2 port map( A1 => n11168, A2 => n25562, A3 => n14060, ZN => 
                           n26889);
   U7475 : XOR2_X1 port map( A1 => n17102, A2 => n17047, Z => n8685);
   U7477 : XOR2_X1 port map( A1 => n10670, A2 => n21926, Z => n1385);
   U7478 : XOR2_X1 port map( A1 => n5520, A2 => n12759, Z => n10670);
   U7484 : NAND2_X1 port map( A1 => n27553, A2 => n11267, ZN => n3267);
   U7485 : NOR3_X1 port map( A1 => n26891, A2 => n23253, A3 => n12364, ZN => 
                           n26890);
   U7499 : NAND3_X2 port map( A1 => n23209, A2 => n23210, A3 => n26027, ZN => 
                           n2252);
   U7502 : NAND3_X1 port map( A1 => n9654, A2 => n21126, A3 => n26952, ZN => 
                           n25256);
   U7509 : NAND2_X1 port map( A1 => n21344, A2 => n27439, ZN => n2453);
   U7515 : XOR2_X1 port map( A1 => n21320, A2 => n21438, Z => n10328);
   U7516 : OAI21_X2 port map( A1 => n6926, A2 => n6925, B => n26892, ZN => 
                           n6921);
   U7518 : NAND2_X2 port map( A1 => n6923, A2 => n6924, ZN => n26892);
   U7520 : NAND2_X2 port map( A1 => n11652, A2 => n26893, ZN => n10378);
   U7522 : NAND2_X1 port map( A1 => n22956, A2 => n23043, ZN => n26893);
   U7529 : NAND2_X2 port map( A1 => n12005, A2 => n20210, ZN => n27882);
   U7530 : XOR2_X1 port map( A1 => n8374, A2 => n19324, Z => n8441);
   U7531 : NOR3_X2 port map( A1 => n25042, A2 => n1704, A3 => n21999, ZN => 
                           n8374);
   U7536 : AOI22_X2 port map( A1 => n16305, A2 => n1362, B1 => n3773, B2 => 
                           n26895, ZN => n7900);
   U7540 : NAND3_X1 port map( A1 => n24072, A2 => n5811, A3 => n24071, ZN => 
                           n27807);
   U7541 : NOR2_X1 port map( A1 => n21713, A2 => n15513, ZN => n26908);
   U7544 : OAI21_X1 port map( A1 => n10388, A2 => n10389, B => n1284, ZN => 
                           n28386);
   U7545 : XOR2_X1 port map( A1 => n26896, A2 => n21650, Z => Ciphertext(169));
   U7556 : OAI22_X1 port map( A1 => n10124, A2 => n21660, B1 => n22743, B2 => 
                           n21655, ZN => n26896);
   U7561 : NAND3_X2 port map( A1 => n10924, A2 => n8716, A3 => n3960, ZN => 
                           n24075);
   U7562 : OR2_X1 port map( A1 => n12494, A2 => n26897, Z => n24645);
   U7566 : BUF_X2 port map( I => n879, Z => n26899);
   U7571 : OAI21_X2 port map( A1 => n26901, A2 => n26900, B => n2973, ZN => 
                           n15226);
   U7573 : NAND2_X2 port map( A1 => n2971, A2 => n15461, ZN => n26900);
   U7577 : OAI21_X2 port map( A1 => n7153, A2 => n11129, B => n11126, ZN => 
                           n13478);
   U7579 : INV_X1 port map( I => n784, ZN => n27785);
   U7580 : OR2_X1 port map( A1 => n784, A2 => n18491, Z => n27784);
   U7582 : NOR2_X2 port map( A1 => n16113, A2 => n1881, ZN => n6713);
   U7583 : AOI21_X2 port map( A1 => n23419, A2 => n10636, B => n6909, ZN => 
                           n6355);
   U7584 : NOR2_X2 port map( A1 => n10595, A2 => n6354, ZN => n6909);
   U7586 : XOR2_X1 port map( A1 => n19083, A2 => n19084, Z => n19649);
   U7587 : XOR2_X1 port map( A1 => n10670, A2 => n21368, Z => n5594);
   U7593 : XOR2_X1 port map( A1 => n21157, A2 => n21158, Z => n21368);
   U7595 : AOI21_X2 port map( A1 => n14896, A2 => n867, B => n26902, ZN => 
                           n20087);
   U7597 : AOI21_X2 port map( A1 => n8887, A2 => n14895, B => n867, ZN => 
                           n26902);
   U7598 : NAND3_X2 port map( A1 => n26903, A2 => n7072, A3 => n18982, ZN => 
                           n23746);
   U7607 : INV_X2 port map( I => n2232, ZN => n25753);
   U7610 : NAND2_X2 port map( A1 => n27042, A2 => n23805, ZN => n2232);
   U7619 : NAND2_X2 port map( A1 => n6487, A2 => n14237, ZN => n6489);
   U7621 : NAND2_X2 port map( A1 => n23291, A2 => n28171, ZN => n6487);
   U7623 : OAI22_X1 port map( A1 => n26092, A2 => n9894, B1 => n1065, B2 => 
                           n6281, ZN => n2407);
   U7630 : OAI21_X2 port map( A1 => n26907, A2 => n26908, B => n12171, ZN => 
                           n9894);
   U7635 : NAND2_X2 port map( A1 => n18761, A2 => n27829, ZN => n27805);
   U7639 : XOR2_X1 port map( A1 => n28312, A2 => n26904, Z => n13170);
   U7640 : XOR2_X1 port map( A1 => n20322, A2 => n20539, Z => n26904);
   U7648 : XOR2_X1 port map( A1 => n26905, A2 => n21557, Z => Ciphertext(152));
   U7650 : AOI22_X1 port map( A1 => n21555, A2 => n21568, B1 => n21556, B2 => 
                           n22789, ZN => n26905);
   U7658 : OAI21_X2 port map( A1 => n2287, A2 => n1464, B => n26906, ZN => 
                           n18097);
   U7660 : NAND3_X2 port map( A1 => n1022, A2 => n9480, A3 => n23645, ZN => 
                           n26906);
   U7662 : AND2_X1 port map( A1 => n17302, A2 => n17193, Z => n24695);
   U7669 : OAI22_X2 port map( A1 => n450, A2 => n5986, B1 => n821, B2 => n18475
                           , ZN => n6913);
   U7670 : NAND2_X2 port map( A1 => n23124, A2 => n21664, ZN => n26907);
   U7672 : NAND2_X2 port map( A1 => n15582, A2 => n26909, ZN => n20535);
   U7675 : NAND2_X2 port map( A1 => n20569, A2 => n22234, ZN => n20436);
   U7676 : NAND2_X2 port map( A1 => n9092, A2 => n25527, ZN => n20569);
   U7678 : XOR2_X1 port map( A1 => n13180, A2 => n26910, Z => n15512);
   U7685 : XOR2_X1 port map( A1 => n13179, A2 => n13178, Z => n26910);
   U7686 : XOR2_X1 port map( A1 => n26911, A2 => n12956, Z => n22718);
   U7688 : XOR2_X1 port map( A1 => n20517, A2 => n20518, Z => n26911);
   U7691 : NAND2_X2 port map( A1 => n7485, A2 => n7484, ZN => n27647);
   U7692 : NAND3_X2 port map( A1 => n26912, A2 => n10759, A3 => n26235, ZN => 
                           n2484);
   U7696 : NAND2_X1 port map( A1 => n2487, A2 => n13455, ZN => n26912);
   U7698 : AOI21_X2 port map( A1 => n1119, A2 => n20110, B => n978, ZN => 
                           n20113);
   U7699 : NAND2_X2 port map( A1 => n20152, A2 => n11519, ZN => n27144);
   U7700 : XOR2_X1 port map( A1 => n25892, A2 => n17970, Z => n27480);
   U7704 : OAI22_X2 port map( A1 => n4972, A2 => n24570, B1 => n4973, B2 => 
                           n4974, ZN => n25892);
   U7705 : AOI22_X1 port map( A1 => n6353, A2 => n7319, B1 => n20610, B2 => 
                           n5195, ZN => n3418);
   U7706 : AOI21_X2 port map( A1 => n8435, A2 => n1222, B => n27287, ZN => 
                           n9965);
   U7707 : XOR2_X1 port map( A1 => n27767, A2 => n21157, Z => n20422);
   U7708 : NAND2_X2 port map( A1 => n6423, A2 => n6422, ZN => n21157);
   U7716 : XOR2_X1 port map( A1 => n13958, A2 => n13960, Z => n18443);
   U7719 : XOR2_X1 port map( A1 => n10072, A2 => n19319, Z => n10069);
   U7721 : NAND2_X1 port map( A1 => n15008, A2 => n18699, ZN => n27515);
   U7724 : BUF_X2 port map( I => n6066, Z => n26913);
   U7725 : NOR2_X2 port map( A1 => n17950, A2 => n17953, ZN => n11488);
   U7726 : NAND2_X2 port map( A1 => n15393, A2 => n15395, ZN => n17953);
   U7728 : OR2_X1 port map( A1 => n8311, A2 => n26914, Z => n5813);
   U7732 : XOR2_X1 port map( A1 => n2595, A2 => n12380, Z => n12655);
   U7734 : NOR2_X2 port map( A1 => n26915, A2 => n27119, ZN => n21561);
   U7735 : NAND2_X2 port map( A1 => n27118, A2 => n27117, ZN => n26915);
   U7737 : NOR2_X2 port map( A1 => n19876, A2 => n23748, ZN => n11836);
   U7738 : XOR2_X1 port map( A1 => n7562, A2 => n14868, Z => n7563);
   U7739 : AOI21_X2 port map( A1 => n26916, A2 => n2385, B => n6041, ZN => 
                           n2382);
   U7740 : OR2_X1 port map( A1 => n27440, A2 => n6042, Z => n26916);
   U7742 : NOR2_X2 port map( A1 => n17436, A2 => n24513, ZN => n8275);
   U7744 : OAI21_X2 port map( A1 => n24185, A2 => n6606, B => n24547, ZN => 
                           n9918);
   U7746 : XOR2_X1 port map( A1 => n2655, A2 => n14604, Z => n8748);
   U7748 : NAND2_X2 port map( A1 => n2513, A2 => n2511, ZN => n2655);
   U7753 : NAND2_X1 port map( A1 => n26919, A2 => n26918, ZN => n8738);
   U7756 : NAND2_X1 port map( A1 => n26921, A2 => n9946, ZN => n26919);
   U7758 : INV_X2 port map( I => n25104, ZN => n26920);
   U7765 : NAND2_X1 port map( A1 => n24524, A2 => n2647, ZN => n26921);
   U7767 : BUF_X2 port map( I => n24107, Z => n26922);
   U7770 : NAND3_X2 port map( A1 => n26925, A2 => n19998, A3 => n19996, ZN => 
                           n1715);
   U7772 : OAI21_X2 port map( A1 => n23073, A2 => n21882, B => n334, ZN => 
                           n26925);
   U7773 : NOR2_X2 port map( A1 => n4040, A2 => n26926, ZN => n26312);
   U7774 : AOI22_X1 port map( A1 => n17573, A2 => n12236, B1 => n3533, B2 => 
                           n17570, ZN => n26926);
   U7778 : NAND3_X2 port map( A1 => n8280, A2 => n21861, A3 => n14054, ZN => 
                           n8293);
   U7779 : NAND2_X2 port map( A1 => n26927, A2 => n4155, ZN => n4383);
   U7780 : NOR2_X1 port map( A1 => n23620, A2 => n23621, ZN => n26927);
   U7781 : INV_X2 port map( I => n14975, ZN => n860);
   U7784 : NAND2_X2 port map( A1 => n15250, A2 => n19804, ZN => n14975);
   U7786 : NAND3_X2 port map( A1 => n15516, A2 => n13917, A3 => n15517, ZN => 
                           n13918);
   U7787 : XOR2_X1 port map( A1 => n26928, A2 => n19385, Z => n18438);
   U7788 : XOR2_X1 port map( A1 => n19330, A2 => n982, Z => n26928);
   U7789 : XNOR2_X1 port map( A1 => n17077, A2 => n8274, ZN => n27103);
   U7790 : NOR2_X2 port map( A1 => n4832, A2 => n167, ZN => n11270);
   U7796 : XOR2_X1 port map( A1 => n26929, A2 => n14597, Z => Ciphertext(94));
   U7797 : NAND3_X1 port map( A1 => n13033, A2 => n13030, A3 => n13031, ZN => 
                           n26929);
   U7798 : NAND2_X1 port map( A1 => n26942, A2 => n1072, ZN => n10630);
   U7800 : INV_X2 port map( I => n26930, ZN => n27749);
   U7801 : NOR2_X2 port map( A1 => n26931, A2 => n4488, ZN => n4487);
   U7803 : NOR2_X2 port map( A1 => n9363, A2 => n16329, ZN => n26931);
   U7809 : INV_X2 port map( I => n26932, ZN => n1403);
   U7810 : NAND2_X2 port map( A1 => n3768, A2 => n3767, ZN => n26932);
   U7813 : OAI21_X2 port map( A1 => n26936, A2 => n12159, B => n24146, ZN => 
                           n8166);
   U7814 : NOR2_X2 port map( A1 => n28443, A2 => n26126, ZN => n22815);
   U7820 : NAND2_X2 port map( A1 => n12033, A2 => n26933, ZN => n15334);
   U7822 : NAND2_X2 port map( A1 => n20245, A2 => n3891, ZN => n35);
   U7826 : XOR2_X1 port map( A1 => n18300, A2 => n18299, Z => n10055);
   U7827 : XOR2_X1 port map( A1 => n28263, A2 => n27624, Z => n2019);
   U7828 : XOR2_X1 port map( A1 => n26934, A2 => n1306, Z => Ciphertext(92));
   U7834 : NAND2_X1 port map( A1 => n26015, A2 => n8543, ZN => n26934);
   U7836 : XOR2_X1 port map( A1 => n27692, A2 => n27691, Z => n22122);
   U7838 : OAI21_X2 port map( A1 => n23471, A2 => n24821, B => n26935, ZN => 
                           n17549);
   U7839 : OAI21_X2 port map( A1 => n17540, A2 => n11857, B => n3980, ZN => 
                           n26935);
   U7841 : NOR2_X2 port map( A1 => n113, A2 => n813, ZN => n26936);
   U7842 : XOR2_X1 port map( A1 => n10378, A2 => n14621, Z => n12321);
   U7848 : XOR2_X1 port map( A1 => n26937, A2 => n23827, Z => n19916);
   U7851 : XOR2_X1 port map( A1 => n19415, A2 => n28067, Z => n26937);
   U7853 : AOI22_X2 port map( A1 => n7524, A2 => n9593, B1 => n17561, B2 => 
                           n17562, ZN => n4070);
   U7858 : OAI22_X2 port map( A1 => n15077, A2 => n17561, B1 => n14061, B2 => 
                           n17559, ZN => n7524);
   U7861 : NAND3_X2 port map( A1 => n26938, A2 => n6092, A3 => n6091, ZN => 
                           n21289);
   U7862 : NAND3_X2 port map( A1 => n26011, A2 => n26010, A3 => n6095, ZN => 
                           n26938);
   U7864 : OR2_X1 port map( A1 => n20154, A2 => n958, Z => n677);
   U7865 : XOR2_X1 port map( A1 => n11100, A2 => n20564, Z => n7467);
   U7867 : XOR2_X1 port map( A1 => n8819, A2 => n17133, Z => n13661);
   U7870 : NOR2_X2 port map( A1 => n14270, A2 => n7806, ZN => n8819);
   U7871 : BUF_X2 port map( I => n23391, Z => n26939);
   U7879 : NAND2_X2 port map( A1 => n18933, A2 => n8683, ZN => n19014);
   U7886 : NAND2_X2 port map( A1 => n26975, A2 => n13954, ZN => n16531);
   U7888 : BUF_X2 port map( I => n21695, Z => n22828);
   U7903 : XOR2_X1 port map( A1 => n19403, A2 => n26940, Z => n23109);
   U7905 : XOR2_X1 port map( A1 => n19173, A2 => n14971, Z => n26940);
   U7907 : XOR2_X1 port map( A1 => n6615, A2 => n6614, Z => n9618);
   U7908 : AOI21_X2 port map( A1 => n16608, A2 => n16605, B => n26941, ZN => 
                           n12275);
   U7909 : OAI22_X2 port map( A1 => n703, A2 => n4059, B1 => n16605, B2 => 
                           n16508, ZN => n26941);
   U7910 : NAND2_X2 port map( A1 => n6998, A2 => n14513, ZN => n13429);
   U7912 : NAND2_X2 port map( A1 => n24145, A2 => n24144, ZN => n6998);
   U7915 : MUX2_X1 port map( I0 => n20956, I1 => n20957, S => n23088, Z => 
                           n20960);
   U7916 : INV_X1 port map( I => n477, ZN => n26942);
   U7918 : NOR2_X2 port map( A1 => n20925, A2 => n20924, ZN => n477);
   U7919 : OR2_X2 port map( A1 => n10497, A2 => n26754, Z => n4797);
   U7920 : XOR2_X1 port map( A1 => n11578, A2 => n20546, Z => n11752);
   U7922 : XOR2_X1 port map( A1 => n26634, A2 => n3506, Z => n11578);
   U7924 : BUF_X2 port map( I => n13752, Z => n27863);
   U7927 : AOI21_X2 port map( A1 => n8989, A2 => n28382, B => n28381, ZN => 
                           n26943);
   U7931 : NAND2_X2 port map( A1 => n26945, A2 => n25965, ZN => n12995);
   U7933 : OAI21_X2 port map( A1 => n12492, A2 => n12491, B => n12659, ZN => 
                           n26945);
   U7934 : NAND2_X2 port map( A1 => n26947, A2 => n26946, ZN => n23686);
   U7935 : NAND2_X2 port map( A1 => n6182, A2 => n21659, ZN => n2766);
   U7937 : XOR2_X1 port map( A1 => n19533, A2 => n19464, Z => n4203);
   U7952 : NAND2_X2 port map( A1 => n22093, A2 => n2676, ZN => n19533);
   U7954 : XOR2_X1 port map( A1 => n9058, A2 => n9124, Z => n23687);
   U7960 : OAI21_X1 port map( A1 => n7698, A2 => n13234, B => n20670, ZN => 
                           n10409);
   U7963 : XOR2_X1 port map( A1 => n27285, A2 => n10084, Z => n5086);
   U7972 : XOR2_X1 port map( A1 => n5082, A2 => n21376, Z => n10084);
   U7977 : XOR2_X1 port map( A1 => n23086, A2 => n15052, Z => n19397);
   U7981 : XOR2_X1 port map( A1 => n7215, A2 => n10071, Z => n19291);
   U7983 : AOI22_X1 port map( A1 => n15435, A2 => n12521, B1 => n22643, B2 => 
                           n15429, ZN => n26949);
   U7985 : NAND2_X2 port map( A1 => n26950, A2 => n3521, ZN => n3479);
   U7986 : XOR2_X1 port map( A1 => n12100, A2 => n19421, Z => n28318);
   U7991 : NOR2_X2 port map( A1 => n5038, A2 => n2108, ZN => n19421);
   U7998 : AOI22_X2 port map( A1 => n13835, A2 => n1101, B1 => n20132, B2 => 
                           n28408, ZN => n3220);
   U8000 : NAND2_X2 port map( A1 => n12656, A2 => n25827, ZN => n27417);
   U8002 : NOR2_X2 port map( A1 => n12659, A2 => n11583, ZN => n12658);
   U8004 : XOR2_X1 port map( A1 => n13811, A2 => n26951, Z => n9641);
   U8005 : XOR2_X1 port map( A1 => n28529, A2 => n28530, Z => n26951);
   U8015 : OR2_X2 port map( A1 => n8032, A2 => n14221, Z => n20173);
   U8019 : XOR2_X1 port map( A1 => n19457, A2 => n26725, Z => n5174);
   U8025 : XOR2_X1 port map( A1 => n19302, A2 => n19274, Z => n19457);
   U8027 : NAND2_X2 port map( A1 => n23602, A2 => n24616, ZN => n5974);
   U8030 : AOI22_X2 port map( A1 => n23819, A2 => n6825, B1 => n8237, B2 => 
                           n6330, ZN => n23602);
   U8034 : NAND2_X2 port map( A1 => n4057, A2 => n21124, ZN => n9654);
   U8044 : AOI21_X2 port map( A1 => n8380, A2 => n17431, B => n26953, ZN => 
                           n8379);
   U8049 : NOR3_X2 port map( A1 => n8263, A2 => n23105, A3 => n17519, ZN => 
                           n26953);
   U8050 : XOR2_X1 port map( A1 => n24275, A2 => n28465, Z => n19326);
   U8056 : XOR2_X1 port map( A1 => n12411, A2 => n4383, Z => n2319);
   U8063 : XOR2_X1 port map( A1 => n15488, A2 => n15487, Z => n1679);
   U8073 : XOR2_X1 port map( A1 => n1397, A2 => n18066, Z => n15487);
   U8075 : OAI22_X2 port map( A1 => n25289, A2 => n5081, B1 => n13481, B2 => 
                           n16732, ZN => n27976);
   U8076 : NAND2_X2 port map( A1 => n5725, A2 => n26280, ZN => n11413);
   U8078 : XOR2_X1 port map( A1 => n26954, A2 => n19270, Z => Ciphertext(154));
   U8083 : NAND2_X2 port map( A1 => n24221, A2 => n26955, ZN => n18217);
   U8087 : OAI21_X2 port map( A1 => n14025, A2 => n8071, B => n23856, ZN => 
                           n26955);
   U8092 : INV_X2 port map( I => n3016, ZN => n25151);
   U8093 : NOR2_X2 port map( A1 => n24147, A2 => n20156, ZN => n3016);
   U8094 : AOI21_X2 port map( A1 => n28218, A2 => n17172, B => n5204, ZN => 
                           n9419);
   U8100 : NAND2_X2 port map( A1 => n11576, A2 => n23905, ZN => n1418);
   U8103 : NOR2_X2 port map( A1 => n19908, A2 => n27303, ZN => n27721);
   U8105 : INV_X2 port map( I => n26956, ZN => n24458);
   U8106 : XOR2_X1 port map( A1 => n4945, A2 => n4947, Z => n26956);
   U8107 : XOR2_X1 port map( A1 => n15007, A2 => n26957, Z => n27141);
   U8108 : XOR2_X1 port map( A1 => n21316, A2 => n26958, Z => n26957);
   U8114 : NAND2_X1 port map( A1 => n19126, A2 => n2617, ZN => n18576);
   U8116 : NAND2_X2 port map( A1 => n25162, A2 => n26281, ZN => n19126);
   U8124 : BUF_X4 port map( I => n5961, Z => n100);
   U8125 : OAI21_X2 port map( A1 => n3547, A2 => n9142, B => n26959, ZN => 
                           n8000);
   U8126 : AOI22_X2 port map( A1 => n24507, A2 => n3544, B1 => n5353, B2 => 
                           n3545, ZN => n26959);
   U8136 : BUF_X2 port map( I => n23146, Z => n26960);
   U8137 : AOI21_X2 port map( A1 => n26994, A2 => n27443, B => n9094, ZN => 
                           n26961);
   U8141 : NOR2_X2 port map( A1 => n11140, A2 => n26674, ZN => n27300);
   U8142 : NAND2_X2 port map( A1 => n22732, A2 => n22789, ZN => n21566);
   U8147 : NAND2_X2 port map( A1 => n27840, A2 => n26964, ZN => n4265);
   U8149 : NAND3_X2 port map( A1 => n22557, A2 => n10872, A3 => n22621, ZN => 
                           n26964);
   U8155 : NAND2_X1 port map( A1 => n27284, A2 => n22237, ZN => n24970);
   U8161 : NOR2_X2 port map( A1 => n26966, A2 => n26965, ZN => n25241);
   U8163 : NAND2_X2 port map( A1 => n28308, A2 => n22789, ZN => n26965);
   U8165 : INV_X1 port map( I => n21565, ZN => n26966);
   U8171 : XOR2_X1 port map( A1 => n21201, A2 => n7813, Z => n26967);
   U8172 : NAND3_X2 port map( A1 => n1799, A2 => n28391, A3 => n630, ZN => 
                           n1869);
   U8173 : XOR2_X1 port map( A1 => n6123, A2 => n18063, Z => n18167);
   U8176 : NAND2_X2 port map( A1 => n23833, A2 => n5828, ZN => n6123);
   U8180 : XOR2_X1 port map( A1 => n1197, A2 => n18249, Z => n18084);
   U8183 : NAND2_X2 port map( A1 => n27605, A2 => n24665, ZN => n1197);
   U8184 : NAND2_X2 port map( A1 => n7421, A2 => n4667, ZN => n21029);
   U8188 : NOR2_X2 port map( A1 => n26968, A2 => n4005, ZN => n16784);
   U8192 : NAND2_X2 port map( A1 => n26357, A2 => n21833, ZN => n26968);
   U8195 : NAND2_X1 port map( A1 => n25524, A2 => n17796, ZN => n27605);
   U8197 : XOR2_X1 port map( A1 => n11989, A2 => n5494, Z => n19651);
   U8201 : AOI22_X2 port map( A1 => n20890, A2 => n26978, B1 => n27689, B2 => 
                           n4742, ZN => n20893);
   U8203 : XOR2_X1 port map( A1 => n5597, A2 => n5596, Z => n5595);
   U8205 : NAND2_X2 port map( A1 => n27198, A2 => n2772, ZN => n5597);
   U8210 : INV_X2 port map( I => n20312, ZN => n26970);
   U8214 : NAND3_X2 port map( A1 => n11517, A2 => n2444, A3 => n26971, ZN => 
                           n20183);
   U8217 : OAI21_X2 port map( A1 => n24855, A2 => n24854, B => n1119, ZN => 
                           n26971);
   U8223 : XOR2_X1 port map( A1 => n23314, A2 => n22778, Z => n15647);
   U8224 : NAND2_X2 port map( A1 => n23141, A2 => n2834, ZN => n23314);
   U8227 : NAND2_X1 port map( A1 => n6622, A2 => n6621, ZN => n6620);
   U8234 : NAND2_X2 port map( A1 => n5353, A2 => n27959, ZN => n17517);
   U8235 : NAND2_X2 port map( A1 => n10264, A2 => n26972, ZN => n24275);
   U8244 : AOI22_X2 port map( A1 => n19141, A2 => n10474, B1 => n25664, B2 => 
                           n13171, ZN => n26972);
   U8246 : OAI21_X2 port map( A1 => n24539, A2 => n1085, B => n26973, ZN => 
                           n5756);
   U8259 : AOI21_X2 port map( A1 => n5753, A2 => n24539, B => n24078, ZN => 
                           n26973);
   U8260 : NAND2_X1 port map( A1 => n14737, A2 => n26491, ZN => n17782);
   U8263 : NAND2_X2 port map( A1 => n11589, A2 => n28036, ZN => n14737);
   U8265 : AOI21_X1 port map( A1 => n12235, A2 => n28165, B => n20667, ZN => 
                           n20669);
   U8269 : AOI22_X2 port map( A1 => n16114, A2 => n9526, B1 => n3262, B2 => 
                           n15921, ZN => n26975);
   U8270 : NAND2_X2 port map( A1 => n26976, A2 => n28368, ZN => n4179);
   U8280 : OAI21_X2 port map( A1 => n2258, A2 => n4542, B => n2257, ZN => 
                           n18921);
   U8295 : NAND2_X2 port map( A1 => n10217, A2 => n6756, ZN => n21228);
   U8307 : NAND2_X2 port map( A1 => n28228, A2 => n28427, ZN => n10217);
   U8312 : XOR2_X1 port map( A1 => n3806, A2 => n26977, Z => n21271);
   U8319 : XOR2_X1 port map( A1 => n14882, A2 => n20481, Z => n26977);
   U8325 : INV_X4 port map( I => n24323, ZN => n27959);
   U8349 : NAND2_X2 port map( A1 => n28205, A2 => n25882, ZN => n3846);
   U8384 : AOI22_X2 port map( A1 => n17205, A2 => n897, B1 => n17409, B2 => 
                           n17206, ZN => n25882);
   U8389 : OAI21_X2 port map( A1 => n3848, A2 => n14357, B => n3847, ZN => 
                           n28205);
   U8399 : BUF_X2 port map( I => n21024, Z => n26978);
   U8401 : NAND2_X2 port map( A1 => n26979, A2 => n1665, ZN => n8820);
   U8403 : NAND2_X2 port map( A1 => n24770, A2 => n16410, ZN => n26979);
   U8406 : XOR2_X1 port map( A1 => n18120, A2 => n18317, Z => n13860);
   U8408 : NAND2_X2 port map( A1 => n15563, A2 => n17805, ZN => n18317);
   U8409 : NAND3_X2 port map( A1 => n13453, A2 => n22291, A3 => n28188, ZN => 
                           n19980);
   U8410 : NAND2_X2 port map( A1 => n986, A2 => n12583, ZN => n23643);
   U8412 : NAND2_X1 port map( A1 => n26980, A2 => n1652, ZN => n27795);
   U8413 : NAND2_X1 port map( A1 => n25252, A2 => n7212, ZN => n26980);
   U8416 : INV_X2 port map( I => n18918, ZN => n18919);
   U8420 : NAND2_X2 port map( A1 => n12195, A2 => n3932, ZN => n18918);
   U8427 : AOI22_X2 port map( A1 => n26981, A2 => n23138, B1 => n19018, B2 => 
                           n19017, ZN => n19536);
   U8431 : XOR2_X1 port map( A1 => n14753, A2 => n16991, Z => n17073);
   U8433 : NAND2_X2 port map( A1 => n27015, A2 => n25425, ZN => n16991);
   U8434 : NAND2_X2 port map( A1 => n9692, A2 => n9694, ZN => n21536);
   U8436 : XOR2_X1 port map( A1 => n21239, A2 => n20361, Z => n9933);
   U8442 : BUF_X2 port map( I => n12507, Z => n26982);
   U8445 : NOR2_X2 port map( A1 => n14193, A2 => n968, ZN => n19544);
   U8447 : INV_X2 port map( I => n3725, ZN => n937);
   U8448 : XOR2_X1 port map( A1 => n5275, A2 => n25092, Z => n25955);
   U8453 : NAND2_X1 port map( A1 => n7950, A2 => n26989, ZN => n14945);
   U8454 : XOR2_X1 port map( A1 => n26983, A2 => n3394, Z => n3353);
   U8455 : XOR2_X1 port map( A1 => n8072, A2 => n20512, Z => n26983);
   U8457 : XOR2_X1 port map( A1 => n19261, A2 => n19527, Z => n19549);
   U8460 : NAND2_X2 port map( A1 => n27917, A2 => n22640, ZN => n19527);
   U8461 : NAND2_X2 port map( A1 => n20329, A2 => n20415, ZN => n26551);
   U8463 : NAND2_X1 port map( A1 => n4111, A2 => n1030, ZN => n13492);
   U8466 : NAND2_X2 port map( A1 => n21279, A2 => n6066, ZN => n3531);
   U8469 : NAND2_X1 port map( A1 => n8754, A2 => n9896, ZN => n26985);
   U8470 : XOR2_X1 port map( A1 => n27396, A2 => n28159, Z => n5772);
   U8478 : INV_X2 port map( I => n20842, ZN => n27751);
   U8484 : XOR2_X1 port map( A1 => n26987, A2 => n3587, Z => n10241);
   U8487 : XOR2_X1 port map( A1 => n25627, A2 => n19356, Z => n26987);
   U8489 : INV_X2 port map( I => n26988, ZN => n28081);
   U8490 : INV_X2 port map( I => n16534, ZN => n26988);
   U8496 : INV_X1 port map( I => n17369, ZN => n26989);
   U8497 : NAND3_X2 port map( A1 => n3678, A2 => n26991, A3 => n26990, ZN => 
                           n4112);
   U8510 : NAND2_X2 port map( A1 => n24707, A2 => n23689, ZN => n28526);
   U8511 : NAND2_X2 port map( A1 => n5353, A2 => n26616, ZN => n25624);
   U8512 : BUF_X2 port map( I => n18535, Z => n26992);
   U8514 : NOR2_X2 port map( A1 => n28333, A2 => n28332, ZN => n3272);
   U8516 : XOR2_X1 port map( A1 => n15053, A2 => n19508, Z => n15052);
   U8518 : XOR2_X1 port map( A1 => n13715, A2 => n27448, Z => n15053);
   U8523 : NAND3_X2 port map( A1 => n5756, A2 => n27147, A3 => n8700, ZN => 
                           n20878);
   U8531 : AOI22_X2 port map( A1 => n26995, A2 => n25063, B1 => n13315, B2 => 
                           n709, ZN => n2347);
   U8532 : NAND2_X2 port map( A1 => n23253, A2 => n12364, ZN => n13864);
   U8536 : NAND2_X2 port map( A1 => n9012, A2 => n7865, ZN => n22237);
   U8540 : NOR2_X2 port map( A1 => n20826, A2 => n27751, ZN => n13072);
   U8547 : XOR2_X1 port map( A1 => n3751, A2 => n26996, Z => n28064);
   U8549 : INV_X2 port map( I => n16914, ZN => n26996);
   U8556 : NOR2_X2 port map( A1 => n16377, A2 => n16376, ZN => n3751);
   U8557 : XOR2_X1 port map( A1 => n7861, A2 => n8484, Z => n9158);
   U8559 : OAI21_X2 port map( A1 => n15996, A2 => n6237, B => n15995, ZN => 
                           n26998);
   U8562 : XOR2_X1 port map( A1 => n11787, A2 => n18113, Z => n18218);
   U8563 : NOR2_X2 port map( A1 => n8535, A2 => n24194, ZN => n18113);
   U8569 : INV_X2 port map( I => n28129, ZN => n21824);
   U8570 : NAND2_X2 port map( A1 => n26999, A2 => n12219, ZN => n14088);
   U8577 : OAI21_X2 port map( A1 => n26129, A2 => n19742, B => n975, ZN => 
                           n26999);
   U8581 : NAND2_X2 port map( A1 => n27708, A2 => n15049, ZN => n20168);
   U8584 : BUF_X4 port map( I => n3553, Z => n28231);
   U8586 : NAND2_X2 port map( A1 => n25956, A2 => n8171, ZN => n27044);
   U8587 : NAND2_X2 port map( A1 => n27000, A2 => n10094, ZN => n20155);
   U8588 : NOR2_X2 port map( A1 => n24720, A2 => n15461, ZN => n20259);
   U8590 : OR2_X2 port map( A1 => n21266, A2 => n11326, Z => n3504);
   U8591 : NAND2_X2 port map( A1 => n27256, A2 => n27003, ZN => n11077);
   U8598 : NOR2_X2 port map( A1 => n24804, A2 => n22109, ZN => n27003);
   U8600 : OR2_X1 port map( A1 => n7029, A2 => n23307, Z => n23644);
   U8601 : XOR2_X1 port map( A1 => n20576, A2 => n20714, Z => n22705);
   U8604 : OAI21_X2 port map( A1 => n11760, A2 => n21629, B => n11759, ZN => 
                           n27004);
   U8607 : NAND2_X1 port map( A1 => n19576, A2 => n5291, ZN => n27062);
   U8611 : XOR2_X1 port map( A1 => n16778, A2 => n16886, Z => n16486);
   U8612 : NOR2_X2 port map( A1 => n1374, A2 => n1373, ZN => n16778);
   U8614 : OAI21_X2 port map( A1 => n26355, A2 => n24179, B => n20122, ZN => 
                           n20124);
   U8616 : NAND4_X2 port map( A1 => n21676, A2 => n21674, A3 => n21673, A4 => 
                           n21675, ZN => n28230);
   U8620 : XOR2_X1 port map( A1 => n13449, A2 => n5742, Z => n13464);
   U8624 : OAI21_X2 port map( A1 => n3072, A2 => n25982, B => n25078, ZN => 
                           n13449);
   U8627 : XOR2_X1 port map( A1 => n24427, A2 => n7701, Z => n7700);
   U8632 : NOR2_X2 port map( A1 => n15041, A2 => n8646, ZN => n3833);
   U8634 : OAI21_X2 port map( A1 => n21098, A2 => n10558, B => n12309, ZN => 
                           n13020);
   U8636 : NAND2_X2 port map( A1 => n19169, A2 => n27006, ZN => n25283);
   U8638 : NAND2_X2 port map( A1 => n27007, A2 => n25276, ZN => n13752);
   U8641 : NAND2_X2 port map( A1 => n2068, A2 => n2549, ZN => n27008);
   U8642 : BUF_X2 port map( I => n9365, Z => n27010);
   U8646 : NAND4_X2 port map( A1 => n20904, A2 => n20903, A3 => n12034, A4 => 
                           n20905, ZN => n20907);
   U8650 : NAND2_X2 port map( A1 => n27011, A2 => n5951, ZN => n20326);
   U8654 : INV_X2 port map( I => n27759, ZN => n22879);
   U8662 : NAND2_X2 port map( A1 => n20329, A2 => n20415, ZN => n22183);
   U8665 : XOR2_X1 port map( A1 => n19176, A2 => n24242, Z => n27792);
   U8666 : XNOR2_X1 port map( A1 => n21257, A2 => n21369, ZN => n13680);
   U8667 : NAND3_X2 port map( A1 => n15194, A2 => n15192, A3 => n13233, ZN => 
                           n21369);
   U8669 : XOR2_X1 port map( A1 => n27012, A2 => n14001, Z => n19672);
   U8670 : XOR2_X1 port map( A1 => n19347, A2 => n12228, Z => n27012);
   U8672 : NOR3_X1 port map( A1 => n12979, A2 => n27631, A3 => n10564, ZN => 
                           n25149);
   U8677 : NAND2_X1 port map( A1 => n3406, A2 => n28343, ZN => n25284);
   U8678 : XOR2_X1 port map( A1 => n25361, A2 => n853, Z => n2306);
   U8680 : NAND2_X2 port map( A1 => n7184, A2 => n2095, ZN => n27290);
   U8681 : NAND2_X2 port map( A1 => n21098, A2 => n12066, ZN => n7184);
   U8683 : NAND2_X2 port map( A1 => n26154, A2 => n11052, ZN => n11400);
   U8684 : INV_X2 port map( I => n13333, ZN => n27013);
   U8685 : NOR2_X2 port map( A1 => n27013, A2 => n2544, ZN => n11398);
   U8686 : XOR2_X1 port map( A1 => n9548, A2 => n27014, Z => n9550);
   U8689 : XOR2_X1 port map( A1 => n20774, A2 => n15651, Z => n27014);
   U8690 : NAND3_X1 port map( A1 => n10891, A2 => n23439, A3 => n7237, ZN => 
                           n27015);
   U8691 : NAND2_X2 port map( A1 => n27016, A2 => n13263, ZN => n14580);
   U8695 : XOR2_X1 port map( A1 => n12114, A2 => n1975, Z => n6087);
   U8698 : NAND2_X2 port map( A1 => n13865, A2 => n13868, ZN => n12114);
   U8699 : OAI21_X2 port map( A1 => n26382, A2 => n8255, B => n19796, ZN => 
                           n19797);
   U8701 : INV_X4 port map( I => n10904, ZN => n18505);
   U8702 : NAND2_X2 port map( A1 => n1435, A2 => n5353, ZN => n12634);
   U8704 : NAND2_X1 port map( A1 => n27522, A2 => n9268, ZN => n7548);
   U8706 : NAND3_X1 port map( A1 => n4574, A2 => n23740, A3 => n21777, ZN => 
                           n28024);
   U8708 : XOR2_X1 port map( A1 => n17029, A2 => n17063, Z => n8705);
   U8712 : XOR2_X1 port map( A1 => n16806, A2 => n1651, Z => n17064);
   U8716 : OAI21_X2 port map( A1 => n23349, A2 => n1048, B => n1991, ZN => 
                           n16806);
   U8721 : AOI21_X2 port map( A1 => n16460, A2 => n13758, B => n27017, ZN => 
                           n16462);
   U8723 : OAI21_X2 port map( A1 => n27018, A2 => n27489, B => n17792, ZN => 
                           n18120);
   U8728 : NAND2_X1 port map( A1 => n9733, A2 => n2605, ZN => n27018);
   U8729 : BUF_X2 port map( I => n14513, Z => n1101);
   U8731 : NAND2_X2 port map( A1 => n12266, A2 => n12265, ZN => n4311);
   U8734 : NAND3_X2 port map( A1 => n28054, A2 => n9654, A3 => n4430, ZN => 
                           n27190);
   U8736 : NOR2_X1 port map( A1 => n28400, A2 => n13739, ZN => n13069);
   U8738 : NAND2_X2 port map( A1 => n8385, A2 => n8384, ZN => n22643);
   U8743 : OAI21_X2 port map( A1 => n6558, A2 => n14784, B => n166, ZN => n8385
                           );
   U8745 : XOR2_X1 port map( A1 => n13712, A2 => n13711, Z => n13710);
   U8746 : XOR2_X1 port map( A1 => n27020, A2 => n4043, Z => n5475);
   U8751 : XOR2_X1 port map( A1 => n19518, A2 => n27039, Z => n27020);
   U8752 : OAI21_X2 port map( A1 => n806, A2 => n9956, B => n8733, ZN => n27021
                           );
   U8754 : XOR2_X1 port map( A1 => n14694, A2 => n20534, Z => n3422);
   U8755 : XOR2_X1 port map( A1 => n20379, A2 => n11389, Z => n14694);
   U8756 : XOR2_X1 port map( A1 => n27022, A2 => n16832, Z => n16846);
   U8762 : XOR2_X1 port map( A1 => n15556, A2 => n6582, Z => n27022);
   U8763 : NAND3_X2 port map( A1 => n18845, A2 => n1813, A3 => n8557, ZN => 
                           n19231);
   U8766 : AOI22_X2 port map( A1 => n856, A2 => n20197, B1 => n733, B2 => 
                           n22807, ZN => n7566);
   U8767 : NAND2_X2 port map( A1 => n27294, A2 => n14443, ZN => n6756);
   U8772 : BUF_X1 port map( I => n19014, Z => n27138);
   U8775 : XOR2_X1 port map( A1 => n18172, A2 => n14026, Z => n18016);
   U8776 : NAND2_X1 port map( A1 => n5450, A2 => n27023, ZN => n7312);
   U8785 : XOR2_X1 port map( A1 => n15272, A2 => n12501, Z => n15273);
   U8786 : INV_X2 port map( I => n27024, ZN => n7289);
   U8789 : AOI21_X2 port map( A1 => n13311, A2 => n26041, B => n27025, ZN => 
                           n27024);
   U8800 : INV_X2 port map( I => n18294, ZN => n27026);
   U8801 : INV_X2 port map( I => n27027, ZN => n18357);
   U8807 : NOR2_X2 port map( A1 => n25592, A2 => n12542, ZN => n19102);
   U8810 : NAND2_X2 port map( A1 => n27028, A2 => n18399, ZN => n12962);
   U8812 : NAND2_X1 port map( A1 => n992, A2 => n26831, ZN => n27028);
   U8813 : OAI21_X2 port map( A1 => n12066, A2 => n12309, B => n21993, ZN => 
                           n23335);
   U8816 : NAND2_X2 port map( A1 => n12338, A2 => n18947, ZN => n19005);
   U8817 : NOR2_X2 port map( A1 => n12735, A2 => n12736, ZN => n12338);
   U8819 : NAND2_X1 port map( A1 => n3233, A2 => n17774, ZN => n17777);
   U8824 : AND2_X1 port map( A1 => n205, A2 => n19400, Z => n28111);
   U8828 : NAND2_X2 port map( A1 => n5282, A2 => n5281, ZN => n413);
   U8832 : NAND3_X1 port map( A1 => n10858, A2 => n26712, A3 => n12836, ZN => 
                           n13272);
   U8837 : NAND2_X1 port map( A1 => n2377, A2 => n14639, ZN => n5409);
   U8840 : AND2_X1 port map( A1 => n3347, A2 => n23245, Z => n24808);
   U8841 : NAND3_X2 port map( A1 => n26731, A2 => n27519, A3 => n27030, ZN => 
                           n20458);
   U8843 : AOI22_X1 port map( A1 => n20232, A2 => n8910, B1 => n20088, B2 => 
                           n14641, ZN => n27030);
   U8844 : XOR2_X1 port map( A1 => n20767, A2 => n21185, Z => n20568);
   U8847 : NAND2_X2 port map( A1 => n20199, A2 => n20198, ZN => n21185);
   U8850 : XOR2_X1 port map( A1 => n8953, A2 => n26429, Z => n6029);
   U8856 : AOI22_X2 port map( A1 => n24816, A2 => n14982, B1 => n14116, B2 => 
                           n17948, ZN => n14981);
   U8860 : XOR2_X1 port map( A1 => n319, A2 => n27031, Z => n5505);
   U8862 : XOR2_X1 port map( A1 => n18356, A2 => n18357, Z => n27031);
   U8863 : XOR2_X1 port map( A1 => n19272, A2 => n21411, Z => n22287);
   U8864 : NAND2_X2 port map( A1 => n18657, A2 => n18656, ZN => n19272);
   U8870 : NOR2_X2 port map( A1 => n27823, A2 => n23782, ZN => n5883);
   U8872 : XOR2_X1 port map( A1 => n20422, A2 => n1589, Z => n1588);
   U8873 : NAND2_X2 port map( A1 => n17716, A2 => n27032, ZN => n10056);
   U8878 : AOI22_X2 port map( A1 => n24330, A2 => n24640, B1 => n14351, B2 => 
                           n17845, ZN => n27032);
   U8879 : NAND2_X1 port map( A1 => n27368, A2 => n11385, ZN => n28087);
   U8881 : NAND3_X2 port map( A1 => n15524, A2 => n13768, A3 => n13052, ZN => 
                           n11385);
   U8883 : NAND3_X2 port map( A1 => n27033, A2 => n2396, A3 => n2399, ZN => 
                           n12697);
   U8884 : NAND3_X2 port map( A1 => n27697, A2 => n2395, A3 => n10323, ZN => 
                           n27033);
   U8887 : NAND2_X2 port map( A1 => n27151, A2 => n24075, ZN => n27034);
   U8888 : XOR2_X1 port map( A1 => n11964, A2 => n27035, Z => n28440);
   U8892 : XOR2_X1 port map( A1 => n22761, A2 => n26656, Z => n27035);
   U8897 : OAI21_X2 port map( A1 => n27724, A2 => n22311, B => n24998, ZN => 
                           n2967);
   U8906 : XOR2_X1 port map( A1 => n7598, A2 => n18286, Z => n18198);
   U8910 : NOR2_X2 port map( A1 => n13944, A2 => n13943, ZN => n7598);
   U8911 : XOR2_X1 port map( A1 => n27036, A2 => n14598, Z => Ciphertext(138));
   U8915 : NAND3_X1 port map( A1 => n21471, A2 => n21470, A3 => n21469, ZN => 
                           n27036);
   U8916 : NAND2_X1 port map( A1 => n27426, A2 => n21063, ZN => n3645);
   U8917 : XOR2_X1 port map( A1 => n3594, A2 => n3595, Z => n27426);
   U8919 : NAND2_X2 port map( A1 => n10841, A2 => n10840, ZN => n8683);
   U8923 : NAND2_X2 port map( A1 => n27037, A2 => n12393, ZN => n2079);
   U8925 : OAI22_X2 port map( A1 => n27038, A2 => n818, B1 => n18965, B2 => 
                           n989, ZN => n18966);
   U8927 : NAND2_X1 port map( A1 => n14683, A2 => n5746, ZN => n26520);
   U8928 : OR2_X1 port map( A1 => n17964, A2 => n23023, Z => n27920);
   U8931 : XOR2_X1 port map( A1 => n12725, A2 => n6707, Z => n6706);
   U8935 : XOR2_X1 port map( A1 => n11794, A2 => n11679, Z => n12725);
   U8943 : INV_X2 port map( I => n21714, ZN => n5396);
   U8945 : XOR2_X1 port map( A1 => n3291, A2 => n4048, Z => n27039);
   U8948 : NAND2_X2 port map( A1 => n10226, A2 => n10222, ZN => n13092);
   U8951 : INV_X2 port map( I => n3812, ZN => n19526);
   U8953 : XNOR2_X1 port map( A1 => n21758, A2 => n11417, ZN => n3812);
   U8959 : XOR2_X1 port map( A1 => n27041, A2 => n24659, Z => n15485);
   U8960 : XOR2_X1 port map( A1 => n14026, A2 => n1970, Z => n27041);
   U8961 : NAND2_X2 port map( A1 => n21297, A2 => n21444, ZN => n27042);
   U8962 : AND2_X1 port map( A1 => n15255, A2 => n7370, Z => n15401);
   U8963 : XOR2_X1 port map( A1 => n4332, A2 => n7815, Z => n5277);
   U8964 : CLKBUF_X4 port map( I => n10061, Z => n10058);
   U8967 : INV_X4 port map( I => n27632, ZN => n26396);
   U8968 : AND2_X1 port map( A1 => n27346, A2 => n24800, Z => n28201);
   U8969 : BUF_X4 port map( I => n19144, Z => n27043);
   U8970 : BUF_X4 port map( I => n15529, Z => n10015);
   U8977 : NAND2_X2 port map( A1 => n23979, A2 => n13235, ZN => n17762);
   U8978 : INV_X2 port map( I => n13473, ZN => n13472);
   U8993 : NAND3_X2 port map( A1 => n11207, A2 => n11209, A3 => n22501, ZN => 
                           n13473);
   U8999 : XOR2_X1 port map( A1 => n28325, A2 => n18209, Z => n7475);
   U9000 : XOR2_X1 port map( A1 => n883, A2 => n18103, Z => n18240);
   U9001 : INV_X2 port map( I => n18337, ZN => n883);
   U9005 : NOR2_X2 port map( A1 => n27961, A2 => n27808, ZN => n18337);
   U9007 : NAND2_X2 port map( A1 => n15888, A2 => n27045, ZN => n16981);
   U9011 : OAI21_X2 port map( A1 => n15613, A2 => n15614, B => n26105, ZN => 
                           n27045);
   U9014 : NAND2_X2 port map( A1 => n12057, A2 => n3481, ZN => n12053);
   U9016 : NAND2_X2 port map( A1 => n25052, A2 => n27046, ZN => n12191);
   U9018 : NAND2_X2 port map( A1 => n27047, A2 => n23831, ZN => n14033);
   U9022 : XOR2_X1 port map( A1 => n15726, A2 => n20440, Z => n24906);
   U9029 : XOR2_X1 port map( A1 => n20566, A2 => n7044, Z => n15726);
   U9034 : INV_X2 port map( I => n25013, ZN => n27048);
   U9036 : NOR2_X2 port map( A1 => n27048, A2 => n24458, ZN => n6903);
   U9039 : INV_X2 port map( I => n15729, ZN => n21058);
   U9042 : XOR2_X1 port map( A1 => n13359, A2 => n14248, Z => n15729);
   U9045 : XNOR2_X1 port map( A1 => n18179, A2 => n18180, ZN => n18284);
   U9046 : XOR2_X1 port map( A1 => n27447, A2 => n6523, Z => n8488);
   U9047 : OR2_X1 port map( A1 => n21456, A2 => n24680, Z => n21587);
   U9048 : NAND3_X1 port map( A1 => n10151, A2 => n5934, A3 => n20312, ZN => 
                           n6096);
   U9052 : OAI21_X2 port map( A1 => n9811, A2 => n9814, B => n9809, ZN => 
                           n10151);
   U9054 : NAND2_X2 port map( A1 => n19748, A2 => n19923, ZN => n19761);
   U9056 : NAND2_X1 port map( A1 => n5396, A2 => n27049, ZN => n27811);
   U9057 : NAND2_X1 port map( A1 => n10588, A2 => n9979, ZN => n27049);
   U9063 : NAND2_X2 port map( A1 => n110, A2 => n3627, ZN => n27368);
   U9064 : OAI21_X1 port map( A1 => n4274, A2 => n2185, B => n20023, ZN => 
                           n3883);
   U9067 : NAND2_X2 port map( A1 => n28426, A2 => n5249, ZN => n4274);
   U9071 : XOR2_X1 port map( A1 => n19501, A2 => n19394, Z => n23130);
   U9072 : NAND2_X2 port map( A1 => n28304, A2 => n6509, ZN => n3983);
   U9077 : OAI21_X2 port map( A1 => n5040, A2 => n22920, B => n27225, ZN => 
                           n5038);
   U9078 : NOR2_X2 port map( A1 => n23322, A2 => n26767, ZN => n10411);
   U9081 : INV_X2 port map( I => n18258, ZN => n5542);
   U9082 : OAI22_X2 port map( A1 => n2900, A2 => n17691, B1 => n2898, B2 => 
                           n23564, ZN => n18258);
   U9087 : NAND3_X1 port map( A1 => n26680, A2 => n23494, A3 => n27648, ZN => 
                           n8667);
   U9092 : NAND2_X1 port map( A1 => n14283, A2 => n10763, ZN => n11001);
   U9101 : NOR2_X1 port map( A1 => n13693, A2 => n13320, ZN => n17473);
   U9114 : NAND2_X2 port map( A1 => n12260, A2 => n12259, ZN => n15220);
   U9119 : NAND2_X2 port map( A1 => n19506, A2 => n19393, ZN => n12260);
   U9122 : XOR2_X1 port map( A1 => n15743, A2 => n5600, Z => n5599);
   U9125 : XOR2_X1 port map( A1 => n18077, A2 => n5602, Z => n15743);
   U9134 : INV_X4 port map( I => n26055, ZN => n26144);
   U9138 : NAND2_X1 port map( A1 => n17348, A2 => n2377, ZN => n3787);
   U9143 : NAND2_X2 port map( A1 => n21538, A2 => n4827, ZN => n21525);
   U9149 : INV_X2 port map( I => n9131, ZN => n21278);
   U9150 : XOR2_X1 port map( A1 => n21299, A2 => n16961, Z => n4260);
   U9154 : NAND3_X2 port map( A1 => n10487, A2 => n12800, A3 => n12802, ZN => 
                           n21299);
   U9155 : XOR2_X1 port map( A1 => n27051, A2 => n20467, Z => Ciphertext(29));
   U9157 : OAI22_X1 port map( A1 => n20465, A2 => n20693, B1 => n20466, B2 => 
                           n8388, ZN => n27051);
   U9159 : NOR2_X2 port map( A1 => n17894, A2 => n26642, ZN => n2751);
   U9160 : XOR2_X1 port map( A1 => n1402, A2 => n16939, Z => n1401);
   U9166 : XOR2_X1 port map( A1 => n2266, A2 => n2265, Z => n16939);
   U9167 : XOR2_X1 port map( A1 => n18208, A2 => n12932, Z => n12095);
   U9170 : AOI22_X2 port map( A1 => n23430, A2 => n18254, B1 => n18253, B2 => 
                           n23138, ZN => n19261);
   U9171 : INV_X4 port map( I => n20339, ZN => n20152);
   U9173 : NAND2_X2 port map( A1 => n19106, A2 => n6778, ZN => n8134);
   U9174 : AND2_X1 port map( A1 => n401, A2 => n10559, Z => n24607);
   U9176 : AOI21_X2 port map( A1 => n14153, A2 => n5047, B => n5049, ZN => 
                           n14152);
   U9183 : NAND3_X2 port map( A1 => n47, A2 => n3346, A3 => n21842, ZN => 
                           n14717);
   U9186 : XOR2_X1 port map( A1 => n10069, A2 => n10070, Z => n13665);
   U9187 : OAI21_X2 port map( A1 => n17575, A2 => n17574, B => n17501, ZN => 
                           n27619);
   U9188 : XOR2_X1 port map( A1 => n1689, A2 => n12555, Z => n11610);
   U9194 : NAND2_X1 port map( A1 => n21499, A2 => n21501, ZN => n27052);
   U9196 : INV_X2 port map( I => n12100, ZN => n23010);
   U9199 : NAND2_X2 port map( A1 => n3267, A2 => n13645, ZN => n12100);
   U9200 : BUF_X4 port map( I => n8383, Z => n28287);
   U9203 : INV_X4 port map( I => n20279, ZN => n858);
   U9207 : NAND2_X2 port map( A1 => n8166, A2 => n8167, ZN => n20279);
   U9209 : NAND3_X2 port map( A1 => n27053, A2 => n27492, A3 => n18833, ZN => 
                           n28216);
   U9210 : NAND2_X2 port map( A1 => n27279, A2 => n21776, ZN => n27053);
   U9211 : XOR2_X1 port map( A1 => n27054, A2 => n11472, Z => Ciphertext(149));
   U9212 : AOI22_X1 port map( A1 => n21537, A2 => n21536, B1 => n6972, B2 => 
                           n9575, ZN => n27054);
   U9215 : NAND2_X2 port map( A1 => n20194, A2 => n20294, ZN => n20146);
   U9217 : NAND2_X2 port map( A1 => n28201, A2 => n8190, ZN => n20194);
   U9218 : XOR2_X1 port map( A1 => n10004, A2 => n23312, Z => n25354);
   U9225 : NOR2_X2 port map( A1 => n13508, A2 => n18541, ZN => n26417);
   U9234 : NOR2_X2 port map( A1 => n348, A2 => n7350, ZN => n18541);
   U9235 : AOI22_X2 port map( A1 => n10808, A2 => n13924, B1 => n12503, B2 => 
                           n26577, ZN => n28195);
   U9237 : NAND2_X2 port map( A1 => n10965, A2 => n12255, ZN => n4793);
   U9238 : AOI22_X2 port map( A1 => n19053, A2 => n24061, B1 => n23931, B2 => 
                           n22346, ZN => n10965);
   U9246 : XOR2_X1 port map( A1 => n9034, A2 => n24176, Z => n13679);
   U9249 : XOR2_X1 port map( A1 => n27996, A2 => n19494, Z => n9034);
   U9251 : AOI22_X2 port map( A1 => n1203, A2 => n6076, B1 => n21842, B2 => 
                           n17864, ZN => n2898);
   U9253 : AOI22_X2 port map( A1 => n28492, A2 => n24693, B1 => n18847, B2 => 
                           n7260, ZN => n15100);
   U9259 : XOR2_X1 port map( A1 => n640, A2 => n8260, Z => n27943);
   U9264 : NAND2_X2 port map( A1 => n27056, A2 => n27055, ZN => n6975);
   U9267 : INV_X2 port map( I => n22646, ZN => n27056);
   U9272 : NAND2_X2 port map( A1 => n2324, A2 => n24514, ZN => n22646);
   U9273 : NAND3_X2 port map( A1 => n27716, A2 => n21499, A3 => n3504, ZN => 
                           n5172);
   U9276 : XOR2_X1 port map( A1 => n27057, A2 => n26793, Z => Ciphertext(132));
   U9280 : AOI22_X1 port map( A1 => n7946, A2 => n10851, B1 => n7945, B2 => 
                           n21455, ZN => n27057);
   U9281 : OR2_X1 port map( A1 => n26754, A2 => n12595, Z => n12639);
   U9285 : NAND2_X2 port map( A1 => n27711, A2 => n5172, ZN => n11492);
   U9291 : XOR2_X1 port map( A1 => n27726, A2 => n17753, Z => n8361);
   U9293 : XOR2_X1 port map( A1 => n25892, A2 => n3701, Z => n17753);
   U9294 : NAND2_X1 port map( A1 => n7312, A2 => n21587, ZN => n27163);
   U9295 : NAND2_X1 port map( A1 => n8205, A2 => n25959, ZN => n8204);
   U9297 : OR2_X1 port map( A1 => n11492, A2 => n12011, Z => n6080);
   U9299 : NAND2_X2 port map( A1 => n14519, A2 => n1271, ZN => n16014);
   U9302 : OR2_X1 port map( A1 => n5541, A2 => n12834, Z => n17326);
   U9306 : NAND2_X2 port map( A1 => n450, A2 => n15623, ZN => n1800);
   U9308 : INV_X4 port map( I => n14180, ZN => n8009);
   U9317 : NAND2_X2 port map( A1 => n24986, A2 => n10231, ZN => n14180);
   U9319 : OR2_X1 port map( A1 => n15986, A2 => n15984, Z => n16022);
   U9320 : OAI22_X1 port map( A1 => n27058, A2 => n9019, B1 => n16736, B2 => 
                           n6955, ZN => n11039);
   U9324 : OAI21_X1 port map( A1 => n16644, A2 => n25766, B => n6058, ZN => 
                           n27058);
   U9325 : NAND2_X2 port map( A1 => n19211, A2 => n19210, ZN => n25006);
   U9329 : NAND3_X2 port map( A1 => n11559, A2 => n19206, A3 => n19203, ZN => 
                           n19211);
   U9330 : NAND2_X2 port map( A1 => n25697, A2 => n1617, ZN => n9630);
   U9333 : NAND2_X2 port map( A1 => n13984, A2 => n25198, ZN => n18799);
   U9337 : NOR2_X2 port map( A1 => n27060, A2 => n6334, ZN => n6339);
   U9339 : NAND3_X2 port map( A1 => n26091, A2 => n6338, A3 => n6336, ZN => 
                           n27060);
   U9348 : NAND2_X2 port map( A1 => n27061, A2 => n27957, ZN => n18813);
   U9350 : NAND2_X2 port map( A1 => n23390, A2 => n23540, ZN => n27061);
   U9351 : NAND2_X2 port map( A1 => n27711, A2 => n5172, ZN => n27431);
   U9353 : XOR2_X1 port map( A1 => n21260, A2 => n11578, Z => n23646);
   U9354 : XOR2_X1 port map( A1 => n19237, A2 => n19556, Z => n18521);
   U9359 : XOR2_X1 port map( A1 => n13906, A2 => n8957, Z => n19556);
   U9360 : OR3_X1 port map( A1 => n9879, A2 => n27161, A3 => n9362, Z => n22489
                           );
   U9361 : BUF_X4 port map( I => n13925, Z => n13924);
   U9363 : XOR2_X1 port map( A1 => n12279, A2 => n3000, Z => n27267);
   U9365 : NAND2_X1 port map( A1 => n8166, A2 => n8167, ZN => n22786);
   U9370 : NOR2_X2 port map( A1 => n27062, A2 => n12472, ZN => n19967);
   U9372 : INV_X1 port map( I => n27063, ZN => n9573);
   U9374 : NAND3_X1 port map( A1 => n24567, A2 => n24560, A3 => n4127, ZN => 
                           n27063);
   U9376 : NAND2_X1 port map( A1 => n10818, A2 => n27276, ZN => n11257);
   U9383 : NOR2_X1 port map( A1 => n22111, A2 => n22112, ZN => n10462);
   U9391 : NAND3_X2 port map( A1 => n18811, A2 => n27138, A3 => n18812, ZN => 
                           n19333);
   U9392 : XNOR2_X1 port map( A1 => n3574, A2 => n12366, ZN => n21926);
   U9394 : AOI22_X2 port map( A1 => n28449, A2 => n20308, B1 => n4491, B2 => 
                           n20307, ZN => n4966);
   U9396 : XOR2_X1 port map( A1 => n20552, A2 => n12181, Z => n21151);
   U9399 : AOI21_X2 port map( A1 => n24481, A2 => n20244, B => n28097, ZN => 
                           n20552);
   U9400 : XOR2_X1 port map( A1 => n16823, A2 => n24956, Z => n7948);
   U9403 : NAND2_X1 port map( A1 => n27065, A2 => n4665, ZN => n11361);
   U9405 : NAND2_X1 port map( A1 => n4664, A2 => n19694, ZN => n27065);
   U9413 : OAI21_X2 port map( A1 => n25927, A2 => n7330, B => n10610, ZN => 
                           n27066);
   U9414 : XOR2_X1 port map( A1 => n8293, A2 => n20467, Z => n5287);
   U9416 : OAI21_X1 port map( A1 => n10673, A2 => n17956, B => n27067, ZN => 
                           n27115);
   U9418 : INV_X2 port map( I => n23542, ZN => n27067);
   U9419 : NOR2_X2 port map( A1 => n13530, A2 => n18003, ZN => n27068);
   U9420 : INV_X1 port map( I => n9175, ZN => n27069);
   U9421 : AND2_X1 port map( A1 => n9450, A2 => n27069, Z => n8235);
   U9422 : NAND2_X2 port map( A1 => n6169, A2 => n4390, ZN => n18331);
   U9423 : NAND2_X2 port map( A1 => n2285, A2 => n6435, ZN => n22485);
   U9424 : NAND2_X2 port map( A1 => n25325, A2 => n8311, ZN => n20750);
   U9427 : OAI21_X2 port map( A1 => n14665, A2 => n6410, B => n22641, ZN => 
                           n25325);
   U9428 : XOR2_X1 port map( A1 => n16981, A2 => n14744, Z => n17082);
   U9429 : NOR2_X2 port map( A1 => n9276, A2 => n9275, ZN => n14744);
   U9431 : AOI22_X2 port map( A1 => n19040, A2 => n22894, B1 => n2726, B2 => 
                           n19041, ZN => n5700);
   U9432 : BUF_X8 port map( I => n25586, Z => n27492);
   U9439 : NOR2_X1 port map( A1 => n19775, A2 => n977, ZN => n19601);
   U9443 : XOR2_X1 port map( A1 => n19333, A2 => n19334, Z => n19504);
   U9444 : XOR2_X1 port map( A1 => n27070, A2 => n1287, Z => Ciphertext(150));
   U9445 : NOR2_X1 port map( A1 => n27112, A2 => n10100, ZN => n27070);
   U9450 : NAND3_X2 port map( A1 => n24749, A2 => n19395, A3 => n27071, ZN => 
                           n20376);
   U9451 : BUF_X2 port map( I => n27599, Z => n27072);
   U9453 : XOR2_X1 port map( A1 => n21979, A2 => n21314, Z => n12070);
   U9454 : AOI22_X2 port map( A1 => n12563, A2 => n6470, B1 => n23374, B2 => 
                           n13694, ZN => n12042);
   U9455 : AOI22_X2 port map( A1 => n16016, A2 => n16146, B1 => n16017, B2 => 
                           n11429, ZN => n21964);
   U9456 : NOR2_X1 port map( A1 => n15835, A2 => n16143, ZN => n11429);
   U9457 : XOR2_X1 port map( A1 => n2850, A2 => n767, Z => n3946);
   U9458 : NAND2_X2 port map( A1 => n7900, A2 => n7899, ZN => n26008);
   U9468 : NAND2_X1 port map( A1 => n24224, A2 => n23990, ZN => n24880);
   U9469 : AND2_X1 port map( A1 => n28546, A2 => n10570, Z => n11873);
   U9480 : AND2_X2 port map( A1 => n27473, A2 => n11094, Z => n24638);
   U9482 : OR2_X1 port map( A1 => n17956, A2 => n27135, Z => n14190);
   U9483 : OAI21_X2 port map( A1 => n21866, A2 => n3956, B => n27075, ZN => 
                           n16602);
   U9484 : AOI22_X2 port map( A1 => n28012, A2 => n28011, B1 => n12274, B2 => 
                           n16013, ZN => n27075);
   U9485 : NAND2_X2 port map( A1 => n25202, A2 => n27076, ZN => n12797);
   U9488 : NAND2_X2 port map( A1 => n23774, A2 => n19151, ZN => n22155);
   U9489 : NAND3_X2 port map( A1 => n28486, A2 => n24124, A3 => n11726, ZN => 
                           n24107);
   U9493 : XOR2_X1 port map( A1 => n22731, A2 => n7329, Z => n383);
   U9494 : NAND2_X1 port map( A1 => n27077, A2 => n8771, ZN => n4328);
   U9501 : NOR2_X1 port map( A1 => n27078, A2 => n6465, ZN => n26604);
   U9503 : NAND2_X1 port map( A1 => n8145, A2 => n14423, ZN => n8144);
   U9505 : XOR2_X1 port map( A1 => n12071, A2 => n27079, Z => n15696);
   U9506 : XOR2_X1 port map( A1 => n12070, A2 => n12069, Z => n27079);
   U9507 : NAND2_X2 port map( A1 => n13902, A2 => n28023, ZN => n27779);
   U9508 : AOI21_X2 port map( A1 => n14872, A2 => n26721, B => n5554, ZN => 
                           n28437);
   U9510 : NOR2_X2 port map( A1 => n26417, A2 => n25118, ZN => n8988);
   U9511 : XOR2_X1 port map( A1 => n10084, A2 => n21187, Z => n20479);
   U9515 : XOR2_X1 port map( A1 => n20448, A2 => n20423, Z => n21187);
   U9524 : NAND2_X2 port map( A1 => n27081, A2 => n27080, ZN => n24594);
   U9527 : INV_X2 port map( I => n16355, ZN => n27081);
   U9533 : XOR2_X1 port map( A1 => n27082, A2 => n20702, Z => Ciphertext(27));
   U9534 : NAND4_X2 port map( A1 => n20699, A2 => n20698, A3 => n20700, A4 => 
                           n20701, ZN => n27082);
   U9535 : INV_X2 port map( I => n5345, ZN => n7350);
   U9537 : XOR2_X1 port map( A1 => n27695, A2 => n13296, Z => n5345);
   U9541 : NAND3_X2 port map( A1 => n17529, A2 => n9989, A3 => n22918, ZN => 
                           n27293);
   U9542 : NAND3_X2 port map( A1 => n5048, A2 => n675, A3 => n5047, ZN => 
                           n12800);
   U9543 : NOR3_X1 port map( A1 => n8227, A2 => n13278, A3 => n15478, ZN => 
                           n28006);
   U9545 : NOR3_X1 port map( A1 => n27083, A2 => n21522, A3 => n6957, ZN => 
                           n28219);
   U9550 : NOR2_X1 port map( A1 => n21521, A2 => n14229, ZN => n27083);
   U9551 : XOR2_X1 port map( A1 => n3356, A2 => n20389, Z => n28133);
   U9556 : XOR2_X1 port map( A1 => n12355, A2 => n20388, Z => n3356);
   U9559 : AOI21_X2 port map( A1 => n9099, A2 => n915, B => n27085, ZN => 
                           n13138);
   U9560 : OAI22_X2 port map( A1 => n9098, A2 => n16320, B1 => n12734, B2 => 
                           n16321, ZN => n27085);
   U9569 : XOR2_X1 port map( A1 => n19326, A2 => n27086, Z => n23482);
   U9574 : XOR2_X1 port map( A1 => n19443, A2 => n19324, Z => n27086);
   U9575 : INV_X4 port map( I => n4827, ZN => n21531);
   U9577 : NAND3_X2 port map( A1 => n5031, A2 => n5029, A3 => n5030, ZN => 
                           n12246);
   U9578 : XOR2_X1 port map( A1 => n26119, A2 => n20378, Z => n20815);
   U9580 : XOR2_X1 port map( A1 => n20334, A2 => n7248, Z => n20378);
   U9581 : BUF_X2 port map( I => n13684, Z => n27087);
   U9588 : CLKBUF_X12 port map( I => n18169, Z => n28355);
   U9589 : XOR2_X1 port map( A1 => n22855, A2 => n11336, Z => n27088);
   U9593 : NOR2_X1 port map( A1 => n1422, A2 => n1424, ZN => n1421);
   U9600 : OAI22_X1 port map( A1 => n12703, A2 => n18124, B1 => n12820, B2 => 
                           n24133, ZN => n12702);
   U9610 : INV_X4 port map( I => n18012, ZN => n27410);
   U9612 : NAND2_X2 port map( A1 => n27940, A2 => n22157, ZN => n4833);
   U9614 : NOR2_X2 port map( A1 => n3271, A2 => n3885, ZN => n27940);
   U9615 : XNOR2_X1 port map( A1 => n16940, A2 => n14023, ZN => n27167);
   U9621 : NAND2_X2 port map( A1 => n9358, A2 => n10015, ZN => n17270);
   U9627 : AOI22_X2 port map( A1 => n21135, A2 => n26773, B1 => n20263, B2 => 
                           n13023, ZN => n27089);
   U9636 : XOR2_X1 port map( A1 => n8244, A2 => n27090, Z => n15349);
   U9637 : XOR2_X1 port map( A1 => n18122, A2 => n13109, Z => n27090);
   U9642 : XOR2_X1 port map( A1 => n20563, A2 => n20762, Z => n24493);
   U9644 : NAND2_X2 port map( A1 => n9775, A2 => n27092, ZN => n8262);
   U9647 : OAI21_X1 port map( A1 => n9778, A2 => n17432, B => n17431, ZN => 
                           n27092);
   U9652 : OAI22_X2 port map( A1 => n12308, A2 => n12307, B1 => n27094, B2 => 
                           n27093, ZN => n21052);
   U9654 : NAND2_X1 port map( A1 => n6962, A2 => n26512, ZN => n27093);
   U9655 : NAND2_X2 port map( A1 => n8215, A2 => n21692, ZN => n1765);
   U9658 : NOR2_X2 port map( A1 => n27095, A2 => n8660, ZN => n10134);
   U9659 : NAND2_X2 port map( A1 => n7324, A2 => n15492, ZN => n27095);
   U9665 : INV_X2 port map( I => n24522, ZN => n18752);
   U9666 : NOR2_X2 port map( A1 => n27096, A2 => n7171, ZN => n9538);
   U9669 : INV_X2 port map( I => n21734, ZN => n27098);
   U9670 : OAI21_X2 port map( A1 => n28242, A2 => n28241, B => n27099, ZN => 
                           n8957);
   U9671 : NAND2_X2 port map( A1 => n25494, A2 => n28143, ZN => n27099);
   U9672 : BUF_X2 port map( I => n28295, Z => n27100);
   U9673 : XOR2_X1 port map( A1 => n2098, A2 => n18072, Z => n15174);
   U9674 : NOR2_X1 port map( A1 => n4657, A2 => n28268, ZN => n19795);
   U9677 : INV_X2 port map( I => n13909, ZN => n28268);
   U9678 : XOR2_X1 port map( A1 => n10390, A2 => n10391, Z => n13909);
   U9681 : BUF_X4 port map( I => n20324, Z => n21772);
   U9683 : OAI21_X2 port map( A1 => n9575, A2 => n21531, B => n30, ZN => n21537
                           );
   U9694 : NAND2_X2 port map( A1 => n8755, A2 => n23644, ZN => n13775);
   U9696 : OAI21_X2 port map( A1 => n20216, A2 => n10221, B => n20214, ZN => 
                           n10026);
   U9697 : BUF_X2 port map( I => n17942, Z => n27101);
   U9699 : XOR2_X1 port map( A1 => n27102, A2 => n302, Z => n27971);
   U9700 : XOR2_X1 port map( A1 => n11539, A2 => n27103, Z => n27102);
   U9701 : NAND2_X2 port map( A1 => n1365, A2 => n13928, ZN => n17935);
   U9702 : NOR2_X2 port map( A1 => n4402, A2 => n3147, ZN => n1365);
   U9703 : NAND2_X1 port map( A1 => n4917, A2 => n28295, ZN => n2781);
   U9705 : NOR2_X2 port map( A1 => n27660, A2 => n1513, ZN => n28295);
   U9707 : XOR2_X1 port map( A1 => n18258, A2 => n18234, Z => n18356);
   U9710 : NAND2_X2 port map( A1 => n27105, A2 => n1457, ZN => n27264);
   U9712 : NAND2_X2 port map( A1 => n946, A2 => n27266, ZN => n27105);
   U9715 : AOI22_X2 port map( A1 => n4161, A2 => n5407, B1 => n3674, B2 => 
                           n7960, ZN => n8638);
   U9716 : AOI22_X2 port map( A1 => n9052, A2 => n887, B1 => n4828, B2 => 
                           n17641, ZN => n26513);
   U9718 : NAND3_X2 port map( A1 => n17429, A2 => n27106, A3 => n22658, ZN => 
                           n17818);
   U9719 : INV_X4 port map( I => n27798, ZN => n24811);
   U9724 : INV_X2 port map( I => n14528, ZN => n23275);
   U9725 : XOR2_X1 port map( A1 => n4375, A2 => n4239, Z => n8795);
   U9726 : NOR2_X2 port map( A1 => n2100, A2 => n2099, ZN => n28370);
   U9727 : NOR2_X2 port map( A1 => n28490, A2 => n28100, ZN => n17007);
   U9729 : INV_X2 port map( I => n12022, ZN => n1024);
   U9737 : OAI21_X2 port map( A1 => n3093, A2 => n3095, B => n3092, ZN => 
                           n12022);
   U9743 : INV_X2 port map( I => n21120, ZN => n13444);
   U9744 : NAND2_X2 port map( A1 => n13445, A2 => n13446, ZN => n21120);
   U9747 : XOR2_X1 port map( A1 => n19510, A2 => n13918, Z => n19464);
   U9751 : XOR2_X1 port map( A1 => n7244, A2 => n17754, Z => n6272);
   U9753 : AOI22_X2 port map( A1 => n26478, A2 => n14826, B1 => n3682, B2 => 
                           n25542, ZN => n7244);
   U9755 : NAND2_X2 port map( A1 => n27107, A2 => n3380, ZN => n10027);
   U9758 : AOI22_X2 port map( A1 => n27837, A2 => n23529, B1 => n13758, B2 => 
                           n9500, ZN => n27107);
   U9761 : NAND2_X2 port map( A1 => n21274, A2 => n21273, ZN => n21276);
   U9762 : NOR2_X2 port map( A1 => n8398, A2 => n14546, ZN => n8923);
   U9763 : XOR2_X1 port map( A1 => n25312, A2 => n18029, Z => n18297);
   U9765 : NAND3_X2 port map( A1 => n17579, A2 => n14717, A3 => n14716, ZN => 
                           n18029);
   U9773 : NAND2_X2 port map( A1 => n19155, A2 => n6889, ZN => n24055);
   U9780 : NOR2_X2 port map( A1 => n18006, A2 => n3496, ZN => n6889);
   U9782 : XOR2_X1 port map( A1 => n21899, A2 => n17057, Z => n24013);
   U9785 : XOR2_X1 port map( A1 => n2994, A2 => n27108, Z => n1622);
   U9787 : NAND2_X2 port map( A1 => n8295, A2 => n27629, ZN => n2994);
   U9801 : XOR2_X1 port map( A1 => n19421, A2 => n19447, Z => n19523);
   U9806 : XOR2_X1 port map( A1 => n16486, A2 => n22698, Z => n2410);
   U9808 : NAND2_X1 port map( A1 => n5798, A2 => n5799, ZN => n26372);
   U9814 : AOI21_X2 port map( A1 => n18568, A2 => n18752, B => n6311, ZN => 
                           n6310);
   U9815 : INV_X1 port map( I => n19124, ZN => n27109);
   U9817 : OR2_X1 port map( A1 => n24743, A2 => n27109, Z => n3054);
   U9818 : NAND2_X2 port map( A1 => n26248, A2 => n27845, ZN => n4355);
   U9819 : NAND2_X2 port map( A1 => n27110, A2 => n2086, ZN => n2085);
   U9827 : OAI21_X2 port map( A1 => n27839, A2 => n24545, B => n1491, ZN => 
                           n27110);
   U9828 : NAND2_X2 port map( A1 => n27111, A2 => n7925, ZN => n23443);
   U9829 : NOR2_X2 port map( A1 => n2911, A2 => n7927, ZN => n27111);
   U9831 : AOI21_X1 port map( A1 => n10103, A2 => n12270, B => n22732, ZN => 
                           n27112);
   U9835 : INV_X1 port map( I => n19451, ZN => n27113);
   U9837 : NOR2_X2 port map( A1 => n26988, A2 => n6766, ZN => n16551);
   U9841 : NAND2_X2 port map( A1 => n19102, A2 => n7018, ZN => n11559);
   U9842 : INV_X1 port map( I => n3983, ZN => n24285);
   U9846 : XOR2_X1 port map( A1 => n18191, A2 => n18190, Z => n18196);
   U9847 : XOR2_X1 port map( A1 => n4288, A2 => n6675, Z => n18190);
   U9848 : NAND3_X2 port map( A1 => n25791, A2 => n20840, A3 => n20838, ZN => 
                           n28387);
   U9850 : OR2_X1 port map( A1 => n7085, A2 => n21563, Z => n27117);
   U9852 : INV_X2 port map( I => n24574, ZN => n27118);
   U9854 : XOR2_X1 port map( A1 => n10379, A2 => n22330, Z => n14291);
   U9856 : XOR2_X1 port map( A1 => n14538, A2 => n26613, Z => n23278);
   U9858 : NOR2_X2 port map( A1 => n17799, A2 => n17981, ZN => n8184);
   U9860 : INV_X2 port map( I => n17799, ZN => n8382);
   U9861 : XOR2_X1 port map( A1 => n28009, A2 => n27120, Z => n27283);
   U9863 : XOR2_X1 port map( A1 => n26012, A2 => n26495, Z => n27120);
   U9869 : AND2_X1 port map( A1 => n7807, A2 => n8468, Z => n8233);
   U9870 : XOR2_X1 port map( A1 => n7809, A2 => n7808, Z => n8246);
   U9872 : NAND2_X2 port map( A1 => n26325, A2 => n27121, ZN => n17125);
   U9874 : AOI22_X1 port map( A1 => n16684, A2 => n16685, B1 => n16686, B2 => 
                           n25994, ZN => n27121);
   U9876 : NAND3_X1 port map( A1 => n26698, A2 => n19768, A3 => n11470, ZN => 
                           n28146);
   U9879 : XOR2_X1 port map( A1 => n27848, A2 => n15038, Z => n16734);
   U9881 : NAND2_X1 port map( A1 => n27122, A2 => n22655, ZN => n28471);
   U9882 : XOR2_X1 port map( A1 => n6878, A2 => n10999, Z => n9244);
   U9884 : NOR2_X2 port map( A1 => n5775, A2 => n5773, ZN => n10999);
   U9885 : NAND2_X2 port map( A1 => n21918, A2 => n13066, ZN => n27821);
   U9891 : NOR2_X1 port map( A1 => n5081, A2 => n11413, ZN => n16535);
   U9892 : INV_X2 port map( I => n24458, ZN => n9879);
   U9895 : BUF_X2 port map( I => n28284, Z => n27123);
   U9899 : AND2_X1 port map( A1 => n713, A2 => n17578, Z => n22247);
   U9902 : XOR2_X1 port map( A1 => n7403, A2 => n22349, Z => n9017);
   U9905 : NAND3_X2 port map( A1 => n25811, A2 => n8401, A3 => n8063, ZN => 
                           n7403);
   U9906 : INV_X2 port map( I => n27124, ZN => n6375);
   U9907 : XOR2_X1 port map( A1 => n6376, A2 => n6377, Z => n27124);
   U9908 : INV_X2 port map( I => n6260, ZN => n11471);
   U9909 : OAI21_X2 port map( A1 => n23756, A2 => n25216, B => n27125, ZN => 
                           n26218);
   U9911 : XOR2_X1 port map( A1 => Plaintext(7), A2 => Key(7), Z => n28284);
   U9912 : NAND2_X2 port map( A1 => n14662, A2 => n18091, ZN => n26478);
   U9914 : NAND2_X2 port map( A1 => n24570, A2 => n28104, ZN => n14662);
   U9915 : XOR2_X1 port map( A1 => n3390, A2 => n11815, Z => n3603);
   U9919 : XOR2_X1 port map( A1 => n27126, A2 => n1297, Z => Ciphertext(74));
   U9921 : INV_X2 port map( I => n15448, ZN => n24870);
   U9923 : XOR2_X1 port map( A1 => n24258, A2 => n18013, Z => n13165);
   U9924 : XOR2_X1 port map( A1 => n13695, A2 => n14091, Z => n507);
   U9925 : XOR2_X1 port map( A1 => n27127, A2 => n10374, Z => n503);
   U9928 : XOR2_X1 port map( A1 => n23463, A2 => n25317, Z => n27127);
   U9929 : XOR2_X1 port map( A1 => n19234, A2 => n13949, Z => n19311);
   U9931 : NOR3_X2 port map( A1 => n1581, A2 => n5491, A3 => n18561, ZN => 
                           n19234);
   U9935 : AOI21_X2 port map( A1 => n5048, A2 => n20205, B => n12362, ZN => 
                           n3815);
   U9940 : NAND2_X2 port map( A1 => n1934, A2 => n27128, ZN => n20107);
   U9941 : NAND2_X1 port map( A1 => n1948, A2 => n6210, ZN => n27128);
   U9943 : INV_X2 port map( I => n12111, ZN => n12113);
   U9944 : NAND2_X2 port map( A1 => n24157, A2 => n24262, ZN => n12111);
   U9947 : BUF_X2 port map( I => n5080, Z => n27129);
   U9951 : NAND2_X2 port map( A1 => n27685, A2 => n12722, ZN => n5949);
   U9952 : NOR3_X2 port map( A1 => n27689, A2 => n708, A3 => n21024, ZN => 
                           n12490);
   U9953 : XOR2_X1 port map( A1 => n26416, A2 => n27130, Z => n8727);
   U9958 : XOR2_X1 port map( A1 => n18278, A2 => n9369, Z => n27130);
   U9959 : NAND2_X2 port map( A1 => n8820, A2 => n10156, ZN => n16819);
   U9961 : XOR2_X1 port map( A1 => n1944, A2 => n3845, Z => n6166);
   U9962 : XOR2_X1 port map( A1 => n25296, A2 => n13850, Z => n18654);
   U9963 : AOI22_X1 port map( A1 => n4022, A2 => n5042, B1 => n22828, B2 => 
                           n21727, ZN => n22522);
   U9965 : NOR2_X2 port map( A1 => n948, A2 => n4122, ZN => n4022);
   U9977 : NOR2_X2 port map( A1 => n22635, A2 => n8555, ZN => n2309);
   U9980 : XOR2_X1 port map( A1 => n27131, A2 => n16720, Z => n534);
   U9988 : XOR2_X1 port map( A1 => n24069, A2 => n16914, Z => n27131);
   U9991 : XNOR2_X1 port map( A1 => n19310, A2 => n14021, ZN => n27159);
   U9994 : NAND2_X2 port map( A1 => n8625, A2 => n8626, ZN => n17950);
   U9999 : XOR2_X1 port map( A1 => n28497, A2 => n14709, Z => n24735);
   U10001 : OAI22_X2 port map( A1 => n21793, A2 => n17409, B1 => n9898, B2 => 
                           n17408, ZN => n17410);
   U10002 : OAI21_X2 port map( A1 => n16505, A2 => n12039, B => n27133, ZN => 
                           n27828);
   U10005 : OAI21_X2 port map( A1 => n26186, A2 => n22712, B => n3874, ZN => 
                           n15645);
   U10009 : NAND2_X2 port map( A1 => n1421, A2 => n1425, ZN => n27573);
   U10011 : XOR2_X1 port map( A1 => n18351, A2 => n24659, Z => n26085);
   U10013 : XOR2_X1 port map( A1 => n27134, A2 => n1292, Z => Ciphertext(40));
   U10014 : NOR3_X1 port map( A1 => n24714, A2 => n21871, A3 => n13365, ZN => 
                           n27134);
   U10015 : XOR2_X1 port map( A1 => n19387, A2 => n1137, Z => n12049);
   U10020 : INV_X4 port map( I => n27135, ZN => n5402);
   U10021 : AND2_X2 port map( A1 => n6966, A2 => n27960, Z => n27135);
   U10022 : AOI21_X1 port map( A1 => n4779, A2 => n10673, B => n23542, ZN => 
                           n27961);
   U10025 : OAI21_X2 port map( A1 => n20710, A2 => n12140, B => n953, ZN => 
                           n24830);
   U10036 : NOR2_X1 port map( A1 => n666, A2 => n664, ZN => n19820);
   U10042 : XOR2_X1 port map( A1 => n26519, A2 => n14780, Z => n15540);
   U10044 : XOR2_X1 port map( A1 => n28325, A2 => n27145, Z => n4189);
   U10046 : XOR2_X1 port map( A1 => n27136, A2 => n17103, Z => n22849);
   U10047 : XOR2_X1 port map( A1 => n13344, A2 => n16868, Z => n17103);
   U10048 : INV_X4 port map( I => n9525, ZN => n13301);
   U10050 : NAND2_X2 port map( A1 => n13539, A2 => n24984, ZN => n9525);
   U10051 : XOR2_X1 port map( A1 => n13761, A2 => n20452, Z => n21240);
   U10052 : NAND2_X2 port map( A1 => n20221, A2 => n13762, ZN => n13761);
   U10058 : INV_X2 port map( I => n27139, ZN => n3880);
   U10059 : XOR2_X1 port map( A1 => n8438, A2 => n19313, Z => n27139);
   U10063 : NAND2_X2 port map( A1 => n13494, A2 => n5070, ZN => n23772);
   U10064 : NOR2_X2 port map( A1 => n12969, A2 => n27278, ZN => n13494);
   U10065 : INV_X2 port map( I => n27141, ZN => n21545);
   U10072 : NOR2_X2 port map( A1 => n27144, A2 => n27143, ZN => n2084);
   U10076 : NAND2_X2 port map( A1 => n2085, A2 => n5057, ZN => n11519);
   U10078 : NOR2_X2 port map( A1 => n22997, A2 => n26097, ZN => n6930);
   U10079 : XOR2_X1 port map( A1 => n3078, A2 => n3107, Z => n12696);
   U10082 : XOR2_X1 port map( A1 => n11183, A2 => n10445, Z => n21181);
   U10083 : INV_X4 port map( I => n9683, ZN => n2481);
   U10088 : AOI22_X2 port map( A1 => n7396, A2 => n20152, B1 => n24085, B2 => 
                           n11519, ZN => n27639);
   U10089 : BUF_X2 port map( I => n17855, Z => n27146);
   U10091 : NOR2_X2 port map( A1 => n3495, A2 => n3494, ZN => n19155);
   U10105 : AOI21_X1 port map( A1 => n2185, A2 => n4021, B => n26206, ZN => 
                           n7978);
   U10108 : INV_X2 port map( I => n7379, ZN => n9167);
   U10114 : INV_X4 port map( I => n26410, ZN => n28419);
   U10117 : NAND2_X2 port map( A1 => n2170, A2 => n2171, ZN => n23146);
   U10118 : AOI22_X2 port map( A1 => n2832, A2 => n183, B1 => n25722, B2 => 
                           n2833, ZN => n22778);
   U10120 : XOR2_X1 port map( A1 => n6761, A2 => n27148, Z => n6760);
   U10122 : XOR2_X1 port map( A1 => n20580, A2 => n27149, Z => n27148);
   U10128 : INV_X1 port map( I => n13859, ZN => n27149);
   U10129 : XOR2_X1 port map( A1 => n6507, A2 => n26398, Z => n4945);
   U10134 : XOR2_X1 port map( A1 => n6490, A2 => n9534, Z => n6507);
   U10136 : INV_X2 port map( I => n26178, ZN => n22381);
   U10146 : INV_X2 port map( I => n18428, ZN => n1168);
   U10150 : NAND2_X2 port map( A1 => n14745, A2 => n18552, ZN => n18428);
   U10157 : NAND2_X2 port map( A1 => n19, A2 => n22735, ZN => n20070);
   U10158 : NAND2_X2 port map( A1 => n19736, A2 => n976, ZN => n4226);
   U10159 : XOR2_X1 port map( A1 => n15485, A2 => n17628, Z => n18552);
   U10161 : AOI22_X2 port map( A1 => n1168, A2 => n18722, B1 => n3886, B2 => 
                           n1184, ZN => n27586);
   U10164 : AOI21_X2 port map( A1 => n17314, A2 => n1234, B => n23956, ZN => 
                           n23819);
   U10168 : NAND2_X2 port map( A1 => n15777, A2 => n15778, ZN => n27367);
   U10177 : OAI22_X2 port map( A1 => n27281, A2 => n14883, B1 => n18675, B2 => 
                           n18676, ZN => n27150);
   U10178 : XOR2_X1 port map( A1 => n16765, A2 => n2363, Z => n5964);
   U10182 : XOR2_X1 port map( A1 => n21995, A2 => n12147, Z => n16765);
   U10189 : OR2_X2 port map( A1 => n27453, A2 => n13896, Z => n18727);
   U10196 : XOR2_X1 port map( A1 => n24719, A2 => n18054, Z => n6364);
   U10197 : NAND3_X2 port map( A1 => n11718, A2 => n8714, A3 => n10924, ZN => 
                           n27151);
   U10204 : OAI22_X2 port map( A1 => n13485, A2 => n1101, B1 => n20132, B2 => 
                           n20319, ZN => n21153);
   U10210 : AOI22_X2 port map( A1 => n20317, A2 => n6998, B1 => n13754, B2 => 
                           n20316, ZN => n20319);
   U10211 : XOR2_X1 port map( A1 => n17109, A2 => n2225, Z => n16907);
   U10213 : NAND2_X2 port map( A1 => n5669, A2 => n23896, ZN => n17109);
   U10220 : XOR2_X1 port map( A1 => n7467, A2 => n4585, Z => n12071);
   U10221 : NAND2_X2 port map( A1 => n25803, A2 => n10043, ZN => n25802);
   U10225 : OAI22_X2 port map( A1 => n11453, A2 => n13646, B1 => n18605, B2 => 
                           n10569, ZN => n10043);
   U10226 : INV_X2 port map( I => n21212, ZN => n22057);
   U10230 : NAND3_X2 port map( A1 => n21178, A2 => n7377, A3 => n10551, ZN => 
                           n21212);
   U10231 : AOI21_X2 port map( A1 => n27155, A2 => n4331, B => n22450, ZN => 
                           n4329);
   U10232 : OAI21_X2 port map( A1 => n784, A2 => n1014, B => n882, ZN => n27155
                           );
   U10244 : XOR2_X1 port map( A1 => n18147, A2 => n6562, Z => n18299);
   U10246 : NAND2_X2 port map( A1 => n25668, A2 => n27667, ZN => n13333);
   U10249 : NAND2_X2 port map( A1 => n6482, A2 => n27156, ZN => n12421);
   U10254 : OAI21_X2 port map( A1 => n28122, A2 => n23706, B => n885, ZN => 
                           n27156);
   U10255 : NOR2_X2 port map( A1 => n4324, A2 => n27064, ZN => n28099);
   U10263 : OR2_X1 port map( A1 => n8723, A2 => n7134, Z => n9845);
   U10269 : XOR2_X1 port map( A1 => n9637, A2 => n26569, Z => n21295);
   U10270 : XOR2_X1 port map( A1 => n15119, A2 => n21183, Z => n13803);
   U10272 : NAND2_X2 port map( A1 => n19578, A2 => n19579, ZN => n21183);
   U10274 : INV_X1 port map( I => n24336, ZN => n22269);
   U10280 : XOR2_X1 port map( A1 => n27159, A2 => n5588, Z => n24336);
   U10281 : BUF_X4 port map( I => n10602, Z => n27484);
   U10293 : NAND2_X2 port map( A1 => n27856, A2 => n19605, ZN => n5838);
   U10295 : BUF_X2 port map( I => n6870, Z => n27161);
   U10298 : OR2_X1 port map( A1 => n28019, A2 => n2869, Z => n6835);
   U10301 : BUF_X2 port map( I => n16111, Z => n27162);
   U10307 : AOI22_X2 port map( A1 => n27163, A2 => n25064, B1 => n12012, B2 => 
                           n8751, ZN => n12011);
   U10309 : NOR2_X2 port map( A1 => n8425, A2 => n18458, ZN => n9097);
   U10310 : NOR2_X2 port map( A1 => n15168, A2 => n26477, ZN => n11249);
   U10311 : AOI22_X2 port map( A1 => n26347, A2 => n27164, B1 => n26671, B2 => 
                           n3347, ZN => n2808);
   U10314 : NAND2_X2 port map( A1 => n27165, A2 => n13140, ZN => n16820);
   U10315 : OAI22_X2 port map( A1 => n27166, A2 => n1558, B1 => n18918, B2 => 
                           n6708, ZN => n26256);
   U10316 : NAND2_X2 port map( A1 => n427, A2 => n869, ZN => n27166);
   U10318 : XOR2_X1 port map( A1 => n27167, A2 => n22146, Z => n27982);
   U10323 : XOR2_X1 port map( A1 => n3862, A2 => n19494, Z => n12580);
   U10325 : AOI22_X1 port map( A1 => n16083, A2 => n16256, B1 => n6605, B2 => 
                           n12035, ZN => n27832);
   U10326 : AND2_X1 port map( A1 => n19923, A2 => n669, Z => n25096);
   U10327 : XOR2_X1 port map( A1 => n13469, A2 => n8605, Z => n12691);
   U10328 : NOR2_X2 port map( A1 => n6472, A2 => n27976, ZN => n13469);
   U10330 : NOR2_X2 port map( A1 => n6766, A2 => n11658, ZN => n16474);
   U10333 : BUF_X2 port map( I => n17442, Z => n27168);
   U10336 : OAI21_X2 port map( A1 => n23534, A2 => n18693, B => n25802, ZN => 
                           n25368);
   U10339 : XOR2_X1 port map( A1 => n19363, A2 => n19224, Z => n9985);
   U10340 : NAND2_X2 port map( A1 => n26392, A2 => n18975, ZN => n19363);
   U10343 : NAND2_X2 port map( A1 => n20279, A2 => n7749, ZN => n13378);
   U10345 : AOI21_X2 port map( A1 => n18869, A2 => n18945, B => n22954, ZN => 
                           n19224);
   U10351 : NOR2_X2 port map( A1 => n28145, A2 => n27948, ZN => n1530);
   U10359 : NAND2_X2 port map( A1 => n27170, A2 => n3893, ZN => n4462);
   U10363 : OAI21_X2 port map( A1 => n16008, A2 => n15990, B => n5362, ZN => 
                           n27170);
   U10364 : XOR2_X1 port map( A1 => n19558, A2 => n19449, Z => n6085);
   U10368 : XOR2_X1 port map( A1 => n8636, A2 => n10358, Z => n19558);
   U10377 : INV_X2 port map( I => n25, ZN => n27171);
   U10383 : INV_X2 port map( I => n17980, ZN => n27172);
   U10385 : XOR2_X1 port map( A1 => n3779, A2 => n3778, Z => n3843);
   U10387 : NAND2_X1 port map( A1 => n21344, A2 => n21347, ZN => n21345);
   U10388 : AND2_X1 port map( A1 => n25736, A2 => n27173, Z => n6493);
   U10389 : NAND2_X2 port map( A1 => n18932, A2 => n11874, ZN => n18847);
   U10390 : NAND2_X2 port map( A1 => n11344, A2 => n1152, ZN => n9374);
   U10393 : NAND2_X2 port map( A1 => n9376, A2 => n18914, ZN => n11344);
   U10395 : NOR2_X2 port map( A1 => n27174, A2 => n13972, ZN => n25704);
   U10400 : NOR2_X2 port map( A1 => n27942, A2 => n27941, ZN => n27174);
   U10411 : NAND2_X2 port map( A1 => n21534, A2 => n27389, ZN => n6798);
   U10412 : XOR2_X1 port map( A1 => n13382, A2 => n19375, Z => n19310);
   U10415 : NAND2_X2 port map( A1 => n10756, A2 => n13594, ZN => n13382);
   U10417 : XOR2_X1 port map( A1 => n19358, A2 => n19457, Z => n28336);
   U10418 : XOR2_X1 port map( A1 => n24202, A2 => n22267, Z => n24522);
   U10420 : XOR2_X1 port map( A1 => n27176, A2 => n21085, Z => Ciphertext(88));
   U10422 : NAND2_X1 port map( A1 => n3319, A2 => n6883, ZN => n27176);
   U10425 : NOR2_X1 port map( A1 => n482, A2 => n4158, ZN => n23436);
   U10431 : NAND2_X2 port map( A1 => n25319, A2 => n27175, ZN => n15704);
   U10436 : XOR2_X1 port map( A1 => n16928, A2 => n28416, Z => n620);
   U10437 : NOR2_X2 port map( A1 => n27179, A2 => n25736, ZN => n15338);
   U10438 : NAND2_X2 port map( A1 => n25766, A2 => n14968, ZN => n27179);
   U10444 : OAI22_X1 port map( A1 => n21282, A2 => n21291, B1 => n21283, B2 => 
                           n21279, ZN => n27596);
   U10445 : NAND2_X1 port map( A1 => n6293, A2 => n8724, ZN => n27181);
   U10457 : OAI21_X1 port map( A1 => n943, A2 => n25298, B => n26156, ZN => 
                           n21992);
   U10459 : INV_X2 port map( I => n21271, ZN => n25298);
   U10460 : NAND2_X2 port map( A1 => n27182, A2 => n12247, ZN => n11389);
   U10462 : NAND2_X2 port map( A1 => n5388, A2 => n1113, ZN => n27182);
   U10467 : AND2_X1 port map( A1 => n6485, A2 => n26649, Z => n7107);
   U10474 : NAND2_X2 port map( A1 => n2231, A2 => n22779, ZN => n20139);
   U10477 : INV_X2 port map( I => n8012, ZN => n15067);
   U10482 : XOR2_X1 port map( A1 => n27183, A2 => n21320, Z => n15007);
   U10485 : XOR2_X1 port map( A1 => n28502, A2 => n21318, Z => n27183);
   U10495 : XOR2_X1 port map( A1 => n23238, A2 => n16842, Z => n8793);
   U10496 : AOI22_X2 port map( A1 => n989, A2 => n4702, B1 => n13812, B2 => 
                           n4705, ZN => n8052);
   U10498 : AOI21_X2 port map( A1 => n1982, A2 => n5874, B => n23861, ZN => 
                           n1977);
   U10499 : OAI21_X2 port map( A1 => n28040, A2 => n20898, B => n20902, ZN => 
                           n26006);
   U10501 : NAND2_X2 port map( A1 => n27184, A2 => n23914, ZN => n20393);
   U10505 : OAI21_X2 port map( A1 => n21808, A2 => n23912, B => n14179, ZN => 
                           n27184);
   U10512 : NAND2_X2 port map( A1 => n28547, A2 => n18999, ZN => n7609);
   U10513 : OAI21_X2 port map( A1 => n1882, A2 => n9304, B => n17929, ZN => 
                           n13185);
   U10515 : XOR2_X1 port map( A1 => n26246, A2 => n17125, Z => n26093);
   U10523 : NAND2_X2 port map( A1 => n6564, A2 => n6565, ZN => n26246);
   U10529 : BUF_X4 port map( I => n25270, Z => n28464);
   U10530 : INV_X2 port map( I => n7256, ZN => n18206);
   U10544 : XOR2_X1 port map( A1 => n12439, A2 => n7256, Z => n10914);
   U10546 : AOI21_X2 port map( A1 => n26630, A2 => n27186, B => n27185, ZN => 
                           n7256);
   U10547 : XOR2_X1 port map( A1 => n18084, A2 => n18181, Z => n12258);
   U10548 : XOR2_X1 port map( A1 => n18353, A2 => n18040, Z => n18181);
   U10550 : XOR2_X1 port map( A1 => n27188, A2 => n27187, Z => n10815);
   U10558 : XOR2_X1 port map( A1 => n18191, A2 => n7625, Z => n27187);
   U10559 : XOR2_X1 port map( A1 => n18053, A2 => n18293, Z => n27188);
   U10561 : XOR2_X1 port map( A1 => n14336, A2 => n16796, Z => n17180);
   U10562 : XOR2_X1 port map( A1 => n3869, A2 => n1094, Z => n274);
   U10564 : XOR2_X1 port map( A1 => n23686, A2 => n21364, Z => n3382);
   U10565 : XOR2_X1 port map( A1 => n19199, A2 => n2457, Z => n25900);
   U10573 : AOI22_X2 port map( A1 => n24597, A2 => n4822, B1 => n20625, B2 => 
                           n15287, ZN => n20627);
   U10574 : NAND3_X2 port map( A1 => n13036, A2 => n7043, A3 => n6651, ZN => 
                           n13056);
   U10586 : AOI21_X2 port map( A1 => n25910, A2 => n24390, B => n28523, ZN => 
                           n4711);
   U10588 : XOR2_X1 port map( A1 => n22847, A2 => n19526, Z => n3456);
   U10601 : XOR2_X1 port map( A1 => n24528, A2 => n4175, Z => n22847);
   U10608 : NAND2_X2 port map( A1 => n22263, A2 => n27189, ZN => n17926);
   U10624 : XOR2_X1 port map( A1 => n27190, A2 => n14360, Z => Ciphertext(96));
   U10658 : NOR2_X2 port map( A1 => n26651, A2 => n15697, ZN => n21361);
   U10666 : XOR2_X1 port map( A1 => n22831, A2 => n13793, Z => n9369);
   U10697 : BUF_X4 port map( I => n21788, Z => n27202);
   U10725 : NAND2_X1 port map( A1 => n27592, A2 => n27336, ZN => n22144);
   U10733 : XOR2_X1 port map( A1 => n27191, A2 => n20692, Z => Ciphertext(25));
   U10735 : NAND3_X1 port map( A1 => n22221, A2 => n3756, A3 => n3755, ZN => 
                           n27191);
   U10736 : AOI22_X2 port map( A1 => n8923, A2 => n1269, B1 => n4841, B2 => 
                           n4926, ZN => n7661);
   U10737 : NOR2_X2 port map( A1 => n8926, A2 => n16120, ZN => n4841);
   U10738 : AOI22_X2 port map( A1 => n10132, A2 => n8658, B1 => n27192, B2 => 
                           n17943, ZN => n10135);
   U10741 : INV_X1 port map( I => n10131, ZN => n27192);
   U10746 : AND2_X1 port map( A1 => n391, A2 => n26312, Z => n2736);
   U10747 : INV_X2 port map( I => n22349, ZN => n980);
   U10748 : XOR2_X1 port map( A1 => n315, A2 => n18111, Z => n18366);
   U10751 : NOR2_X2 port map( A1 => n25894, A2 => n27965, ZN => n27790);
   U10754 : INV_X2 port map( I => n19191, ZN => n27965);
   U10757 : NOR2_X2 port map( A1 => n18616, A2 => n8697, ZN => n19191);
   U10759 : XOR2_X1 port map( A1 => n27193, A2 => n21037, Z => Ciphertext(79));
   U10761 : XOR2_X1 port map( A1 => n18129, A2 => n13468, Z => n14709);
   U10762 : NAND3_X1 port map( A1 => n1112, A2 => n5931, A3 => n10151, ZN => 
                           n20001);
   U10763 : NAND2_X2 port map( A1 => n4739, A2 => n27194, ZN => n20332);
   U10770 : XOR2_X1 port map( A1 => n26342, A2 => n24741, Z => n25450);
   U10775 : NAND2_X2 port map( A1 => n847, A2 => n26913, ZN => n26011);
   U10780 : XOR2_X1 port map( A1 => n27196, A2 => n3869, Z => n22674);
   U10781 : NOR2_X2 port map( A1 => n1358, A2 => n1357, ZN => n3869);
   U10782 : XOR2_X1 port map( A1 => n21235, A2 => n14558, Z => n27196);
   U10785 : XOR2_X1 port map( A1 => n17138, A2 => n14058, Z => n25428);
   U10786 : AOI21_X1 port map( A1 => n21023, A2 => n21043, B => n21035, ZN => 
                           n21032);
   U10787 : XNOR2_X1 port map( A1 => n6218, A2 => n5398, ZN => n28377);
   U10788 : NOR2_X2 port map( A1 => n18810, A2 => n23126, ZN => n18934);
   U10790 : NAND2_X2 port map( A1 => n10673, A2 => n17956, ZN => n13615);
   U10793 : OR2_X1 port map( A1 => n14450, A2 => n21501, Z => n5171);
   U10802 : OR2_X1 port map( A1 => n19720, A2 => n12467, Z => n19824);
   U10803 : XNOR2_X1 port map( A1 => n10749, A2 => n11550, ZN => n10501);
   U10804 : XOR2_X1 port map( A1 => n12697, A2 => n19071, Z => n11550);
   U10805 : NAND2_X2 port map( A1 => n28328, A2 => n28327, ZN => n27198);
   U10806 : XOR2_X1 port map( A1 => n16945, A2 => n16946, Z => n16948);
   U10807 : XOR2_X1 port map( A1 => n15637, A2 => n1237, Z => n16946);
   U10810 : NAND2_X2 port map( A1 => n20804, A2 => n20803, ZN => n20801);
   U10813 : AOI21_X2 port map( A1 => n27227, A2 => n14991, B => n27197, ZN => 
                           n20105);
   U10816 : OAI21_X1 port map( A1 => n26852, A2 => n26081, B => n17514, ZN => 
                           n24878);
   U10819 : NAND2_X2 port map( A1 => n4898, A2 => n14792, ZN => n17740);
   U10826 : XOR2_X1 port map( A1 => n10202, A2 => n27364, Z => n3663);
   U10827 : NAND2_X2 port map( A1 => n8895, A2 => n8893, ZN => n10202);
   U10828 : NAND2_X1 port map( A1 => n25297, A2 => n23017, ZN => n27938);
   U10829 : INV_X2 port map( I => n27199, ZN => n25497);
   U10832 : XOR2_X1 port map( A1 => n16768, A2 => n9027, Z => n27199);
   U10833 : BUF_X2 port map( I => n8199, Z => n27200);
   U10834 : INV_X2 port map( I => n12042, ZN => n21979);
   U10836 : XOR2_X1 port map( A1 => n18097, A2 => n18147, Z => n18129);
   U10838 : NOR2_X2 port map( A1 => n5753, A2 => n28014, ZN => n13352);
   U10839 : NAND2_X2 port map( A1 => n5936, A2 => n10013, ZN => n7533);
   U10841 : NAND2_X2 port map( A1 => n2445, A2 => n22518, ZN => n9923);
   U10844 : XOR2_X1 port map( A1 => n19493, A2 => n19323, Z => n24910);
   U10845 : XOR2_X1 port map( A1 => n10828, A2 => n19462, Z => n19323);
   U10847 : XOR2_X1 port map( A1 => n27203, A2 => n21570, Z => Ciphertext(155))
                           ;
   U10848 : AOI22_X1 port map( A1 => n9220, A2 => n22732, B1 => n24574, B2 => 
                           n21569, ZN => n27203);
   U10850 : BUF_X2 port map( I => n755, Z => n27204);
   U10852 : INV_X2 port map( I => n10488, ZN => n3255);
   U10853 : NOR3_X2 port map( A1 => n27206, A2 => n27205, A3 => n5639, ZN => 
                           n27973);
   U10854 : NOR2_X1 port map( A1 => n17513, A2 => n26081, ZN => n27205);
   U10855 : NOR2_X2 port map( A1 => n24018, A2 => n26628, ZN => n27206);
   U10863 : NOR2_X2 port map( A1 => n5805, A2 => n18776, ZN => n11280);
   U10864 : NAND2_X2 port map( A1 => n18535, A2 => n4410, ZN => n5805);
   U10865 : NAND3_X2 port map( A1 => n1185, A2 => n18698, A3 => n18610, ZN => 
                           n27207);
   U10866 : OAI21_X2 port map( A1 => n15718, A2 => n11196, B => n11197, ZN => 
                           n10842);
   U10868 : XOR2_X1 port map( A1 => n24095, A2 => n21421, Z => n15372);
   U10874 : AND3_X1 port map( A1 => n20186, A2 => n11961, A3 => n5931, Z => 
                           n27215);
   U10875 : NOR2_X2 port map( A1 => n3121, A2 => n27208, ZN => n24787);
   U10879 : NOR3_X1 port map( A1 => n972, A2 => n27905, A3 => n19748, ZN => 
                           n27208);
   U10882 : NAND2_X1 port map( A1 => n11001, A2 => n27209, ZN => n22060);
   U10884 : NAND3_X1 port map( A1 => n26422, A2 => n8672, A3 => n21711, ZN => 
                           n27209);
   U10893 : NOR2_X1 port map( A1 => n23624, A2 => n12682, ZN => n10493);
   U10895 : XOR2_X1 port map( A1 => n27210, A2 => n18109, Z => n4055);
   U10898 : XOR2_X1 port map( A1 => n24363, A2 => n22135, Z => n27210);
   U10899 : AND2_X1 port map( A1 => n13472, A2 => n21124, Z => n27579);
   U10900 : NAND2_X2 port map( A1 => n17894, A2 => n22253, ZN => n27211);
   U10903 : XOR2_X1 port map( A1 => n20446, A2 => n27212, Z => n21063);
   U10904 : XOR2_X1 port map( A1 => n22402, A2 => n2319, Z => n27212);
   U10905 : NOR2_X2 port map( A1 => n1684, A2 => n1683, ZN => n20072);
   U10908 : XOR2_X1 port map( A1 => n27767, A2 => n20480, Z => n21201);
   U10909 : NOR2_X2 port map( A1 => n17491, A2 => n14504, ZN => n3839);
   U10911 : AOI22_X2 port map( A1 => n17363, A2 => n17362, B1 => n17489, B2 => 
                           n25971, ZN => n17491);
   U10912 : INV_X2 port map( I => n5511, ZN => n1149);
   U10914 : XOR2_X1 port map( A1 => n538, A2 => n17095, Z => n22313);
   U10919 : XOR2_X1 port map( A1 => n2850, A2 => n9902, Z => n17095);
   U10922 : NAND2_X1 port map( A1 => n21087, A2 => n6473, ZN => n27213);
   U10924 : NOR2_X2 port map( A1 => n19110, A2 => n28547, ZN => n19113);
   U10925 : AOI22_X1 port map( A1 => n2271, A2 => n27862, B1 => n17586, B2 => 
                           n8882, ZN => n27845);
   U10929 : XOR2_X1 port map( A1 => n21784, A2 => n451, Z => n640);
   U10930 : NOR2_X2 port map( A1 => n454, A2 => n15646, ZN => n3096);
   U10934 : OR2_X1 port map( A1 => n18426, A2 => n19147, Z => n10159);
   U10939 : NOR3_X2 port map( A1 => n27215, A2 => n24173, A3 => n27214, ZN => 
                           n24172);
   U10940 : XOR2_X1 port map( A1 => n27216, A2 => n1318, Z => Ciphertext(32));
   U10943 : OAI22_X1 port map( A1 => n6054, A2 => n6053, B1 => n20743, B2 => 
                           n20749, ZN => n27216);
   U10944 : AND2_X1 port map( A1 => n27419, A2 => n26882, Z => n21549);
   U10947 : OAI21_X1 port map( A1 => n6485, A2 => n26649, B => n21080, ZN => 
                           n9864);
   U10948 : INV_X2 port map( I => n7126, ZN => n370);
   U10949 : OAI21_X2 port map( A1 => n18893, A2 => n22967, B => n26503, ZN => 
                           n7126);
   U10950 : AOI21_X2 port map( A1 => n9450, A2 => n12477, B => n20125, ZN => 
                           n8268);
   U10961 : INV_X2 port map( I => n2544, ZN => n25465);
   U10962 : NAND2_X2 port map( A1 => n10920, A2 => n10566, ZN => n26356);
   U10967 : NOR2_X2 port map( A1 => n25828, A2 => n18752, ZN => n10267);
   U10969 : INV_X2 port map( I => n27218, ZN => n19008);
   U10970 : AOI21_X2 port map( A1 => n5320, A2 => n15142, B => n15143, ZN => 
                           n27218);
   U10973 : BUF_X4 port map( I => n7652, Z => n25542);
   U10976 : NAND2_X1 port map( A1 => n26551, A2 => n23929, ZN => n12847);
   U10977 : NAND2_X2 port map( A1 => n10764, A2 => n14213, ZN => n20329);
   U10979 : BUF_X2 port map( I => n7134, Z => n27219);
   U10987 : NAND3_X2 port map( A1 => n27220, A2 => n21324, A3 => n25739, ZN => 
                           n22990);
   U10989 : NAND2_X1 port map( A1 => n21325, A2 => n21278, ZN => n27220);
   U10992 : XOR2_X1 port map( A1 => n27221, A2 => n14505, Z => Ciphertext(111))
                           ;
   U10994 : XOR2_X1 port map( A1 => n27222, A2 => n20949, Z => Ciphertext(62));
   U10995 : NAND2_X1 port map( A1 => n14466, A2 => n14465, ZN => n27222);
   U10997 : BUF_X4 port map( I => n5305, Z => n25);
   U11001 : OR2_X1 port map( A1 => n21924, A2 => n20921, Z => n5798);
   U11003 : NAND2_X1 port map( A1 => n22905, A2 => n1003, ZN => n27552);
   U11009 : AOI21_X2 port map( A1 => n17228, A2 => n23787, B => n27223, ZN => 
                           n22202);
   U11011 : AOI21_X2 port map( A1 => n13319, A2 => n23019, B => n17185, ZN => 
                           n27223);
   U11013 : NOR2_X2 port map( A1 => n944, A2 => n25298, ZN => n12310);
   U11017 : OAI22_X2 port map( A1 => n8950, A2 => n8951, B1 => n8949, B2 => 
                           n4657, ZN => n28266);
   U11026 : OAI21_X2 port map( A1 => n10046, A2 => n26255, B => n27224, ZN => 
                           n8174);
   U11027 : NAND2_X2 port map( A1 => n26255, A2 => n898, ZN => n27224);
   U11028 : NOR2_X1 port map( A1 => n18608, A2 => n11452, ZN => n7080);
   U11034 : AOI21_X2 port map( A1 => n28122, A2 => n17638, B => n17822, ZN => 
                           n8535);
   U11036 : NOR2_X2 port map( A1 => n2084, A2 => n22965, ZN => n6423);
   U11038 : NAND2_X1 port map( A1 => n25318, A2 => n20618, ZN => n13622);
   U11040 : NAND2_X1 port map( A1 => n2622, A2 => n22522, ZN => n25318);
   U11045 : INV_X2 port map( I => n7326, ZN => n27445);
   U11047 : OAI21_X1 port map( A1 => n1410, A2 => n8197, B => n14663, ZN => 
                           n27475);
   U11051 : NAND3_X1 port map( A1 => n22338, A2 => n25586, A3 => n19163, ZN => 
                           n27225);
   U11057 : XOR2_X1 port map( A1 => n27226, A2 => n1301, Z => Ciphertext(68));
   U11058 : AOI22_X1 port map( A1 => n27570, A2 => n27571, B1 => n1825, B2 => 
                           n928, ZN => n27226);
   U11060 : BUF_X2 port map( I => n22598, Z => n27227);
   U11061 : NAND2_X2 port map( A1 => n26668, A2 => n1130, ZN => n6981);
   U11062 : INV_X2 port map( I => n27228, ZN => n13121);
   U11068 : XOR2_X1 port map( A1 => n10201, A2 => n27789, Z => n27228);
   U11072 : NAND2_X2 port map( A1 => n26627, A2 => n21059, ZN => n26220);
   U11073 : NAND2_X1 port map( A1 => n26219, A2 => n26221, ZN => n11018);
   U11075 : INV_X1 port map( I => n13121, ZN => n25614);
   U11077 : NAND2_X2 port map( A1 => n27229, A2 => n23889, ZN => n28472);
   U11078 : NAND2_X2 port map( A1 => n18409, A2 => n22031, ZN => n27229);
   U11079 : NAND2_X2 port map( A1 => n27230, A2 => n25449, ZN => n17751);
   U11080 : NAND3_X2 port map( A1 => n27231, A2 => n4668, A3 => n23264, ZN => 
                           n6959);
   U11081 : OR2_X1 port map( A1 => n10061, A2 => n17992, Z => n10059);
   U11082 : OAI21_X2 port map( A1 => n17231, A2 => n14061, B => n27232, ZN => 
                           n17869);
   U11083 : AOI22_X2 port map( A1 => n10432, A2 => n25786, B1 => n10692, B2 => 
                           n17561, ZN => n27232);
   U11085 : NOR2_X2 port map( A1 => n27200, A2 => n27989, ZN => n16376);
   U11089 : NOR2_X2 port map( A1 => n1271, A2 => n12272, ZN => n15866);
   U11098 : NAND2_X1 port map( A1 => n27233, A2 => n25961, ZN => n20940);
   U11101 : NAND2_X1 port map( A1 => n25963, A2 => n1072, ZN => n27233);
   U11102 : XOR2_X1 port map( A1 => n6384, A2 => n6386, Z => n28075);
   U11104 : INV_X2 port map( I => n27234, ZN => n23004);
   U11105 : XNOR2_X1 port map( A1 => n8681, A2 => n8682, ZN => n27234);
   U11106 : NAND2_X2 port map( A1 => n18836, A2 => n28216, ZN => n8657);
   U11108 : NAND3_X1 port map( A1 => n27235, A2 => n25959, A3 => n20277, ZN => 
                           n10631);
   U11109 : OR2_X2 port map( A1 => n1995, A2 => n8937, Z => n9361);
   U11110 : XOR2_X1 port map( A1 => n1743, A2 => n1741, Z => n1995);
   U11111 : NAND2_X2 port map( A1 => n7890, A2 => n12463, ZN => n21455);
   U11114 : AOI22_X2 port map( A1 => n21511, A2 => n21543, B1 => n21513, B2 => 
                           n21440, ZN => n7890);
   U11115 : NAND3_X1 port map( A1 => n3736, A2 => n6683, A3 => n6879, ZN => 
                           n25086);
   U11116 : INV_X2 port map( I => n27237, ZN => n18739);
   U11126 : XNOR2_X1 port map( A1 => n27533, A2 => n9241, ZN => n27237);
   U11133 : INV_X2 port map( I => n14456, ZN => n3771);
   U11135 : INV_X2 port map( I => n27238, ZN => n2404);
   U11139 : XOR2_X1 port map( A1 => Plaintext(29), A2 => Key(29), Z => n27238);
   U11144 : BUF_X2 port map( I => n16565, Z => n27239);
   U11149 : NOR2_X2 port map( A1 => n914, A2 => n27240, ZN => n15953);
   U11150 : INV_X2 port map( I => n338, ZN => n27240);
   U11153 : NAND2_X2 port map( A1 => n19640, A2 => n19641, ZN => n27667);
   U11155 : XOR2_X1 port map( A1 => n15221, A2 => n12233, Z => n7201);
   U11157 : BUF_X2 port map( I => n25609, Z => n27241);
   U11164 : OAI21_X2 port map( A1 => n15207, A2 => n14239, B => n28446, ZN => 
                           n12259);
   U11167 : NAND2_X1 port map( A1 => n27544, A2 => n28227, ZN => n6958);
   U11172 : INV_X2 port map( I => n17325, ZN => n15037);
   U11176 : XOR2_X1 port map( A1 => n1401, A2 => n27242, Z => n17325);
   U11178 : AOI21_X2 port map( A1 => n6354, A2 => n23653, B => n27618, ZN => 
                           n27617);
   U11183 : BUF_X2 port map( I => n17147, Z => n27243);
   U11187 : NAND2_X1 port map( A1 => n7912, A2 => n900, ZN => n4254);
   U11190 : AOI21_X2 port map( A1 => n15211, A2 => n15210, B => n27244, ZN => 
                           n12974);
   U11191 : OAI22_X1 port map( A1 => n15882, A2 => n7910, B1 => n2331, B2 => 
                           n16193, ZN => n27244);
   U11194 : BUF_X2 port map( I => n18205, Z => n27245);
   U11196 : NAND2_X2 port map( A1 => n16508, A2 => n1054, ZN => n23828);
   U11197 : NAND2_X2 port map( A1 => n16055, A2 => n16604, ZN => n16508);
   U11198 : XOR2_X1 port map( A1 => n23917, A2 => n19272, Z => n14002);
   U11203 : INV_X4 port map( I => n17546, ZN => n765);
   U11206 : XOR2_X1 port map( A1 => n25941, A2 => n19250, Z => n3615);
   U11207 : XOR2_X1 port map( A1 => n21240, A2 => n21241, Z => n84);
   U11212 : AOI21_X2 port map( A1 => n3766, A2 => n1167, B => n27246, ZN => 
                           n3764);
   U11215 : NOR2_X2 port map( A1 => n4883, A2 => n18455, ZN => n27246);
   U11220 : OAI21_X2 port map( A1 => n19596, A2 => n1128, B => n27247, ZN => 
                           n4191);
   U11221 : AOI22_X2 port map( A1 => n27844, A2 => n19847, B1 => n19846, B2 => 
                           n19595, ZN => n27247);
   U11222 : INV_X4 port map( I => n17518, ZN => n1029);
   U11223 : OR2_X1 port map( A1 => n25380, A2 => n7912, Z => n4250);
   U11229 : INV_X2 port map( I => n11789, ZN => n19965);
   U11234 : AND2_X2 port map( A1 => n11732, A2 => n12599, Z => n2469);
   U11239 : INV_X4 port map( I => n21724, ZN => n28027);
   U11241 : NAND2_X2 port map( A1 => n26287, A2 => n26288, ZN => n26055);
   U11244 : XOR2_X1 port map( A1 => n11999, A2 => n18115, Z => n6062);
   U11245 : XOR2_X1 port map( A1 => n18262, A2 => n1970, Z => n18115);
   U11249 : XOR2_X1 port map( A1 => n27249, A2 => n7725, Z => n17334);
   U11252 : XOR2_X1 port map( A1 => n7729, A2 => n15097, Z => n27249);
   U11253 : NOR3_X1 port map( A1 => n1214, A2 => n3929, A3 => n17724, ZN => 
                           n26266);
   U11259 : NAND2_X2 port map( A1 => n17712, A2 => n24807, ZN => n24155);
   U11260 : NAND2_X2 port map( A1 => n21998, A2 => n27029, ZN => n17712);
   U11266 : NAND2_X2 port map( A1 => n2167, A2 => n27250, ZN => n26319);
   U11267 : NOR2_X2 port map( A1 => n27252, A2 => n27251, ZN => n27250);
   U11270 : NOR2_X1 port map( A1 => n14502, A2 => n24190, ZN => n27251);
   U11272 : INV_X2 port map( I => n14925, ZN => n27252);
   U11274 : NOR2_X2 port map( A1 => n5707, A2 => n14459, ZN => n19862);
   U11277 : INV_X2 port map( I => n19649, ZN => n5707);
   U11279 : NOR3_X2 port map( A1 => n26212, A2 => n26703, A3 => n21965, ZN => 
                           n8630);
   U11280 : NAND2_X2 port map( A1 => n27253, A2 => n23167, ZN => n20339);
   U11284 : NAND2_X1 port map( A1 => n19745, A2 => n10557, ZN => n27253);
   U11285 : AND3_X1 port map( A1 => n16700, A2 => n10868, A3 => n27572, Z => 
                           n1422);
   U11286 : XOR2_X1 port map( A1 => n18099, A2 => n27254, Z => n18282);
   U11289 : NAND2_X1 port map( A1 => n14169, A2 => n2209, ZN => n2208);
   U11290 : INV_X1 port map( I => n27574, ZN => n21753);
   U11292 : OR2_X1 port map( A1 => n27574, A2 => n17941, Z => n17945);
   U11300 : AOI21_X1 port map( A1 => n4328, A2 => n27407, B => n4326, ZN => 
                           n27892);
   U11306 : INV_X2 port map( I => n27255, ZN => n6672);
   U11308 : XNOR2_X1 port map( A1 => n6673, A2 => n4524, ZN => n27255);
   U11310 : NAND2_X2 port map( A1 => n3398, A2 => n4824, ZN => n19498);
   U11311 : XOR2_X1 port map( A1 => n7413, A2 => n13891, Z => n12146);
   U11312 : NAND2_X2 port map( A1 => n15682, A2 => n15681, ZN => n7413);
   U11315 : AND2_X1 port map( A1 => n18557, A2 => n27436, Z => n3697);
   U11317 : NOR2_X2 port map( A1 => n8837, A2 => n8835, ZN => n27256);
   U11321 : XOR2_X1 port map( A1 => n16780, A2 => n14675, Z => n2236);
   U11323 : XOR2_X1 port map( A1 => n16950, A2 => n3477, Z => n16780);
   U11327 : AND2_X1 port map( A1 => n21062, A2 => n15729, Z => n27270);
   U11331 : XOR2_X1 port map( A1 => n20510, A2 => n20509, Z => n5755);
   U11332 : INV_X1 port map( I => n28110, ZN => n27583);
   U11334 : AOI21_X2 port map( A1 => n974, A2 => n13387, B => n19830, ZN => 
                           n27257);
   U11336 : NAND2_X1 port map( A1 => n26669, A2 => n10210, ZN => n6410);
   U11341 : AND2_X1 port map( A1 => n25368, A2 => n19150, Z => n22471);
   U11342 : XOR2_X1 port map( A1 => n27259, A2 => n4183, Z => n7966);
   U11343 : XOR2_X1 port map( A1 => n4184, A2 => n18128, Z => n27259);
   U11351 : OAI21_X2 port map( A1 => n17862, A2 => n713, B => n17861, ZN => 
                           n17866);
   U11361 : NOR2_X2 port map( A1 => n25607, A2 => n26312, ZN => n17862);
   U11367 : INV_X4 port map( I => n4790, ZN => n20171);
   U11368 : NAND2_X2 port map( A1 => n27990, A2 => n6548, ZN => n4790);
   U11372 : OAI22_X2 port map( A1 => n27261, A2 => n27260, B1 => n20588, B2 => 
                           n8823, ZN => n12235);
   U11375 : NAND2_X2 port map( A1 => n24170, A2 => n21915, ZN => n18936);
   U11378 : XOR2_X1 port map( A1 => n21181, A2 => n20529, Z => n2367);
   U11380 : XOR2_X1 port map( A1 => n26537, A2 => n12533, Z => n20529);
   U11382 : AOI22_X2 port map( A1 => n19627, A2 => n19754, B1 => n26382, B2 => 
                           n19626, ZN => n24245);
   U11383 : NAND3_X1 port map( A1 => n27056, A2 => n27458, A3 => n23923, ZN => 
                           n17689);
   U11384 : XOR2_X1 port map( A1 => n22802, A2 => n21262, Z => n27262);
   U11390 : NAND2_X2 port map( A1 => n17761, A2 => n13235, ZN => n17964);
   U11391 : NAND3_X2 port map( A1 => n24594, A2 => n2047, A3 => n27263, ZN => 
                           n6687);
   U11392 : XOR2_X1 port map( A1 => n2467, A2 => n22793, Z => n27292);
   U11393 : NAND2_X2 port map( A1 => n11154, A2 => n11155, ZN => n22793);
   U11394 : INV_X2 port map( I => n17084, ZN => n17025);
   U11397 : OR2_X1 port map( A1 => n14975, A2 => n23817, Z => n23954);
   U11402 : NAND2_X2 port map( A1 => n18873, A2 => n26831, ZN => n18875);
   U11404 : NAND2_X2 port map( A1 => n27264, A2 => n5141, ZN => n1455);
   U11405 : INV_X2 port map( I => n20263, ZN => n27265);
   U11406 : INV_X2 port map( I => n12287, ZN => n27266);
   U11417 : XOR2_X1 port map( A1 => n18227, A2 => n20396, Z => n5090);
   U11418 : NOR2_X2 port map( A1 => n10211, A2 => n26364, ZN => n18227);
   U11420 : XOR2_X1 port map( A1 => n27267, A2 => n12277, Z => n3216);
   U11421 : INV_X2 port map( I => n27268, ZN => n19908);
   U11426 : NAND4_X2 port map( A1 => n19912, A2 => n19911, A3 => n27479, A4 => 
                           n27268, ZN => n24533);
   U11430 : NAND2_X2 port map( A1 => n26654, A2 => n26948, ZN => n27268);
   U11431 : NAND3_X1 port map( A1 => n25256, A2 => n21121, A3 => n7313, ZN => 
                           n27504);
   U11432 : INV_X4 port map( I => n6672, ZN => n17490);
   U11433 : XOR2_X1 port map( A1 => n27358, A2 => n19305, Z => n23638);
   U11434 : NAND2_X2 port map( A1 => n11997, A2 => n11996, ZN => n27358);
   U11438 : XOR2_X1 port map( A1 => n2914, A2 => n26718, Z => n2912);
   U11440 : NAND2_X2 port map( A1 => n11425, A2 => n14683, ZN => n14417);
   U11442 : NAND2_X1 port map( A1 => n22517, A2 => n11499, ZN => n28374);
   U11446 : NOR2_X1 port map( A1 => n28374, A2 => n23205, ZN => n23204);
   U11453 : XOR2_X1 port map( A1 => n27269, A2 => n28342, Z => Ciphertext(137))
                           ;
   U11454 : AOI22_X1 port map( A1 => n13798, A2 => n23579, B1 => n27866, B2 => 
                           n13799, ZN => n27269);
   U11455 : XOR2_X1 port map( A1 => n6523, A2 => n6996, Z => n25174);
   U11456 : XOR2_X1 port map( A1 => n5283, A2 => n8490, Z => n27416);
   U11459 : XOR2_X1 port map( A1 => n8488, A2 => n8489, Z => n5283);
   U11462 : XOR2_X1 port map( A1 => n19250, A2 => n6275, Z => n12948);
   U11463 : NOR2_X2 port map( A1 => n14272, A2 => n18966, ZN => n19250);
   U11464 : OAI21_X2 port map( A1 => n11334, A2 => n6861, B => n19731, ZN => 
                           n8387);
   U11465 : INV_X1 port map( I => n25173, ZN => n27271);
   U11467 : NAND3_X2 port map( A1 => n3293, A2 => n21102, A3 => n27272, ZN => 
                           n24858);
   U11468 : AOI22_X1 port map( A1 => n11521, A2 => n21113, B1 => n11522, B2 => 
                           n13021, ZN => n27272);
   U11469 : XOR2_X1 port map( A1 => n11098, A2 => n27273, Z => n12286);
   U11470 : XOR2_X1 port map( A1 => n11253, A2 => n19409, Z => n27273);
   U11472 : XOR2_X1 port map( A1 => n19253, A2 => n19252, Z => n19254);
   U11474 : NAND3_X2 port map( A1 => n8493, A2 => n3132, A3 => n7000, ZN => 
                           n28176);
   U11477 : XNOR2_X1 port map( A1 => n18133, A2 => n18158, ZN => n27274);
   U11479 : BUF_X4 port map( I => n24283, Z => n27345);
   U11483 : XOR2_X1 port map( A1 => n698, A2 => n1309, Z => n5314);
   U11484 : NAND2_X2 port map( A1 => n23776, A2 => n4613, ZN => n698);
   U11489 : XOR2_X1 port map( A1 => n3597, A2 => n27274, Z => n25609);
   U11491 : INV_X2 port map( I => n26647, ZN => n26092);
   U11492 : OAI21_X2 port map( A1 => n14565, A2 => n19658, B => n8754, ZN => 
                           n8950);
   U11494 : NOR2_X1 port map( A1 => n8934, A2 => n23484, ZN => n27275);
   U11495 : XNOR2_X1 port map( A1 => n20770, A2 => n20489, ZN => n2201);
   U11499 : XOR2_X1 port map( A1 => n27352, A2 => n13437, Z => n4026);
   U11501 : NAND3_X2 port map( A1 => n24449, A2 => n4028, A3 => n24450, ZN => 
                           n13437);
   U11507 : OR2_X1 port map( A1 => n20078, A2 => n19999, Z => n4269);
   U11509 : XOR2_X1 port map( A1 => n13916, A2 => n16746, Z => n11339);
   U11514 : AOI21_X2 port map( A1 => n12329, A2 => n10710, B => n12328, ZN => 
                           n13916);
   U11515 : XOR2_X1 port map( A1 => n8776, A2 => n10773, Z => n17029);
   U11519 : NAND2_X2 port map( A1 => n25626, A2 => n12214, ZN => n8776);
   U11524 : AND2_X1 port map( A1 => n15859, A2 => n26434, Z => n16164);
   U11525 : BUF_X2 port map( I => n18798, Z => n23672);
   U11530 : NAND2_X2 port map( A1 => n7478, A2 => n26694, ZN => n23905);
   U11538 : XOR2_X1 port map( A1 => n15537, A2 => n13834, Z => n11811);
   U11543 : NAND2_X2 port map( A1 => n23617, A2 => n22696, ZN => n15537);
   U11544 : NAND3_X2 port map( A1 => n22494, A2 => n17750, A3 => n12590, ZN => 
                           n15682);
   U11546 : NOR3_X2 port map( A1 => n8935, A2 => n5195, A3 => n14750, ZN => 
                           n23484);
   U11547 : INV_X2 port map( I => n26647, ZN => n21739);
   U11551 : NOR3_X1 port map( A1 => n13467, A2 => n18687, A3 => n5523, ZN => 
                           n27278);
   U11553 : XOR2_X1 port map( A1 => n19377, A2 => n22768, Z => n3862);
   U11554 : NAND2_X2 port map( A1 => n3480, A2 => n22746, ZN => n19377);
   U11556 : NAND2_X2 port map( A1 => n14750, A2 => n5578, ZN => n6433);
   U11561 : NAND2_X2 port map( A1 => n9894, A2 => n26647, ZN => n8771);
   U11563 : NAND2_X1 port map( A1 => n12465, A2 => n7354, ZN => n27998);
   U11567 : XOR2_X1 port map( A1 => n356, A2 => n27585, Z => n7354);
   U11568 : XOR2_X1 port map( A1 => n20038, A2 => n20488, Z => n21320);
   U11571 : NAND3_X2 port map( A1 => n22679, A2 => n20037, A3 => n20036, ZN => 
                           n20488);
   U11572 : NAND2_X1 port map( A1 => n26553, A2 => n26552, ZN => n28427);
   U11574 : XOR2_X1 port map( A1 => n27280, A2 => n14640, Z => Ciphertext(124))
                           ;
   U11575 : NAND2_X2 port map( A1 => n27282, A2 => n26160, ZN => n3496);
   U11577 : XOR2_X1 port map( A1 => n10369, A2 => n5517, Z => n21548);
   U11583 : XOR2_X1 port map( A1 => n27283, A2 => n23576, Z => n25503);
   U11589 : NAND2_X1 port map( A1 => n25161, A2 => n15502, ZN => n27284);
   U11593 : XOR2_X1 port map( A1 => n28222, A2 => n21185, Z => n27285);
   U11595 : XOR2_X1 port map( A1 => n19340, A2 => n11004, Z => n6274);
   U11599 : XOR2_X1 port map( A1 => n6273, A2 => n6275, Z => n19340);
   U11600 : NOR2_X2 port map( A1 => n24998, A2 => n19978, ZN => n28002);
   U11601 : NAND2_X2 port map( A1 => n28002, A2 => n27286, ZN => n24677);
   U11602 : INV_X2 port map( I => n17291, ZN => n27287);
   U11609 : NAND2_X2 port map( A1 => n10580, A2 => n26198, ZN => n17291);
   U11610 : AOI22_X2 port map( A1 => n4881, A2 => n1987, B1 => n13742, B2 => 
                           n4750, ZN => n4880);
   U11611 : AND2_X1 port map( A1 => n18597, A2 => n4679, Z => n12671);
   U11613 : NAND2_X2 port map( A1 => n21722, A2 => n21721, ZN => n6338);
   U11614 : NAND2_X2 port map( A1 => n6415, A2 => n17664, ZN => n3695);
   U11616 : NOR2_X1 port map( A1 => n28300, A2 => n13050, ZN => n9004);
   U11617 : NOR2_X1 port map( A1 => n21736, A2 => n21735, ZN => n26326);
   U11624 : XOR2_X1 port map( A1 => n27289, A2 => n5212, Z => n1527);
   U11625 : XOR2_X1 port map( A1 => n3, A2 => n15038, Z => n27289);
   U11632 : OR2_X1 port map( A1 => n17927, A2 => n4814, Z => n17774);
   U11634 : OAI22_X2 port map( A1 => n19862, A2 => n19914, B1 => n12614, B2 => 
                           n204, ZN => n27990);
   U11636 : AOI21_X2 port map( A1 => n9446, A2 => n9264, B => n9175, ZN => 
                           n9447);
   U11637 : AOI22_X1 port map( A1 => n27315, A2 => n802, B1 => n11640, B2 => 
                           n22753, ZN => n27903);
   U11638 : NOR2_X2 port map( A1 => n27528, A2 => n14260, ZN => n5188);
   U11639 : INV_X2 port map( I => n15709, ZN => n14260);
   U11644 : XOR2_X1 port map( A1 => n2855, A2 => n9451, Z => n15709);
   U11647 : NAND2_X2 port map( A1 => n27330, A2 => n17755, ZN => n26364);
   U11648 : NOR2_X2 port map( A1 => n19101, A2 => n7018, ZN => n18991);
   U11653 : NAND2_X2 port map( A1 => n23428, A2 => n23302, ZN => n7018);
   U11655 : NAND2_X2 port map( A1 => n7566, A2 => n11059, ZN => n20564);
   U11656 : OAI21_X2 port map( A1 => n17296, A2 => n2966, B => n1229, ZN => 
                           n2566);
   U11660 : XOR2_X1 port map( A1 => n19404, A2 => n27292, Z => n7640);
   U11663 : NAND2_X2 port map( A1 => n17869, A2 => n7321, ZN => n6038);
   U11664 : BUF_X4 port map( I => n17202, Z => n17510);
   U11666 : XOR2_X1 port map( A1 => n19368, A2 => n8322, Z => n9656);
   U11669 : NAND3_X2 port map( A1 => n18993, A2 => n9657, A3 => n18992, ZN => 
                           n19368);
   U11672 : NAND3_X2 port map( A1 => n28392, A2 => n17272, A3 => n27293, ZN => 
                           n25214);
   U11674 : NOR3_X1 port map( A1 => n22385, A2 => n114, A3 => n28237, ZN => 
                           n8127);
   U11675 : XOR2_X1 port map( A1 => n22126, A2 => n275, Z => n633);
   U11679 : INV_X2 port map( I => n12034, ZN => n27376);
   U11680 : XOR2_X1 port map( A1 => n11768, A2 => n10075, Z => n10076);
   U11681 : XOR2_X1 port map( A1 => n7200, A2 => n16845, Z => n10075);
   U11682 : NOR2_X2 port map( A1 => n2213, A2 => n1541, ZN => n27294);
   U11686 : AOI22_X2 port map( A1 => n27295, A2 => n21759, B1 => n20249, B2 => 
                           n20141, ZN => n21386);
   U11687 : NAND2_X2 port map( A1 => n35, A2 => n26960, ZN => n27295);
   U11691 : NOR2_X1 port map( A1 => n27583, A2 => n27582, ZN => n22528);
   U11693 : XOR2_X1 port map( A1 => n25183, A2 => n11768, Z => n27296);
   U11696 : NAND3_X1 port map( A1 => n27552, A2 => n3215, A3 => n27440, ZN => 
                           n28171);
   U11699 : AND2_X1 port map( A1 => n4644, A2 => n27019, Z => n22908);
   U11700 : XOR2_X1 port map( A1 => n27297, A2 => n6983, Z => n7571);
   U11706 : XOR2_X1 port map( A1 => n17062, A2 => n28070, Z => n27297);
   U11707 : AOI22_X2 port map( A1 => n11402, A2 => n26154, B1 => n11398, B2 => 
                           n10764, ZN => n11401);
   U11708 : NAND2_X2 port map( A1 => n24188, A2 => n778, ZN => n10665);
   U11709 : BUF_X4 port map( I => n17996, Z => n27640);
   U11710 : AOI22_X2 port map( A1 => n27547, A2 => n25542, B1 => n4192, B2 => 
                           n1211, ZN => n25982);
   U11713 : NAND2_X2 port map( A1 => n21734, A2 => n21737, ZN => n21741);
   U11714 : NAND2_X2 port map( A1 => n27298, A2 => n4016, ZN => n7103);
   U11719 : AOI21_X1 port map( A1 => n4015, A2 => n4013, B => n24087, ZN => 
                           n27298);
   U11723 : BUF_X4 port map( I => n24147, Z => n26009);
   U11727 : XOR2_X1 port map( A1 => n16800, A2 => n16852, Z => n16804);
   U11732 : NAND2_X2 port map( A1 => n10422, A2 => n16433, ZN => n16410);
   U11738 : OAI21_X2 port map( A1 => n27299, A2 => n24371, B => n24335, ZN => 
                           n3976);
   U11740 : NOR2_X2 port map( A1 => n27300, A2 => n12490, ZN => n11138);
   U11746 : INV_X2 port map( I => n27301, ZN => n26615);
   U11750 : XOR2_X1 port map( A1 => n10396, A2 => n22347, Z => n27301);
   U11754 : NAND2_X1 port map( A1 => n19033, A2 => n8290, ZN => n6722);
   U11755 : XOR2_X1 port map( A1 => n3869, A2 => n27302, Z => n28041);
   U11756 : XOR2_X1 port map( A1 => n19414, A2 => n19493, Z => n10413);
   U11757 : XOR2_X1 port map( A1 => n19490, A2 => n12739, Z => n19414);
   U11758 : NAND2_X1 port map( A1 => n26773, A2 => n12287, ZN => n68);
   U11759 : XOR2_X1 port map( A1 => n11677, A2 => n27306, Z => n615);
   U11761 : XOR2_X1 port map( A1 => n12857, A2 => n26664, Z => n27306);
   U11762 : NOR2_X2 port map( A1 => n22312, A2 => n23542, ZN => n27307);
   U11765 : XOR2_X1 port map( A1 => n13497, A2 => n27308, Z => n17891);
   U11768 : XOR2_X1 port map( A1 => n23574, A2 => n9832, Z => n27308);
   U11776 : BUF_X4 port map( I => n12079, Z => n10963);
   U11778 : OR2_X1 port map( A1 => n19468, A2 => n3083, Z => n3099);
   U11779 : OAI21_X2 port map( A1 => n2804, A2 => n2805, B => n27309, ZN => 
                           n2800);
   U11782 : AOI22_X1 port map( A1 => n2802, A2 => n952, B1 => n5950, B2 => 
                           n5721, ZN => n27309);
   U11791 : BUF_X2 port map( I => n14961, Z => n23036);
   U11792 : NAND2_X2 port map( A1 => n6245, A2 => n27310, ZN => n6447);
   U11795 : AOI22_X2 port map( A1 => n18547, A2 => n2445, B1 => n18626, B2 => 
                           n18546, ZN => n27310);
   U11796 : AND2_X1 port map( A1 => n6881, A2 => n21082, Z => n27311);
   U11805 : AOI21_X2 port map( A1 => n19592, A2 => n19871, B => n27312, ZN => 
                           n20064);
   U11806 : AOI21_X2 port map( A1 => n28192, A2 => n28193, B => n6503, ZN => 
                           n6502);
   U11807 : XOR2_X1 port map( A1 => n27573, A2 => n7973, Z => n14675);
   U11813 : NAND2_X2 port map( A1 => n22309, A2 => n3063, ZN => n7973);
   U11829 : INV_X2 port map( I => n13104, ZN => n809);
   U11830 : NAND2_X2 port map( A1 => n5301, A2 => n23846, ZN => n13104);
   U11832 : NOR2_X2 port map( A1 => n1084, A2 => n23036, ZN => n22106);
   U11835 : XOR2_X1 port map( A1 => n23572, A2 => n25098, Z => n19059);
   U11836 : NOR2_X2 port map( A1 => n23276, A2 => n17478, ZN => n27313);
   U11838 : XOR2_X1 port map( A1 => n27314, A2 => n8677, Z => n25606);
   U11839 : XOR2_X1 port map( A1 => n8675, A2 => n26724, Z => n27314);
   U11841 : XOR2_X1 port map( A1 => n13344, A2 => n16924, Z => n17046);
   U11843 : NOR2_X2 port map( A1 => n15381, A2 => n14172, ZN => n13344);
   U11848 : NAND2_X2 port map( A1 => n24566, A2 => n14639, ZN => n17570);
   U11849 : XOR2_X1 port map( A1 => n12681, A2 => n18302, Z => n3840);
   U11851 : XOR2_X1 port map( A1 => n14345, A2 => n25351, Z => n18302);
   U11853 : NOR2_X2 port map( A1 => n9381, A2 => n7379, ZN => n15752);
   U11856 : INV_X2 port map( I => n27316, ZN => n26434);
   U11857 : XOR2_X1 port map( A1 => Plaintext(110), A2 => Key(110), Z => n27316
                           );
   U11859 : NOR2_X1 port map( A1 => n21415, A2 => n21409, ZN => n27318);
   U11863 : XOR2_X1 port map( A1 => n6554, A2 => n26815, Z => n18323);
   U11864 : NOR2_X2 port map( A1 => n28187, A2 => n25278, ZN => n6554);
   U11865 : XOR2_X1 port map( A1 => n1679, A2 => n22121, Z => n643);
   U11866 : XOR2_X1 port map( A1 => n17068, A2 => n13344, Z => n25036);
   U11868 : NOR2_X2 port map( A1 => n12553, A2 => n12554, ZN => n27324);
   U11870 : NAND3_X2 port map( A1 => n6840, A2 => n9967, A3 => n15970, ZN => 
                           n6839);
   U11871 : XOR2_X1 port map( A1 => n27319, A2 => n27382, Z => n22524);
   U11873 : OAI21_X1 port map( A1 => n11645, A2 => n13944, B => n2261, ZN => 
                           n27319);
   U11874 : NAND2_X2 port map( A1 => n20147, A2 => n23817, ZN => n22782);
   U11876 : NOR2_X2 port map( A1 => n12673, A2 => n19959, ZN => n27858);
   U11881 : XOR2_X1 port map( A1 => n19540, A2 => n370, Z => n11990);
   U11882 : NAND3_X2 port map( A1 => n18892, A2 => n13212, A3 => n10170, ZN => 
                           n19540);
   U11883 : NOR2_X2 port map( A1 => n12177, A2 => n20183, ZN => n2472);
   U11887 : XOR2_X1 port map( A1 => n18038, A2 => n15339, Z => n27320);
   U11889 : NAND2_X2 port map( A1 => n15101, A2 => n23665, ZN => n19487);
   U11891 : XOR2_X1 port map( A1 => n27321, A2 => n20621, Z => Ciphertext(8));
   U11893 : NAND2_X1 port map( A1 => n10273, A2 => n23260, ZN => n27321);
   U11894 : OAI21_X2 port map( A1 => n21290, A2 => n21286, B => n3531, ZN => 
                           n21293);
   U11895 : OAI21_X2 port map( A1 => n18472, A2 => n14408, B => n18602, ZN => 
                           n18166);
   U11896 : XOR2_X1 port map( A1 => n27322, A2 => n19418, Z => n9088);
   U11898 : INV_X1 port map( I => n4026, ZN => n27322);
   U11900 : NAND2_X2 port map( A1 => n3279, A2 => n6113, ZN => n19035);
   U11904 : XOR2_X1 port map( A1 => n12739, A2 => n19214, Z => n12242);
   U11908 : NAND2_X2 port map( A1 => n13883, A2 => n13882, ZN => n12739);
   U11909 : AOI22_X2 port map( A1 => n25071, A2 => n16206, B1 => n23270, B2 => 
                           n25072, ZN => n16429);
   U11912 : NAND2_X2 port map( A1 => n23561, A2 => n8921, ZN => n28237);
   U11914 : NOR2_X1 port map( A1 => n28399, A2 => n22598, ZN => n7935);
   U11916 : NAND2_X2 port map( A1 => n14751, A2 => n3336, ZN => n22598);
   U11917 : XOR2_X1 port map( A1 => n16792, A2 => n16791, Z => n22969);
   U11921 : XOR2_X1 port map( A1 => n15708, A2 => n94, Z => n16791);
   U11926 : XOR2_X1 port map( A1 => n5499, A2 => n11684, Z => n16792);
   U11929 : INV_X2 port map( I => n20286, ZN => n20190);
   U11930 : NAND3_X2 port map( A1 => n28272, A2 => n14075, A3 => n20111, ZN => 
                           n20286);
   U11936 : XOR2_X1 port map( A1 => n15447, A2 => n18225, Z => n18276);
   U11937 : NAND3_X2 port map( A1 => n17859, A2 => n17858, A3 => n17860, ZN => 
                           n15447);
   U11941 : NAND2_X2 port map( A1 => n4953, A2 => n11485, ZN => n12896);
   U11947 : AND2_X1 port map( A1 => n1459, A2 => n26620, Z => n19622);
   U11950 : XOR2_X1 port map( A1 => n27999, A2 => n25867, Z => n26536);
   U11952 : NAND2_X1 port map( A1 => n2897, A2 => n2895, ZN => n27323);
   U11956 : NOR2_X2 port map( A1 => n24474, A2 => n3954, ZN => n4362);
   U11957 : NOR2_X2 port map( A1 => n28156, A2 => n28157, ZN => n28155);
   U11965 : NAND2_X2 port map( A1 => n27324, A2 => n12551, ZN => n17855);
   U11966 : BUF_X2 port map( I => n3353, Z => n5796);
   U11967 : NAND2_X2 port map( A1 => n11307, A2 => n23872, ZN => n11318);
   U11972 : NAND2_X2 port map( A1 => n27987, A2 => n27986, ZN => n11307);
   U11977 : INV_X2 port map( I => n5961, ZN => n9344);
   U11978 : OAI22_X2 port map( A1 => n4888, A2 => n27886, B1 => n4253, B2 => 
                           n4252, ZN => n5961);
   U11981 : NAND3_X2 port map( A1 => n27785, A2 => n28184, A3 => n882, ZN => 
                           n27614);
   U11984 : XOR2_X1 port map( A1 => n16922, A2 => n8413, Z => n4674);
   U11988 : AOI22_X2 port map( A1 => n23592, A2 => n1102, B1 => n20068, B2 => 
                           n20270, ZN => n3872);
   U11989 : NOR2_X2 port map( A1 => n24554, A2 => n27377, ZN => n20068);
   U11990 : NOR2_X2 port map( A1 => n27326, A2 => n22104, ZN => n27919);
   U11992 : NOR3_X1 port map( A1 => n1342, A2 => n23311, A3 => n13235, ZN => 
                           n27326);
   U11996 : NOR2_X2 port map( A1 => n15538, A2 => n27327, ZN => n16944);
   U11999 : OAI21_X2 port map( A1 => n16667, A2 => n16668, B => n16670, ZN => 
                           n27327);
   U12000 : XOR2_X1 port map( A1 => n27329, A2 => n26566, Z => Ciphertext(54));
   U12002 : AOI22_X1 port map( A1 => n22729, A2 => n7907, B1 => n7906, B2 => 
                           n20915, ZN => n27329);
   U12007 : NAND2_X2 port map( A1 => n28442, A2 => n25161, ZN => n21846);
   U12008 : INV_X2 port map( I => n7969, ZN => n1104);
   U12009 : NAND3_X2 port map( A1 => n4112, A2 => n11033, A3 => n7667, ZN => 
                           n7969);
   U12010 : BUF_X4 port map( I => n19280, Z => n19890);
   U12016 : OAI21_X2 port map( A1 => n6782, A2 => n20082, B => n27398, ZN => 
                           n26599);
   U12022 : NOR2_X2 port map( A1 => n21759, A2 => n27414, ZN => n20082);
   U12033 : NAND3_X2 port map( A1 => n10823, A2 => n17956, A3 => n10673, ZN => 
                           n27330);
   U12034 : OAI21_X2 port map( A1 => n17952, A2 => n28495, B => n11488, ZN => 
                           n11359);
   U12036 : NOR2_X2 port map( A1 => n25831, A2 => n2198, ZN => n25830);
   U12037 : INV_X2 port map( I => n27331, ZN => n28538);
   U12040 : XOR2_X1 port map( A1 => n4764, A2 => n24805, Z => n27331);
   U12041 : NAND2_X2 port map( A1 => n11872, A2 => n17727, ZN => n17632);
   U12042 : AND2_X2 port map( A1 => n17244, A2 => n13693, Z => n17471);
   U12045 : AOI22_X2 port map( A1 => n946, A2 => n21136, B1 => n13600, B2 => 
                           n20263, ZN => n11013);
   U12047 : XOR2_X1 port map( A1 => n27334, A2 => n27333, Z => n8337);
   U12052 : INV_X2 port map( I => n19427, ZN => n27333);
   U12053 : XOR2_X1 port map( A1 => n7776, A2 => n20694, Z => n27334);
   U12055 : NAND2_X2 port map( A1 => n4783, A2 => n4311, ZN => n27486);
   U12063 : NAND2_X2 port map( A1 => n12267, A2 => n4859, ZN => n4783);
   U12066 : OAI21_X1 port map( A1 => n1577, A2 => n6090, B => n18953, ZN => 
                           n27562);
   U12068 : XOR2_X1 port map( A1 => n20480, A2 => n23648, Z => n20776);
   U12069 : AOI22_X2 port map( A1 => n21875, A2 => n10635, B1 => n9422, B2 => 
                           n21052, ZN => n21051);
   U12070 : XOR2_X1 port map( A1 => n21180, A2 => n27335, Z => n27922);
   U12071 : XOR2_X1 port map( A1 => n6523, A2 => n7848, Z => n27335);
   U12078 : NAND2_X1 port map( A1 => n735, A2 => n27588, ZN => n6211);
   U12079 : XOR2_X1 port map( A1 => n1943, A2 => n25271, Z => n27588);
   U12083 : NAND2_X2 port map( A1 => n27337, A2 => n8498, ZN => n5243);
   U12085 : NAND3_X1 port map( A1 => n27841, A2 => n6658, A3 => n25917, ZN => 
                           n27337);
   U12091 : NOR2_X2 port map( A1 => n27338, A2 => n5346, ZN => n23466);
   U12093 : NOR2_X1 port map( A1 => n17168, A2 => n17169, ZN => n27338);
   U12094 : INV_X4 port map( I => n17653, ZN => n10823);
   U12095 : NAND2_X2 port map( A1 => n17357, A2 => n27682, ZN => n17653);
   U12103 : NOR2_X2 port map( A1 => n24453, A2 => n17210, ZN => n24304);
   U12107 : AND2_X1 port map( A1 => n4611, A2 => n27339, Z => n23776);
   U12108 : NAND2_X2 port map( A1 => n27340, A2 => n7789, ZN => n7569);
   U12109 : BUF_X2 port map( I => n24513, Z => n27341);
   U12112 : NOR2_X2 port map( A1 => n27056, A2 => n17887, ZN => n17801);
   U12114 : NAND2_X2 port map( A1 => n5764, A2 => n5763, ZN => n18081);
   U12118 : XOR2_X1 port map( A1 => n19317, A2 => n13299, Z => n27343);
   U12119 : XOR2_X1 port map( A1 => n16829, A2 => n17152, Z => n7506);
   U12120 : XOR2_X1 port map( A1 => n8274, A2 => n16958, Z => n17152);
   U12123 : NAND2_X2 port map( A1 => n14037, A2 => n12111, ZN => n12139);
   U12124 : OAI22_X2 port map( A1 => n24874, A2 => n2232, B1 => n21344, B2 => 
                           n21347, ZN => n21356);
   U12125 : NAND3_X2 port map( A1 => n14902, A2 => n1703, A3 => n15378, ZN => 
                           n492);
   U12128 : INV_X4 port map( I => n15209, ZN => n21387);
   U12132 : BUF_X4 port map( I => n12946, Z => n28091);
   U12135 : AOI22_X2 port map( A1 => n18899, A2 => n27432, B1 => n18898, B2 => 
                           n817, ZN => n2906);
   U12136 : INV_X4 port map( I => n9583, ZN => n9644);
   U12138 : OAI21_X2 port map( A1 => n16397, A2 => n23749, B => n16572, ZN => 
                           n2852);
   U12154 : INV_X2 port map( I => n6487, ZN => n22634);
   U12155 : OR2_X1 port map( A1 => n23474, A2 => n28141, Z => n9907);
   U12157 : INV_X4 port map( I => n19809, ZN => n28285);
   U12160 : NAND2_X2 port map( A1 => n26302, A2 => n18683, ZN => n26209);
   U12162 : INV_X1 port map( I => n9652, ZN => n27344);
   U12164 : INV_X1 port map( I => n9652, ZN => n28141);
   U12166 : INV_X2 port map( I => n19691, ZN => n19830);
   U12167 : OR2_X2 port map( A1 => n19691, A2 => n14685, Z => n19947);
   U12173 : INV_X1 port map( I => n5573, ZN => n1106);
   U12179 : NAND2_X2 port map( A1 => n9186, A2 => n27634, ZN => n27347);
   U12182 : OR2_X1 port map( A1 => n24534, A2 => n27347, Z => n23210);
   U12183 : NOR2_X1 port map( A1 => n9522, A2 => n9523, ZN => n25792);
   U12184 : NAND2_X1 port map( A1 => n14474, A2 => n25158, ZN => n18324);
   U12185 : OR2_X1 port map( A1 => n15366, A2 => n5919, Z => n18658);
   U12187 : NAND2_X1 port map( A1 => n11579, A2 => n7017, ZN => n22895);
   U12203 : NOR2_X1 port map( A1 => n11579, A2 => n7017, ZN => n27582);
   U12205 : INV_X2 port map( I => n3644, ZN => n27349);
   U12208 : INV_X1 port map( I => n3644, ZN => n4393);
   U12211 : OAI21_X1 port map( A1 => n17573, A2 => n10603, B => n25265, ZN => 
                           n4040);
   U12215 : CLKBUF_X4 port map( I => n14414, Z => n13969);
   U12217 : OAI22_X1 port map( A1 => n2811, A2 => n9141, B1 => n12810, B2 => 
                           n8351, ZN => n28021);
   U12223 : AND2_X1 port map( A1 => n10150, A2 => n14509, Z => n7155);
   U12225 : OAI22_X1 port map( A1 => n14900, A2 => n8996, B1 => n14509, B2 => 
                           n10875, ZN => n10952);
   U12227 : INV_X1 port map( I => n22446, ZN => n8651);
   U12229 : OR2_X2 port map( A1 => n22819, A2 => n22446, Z => n18467);
   U12235 : INV_X2 port map( I => n2869, ZN => n24573);
   U12238 : OAI21_X1 port map( A1 => n17646, A2 => n25724, B => n3119, ZN => 
                           n6656);
   U12239 : CLKBUF_X2 port map( I => n18331, Z => n28269);
   U12241 : OAI22_X1 port map( A1 => n8301, A2 => n18797, B1 => n18522, B2 => 
                           n13349, ZN => n18524);
   U12246 : INV_X1 port map( I => n26640, ZN => n19092);
   U12249 : INV_X1 port map( I => n1129, ZN => n27350);
   U12250 : BUF_X2 port map( I => n3600, Z => n3563);
   U12251 : AOI21_X1 port map( A1 => n3563, A2 => n19689, B => n8794, ZN => 
                           n19690);
   U12252 : NOR2_X1 port map( A1 => n9051, A2 => n26491, ZN => n9107);
   U12275 : NOR2_X1 port map( A1 => n15268, A2 => n15560, ZN => n23035);
   U12279 : NOR2_X1 port map( A1 => n20926, A2 => n20981, ZN => n27824);
   U12282 : NAND3_X1 port map( A1 => n20977, A2 => n20981, A3 => n12465, ZN => 
                           n20984);
   U12294 : AOI21_X1 port map( A1 => n25298, A2 => n944, B => n21992, ZN => 
                           n3658);
   U12304 : INV_X1 port map( I => n17486, ZN => n27351);
   U12310 : BUF_X2 port map( I => n16722, Z => n17560);
   U12315 : INV_X2 port map( I => n15030, ZN => n13532);
   U12324 : CLKBUF_X2 port map( I => n15030, Z => n10958);
   U12325 : NOR2_X1 port map( A1 => n13815, A2 => n5244, ZN => n15481);
   U12326 : AOI22_X1 port map( A1 => n16680, A2 => n13815, B1 => n24727, B2 => 
                           n16681, ZN => n9871);
   U12332 : NAND2_X1 port map( A1 => n5244, A2 => n13815, ZN => n15992);
   U12343 : NAND2_X1 port map( A1 => n27404, A2 => n15469, ZN => n12399);
   U12346 : AOI21_X2 port map( A1 => n8083, A2 => n8082, B => n25259, ZN => 
                           n27352);
   U12349 : AOI21_X1 port map( A1 => n8083, A2 => n8082, B => n25259, ZN => 
                           n19535);
   U12361 : NOR2_X1 port map( A1 => n7668, A2 => n16497, ZN => n27353);
   U12362 : INV_X1 port map( I => n17493, ZN => n27354);
   U12366 : INV_X1 port map( I => n27354, ZN => n27355);
   U12367 : NOR2_X1 port map( A1 => n7668, A2 => n16497, ZN => n13528);
   U12372 : INV_X2 port map( I => n13415, ZN => n7668);
   U12378 : NAND2_X1 port map( A1 => n15270, A2 => n27627, ZN => n27404);
   U12379 : OAI21_X1 port map( A1 => n21987, A2 => n9094, B => n24336, ZN => 
                           n3465);
   U12382 : NOR2_X2 port map( A1 => n14584, A2 => n16123, ZN => n15766);
   U12385 : INV_X2 port map( I => n26317, ZN => n784);
   U12388 : NOR2_X1 port map( A1 => n26317, A2 => n13372, ZN => n22459);
   U12409 : NAND2_X1 port map( A1 => n26317, A2 => n18719, ZN => n11240);
   U12412 : NOR2_X1 port map( A1 => n20431, A2 => n20430, ZN => n4925);
   U12421 : NOR3_X1 port map( A1 => n17729, A2 => n17727, A3 => n17728, ZN => 
                           n28187);
   U12426 : OR2_X2 port map( A1 => n14750, A2 => n7319, Z => n14749);
   U12427 : OR2_X1 port map( A1 => n15227, A2 => n7087, Z => n13455);
   U12428 : CLKBUF_X1 port map( I => n7403, Z => n27388);
   U12430 : NOR2_X1 port map( A1 => n20022, A2 => n4274, ZN => n7063);
   U12431 : INV_X1 port map( I => n3878, ZN => n24707);
   U12433 : INV_X1 port map( I => n25324, ZN => n28165);
   U12436 : NOR2_X1 port map( A1 => n6392, A2 => n19845, ZN => n23626);
   U12437 : OAI21_X1 port map( A1 => n4401, A2 => n3824, B => n2254, ZN => 
                           n28536);
   U12438 : NAND2_X1 port map( A1 => n574, A2 => n27123, ZN => n13457);
   U12446 : OAI21_X1 port map( A1 => n16076, A2 => n574, B => n24132, ZN => 
                           n15761);
   U12451 : AND2_X2 port map( A1 => n574, A2 => n15905, Z => n16219);
   U12452 : OAI21_X1 port map( A1 => n3763, A2 => n877, B => n18455, ZN => 
                           n3762);
   U12461 : AOI22_X1 port map( A1 => n17248, A2 => n10150, B1 => n1223, B2 => 
                           n14900, ZN => n10165);
   U12462 : AND2_X1 port map( A1 => n735, A2 => n4263, Z => n23075);
   U12464 : INV_X2 port map( I => n9131, ZN => n27356);
   U12468 : AND2_X1 port map( A1 => n21328, A2 => n27356, Z => n5483);
   U12469 : NOR2_X1 port map( A1 => n10188, A2 => n10189, ZN => n9822);
   U12470 : CLKBUF_X12 port map( I => n666, Z => n174);
   U12472 : NAND2_X2 port map( A1 => n18836, A2 => n28216, ZN => n27357);
   U12474 : INV_X1 port map( I => n23105, ZN => n2756);
   U12478 : NAND2_X1 port map( A1 => n734, A2 => n9087, ZN => n25420);
   U12487 : NOR2_X1 port map( A1 => n18487, A2 => n24870, ZN => n24050);
   U12492 : CLKBUF_X2 port map( I => n15448, Z => n27497);
   U12493 : INV_X1 port map( I => n21066, ZN => n3344);
   U12497 : AOI21_X1 port map( A1 => n23309, A2 => n1260, B => n16164, ZN => 
                           n11712);
   U12498 : AOI21_X1 port map( A1 => n3573, A2 => n3571, B => n16164, ZN => 
                           n3570);
   U12500 : NAND2_X1 port map( A1 => n11997, A2 => n11996, ZN => n11501);
   U12501 : OR2_X2 port map( A1 => n17391, A2 => n791, Z => n8625);
   U12504 : AOI21_X2 port map( A1 => n4371, A2 => n13732, B => n21834, ZN => 
                           n27360);
   U12506 : NOR2_X1 port map( A1 => n25530, A2 => n17757, ZN => n24785);
   U12507 : NAND2_X1 port map( A1 => n11157, A2 => n17757, ZN => n2326);
   U12508 : INV_X2 port map( I => n23978, ZN => n11411);
   U12513 : INV_X1 port map( I => n12533, ZN => n28531);
   U12517 : NAND2_X1 port map( A1 => n15279, A2 => n14975, ZN => n14217);
   U12518 : AOI21_X2 port map( A1 => n20861, A2 => n20899, B => n13879, ZN => 
                           n13574);
   U12521 : NAND2_X1 port map( A1 => n10978, A2 => n7682, ZN => n14169);
   U12522 : NAND3_X2 port map( A1 => n2034, A2 => n19761, A3 => n2492, ZN => 
                           n26005);
   U12525 : NAND3_X1 port map( A1 => n18982, A2 => n19079, A3 => n11983, ZN => 
                           n18838);
   U12528 : NAND3_X1 port map( A1 => n17722, A2 => n6794, A3 => n11112, ZN => 
                           n9495);
   U12529 : OAI21_X1 port map( A1 => n1617, A2 => n17722, B => n6629, ZN => 
                           n6591);
   U12530 : XOR2_X1 port map( A1 => n27474, A2 => n10711, Z => n27361);
   U12533 : OR3_X1 port map( A1 => n2309, A2 => n8552, A3 => n8553, Z => n27362
                           );
   U12535 : NOR2_X1 port map( A1 => n8557, A2 => n18977, ZN => n8552);
   U12545 : INV_X2 port map( I => n631, ZN => n5639);
   U12547 : AOI21_X1 port map( A1 => n14153, A2 => n5163, B => n5047, ZN => 
                           n9949);
   U12551 : NAND2_X1 port map( A1 => n12524, A2 => n5047, ZN => n11212);
   U12553 : XNOR2_X1 port map( A1 => n21247, A2 => n21302, ZN => n28323);
   U12554 : INV_X2 port map( I => n14513, ZN => n23674);
   U12555 : CLKBUF_X4 port map( I => n13628, Z => n4122);
   U12556 : INV_X2 port map( I => n24094, ZN => n6764);
   U12557 : NAND3_X1 port map( A1 => n4852, A2 => n4850, A3 => n4849, ZN => 
                           n4848);
   U12560 : INV_X1 port map( I => n21457, ZN => n11248);
   U12562 : CLKBUF_X4 port map( I => n19472, Z => n19952);
   U12564 : INV_X2 port map( I => n16728, ZN => n794);
   U12569 : NAND2_X1 port map( A1 => n237, A2 => n17941, ZN => n10131);
   U12572 : NAND2_X1 port map( A1 => n25009, A2 => n20938, ZN => n8029);
   U12576 : INV_X1 port map( I => n5009, ZN => n27363);
   U12582 : CLKBUF_X1 port map( I => n3751, Z => n27745);
   U12585 : AOI21_X1 port map( A1 => n21451, A2 => n21452, B => n12466, ZN => 
                           n13929);
   U12589 : OAI21_X1 port map( A1 => n10851, A2 => n6080, B => n13780, ZN => 
                           n12466);
   U12591 : NAND3_X1 port map( A1 => n20975, A2 => n24470, A3 => n25841, ZN => 
                           n15335);
   U12595 : NAND2_X1 port map( A1 => n20975, A2 => n21020, ZN => n13847);
   U12597 : INV_X1 port map( I => n12598, ZN => n20975);
   U12603 : INV_X1 port map( I => n21168, ZN => n13822);
   U12607 : AOI22_X1 port map( A1 => n3990, A2 => n859, B1 => n4791, B2 => 
                           n4783, ZN => n27364);
   U12608 : AOI22_X1 port map( A1 => n3990, A2 => n859, B1 => n4791, B2 => 
                           n4783, ZN => n10339);
   U12609 : OR2_X1 port map( A1 => n18487, A2 => n23004, Z => n2945);
   U12610 : NAND3_X1 port map( A1 => n27345, A2 => n22025, A3 => n15544, ZN => 
                           n28500);
   U12622 : XOR2_X1 port map( A1 => n27357, A2 => n19412, Z => n27365);
   U12624 : OAI22_X2 port map( A1 => n23143, A2 => n20310, B1 => n9447, B2 => 
                           n23913, ZN => n27366);
   U12638 : OAI22_X1 port map( A1 => n23143, A2 => n20310, B1 => n9447, B2 => 
                           n23913, ZN => n9445);
   U12641 : CLKBUF_X12 port map( I => Key(122), Z => n20519);
   U12643 : OAI21_X1 port map( A1 => n27630, A2 => n12973, B => n25557, ZN => 
                           n13075);
   U12644 : CLKBUF_X4 port map( I => n8262, Z => n21779);
   U12647 : NOR2_X1 port map( A1 => n27988, A2 => n20932, ZN => n27987);
   U12651 : NAND2_X1 port map( A1 => n10484, A2 => n20932, ZN => n10483);
   U12653 : AOI22_X1 port map( A1 => n16680, A2 => n4281, B1 => n4462, B2 => 
                           n5244, ZN => n28275);
   U12654 : NAND2_X2 port map( A1 => n2556, A2 => n2555, ZN => n15778);
   U12664 : NAND2_X1 port map( A1 => n2051, A2 => n5305, ZN => n17795);
   U12666 : NAND2_X1 port map( A1 => n2391, A2 => n14451, ZN => n16394);
   U12668 : CLKBUF_X4 port map( I => n19019, Z => n23138);
   U12671 : OR2_X2 port map( A1 => n2404, A2 => n338, Z => n2406);
   U12672 : CLKBUF_X2 port map( I => n10241, Z => n3584);
   U12674 : NAND2_X1 port map( A1 => n9315, A2 => n9314, ZN => n10395);
   U12679 : OAI22_X1 port map( A1 => n7983, A2 => n7985, B1 => n8070, B2 => 
                           n7986, ZN => n7982);
   U12681 : AOI21_X1 port map( A1 => n22950, A2 => n12018, B => n9929, ZN => 
                           n9928);
   U12683 : INV_X1 port map( I => n13303, ZN => n821);
   U12684 : NAND2_X1 port map( A1 => n13330, A2 => n19991, ZN => n21261);
   U12687 : NAND2_X1 port map( A1 => n26140, A2 => n855, ZN => n12475);
   U12688 : OR2_X1 port map( A1 => n4679, A2 => n22429, Z => n4706);
   U12689 : NAND3_X1 port map( A1 => n8935, A2 => n927, A3 => n4315, ZN => 
                           n20599);
   U12691 : AOI22_X1 port map( A1 => n6353, A2 => n6433, B1 => n14749, B2 => 
                           n6432, ZN => n15090);
   U12694 : NAND2_X2 port map( A1 => n25823, A2 => n18882, ZN => n27369);
   U12695 : AND2_X2 port map( A1 => n27940, A2 => n22157, Z => n27370);
   U12696 : NAND2_X2 port map( A1 => n20282, A2 => n20281, ZN => n27371);
   U12702 : NAND2_X1 port map( A1 => n20282, A2 => n20281, ZN => n20553);
   U12705 : NOR2_X1 port map( A1 => n11089, A2 => n21208, ZN => n10621);
   U12706 : AND2_X1 port map( A1 => n20703, A2 => n22730, Z => n20697);
   U12710 : OAI22_X1 port map( A1 => n27859, A2 => n21008, B1 => n21004, B2 => 
                           n13395, ZN => n15678);
   U12711 : AND2_X2 port map( A1 => n16098, A2 => n16097, Z => n27372);
   U12714 : NAND3_X1 port map( A1 => n28536, A2 => n20648, A3 => n20649, ZN => 
                           n56);
   U12721 : NOR3_X1 port map( A1 => n540, A2 => n2527, A3 => n2831, ZN => 
                           n11295);
   U12727 : OAI22_X1 port map( A1 => n17187, A2 => n2831, B1 => n17311, B2 => 
                           n2527, ZN => n24791);
   U12730 : AOI21_X1 port map( A1 => n17311, A2 => n3360, B => n2831, ZN => 
                           n23507);
   U12735 : NOR2_X1 port map( A1 => n21324, A2 => n9131, ZN => n7131);
   U12736 : CLKBUF_X12 port map( I => n12653, Z => n5009);
   U12741 : NAND2_X2 port map( A1 => n1606, A2 => n1607, ZN => n27563);
   U12748 : NAND2_X1 port map( A1 => n5609, A2 => n5213, ZN => n27373);
   U12749 : NAND2_X1 port map( A1 => n5609, A2 => n5213, ZN => n6809);
   U12757 : INV_X2 port map( I => n6089, ZN => n7565);
   U12758 : NAND2_X1 port map( A1 => n23253, A2 => n12644, ZN => n27602);
   U12759 : AND2_X2 port map( A1 => n20736, A2 => n20783, Z => n21936);
   U12761 : OR2_X1 port map( A1 => n6999, A2 => n9050, Z => n27810);
   U12763 : NAND2_X1 port map( A1 => n19676, A2 => n6861, ZN => n8208);
   U12764 : INV_X2 port map( I => n10062, ZN => n18580);
   U12769 : NOR3_X1 port map( A1 => n18581, A2 => n18580, A3 => n10537, ZN => 
                           n18582);
   U12774 : AOI21_X1 port map( A1 => n26030, A2 => n3160, B => n18432, ZN => 
                           n8026);
   U12778 : NAND2_X2 port map( A1 => n6502, A2 => n24596, ZN => n27374);
   U12790 : NOR2_X1 port map( A1 => n9450, A2 => n12477, ZN => n9449);
   U12794 : NOR2_X1 port map( A1 => n28432, A2 => n21668, ZN => n28431);
   U12795 : NAND2_X1 port map( A1 => n28365, A2 => n28366, ZN => n7837);
   U12797 : NOR2_X1 port map( A1 => n6046, A2 => n21692, ZN => n8217);
   U12803 : CLKBUF_X2 port map( I => n12531, Z => n23463);
   U12805 : AOI22_X1 port map( A1 => n12187, A2 => n26712, B1 => n21001, B2 => 
                           n12559, ZN => n27995);
   U12806 : INV_X1 port map( I => n13095, ZN => n27375);
   U12808 : INV_X2 port map( I => n13095, ZN => n935);
   U12809 : BUF_X2 port map( I => n24533, Z => n253);
   U12810 : INV_X1 port map( I => n18182, ZN => n4517);
   U12815 : NOR2_X1 port map( A1 => n14096, A2 => n7791, ZN => n5245);
   U12820 : NAND3_X1 port map( A1 => n5582, A2 => n14096, A3 => n7791, ZN => 
                           n14095);
   U12822 : NAND2_X1 port map( A1 => n19944, A2 => n19943, ZN => n27377);
   U12826 : AOI22_X1 port map( A1 => n12675, A2 => n22762, B1 => n6181, B2 => 
                           n21659, ZN => n21660);
   U12833 : NAND2_X1 port map( A1 => n10058, A2 => n6642, ZN => n17993);
   U12836 : OR2_X1 port map( A1 => n8514, A2 => n23161, Z => n18856);
   U12838 : INV_X1 port map( I => n12653, ZN => n10732);
   U12839 : INV_X2 port map( I => n13386, ZN => n19827);
   U12843 : NOR2_X1 port map( A1 => n19951, A2 => n19827, ZN => n19717);
   U12849 : NAND3_X2 port map( A1 => n14889, A2 => n28317, A3 => n28316, ZN => 
                           n27378);
   U12850 : CLKBUF_X12 port map( I => n13491, Z => n27379);
   U12851 : INV_X1 port map( I => n27518, ZN => n13769);
   U12853 : CLKBUF_X1 port map( I => n16496, Z => n28172);
   U12855 : NAND2_X1 port map( A1 => n16496, A2 => n5442, ZN => n16540);
   U12860 : INV_X1 port map( I => n16496, ZN => n16615);
   U12864 : NAND2_X1 port map( A1 => n7759, A2 => n22529, ZN => n10425);
   U12866 : AND2_X2 port map( A1 => n6841, A2 => n6839, Z => n27381);
   U12867 : OAI21_X1 port map( A1 => n708, A2 => n1082, B => n4667, ZN => n4846
                           );
   U12868 : INV_X2 port map( I => n4667, ZN => n4742);
   U12870 : CLKBUF_X12 port map( I => n4355, Z => n27382);
   U12873 : AOI21_X1 port map( A1 => n5292, A2 => n253, B => n4393, ZN => 
                           n22437);
   U12875 : NAND3_X1 port map( A1 => n978, A2 => n26155, A3 => n2925, ZN => 
                           n11517);
   U12880 : INV_X2 port map( I => n15703, ZN => n20141);
   U12881 : NAND3_X1 port map( A1 => n21222, A2 => n21221, A3 => n22027, ZN => 
                           n6830);
   U12886 : INV_X1 port map( I => n20534, ZN => n4478);
   U12892 : CLKBUF_X12 port map( I => n13793, Z => n28148);
   U12893 : AOI21_X1 port map( A1 => n8049, A2 => n1163, B => n19190, ZN => 
                           n8416);
   U12896 : OR2_X2 port map( A1 => n11024, A2 => n15025, Z => n11023);
   U12897 : INV_X1 port map( I => n13879, ZN => n2184);
   U12899 : NAND3_X1 port map( A1 => n26601, A2 => n26667, A3 => n19846, ZN => 
                           n13522);
   U12902 : INV_X1 port map( I => n936, ZN => n27427);
   U12904 : OAI21_X1 port map( A1 => n1260, A2 => n28032, B => n6427, ZN => 
                           n6658);
   U12914 : CLKBUF_X4 port map( I => n2588, Z => n2587);
   U12922 : AND3_X1 port map( A1 => n936, A2 => n21174, A3 => n21166, Z => 
                           n15656);
   U12923 : OR2_X1 port map( A1 => n21174, A2 => n11107, Z => n4541);
   U12924 : NAND2_X1 port map( A1 => n14806, A2 => n20897, ZN => n7881);
   U12925 : NAND2_X2 port map( A1 => n25789, A2 => n5236, ZN => n27384);
   U12929 : NAND2_X1 port map( A1 => n25789, A2 => n5236, ZN => n18239);
   U12930 : AND2_X1 port map( A1 => n21623, A2 => n21622, Z => n24548);
   U12931 : INV_X1 port map( I => n868, ZN => n28208);
   U12934 : OAI21_X1 port map( A1 => n13986, A2 => n12508, B => n13934, ZN => 
                           n27866);
   U12935 : CLKBUF_X4 port map( I => n5475, Z => n21788);
   U12936 : NAND2_X1 port map( A1 => n18660, A2 => n14420, ZN => n13191);
   U12937 : INV_X1 port map( I => n9087, ZN => n27385);
   U12938 : NAND2_X2 port map( A1 => n22205, A2 => n22204, ZN => n28274);
   U12939 : OAI21_X1 port map( A1 => n7836, A2 => n6037, B => n1070, ZN => 
                           n28366);
   U12942 : AOI21_X1 port map( A1 => n21395, A2 => n21445, B => n14281, ZN => 
                           n15606);
   U12946 : INV_X2 port map( I => n8262, ZN => n12964);
   U12948 : CLKBUF_X4 port map( I => n5797, Z => n5753);
   U12951 : INV_X1 port map( I => n8890, ZN => n27691);
   U12954 : INV_X1 port map( I => n16215, ZN => n21959);
   U12960 : INV_X1 port map( I => n16980, ZN => n27513);
   U12962 : INV_X1 port map( I => n20100, ZN => n20090);
   U12964 : NAND2_X1 port map( A1 => n24562, A2 => n22753, ZN => n8162);
   U12965 : NAND2_X1 port map( A1 => n2670, A2 => n10764, ZN => n19983);
   U12969 : NAND2_X1 port map( A1 => n1977, A2 => n1980, ZN => n27387);
   U12978 : NOR2_X1 port map( A1 => n21620, A2 => n21586, ZN => n24261);
   U12980 : NAND2_X2 port map( A1 => n22691, A2 => n28007, ZN => n27389);
   U12981 : NOR2_X1 port map( A1 => n8425, A2 => n18474, ZN => n28423);
   U12982 : OAI21_X1 port map( A1 => n18460, A2 => n18458, B => n8425, ZN => 
                           n14407);
   U12983 : NAND2_X1 port map( A1 => n21136, A2 => n20263, ZN => n21137);
   U12990 : NOR2_X2 port map( A1 => n21094, A2 => n15451, ZN => n15450);
   U12992 : OAI21_X1 port map( A1 => n1117, A2 => n19866, B => n19865, ZN => 
                           n27719);
   U12994 : NAND2_X1 port map( A1 => n21627, A2 => n13426, ZN => n13097);
   U12995 : INV_X2 port map( I => n9993, ZN => n15560);
   U13003 : NAND2_X2 port map( A1 => n13994, A2 => n24738, ZN => n27390);
   U13006 : NAND2_X2 port map( A1 => n13993, A2 => n13992, ZN => n24738);
   U13012 : CLKBUF_X4 port map( I => n21016, Z => n14341);
   U13019 : NAND2_X2 port map( A1 => n21929, A2 => n27688, ZN => n27391);
   U13025 : NAND2_X1 port map( A1 => n21929, A2 => n27688, ZN => n9049);
   U13026 : INV_X2 port map( I => n28113, ZN => n23935);
   U13033 : OAI21_X1 port map( A1 => n10469, A2 => n10470, B => n9561, ZN => 
                           n26060);
   U13035 : INV_X1 port map( I => n5206, ZN => n8167);
   U13037 : OAI21_X2 port map( A1 => n5839, A2 => n19785, B => n14522, ZN => 
                           n15373);
   U13043 : OR2_X2 port map( A1 => n6047, A2 => n21916, Z => n6885);
   U13044 : BUF_X2 port map( I => n20559, Z => n21059);
   U13049 : NAND2_X1 port map( A1 => n21016, A2 => n20559, ZN => n25173);
   U13053 : NAND2_X1 port map( A1 => n3481, A2 => n12057, ZN => n27392);
   U13056 : BUF_X2 port map( I => n11224, Z => n23719);
   U13057 : INV_X2 port map( I => n11224, ZN => n25415);
   U13066 : INV_X1 port map( I => n18144, ZN => n27702);
   U13067 : NOR2_X1 port map( A1 => n11213, A2 => n19930, ZN => n10139);
   U13072 : NAND3_X1 port map( A1 => n11213, A2 => n10041, A3 => n754, ZN => 
                           n19571);
   U13077 : INV_X1 port map( I => n14033, ZN => n27603);
   U13088 : NAND2_X1 port map( A1 => n20751, A2 => n14352, ZN => n20752);
   U13090 : NAND2_X1 port map( A1 => n8910, A2 => n25879, ZN => n10794);
   U13091 : INV_X1 port map( I => n25879, ZN => n26028);
   U13094 : NAND2_X1 port map( A1 => n20866, A2 => n5367, ZN => n20457);
   U13101 : NOR2_X1 port map( A1 => n10904, A2 => n13619, ZN => n1997);
   U13105 : AOI22_X1 port map( A1 => n7199, A2 => n13741, B1 => n21413, B2 => 
                           n25369, ZN => n21416);
   U13106 : INV_X1 port map( I => n13741, ZN => n13756);
   U13107 : INV_X2 port map( I => n10639, ZN => n10484);
   U13112 : AOI21_X1 port map( A1 => n20933, A2 => n10639, B => n28059, ZN => 
                           n20936);
   U13114 : NAND2_X1 port map( A1 => n10639, A2 => n20938, ZN => n27986);
   U13116 : CLKBUF_X4 port map( I => n722, Z => n1383);
   U13123 : NAND2_X1 port map( A1 => n21168, A2 => n21174, ZN => n25784);
   U13124 : NAND2_X1 port map( A1 => n12287, A2 => n21175, ZN => n1457);
   U13127 : INV_X2 port map( I => n14917, ZN => n1033);
   U13129 : AOI21_X2 port map( A1 => n14390, A2 => n22516, B => n21720, ZN => 
                           n27395);
   U13136 : NAND2_X1 port map( A1 => n1121, A2 => n4364, ZN => n6585);
   U13138 : NOR2_X1 port map( A1 => n4364, A2 => n3953, ZN => n27517);
   U13140 : INV_X2 port map( I => n598, ZN => n4364);
   U13141 : NAND2_X1 port map( A1 => n5159, A2 => n5161, ZN => n27393);
   U13144 : NAND2_X1 port map( A1 => n5159, A2 => n5161, ZN => n27394);
   U13145 : NAND2_X1 port map( A1 => n5159, A2 => n5161, ZN => n14145);
   U13146 : OAI21_X2 port map( A1 => n25430, A2 => n25429, B => n14579, ZN => 
                           n5161);
   U13150 : NAND2_X2 port map( A1 => n21696, A2 => n15307, ZN => n14390);
   U13153 : AOI21_X1 port map( A1 => n1163, A2 => n19191, B => n18949, ZN => 
                           n6534);
   U13154 : AND3_X2 port map( A1 => n6928, A2 => n6927, A3 => n6931, Z => 
                           n27397);
   U13156 : NAND2_X1 port map( A1 => n8723, A2 => n19975, ZN => n2730);
   U13160 : NAND2_X1 port map( A1 => n27630, A2 => n19975, ZN => n25557);
   U13162 : CLKBUF_X1 port map( I => n19975, Z => n22943);
   U13165 : XOR2_X1 port map( A1 => n21298, A2 => n1611, Z => n27399);
   U13166 : NAND2_X1 port map( A1 => n28262, A2 => n28211, ZN => n28261);
   U13170 : INV_X4 port map( I => n13824, ZN => n26382);
   U13175 : OAI21_X1 port map( A1 => n3759, A2 => n20703, B => n28376, ZN => 
                           n22221);
   U13178 : INV_X1 port map( I => n2292, ZN => n954);
   U13180 : XOR2_X1 port map( A1 => n24377, A2 => n1671, Z => n27402);
   U13182 : XOR2_X1 port map( A1 => n25747, A2 => n6291, Z => n27403);
   U13187 : INV_X1 port map( I => n7918, ZN => n7960);
   U13191 : CLKBUF_X2 port map( I => n7918, Z => n5407);
   U13192 : NAND2_X1 port map( A1 => n5488, A2 => n17460, ZN => n17461);
   U13197 : CLKBUF_X12 port map( I => n7651, Z => n5488);
   U13202 : INV_X1 port map( I => n935, ZN => n27405);
   U13203 : XNOR2_X1 port map( A1 => n5648, A2 => n5646, ZN => n27406);
   U13204 : AND3_X2 port map( A1 => n7105, A2 => n7537, A3 => n10394, Z => 
                           n27407);
   U13210 : NAND2_X2 port map( A1 => n10405, A2 => n3983, ZN => n7105);
   U13212 : INV_X1 port map( I => n27406, ZN => n28305);
   U13213 : NOR2_X1 port map( A1 => n21100, A2 => n13461, ZN => n20968);
   U13216 : OAI21_X1 port map( A1 => n13461, A2 => n26512, B => n10558, ZN => 
                           n21994);
   U13220 : NAND2_X1 port map( A1 => n18398, A2 => n12980, ZN => n23147);
   U13232 : NOR2_X1 port map( A1 => n11323, A2 => n27822, ZN => n12044);
   U13236 : INV_X2 port map( I => n21501, ZN => n1074);
   U13241 : OAI21_X1 port map( A1 => n2307, A2 => n14583, B => n3725, ZN => 
                           n3737);
   U13247 : AOI22_X1 port map( A1 => n22216, A2 => n20128, B1 => n11372, B2 => 
                           n26944, ZN => n27408);
   U13249 : AND2_X1 port map( A1 => n21394, A2 => n21406, Z => n5360);
   U13254 : NAND3_X1 port map( A1 => n21685, A2 => n25314, A3 => n9047, ZN => 
                           n21674);
   U13259 : INV_X1 port map( I => n6237, ZN => n26017);
   U13260 : OAI21_X1 port map( A1 => n25697, A2 => n17723, B => n25926, ZN => 
                           n5630);
   U13274 : INV_X1 port map( I => n12532, ZN => n14123);
   U13275 : XNOR2_X1 port map( A1 => Plaintext(152), A2 => Key(152), ZN => 
                           n16065);
   U13278 : XOR2_X1 port map( A1 => n23047, A2 => n11322, Z => n27409);
   U13281 : XNOR2_X1 port map( A1 => n10986, A2 => n20399, ZN => n1353);
   U13287 : AOI21_X1 port map( A1 => n19633, A2 => n8255, B => n26382, ZN => 
                           n2635);
   U13295 : NAND3_X1 port map( A1 => n8192, A2 => n28121, A3 => n26382, ZN => 
                           n7458);
   U13299 : OR2_X1 port map( A1 => n16065, A2 => n16066, Z => n16100);
   U13300 : NAND2_X1 port map( A1 => n4712, A2 => n12206, ZN => n4150);
   U13302 : NAND2_X1 port map( A1 => n18763, A2 => n14022, ZN => n22557);
   U13305 : INV_X2 port map( I => n10210, ZN => n1073);
   U13312 : NAND2_X1 port map( A1 => n9807, A2 => n9805, ZN => n27411);
   U13313 : NAND2_X1 port map( A1 => n9807, A2 => n9805, ZN => n27412);
   U13314 : NAND2_X1 port map( A1 => n9807, A2 => n9805, ZN => n12675);
   U13316 : NOR2_X1 port map( A1 => n21737, A2 => n27471, ZN => n28347);
   U13321 : NOR2_X1 port map( A1 => n21734, A2 => n21737, ZN => n21736);
   U13327 : CLKBUF_X4 port map( I => n20336, Z => n7457);
   U13329 : AOI21_X1 port map( A1 => n21059, A2 => n21096, B => n21062, ZN => 
                           n14508);
   U13330 : NOR2_X1 port map( A1 => n12503, A2 => n20200, ZN => n14514);
   U13332 : OAI21_X1 port map( A1 => n23128, A2 => n16711, B => n22529, ZN => 
                           n10155);
   U13346 : CLKBUF_X4 port map( I => n16711, Z => n11503);
   U13350 : CLKBUF_X12 port map( I => n21714, Z => n27413);
   U13351 : INV_X1 port map( I => n9056, ZN => n27618);
   U13352 : CLKBUF_X4 port map( I => n10474, Z => n24442);
   U13354 : OAI21_X1 port map( A1 => n1121, A2 => n19781, B => n3954, ZN => 
                           n19568);
   U13359 : AND2_X1 port map( A1 => n19114, A2 => n28547, Z => n8027);
   U13374 : NOR2_X1 port map( A1 => n25770, A2 => n28547, ZN => n76);
   U13376 : INV_X2 port map( I => n2041, ZN => n9865);
   U13380 : NAND2_X1 port map( A1 => n9865, A2 => n17036, ZN => n4111);
   U13384 : INV_X2 port map( I => n9865, ZN => n13674);
   U13385 : OAI21_X1 port map( A1 => n17036, A2 => n9865, B => n17204, ZN => 
                           n6367);
   U13388 : OAI21_X1 port map( A1 => n619, A2 => n9865, B => n15699, ZN => 
                           n4267);
   U13391 : NAND2_X1 port map( A1 => n2079, A2 => n28339, ZN => n27414);
   U13392 : INV_X1 port map( I => n17202, ZN => n17514);
   U13396 : NOR2_X1 port map( A1 => n19090, A2 => n6906, ZN => n27870);
   U13397 : INV_X2 port map( I => n6473, ZN => n25952);
   U13398 : OAI22_X2 port map( A1 => n22629, A2 => n23835, B1 => n18923, B2 => 
                           n19009, ZN => n27415);
   U13399 : OAI22_X1 port map( A1 => n22629, A2 => n23835, B1 => n18923, B2 => 
                           n19009, ZN => n19373);
   U13400 : AND2_X2 port map( A1 => n9236, A2 => n18953, Z => n22629);
   U13402 : CLKBUF_X12 port map( I => n26494, Z => n25499);
   U13405 : INV_X1 port map( I => n797, ZN => n1261);
   U13409 : NAND2_X1 port map( A1 => n12066, A2 => n12309, ZN => n20923);
   U13410 : INV_X2 port map( I => n21455, ZN => n15345);
   U13418 : INV_X2 port map( I => n16493, ZN => n23236);
   U13429 : NOR2_X1 port map( A1 => n910, A2 => n16493, ZN => n16438);
   U13434 : INV_X2 port map( I => n14641, ZN => n26027);
   U13435 : INV_X1 port map( I => n7832, ZN => n481);
   U13436 : INV_X1 port map( I => n14401, ZN => n25766);
   U13439 : OR2_X2 port map( A1 => n14401, A2 => n6859, Z => n14967);
   U13442 : OR2_X1 port map( A1 => n27409, A2 => n7181, Z => n19643);
   U13450 : NAND2_X1 port map( A1 => n4212, A2 => n6999, ZN => n3165);
   U13455 : INV_X2 port map( I => n1699, ZN => n14334);
   U13468 : INV_X1 port map( I => n5008, ZN => n12219);
   U13477 : OR2_X1 port map( A1 => n329, A2 => n5008, Z => n12892);
   U13483 : NAND2_X2 port map( A1 => n12656, A2 => n25827, ZN => n27418);
   U13490 : NAND2_X2 port map( A1 => n13541, A2 => n25779, ZN => n25827);
   U13494 : AND2_X2 port map( A1 => n4370, A2 => n20245, Z => n21834);
   U13495 : OAI21_X1 port map( A1 => n20245, A2 => n15076, B => n20248, ZN => 
                           n4371);
   U13500 : NAND2_X1 port map( A1 => n23283, A2 => n23891, ZN => n18238);
   U13506 : INV_X2 port map( I => n7904, ZN => n20976);
   U13508 : NAND2_X1 port map( A1 => n20100, A2 => n13925, ZN => n15151);
   U13518 : OAI22_X1 port map( A1 => n20484, A2 => n21722, B1 => n15307, B2 => 
                           n28027, ZN => n10284);
   U13521 : NAND2_X1 port map( A1 => n20657, A2 => n4766, ZN => n8560);
   U13523 : INV_X2 port map( I => n27419, ZN => n21590);
   U13525 : XNOR2_X1 port map( A1 => n21377, A2 => n21378, ZN => n27420);
   U13526 : NAND3_X2 port map( A1 => n5751, A2 => n12817, A3 => n11646, ZN => 
                           n27421);
   U13529 : NAND3_X1 port map( A1 => n5751, A2 => n12817, A3 => n11646, ZN => 
                           n19180);
   U13530 : INV_X1 port map( I => n9902, ZN => n9903);
   U13531 : NAND2_X1 port map( A1 => n11992, A2 => n10081, ZN => n28270);
   U13540 : NAND2_X1 port map( A1 => n10081, A2 => n10985, ZN => n12706);
   U13545 : OAI21_X1 port map( A1 => n10081, A2 => n11992, B => n13380, ZN => 
                           n10082);
   U13546 : NOR3_X1 port map( A1 => n10081, A2 => n27648, A3 => n11992, ZN => 
                           n11366);
   U13558 : INV_X1 port map( I => n19188, ZN => n27503);
   U13559 : OAI21_X1 port map( A1 => n14062, A2 => n6681, B => n17230, ZN => 
                           n23287);
   U13560 : NAND2_X1 port map( A1 => n14062, A2 => n6681, ZN => n23339);
   U13565 : NOR2_X1 port map( A1 => n24299, A2 => n6681, ZN => n3921);
   U13583 : OAI21_X1 port map( A1 => n6681, A2 => n17558, B => n740, ZN => 
                           n3648);
   U13592 : AOI22_X1 port map( A1 => n27419, A2 => n21507, B1 => n14679, B2 => 
                           n951, ZN => n12649);
   U13602 : AOI21_X1 port map( A1 => n951, A2 => n21590, B => n21507, ZN => 
                           n21508);
   U13609 : INV_X2 port map( I => n1017, ZN => n3674);
   U13610 : INV_X2 port map( I => n14103, ZN => n17525);
   U13611 : BUF_X2 port map( I => n14103, Z => n25733);
   U13613 : INV_X1 port map( I => n11785, ZN => n15268);
   U13617 : OR2_X2 port map( A1 => n25283, A2 => n10650, Z => n27423);
   U13623 : AND2_X2 port map( A1 => n20239, A2 => n20183, Z => n10650);
   U13627 : BUF_X2 port map( I => n19978, Z => n183);
   U13628 : NAND2_X1 port map( A1 => n22887, A2 => n1416, ZN => n28463);
   U13630 : INV_X2 port map( I => n4309, ZN => n18424);
   U13634 : NAND2_X1 port map( A1 => n28205, A2 => n25882, ZN => n27424);
   U13635 : NOR2_X1 port map( A1 => n22057, A2 => n9494, ZN => n21226);
   U13637 : OR2_X2 port map( A1 => n21212, A2 => n9494, Z => n9493);
   U13642 : INV_X1 port map( I => n9494, ZN => n22027);
   U13644 : NOR2_X1 port map( A1 => n2377, A2 => n1037, ZN => n28065);
   U13645 : XNOR2_X1 port map( A1 => n12481, A2 => n16938, ZN => n24154);
   U13647 : NAND2_X2 port map( A1 => n4912, A2 => n4911, ZN => n27425);
   U13648 : XOR2_X1 port map( A1 => n15213, A2 => n27735, Z => n27428);
   U13659 : OAI22_X1 port map( A1 => n21479, A2 => n21483, B1 => n11624, B2 => 
                           n11623, ZN => n27554);
   U13660 : INV_X1 port map( I => n13610, ZN => n15003);
   U13661 : INV_X2 port map( I => n13056, ZN => n28213);
   U13665 : NAND2_X1 port map( A1 => n21446, A2 => n15094, ZN => n27518);
   U13667 : NAND3_X1 port map( A1 => n25277, A2 => n3549, A3 => n21446, ZN => 
                           n7377);
   U13668 : NAND2_X1 port map( A1 => n18581, A2 => n18580, ZN => n27712);
   U13672 : NOR2_X1 port map( A1 => n18791, A2 => n12584, ZN => n18889);
   U13674 : NOR2_X1 port map( A1 => n19163, A2 => n19164, ZN => n28309);
   U13677 : NOR2_X1 port map( A1 => n17513, A2 => n17514, ZN => n7245);
   U13682 : NAND2_X1 port map( A1 => n6181, A2 => n6182, ZN => n14032);
   U13683 : NOR2_X1 port map( A1 => n952, A2 => n5721, ZN => n2570);
   U13689 : NOR2_X1 port map( A1 => n15314, A2 => n20408, ZN => n2321);
   U13690 : XNOR2_X1 port map( A1 => n6241, A2 => n18019, ZN => n27430);
   U13691 : NAND2_X1 port map( A1 => n22129, A2 => n27373, ZN => n2519);
   U13692 : BUF_X2 port map( I => n12711, Z => n5192);
   U13698 : INV_X1 port map( I => n26001, ZN => n20981);
   U13702 : AOI21_X1 port map( A1 => n7364, A2 => n334, B => n12712, ZN => 
                           n20495);
   U13704 : INV_X1 port map( I => n26059, ZN => n26333);
   U13705 : NAND2_X1 port map( A1 => n12206, A2 => n27091, ZN => n5292);
   U13706 : CLKBUF_X4 port map( I => n14501, Z => n24243);
   U13710 : NAND2_X1 port map( A1 => n27013, A2 => n2544, ZN => n20328);
   U13712 : AOI21_X1 port map( A1 => n14358, A2 => n22019, B => n10480, ZN => 
                           n11841);
   U13713 : XOR2_X1 port map( A1 => n9332, A2 => n644, Z => n27433);
   U13715 : NAND2_X1 port map( A1 => n20143, A2 => n20107, ZN => n20206);
   U13718 : NOR2_X1 port map( A1 => n21700, A2 => n945, ZN => n15627);
   U13720 : NAND2_X1 port map( A1 => n14892, A2 => n25368, ZN => n1819);
   U13721 : AOI21_X1 port map( A1 => n19152, A2 => n14925, B => n25368, ZN => 
                           n15621);
   U13725 : INV_X1 port map( I => n20979, ZN => n20977);
   U13730 : NAND2_X1 port map( A1 => n11553, A2 => n18798, ZN => n27775);
   U13732 : AND2_X1 port map( A1 => n7067, A2 => n8963, Z => n20864);
   U13733 : AOI21_X1 port map( A1 => n14545, A2 => n6778, B => n19106, ZN => 
                           n22514);
   U13738 : NAND2_X1 port map( A1 => n14580, A2 => n6906, ZN => n18997);
   U13750 : NAND3_X1 port map( A1 => n9354, A2 => n14580, A3 => n19090, ZN => 
                           n27817);
   U13752 : CLKBUF_X2 port map( I => n14580, Z => n24306);
   U13754 : OR3_X2 port map( A1 => n17873, A2 => n22253, A3 => n26643, Z => 
                           n10073);
   U13757 : NOR2_X1 port map( A1 => n26643, A2 => n22253, ZN => n2725);
   U13761 : INV_X1 port map( I => n26643, ZN => n13187);
   U13765 : NAND2_X1 port map( A1 => n8656, A2 => n1699, ZN => n24209);
   U13767 : NOR2_X1 port map( A1 => n15287, A2 => n4822, ZN => n13086);
   U13768 : AND2_X2 port map( A1 => n19100, A2 => n11692, Z => n27434);
   U13770 : NAND2_X1 port map( A1 => n18924, A2 => n14502, ZN => n1818);
   U13771 : NOR2_X1 port map( A1 => n27404, A2 => n9611, ZN => n13922);
   U13773 : CLKBUF_X4 port map( I => n7582, Z => n204);
   U13774 : NAND2_X1 port map( A1 => n22385, A2 => n28237, ZN => n19081);
   U13779 : AOI21_X1 port map( A1 => n10488, A2 => n11205, B => n24146, ZN => 
                           n5206);
   U13780 : INV_X2 port map( I => n21406, ZN => n21409);
   U13781 : INV_X1 port map( I => n19535, ZN => n1359);
   U13792 : NOR2_X1 port map( A1 => n2701, A2 => n9050, ZN => n1446);
   U13794 : NAND2_X1 port map( A1 => n25809, A2 => n28176, ZN => n10000);
   U13797 : NAND2_X1 port map( A1 => n27667, A2 => n25668, ZN => n27435);
   U13799 : NAND2_X1 port map( A1 => n17560, A2 => n17559, ZN => n3225);
   U13808 : NAND2_X1 port map( A1 => n13607, A2 => n17560, ZN => n17366);
   U13809 : CLKBUF_X4 port map( I => n8386, Z => n7904);
   U13811 : AND2_X2 port map( A1 => n16538, A2 => n16493, Z => n25397);
   U13812 : XOR2_X1 port map( A1 => n3331, A2 => n8450, Z => n27436);
   U13813 : OAI21_X2 port map( A1 => n14646, A2 => n8508, B => n8506, ZN => 
                           n27437);
   U13814 : OAI21_X1 port map( A1 => n14646, A2 => n8508, B => n8506, ZN => 
                           n5623);
   U13818 : NOR2_X2 port map( A1 => n24691, A2 => n13652, ZN => n27438);
   U13819 : NAND2_X1 port map( A1 => n21087, A2 => n21083, ZN => n21084);
   U13820 : AND2_X2 port map( A1 => n15891, A2 => n25224, Z => n10728);
   U13833 : CLKBUF_X12 port map( I => n15891, Z => n22454);
   U13835 : NAND3_X1 port map( A1 => n19821, A2 => n11175, A3 => n11110, ZN => 
                           n9266);
   U13836 : NAND2_X1 port map( A1 => n964, A2 => n11110, ZN => n7042);
   U13839 : NAND2_X2 port map( A1 => n26580, A2 => n11560, ZN => n7296);
   U13841 : AND3_X1 port map( A1 => n25526, A2 => n15002, A3 => n25525, Z => 
                           n27441);
   U13843 : NAND2_X1 port map( A1 => n2346, A2 => n4549, ZN => n15326);
   U13844 : INV_X1 port map( I => n21498, ZN => n27442);
   U13846 : INV_X1 port map( I => n7463, ZN => n3835);
   U13850 : CLKBUF_X12 port map( I => n22202, Z => n21998);
   U13854 : INV_X4 port map( I => n28225, ZN => n27443);
   U13855 : NAND2_X1 port map( A1 => n615, A2 => n7269, ZN => n2713);
   U13857 : NAND2_X1 port map( A1 => n10981, A2 => n16556, ZN => n12329);
   U13867 : OAI22_X2 port map( A1 => n8829, A2 => n19031, B1 => n8828, B2 => 
                           n19032, ZN => n27444);
   U13871 : OAI22_X1 port map( A1 => n8829, A2 => n19031, B1 => n8828, B2 => 
                           n19032, ZN => n12939);
   U13878 : NAND2_X1 port map( A1 => n15986, A2 => n15983, ZN => n15985);
   U13882 : NAND2_X2 port map( A1 => n21620, A2 => n26435, ZN => n11738);
   U13886 : NOR2_X1 port map( A1 => n21456, A2 => n21619, ZN => n12476);
   U13892 : XOR2_X1 port map( A1 => n23010, A2 => n9650, Z => n27446);
   U13893 : NOR2_X2 port map( A1 => n24709, A2 => n22596, ZN => n27447);
   U13897 : OAI22_X2 port map( A1 => n18840, A2 => n18839, B1 => n18896, B2 => 
                           n11577, ZN => n27448);
   U13899 : CLKBUF_X12 port map( I => n12208, Z => n357);
   U13903 : INV_X1 port map( I => n23779, ZN => n27449);
   U13905 : NOR2_X1 port map( A1 => n13674, A2 => n17036, ZN => n5579);
   U13906 : OAI21_X1 port map( A1 => n17036, A2 => n9865, B => n17413, ZN => 
                           n10912);
   U13907 : INV_X2 port map( I => n17036, ZN => n17315);
   U13908 : XOR2_X1 port map( A1 => n18061, A2 => n5413, Z => n27451);
   U13909 : NAND3_X2 port map( A1 => n18102, A2 => n14984, A3 => n17760, ZN => 
                           n5413);
   U13915 : INV_X2 port map( I => n6485, ZN => n11923);
   U13919 : INV_X1 port map( I => n19254, ZN => n13167);
   U13925 : CLKBUF_X2 port map( I => n19254, Z => n19730);
   U13930 : INV_X2 port map( I => n8646, ZN => n14188);
   U13941 : CLKBUF_X12 port map( I => n19932, Z => n27452);
   U13944 : BUF_X1 port map( I => n4518, Z => n162);
   U13952 : XOR2_X1 port map( A1 => n13370, A2 => n18266, Z => n27453);
   U13953 : NAND2_X1 port map( A1 => n12046, A2 => n12186, ZN => n20999);
   U13959 : INV_X2 port map( I => n19116, ZN => n25770);
   U13960 : NAND2_X1 port map( A1 => n17867, A2 => n7321, ZN => n14167);
   U13962 : OAI21_X1 port map( A1 => n23357, A2 => n23356, B => n7321, ZN => 
                           n23475);
   U13963 : INV_X1 port map( I => n2404, ZN => n27456);
   U13966 : NOR2_X1 port map( A1 => n18793, A2 => n23305, ZN => n23793);
   U13968 : CLKBUF_X2 port map( I => n18793, Z => n992);
   U13970 : NAND2_X2 port map( A1 => n18793, A2 => n18396, ZN => n18795);
   U13975 : INV_X1 port map( I => n10640, ZN => n27457);
   U13981 : NOR3_X1 port map( A1 => n725, A2 => n9040, A3 => n17766, ZN => 
                           n17702);
   U13983 : NAND2_X1 port map( A1 => n9040, A2 => n17766, ZN => n17264);
   U13986 : AND2_X2 port map( A1 => n26476, A2 => n26197, Z => n27458);
   U13990 : OR2_X2 port map( A1 => n28248, A2 => n27647, Z => n22949);
   U14001 : CLKBUF_X12 port map( I => n15353, Z => n2813);
   U14003 : NAND2_X1 port map( A1 => n20088, A2 => n27347, ZN => n10028);
   U14006 : NAND2_X1 port map( A1 => n27367, A2 => n16707, ZN => n16705);
   U14012 : AND2_X1 port map( A1 => n13411, A2 => n8546, Z => n17416);
   U14013 : CLKBUF_X12 port map( I => n13411, Z => n193);
   U14014 : BUF_X2 port map( I => n18660, Z => n8022);
   U14029 : INV_X1 port map( I => n18660, ZN => n26292);
   U14034 : NAND2_X2 port map( A1 => n28469, A2 => n28351, ZN => n27460);
   U14041 : NAND2_X1 port map( A1 => n12191, A2 => n21166, ZN => n21169);
   U14043 : NAND2_X1 port map( A1 => n936, A2 => n21166, ZN => n4307);
   U14052 : AND2_X1 port map( A1 => n562, A2 => n15964, Z => n16256);
   U14057 : AND2_X2 port map( A1 => n18715, A2 => n15366, Z => n4290);
   U14074 : INV_X1 port map( I => n15624, ZN => n21725);
   U14076 : XNOR2_X1 port map( A1 => n12242, A2 => n12771, ZN => n27461);
   U14077 : NAND2_X1 port map( A1 => n26720, A2 => n23772, ZN => n7814);
   U14078 : BUF_X2 port map( I => n26001, Z => n24040);
   U14082 : NAND2_X1 port map( A1 => n11983, A2 => n5511, ZN => n10229);
   U14086 : NOR2_X1 port map( A1 => n7568, A2 => n6778, ZN => n26167);
   U14093 : NAND2_X1 port map( A1 => n8226, A2 => n6778, ZN => n27522);
   U14111 : NOR2_X1 port map( A1 => n7908, A2 => n7749, ZN => n1410);
   U14114 : OAI22_X1 port map( A1 => n9288, A2 => n25255, B1 => n9726, B2 => 
                           n16587, ZN => n27462);
   U14119 : OAI22_X1 port map( A1 => n9288, A2 => n25255, B1 => n9726, B2 => 
                           n16587, ZN => n27463);
   U14125 : OAI22_X1 port map( A1 => n9288, A2 => n25255, B1 => n9726, B2 => 
                           n16587, ZN => n10187);
   U14126 : INV_X1 port map( I => n7965, ZN => n10579);
   U14127 : CLKBUF_X12 port map( I => n7965, Z => n288);
   U14131 : NAND2_X1 port map( A1 => n3852, A2 => n5131, ZN => n27464);
   U14133 : NAND2_X1 port map( A1 => n3852, A2 => n5131, ZN => n27465);
   U14141 : NAND2_X1 port map( A1 => n3852, A2 => n5131, ZN => n19114);
   U14144 : NOR2_X1 port map( A1 => n26140, A2 => n20072, ZN => n1956);
   U14146 : CLKBUF_X12 port map( I => n12571, Z => n23920);
   U14152 : XOR2_X1 port map( A1 => n7598, A2 => n8608, Z => n27466);
   U14156 : XOR2_X1 port map( A1 => n4965, A2 => n23589, Z => n27467);
   U14159 : NAND2_X2 port map( A1 => n26004, A2 => n13554, ZN => n27468);
   U14163 : NAND2_X2 port map( A1 => n20854, A2 => n20855, ZN => n13554);
   U14165 : XNOR2_X1 port map( A1 => n1801, A2 => Plaintext(19), ZN => n27469);
   U14166 : XOR2_X1 port map( A1 => n25166, A2 => n5698, Z => n27470);
   U14167 : INV_X2 port map( I => Key(19), ZN => n1801);
   U14170 : OR3_X2 port map( A1 => n8896, A2 => n24278, A3 => n10598, Z => 
                           n27471);
   U14174 : NAND3_X1 port map( A1 => n7342, A2 => n28176, A3 => n13234, ZN => 
                           n20681);
   U14175 : NAND3_X1 port map( A1 => n20145, A2 => n23212, A3 => n19, ZN => 
                           n6969);
   U14189 : NAND2_X1 port map( A1 => n19, A2 => n23212, ZN => n9919);
   U14191 : INV_X2 port map( I => n23212, ZN => n20071);
   U14193 : AND2_X2 port map( A1 => n6185, A2 => n27662, Z => n6183);
   U14194 : NAND2_X1 port map( A1 => n13528, A2 => n16572, ZN => n1761);
   U14196 : NAND2_X1 port map( A1 => n16573, A2 => n16572, ZN => n13605);
   U14197 : NOR3_X1 port map( A1 => n14974, A2 => n20196, A3 => n14975, ZN => 
                           n14973);
   U14204 : NAND2_X1 port map( A1 => n15732, A2 => n20286, ZN => n24496);
   U14205 : NAND2_X1 port map( A1 => n15732, A2 => n19989, ZN => n19987);
   U14211 : NOR2_X1 port map( A1 => n25738, A2 => n8000, ZN => n2271);
   U14212 : AOI22_X1 port map( A1 => n3724, A2 => n1431, B1 => n25003, B2 => 
                           n3725, ZN => n3406);
   U14213 : NAND3_X1 port map( A1 => n937, A2 => n13395, A3 => n14583, ZN => 
                           n2007);
   U14216 : OAI22_X2 port map( A1 => n18944, A2 => n4212, B1 => n18943, B2 => 
                           n12896, ZN => n25259);
   U14218 : NAND3_X1 port map( A1 => n27901, A2 => n5353, A3 => n26227, ZN => 
                           n28391);
   U14221 : XOR2_X1 port map( A1 => n18212, A2 => n4777, Z => n3581);
   U14223 : XOR2_X1 port map( A1 => n4901, A2 => n18085, Z => n13960);
   U14224 : AND3_X2 port map( A1 => n16044, A2 => n16042, A3 => n16043, Z => 
                           n27472);
   U14227 : AOI22_X2 port map( A1 => n24847, A2 => n4661, B1 => n28481, B2 => 
                           n13963, ZN => n7737);
   U14228 : AOI21_X2 port map( A1 => n4537, A2 => n859, B => n20171, ZN => 
                           n28333);
   U14229 : XOR2_X1 port map( A1 => n6528, A2 => n13752, Z => n19518);
   U14230 : NAND2_X2 port map( A1 => n9215, A2 => n7994, ZN => n6528);
   U14240 : NAND3_X1 port map( A1 => n25087, A2 => n11092, A3 => n11093, ZN => 
                           n27473);
   U14241 : XOR2_X1 port map( A1 => n21298, A2 => n1611, Z => n20334);
   U14251 : AOI22_X2 port map( A1 => n24102, A2 => n28068, B1 => n19862, B2 => 
                           n19914, ZN => n23159);
   U14259 : XOR2_X1 port map( A1 => n27474, A2 => n10711, Z => n14065);
   U14263 : XOR2_X1 port map( A1 => n18198, A2 => n18197, Z => n27474);
   U14266 : XOR2_X1 port map( A1 => n18331, A2 => n18123, Z => n4681);
   U14276 : AOI22_X2 port map( A1 => n17777, A2 => n17776, B1 => n17775, B2 => 
                           n23915, ZN => n18123);
   U14279 : AOI22_X2 port map( A1 => n20586, A2 => n20781, B1 => n21936, B2 => 
                           n15689, ZN => n9074);
   U14280 : NOR2_X2 port map( A1 => n13188, A2 => n24575, ZN => n20586);
   U14287 : NAND2_X1 port map( A1 => n27958, A2 => n17515, ZN => n27901);
   U14290 : NAND2_X2 port map( A1 => n1408, A2 => n27475, ZN => n20282);
   U14291 : NAND2_X2 port map( A1 => n19008, A2 => n22391, ZN => n9236);
   U14292 : NAND2_X2 port map( A1 => n27499, A2 => n24864, ZN => n22391);
   U14297 : XOR2_X1 port map( A1 => n27476, A2 => n21430, Z => n5550);
   U14299 : XOR2_X1 port map( A1 => n9125, A2 => n25748, Z => n27476);
   U14303 : INV_X2 port map( I => n10574, ZN => n9994);
   U14305 : XOR2_X1 port map( A1 => n6664, A2 => n11709, Z => n10574);
   U14314 : NOR2_X2 port map( A1 => n27477, A2 => n20157, ZN => n8366);
   U14318 : NOR2_X1 port map( A1 => n14399, A2 => n14398, ZN => n27477);
   U14319 : NOR2_X2 port map( A1 => n27478, A2 => n11366, ZN => n5229);
   U14326 : XOR2_X1 port map( A1 => n14659, A2 => n4204, Z => n5868);
   U14327 : NAND2_X2 port map( A1 => n21986, A2 => n7381, ZN => n4204);
   U14334 : XOR2_X1 port map( A1 => n18047, A2 => n3613, Z => n18136);
   U14335 : NAND2_X2 port map( A1 => n5894, A2 => n5896, ZN => n18047);
   U14338 : NOR3_X2 port map( A1 => n11223, A2 => n14695, A3 => n22798, ZN => 
                           n2561);
   U14340 : AOI22_X2 port map( A1 => n6368, A2 => n9132, B1 => n1030, B2 => 
                           n6367, ZN => n5305);
   U14351 : INV_X2 port map( I => n4119, ZN => n4246);
   U14358 : XOR2_X1 port map( A1 => n15213, A2 => n27735, Z => n4119);
   U14361 : NAND3_X2 port map( A1 => n28130, A2 => n19906, A3 => n19907, ZN => 
                           n27479);
   U14364 : NAND2_X2 port map( A1 => n27485, A2 => n13186, ZN => n4683);
   U14367 : INV_X4 port map( I => n7652, ZN => n28104);
   U14369 : INV_X2 port map( I => n27480, ZN => n4901);
   U14370 : OAI21_X2 port map( A1 => n10114, A2 => n24657, B => n10112, ZN => 
                           n2225);
   U14373 : XOR2_X1 port map( A1 => n23567, A2 => n27481, Z => n17160);
   U14378 : XOR2_X1 port map( A1 => n10191, A2 => n16982, Z => n27481);
   U14383 : NAND2_X2 port map( A1 => n27482, A2 => n23067, ZN => n3725);
   U14389 : OAI21_X2 port map( A1 => n20558, A2 => n20557, B => n7341, ZN => 
                           n27482);
   U14397 : NOR2_X2 port map( A1 => n23542, A2 => n27483, ZN => n14035);
   U14400 : OAI22_X2 port map( A1 => n7631, A2 => n9769, B1 => n16241, B2 => 
                           n16312, ZN => n27485);
   U14402 : NOR2_X2 port map( A1 => n27487, A2 => n27486, ZN => n25084);
   U14413 : XOR2_X1 port map( A1 => n18071, A2 => n7764, Z => n23359);
   U14416 : NAND2_X2 port map( A1 => n1428, A2 => n23232, ZN => n7764);
   U14422 : XOR2_X1 port map( A1 => n17110, A2 => n27488, Z => n17112);
   U14430 : XOR2_X1 port map( A1 => n11124, A2 => n17109, Z => n27488);
   U14431 : OAI22_X2 port map( A1 => n14022, A2 => n5115, B1 => n27871, B2 => 
                           n18645, ZN => n18761);
   U14432 : AOI21_X2 port map( A1 => n14735, A2 => n14734, B => n4929, ZN => 
                           n4928);
   U14434 : NAND2_X2 port map( A1 => n26687, A2 => n26231, ZN => n14735);
   U14435 : NAND3_X1 port map( A1 => n15398, A2 => n15397, A3 => n18705, ZN => 
                           n27616);
   U14438 : XOR2_X1 port map( A1 => n13890, A2 => n18282, Z => n9292);
   U14439 : NOR3_X1 port map( A1 => n14427, A2 => n11262, A3 => n18432, ZN => 
                           n25066);
   U14452 : INV_X2 port map( I => n25955, ZN => n18432);
   U14453 : OAI22_X2 port map( A1 => n1084, A2 => n21160, B1 => n9005, B2 => 
                           n11905, ZN => n28260);
   U14454 : XOR2_X1 port map( A1 => n27490, A2 => n14800, Z => n2311);
   U14456 : XOR2_X1 port map( A1 => n27243, A2 => n25933, Z => n27490);
   U14458 : NAND2_X1 port map( A1 => n27491, A2 => n21047, ZN => n14954);
   U14463 : INV_X1 port map( I => n21045, ZN => n27491);
   U14464 : NOR2_X2 port map( A1 => n21040, A2 => n22797, ZN => n21045);
   U14467 : XOR2_X1 port map( A1 => n4204, A2 => n18066, Z => n18335);
   U14468 : OAI21_X2 port map( A1 => n7894, A2 => n8307, B => n27493, ZN => 
                           n24862);
   U14470 : AOI22_X2 port map( A1 => n23075, A2 => n7793, B1 => n7893, B2 => 
                           n724, ZN => n27493);
   U14483 : BUF_X2 port map( I => n10007, Z => n27494);
   U14486 : XOR2_X1 port map( A1 => n27495, A2 => n28344, Z => n421);
   U14487 : XOR2_X1 port map( A1 => n18229, A2 => n25681, Z => n27495);
   U14491 : INV_X2 port map( I => n20847, ZN => n20827);
   U14492 : NAND3_X2 port map( A1 => n20813, A2 => n20812, A3 => n27584, ZN => 
                           n20847);
   U14494 : XOR2_X1 port map( A1 => n4920, A2 => n4918, Z => n24228);
   U14496 : AOI22_X1 port map( A1 => n28409, A2 => n22427, B1 => n10664, B2 => 
                           n13161, ZN => n27511);
   U14497 : NAND2_X2 port map( A1 => n27496, A2 => n26387, ZN => n5395);
   U14501 : OAI22_X2 port map( A1 => n17871, A2 => n17898, B1 => n21768, B2 => 
                           n14278, ZN => n17900);
   U14502 : NAND2_X2 port map( A1 => n12852, A2 => n12851, ZN => n12046);
   U14506 : AOI22_X2 port map( A1 => n3344, A2 => n1090, B1 => n20976, B2 => 
                           n10661, ZN => n12851);
   U14507 : NAND2_X2 port map( A1 => n28163, A2 => n12843, ZN => n27498);
   U14508 : NAND3_X1 port map( A1 => n7578, A2 => n7577, A3 => n26031, ZN => 
                           n27499);
   U14513 : NAND2_X1 port map( A1 => n10430, A2 => n20604, ZN => n25675);
   U14515 : NOR2_X2 port map( A1 => n27500, A2 => n19474, ZN => n7183);
   U14522 : INV_X2 port map( I => n27501, ZN => n8546);
   U14523 : XOR2_X1 port map( A1 => n8548, A2 => n8549, Z => n27501);
   U14527 : XOR2_X1 port map( A1 => n26761, A2 => n17049, Z => n17096);
   U14531 : AOI21_X2 port map( A1 => n24583, A2 => n16760, B => n465, ZN => 
                           n17049);
   U14533 : XOR2_X1 port map( A1 => n27502, A2 => n19456, Z => n27796);
   U14535 : XOR2_X1 port map( A1 => n27615, A2 => n27503, Z => n27502);
   U14536 : XOR2_X1 port map( A1 => n27504, A2 => n21367, Z => Ciphertext(100))
                           ;
   U14541 : XOR2_X1 port map( A1 => n26469, A2 => n7409, Z => n24035);
   U14543 : NAND2_X2 port map( A1 => n12711, A2 => n11160, ZN => n13726);
   U14554 : OAI21_X2 port map( A1 => n27505, A2 => n21841, B => n874, ZN => 
                           n13239);
   U14556 : NOR2_X2 port map( A1 => n1158, A2 => n11718, ZN => n27505);
   U14559 : XOR2_X1 port map( A1 => n13449, A2 => n14619, Z => n18036);
   U14560 : OAI21_X2 port map( A1 => n27507, A2 => n5621, B => n18672, ZN => 
                           n19110);
   U14562 : AOI21_X2 port map( A1 => n9205, A2 => n9204, B => n27508, ZN => 
                           n9203);
   U14569 : XOR2_X1 port map( A1 => n6582, A2 => n10191, Z => n7949);
   U14572 : OAI22_X2 port map( A1 => n9822, A2 => n767, B1 => n62, B2 => n17026
                           , ZN => n6582);
   U14577 : NAND2_X2 port map( A1 => n12872, A2 => n27509, ZN => n14601);
   U14580 : XOR2_X1 port map( A1 => n27511, A2 => n21594, Z => Ciphertext(156))
                           ;
   U14581 : BUF_X2 port map( I => n20976, Z => n27512);
   U14589 : XOR2_X1 port map( A1 => n18353, A2 => n7338, Z => n18316);
   U14590 : XOR2_X1 port map( A1 => n27513, A2 => n17077, Z => n13658);
   U14592 : NAND2_X2 port map( A1 => n16033, A2 => n16032, ZN => n17077);
   U14594 : OR3_X1 port map( A1 => n26001, A2 => n15004, A3 => n26924, Z => 
                           n27977);
   U14595 : XOR2_X1 port map( A1 => n17067, A2 => n27514, Z => n13519);
   U14611 : XOR2_X1 port map( A1 => n17068, A2 => n2265, Z => n27514);
   U14612 : NAND2_X2 port map( A1 => n27515, A2 => n26331, ZN => n11553);
   U14614 : XOR2_X1 port map( A1 => n26279, A2 => n19228, Z => n25005);
   U14628 : XOR2_X1 port map( A1 => n19334, A2 => n19482, Z => n19228);
   U14630 : XOR2_X1 port map( A1 => n17038, A2 => n7786, Z => n25184);
   U14632 : NOR2_X2 port map( A1 => n16416, A2 => n14698, ZN => n17038);
   U14633 : NAND3_X1 port map( A1 => n21002, A2 => n21005, A3 => n13961, ZN => 
                           n14458);
   U14639 : INV_X2 port map( I => n24764, ZN => n21005);
   U14640 : NAND2_X2 port map( A1 => n24765, A2 => n20562, ZN => n24764);
   U14641 : NAND2_X1 port map( A1 => n9202, A2 => n16535, ZN => n5915);
   U14642 : XOR2_X1 port map( A1 => n27516, A2 => n657, Z => n14391);
   U14644 : XOR2_X1 port map( A1 => n22750, A2 => n5852, Z => n27516);
   U14649 : NOR2_X2 port map( A1 => n23923, A2 => n17687, ZN => n13621);
   U14651 : NAND2_X2 port map( A1 => n15406, A2 => n15407, ZN => n13515);
   U14661 : XOR2_X1 port map( A1 => n22849, A2 => n17104, Z => n15190);
   U14662 : AOI22_X2 port map( A1 => n9792, A2 => n16136, B1 => n16134, B2 => 
                           n16135, ZN => n10457);
   U14667 : INV_X1 port map( I => n27517, ZN => n6586);
   U14670 : NAND3_X2 port map( A1 => n27587, A2 => n12376, A3 => n8574, ZN => 
                           n8573);
   U14672 : XOR2_X1 port map( A1 => n19498, A2 => n19449, Z => n25618);
   U14673 : XOR2_X1 port map( A1 => n17028, A2 => n17084, Z => n16936);
   U14674 : OAI22_X2 port map( A1 => n16714, A2 => n16432, B1 => n28039, B2 => 
                           n3297, ZN => n17084);
   U14676 : XOR2_X1 port map( A1 => n27520, A2 => n21336, Z => Ciphertext(120))
                           ;
   U14681 : NAND2_X1 port map( A1 => n14927, A2 => n14225, ZN => n27520);
   U14686 : NAND3_X2 port map( A1 => n25714, A2 => n26023, A3 => n15310, ZN => 
                           n4366);
   U14687 : INV_X1 port map( I => n18336, ZN => n27770);
   U14692 : OAI22_X2 port map( A1 => n5195, A2 => n25315, B1 => n842, B2 => 
                           n20609, ZN => n6353);
   U14694 : INV_X2 port map( I => n20608, ZN => n842);
   U14696 : NAND2_X2 port map( A1 => n6355, A2 => n13310, ZN => n20608);
   U14698 : OR2_X1 port map( A1 => n16602, A2 => n16604, Z => n4059);
   U14699 : NAND2_X2 port map( A1 => n27523, A2 => n26362, ZN => n17277);
   U14701 : NOR2_X2 port map( A1 => n26361, A2 => n1224, ZN => n27523);
   U14706 : NAND2_X2 port map( A1 => n27586, A2 => n3887, ZN => n28547);
   U14708 : XOR2_X1 port map( A1 => n27524, A2 => n21211, Z => Ciphertext(108))
                           ;
   U14714 : AOI22_X1 port map( A1 => n24973, A2 => n10217, B1 => n26311, B2 => 
                           n5350, ZN => n27524);
   U14715 : OAI21_X2 port map( A1 => n10009, A2 => n18625, B => n14308, ZN => 
                           n10008);
   U14716 : NOR2_X1 port map( A1 => n1440, A2 => n18527, ZN => n18625);
   U14717 : OR2_X1 port map( A1 => n14442, A2 => n16273, Z => n2495);
   U14718 : OAI21_X2 port map( A1 => n22373, A2 => n26054, B => n27525, ZN => 
                           n12365);
   U14723 : XOR2_X1 port map( A1 => n20371, A2 => n20370, Z => n25502);
   U14724 : OR2_X1 port map( A1 => n19468, A2 => n19827, Z => n19685);
   U14725 : XOR2_X1 port map( A1 => n14856, A2 => n15173, Z => n24379);
   U14729 : INV_X4 port map( I => n27972, ZN => n18953);
   U14732 : XOR2_X1 port map( A1 => n7831, A2 => n27526, Z => n9911);
   U14734 : XOR2_X1 port map( A1 => n7833, A2 => n7830, Z => n27526);
   U14736 : NOR2_X2 port map( A1 => n27527, A2 => n14702, ZN => n28042);
   U14738 : NAND2_X2 port map( A1 => n1158, A2 => n11718, ZN => n27527);
   U14748 : XOR2_X1 port map( A1 => n18074, A2 => n5742, Z => n9274);
   U14751 : NAND2_X2 port map( A1 => n5349, A2 => n25476, ZN => n18074);
   U14752 : XOR2_X1 port map( A1 => n6275, A2 => n3372, Z => n8);
   U14753 : OR2_X1 port map( A1 => n5752, A2 => n22718, Z => n11309);
   U14755 : XOR2_X1 port map( A1 => n18276, A2 => n27529, Z => n2029);
   U14761 : XOR2_X1 port map( A1 => n2031, A2 => n18071, Z => n27529);
   U14762 : INV_X2 port map( I => n27867, ZN => n647);
   U14763 : NOR2_X2 port map( A1 => n17185, A2 => n17345, ZN => n17575);
   U14766 : OR2_X1 port map( A1 => n11982, A2 => n28309, Z => n23936);
   U14769 : INV_X2 port map( I => n4315, ZN => n20609);
   U14770 : NAND2_X2 port map( A1 => n9973, A2 => n9972, ZN => n4315);
   U14773 : XOR2_X1 port map( A1 => n15069, A2 => n25075, Z => n25547);
   U14780 : BUF_X2 port map( I => n25338, Z => n27530);
   U14792 : XOR2_X1 port map( A1 => n27531, A2 => n21709, Z => Ciphertext(184))
                           ;
   U14794 : NOR2_X2 port map( A1 => n11216, A2 => n11217, ZN => n26110);
   U14795 : NAND2_X2 port map( A1 => n15122, A2 => n15121, ZN => n11216);
   U14797 : NOR3_X2 port map( A1 => n1658, A2 => n2356, A3 => n14545, ZN => 
                           n23183);
   U14798 : OR2_X2 port map( A1 => n11809, A2 => n14501, Z => n10642);
   U14799 : OAI22_X1 port map( A1 => n20988, A2 => n27822, B1 => n11345, B2 => 
                           n21001, ZN => n24276);
   U14801 : NAND2_X2 port map( A1 => n27532, A2 => n3877, ZN => n18066);
   U14805 : NAND2_X2 port map( A1 => n2388, A2 => n17713, ZN => n27532);
   U14806 : XOR2_X1 port map( A1 => n6175, A2 => n2311, Z => n22620);
   U14807 : NOR2_X2 port map( A1 => n13167, A2 => n27445, ZN => n19845);
   U14808 : XOR2_X1 port map( A1 => n28084, A2 => n18309, Z => n27533);
   U14809 : XOR2_X1 port map( A1 => n9357, A2 => n18240, Z => n1649);
   U14811 : NAND2_X1 port map( A1 => n815, A2 => n7182, ZN => n8359);
   U14812 : NOR2_X2 port map( A1 => n8854, A2 => n8852, ZN => n27534);
   U14816 : NAND2_X2 port map( A1 => n27535, A2 => n23732, ZN => n11997);
   U14818 : AOI21_X2 port map( A1 => n4471, A2 => n24664, B => n27536, ZN => 
                           n27535);
   U14821 : NAND3_X1 port map( A1 => n8658, A2 => n17942, A3 => n237, ZN => 
                           n12943);
   U14824 : NAND2_X2 port map( A1 => n19835, A2 => n811, ZN => n27537);
   U14827 : NOR3_X2 port map( A1 => n21961, A2 => n27538, A3 => n8463, ZN => 
                           n14554);
   U14828 : NOR3_X1 port map( A1 => n811, A2 => n11078, A3 => n14343, ZN => 
                           n27538);
   U14829 : NAND2_X2 port map( A1 => n4731, A2 => n27539, ZN => n19477);
   U14833 : NAND2_X2 port map( A1 => n27541, A2 => n27540, ZN => n17974);
   U14837 : NAND2_X1 port map( A1 => n8108, A2 => n8107, ZN => n27541);
   U14842 : XOR2_X1 port map( A1 => n12926, A2 => n20459, Z => n21179);
   U14849 : NOR2_X2 port map( A1 => n12812, A2 => n28385, ZN => n12926);
   U14850 : XOR2_X1 port map( A1 => n27357, A2 => n19412, Z => n19441);
   U14851 : NAND2_X1 port map( A1 => n23709, A2 => n23782, ZN => n27542);
   U14852 : NAND2_X1 port map( A1 => n19063, A2 => n8998, ZN => n27544);
   U14853 : AND2_X1 port map( A1 => n28019, A2 => n18879, Z => n26014);
   U14857 : OAI21_X1 port map( A1 => n7525, A2 => n7735, B => n25873, ZN => 
                           n2345);
   U14858 : XOR2_X1 port map( A1 => n17129, A2 => n8997, Z => n295);
   U14859 : NOR3_X2 port map( A1 => n27852, A2 => n4812, A3 => n17925, ZN => 
                           n27545);
   U14869 : NOR2_X2 port map( A1 => n25374, A2 => n8423, ZN => n17208);
   U14870 : NAND2_X2 port map( A1 => n27546, A2 => n11907, ZN => n11906);
   U14872 : NAND2_X2 port map( A1 => n1020, A2 => n27640, ZN => n27547);
   U14873 : INV_X1 port map( I => n1824, ZN => n27571);
   U14879 : NOR2_X2 port map( A1 => n27549, A2 => n7328, ZN => n8280);
   U14880 : NOR2_X1 port map( A1 => n14377, A2 => n12712, ZN => n27549);
   U14882 : BUF_X2 port map( I => n24127, Z => n27550);
   U14884 : AOI21_X2 port map( A1 => n27918, A2 => n13872, B => n27551, ZN => 
                           n27917);
   U14885 : NOR2_X2 port map( A1 => n13872, A2 => n19135, ZN => n27551);
   U14889 : NAND2_X1 port map( A1 => n11471, A2 => n10291, ZN => n11236);
   U14891 : XOR2_X1 port map( A1 => n12414, A2 => n26517, Z => n6014);
   U14895 : XOR2_X1 port map( A1 => n25353, A2 => n2510, Z => n2509);
   U14896 : NAND2_X2 port map( A1 => n20113, A2 => n20112, ZN => n28272);
   U14904 : XOR2_X1 port map( A1 => n27554, A2 => n14492, Z => Ciphertext(141))
                           ;
   U14905 : XOR2_X1 port map( A1 => n19505, A2 => n27555, Z => n15156);
   U14908 : XOR2_X1 port map( A1 => n9985, A2 => n4303, Z => n27555);
   U14909 : OR2_X1 port map( A1 => n15462, A2 => n27556, Z => n17677);
   U14925 : BUF_X2 port map( I => n15268, Z => n27557);
   U14926 : BUF_X2 port map( I => n24190, Z => n27558);
   U14927 : OAI22_X2 port map( A1 => n10972, A2 => n17294, B1 => n25246, B2 => 
                           n195, ZN => n8472);
   U14928 : XOR2_X1 port map( A1 => n18297, A2 => n27559, Z => n22393);
   U14929 : XOR2_X1 port map( A1 => n6129, A2 => n27410, Z => n27559);
   U14930 : INV_X2 port map( I => n27560, ZN => n10206);
   U14931 : XNOR2_X1 port map( A1 => n23319, A2 => n6736, ZN => n27560);
   U14935 : NAND2_X1 port map( A1 => n20078, A2 => n9365, ZN => n20137);
   U14936 : NAND3_X2 port map( A1 => n15373, A2 => n28029, A3 => n19699, ZN => 
                           n20078);
   U14939 : NAND2_X1 port map( A1 => n22598, A2 => n22374, ZN => n2373);
   U14944 : XOR2_X1 port map( A1 => n25442, A2 => n18131, Z => n22659);
   U14945 : XOR2_X1 port map( A1 => n5868, A2 => n27410, Z => n18131);
   U14947 : XOR2_X1 port map( A1 => n18071, A2 => n28370, Z => n18334);
   U14948 : OAI21_X2 port map( A1 => n24091, A2 => n24566, B => n1037, ZN => 
                           n27561);
   U14953 : XOR2_X1 port map( A1 => n21432, A2 => n1912, Z => n20563);
   U14958 : NOR2_X2 port map( A1 => n24877, A2 => n20432, ZN => n21432);
   U14960 : NAND3_X2 port map( A1 => n17172, A2 => n3533, A3 => n894, ZN => 
                           n24007);
   U14966 : NAND3_X1 port map( A1 => n14945, A2 => n10461, A3 => n8125, ZN => 
                           n8804);
   U14967 : NOR2_X1 port map( A1 => n15916, A2 => n16306, ZN => n13877);
   U14975 : NAND3_X2 port map( A1 => n12157, A2 => n1118, A3 => n19802, ZN => 
                           n28493);
   U14977 : INV_X2 port map( I => n27563, ZN => n21863);
   U14993 : NAND2_X2 port map( A1 => n18694, A2 => n27361, ZN => n9198);
   U15001 : NOR2_X2 port map( A1 => n10388, A2 => n10389, ZN => n9952);
   U15004 : AOI21_X2 port map( A1 => n16154, A2 => n16701, B => n27565, ZN => 
                           n1763);
   U15005 : NOR2_X2 port map( A1 => n16467, A2 => n16469, ZN => n27565);
   U15008 : XNOR2_X1 port map( A1 => n3810, A2 => n16580, ZN => n28283);
   U15014 : OAI21_X2 port map( A1 => n12977, A2 => n12976, B => n27566, ZN => 
                           n23435);
   U15016 : NAND2_X2 port map( A1 => n10882, A2 => n7282, ZN => n27566);
   U15017 : NOR2_X2 port map( A1 => n27567, A2 => n22617, ZN => n26140);
   U15018 : INV_X2 port map( I => n23159, ZN => n27567);
   U15022 : INV_X2 port map( I => n27568, ZN => n16203);
   U15025 : XNOR2_X1 port map( A1 => n23845, A2 => Key(84), ZN => n27568);
   U15026 : XOR2_X1 port map( A1 => n19224, A2 => n4789, Z => n19093);
   U15032 : NAND2_X2 port map( A1 => n27966, A2 => n6533, ZN => n4789);
   U15033 : AND2_X1 port map( A1 => n20058, A2 => n6969, Z => n10168);
   U15034 : XOR2_X1 port map( A1 => n3688, A2 => n3684, Z => n27662);
   U15035 : BUF_X2 port map( I => n7030, Z => n27569);
   U15036 : OR2_X1 port map( A1 => n26712, A2 => n12046, Z => n27570);
   U15038 : NOR2_X1 port map( A1 => n28503, A2 => n28504, ZN => n14263);
   U15040 : NAND2_X2 port map( A1 => n20277, A2 => n287, ZN => n20217);
   U15041 : OAI21_X2 port map( A1 => n9452, A2 => n24026, B => n9453, ZN => 
                           n287);
   U15042 : NAND2_X2 port map( A1 => n17942, A2 => n4531, ZN => n27574);
   U15043 : NAND2_X2 port map( A1 => n11434, A2 => n11699, ZN => n17942);
   U15046 : AOI22_X2 port map( A1 => n10586, A2 => n950, B1 => n25326, B2 => 
                           n11306, ZN => n23872);
   U15048 : XOR2_X1 port map( A1 => n27575, A2 => n8890, Z => n5722);
   U15052 : XOR2_X1 port map( A1 => n2769, A2 => n7467, Z => n27575);
   U15055 : XOR2_X1 port map( A1 => n8848, A2 => n5771, Z => n3466);
   U15065 : NOR2_X2 port map( A1 => n27576, A2 => n25688, ZN => n12935);
   U15072 : AOI21_X2 port map( A1 => n5218, A2 => n3846, B => n27577, ZN => 
                           n27576);
   U15073 : XOR2_X1 port map( A1 => n28259, A2 => n17134, Z => n27655);
   U15076 : NAND2_X2 port map( A1 => n2597, A2 => n2596, ZN => n17134);
   U15078 : AOI21_X2 port map( A1 => n15548, A2 => n9202, B => n9517, ZN => 
                           n27599);
   U15083 : NAND3_X2 port map( A1 => n23671, A2 => n21510, A3 => n5509, ZN => 
                           n21538);
   U15085 : NAND3_X2 port map( A1 => n28091, A2 => n20308, A3 => n26365, ZN => 
                           n20003);
   U15088 : INV_X2 port map( I => n21124, ZN => n24951);
   U15093 : NAND2_X2 port map( A1 => n23728, A2 => n14870, ZN => n21124);
   U15097 : OAI21_X1 port map( A1 => n27579, A2 => n27578, B => n4428, ZN => 
                           n22585);
   U15098 : NOR2_X1 port map( A1 => n23976, A2 => n13472, ZN => n27578);
   U15101 : AOI22_X2 port map( A1 => n25008, A2 => n1687, B1 => n27581, B2 => 
                           n19925, ZN => n23212);
   U15103 : NAND3_X2 port map( A1 => n5731, A2 => n16428, A3 => n265, ZN => 
                           n5730);
   U15104 : XOR2_X1 port map( A1 => n16886, A2 => n24077, Z => n16759);
   U15107 : XOR2_X1 port map( A1 => n27921, A2 => n19515, Z => n11098);
   U15110 : XOR2_X1 port map( A1 => n11026, A2 => n206, Z => n12413);
   U15111 : NOR2_X1 port map( A1 => n2484, A2 => n12667, ZN => n28174);
   U15115 : NOR2_X1 port map( A1 => n3326, A2 => n8472, ZN => n23311);
   U15119 : NAND3_X1 port map( A1 => n2452, A2 => n2453, A3 => n25753, ZN => 
                           n28183);
   U15122 : XOR2_X1 port map( A1 => n11575, A2 => n19349, Z => n19449);
   U15129 : NOR2_X1 port map( A1 => n6889, A2 => n19155, ZN => n14395);
   U15136 : NAND3_X1 port map( A1 => n20811, A2 => n20810, A3 => n27332, ZN => 
                           n27584);
   U15138 : NAND2_X2 port map( A1 => n13515, A2 => n10823, ZN => n27836);
   U15141 : XOR2_X1 port map( A1 => n15723, A2 => n609, Z => n27585);
   U15143 : XOR2_X1 port map( A1 => n25445, A2 => n28466, Z => n27999);
   U15147 : NAND3_X2 port map( A1 => n1006, A2 => n12375, A3 => n5801, ZN => 
                           n27587);
   U15151 : XOR2_X1 port map( A1 => n2978, A2 => n18231, Z => n25227);
   U15157 : XNOR2_X1 port map( A1 => n25445, A2 => n13851, ZN => n18231);
   U15159 : XOR2_X1 port map( A1 => n27700, A2 => n25865, Z => n2978);
   U15163 : XOR2_X1 port map( A1 => n18215, A2 => n6718, Z => n18175);
   U15165 : NAND2_X2 port map( A1 => n6719, A2 => n27836, ZN => n18215);
   U15167 : NAND2_X1 port map( A1 => n6042, A2 => n24429, ZN => n18672);
   U15171 : OAI21_X2 port map( A1 => n5227, A2 => n16657, B => n16512, ZN => 
                           n10989);
   U15174 : XOR2_X1 port map( A1 => n19274, A2 => n27589, Z => n24669);
   U15181 : INV_X1 port map( I => n14590, ZN => n27589);
   U15183 : NOR2_X2 port map( A1 => n15424, A2 => n14582, ZN => n19274);
   U15189 : INV_X2 port map( I => n27590, ZN => n8102);
   U15193 : XOR2_X1 port map( A1 => n18246, A2 => n14139, Z => n27694);
   U15194 : NOR2_X2 port map( A1 => n12488, A2 => n17613, ZN => n18246);
   U15195 : NOR2_X1 port map( A1 => n15892, A2 => n15891, ZN => n6314);
   U15196 : XOR2_X1 port map( A1 => Plaintext(5), A2 => Key(5), Z => n15891);
   U15197 : XOR2_X1 port map( A1 => n11034, A2 => n28350, Z => n15030);
   U15199 : XOR2_X1 port map( A1 => n24107, A2 => n27591, Z => n17100);
   U15204 : NAND2_X1 port map( A1 => n19837, A2 => n27202, ZN => n27592);
   U15205 : OAI22_X2 port map( A1 => n13105, A2 => n12889, B1 => n12888, B2 => 
                           n18971, ZN => n19532);
   U15207 : XOR2_X1 port map( A1 => n9985, A2 => n608, Z => n3358);
   U15211 : NAND2_X2 port map( A1 => n11800, A2 => n13106, ZN => n21035);
   U15214 : NAND2_X1 port map( A1 => n14319, A2 => n4386, ZN => n27593);
   U15220 : INV_X2 port map( I => n25316, ZN => n11803);
   U15223 : NAND2_X2 port map( A1 => n1084, A2 => n13050, ZN => n25316);
   U15227 : NOR2_X1 port map( A1 => n27838, A2 => n12593, ZN => n13682);
   U15234 : XOR2_X1 port map( A1 => n15088, A2 => n21201, Z => n4834);
   U15238 : XOR2_X1 port map( A1 => n27595, A2 => n2423, Z => Ciphertext(75));
   U15239 : NOR2_X1 port map( A1 => n2425, A2 => n28424, ZN => n27595);
   U15242 : XOR2_X1 port map( A1 => n27596, A2 => n11152, Z => Ciphertext(116))
                           ;
   U15255 : OAI21_X1 port map( A1 => n21457, A2 => n21441, B => n24538, ZN => 
                           n5214);
   U15259 : INV_X4 port map( I => n27597, ZN => n12521);
   U15260 : AND2_X2 port map( A1 => n23201, A2 => n8436, Z => n27597);
   U15261 : NAND2_X2 port map( A1 => n25841, A2 => n21020, ZN => n21066);
   U15268 : AOI22_X2 port map( A1 => n27598, A2 => n17785, B1 => n9062, B2 => 
                           n22312, ZN => n18237);
   U15273 : OAI22_X2 port map( A1 => n22312, A2 => n8117, B1 => n23542, B2 => 
                           n10823, ZN => n27598);
   U15278 : NAND2_X2 port map( A1 => n10842, A2 => n10668, ZN => n18933);
   U15292 : XOR2_X1 port map( A1 => n28253, A2 => n20726, Z => n10460);
   U15294 : XOR2_X1 port map( A1 => n22806, A2 => n20543, Z => n20726);
   U15296 : NAND3_X2 port map( A1 => n27601, A2 => n8617, A3 => n27600, ZN => 
                           n14382);
   U15300 : NAND2_X1 port map( A1 => n8616, A2 => n8619, ZN => n27601);
   U15301 : XOR2_X1 port map( A1 => n26548, A2 => n18229, Z => n12484);
   U15302 : OAI22_X2 port map( A1 => n28264, A2 => n11454, B1 => n23533, B2 => 
                           n27606, ZN => n23355);
   U15303 : XOR2_X1 port map( A1 => n19509, A2 => n15053, Z => n13714);
   U15306 : XOR2_X1 port map( A1 => n14979, A2 => n26723, Z => n27764);
   U15309 : NAND2_X2 port map( A1 => n27603, A2 => n17653, ZN => n17755);
   U15319 : XOR2_X1 port map( A1 => n19488, A2 => n26728, Z => n26589);
   U15322 : XOR2_X1 port map( A1 => n12527, A2 => n19312, Z => n19488);
   U15328 : XOR2_X1 port map( A1 => n18058, A2 => n18204, Z => n24498);
   U15329 : XOR2_X1 port map( A1 => n23681, A2 => n10149, Z => n18204);
   U15330 : INV_X2 port map( I => n14929, ZN => n27606);
   U15336 : INV_X2 port map( I => n674, ZN => n27607);
   U15337 : XOR2_X1 port map( A1 => n24094, A2 => n10202, Z => n20363);
   U15338 : NAND2_X1 port map( A1 => n16517, A2 => n10543, ZN => n4983);
   U15342 : AOI22_X2 port map( A1 => n4954, A2 => n5884, B1 => n9966, B2 => 
                           n15809, ZN => n10543);
   U15345 : NOR2_X2 port map( A1 => n14649, A2 => n18782, ZN => n6558);
   U15348 : BUF_X4 port map( I => n10538, Z => n27848);
   U15353 : XOR2_X1 port map( A1 => n27609, A2 => n13497, Z => n24329);
   U15354 : XOR2_X1 port map( A1 => n24506, A2 => n13109, Z => n27609);
   U15361 : NAND2_X2 port map( A1 => n4234, A2 => n27610, ZN => n12276);
   U15365 : XOR2_X1 port map( A1 => n27611, A2 => n21902, Z => n23568);
   U15369 : XOR2_X1 port map( A1 => n18039, A2 => n28287, Z => n27611);
   U15371 : NAND2_X2 port map( A1 => n8326, A2 => n27607, ZN => n23533);
   U15373 : INV_X2 port map( I => n27612, ZN => n18694);
   U15374 : XNOR2_X1 port map( A1 => n18196, A2 => n25138, ZN => n27612);
   U15382 : XOR2_X1 port map( A1 => n9932, A2 => n9933, Z => n20367);
   U15383 : AND2_X2 port map( A1 => n8564, A2 => n26415, Z => n19683);
   U15384 : XOR2_X1 port map( A1 => n19564, A2 => n19182, Z => n7660);
   U15392 : XOR2_X1 port map( A1 => n19481, A2 => n26178, Z => n19564);
   U15408 : XOR2_X1 port map( A1 => n20399, A2 => n11811, Z => n2776);
   U15409 : XOR2_X1 port map( A1 => n21299, A2 => n15547, Z => n20399);
   U15412 : NAND2_X2 port map( A1 => n4329, A2 => n27614, ZN => n8290);
   U15413 : NAND2_X2 port map( A1 => n2251, A2 => n2252, ZN => n3574);
   U15415 : AOI22_X2 port map( A1 => n3113, A2 => n23725, B1 => n20088, B2 => 
                           n11991, ZN => n2251);
   U15417 : XOR2_X1 port map( A1 => n9674, A2 => n1496, Z => n19188);
   U15419 : INV_X1 port map( I => n6912, ZN => n27615);
   U15426 : NAND2_X2 port map( A1 => n27616, A2 => n27717, ZN => n19150);
   U15427 : NOR2_X2 port map( A1 => n19889, A2 => n19850, ZN => n3878);
   U15432 : XOR2_X1 port map( A1 => n19444, A2 => n15639, Z => n28067);
   U15433 : NAND2_X2 port map( A1 => n27617, A2 => n28123, ZN => n28469);
   U15434 : INV_X4 port map( I => n19011, ZN => n1159);
   U15436 : NAND2_X2 port map( A1 => n2132, A2 => n27628, ZN => n19011);
   U15439 : INV_X1 port map( I => n18714, ZN => n27657);
   U15440 : XOR2_X1 port map( A1 => n27936, A2 => n17109, Z => n14797);
   U15457 : XOR2_X1 port map( A1 => n27620, A2 => n5823, Z => n25985);
   U15471 : XOR2_X1 port map( A1 => n18292, A2 => n18293, Z => n27620);
   U15477 : INV_X2 port map( I => n21008, ZN => n1431);
   U15478 : NAND2_X2 port map( A1 => n9396, A2 => n27621, ZN => n13001);
   U15485 : NAND2_X2 port map( A1 => n27790, A2 => n14959, ZN => n27621);
   U15486 : XOR2_X1 port map( A1 => n10906, A2 => n2025, Z => n2026);
   U15493 : AOI22_X2 port map( A1 => n16733, A2 => n10518, B1 => n10517, B2 => 
                           n16474, ZN => n10906);
   U15500 : NAND3_X2 port map( A1 => n13005, A2 => n25662, A3 => n27622, ZN => 
                           n25559);
   U15502 : NAND3_X1 port map( A1 => n18446, A2 => n3674, A3 => n18534, ZN => 
                           n27622);
   U15507 : XOR2_X1 port map( A1 => n14294, A2 => n27661, Z => n2235);
   U15509 : NOR2_X2 port map( A1 => n15012, A2 => n15013, ZN => n27661);
   U15516 : BUF_X2 port map( I => n14754, Z => n27623);
   U15517 : NAND2_X1 port map( A1 => n8135, A2 => n8810, ZN => n19812);
   U15524 : NAND3_X1 port map( A1 => n461, A2 => n10081, A3 => n17452, ZN => 
                           n17004);
   U15528 : XOR2_X1 port map( A1 => n27625, A2 => n21597, Z => Ciphertext(157))
                           ;
   U15534 : NAND2_X2 port map( A1 => n27687, A2 => n16590, ZN => n17039);
   U15535 : OAI21_X2 port map( A1 => n17961, A2 => n5449, B => n17960, ZN => 
                           n18205);
   U15536 : XOR2_X1 port map( A1 => n21421, A2 => n20718, Z => n5724);
   U15537 : XOR2_X1 port map( A1 => n5446, A2 => n21183, Z => n21421);
   U15540 : NAND2_X2 port map( A1 => n15270, A2 => n27627, ZN => n15470);
   U15542 : OAI21_X2 port map( A1 => n5311, A2 => n1076, B => n1079, ZN => 
                           n27627);
   U15543 : XOR2_X1 port map( A1 => n26038, A2 => n4656, Z => n16545);
   U15545 : XOR2_X1 port map( A1 => n22788, A2 => n27425, Z => n11630);
   U15551 : NAND2_X2 port map( A1 => n14855, A2 => n14854, ZN => n22788);
   U15552 : NAND2_X1 port map( A1 => n2135, A2 => n2136, ZN => n27628);
   U15555 : XOR2_X1 port map( A1 => n8424, A2 => n7988, Z => n25797);
   U15558 : INV_X1 port map( I => n1995, ZN => n11225);
   U15559 : NAND2_X1 port map( A1 => n12256, A2 => n1995, ZN => n4664);
   U15563 : AOI22_X2 port map( A1 => n24806, A2 => n14866, B1 => n15490, B2 => 
                           n10142, ZN => n27629);
   U15564 : NAND2_X2 port map( A1 => n25233, A2 => n22047, ZN => n6216);
   U15566 : XOR2_X1 port map( A1 => n19555, A2 => n19558, Z => n10391);
   U15576 : NAND2_X2 port map( A1 => n2328, A2 => n2329, ZN => n18286);
   U15577 : AND3_X1 port map( A1 => n24697, A2 => n15596, A3 => n24696, Z => 
                           n27632);
   U15581 : AOI22_X2 port map( A1 => n18600, A2 => n18602, B1 => n18458, B2 => 
                           n18599, ZN => n5424);
   U15582 : NOR2_X2 port map( A1 => n13788, A2 => n5325, ZN => n15641);
   U15583 : NAND2_X2 port map( A1 => n27641, A2 => n22142, ZN => n20550);
   U15586 : NOR2_X2 port map( A1 => n22672, A2 => n20314, ZN => n26514);
   U15587 : NAND2_X2 port map( A1 => n11154, A2 => n11155, ZN => n10038);
   U15590 : OAI21_X2 port map( A1 => n23034, A2 => n23035, B => n11175, ZN => 
                           n27634);
   U15595 : NAND2_X1 port map( A1 => n26234, A2 => n23488, ZN => n3801);
   U15603 : NOR2_X2 port map( A1 => n23129, A2 => n7771, ZN => n23488);
   U15607 : NAND2_X2 port map( A1 => n27635, A2 => n24405, ZN => n9978);
   U15609 : NAND2_X1 port map( A1 => n23165, A2 => n10001, ZN => n27635);
   U15613 : NAND2_X2 port map( A1 => n22277, A2 => n27636, ZN => n16853);
   U15614 : OAI21_X2 port map( A1 => n12504, A2 => n13305, B => n912, ZN => 
                           n27636);
   U15617 : NAND2_X2 port map( A1 => n27637, A2 => n17894, ZN => n11959);
   U15619 : NAND2_X2 port map( A1 => n26643, A2 => n22253, ZN => n27637);
   U15620 : INV_X1 port map( I => n19124, ZN => n27736);
   U15623 : NAND2_X2 port map( A1 => n27795, A2 => n18567, ZN => n19124);
   U15626 : INV_X1 port map( I => n19527, ZN => n19200);
   U15634 : OAI21_X1 port map( A1 => n15243, A2 => n6767, B => n13662, ZN => 
                           n5456);
   U15640 : OR2_X1 port map( A1 => n25769, A2 => n10537, Z => n18080);
   U15645 : NOR2_X2 port map( A1 => n13872, A2 => n990, ZN => n5818);
   U15648 : OAI22_X2 port map( A1 => n27638, A2 => n4397, B1 => n5984, B2 => 
                           n19120, ZN => n8777);
   U15649 : NOR2_X2 port map( A1 => n8814, A2 => n28548, ZN => n27638);
   U15653 : NAND3_X2 port map( A1 => n25526, A2 => n15002, A3 => n25525, ZN => 
                           n19435);
   U15654 : NAND2_X2 port map( A1 => n24622, A2 => n27639, ZN => n12816);
   U15657 : OAI21_X2 port map( A1 => n16424, A2 => n16687, B => n11951, ZN => 
                           n28517);
   U15658 : NOR2_X2 port map( A1 => n26514, A2 => n24445, ZN => n27641);
   U15664 : NOR3_X2 port map( A1 => n20220, A2 => n27642, A3 => n26706, ZN => 
                           n20221);
   U15668 : OR2_X1 port map( A1 => n14726, A2 => n19846, Z => n28375);
   U15669 : XOR2_X1 port map( A1 => n507, A2 => n27644, Z => n11619);
   U15670 : XOR2_X1 port map( A1 => n8224, A2 => n7267, Z => n27644);
   U15673 : NAND2_X1 port map( A1 => n6257, A2 => n6255, ZN => n28458);
   U15674 : NOR2_X2 port map( A1 => n20090, A2 => n20288, ZN => n20431);
   U15675 : NAND2_X2 port map( A1 => n14660, A2 => n14661, ZN => n20100);
   U15676 : NAND3_X2 port map( A1 => n24645, A2 => n25061, A3 => n1906, ZN => 
                           n7832);
   U15678 : NAND2_X2 port map( A1 => n27645, A2 => n1793, ZN => n8915);
   U15679 : NOR2_X2 port map( A1 => n26690, A2 => n2481, ZN => n27645);
   U15680 : NOR2_X2 port map( A1 => n27646, A2 => n6887, ZN => n19496);
   U15681 : NAND2_X2 port map( A1 => n28505, A2 => n3220, ZN => n13834);
   U15682 : XOR2_X1 port map( A1 => n18357, A2 => n1680, Z => n1676);
   U15690 : XOR2_X1 port map( A1 => n25631, A2 => n6718, Z => n1680);
   U15702 : NAND2_X2 port map( A1 => n19468, A2 => n19949, ZN => n11973);
   U15703 : XOR2_X1 port map( A1 => n16786, A2 => n4659, Z => n16790);
   U15707 : XOR2_X1 port map( A1 => n23754, A2 => n7973, Z => n16786);
   U15712 : XOR2_X1 port map( A1 => n15546, A2 => n5937, Z => n5543);
   U15714 : INV_X2 port map( I => n10985, ZN => n27648);
   U15716 : OAI21_X2 port map( A1 => n27651, A2 => n27650, B => n27649, ZN => 
                           n853);
   U15717 : INV_X2 port map( I => n8976, ZN => n27651);
   U15735 : NAND2_X2 port map( A1 => n2208, A2 => n27652, ZN => n5231);
   U15739 : XOR2_X1 port map( A1 => n27654, A2 => n18237, Z => n18194);
   U15740 : INV_X2 port map( I => n6024, ZN => n27654);
   U15745 : XOR2_X1 port map( A1 => n27655, A2 => n13223, Z => n167);
   U15746 : OAI21_X2 port map( A1 => n24149, A2 => n9784, B => n26992, ZN => 
                           n28307);
   U15754 : NOR3_X1 port map( A1 => n18294, A2 => n1618, A3 => n25968, ZN => 
                           n27656);
   U15757 : BUF_X2 port map( I => n22085, Z => n27658);
   U15758 : XOR2_X1 port map( A1 => n22487, A2 => n27659, Z => n2914);
   U15759 : XOR2_X1 port map( A1 => n27459, A2 => n11502, Z => n27659);
   U15765 : XOR2_X1 port map( A1 => n7679, A2 => n25408, Z => n7681);
   U15766 : OAI21_X1 port map( A1 => n8897, A2 => n10797, B => n27776, ZN => 
                           n8896);
   U15773 : NOR3_X1 port map( A1 => n23488, A2 => n26234, A3 => n875, ZN => 
                           n18561);
   U15774 : NAND2_X2 port map( A1 => n24007, A2 => n24006, ZN => n27660);
   U15776 : NAND2_X2 port map( A1 => n10662, A2 => n27663, ZN => n15679);
   U15779 : OAI21_X2 port map( A1 => n3661, A2 => n14017, B => n27665, ZN => 
                           n13888);
   U15780 : AOI22_X2 port map( A1 => n5627, A2 => n849, B1 => n5626, B2 => 
                           n14281, ZN => n27665);
   U15782 : NAND2_X2 port map( A1 => n2232, A2 => n21342, ZN => n21343);
   U15784 : NAND2_X1 port map( A1 => n27666, A2 => n16283, ZN => n12510);
   U15791 : XOR2_X1 port map( A1 => n3358, A2 => n9324, Z => n7186);
   U15793 : BUF_X2 port map( I => n2706, Z => n27668);
   U15798 : XOR2_X1 port map( A1 => n28182, A2 => n11630, Z => n215);
   U15809 : XOR2_X1 port map( A1 => n19214, A2 => n22349, Z => n19493);
   U15811 : NOR2_X2 port map( A1 => n18637, A2 => n18638, ZN => n19214);
   U15817 : AND2_X1 port map( A1 => n20023, A2 => n4021, Z => n28331);
   U15823 : BUF_X2 port map( I => n17353, Z => n27670);
   U15830 : NAND3_X2 port map( A1 => n26300, A2 => n27672, A3 => n27671, ZN => 
                           n6928);
   U15832 : BUF_X2 port map( I => n14876, Z => n27673);
   U15840 : BUF_X2 port map( I => n20044, Z => n27674);
   U15847 : NAND2_X2 port map( A1 => n27675, A2 => n2745, ZN => n10175);
   U15851 : XOR2_X1 port map( A1 => n9774, A2 => n16806, Z => n4334);
   U15853 : NAND2_X2 port map( A1 => n22959, A2 => n28074, ZN => n9774);
   U15858 : XOR2_X1 port map( A1 => n19445, A2 => n4076, Z => n19276);
   U15864 : NAND2_X2 port map( A1 => n3646, A2 => n3647, ZN => n4076);
   U15866 : XOR2_X1 port map( A1 => n16894, A2 => n27676, Z => n10333);
   U15867 : XOR2_X1 port map( A1 => n27677, A2 => n17049, Z => n27676);
   U15872 : INV_X1 port map( I => n16809, ZN => n27677);
   U15873 : XOR2_X1 port map( A1 => n3834, A2 => n12674, Z => n26305);
   U15874 : NOR2_X2 port map( A1 => n24065, A2 => n24064, ZN => n3834);
   U15875 : NAND2_X2 port map( A1 => n2253, A2 => n7769, ZN => n8213);
   U15876 : XOR2_X1 port map( A1 => n16886, A2 => n17094, Z => n27861);
   U15882 : AOI22_X2 port map( A1 => n5559, A2 => n28083, B1 => n7265, B2 => 
                           n10893, ZN => n16886);
   U15884 : XOR2_X1 port map( A1 => n22760, A2 => n19512, Z => n19411);
   U15887 : NAND2_X2 port map( A1 => n18911, A2 => n14438, ZN => n19512);
   U15893 : NOR3_X2 port map( A1 => n28126, A2 => n16474, A3 => n28125, ZN => 
                           n6472);
   U15898 : NAND2_X2 port map( A1 => n10117, A2 => n10119, ZN => n17141);
   U15905 : NOR2_X1 port map( A1 => n27454, A2 => n28151, ZN => n25833);
   U15906 : NOR2_X2 port map( A1 => n9653, A2 => n12056, ZN => n22797);
   U15908 : XOR2_X1 port map( A1 => n27678, A2 => n19548, Z => n7181);
   U15909 : XOR2_X1 port map( A1 => n22423, A2 => n19287, Z => n27678);
   U15911 : BUF_X2 port map( I => n8100, Z => n27679);
   U15913 : NAND2_X1 port map( A1 => n739, A2 => n6076, ZN => n4104);
   U15916 : NAND3_X1 port map( A1 => n17508, A2 => n8165, A3 => n16846, ZN => 
                           n25392);
   U15919 : XOR2_X1 port map( A1 => n3020, A2 => n27680, Z => n3019);
   U15922 : XOR2_X1 port map( A1 => n23973, A2 => n3022, Z => n27680);
   U15924 : INV_X1 port map( I => n3645, ZN => n21983);
   U15930 : NAND2_X1 port map( A1 => n19976, A2 => n12973, ZN => n28188);
   U15932 : NAND2_X2 port map( A1 => n15679, A2 => n9115, ZN => n2352);
   U15935 : NAND3_X2 port map( A1 => n15046, A2 => n23869, A3 => n25103, ZN => 
                           n27681);
   U15936 : NAND2_X1 port map( A1 => n21689, A2 => n21730, ZN => n13398);
   U15949 : NAND2_X2 port map( A1 => n19974, A2 => n3535, ZN => n3534);
   U15951 : NAND2_X1 port map( A1 => n17354, A2 => n17355, ZN => n27682);
   U15952 : NAND2_X2 port map( A1 => n19227, A2 => n19226, ZN => n19366);
   U15954 : NAND2_X2 port map( A1 => n26722, A2 => n2178, ZN => n19227);
   U15959 : OR2_X2 port map( A1 => n22478, A2 => n24990, Z => n21140);
   U15961 : OR3_X1 port map( A1 => n20817, A2 => n23284, A3 => n6375, Z => 
                           n8198);
   U15972 : NAND2_X2 port map( A1 => n11262, A2 => n18432, ZN => n8025);
   U15986 : XOR2_X1 port map( A1 => n12036, A2 => n27683, Z => n18575);
   U15987 : XOR2_X1 port map( A1 => n17746, A2 => n18326, Z => n27683);
   U15992 : NAND2_X1 port map( A1 => n1880, A2 => n8230, ZN => n27723);
   U15994 : XOR2_X1 port map( A1 => n27684, A2 => n14573, Z => Ciphertext(15));
   U15996 : NAND2_X1 port map( A1 => n23820, A2 => n25258, ZN => n27684);
   U16001 : OAI21_X2 port map( A1 => n22921, A2 => n25833, B => n6264, ZN => 
                           n27685);
   U16004 : XOR2_X1 port map( A1 => n23917, A2 => n27944, Z => n19534);
   U16006 : OAI21_X2 port map( A1 => n25560, A2 => n25561, B => n23421, ZN => 
                           n4816);
   U16009 : XOR2_X1 port map( A1 => n10072, A2 => n14166, Z => n26083);
   U16013 : XOR2_X1 port map( A1 => n23010, A2 => n9650, Z => n10072);
   U16014 : XOR2_X1 port map( A1 => n10798, A2 => n1094, Z => n27686);
   U16015 : AOI22_X2 port map( A1 => n22201, A2 => n16584, B1 => n7115, B2 => 
                           n1697, ZN => n27687);
   U16024 : AOI22_X2 port map( A1 => n28175, A2 => n8268, B1 => n8265, B2 => 
                           n8267, ZN => n27688);
   U16025 : XOR2_X1 port map( A1 => n2224, A2 => n20012, Z => n21974);
   U16029 : NOR3_X2 port map( A1 => n8026, A2 => n10677, A3 => n18669, ZN => 
                           n19116);
   U16032 : XOR2_X1 port map( A1 => n13966, A2 => n19345, Z => n22463);
   U16038 : XOR2_X1 port map( A1 => n11054, A2 => n19445, Z => n13966);
   U16039 : XOR2_X1 port map( A1 => n13904, A2 => n13357, Z => n12480);
   U16043 : NAND2_X2 port map( A1 => n4448, A2 => n4447, ZN => n13904);
   U16045 : XOR2_X1 port map( A1 => n15801, A2 => Key(162), Z => n27877);
   U16048 : XOR2_X1 port map( A1 => n23248, A2 => n2887, Z => n27692);
   U16051 : INV_X2 port map( I => n27694, ZN => n24659);
   U16054 : NAND2_X2 port map( A1 => n22282, A2 => n22561, ZN => n19161);
   U16055 : XOR2_X1 port map( A1 => n19336, A2 => n599, Z => n13863);
   U16058 : NOR2_X1 port map( A1 => n10111, A2 => n8632, ZN => n10114);
   U16060 : XOR2_X1 port map( A1 => n8225, A2 => n27732, Z => n27695);
   U16068 : AND2_X1 port map( A1 => n14718, A2 => n8668, Z => n28509);
   U16070 : NAND2_X2 port map( A1 => n11027, A2 => n11028, ZN => n13357);
   U16071 : XOR2_X1 port map( A1 => n11811, A2 => n14227, Z => n21300);
   U16074 : NAND2_X1 port map( A1 => n2023, A2 => n2656, ZN => n27696);
   U16075 : XOR2_X1 port map( A1 => n12095, A2 => n12093, Z => n27797);
   U16076 : OAI21_X1 port map( A1 => n12836, A2 => n10858, B => n27822, ZN => 
                           n24734);
   U16077 : NAND2_X2 port map( A1 => n11138, A2 => n10658, ZN => n27822);
   U16078 : INV_X2 port map( I => n2394, ZN => n27697);
   U16081 : NAND3_X2 port map( A1 => n17703, A2 => n26714, A3 => n22962, ZN => 
                           n27759);
   U16083 : NAND2_X2 port map( A1 => n17281, A2 => n7120, ZN => n17703);
   U16087 : XOR2_X1 port map( A1 => n27698, A2 => n18123, Z => n10641);
   U16089 : NAND2_X1 port map( A1 => n17865, A2 => n17866, ZN => n27698);
   U16093 : NAND2_X1 port map( A1 => n1497, A2 => n22727, ZN => n1494);
   U16100 : NAND2_X2 port map( A1 => n23878, A2 => n8281, ZN => n22727);
   U16104 : BUF_X2 port map( I => n17470, Z => n27699);
   U16106 : OAI21_X2 port map( A1 => n24615, A2 => n2958, B => n2956, ZN => 
                           n25865);
   U16107 : OAI22_X2 port map( A1 => n1650, A2 => n7228, B1 => n20556, B2 => 
                           n1090, ZN => n1891);
   U16110 : AND2_X1 port map( A1 => n3855, A2 => n15500, Z => n12446);
   U16113 : AOI22_X2 port map( A1 => n19794, A2 => n19795, B1 => n12982, B2 => 
                           n13775, ZN => n20291);
   U16119 : INV_X1 port map( I => n17157, ZN => n27773);
   U16121 : NAND2_X2 port map( A1 => n19100, A2 => n11692, ZN => n13719);
   U16123 : NAND2_X2 port map( A1 => n12749, A2 => n25847, ZN => n19100);
   U16124 : BUF_X2 port map( I => n25592, Z => n27701);
   U16126 : OAI21_X2 port map( A1 => n8027, A2 => n3156, B => n25468, ZN => 
                           n27703);
   U16128 : NAND2_X2 port map( A1 => n8187, A2 => n17705, ZN => n18172);
   U16129 : XOR2_X1 port map( A1 => n16944, A2 => n13443, Z => n16767);
   U16132 : NOR2_X2 port map( A1 => n27706, A2 => n12755, ZN => n12754);
   U16133 : NOR2_X2 port map( A1 => n20102, A2 => n1580, ZN => n27706);
   U16134 : BUF_X4 port map( I => n12718, Z => n28233);
   U16135 : OAI21_X2 port map( A1 => n8180, A2 => n3961, B => n27707, ZN => 
                           n17253);
   U16136 : NAND2_X2 port map( A1 => n8180, A2 => n17251, ZN => n27707);
   U16137 : OAI21_X2 port map( A1 => n18800, A2 => n27701, B => n27709, ZN => 
                           n5652);
   U16139 : NOR2_X2 port map( A1 => n18991, A2 => n27704, ZN => n27709);
   U16142 : NAND2_X1 port map( A1 => n27710, A2 => n3433, ZN => n18714);
   U16147 : XOR2_X1 port map( A1 => n3331, A2 => n8450, Z => n3433);
   U16160 : NAND2_X1 port map( A1 => n6081, A2 => n6082, ZN => n27711);
   U16161 : NAND2_X2 port map( A1 => n24723, A2 => n4445, ZN => n8467);
   U16163 : XOR2_X1 port map( A1 => n23720, A2 => n6545, Z => n6968);
   U16165 : XOR2_X1 port map( A1 => n6985, A2 => n22198, Z => n7029);
   U16169 : NAND3_X2 port map( A1 => n11390, A2 => n11424, A3 => n16445, ZN => 
                           n12434);
   U16171 : NAND2_X2 port map( A1 => n13438, A2 => n24227, ZN => n11390);
   U16176 : NAND2_X2 port map( A1 => n1211, A2 => n17996, ZN => n18091);
   U16177 : AOI22_X2 port map( A1 => n22411, A2 => n24580, B1 => n12669, B2 => 
                           n2390, ZN => n8206);
   U16181 : INV_X2 port map( I => n9855, ZN => n5954);
   U16182 : NAND2_X2 port map( A1 => n27714, A2 => n18101, ZN => n9855);
   U16187 : INV_X2 port map( I => n6770, ZN => n27714);
   U16195 : AOI22_X2 port map( A1 => n6917, A2 => n14826, B1 => n6916, B2 => 
                           n4976, ZN => n27883);
   U16202 : NOR2_X2 port map( A1 => n28105, A2 => n28104, ZN => n6917);
   U16203 : XOR2_X1 port map( A1 => n28077, A2 => n19554, Z => n8654);
   U16204 : NAND2_X2 port map( A1 => n18450, A2 => n18449, ZN => n28384);
   U16207 : XOR2_X1 port map( A1 => n26559, A2 => n24530, Z => n598);
   U16208 : NAND2_X1 port map( A1 => n19955, A2 => n19828, ZN => n19473);
   U16211 : NAND3_X2 port map( A1 => n25908, A2 => n13736, A3 => n24589, ZN => 
                           n13759);
   U16214 : BUF_X4 port map( I => n4683, Z => n27734);
   U16215 : NAND3_X2 port map( A1 => n9289, A2 => n3745, A3 => n3744, ZN => 
                           n27818);
   U16221 : NAND2_X2 port map( A1 => n3697, A2 => n18556, ZN => n9289);
   U16222 : NAND2_X2 port map( A1 => n1074, A2 => n14634, ZN => n27716);
   U16236 : INV_X1 port map( I => n5231, ZN => n20088);
   U16239 : AND2_X1 port map( A1 => n27873, A2 => n5231, Z => n20232);
   U16240 : XOR2_X1 port map( A1 => n9338, A2 => n27718, Z => n10319);
   U16244 : INV_X1 port map( I => n8224, ZN => n27718);
   U16246 : AOI22_X1 port map( A1 => n27344, A2 => n8530, B1 => n23474, B2 => 
                           n8534, ZN => n1858);
   U16248 : AOI22_X2 port map( A1 => n24413, A2 => n23169, B1 => n13345, B2 => 
                           n4241, ZN => n22835);
   U16251 : NAND2_X2 port map( A1 => n12892, A2 => n865, ZN => n24413);
   U16257 : OAI22_X2 port map( A1 => n5288, A2 => n28311, B1 => n817, B2 => 
                           n27720, ZN => n7776);
   U16258 : AOI21_X1 port map( A1 => n28311, A2 => n27432, B => n19167, ZN => 
                           n27720);
   U16259 : NOR2_X2 port map( A1 => n27721, A2 => n13649, ZN => n24147);
   U16264 : NAND2_X2 port map( A1 => n11874, A2 => n11376, ZN => n18827);
   U16266 : INV_X2 port map( I => n27722, ZN => n17463);
   U16273 : XNOR2_X1 port map( A1 => n14485, A2 => n16921, ZN => n27722);
   U16274 : XOR2_X1 port map( A1 => n21386, A2 => n20458, Z => n4585);
   U16282 : NAND2_X2 port map( A1 => n27723, A2 => n28398, ZN => n23753);
   U16284 : NOR2_X2 port map( A1 => n28144, A2 => n12767, ZN => n12766);
   U16285 : NOR2_X2 port map( A1 => n22066, A2 => n27219, ZN => n27724);
   U16287 : XOR2_X1 port map( A1 => n27725, A2 => n20524, Z => n6376);
   U16291 : XOR2_X1 port map( A1 => n20565, A2 => n25023, Z => n27725);
   U16292 : INV_X4 port map( I => n12836, ZN => n20998);
   U16303 : AND2_X1 port map( A1 => n13873, A2 => n24937, Z => n26223);
   U16305 : NAND2_X1 port map( A1 => n21457, A2 => n21441, ZN => n11562);
   U16309 : XOR2_X1 port map( A1 => n25000, A2 => n27348, Z => n27726);
   U16310 : XOR2_X1 port map( A1 => n27727, A2 => n19554, Z => n606);
   U16311 : XOR2_X1 port map( A1 => n19311, A2 => n27997, Z => n27727);
   U16321 : NOR2_X2 port map( A1 => n5121, A2 => n27728, ZN => n16636);
   U16322 : AOI22_X2 port map( A1 => n24916, A2 => n4730, B1 => n9675, B2 => 
                           n17807, ZN => n24863);
   U16324 : NAND2_X2 port map( A1 => n27729, A2 => n12348, ZN => n12346);
   U16327 : BUF_X4 port map( I => n17917, Z => n24563);
   U16328 : AOI21_X2 port map( A1 => n26089, A2 => n27731, B => n28313, ZN => 
                           n2292);
   U16331 : NAND2_X1 port map( A1 => n14104, A2 => n20131, ZN => n27731);
   U16333 : XOR2_X1 port map( A1 => n481, A2 => n7951, Z => n8225);
   U16334 : OAI21_X2 port map( A1 => n14120, A2 => n14121, B => n758, ZN => 
                           n27733);
   U16336 : XOR2_X1 port map( A1 => n7422, A2 => n7424, Z => n9993);
   U16337 : XOR2_X1 port map( A1 => n12635, A2 => n26056, Z => n27735);
   U16344 : OR2_X1 port map( A1 => n822, A2 => n18683, Z => n22668);
   U16346 : XOR2_X1 port map( A1 => n7546, A2 => n7545, Z => n28135);
   U16348 : XOR2_X1 port map( A1 => n4398, A2 => n7547, Z => n7546);
   U16352 : XOR2_X1 port map( A1 => n19258, A2 => n19257, Z => n19593);
   U16354 : XOR2_X1 port map( A1 => n17840, A2 => n24318, Z => n18058);
   U16357 : XOR2_X1 port map( A1 => n27911, A2 => n15039, Z => n3462);
   U16362 : NAND2_X2 port map( A1 => n27738, A2 => n21327, ZN => n21330);
   U16365 : NAND2_X2 port map( A1 => n28209, A2 => n2661, ZN => n9314);
   U16367 : INV_X2 port map( I => n13685, ZN => n14059);
   U16384 : NAND2_X2 port map( A1 => n12459, A2 => n161, ZN => n13685);
   U16386 : XOR2_X1 port map( A1 => n16913, A2 => n16914, Z => n26579);
   U16387 : NAND2_X2 port map( A1 => n26057, A2 => n16441, ZN => n16914);
   U16393 : NOR2_X2 port map( A1 => n21500, A2 => n21495, ZN => n21465);
   U16398 : INV_X1 port map( I => n27780, ZN => n21495);
   U16399 : XOR2_X1 port map( A1 => n84, A2 => n3348, Z => n27780);
   U16401 : AOI21_X1 port map( A1 => n7841, A2 => n4780, B => n2202, ZN => 
                           n18365);
   U16403 : NAND2_X2 port map( A1 => n24847, A2 => n24846, ZN => n2202);
   U16406 : AOI21_X2 port map( A1 => n19847, A2 => n19848, B => n1116, ZN => 
                           n14661);
   U16410 : INV_X2 port map( I => n27740, ZN => n24643);
   U16412 : XNOR2_X1 port map( A1 => Plaintext(25), A2 => Key(25), ZN => n27740
                           );
   U16413 : XOR2_X1 port map( A1 => n27741, A2 => n27742, Z => n24120);
   U16415 : XOR2_X1 port map( A1 => n1859, A2 => n16931, Z => n27742);
   U16419 : NAND2_X2 port map( A1 => n10249, A2 => n12323, ZN => n19073);
   U16423 : AOI22_X2 port map( A1 => n18630, A2 => n21783, B1 => n14138, B2 => 
                           n12324, ZN => n12323);
   U16424 : NOR3_X2 port map( A1 => n24898, A2 => n27743, A3 => n5371, ZN => 
                           n16711);
   U16426 : XOR2_X1 port map( A1 => n5646, A2 => n5648, Z => n6509);
   U16428 : AOI21_X2 port map( A1 => n12020, A2 => n8864, B => n27744, ZN => 
                           n21182);
   U16449 : NOR2_X1 port map( A1 => n20473, A2 => n20226, ZN => n27744);
   U16453 : OAI21_X2 port map( A1 => n25987, A2 => n3373, B => n27746, ZN => 
                           n23129);
   U16454 : NOR2_X2 port map( A1 => n5704, A2 => n737, ZN => n27747);
   U16457 : OAI22_X2 port map( A1 => n23479, A2 => n4158, B1 => n3122, B2 => 
                           n11783, ZN => n7030);
   U16461 : XOR2_X1 port map( A1 => n21240, A2 => n20501, Z => n5648);
   U16462 : NAND2_X1 port map( A1 => n27899, A2 => n27748, ZN => n22575);
   U16465 : OR2_X1 port map( A1 => n7238, A2 => n19750, Z => n27748);
   U16471 : INV_X4 port map( I => n27749, ZN => n4192);
   U16472 : NAND2_X1 port map( A1 => n27752, A2 => n27750, ZN => n11320);
   U16473 : NAND2_X1 port map( A1 => n11321, A2 => n20842, ZN => n27752);
   U16481 : NOR2_X1 port map( A1 => n23938, A2 => n13084, ZN => n28094);
   U16483 : XOR2_X1 port map( A1 => n4789, A2 => n13904, Z => n11493);
   U16488 : XOR2_X1 port map( A1 => n9284, A2 => n9281, Z => n10550);
   U16489 : NAND2_X2 port map( A1 => n9029, A2 => n9030, ZN => n13095);
   U16494 : NAND2_X1 port map( A1 => n21793, A2 => n17463, ZN => n6332);
   U16496 : XOR2_X1 port map( A1 => n16917, A2 => n21890, Z => n14485);
   U16497 : XOR2_X1 port map( A1 => n22926, A2 => n27394, Z => n16917);
   U16498 : XOR2_X1 port map( A1 => n6309, A2 => n19272, Z => n15073);
   U16500 : OAI22_X2 port map( A1 => n18936, A2 => n444, B1 => n5711, B2 => 
                           n18934, ZN => n6309);
   U16501 : NAND2_X2 port map( A1 => n27753, A2 => n28161, ZN => n12667);
   U16503 : NAND2_X1 port map( A1 => n11142, A2 => n1005, ZN => n27753);
   U16504 : AOI22_X1 port map( A1 => n23557, A2 => n23556, B1 => n17286, B2 => 
                           n6762, ZN => n23486);
   U16506 : XOR2_X1 port map( A1 => n9597, A2 => n20513, Z => n20285);
   U16509 : XOR2_X1 port map( A1 => n20765, A2 => n20764, Z => n25474);
   U16514 : XOR2_X1 port map( A1 => n27754, A2 => n27384, Z => n26118);
   U16515 : XOR2_X1 port map( A1 => n18110, A2 => n12439, Z => n27754);
   U16516 : XOR2_X1 port map( A1 => n28517, A2 => n27854, Z => n9102);
   U16519 : AOI22_X2 port map( A1 => n12200, A2 => n1010, B1 => n12573, B2 => 
                           n23761, ZN => n23960);
   U16520 : XOR2_X1 port map( A1 => n6445, A2 => n23818, Z => n18928);
   U16521 : NAND2_X2 port map( A1 => n25161, A2 => n22237, ZN => n3279);
   U16524 : NAND2_X2 port map( A1 => n25262, A2 => n6115, ZN => n25161);
   U16529 : NAND2_X2 port map( A1 => n16452, A2 => n16451, ZN => n28363);
   U16530 : NOR2_X2 port map( A1 => n27756, A2 => n27755, ZN => n17588);
   U16536 : NAND2_X1 port map( A1 => n26110, A2 => n22646, ZN => n27755);
   U16538 : XOR2_X1 port map( A1 => n27084, A2 => n12523, Z => n16859);
   U16544 : AOI21_X2 port map( A1 => n16246, A2 => n24996, B => n9473, ZN => 
                           n12523);
   U16550 : XOR2_X1 port map( A1 => n5727, A2 => n27757, Z => n20935);
   U16551 : XOR2_X1 port map( A1 => n20726, A2 => n8024, Z => n27757);
   U16552 : NOR2_X1 port map( A1 => n19073, A2 => n25559, ZN => n10565);
   U16563 : XOR2_X1 port map( A1 => n18112, A2 => n18061, Z => n13109);
   U16566 : XOR2_X1 port map( A1 => n27758, A2 => n21303, Z => n28273);
   U16567 : XOR2_X1 port map( A1 => n15130, A2 => n21302, Z => n27758);
   U16570 : NAND2_X2 port map( A1 => n6687, A2 => n6688, ZN => n16413);
   U16574 : NAND2_X2 port map( A1 => n18712, A2 => n13375, ZN => n13873);
   U16575 : INV_X2 port map( I => n27760, ZN => n21924);
   U16581 : XOR2_X1 port map( A1 => n3705, A2 => n3702, Z => n27760);
   U16585 : INV_X2 port map( I => n27761, ZN => n24978);
   U16586 : XOR2_X1 port map( A1 => n14916, A2 => n14915, Z => n27761);
   U16590 : XOR2_X1 port map( A1 => n11862, A2 => n27762, Z => n20526);
   U16591 : XOR2_X1 port map( A1 => n20524, A2 => n20525, Z => n27762);
   U16600 : NAND3_X2 port map( A1 => n22407, A2 => n26372, A3 => n25116, ZN => 
                           n20965);
   U16601 : NAND2_X2 port map( A1 => n2995, A2 => n27670, ZN => n10414);
   U16603 : NAND2_X2 port map( A1 => n13766, A2 => n10141, ZN => n2995);
   U16608 : INV_X2 port map( I => n27764, ZN => n18535);
   U16618 : NAND2_X2 port map( A1 => n23564, A2 => n27763, ZN => n27766);
   U16619 : XOR2_X1 port map( A1 => n8374, A2 => n22804, Z => n19374);
   U16622 : NAND2_X2 port map( A1 => n22887, A2 => n1416, ZN => n22804);
   U16627 : INV_X2 port map( I => n3006, ZN => n27905);
   U16636 : XOR2_X1 port map( A1 => n22341, A2 => n3007, Z => n3006);
   U16639 : NAND2_X2 port map( A1 => n13330, A2 => n19991, ZN => n27767);
   U16642 : NOR2_X1 port map( A1 => n1004, A2 => n24870, ZN => n14923);
   U16645 : NAND3_X2 port map( A1 => n14521, A2 => n11631, A3 => n20019, ZN => 
                           n14854);
   U16647 : NAND2_X2 port map( A1 => n14926, A2 => n18390, ZN => n14502);
   U16652 : XOR2_X1 port map( A1 => n27771, A2 => n27769, Z => n28102);
   U16653 : XOR2_X1 port map( A1 => n27770, A2 => n18335, Z => n27769);
   U16654 : XOR2_X1 port map( A1 => n18338, A2 => n12548, Z => n27771);
   U16655 : OAI22_X2 port map( A1 => n27772, A2 => n3929, B1 => n17632, B2 => 
                           n17729, ZN => n25278);
   U16657 : AOI22_X2 port map( A1 => n2377, A2 => n25206, B1 => n17232, B2 => 
                           n1037, ZN => n23547);
   U16660 : NOR2_X2 port map( A1 => n6657, A2 => n6656, ZN => n13851);
   U16663 : NAND2_X1 port map( A1 => n11739, A2 => n12077, ZN => n407);
   U16664 : XOR2_X1 port map( A1 => n8319, A2 => n8318, Z => n13507);
   U16667 : XOR2_X1 port map( A1 => n9549, A2 => n20772, Z => n9548);
   U16675 : XOR2_X1 port map( A1 => n27673, A2 => n21435, Z => n20772);
   U16679 : OAI22_X2 port map( A1 => n21793, A2 => n17295, B1 => n3752, B2 => 
                           n9459, ZN => n3286);
   U16684 : OR2_X1 port map( A1 => n14392, A2 => n27773, Z => n17251);
   U16693 : INV_X2 port map( I => n27774, ZN => n28545);
   U16694 : NAND2_X2 port map( A1 => n3698, A2 => n9289, ZN => n27774);
   U16695 : NAND2_X1 port map( A1 => n5950, A2 => n27379, ZN => n27776);
   U16696 : OAI21_X2 port map( A1 => n2823, A2 => n26155, B => n27777, ZN => 
                           n2890);
   U16697 : OAI21_X2 port map( A1 => n25489, A2 => n24670, B => n2925, ZN => 
                           n27777);
   U16704 : NAND2_X2 port map( A1 => n19133, A2 => n25412, ZN => n19132);
   U16721 : AOI21_X2 port map( A1 => n25048, A2 => n23700, B => n27778, ZN => 
                           n3047);
   U16722 : NOR2_X1 port map( A1 => n23450, A2 => n20217, ZN => n10932);
   U16723 : XNOR2_X1 port map( A1 => n19188, A2 => n18951, ZN => n27789);
   U16724 : AOI22_X2 port map( A1 => n1923, A2 => n992, B1 => n26395, B2 => 
                           n1924, ZN => n1922);
   U16730 : NAND3_X2 port map( A1 => n27779, A2 => n26683, A3 => n13903, ZN => 
                           n10061);
   U16740 : XOR2_X1 port map( A1 => n640, A2 => n26003, Z => n27782);
   U16743 : NAND2_X2 port map( A1 => n27805, A2 => n27783, ZN => n13573);
   U16752 : NAND2_X2 port map( A1 => n18764, A2 => n26697, ZN => n27783);
   U16758 : BUF_X2 port map( I => n28299, Z => n27787);
   U16762 : BUF_X2 port map( I => n23214, Z => n27788);
   U16763 : OAI21_X1 port map( A1 => n13, A2 => n25559, B => n12521, ZN => 
                           n28242);
   U16764 : NAND2_X2 port map( A1 => n2405, A2 => n2406, ZN => n16215);
   U16768 : XOR2_X1 port map( A1 => n8150, A2 => n25633, Z => n4157);
   U16772 : XOR2_X1 port map( A1 => n12674, A2 => n2437, Z => n8150);
   U16773 : NOR2_X2 port map( A1 => n24653, A2 => n25212, ZN => n18040);
   U16774 : NOR2_X2 port map( A1 => n15650, A2 => n15649, ZN => n10773);
   U16777 : XOR2_X1 port map( A1 => n3107, A2 => n27791, Z => n25616);
   U16783 : XOR2_X1 port map( A1 => n13808, A2 => n6523, Z => n27791);
   U16786 : XOR2_X1 port map( A1 => n9670, A2 => n2986, Z => n2279);
   U16788 : XOR2_X1 port map( A1 => n6773, A2 => n27792, Z => n19734);
   U16790 : XOR2_X1 port map( A1 => n21433, A2 => n27793, Z => n23565);
   U16794 : XOR2_X1 port map( A1 => n13361, A2 => n7848, Z => n27793);
   U16795 : NAND2_X2 port map( A1 => n25951, A2 => n2121, ZN => n2185);
   U16798 : XOR2_X1 port map( A1 => n27794, A2 => n21613, Z => Ciphertext(161))
                           ;
   U16805 : OAI22_X1 port map( A1 => n21611, A2 => n21612, B1 => n21610, B2 => 
                           n24044, ZN => n27794);
   U16807 : NAND2_X1 port map( A1 => n1191, A2 => n13564, ZN => n4959);
   U16812 : INV_X2 port map( I => n27796, ZN => n19949);
   U16816 : OAI21_X2 port map( A1 => n27800, A2 => n27799, B => n8738, ZN => 
                           n13949);
   U16818 : INV_X2 port map( I => n8740, ZN => n27799);
   U16820 : INV_X2 port map( I => n4397, ZN => n27800);
   U16830 : AOI21_X2 port map( A1 => n6788, A2 => n1084, B => n27801, ZN => 
                           n6786);
   U16833 : NOR3_X2 port map( A1 => n1084, A2 => n27594, A3 => n13050, ZN => 
                           n27801);
   U16836 : XOR2_X1 port map( A1 => n27803, A2 => n4293, Z => n15234);
   U16840 : XOR2_X1 port map( A1 => n26192, A2 => n21926, Z => n27803);
   U16841 : XOR2_X1 port map( A1 => n21424, A2 => n103, Z => n24886);
   U16848 : NAND2_X2 port map( A1 => n11750, A2 => n11748, ZN => n21424);
   U16849 : AOI21_X2 port map( A1 => n17785, A2 => n10823, B => n27806, ZN => 
                           n10211);
   U16851 : NAND2_X2 port map( A1 => n9430, A2 => n11958, ZN => n1397);
   U16854 : AND2_X1 port map( A1 => n13473, A2 => n25342, Z => n10663);
   U16864 : NAND3_X2 port map( A1 => n13755, A2 => n14845, A3 => n19620, ZN => 
                           n13754);
   U16866 : NAND2_X2 port map( A1 => n19621, A2 => n25230, ZN => n13755);
   U16873 : NAND2_X2 port map( A1 => n20571, A2 => n20573, ZN => n22234);
   U16874 : NAND3_X2 port map( A1 => n4760, A2 => n13709, A3 => n10672, ZN => 
                           n2346);
   U16875 : NAND2_X2 port map( A1 => n21825, A2 => n13963, ZN => n13709);
   U16882 : INV_X2 port map( I => n11522, ZN => n23274);
   U16886 : XOR2_X1 port map( A1 => n27807, A2 => n14623, Z => Ciphertext(34));
   U16891 : AOI21_X2 port map( A1 => n17755, A2 => n13615, B => n17785, ZN => 
                           n27808);
   U16899 : XOR2_X1 port map( A1 => n27809, A2 => n20765, Z => n248);
   U16907 : XOR2_X1 port map( A1 => n8579, A2 => n13599, Z => n27809);
   U16908 : AOI22_X2 port map( A1 => n13663, A2 => n27810, B1 => n18904, B2 => 
                           n28412, ZN => n14608);
   U16909 : OAI22_X2 port map( A1 => n20971, A2 => n20973, B1 => n15450, B2 => 
                           n21097, ZN => n12836);
   U16919 : NAND2_X2 port map( A1 => n23512, A2 => n23334, ZN => n20804);
   U16921 : OAI21_X2 port map( A1 => n11303, A2 => n19574, B => n23159, ZN => 
                           n22735);
   U16923 : NOR2_X2 port map( A1 => n10847, A2 => n8831, ZN => n27812);
   U16928 : BUF_X2 port map( I => n19189, Z => n27813);
   U16938 : XOR2_X1 port map( A1 => n27814, A2 => n21090, Z => Ciphertext(89));
   U16939 : OAI22_X1 port map( A1 => n1339, A2 => n21081, B1 => n25953, B2 => 
                           n25952, ZN => n27814);
   U16940 : OAI21_X2 port map( A1 => n20219, A2 => n20138, B => n27815, ZN => 
                           n13694);
   U16941 : BUF_X4 port map( I => n7168, Z => n28481);
   U16943 : BUF_X2 port map( I => n18027, Z => n27816);
   U16946 : XNOR2_X1 port map( A1 => n19142, A2 => n21988, ZN => n28217);
   U16947 : XOR2_X1 port map( A1 => n5082, A2 => n21341, Z => n24623);
   U16951 : XOR2_X1 port map( A1 => n21433, A2 => n21431, Z => n28150);
   U16959 : INV_X2 port map( I => n7563, ZN => n21431);
   U16960 : AOI21_X1 port map( A1 => n23706, A2 => n885, B => n11967, ZN => 
                           n4608);
   U16969 : NAND2_X2 port map( A1 => n13380, A2 => n17452, ZN => n8538);
   U16981 : NAND2_X2 port map( A1 => n27818, A2 => n3742, ZN => n3960);
   U16982 : NAND2_X2 port map( A1 => n22691, A2 => n28007, ZN => n21529);
   U16987 : XOR2_X1 port map( A1 => n17031, A2 => n16992, Z => n5819);
   U16988 : XOR2_X1 port map( A1 => n10107, A2 => n18359, Z => n22487);
   U16993 : OAI22_X2 port map( A1 => n9165, A2 => n23087, B1 => n6877, B2 => 
                           n10587, ZN => n10107);
   U16994 : NAND2_X2 port map( A1 => n27819, A2 => n27991, ZN => n25412);
   U17002 : NAND2_X1 port map( A1 => n4300, A2 => n18756, ZN => n27819);
   U17009 : NAND3_X2 port map( A1 => n24790, A2 => n21504, A3 => n25424, ZN => 
                           n21534);
   U17013 : XOR2_X1 port map( A1 => n7896, A2 => n10299, Z => n5688);
   U17015 : XOR2_X1 port map( A1 => n15226, A2 => n4383, Z => n10299);
   U17017 : NOR2_X2 port map( A1 => n28252, A2 => n27458, ZN => n116);
   U17019 : OAI22_X2 port map( A1 => n7503, A2 => n7502, B1 => n23161, B2 => 
                           n27821, ZN => n12209);
   U17020 : NAND2_X1 port map( A1 => n14843, A2 => n10269, ZN => n12560);
   U17022 : NOR2_X2 port map( A1 => n27824, A2 => n15603, ZN => n26004);
   U17023 : XOR2_X1 port map( A1 => n3862, A2 => n3864, Z => n14495);
   U17026 : AOI21_X2 port map( A1 => n17238, A2 => n886, B => n27825, ZN => 
                           n6675);
   U17029 : NOR2_X2 port map( A1 => n14920, A2 => n14921, ZN => n19236);
   U17033 : INV_X2 port map( I => n20852, ZN => n28198);
   U17037 : INV_X2 port map( I => n27826, ZN => n17343);
   U17038 : XOR2_X1 port map( A1 => n3636, A2 => n3639, Z => n27826);
   U17039 : NAND3_X1 port map( A1 => n24419, A2 => n2527, A3 => n11581, ZN => 
                           n22380);
   U17040 : NOR2_X2 port map( A1 => n16349, A2 => n11330, ZN => n3088);
   U17042 : INV_X2 port map( I => n16347, ZN => n11330);
   U17043 : NOR2_X2 port map( A1 => n27123, A2 => n574, ZN => n16347);
   U17046 : XOR2_X1 port map( A1 => n27827, A2 => n11524, Z => n4744);
   U17050 : XOR2_X1 port map( A1 => n1593, A2 => n24033, Z => n27827);
   U17054 : NOR2_X2 port map( A1 => n27828, A2 => n28434, ZN => n28293);
   U17055 : INV_X2 port map( I => n27831, ZN => n14097);
   U17067 : NAND3_X1 port map( A1 => n3787, A2 => n3786, A3 => n12236, ZN => 
                           n3783);
   U17071 : XOR2_X1 port map( A1 => n13119, A2 => n18243, Z => n18326);
   U17075 : NAND2_X2 port map( A1 => n14705, A2 => n17741, ZN => n18243);
   U17078 : OAI21_X2 port map( A1 => n8180, A2 => n3741, B => n17251, ZN => 
                           n25869);
   U17080 : NOR2_X1 port map( A1 => n22303, A2 => n8898, ZN => n22302);
   U17082 : XOR2_X1 port map( A1 => n17125, A2 => n16951, Z => n17031);
   U17091 : NAND2_X2 port map( A1 => n12686, A2 => n14761, ZN => n16951);
   U17095 : AOI21_X2 port map( A1 => n24334, A2 => n27381, B => n13211, ZN => 
                           n415);
   U17100 : NAND2_X2 port map( A1 => n28411, A2 => n27832, ZN => n6766);
   U17103 : XOR2_X1 port map( A1 => n883, A2 => n17754, Z => n4777);
   U17105 : NOR2_X1 port map( A1 => n18694, A2 => n9248, ZN => n18201);
   U17106 : NOR2_X2 port map( A1 => n27833, A2 => n25496, ZN => n18099);
   U17108 : AOI21_X2 port map( A1 => n17640, A2 => n14446, B => n25929, ZN => 
                           n27833);
   U17109 : OAI21_X2 port map( A1 => n4819, A2 => n17249, B => n27834, ZN => 
                           n4814);
   U17112 : AOI22_X2 port map( A1 => n26153, A2 => n10577, B1 => n17370, B2 => 
                           n17248, ZN => n27834);
   U17115 : INV_X1 port map( I => n11854, ZN => n27835);
   U17119 : NAND2_X2 port map( A1 => n2215, A2 => n11856, ZN => n11854);
   U17129 : XOR2_X1 port map( A1 => n20422, A2 => n10986, Z => n7653);
   U17131 : XOR2_X1 port map( A1 => n12320, A2 => n9789, Z => n10986);
   U17134 : NOR2_X2 port map( A1 => n18813, A2 => n18814, ZN => n8646);
   U17138 : XOR2_X1 port map( A1 => n16957, A2 => n17077, Z => n16627);
   U17139 : AOI21_X2 port map( A1 => n22197, A2 => n14180, B => n17935, ZN => 
                           n7602);
   U17140 : NOR2_X2 port map( A1 => n3981, A2 => n2976, ZN => n27837);
   U17143 : INV_X4 port map( I => n4192, ZN => n4976);
   U17148 : OAI22_X2 port map( A1 => n34, A2 => n10593, B1 => n12145, B2 => 
                           n12863, ZN => n19920);
   U17150 : NAND2_X2 port map( A1 => n15334, A2 => n1114, ZN => n20245);
   U17151 : XOR2_X1 port map( A1 => n6572, A2 => n5610, Z => n6575);
   U17161 : XOR2_X1 port map( A1 => n17047, A2 => n6573, Z => n6572);
   U17165 : XOR2_X1 port map( A1 => n12361, A2 => n26662, Z => n7320);
   U17169 : XOR2_X1 port map( A1 => n9727, A2 => n18088, Z => n12361);
   U17175 : NOR2_X1 port map( A1 => n13278, A2 => n7793, ZN => n27839);
   U17176 : NOR2_X2 port map( A1 => n26044, A2 => n25567, ZN => n27840);
   U17179 : NAND2_X1 port map( A1 => n15860, A2 => n16292, ZN => n27841);
   U17183 : OAI21_X2 port map( A1 => n28001, A2 => n5400, B => n27842, ZN => 
                           n9731);
   U17184 : NAND3_X2 port map( A1 => n28285, A2 => n7767, A3 => n9701, ZN => 
                           n27842);
   U17203 : NAND2_X2 port map( A1 => n2523, A2 => n27843, ZN => n2591);
   U17204 : AOI21_X1 port map( A1 => n914, A2 => n24643, B => n7226, ZN => 
                           n27843);
   U17205 : NOR2_X2 port map( A1 => n26271, A2 => n19731, ZN => n27844);
   U17206 : XOR2_X1 port map( A1 => n20763, A2 => n5537, Z => n11643);
   U17207 : OAI22_X2 port map( A1 => n10901, A2 => n9103, B1 => n20032, B2 => 
                           n806, ZN => n20763);
   U17211 : NAND2_X1 port map( A1 => n28112, A2 => n14070, ZN => n8283);
   U17212 : XOR2_X1 port map( A1 => n27847, A2 => n18257, Z => n13895);
   U17213 : INV_X2 port map( I => n12146, ZN => n27847);
   U17215 : XOR2_X1 port map( A1 => n3834, A2 => n13840, Z => n18257);
   U17219 : INV_X2 port map( I => n27849, ZN => n7561);
   U17221 : XNOR2_X1 port map( A1 => n7559, A2 => n7560, ZN => n27849);
   U17228 : NOR2_X2 port map( A1 => n10865, A2 => n27850, ZN => n3486);
   U17232 : NOR3_X2 port map( A1 => n1271, A2 => n12272, A3 => n14519, ZN => 
                           n27850);
   U17233 : XOR2_X1 port map( A1 => n22050, A2 => n26216, Z => n3810);
   U17235 : NAND2_X2 port map( A1 => n1763, A2 => n16153, ZN => n26216);
   U17238 : XOR2_X1 port map( A1 => n27851, A2 => n14518, Z => Ciphertext(51));
   U17240 : BUF_X2 port map( I => n23011, Z => n27852);
   U17244 : INV_X1 port map( I => n11869, ZN => n27853);
   U17245 : NAND2_X2 port map( A1 => n26004, A2 => n13554, ZN => n11869);
   U17259 : XOR2_X1 port map( A1 => n15226, A2 => n28405, Z => n9655);
   U17260 : OAI21_X2 port map( A1 => n11812, A2 => n10951, B => n10611, ZN => 
                           n10980);
   U17267 : NOR2_X2 port map( A1 => n19689, A2 => n3563, ZN => n10951);
   U17268 : NAND2_X2 port map( A1 => n6604, A2 => n13185, ZN => n28371);
   U17273 : NAND2_X1 port map( A1 => n24323, A2 => n16935, ZN => n26227);
   U17287 : XOR2_X1 port map( A1 => n20543, A2 => n7065, Z => n21260);
   U17289 : NAND2_X2 port map( A1 => n26637, A2 => n857, ZN => n28063);
   U17290 : NOR3_X2 port map( A1 => n3473, A2 => n266, A3 => n5880, ZN => n5877
                           );
   U17308 : XOR2_X1 port map( A1 => n27855, A2 => n21358, Z => Ciphertext(125))
                           ;
   U17312 : AOI22_X1 port map( A1 => n21354, A2 => n2232, B1 => n21356, B2 => 
                           n2448, ZN => n27855);
   U17316 : NOR2_X1 port map( A1 => n8876, A2 => n8875, ZN => n5462);
   U17317 : XOR2_X1 port map( A1 => n27857, A2 => n13982, Z => n25531);
   U17322 : XOR2_X1 port map( A1 => n15329, A2 => n19274, Z => n27857);
   U17325 : NOR2_X1 port map( A1 => n4131, A2 => n18580, ZN => n10660);
   U17331 : INV_X2 port map( I => n16413, ZN => n2857);
   U17333 : AND2_X1 port map( A1 => n24764, A2 => n27859, Z => n3724);
   U17334 : XOR2_X1 port map( A1 => n27860, A2 => n7664, Z => n8724);
   U17346 : XOR2_X1 port map( A1 => n617, A2 => n24148, Z => n27860);
   U17359 : INV_X2 port map( I => n27861, ZN => n24582);
   U17362 : XOR2_X1 port map( A1 => n19518, A2 => n19325, Z => n2881);
   U17363 : OAI21_X2 port map( A1 => n1874, A2 => n467, B => n27928, ZN => 
                           n11874);
   U17364 : XOR2_X1 port map( A1 => n27864, A2 => n21256, Z => n13702);
   U17365 : XOR2_X1 port map( A1 => n28502, A2 => n21258, Z => n27864);
   U17367 : NAND2_X1 port map( A1 => n21467, A2 => n7940, ZN => n6082);
   U17368 : NOR3_X1 port map( A1 => n11147, A2 => n6323, A3 => n27405, ZN => 
                           n21871);
   U17373 : INV_X2 port map( I => n20799, ZN => n11147);
   U17374 : NAND2_X2 port map( A1 => n5302, A2 => n9031, ZN => n20799);
   U17382 : NAND3_X2 port map( A1 => n13726, A2 => n11161, A3 => n15448, ZN => 
                           n27865);
   U17384 : AOI22_X2 port map( A1 => n9402, A2 => n21026, B1 => n20541, B2 => 
                           n12160, ZN => n21004);
   U17386 : OAI22_X2 port map( A1 => n4742, A2 => n1082, B1 => n8050, B2 => 
                           n21024, ZN => n9402);
   U17390 : BUF_X2 port map( I => n23538, Z => n27867);
   U17392 : NAND2_X1 port map( A1 => n18920, A2 => n27869, ZN => n12807);
   U17395 : NOR2_X1 port map( A1 => n27870, A2 => n26641, ZN => n27869);
   U17396 : NAND2_X1 port map( A1 => n24032, A2 => n27871, ZN => n22621);
   U17398 : XOR2_X1 port map( A1 => n3463, A2 => n13810, Z => n24032);
   U17408 : NOR2_X1 port map( A1 => n10797, A2 => n27403, ZN => n2802);
   U17413 : OAI21_X2 port map( A1 => n27872, A2 => n21686, B => n21685, ZN => 
                           n6150);
   U17420 : NOR2_X2 port map( A1 => n2778, A2 => n933, ZN => n27872);
   U17429 : NAND2_X2 port map( A1 => n3578, A2 => n359, ZN => n27873);
   U17431 : AOI22_X2 port map( A1 => n2045, A2 => n16571, B1 => n6373, B2 => 
                           n12039, ZN => n28039);
   U17441 : XOR2_X1 port map( A1 => n10122, A2 => n27874, Z => n1890);
   U17461 : XOR2_X1 port map( A1 => n17026, A2 => n17025, Z => n27874);
   U17464 : INV_X2 port map( I => n27875, ZN => n5986);
   U17467 : XOR2_X1 port map( A1 => n5989, A2 => n5987, Z => n27875);
   U17472 : NAND4_X1 port map( A1 => n12493, A2 => n14926, A3 => n18388, A4 => 
                           n18390, ZN => n18392);
   U17474 : OR2_X1 port map( A1 => n8135, A2 => n8810, Z => n14602);
   U17476 : NAND2_X1 port map( A1 => n13829, A2 => n13830, ZN => n27876);
   U17478 : NAND2_X2 port map( A1 => n14641, A2 => n25879, ZN => n12933);
   U17480 : XOR2_X1 port map( A1 => n18519, A2 => n18518, Z => n18520);
   U17482 : XOR2_X1 port map( A1 => n9414, A2 => n4793, Z => n7423);
   U17485 : OAI22_X2 port map( A1 => n26262, A2 => n8722, B1 => n8512, B2 => 
                           n7964, ZN => n7963);
   U17488 : NAND2_X2 port map( A1 => n1877, A2 => n2627, ZN => n7964);
   U17489 : NOR2_X1 port map( A1 => n22817, A2 => n17687, ZN => n13620);
   U17492 : NAND2_X2 port map( A1 => n26476, A2 => n26197, ZN => n17687);
   U17493 : NAND2_X2 port map( A1 => n10959, A2 => n1996, ZN => n7390);
   U17494 : XOR2_X1 port map( A1 => n27954, A2 => n8308, Z => n616);
   U17497 : XOR2_X1 port map( A1 => n8372, A2 => n9463, Z => n8371);
   U17498 : AND2_X1 port map( A1 => n13387, A2 => n27428, Z => n9190);
   U17507 : AOI21_X2 port map( A1 => n27879, A2 => n18504, B => n26072, ZN => 
                           n23561);
   U17512 : AOI21_X2 port map( A1 => n166, A2 => n14128, B => n6031, ZN => 
                           n27879);
   U17513 : AOI21_X2 port map( A1 => n18648, A2 => n27457, B => n27880, ZN => 
                           n13263);
   U17514 : NOR2_X2 port map( A1 => n3106, A2 => n10904, ZN => n18648);
   U17515 : NOR2_X2 port map( A1 => n27882, A2 => n12007, ZN => n12003);
   U17522 : OAI21_X2 port map( A1 => n24766, A2 => n23692, B => n27883, ZN => 
                           n17840);
   U17526 : AND2_X1 port map( A1 => n19827, A2 => n19684, Z => n19612);
   U17535 : XOR2_X1 port map( A1 => n2129, A2 => n2126, Z => n7965);
   U17537 : XOR2_X1 port map( A1 => n27884, A2 => n14526, Z => Ciphertext(171))
                           ;
   U17538 : NAND2_X2 port map( A1 => n21793, A2 => n6294, ZN => n10897);
   U17547 : NOR2_X2 port map( A1 => n100, A2 => n18101, ZN => n28069);
   U17548 : XOR2_X1 port map( A1 => n14372, A2 => n21315, Z => n10966);
   U17554 : XOR2_X1 port map( A1 => n20770, A2 => n12099, Z => n21315);
   U17557 : NAND3_X2 port map( A1 => n27888, A2 => n14648, A3 => n27887, ZN => 
                           n12376);
   U17559 : INV_X2 port map( I => n24092, ZN => n27888);
   U17564 : NOR2_X2 port map( A1 => n3046, A2 => n13352, ZN => n22803);
   U17567 : OAI22_X2 port map( A1 => n4244, A2 => n20920, B1 => n22785, B2 => 
                           n26660, ZN => n3046);
   U17568 : NAND2_X2 port map( A1 => n12003, A2 => n12009, ZN => n12382);
   U17570 : OAI21_X2 port map( A1 => n447, A2 => n6725, B => n19033, ZN => 
                           n2733);
   U17574 : XOR2_X1 port map( A1 => n18118, A2 => n27890, Z => n26348);
   U17577 : XOR2_X1 port map( A1 => n27904, A2 => n27891, Z => n27890);
   U17579 : XOR2_X1 port map( A1 => n16959, A2 => n17035, Z => n16977);
   U17580 : AOI21_X2 port map( A1 => n16716, A2 => n14055, B => n26050, ZN => 
                           n16959);
   U17589 : XOR2_X1 port map( A1 => n24264, A2 => n2858, Z => n28353);
   U17595 : XOR2_X1 port map( A1 => n27892, A2 => n1303, Z => Ciphertext(186));
   U17598 : NOR3_X1 port map( A1 => n272, A2 => n693, A3 => n3442, ZN => n23211
                           );
   U17600 : XOR2_X1 port map( A1 => n5026, A2 => n4174, Z => n356);
   U17601 : XOR2_X1 port map( A1 => n13855, A2 => n12246, Z => n5026);
   U17604 : NOR2_X2 port map( A1 => n3170, A2 => n6836, ZN => n22349);
   U17613 : NAND2_X2 port map( A1 => n23029, A2 => n5424, ZN => n28019);
   U17624 : XOR2_X1 port map( A1 => n18136, A2 => n18279, Z => n13748);
   U17630 : XOR2_X1 port map( A1 => n12276, A2 => n14203, Z => n18279);
   U17635 : INV_X2 port map( I => n27893, ZN => n24674);
   U17645 : NOR2_X2 port map( A1 => n13824, A2 => n8192, ZN => n27893);
   U17650 : XOR2_X1 port map( A1 => n26884, A2 => n20481, Z => n15308);
   U17653 : XOR2_X1 port map( A1 => n14653, A2 => n20553, Z => n20482);
   U17656 : INV_X2 port map( I => n26717, ZN => n8260);
   U17658 : XOR2_X1 port map( A1 => n17038, A2 => n10538, Z => n16985);
   U17661 : NOR2_X2 port map( A1 => n7755, A2 => n9483, ZN => n10538);
   U17665 : XOR2_X1 port map( A1 => n13524, A2 => n13916, Z => n17067);
   U17666 : NAND2_X1 port map( A1 => n12026, A2 => n12434, ZN => n13897);
   U17670 : AOI21_X2 port map( A1 => n18906, A2 => n9073, B => n23672, ZN => 
                           n26330);
   U17676 : NAND2_X2 port map( A1 => n25592, A2 => n27704, ZN => n9073);
   U17677 : XOR2_X1 port map( A1 => n4656, A2 => n28293, Z => n4707);
   U17682 : NAND2_X2 port map( A1 => n24781, A2 => n25793, ZN => n4656);
   U17684 : NOR2_X2 port map( A1 => n14263, A2 => n14407, ZN => n4549);
   U17685 : INV_X2 port map( I => n3466, ZN => n24576);
   U17688 : XOR2_X1 port map( A1 => n27897, A2 => n21141, Z => Ciphertext(69));
   U17691 : NAND3_X1 port map( A1 => n20993, A2 => n20994, A3 => n20995, ZN => 
                           n27897);
   U17694 : XOR2_X1 port map( A1 => n16932, A2 => n27898, Z => n4302);
   U17697 : XOR2_X1 port map( A1 => n11193, A2 => n16957, Z => n27898);
   U17703 : OAI21_X2 port map( A1 => n10232, A2 => n26666, B => n24387, ZN => 
                           n10231);
   U17710 : NAND2_X2 port map( A1 => n21024, A2 => n21027, ZN => n8059);
   U17711 : NAND2_X2 port map( A1 => n12711, A2 => n13969, ZN => n28251);
   U17731 : INV_X2 port map( I => n2391, ZN => n22453);
   U17733 : INV_X4 port map( I => n27704, ZN => n781);
   U17735 : NAND3_X1 port map( A1 => n14424, A2 => n14594, A3 => n27453, ZN => 
                           n28112);
   U17736 : XOR2_X1 port map( A1 => n8789, A2 => n3474, Z => n10564);
   U17738 : AOI22_X2 port map( A1 => n27492, A2 => n19161, B1 => n8611, B2 => 
                           n18894, ZN => n26503);
   U17741 : OR2_X1 port map( A1 => n4386, A2 => n27428, Z => n22995);
   U17743 : XOR2_X1 port map( A1 => n4262, A2 => n12108, Z => n4386);
   U17747 : NOR2_X1 port map( A1 => n9718, A2 => n10041, ZN => n27899);
   U17752 : NAND3_X2 port map( A1 => n19246, A2 => n27900, A3 => n19247, ZN => 
                           n8810);
   U17756 : NAND3_X1 port map( A1 => n19243, A2 => n19244, A3 => n10041, ZN => 
                           n27900);
   U17760 : OAI21_X2 port map( A1 => n12670, A2 => n725, B => n17701, ZN => 
                           n17266);
   U17761 : NOR2_X2 port map( A1 => n14509, A2 => n10577, ZN => n4472);
   U17762 : INV_X2 port map( I => n7371, ZN => n10577);
   U17764 : XOR2_X1 port map( A1 => n9539, A2 => n9541, Z => n7371);
   U17768 : INV_X4 port map( I => n2549, ZN => n6910);
   U17773 : NAND2_X2 port map( A1 => n28276, A2 => n3976, ZN => n2549);
   U17774 : NOR2_X2 port map( A1 => n27902, A2 => n5381, ZN => n23669);
   U17777 : XOR2_X1 port map( A1 => n27903, A2 => n11975, Z => Ciphertext(50));
   U17781 : AOI21_X1 port map( A1 => n22753, A2 => n20878, B => n20879, ZN => 
                           n7839);
   U17786 : BUF_X2 port map( I => n18286, Z => n27904);
   U17787 : XOR2_X1 port map( A1 => n19350, A2 => n22770, Z => n23539);
   U17790 : NOR2_X2 port map( A1 => n27907, A2 => n27906, ZN => n22770);
   U17792 : AOI22_X2 port map( A1 => n27908, A2 => n19568, B1 => n27064, B2 => 
                           n4480, ZN => n10007);
   U17793 : OAI22_X2 port map( A1 => n15027, A2 => n7129, B1 => n4364, B2 => 
                           n15028, ZN => n27908);
   U17796 : NOR2_X2 port map( A1 => n26653, A2 => n9701, ZN => n6232);
   U17800 : INV_X2 port map( I => n20435, ZN => n25564);
   U17808 : OAI22_X2 port map( A1 => n7635, A2 => n3290, B1 => n7634, B2 => 
                           n11519, ZN => n20435);
   U17809 : XOR2_X1 port map( A1 => n18301, A2 => n27909, Z => n28498);
   U17811 : XOR2_X1 port map( A1 => n2704, A2 => n14622, Z => n27909);
   U17814 : NAND2_X1 port map( A1 => n27910, A2 => n22800, ZN => n26560);
   U17821 : OAI21_X1 port map( A1 => n21702, A2 => n13432, B => n8668, ZN => 
                           n27910);
   U17822 : OAI22_X2 port map( A1 => n5556, A2 => n5557, B1 => n15186, B2 => 
                           n16600, ZN => n21949);
   U17824 : NAND2_X2 port map( A1 => n5861, A2 => n26814, ZN => n16600);
   U17830 : INV_X1 port map( I => n20703, ZN => n20693);
   U17831 : NAND3_X2 port map( A1 => n26303, A2 => n20463, A3 => n20464, ZN => 
                           n20703);
   U17832 : NAND2_X2 port map( A1 => n3700, A2 => n16973, ZN => n17733);
   U17839 : NAND2_X2 port map( A1 => n17563, A2 => n17335, ZN => n3700);
   U17840 : XOR2_X1 port map( A1 => n18211, A2 => n4970, Z => n18109);
   U17842 : NAND3_X2 port map( A1 => n6208, A2 => n6207, A3 => n6206, ZN => 
                           n18211);
   U17843 : XOR2_X1 port map( A1 => n20517, A2 => n20454, Z => n27911);
   U17846 : NOR2_X1 port map( A1 => n11110, A2 => n7025, ZN => n13213);
   U17853 : INV_X1 port map( I => n12186, ZN => n12045);
   U17855 : NOR2_X2 port map( A1 => n22993, A2 => n26677, ZN => n25126);
   U17859 : NOR2_X2 port map( A1 => n28048, A2 => n27912, ZN => n11087);
   U17862 : NOR2_X2 port map( A1 => n18512, A2 => n13341, ZN => n27912);
   U17871 : AND2_X1 port map( A1 => n9606, A2 => n17751, Z => n12518);
   U17880 : NAND2_X2 port map( A1 => n9607, A2 => n9608, ZN => n9606);
   U17887 : NAND2_X2 port map( A1 => n18696, A2 => n1185, ZN => n22329);
   U17893 : XOR2_X1 port map( A1 => n7103, A2 => n13119, Z => n11644);
   U17896 : INV_X1 port map( I => n7423, ZN => n27996);
   U17897 : NAND3_X1 port map( A1 => n27913, A2 => n26527, A3 => n8330, ZN => 
                           n19854);
   U17904 : NAND3_X1 port map( A1 => n3070, A2 => n27915, A3 => n27914, ZN => 
                           n3067);
   U17906 : INV_X1 port map( I => n22453, ZN => n27914);
   U17907 : NAND2_X2 port map( A1 => n16511, A2 => n8181, ZN => n27915);
   U17913 : NAND2_X2 port map( A1 => n23046, A2 => n3657, ZN => n7134);
   U17914 : NAND2_X2 port map( A1 => n6233, A2 => n6234, ZN => n23046);
   U17918 : AND2_X1 port map( A1 => n21571, A2 => n21572, Z => n26585);
   U17924 : INV_X1 port map( I => n19136, ZN => n27918);
   U17929 : OAI22_X2 port map( A1 => n4491, A2 => n26009, B1 => n20215, B2 => 
                           n26365, ZN => n20157);
   U17935 : NAND2_X2 port map( A1 => n28091, A2 => n10221, ZN => n20215);
   U17938 : INV_X4 port map( I => n9606, ZN => n12611);
   U17939 : XOR2_X1 port map( A1 => n13299, A2 => n19302, Z => n27921);
   U17944 : XOR2_X1 port map( A1 => n27922, A2 => n11105, Z => n21101);
   U17949 : AND2_X1 port map( A1 => n7033, A2 => n5639, Z => n27974);
   U17953 : XNOR2_X1 port map( A1 => n12932, A2 => n14670, ZN => n28089);
   U17955 : NAND2_X2 port map( A1 => n25666, A2 => n27925, ZN => n18041);
   U17961 : BUF_X2 port map( I => n15282, Z => n27926);
   U17963 : AOI21_X2 port map( A1 => n13845, A2 => n27512, B => n1891, ZN => 
                           n21008);
   U17965 : INV_X2 port map( I => n3223, ZN => n7908);
   U17971 : NAND2_X2 port map( A1 => n8152, A2 => n24245, ZN => n3223);
   U17972 : OR2_X1 port map( A1 => n25798, A2 => n27927, Z => n8301);
   U17978 : OAI21_X2 port map( A1 => n26657, A2 => n25275, B => n467, ZN => 
                           n27928);
   U17985 : NAND2_X1 port map( A1 => n13719, A2 => n13853, ZN => n27929);
   U17988 : NOR2_X2 port map( A1 => n14697, A2 => n17268, ZN => n27931);
   U17990 : NAND2_X2 port map( A1 => n5817, A2 => n8147, ZN => n9650);
   U17992 : AOI21_X2 port map( A1 => n27932, A2 => n11792, B => n22398, ZN => 
                           n22987);
   U17998 : XOR2_X1 port map( A1 => n1436, A2 => n13825, Z => n19409);
   U18000 : OAI21_X2 port map( A1 => n8730, A2 => n18767, B => n8728, ZN => 
                           n13825);
   U18008 : NOR2_X1 port map( A1 => n11204, A2 => n16512, ZN => n27934);
   U18020 : XOR2_X1 port map( A1 => n27935, A2 => n20554, Z => n13201);
   U18021 : XOR2_X1 port map( A1 => n446, A2 => n13971, Z => n27935);
   U18024 : INV_X2 port map( I => n4355, ZN => n451);
   U18032 : NAND2_X2 port map( A1 => n10541, A2 => n852, ZN => n21513);
   U18035 : OAI21_X2 port map( A1 => n10016, A2 => n20260, B => n20098, ZN => 
                           n8854);
   U18046 : INV_X2 port map( I => n27937, ZN => n28541);
   U18049 : XOR2_X1 port map( A1 => n18074, A2 => n22938, Z => n27937);
   U18050 : NOR2_X2 port map( A1 => n27939, A2 => n18524, ZN => n25270);
   U18051 : AOI21_X2 port map( A1 => n28372, A2 => n18523, B => n15246, ZN => 
                           n27939);
   U18054 : NOR2_X2 port map( A1 => n24282, A2 => n6421, ZN => n9789);
   U18071 : XOR2_X1 port map( A1 => n23686, A2 => n20527, Z => n5876);
   U18072 : INV_X2 port map( I => n27175, ZN => n27941);
   U18077 : INV_X2 port map( I => n19052, ZN => n27942);
   U18079 : XOR2_X1 port map( A1 => n27943, A2 => n11886, Z => n14321);
   U18080 : NAND2_X2 port map( A1 => n7296, A2 => n492, ZN => n2447);
   U18087 : NAND3_X1 port map( A1 => n6051, A2 => n20744, A3 => n20751, ZN => 
                           n7515);
   U18088 : XOR2_X1 port map( A1 => n18362, A2 => n18056, Z => n17661);
   U18093 : XOR2_X1 port map( A1 => n18241, A2 => n12230, Z => n18362);
   U18095 : INV_X2 port map( I => n27944, ZN => n985);
   U18103 : XOR2_X1 port map( A1 => n19278, A2 => n19447, Z => n19505);
   U18106 : XOR2_X1 port map( A1 => n8912, A2 => n19350, Z => n19278);
   U18107 : XOR2_X1 port map( A1 => n28243, A2 => n6155, Z => n6780);
   U18109 : NAND2_X1 port map( A1 => n23954, A2 => n22782, ZN => n20295);
   U18117 : XOR2_X1 port map( A1 => n16915, A2 => n16895, Z => n6891);
   U18126 : NAND3_X1 port map( A1 => n20997, A2 => n21000, A3 => n10858, ZN => 
                           n8759);
   U18128 : AND2_X1 port map( A1 => n17559, A2 => n26374, Z => n10692);
   U18137 : AOI21_X2 port map( A1 => n26661, A2 => n4480, B => n4362, ZN => 
                           n4361);
   U18148 : NAND3_X2 port map( A1 => n27946, A2 => n764, A3 => n27945, ZN => 
                           n7324);
   U18149 : INV_X1 port map( I => n27530, ZN => n27945);
   U18152 : XOR2_X1 port map( A1 => n24205, A2 => n24033, Z => n10360);
   U18154 : BUF_X2 port map( I => n3326, Z => n27947);
   U18155 : NAND2_X2 port map( A1 => n5285, A2 => n8554, ZN => n15224);
   U18157 : XOR2_X1 port map( A1 => n4834, A2 => n27949, Z => n21202);
   U18160 : XOR2_X1 port map( A1 => n21200, A2 => n4836, Z => n27949);
   U18163 : XOR2_X1 port map( A1 => n22613, A2 => n27950, Z => n8051);
   U18166 : XOR2_X1 port map( A1 => n20540, A2 => n2474, Z => n27950);
   U18174 : NAND2_X1 port map( A1 => n875, A2 => n23488, ZN => n14461);
   U18177 : OAI21_X1 port map( A1 => n27952, A2 => n24679, B => n6393, ZN => 
                           n5951);
   U18179 : NOR2_X1 port map( A1 => n9401, A2 => n13194, ZN => n27952);
   U18185 : NOR2_X2 port map( A1 => n24495, A2 => n27953, ZN => n21191);
   U18186 : OAI21_X2 port map( A1 => n6813, A2 => n21886, B => n1617, ZN => 
                           n25637);
   U18196 : XOR2_X1 port map( A1 => n17096, A2 => n27955, Z => n27954);
   U18197 : XOR2_X1 port map( A1 => n27956, A2 => n7886, Z => n28238);
   U18209 : NOR2_X2 port map( A1 => n11051, A2 => n23877, ZN => n11049);
   U18211 : NAND3_X2 port map( A1 => n18585, A2 => n7190, A3 => n18583, ZN => 
                           n27957);
   U18219 : INV_X2 port map( I => n19750, ZN => n23869);
   U18220 : AND2_X1 port map( A1 => n19750, A2 => n10041, Z => n10140);
   U18221 : AOI21_X1 port map( A1 => n1017, A2 => n26992, B => n4161, ZN => 
                           n8641);
   U18222 : NAND3_X1 port map( A1 => n28207, A2 => n19903, A3 => n19907, ZN => 
                           n19912);
   U18224 : XOR2_X1 port map( A1 => n10191, A2 => n16936, Z => n2700);
   U18227 : OAI21_X2 port map( A1 => n11793, A2 => n9109, B => n22657, ZN => 
                           n24318);
   U18234 : INV_X2 port map( I => n26297, ZN => n674);
   U18238 : XOR2_X1 port map( A1 => n22693, A2 => n489, Z => n26297);
   U18244 : NAND2_X2 port map( A1 => n25126, A2 => n23092, ZN => n25176);
   U18247 : OAI21_X1 port map( A1 => n10941, A2 => n5345, B => n28546, ZN => 
                           n9738);
   U18249 : NAND2_X2 port map( A1 => n5145, A2 => n5956, ZN => n2434);
   U18251 : NAND2_X2 port map( A1 => n28069, A2 => n5957, ZN => n5145);
   U18252 : NAND2_X2 port map( A1 => n27962, A2 => n5332, ZN => n19880);
   U18259 : XOR2_X1 port map( A1 => n18284, A2 => n26663, Z => n26517);
   U18261 : NOR2_X2 port map( A1 => n24345, A2 => n27963, ZN => n14211);
   U18262 : OAI22_X2 port map( A1 => n10515, A2 => n23677, B1 => n20645, B2 => 
                           n27413, ZN => n4934);
   U18266 : INV_X2 port map( I => n28543, ZN => n28160);
   U18275 : XNOR2_X1 port map( A1 => n8200, A2 => n8202, ZN => n28543);
   U18278 : OAI21_X1 port map( A1 => n9550, A2 => n20852, B => n15724, ZN => 
                           n20980);
   U18291 : AOI21_X2 port map( A1 => n26635, A2 => n20203, B => n14991, ZN => 
                           n24709);
   U18295 : NOR2_X2 port map( A1 => n16730, A2 => n5502, ZN => n14891);
   U18296 : NOR2_X2 port map( A1 => n9262, A2 => n11461, ZN => n16730);
   U18300 : NOR2_X2 port map( A1 => n6231, A2 => n6232, ZN => n3657);
   U18302 : OAI22_X2 port map( A1 => n15825, A2 => n15826, B1 => n15827, B2 => 
                           n16020, ZN => n16649);
   U18304 : NAND2_X1 port map( A1 => n16524, A2 => n6911, ZN => n4839);
   U18306 : NAND2_X2 port map( A1 => n4487, A2 => n4490, ZN => n16524);
   U18310 : NAND2_X2 port map( A1 => n3695, A2 => n27964, ZN => n3694);
   U18311 : NAND3_X2 port map( A1 => n28288, A2 => n17664, A3 => n1209, ZN => 
                           n27964);
   U18312 : XOR2_X1 port map( A1 => n20523, A2 => n23825, Z => n5102);
   U18313 : OAI21_X2 port map( A1 => n1887, A2 => n25294, B => n1954, ZN => 
                           n23825);
   U18318 : XOR2_X1 port map( A1 => n4825, A2 => n4823, Z => n5521);
   U18330 : XOR2_X1 port map( A1 => n11493, A2 => n19497, Z => n4825);
   U18333 : AOI22_X2 port map( A1 => n9554, A2 => n1163, B1 => n18949, B2 => 
                           n21757, ZN => n27966);
   U18335 : XOR2_X1 port map( A1 => n27967, A2 => n13852, Z => n3686);
   U18340 : NAND2_X2 port map( A1 => n11341, A2 => n11343, ZN => n13852);
   U18341 : INV_X2 port map( I => n6878, ZN => n27967);
   U18342 : XOR2_X1 port map( A1 => n5065, A2 => n5063, Z => n7793);
   U18354 : NAND2_X2 port map( A1 => n25752, A2 => n6388, ZN => n18249);
   U18355 : OAI21_X2 port map( A1 => n11712, A2 => n16041, B => n25773, ZN => 
                           n1519);
   U18356 : OAI21_X2 port map( A1 => n17688, A2 => n17801, B => n10871, ZN => 
                           n17690);
   U18357 : OAI21_X2 port map( A1 => n5257, A2 => n5258, B => n27288, ZN => 
                           n16994);
   U18358 : XOR2_X1 port map( A1 => n28013, A2 => n13067, Z => n28438);
   U18364 : XOR2_X1 port map( A1 => n18169, A2 => n18038, Z => n12932);
   U18365 : NAND2_X2 port map( A1 => n28371, A2 => n12085, ZN => n18169);
   U18366 : NAND2_X2 port map( A1 => n17552, A2 => n17551, ZN => n17912);
   U18375 : NAND2_X2 port map( A1 => n27968, A2 => n1546, ZN => n1543);
   U18376 : NAND2_X2 port map( A1 => n28324, A2 => n1055, ZN => n27968);
   U18388 : NAND2_X2 port map( A1 => n11085, A2 => n23791, ZN => n3932);
   U18392 : XOR2_X1 port map( A1 => n25306, A2 => n25445, Z => n18269);
   U18399 : NOR2_X2 port map( A1 => n22528, A2 => n8782, ZN => n25306);
   U18400 : XOR2_X1 port map( A1 => n20483, A2 => n7077, Z => n7076);
   U18408 : NAND3_X1 port map( A1 => n19362, A2 => n19361, A3 => n20235, ZN => 
                           n24749);
   U18409 : NAND2_X2 port map( A1 => n7497, A2 => n7495, ZN => n12934);
   U18413 : NAND2_X2 port map( A1 => n17586, A2 => n25688, ZN => n7497);
   U18418 : BUF_X2 port map( I => n24343, Z => n27969);
   U18419 : BUF_X2 port map( I => n6294, Z => n27970);
   U18420 : INV_X2 port map( I => n27971, ZN => n4832);
   U18421 : XOR2_X1 port map( A1 => n26403, A2 => n12114, Z => n26402);
   U18426 : NOR3_X2 port map( A1 => n18422, A2 => n18420, A3 => n18421, ZN => 
                           n27972);
   U18430 : OAI21_X2 port map( A1 => n27974, A2 => n27973, B => n5887, ZN => 
                           n4610);
   U18433 : NAND2_X1 port map( A1 => n15106, A2 => n16102, ZN => n9020);
   U18437 : OAI21_X2 port map( A1 => n27978, A2 => n22150, B => n14943, ZN => 
                           n14878);
   U18441 : NAND3_X2 port map( A1 => n27979, A2 => n10745, A3 => n23322, ZN => 
                           n13042);
   U18444 : INV_X1 port map( I => n22056, ZN => n27979);
   U18448 : XOR2_X1 port map( A1 => n19224, A2 => n1975, Z => n19351);
   U18458 : NAND3_X2 port map( A1 => n1896, A2 => n1898, A3 => n1895, ZN => 
                           n1975);
   U18459 : NAND2_X1 port map( A1 => n27980, A2 => n7442, ZN => n25007);
   U18466 : NOR2_X1 port map( A1 => n7440, A2 => n7441, ZN => n27980);
   U18469 : XOR2_X1 port map( A1 => n3251, A2 => n27981, Z => n19666);
   U18473 : XOR2_X1 port map( A1 => n19530, A2 => n14496, Z => n27981);
   U18476 : BUF_X4 port map( I => n19615, Z => n19889);
   U18477 : XOR2_X1 port map( A1 => n18269, A2 => n18267, Z => n5129);
   U18478 : NOR2_X2 port map( A1 => n12584, A2 => n23575, ZN => n24743);
   U18493 : NAND2_X2 port map( A1 => n14767, A2 => n26309, ZN => n23575);
   U18494 : INV_X2 port map( I => n27982, ZN => n15255);
   U18498 : NAND3_X1 port map( A1 => n16203, A2 => n24581, A3 => n16201, ZN => 
                           n15643);
   U18499 : NAND3_X1 port map( A1 => n9698, A2 => n9358, A3 => n17527, ZN => 
                           n9697);
   U18503 : OAI21_X2 port map( A1 => n10015, A2 => n14324, B => n17421, ZN => 
                           n9698);
   U18505 : AOI21_X2 port map( A1 => n11616, A2 => n27985, B => n22758, ZN => 
                           n11543);
   U18506 : NAND2_X1 port map( A1 => n4782, A2 => n4311, ZN => n27985);
   U18507 : NAND2_X2 port map( A1 => n1798, A2 => n1797, ZN => n23231);
   U18508 : NOR2_X2 port map( A1 => n20938, A2 => n20933, ZN => n27988);
   U18509 : NAND2_X2 port map( A1 => n2566, A2 => n2567, ZN => n17766);
   U18510 : OR2_X2 port map( A1 => n15255, A2 => n26615, Z => n17528);
   U18514 : OAI22_X1 port map( A1 => n1986, A2 => n4647, B1 => n15943, B2 => 
                           n1987, ZN => n23647);
   U18516 : XOR2_X1 port map( A1 => n4423, A2 => n4425, Z => n7854);
   U18517 : OR2_X1 port map( A1 => n13786, A2 => n16426, Z => n27989);
   U18519 : NAND2_X1 port map( A1 => n26202, A2 => n18759, ZN => n27991);
   U18521 : AND2_X1 port map( A1 => n25381, A2 => n2346, Z => n28043);
   U18523 : OAI21_X1 port map( A1 => n3980, A2 => n17540, B => n24821, ZN => 
                           n15395);
   U18526 : AOI22_X2 port map( A1 => n27992, A2 => n4452, B1 => n2894, B2 => 
                           n24454, ZN => n18882);
   U18530 : NOR2_X2 port map( A1 => n24454, A2 => n24573, ZN => n27992);
   U18532 : NAND2_X2 port map( A1 => n20173, A2 => n20267, ZN => n27993);
   U18542 : XOR2_X1 port map( A1 => n14166, A2 => n9673, Z => n26334);
   U18545 : XOR2_X1 port map( A1 => n9952, A2 => n9650, Z => n9673);
   U18548 : XOR2_X1 port map( A1 => n3594, A2 => n3595, Z => n5403);
   U18554 : NAND2_X1 port map( A1 => n15105, A2 => n27994, ZN => n1616);
   U18564 : AOI21_X1 port map( A1 => n16239, A2 => n9768, B => n16316, ZN => 
                           n27994);
   U18570 : XOR2_X1 port map( A1 => n27995, A2 => n22315, Z => Ciphertext(71));
   U18572 : XOR2_X1 port map( A1 => n4966, A2 => n9445, Z => n10248);
   U18574 : XOR2_X1 port map( A1 => n19444, A2 => n18591, Z => n27997);
   U18575 : XOR2_X1 port map( A1 => n19556, A2 => n23667, Z => n9281);
   U18600 : XOR2_X1 port map( A1 => n21305, A2 => n21249, Z => n20438);
   U18613 : AOI21_X2 port map( A1 => n8774, A2 => n13864, B => n8773, ZN => 
                           n21305);
   U18625 : XOR2_X1 port map( A1 => n13585, A2 => n15242, Z => n3224);
   U18628 : NAND2_X2 port map( A1 => n23204, A2 => n23808, ZN => n13585);
   U18637 : XOR2_X1 port map( A1 => n25311, A2 => n21152, Z => n20765);
   U18639 : NAND2_X2 port map( A1 => n26643, A2 => n17766, ZN => n12670);
   U18640 : NAND2_X2 port map( A1 => n25095, A2 => n6635, ZN => n6373);
   U18650 : NAND2_X2 port map( A1 => n11861, A2 => n12594, ZN => n20018);
   U18654 : NOR2_X2 port map( A1 => n23355, A2 => n278, ZN => n11861);
   U18655 : XOR2_X1 port map( A1 => n28000, A2 => n13982, Z => n6251);
   U18660 : XOR2_X1 port map( A1 => n13354, A2 => n6025, Z => n28000);
   U18664 : NOR2_X2 port map( A1 => n2868, A2 => n9701, ZN => n28001);
   U18668 : XOR2_X1 port map( A1 => n7589, A2 => n7588, Z => n28115);
   U18669 : NAND3_X2 port map( A1 => n12487, A2 => n20884, A3 => n20883, ZN => 
                           n12486);
   U18672 : NAND2_X1 port map( A1 => n18739, A2 => n18741, ZN => n18565);
   U18678 : OR3_X1 port map( A1 => n19126, A2 => n19124, A3 => n2617, Z => 
                           n24489);
   U18690 : NAND2_X2 port map( A1 => n11937, A2 => n14737, ZN => n28005);
   U18695 : XOR2_X1 port map( A1 => n9655, A2 => n13253, Z => n20446);
   U18697 : NOR2_X2 port map( A1 => n21905, A2 => n11937, ZN => n13423);
   U18702 : INV_X2 port map( I => n16678, ZN => n28008);
   U18703 : NAND2_X2 port map( A1 => n1049, A2 => n13758, ZN => n4169);
   U18704 : XOR2_X1 port map( A1 => n28010, A2 => n1305, Z => Ciphertext(70));
   U18708 : AOI22_X1 port map( A1 => n12540, A2 => n24734, B1 => n928, B2 => 
                           n12538, ZN => n28010);
   U18709 : XOR2_X1 port map( A1 => n2264, A2 => n16985, Z => n4988);
   U18711 : XOR2_X1 port map( A1 => n16784, A2 => n24343, Z => n2264);
   U18712 : NOR2_X2 port map( A1 => n11373, A2 => n7102, ZN => n7599);
   U18720 : NAND2_X2 port map( A1 => n8750, A2 => n8749, ZN => n7102);
   U18726 : NAND3_X1 port map( A1 => n24936, A2 => n24935, A3 => n1159, ZN => 
                           n28506);
   U18727 : OR2_X2 port map( A1 => n13411, A2 => n3389, Z => n11763);
   U18728 : XOR2_X1 port map( A1 => n15593, A2 => n24254, Z => n13411);
   U18734 : XOR2_X1 port map( A1 => n11046, A2 => n27366, Z => n20512);
   U18735 : NAND3_X2 port map( A1 => n12847, A2 => n7048, A3 => n20332, ZN => 
                           n11046);
   U18741 : NAND2_X2 port map( A1 => n22192, A2 => n18864, ZN => n8636);
   U18747 : NAND2_X2 port map( A1 => n26211, A2 => n11309, ZN => n12180);
   U18752 : BUF_X2 port map( I => n3179, Z => n28013);
   U18754 : NAND3_X1 port map( A1 => n23771, A2 => n9899, A3 => n27454, ZN => 
                           n19395);
   U18759 : NAND2_X2 port map( A1 => n28016, A2 => n28015, ZN => n28014);
   U18780 : INV_X2 port map( I => n24539, ZN => n28015);
   U18782 : OAI21_X1 port map( A1 => n28019, A2 => n18879, B => n23488, ZN => 
                           n28227);
   U18788 : OR2_X1 port map( A1 => n11318, A2 => n13056, Z => n20836);
   U18793 : BUF_X2 port map( I => n10588, Z => n28017);
   U18798 : XOR2_X1 port map( A1 => n19444, A2 => n19443, Z => n28018);
   U18802 : OAI21_X2 port map( A1 => n21509, A2 => n21507, B => n28020, ZN => 
                           n8816);
   U18808 : XOR2_X1 port map( A1 => n28021, A2 => n20208, Z => Ciphertext(176))
                           ;
   U18809 : AOI22_X2 port map( A1 => n9725, A2 => n16587, B1 => n16585, B2 => 
                           n16584, ZN => n9288);
   U18812 : NAND2_X2 port map( A1 => n19718, A2 => n11973, ZN => n9579);
   U18813 : NOR2_X2 port map( A1 => n21663, A2 => n27395, ZN => n9140);
   U18814 : NAND2_X2 port map( A1 => n22653, A2 => n22652, ZN => n21663);
   U18815 : INV_X2 port map( I => n28022, ZN => n24916);
   U18817 : INV_X2 port map( I => n237, ZN => n28022);
   U18819 : NAND2_X2 port map( A1 => n25685, A2 => n1247, ZN => n16669);
   U18823 : AOI21_X2 port map( A1 => n10015, A2 => n26615, B => n17421, ZN => 
                           n28023);
   U18830 : NAND3_X2 port map( A1 => n28024, A2 => n18635, A3 => n18634, ZN => 
                           n23546);
   U18831 : XOR2_X1 port map( A1 => n6559, A2 => n26052, Z => n25407);
   U18832 : INV_X4 port map( I => n20268, ZN => n806);
   U18837 : NAND2_X2 port map( A1 => n19944, A2 => n19943, ZN => n20268);
   U18851 : INV_X4 port map( I => n12053, ZN => n21040);
   U18855 : BUF_X4 port map( I => n103, Z => n28186);
   U18856 : NAND2_X2 port map( A1 => n11049, A2 => n2876, ZN => n20489);
   U18858 : XOR2_X1 port map( A1 => n25343, A2 => n5420, Z => n28474);
   U18863 : AOI21_X2 port map( A1 => n3906, A2 => n3905, B => n18789, ZN => 
                           n25343);
   U18868 : AOI22_X1 port map( A1 => n21599, A2 => n21608, B1 => n21603, B2 => 
                           n15475, ZN => n24432);
   U18873 : XOR2_X1 port map( A1 => n22130, A2 => n6597, Z => n5401);
   U18885 : AOI21_X2 port map( A1 => n13604, A2 => n13605, B => n13606, ZN => 
                           n1651);
   U18891 : OAI21_X1 port map( A1 => n4082, A2 => n20964, B => n20957, ZN => 
                           n139);
   U18892 : NAND2_X2 port map( A1 => n20964, A2 => n4413, ZN => n20957);
   U18906 : NAND3_X2 port map( A1 => n25602, A2 => n25603, A3 => n13422, ZN => 
                           n23181);
   U18909 : OR2_X2 port map( A1 => n3433, A2 => n5226, Z => n13662);
   U18910 : OAI21_X2 port map( A1 => n14618, A2 => n26103, B => n22660, ZN => 
                           n2853);
   U18911 : NOR2_X2 port map( A1 => n28028, A2 => n9743, ZN => n28518);
   U18914 : NAND2_X2 port map( A1 => n19814, A2 => n19815, ZN => n21257);
   U18916 : XOR2_X1 port map( A1 => n19200, A2 => n7050, Z => n7309);
   U18918 : XOR2_X1 port map( A1 => n19549, A2 => n19485, Z => n8503);
   U18921 : INV_X1 port map( I => n23488, ZN => n8998);
   U18923 : XOR2_X1 port map( A1 => n20565, A2 => n22791, Z => n20762);
   U18928 : XOR2_X1 port map( A1 => n8150, A2 => n18214, Z => n3580);
   U18931 : NAND2_X2 port map( A1 => n22776, A2 => n20064, ZN => n11583);
   U18932 : XOR2_X1 port map( A1 => n9228, A2 => n28030, Z => n28350);
   U18934 : XOR2_X1 port map( A1 => n28466, A2 => n14537, Z => n28030);
   U18935 : NAND3_X2 port map( A1 => n15288, A2 => n24136, A3 => n20487, ZN => 
                           n20626);
   U18949 : INV_X2 port map( I => n22873, ZN => n28031);
   U18950 : INV_X1 port map( I => n3573, ZN => n4942);
   U18952 : INV_X1 port map( I => n15859, ZN => n28032);
   U18953 : OAI21_X2 port map( A1 => n16934, A2 => n17409, B => n28034, ZN => 
                           n9485);
   U18958 : OAI21_X2 port map( A1 => n24779, A2 => n8335, B => n28035, ZN => 
                           n28034);
   U18959 : INV_X2 port map( I => n6294, ZN => n28035);
   U18960 : NAND3_X2 port map( A1 => n22537, A2 => n25559, A3 => n13, ZN => 
                           n25242);
   U18966 : NOR3_X2 port map( A1 => n27345, A2 => n26410, A3 => n20314, ZN => 
                           n13399);
   U18967 : XOR2_X1 port map( A1 => n20529, A2 => n28041, Z => n9514);
   U18970 : NAND3_X1 port map( A1 => n7566, A2 => n11059, A3 => n14631, ZN => 
                           n4907);
   U18972 : XOR2_X1 port map( A1 => n2370, A2 => n23007, Z => n2369);
   U18974 : XOR2_X1 port map( A1 => n2979, A2 => n13116, Z => n15573);
   U18976 : NAND2_X1 port map( A1 => n8100, A2 => n9899, ZN => n12603);
   U18978 : NAND2_X2 port map( A1 => n22195, A2 => n2314, ZN => n8100);
   U18980 : OAI21_X2 port map( A1 => n28042, A2 => n18340, B => n18339, ZN => 
                           n19305);
   U18982 : INV_X2 port map( I => n5445, ZN => n28224);
   U18987 : NAND2_X2 port map( A1 => n9571, A2 => n9568, ZN => n7321);
   U18991 : XOR2_X1 port map( A1 => n9832, A2 => n28044, Z => n6631);
   U18993 : XOR2_X1 port map( A1 => n18061, A2 => n25946, Z => n28044);
   U18994 : XOR2_X1 port map( A1 => n18103, A2 => n18217, Z => n9832);
   U18997 : XOR2_X1 port map( A1 => n14962, A2 => n28045, Z => n8710);
   U18998 : XOR2_X1 port map( A1 => n24528, A2 => n19412, Z => n28045);
   U19009 : OAI21_X2 port map( A1 => n22929, A2 => n28046, B => n4555, ZN => 
                           n16642);
   U19014 : NOR2_X1 port map( A1 => n16639, A2 => n16640, ZN => n28046);
   U19015 : OAI22_X2 port map( A1 => n16014, A2 => n16011, B1 => n16010, B2 => 
                           n16009, ZN => n26205);
   U19017 : AND2_X1 port map( A1 => n23437, A2 => n17726, Z => n6179);
   U19026 : NAND2_X2 port map( A1 => n9419, A2 => n23547, ZN => n23437);
   U19033 : NOR2_X2 port map( A1 => n28047, A2 => n1769, ZN => n21647);
   U19034 : NAND2_X2 port map( A1 => n1768, A2 => n1767, ZN => n28047);
   U19046 : NOR3_X2 port map( A1 => n25935, A2 => n758, A3 => n879, ZN => 
                           n28048);
   U19055 : NAND2_X2 port map( A1 => n2482, A2 => n2483, ZN => n9683);
   U19062 : XOR2_X1 port map( A1 => n28049, A2 => n9054, Z => n2041);
   U19063 : XOR2_X1 port map( A1 => n26278, A2 => n1947, Z => n28049);
   U19065 : XOR2_X1 port map( A1 => n4633, A2 => n17031, Z => n23703);
   U19066 : XNOR2_X1 port map( A1 => n14753, A2 => n26246, ZN => n4633);
   U19076 : XOR2_X1 port map( A1 => n19345, A2 => n28050, Z => n23343);
   U19081 : XOR2_X1 port map( A1 => n24275, A2 => n10331, Z => n28050);
   U19083 : XOR2_X1 port map( A1 => n17008, A2 => n17092, Z => n3038);
   U19097 : XOR2_X1 port map( A1 => n22926, A2 => n3039, Z => n17092);
   U19099 : INV_X1 port map( I => n20569, ZN => n20574);
   U19107 : NOR2_X2 port map( A1 => n28051, A2 => n12566, ZN => n19552);
   U19108 : AOI21_X2 port map( A1 => n25109, A2 => n13490, B => n12978, ZN => 
                           n28051);
   U19113 : XOR2_X1 port map( A1 => n17780, A2 => n28052, Z => n23841);
   U19116 : XOR2_X1 port map( A1 => n13807, A2 => n18242, Z => n28052);
   U19117 : AOI22_X2 port map( A1 => n28053, A2 => n1158, B1 => n447, B2 => 
                           n14419, ZN => n5900);
   U19118 : NAND2_X1 port map( A1 => n4058, A2 => n22783, ZN => n28054);
   U19126 : NOR2_X2 port map( A1 => n25940, A2 => n16380, ZN => n16686);
   U19130 : OAI21_X2 port map( A1 => n15867, A2 => n9443, B => n26388, ZN => 
                           n16380);
   U19133 : NAND2_X2 port map( A1 => n20430, A2 => n14611, ZN => n20102);
   U19136 : NAND2_X2 port map( A1 => n19853, A2 => n19854, ZN => n14611);
   U19140 : XOR2_X1 port map( A1 => n19233, A2 => n27421, Z => n19358);
   U19152 : NAND2_X2 port map( A1 => n5900, A2 => n13239, ZN => n19233);
   U19155 : NAND3_X1 port map( A1 => n13928, A2 => n1365, A3 => n10181, ZN => 
                           n28056);
   U19156 : INV_X1 port map( I => n9634, ZN => n28057);
   U19163 : BUF_X2 port map( I => n22050, Z => n28058);
   U19164 : OAI21_X2 port map( A1 => n28061, A2 => n28060, B => n6642, ZN => 
                           n12618);
   U19166 : NOR2_X1 port map( A1 => n21791, A2 => n14342, ZN => n28060);
   U19170 : INV_X1 port map( I => n23020, ZN => n28061);
   U19171 : XOR2_X1 port map( A1 => n28062, A2 => n7010, Z => n10542);
   U19177 : XOR2_X1 port map( A1 => n27847, A2 => n25039, Z => n28062);
   U19178 : NAND3_X2 port map( A1 => n28063, A2 => n15285, A3 => n24130, ZN => 
                           n20447);
   U19179 : OR2_X1 port map( A1 => n18739, A2 => n23538, Z => n28082);
   U19184 : INV_X1 port map( I => n24038, ZN => n9434);
   U19185 : XOR2_X1 port map( A1 => n28064, A2 => n16791, Z => n1392);
   U19189 : AND2_X1 port map( A1 => n17594, A2 => n3929, Z => n26267);
   U19191 : OAI21_X2 port map( A1 => n28066, A2 => n28065, B => n3533, ZN => 
                           n23951);
   U19207 : NOR2_X1 port map( A1 => n10603, A2 => n27662, ZN => n28066);
   U19215 : NAND2_X2 port map( A1 => n9854, A2 => n7002, ZN => n14980);
   U19230 : OAI21_X2 port map( A1 => n5954, A2 => n4461, B => n17830, ZN => 
                           n7002);
   U19260 : INV_X4 port map( I => n13502, ZN => n28492);
   U19267 : BUF_X2 port map( I => n14459, Z => n28068);
   U19268 : XOR2_X1 port map( A1 => n21148, A2 => n9397, Z => n20534);
   U19272 : NAND2_X1 port map( A1 => n13349, A2 => n988, ZN => n19036);
   U19273 : XOR2_X1 port map( A1 => n28072, A2 => n7201, Z => n25133);
   U19276 : XOR2_X1 port map( A1 => n25634, A2 => n28073, Z => n28072);
   U19277 : INV_X2 port map( I => n28075, ZN => n2631);
   U19279 : NAND2_X2 port map( A1 => n28394, A2 => n14274, ZN => n10513);
   U19280 : INV_X4 port map( I => n4813, ZN => n4812);
   U19283 : NAND2_X2 port map( A1 => n4816, A2 => n17246, ZN => n4813);
   U19285 : XOR2_X1 port map( A1 => n18263, A2 => n25901, Z => n18264);
   U19289 : XOR2_X1 port map( A1 => n3706, A2 => n5876, Z => n3705);
   U19296 : XOR2_X1 port map( A1 => n28076, A2 => n16964, Z => n7914);
   U19298 : XOR2_X1 port map( A1 => n27936, A2 => n28510, Z => n28076);
   U19302 : NAND2_X1 port map( A1 => n10497, A2 => n23684, ZN => n17533);
   U19305 : XOR2_X1 port map( A1 => n28117, A2 => n7279, Z => n28077);
   U19310 : NAND3_X1 port map( A1 => n20997, A2 => n20998, A3 => n12045, ZN => 
                           n20993);
   U19311 : XOR2_X1 port map( A1 => n16894, A2 => n16893, Z => n28103);
   U19315 : XOR2_X1 port map( A1 => n25785, A2 => n11680, Z => n16894);
   U19316 : NOR2_X2 port map( A1 => n8181, A2 => n12434, ZN => n24351);
   U19322 : AOI21_X1 port map( A1 => n13395, A2 => n21007, B => n1431, ZN => 
                           n12613);
   U19324 : AOI22_X1 port map( A1 => n3583, A2 => n21174, B1 => n2230, B2 => 
                           n22751, ZN => n23383);
   U19325 : XOR2_X1 port map( A1 => n22939, A2 => n28078, Z => n21839);
   U19329 : INV_X1 port map( I => n14593, ZN => n28078);
   U19330 : NAND2_X2 port map( A1 => n28079, A2 => n2891, ZN => n14075);
   U19335 : INV_X2 port map( I => n20112, ZN => n28079);
   U19338 : NAND2_X2 port map( A1 => n1133, A2 => n10613, ZN => n20112);
   U19343 : NAND2_X2 port map( A1 => n28080, A2 => n25845, ZN => n10443);
   U19344 : NOR2_X1 port map( A1 => n9753, A2 => n9754, ZN => n28080);
   U19345 : OAI21_X2 port map( A1 => n28297, A2 => n23626, B => n6391, ZN => 
                           n26206);
   U19349 : OAI22_X2 port map( A1 => n10874, A2 => n27830, B1 => n25355, B2 => 
                           n10873, ZN => n12735);
   U19350 : XOR2_X1 port map( A1 => n5351, A2 => n27422, Z => n14011);
   U19356 : NAND2_X2 port map( A1 => n3150, A2 => n5467, ZN => n28446);
   U19357 : NOR2_X2 port map( A1 => n22910, A2 => n15970, ZN => n15808);
   U19359 : INV_X2 port map( I => n14542, ZN => n15970);
   U19362 : XOR2_X1 port map( A1 => Plaintext(183), A2 => Key(183), Z => n14542
                           );
   U19369 : NAND2_X2 port map( A1 => n4880, A2 => n25300, ZN => n4518);
   U19370 : AOI21_X2 port map( A1 => n7288, A2 => n28082, B => n14498, ZN => 
                           n6908);
   U19374 : XOR2_X1 port map( A1 => n761, A2 => n18237, Z => n28084);
   U19377 : NOR2_X2 port map( A1 => n28085, A2 => n10685, ZN => n14617);
   U19382 : NOR2_X1 port map( A1 => n9892, A2 => n10453, ZN => n28085);
   U19384 : NAND2_X2 port map( A1 => n28260, A2 => n10444, ZN => n13768);
   U19386 : OAI21_X2 port map( A1 => n5926, A2 => n12611, B => n28086, ZN => 
                           n15182);
   U19389 : AOI22_X2 port map( A1 => n25532, A2 => n17159, B1 => n3943, B2 => 
                           n17986, ZN => n28086);
   U19390 : XOR2_X1 port map( A1 => n10285, A2 => n28089, Z => n28362);
   U19394 : XOR2_X1 port map( A1 => n8132, A2 => n10358, Z => n19492);
   U19396 : NOR2_X2 port map( A1 => n8120, A2 => n8121, ZN => n10358);
   U19401 : XOR2_X1 port map( A1 => n14428, A2 => n16749, Z => n13557);
   U19407 : XOR2_X1 port map( A1 => n21974, A2 => n23967, Z => n9756);
   U19408 : NAND2_X2 port map( A1 => n5139, A2 => n14542, ZN => n16267);
   U19412 : BUF_X2 port map( I => n18639, Z => n28090);
   U19435 : AOI22_X2 port map( A1 => n28092, A2 => n27885, B1 => n21464, B2 => 
                           n21465, ZN => n21481);
   U19436 : OAI21_X2 port map( A1 => n23741, A2 => n21463, B => n21462, ZN => 
                           n28092);
   U19437 : OR2_X1 port map( A1 => n7379, A2 => n2706, Z => n9168);
   U19439 : XOR2_X1 port map( A1 => n28093, A2 => n6164, Z => n8656);
   U19442 : XOR2_X1 port map( A1 => n9597, A2 => n26122, Z => n28093);
   U19448 : XOR2_X1 port map( A1 => n28094, A2 => n13082, Z => Ciphertext(9));
   U19452 : BUF_X2 port map( I => n10291, Z => n28095);
   U19456 : XOR2_X1 port map( A1 => n13089, A2 => n28096, Z => n28149);
   U19458 : OR2_X1 port map( A1 => n25455, A2 => n2706, Z => n28098);
   U19459 : OAI21_X2 port map( A1 => n7129, A2 => n19783, B => n28099, ZN => 
                           n25668);
   U19460 : NOR2_X2 port map( A1 => n14314, A2 => n14313, ZN => n9455);
   U19463 : NAND2_X2 port map( A1 => n9373, A2 => n9372, ZN => n14314);
   U19471 : INV_X2 port map( I => n28100, ZN => n9370);
   U19472 : XNOR2_X1 port map( A1 => n2666, A2 => n25741, ZN => n28100);
   U19473 : XOR2_X1 port map( A1 => n28101, A2 => n20952, Z => Ciphertext(63));
   U19474 : NAND2_X1 port map( A1 => n4606, A2 => n23980, ZN => n28101);
   U19477 : NAND2_X2 port map( A1 => n5614, A2 => n15939, ZN => n28113);
   U19488 : INV_X2 port map( I => n20224, ZN => n5198);
   U19489 : NAND2_X2 port map( A1 => n22916, A2 => n22376, ZN => n20224);
   U19492 : AOI22_X1 port map( A1 => n20655, A2 => n4766, B1 => n23119, B2 => 
                           n20656, ZN => n25258);
   U19502 : INV_X2 port map( I => n28102, ZN => n15448);
   U19504 : NAND2_X2 port map( A1 => n25024, A2 => n2150, ZN => n24190);
   U19508 : XOR2_X1 port map( A1 => n883, A2 => n9250, Z => n12548);
   U19510 : OR2_X1 port map( A1 => n11404, A2 => n25955, Z => n18723);
   U19513 : XOR2_X1 port map( A1 => n19313, A2 => n6445, Z => n19325);
   U19522 : AOI22_X1 port map( A1 => n6897, A2 => n21736, B1 => n2407, B2 => 
                           n8771, ZN => n28226);
   U19530 : XOR2_X1 port map( A1 => n17106, A2 => n16964, Z => n16968);
   U19532 : XOR2_X1 port map( A1 => n10943, A2 => n28103, Z => n17217);
   U19533 : INV_X2 port map( I => n26218, ZN => n28105);
   U19540 : BUF_X2 port map( I => n1177, Z => n28106);
   U19541 : XOR2_X1 port map( A1 => n5914, A2 => n21255, Z => n20513);
   U19551 : NAND2_X2 port map( A1 => n24553, A2 => n8032, ZN => n9956);
   U19552 : NAND2_X2 port map( A1 => n28108, A2 => n28107, ZN => n9667);
   U19556 : NAND3_X2 port map( A1 => n2202, A2 => n2203, A3 => n7165, ZN => 
                           n4760);
   U19557 : NAND2_X2 port map( A1 => n12689, A2 => n28109, ZN => n7379);
   U19565 : OAI21_X2 port map( A1 => n10700, A2 => n14568, B => n19632, ZN => 
                           n28109);
   U19570 : NAND2_X1 port map( A1 => n8611, A2 => n24811, ZN => n13920);
   U19572 : XOR2_X1 port map( A1 => n19552, A2 => n4768, Z => n19219);
   U19581 : NAND2_X2 port map( A1 => n23331, A2 => n4759, ZN => n4768);
   U19591 : OAI21_X1 port map( A1 => n9877, A2 => n20314, B => n15544, ZN => 
                           n14811);
   U19593 : INV_X1 port map( I => n23146, ZN => n957);
   U19600 : OR2_X1 port map( A1 => n23146, A2 => n2231, Z => n3967);
   U19602 : XOR2_X1 port map( A1 => n28114, A2 => n7362, Z => Ciphertext(159));
   U19606 : INV_X2 port map( I => n28115, ZN => n7587);
   U19610 : NAND3_X2 port map( A1 => n28116, A2 => n8029, A3 => n8030, ZN => 
                           n4890);
   U19611 : NAND3_X2 port map( A1 => n28200, A2 => n950, A3 => n13440, ZN => 
                           n28116);
   U19627 : XOR2_X1 port map( A1 => n16980, A2 => n21449, Z => n442);
   U19631 : NAND3_X2 port map( A1 => n28329, A2 => n5915, A3 => n13495, ZN => 
                           n16980);
   U19632 : XOR2_X1 port map( A1 => n25853, A2 => n19324, Z => n28117);
   U19636 : BUF_X2 port map( I => n17818, Z => n28118);
   U19637 : INV_X2 port map( I => n16461, ZN => n1049);
   U19638 : NAND2_X2 port map( A1 => n10450, A2 => n15772, ZN => n16461);
   U19639 : NAND3_X2 port map( A1 => n5750, A2 => n323, A3 => n322, ZN => n9216
                           );
   U19642 : XOR2_X1 port map( A1 => n22254, A2 => n4427, Z => n4140);
   U19647 : NAND3_X1 port map( A1 => n10870, A2 => n12358, A3 => n12272, ZN => 
                           n10869);
   U19648 : OAI22_X2 port map( A1 => n28119, A2 => n10522, B1 => n24431, B2 => 
                           n10521, ZN => n19978);
   U19650 : XOR2_X1 port map( A1 => n28120, A2 => n15519, Z => Ciphertext(189))
                           ;
   U19652 : NOR2_X1 port map( A1 => n15520, A2 => n26326, ZN => n28120);
   U19654 : NOR2_X2 port map( A1 => n17895, A2 => n17766, ZN => n17873);
   U19655 : BUF_X2 port map( I => n2910, Z => n28122);
   U19656 : NAND2_X1 port map( A1 => n27401, A2 => n2492, ZN => n21801);
   U19657 : XOR2_X1 port map( A1 => n27421, A2 => n12648, Z => n14091);
   U19660 : NAND2_X2 port map( A1 => n9350, A2 => n9349, ZN => n12648);
   U19666 : NAND2_X1 port map( A1 => n9057, A2 => n21716, ZN => n28123);
   U19671 : OR2_X1 port map( A1 => n7870, A2 => n7587, Z => n4548);
   U19673 : NAND2_X2 port map( A1 => n28124, A2 => n18858, ZN => n19388);
   U19674 : NOR2_X2 port map( A1 => n469, A2 => n23760, ZN => n18914);
   U19676 : NOR2_X2 port map( A1 => n835, A2 => n5081, ZN => n28125);
   U19679 : INV_X2 port map( I => n13481, ZN => n28126);
   U19681 : XOR2_X1 port map( A1 => n19505, A2 => n28127, Z => n28301);
   U19684 : XOR2_X1 port map( A1 => n2430, A2 => n28128, Z => n28127);
   U19685 : NOR2_X2 port map( A1 => n21824, A2 => n3964, ZN => n26062);
   U19687 : NAND2_X2 port map( A1 => n24774, A2 => n1892, ZN => n28129);
   U19688 : NAND2_X2 port map( A1 => n28131, A2 => n13979, ZN => n5452);
   U19693 : XOR2_X1 port map( A1 => n18280, A2 => n8432, Z => n15488);
   U19694 : NAND2_X2 port map( A1 => n17451, A2 => n14106, ZN => n9691);
   U19696 : XOR2_X1 port map( A1 => n21158, A2 => n21424, Z => n20725);
   U19701 : XOR2_X1 port map( A1 => n4674, A2 => n28132, Z => n8193);
   U19702 : XOR2_X1 port map( A1 => n17045, A2 => n4673, Z => n28132);
   U19705 : NAND3_X1 port map( A1 => n24044, A2 => n15475, A3 => n21606, ZN => 
                           n13831);
   U19711 : NOR3_X1 port map( A1 => n16132, A2 => n15923, A3 => n15981, ZN => 
                           n10685);
   U19712 : AOI21_X2 port map( A1 => n19094, A2 => n3619, B => n8122, ZN => 
                           n8132);
   U19717 : INV_X2 port map( I => n28133, ZN => n28553);
   U19718 : XOR2_X1 port map( A1 => n8885, A2 => n21553, Z => n22684);
   U19721 : AOI22_X2 port map( A1 => n1478, A2 => n26065, B1 => n50, B2 => 
                           n20209, ZN => n8885);
   U19723 : INV_X2 port map( I => n28135, ZN => n28542);
   U19727 : BUF_X2 port map( I => n12667, Z => n28136);
   U19736 : NAND2_X2 port map( A1 => n3974, A2 => n28137, ZN => n12055);
   U19738 : NAND2_X1 port map( A1 => n28139, A2 => n28138, ZN => n28137);
   U19742 : NOR2_X1 port map( A1 => n21016, A2 => n15728, ZN => n28138);
   U19746 : INV_X2 port map( I => n20972, ZN => n28139);
   U19747 : NAND2_X2 port map( A1 => n194, A2 => n14947, ZN => n22374);
   U19757 : NAND2_X2 port map( A1 => n9825, A2 => n28140, ZN => n8723);
   U19764 : AOI22_X2 port map( A1 => n19631, A2 => n19774, B1 => n28268, B2 => 
                           n9896, ZN => n28140);
   U19766 : XOR2_X1 port map( A1 => n21190, A2 => n27437, Z => n21150);
   U19770 : NOR2_X1 port map( A1 => n7446, A2 => n12221, ZN => n12832);
   U19772 : NAND2_X2 port map( A1 => n28518, A2 => n6768, ZN => n19350);
   U19782 : NOR2_X2 port map( A1 => n14212, A2 => n13197, ZN => n23923);
   U19793 : XOR2_X1 port map( A1 => n28142, A2 => n925, Z => Ciphertext(191));
   U19798 : AOI22_X1 port map( A1 => n25645, A2 => n24685, B1 => n2407, B2 => 
                           n9458, ZN => n28142);
   U19801 : XOR2_X1 port map( A1 => n19291, A2 => n15493, Z => n19679);
   U19807 : NOR2_X2 port map( A1 => n16556, A2 => n4938, ZN => n1595);
   U19808 : OAI21_X2 port map( A1 => n15040, A2 => n14654, B => n15435, ZN => 
                           n28143);
   U19812 : AOI21_X2 port map( A1 => n15862, A2 => n16034, B => n16303, ZN => 
                           n28144);
   U19817 : NAND2_X2 port map( A1 => n16471, A2 => n4518, ZN => n16556);
   U19825 : NOR2_X2 port map( A1 => n22260, A2 => n15223, ZN => n28145);
   U19826 : XOR2_X1 port map( A1 => n5432, A2 => n13412, Z => n9001);
   U19831 : NAND2_X2 port map( A1 => n18827, A2 => n4381, ZN => n28453);
   U19837 : NAND2_X2 port map( A1 => n28146, A2 => n28522, ZN => n10810);
   U19841 : BUF_X2 port map( I => n19148, Z => n28147);
   U19843 : OAI22_X2 port map( A1 => n11, A2 => n11325, B1 => n16077, B2 => 
                           n16076, ZN => n16346);
   U19844 : INV_X1 port map( I => n15905, ZN => n11325);
   U19846 : XOR2_X1 port map( A1 => Key(11), A2 => Plaintext(11), Z => n15905);
   U19849 : OAI21_X2 port map( A1 => n2626, A2 => n1878, B => n2523, ZN => 
                           n1877);
   U19853 : OAI21_X2 port map( A1 => n10461, A2 => n8125, B => n24560, ZN => 
                           n9570);
   U19855 : OAI21_X1 port map( A1 => n18718, A2 => n18719, B => n18658, ZN => 
                           n22430);
   U19856 : XOR2_X1 port map( A1 => n28150, A2 => n21934, Z => n23258);
   U19859 : INV_X2 port map( I => n8100, ZN => n28151);
   U19862 : NOR2_X2 port map( A1 => n887, A2 => n24316, ZN => n11858);
   U19863 : BUF_X2 port map( I => n5140, Z => n28152);
   U19869 : NAND2_X2 port map( A1 => n28155, A2 => n28153, ZN => n15147);
   U19886 : NAND2_X1 port map( A1 => n28154, A2 => n334, ZN => n28153);
   U19895 : NAND2_X2 port map( A1 => n26807, A2 => n21772, ZN => n28156);
   U19904 : NOR2_X1 port map( A1 => n334, A2 => n20323, ZN => n28157);
   U19912 : XOR2_X1 port map( A1 => n4075, A2 => n28158, Z => n4268);
   U19918 : XOR2_X1 port map( A1 => n22556, A2 => n18305, Z => n28158);
   U19927 : INV_X4 port map( I => n1711, ZN => n28225);
   U19929 : NOR2_X1 port map( A1 => n1111, A2 => n5198, ZN => n8462);
   U19933 : INV_X2 port map( I => n12079, ZN => n1111);
   U19962 : NOR3_X2 port map( A1 => n10864, A2 => n10863, A3 => n19690, ZN => 
                           n12079);
   U19965 : NAND2_X1 port map( A1 => n18777, A2 => n7960, ZN => n28161);
   U19967 : AOI21_X2 port map( A1 => n28162, A2 => n17264, B => n24479, ZN => 
                           n17267);
   U19975 : NAND2_X1 port map( A1 => n13187, A2 => n22253, ZN => n28162);
   U19976 : INV_X2 port map( I => n28164, ZN => n21715);
   U19980 : XNOR2_X1 port map( A1 => n9679, A2 => n9682, ZN => n28164);
   U19981 : XOR2_X1 port map( A1 => n8225, A2 => n21911, Z => n5127);
   U19982 : NAND2_X2 port map( A1 => n17494, A2 => n14062, ZN => n13928);
   U19990 : BUF_X4 port map( I => n1637, Z => n28166);
   U20000 : NAND3_X2 port map( A1 => n2449, A2 => n28183, A3 => n2454, ZN => 
                           n26549);
   U20006 : XOR2_X1 port map( A1 => n23779, A2 => n7408, Z => n24625);
   U20008 : AOI21_X1 port map( A1 => n3193, A2 => n16341, B => n16340, ZN => 
                           n15712);
   U20016 : INV_X2 port map( I => n21408, ZN => n21415);
   U20031 : NAND2_X2 port map( A1 => n21362, A2 => n24433, ZN => n21408);
   U20033 : XOR2_X1 port map( A1 => n23779, A2 => n17139, Z => n6746);
   U20035 : INV_X4 port map( I => n25975, ZN => n23779);
   U20038 : AOI22_X2 port map( A1 => n12464, A2 => n16690, B1 => n23277, B2 => 
                           n24182, ZN => n25975);
   U20039 : OR2_X1 port map( A1 => n24286, A2 => n7769, Z => n28503);
   U20041 : XOR2_X1 port map( A1 => n7520, A2 => n28167, Z => n965);
   U20042 : XOR2_X1 port map( A1 => n4995, A2 => n8242, Z => n28167);
   U20046 : BUF_X2 port map( I => n9472, Z => n28168);
   U20051 : INV_X1 port map( I => n28318, ZN => n7215);
   U20057 : XOR2_X1 port map( A1 => n28169, A2 => n884, Z => n5969);
   U20060 : XOR2_X1 port map( A1 => n5542, A2 => n18215, Z => n28169);
   U20064 : NAND2_X2 port map( A1 => n7846, A2 => n7845, ZN => n28276);
   U20070 : AND2_X1 port map( A1 => n13873, A2 => n8467, Z => n4736);
   U20071 : NAND2_X1 port map( A1 => n7420, A2 => n7980, ZN => n28170);
   U20073 : INV_X1 port map( I => n9943, ZN => n8444);
   U20077 : NOR2_X2 port map( A1 => n23923, A2 => n21901, ZN => n28252);
   U20080 : NAND2_X1 port map( A1 => n934, A2 => n9563, ZN => n2322);
   U20087 : INV_X2 port map( I => n24821, ZN => n17393);
   U20093 : NOR2_X2 port map( A1 => n17244, A2 => n25338, ZN => n24821);
   U20097 : AOI22_X2 port map( A1 => n28174, A2 => n28173, B1 => n14664, B2 => 
                           n3009, ZN => n128);
   U20109 : NAND2_X2 port map( A1 => n23642, A2 => n24179, ZN => n28175);
   U20110 : XOR2_X1 port map( A1 => n15360, A2 => n10854, Z => n15359);
   U20134 : NAND3_X1 port map( A1 => n28178, A2 => n28177, A3 => n28176, ZN => 
                           n15034);
   U20140 : NAND2_X1 port map( A1 => n12235, A2 => n20680, ZN => n28177);
   U20151 : INV_X1 port map( I => n20670, ZN => n28178);
   U20152 : OAI22_X2 port map( A1 => n2945, A2 => n24870, B1 => n13726, B2 => 
                           n15448, ZN => n2944);
   U20154 : INV_X1 port map( I => n26096, ZN => n28192);
   U20155 : NAND2_X2 port map( A1 => n1602, A2 => n28179, ZN => n2507);
   U20162 : NOR2_X2 port map( A1 => n24972, A2 => n28180, ZN => n10019);
   U20163 : OAI22_X2 port map( A1 => n16132, A2 => n14150, B1 => n6278, B2 => 
                           n10453, ZN => n16137);
   U20164 : XOR2_X1 port map( A1 => n28181, A2 => n10876, Z => n26049);
   U20172 : XOR2_X1 port map( A1 => n17115, A2 => n12120, Z => n28181);
   U20178 : XOR2_X1 port map( A1 => n4910, A2 => n23173, Z => n28182);
   U20179 : AND2_X2 port map( A1 => n14446, A2 => n23011, Z => n28540);
   U20188 : XOR2_X1 port map( A1 => n15647, A2 => n8486, Z => n2370);
   U20189 : XOR2_X1 port map( A1 => n28185, A2 => n20378, Z => n15453);
   U20196 : XOR2_X1 port map( A1 => n1613, A2 => n20497, Z => n28185);
   U20203 : XOR2_X1 port map( A1 => n17029, A2 => n17136, Z => n8018);
   U20204 : XOR2_X1 port map( A1 => n16806, A2 => n16938, Z => n17136);
   U20205 : OAI22_X2 port map( A1 => n14071, A2 => n796, B1 => n24008, B2 => 
                           n23259, ZN => n9652);
   U20206 : NAND2_X2 port map( A1 => n7158, A2 => n5464, ZN => n24008);
   U20207 : XOR2_X1 port map( A1 => n3598, A2 => n12602, Z => n8857);
   U20208 : XOR2_X1 port map( A1 => n23041, A2 => n22839, Z => n3598);
   U20215 : NOR2_X1 port map( A1 => n281, A2 => n28189, ZN => n2358);
   U20227 : NAND2_X1 port map( A1 => n26482, A2 => n1017, ZN => n28189);
   U20228 : OAI21_X2 port map( A1 => n23171, A2 => n17338, B => n17335, ZN => 
                           n17341);
   U20231 : XOR2_X1 port map( A1 => n19565, A2 => n14608, Z => n19385);
   U20234 : XOR2_X1 port map( A1 => n9904, A2 => n13064, Z => n8114);
   U20236 : XOR2_X1 port map( A1 => n3351, A2 => n4680, Z => n4679);
   U20237 : XOR2_X1 port map( A1 => n28190, A2 => n10880, Z => n11404);
   U20242 : XOR2_X1 port map( A1 => n18059, A2 => n18323, Z => n28190);
   U20243 : NAND3_X2 port map( A1 => n28191, A2 => n17297, A3 => n17298, ZN => 
                           n3326);
   U20253 : NOR2_X2 port map( A1 => n27787, A2 => n26098, ZN => n28193);
   U20278 : NOR2_X2 port map( A1 => n20932, A2 => n20938, ZN => n20885);
   U20283 : NAND2_X2 port map( A1 => n6405, A2 => n24186, ZN => n6052);
   U20287 : OAI22_X2 port map( A1 => n15733, A2 => n15732, B1 => n26710, B2 => 
                           n13104, ZN => n20193);
   U20290 : XOR2_X1 port map( A1 => n3753, A2 => n3754, Z => n10105);
   U20292 : XOR2_X1 port map( A1 => n13695, A2 => n19359, Z => n19083);
   U20299 : NAND2_X1 port map( A1 => n28236, A2 => n19571, ZN => n4228);
   U20302 : BUF_X2 port map( I => n28302, Z => n28194);
   U20305 : NAND2_X2 port map( A1 => n6283, A2 => n28195, ZN => n20449);
   U20307 : XOR2_X1 port map( A1 => n18240, A2 => n28196, Z => n26519);
   U20308 : XOR2_X1 port map( A1 => n11787, A2 => n4204, Z => n28196);
   U20313 : INV_X1 port map( I => n23214, ZN => n17174);
   U20315 : NAND2_X1 port map( A1 => n17173, A2 => n1565, ZN => n23214);
   U20330 : INV_X1 port map( I => n15004, ZN => n28197);
   U20339 : NAND2_X1 port map( A1 => n11318, A2 => n28213, ZN => n28212);
   U20352 : NAND3_X1 port map( A1 => n28215, A2 => n27751, A3 => n28212, ZN => 
                           n28211);
   U20357 : INV_X4 port map( I => n9485, ZN => n5584);
   U20358 : NAND2_X2 port map( A1 => n17845, A2 => n17992, ZN => n17991);
   U20361 : OAI21_X2 port map( A1 => n28203, A2 => n28202, B => n18595, ZN => 
                           n19189);
   U20362 : NOR2_X2 port map( A1 => n14154, A2 => n18592, ZN => n28203);
   U20371 : XOR2_X1 port map( A1 => n1389, A2 => n28204, Z => n645);
   U20372 : XOR2_X1 port map( A1 => n2978, A2 => n22077, Z => n28204);
   U20373 : NAND2_X1 port map( A1 => n23154, A2 => n21646, ZN => n23069);
   U20381 : NAND2_X2 port map( A1 => n9464, A2 => n22814, ZN => n18621);
   U20382 : XOR2_X1 port map( A1 => n28206, A2 => n14432, Z => Ciphertext(87));
   U20385 : NAND2_X2 port map( A1 => n27344, A2 => n23255, ZN => n13593);
   U20386 : NAND2_X2 port map( A1 => n7014, A2 => n7015, ZN => n14071);
   U20387 : XOR2_X1 port map( A1 => n9656, A2 => n19367, Z => n9257);
   U20389 : XOR2_X1 port map( A1 => n19540, A2 => n19299, Z => n19367);
   U20393 : NAND2_X2 port map( A1 => n7372, A2 => n23239, ZN => n12527);
   U20397 : BUF_X2 port map( I => n7611, Z => n28207);
   U20398 : XOR2_X1 port map( A1 => n28208, A2 => n28460, Z => n25080);
   U20400 : AND2_X1 port map( A1 => n24089, A2 => n26254, Z => n23256);
   U20401 : XOR2_X1 port map( A1 => n22169, A2 => n14608, Z => n26177);
   U20402 : OAI21_X2 port map( A1 => n25234, A2 => n25235, B => n12035, ZN => 
                           n28209);
   U20404 : NOR3_X1 port map( A1 => n13786, A2 => n16516, A3 => n3470, ZN => 
                           n23070);
   U20417 : NAND2_X2 port map( A1 => n1403, A2 => n3769, ZN => n3470);
   U20424 : XOR2_X1 port map( A1 => n18073, A2 => n28210, Z => n28310);
   U20427 : INV_X2 port map( I => n18184, ZN => n28210);
   U20438 : XOR2_X1 port map( A1 => n15237, A2 => n18072, Z => n18184);
   U20448 : NAND2_X2 port map( A1 => n7968, A2 => n23166, ZN => n2391);
   U20449 : INV_X2 port map( I => n20842, ZN => n28214);
   U20450 : OR2_X1 port map( A1 => n11318, A2 => n8760, Z => n28215);
   U20459 : OR2_X1 port map( A1 => n26317, A2 => n13372, Z => n11241);
   U20466 : XOR2_X1 port map( A1 => n23130, A2 => n28217, Z => n24788);
   U20468 : XNOR2_X1 port map( A1 => n20550, A2 => n5949, ZN => n11672);
   U20478 : NAND2_X2 port map( A1 => n11773, A2 => n17277, ZN => n14278);
   U20479 : INV_X2 port map( I => n14451, ZN => n16657);
   U20483 : NAND3_X2 port map( A1 => n14561, A2 => n5178, A3 => n5179, ZN => 
                           n14451);
   U20487 : AOI22_X1 port map( A1 => n25646, A2 => n15580, B1 => n20653, B2 => 
                           n4766, ZN => n28223);
   U20511 : XOR2_X1 port map( A1 => n28219, A2 => n1278, Z => Ciphertext(146));
   U20519 : XOR2_X1 port map( A1 => n28220, A2 => n3899, Z => n360);
   U20521 : XOR2_X1 port map( A1 => n3898, A2 => n3897, Z => n28220);
   U20530 : XOR2_X1 port map( A1 => n3667, A2 => n16763, Z => n25622);
   U20535 : AOI21_X2 port map( A1 => n17772, A2 => n22307, B => n28221, ZN => 
                           n18270);
   U20544 : OAI22_X2 port map( A1 => n3910, A2 => n28322, B1 => n22307, B2 => 
                           n6038, ZN => n28221);
   U20547 : NAND2_X2 port map( A1 => n21534, A2 => n12625, ZN => n30);
   U20556 : XOR2_X1 port map( A1 => n23865, A2 => n473, Z => n3389);
   U20562 : NAND2_X2 port map( A1 => n4735, A2 => n13371, ZN => n4624);
   U20563 : XOR2_X1 port map( A1 => n28223, A2 => n13678, Z => Ciphertext(14));
   U20577 : XOR2_X1 port map( A1 => n2065, A2 => n25485, Z => n25338);
   U20580 : XOR2_X1 port map( A1 => n14733, A2 => n13284, Z => n2065);
   U20582 : XOR2_X1 port map( A1 => n21260, A2 => n26238, Z => n1734);
   U20585 : INV_X2 port map( I => n20078, ZN => n12143);
   U20588 : NAND2_X2 port map( A1 => n28225, A2 => n28224, ZN => n24337);
   U20596 : NOR2_X2 port map( A1 => n6727, A2 => n6728, ZN => n20850);
   U20619 : AOI21_X2 port map( A1 => n20809, A2 => n1726, B => n20899, ZN => 
                           n6727);
   U20623 : XOR2_X1 port map( A1 => n28226, A2 => n1289, Z => Ciphertext(187));
   U20627 : NAND2_X1 port map( A1 => n4327, A2 => n21740, ZN => n4326);
   U20629 : OAI21_X2 port map( A1 => n5252, A2 => n22212, B => n5251, ZN => 
                           n28228);
   U20631 : XOR2_X1 port map( A1 => n13858, A2 => n8111, Z => n8003);
   U20638 : XOR2_X1 port map( A1 => n18144, A2 => n1197, Z => n8111);
   U20643 : XOR2_X1 port map( A1 => n20527, A2 => n27373, Z => n20012);
   U20648 : NOR3_X1 port map( A1 => n18953, A2 => n18426, A3 => n22391, ZN => 
                           n24425);
   U20660 : NAND2_X2 port map( A1 => n21061, A2 => n21059, ZN => n20971);
   U20662 : NOR2_X1 port map( A1 => n17408, A2 => n6293, ZN => n17206);
   U20667 : INV_X2 port map( I => n7651, ZN => n17408);
   U20669 : XOR2_X1 port map( A1 => n25674, A2 => n620, Z => n7651);
   U20673 : AOI21_X2 port map( A1 => n28229, A2 => n18968, B => n1159, ZN => 
                           n25861);
   U20674 : NAND2_X2 port map( A1 => n4735, A2 => n19134, ZN => n28229);
   U20682 : XOR2_X1 port map( A1 => n28230, A2 => n14622, Z => Ciphertext(174))
                           ;
   U20701 : NAND3_X1 port map( A1 => n10081, A2 => n7498, A3 => n10985, ZN => 
                           n17005);
   U20702 : AND2_X1 port map( A1 => n11497, A2 => n6910, Z => n11498);
   U20706 : XOR2_X1 port map( A1 => n14601, A2 => n5682, Z => n4107);
   U20709 : NAND3_X1 port map( A1 => n13973, A2 => n13974, A3 => n7944, ZN => 
                           n13976);
   U20718 : OAI21_X1 port map( A1 => n10937, A2 => n674, B => n1129, ZN => 
                           n1806);
   U20731 : XOR2_X1 port map( A1 => n25631, A2 => n28232, Z => n5972);
   U20737 : NAND2_X1 port map( A1 => n4238, A2 => n4236, ZN => n28232);
   U20742 : XOR2_X1 port map( A1 => n6572, A2 => n5610, Z => n25380);
   U20744 : OAI22_X2 port map( A1 => n25538, A2 => n21513, B1 => n21511, B2 => 
                           n21512, ZN => n12625);
   U20745 : NAND2_X2 port map( A1 => n25059, A2 => n15128, ZN => n16768);
   U20747 : OAI21_X2 port map( A1 => n8914, A2 => n23931, B => n8913, ZN => 
                           n8912);
   U20750 : INV_X2 port map( I => n28380, ZN => n28548);
   U20756 : BUF_X2 port map( I => n25856, Z => n28234);
   U20758 : OAI21_X2 port map( A1 => n12649, A2 => n21593, B => n28235, ZN => 
                           n9611);
   U20766 : AOI21_X2 port map( A1 => n3096, A2 => n21592, B => n21591, ZN => 
                           n28235);
   U20770 : NAND2_X1 port map( A1 => n19572, A2 => n19573, ZN => n28236);
   U20774 : MUX2_X1 port map( I0 => n20847, I1 => n25360, S => n20850, Z => 
                           n20830);
   U20778 : NAND2_X2 port map( A1 => n5974, A2 => n9285, ZN => n6435);
   U20780 : INV_X2 port map( I => n28238, ZN => n28552);
   U20784 : NAND2_X2 port map( A1 => n6496, A2 => n6495, ZN => n9534);
   U20787 : XOR2_X1 port map( A1 => n4025, A2 => n503, Z => n4123);
   U20791 : INV_X2 port map( I => n26006, ZN => n846);
   U20799 : NOR2_X2 port map( A1 => n22537, A2 => n19165, ZN => n28241);
   U20800 : XOR2_X1 port map( A1 => n6157, A2 => n10088, Z => n28243);
   U20808 : INV_X1 port map( I => n14166, ZN => n19461);
   U20822 : XOR2_X1 port map( A1 => n19306, A2 => n19365, Z => n14166);
   U20825 : NAND2_X2 port map( A1 => n14835, A2 => n14833, ZN => n25332);
   U20828 : AOI22_X2 port map( A1 => n25245, A2 => n14837, B1 => n19108, B2 => 
                           n9268, ZN => n14835);
   U20835 : XOR2_X1 port map( A1 => n6455, A2 => n25648, Z => n17261);
   U20842 : XOR2_X1 port map( A1 => n9338, A2 => n19530, Z => n1743);
   U20858 : NAND2_X2 port map( A1 => n13778, A2 => n15054, ZN => n9338);
   U20863 : NOR3_X2 port map( A1 => n28244, A2 => n17208, A3 => n748, ZN => 
                           n17210);
   U20864 : XOR2_X1 port map( A1 => n16744, A2 => n4958, Z => n4957);
   U20865 : NOR3_X1 port map( A1 => n21528, A2 => n21531, A3 => n21529, ZN => 
                           n21522);
   U20879 : XOR2_X1 port map( A1 => n17083, A2 => n6137, Z => n3639);
   U20888 : XOR2_X1 port map( A1 => n8819, A2 => n4876, Z => n17083);
   U20903 : OR2_X1 port map( A1 => n540, A2 => n17343, Z => n3360);
   U20913 : AOI21_X2 port map( A1 => n1383, A2 => n12752, B => n28245, ZN => 
                           n2359);
   U20920 : OAI22_X2 port map( A1 => n12374, A2 => n21780, B1 => n1383, B2 => 
                           n12373, ZN => n28245);
   U20921 : NAND2_X2 port map( A1 => n13593, A2 => n13592, ZN => n14294);
   U20931 : AOI22_X2 port map( A1 => n5666, A2 => n11702, B1 => n16668, B2 => 
                           n16488, ZN => n13592);
   U20934 : NAND2_X1 port map( A1 => n28246, A2 => n74, ZN => n22128);
   U20945 : NAND2_X1 port map( A1 => n18670, A2 => n25770, ZN => n28246);
   U20946 : BUF_X2 port map( I => n25214, Z => n28247);
   U20949 : OAI21_X2 port map( A1 => n28118, A2 => n21779, B => n9804, ZN => 
                           n1428);
   U20953 : NAND2_X2 port map( A1 => n28249, A2 => n11198, ZN => n23679);
   U20954 : NAND2_X2 port map( A1 => n28250, A2 => n3059, ZN => n28249);
   U20964 : NAND2_X2 port map( A1 => n21623, A2 => n21624, ZN => n3059);
   U20969 : INV_X2 port map( I => n21628, ZN => n28250);
   U20972 : OAI21_X2 port map( A1 => n448, A2 => n13969, B => n28251, ZN => 
                           n13376);
   U20973 : NOR2_X2 port map( A1 => n5837, A2 => n5836, ZN => n10602);
   U20977 : XOR2_X1 port map( A1 => n18132, A2 => n18236, Z => n18274);
   U20980 : OAI22_X2 port map( A1 => n22630, A2 => n17952, B1 => n5765, B2 => 
                           n762, ZN => n18132);
   U20984 : XOR2_X1 port map( A1 => n7248, A2 => n14645, Z => n28253);
   U20987 : XOR2_X1 port map( A1 => n18335, A2 => n21893, Z => n5275);
   U20989 : OAI22_X2 port map( A1 => n20818, A2 => n14113, B1 => n732, B2 => 
                           n7518, ZN => n8470);
   U20990 : NAND2_X2 port map( A1 => n28254, A2 => n19771, ZN => n20323);
   U20992 : NAND2_X1 port map( A1 => n11237, A2 => n11235, ZN => n28254);
   U21000 : XOR2_X1 port map( A1 => n20535, A2 => n20344, Z => n23585);
   U21001 : NAND2_X2 port map( A1 => n4163, A2 => n28256, ZN => n16822);
   U21014 : NAND3_X2 port map( A1 => n4169, A2 => n4168, A3 => n4162, ZN => 
                           n28256);
   U21015 : BUF_X2 port map( I => n16461, Z => n28257);
   U21021 : XOR2_X1 port map( A1 => n28258, A2 => n4049, Z => n24728);
   U21022 : XOR2_X1 port map( A1 => n16764, A2 => n28259, Z => n28258);
   U21028 : INV_X2 port map( I => n24193, ZN => n28259);
   U21029 : NOR2_X2 port map( A1 => n17236, A2 => n17235, ZN => n28302);
   U21031 : XOR2_X1 port map( A1 => n16881, A2 => n3477, Z => n25293);
   U21040 : NAND2_X2 port map( A1 => n14246, A2 => n10531, ZN => n16881);
   U21046 : OR2_X1 port map( A1 => n12413, A2 => n21578, Z => n22227);
   U21070 : XOR2_X1 port map( A1 => n6138, A2 => n23294, Z => n15432);
   U21075 : NAND2_X2 port map( A1 => n7795, A2 => n6776, ZN => n20523);
   U21089 : XOR2_X1 port map( A1 => n28261, A2 => n14624, Z => Ciphertext(44));
   U21099 : NAND2_X1 port map( A1 => n20830, A2 => n20842, ZN => n28262);
   U21103 : NAND2_X2 port map( A1 => n23399, A2 => n27715, ZN => n18737);
   U21107 : OAI22_X2 port map( A1 => n15962, A2 => n4841, B1 => n15961, B2 => 
                           n8925, ZN => n25875);
   U21113 : NOR2_X2 port map( A1 => n25067, A2 => n25066, ZN => n24864);
   U21115 : XOR2_X1 port map( A1 => n19555, A2 => n10213, Z => n8821);
   U21116 : AND2_X1 port map( A1 => n16132, A2 => n15923, Z => n15830);
   U21117 : BUF_X2 port map( I => n18314, Z => n28265);
   U21118 : NAND2_X2 port map( A1 => n2592, A2 => n13055, ZN => n4486);
   U21120 : NOR2_X2 port map( A1 => n5471, A2 => n28266, ZN => n24283);
   U21129 : NAND2_X2 port map( A1 => n16466, A2 => n3479, ZN => n28356);
   U21134 : NAND2_X2 port map( A1 => n11829, A2 => n11828, ZN => n16466);
   U21137 : XOR2_X1 port map( A1 => n2410, A2 => n28267, Z => n13048);
   U21138 : XOR2_X1 port map( A1 => n16922, A2 => n2409, Z => n28267);
   U21143 : OAI21_X2 port map( A1 => n4081, A2 => n20936, B => n20939, ZN => 
                           n4413);
   U21153 : XOR2_X1 port map( A1 => n28273, A2 => n21308, Z => n4384);
   U21154 : AND2_X1 port map( A1 => n20217, A2 => n10810, Z => n23222);
   U21155 : NAND2_X2 port map( A1 => n5182, A2 => n5761, ZN => n7044);
   U21156 : OAI21_X2 port map( A1 => n14261, A2 => n6716, B => n3505, ZN => 
                           n20543);
   U21157 : XOR2_X1 port map( A1 => n20581, A2 => n21190, Z => n21428);
   U21159 : NOR2_X2 port map( A1 => n5014, A2 => n20118, ZN => n20581);
   U21162 : NAND2_X2 port map( A1 => n4279, A2 => n28275, ZN => n6932);
   U21168 : BUF_X2 port map( I => n23253, Z => n28277);
   U21170 : NAND2_X2 port map( A1 => n28279, A2 => n13813, ZN => n11733);
   U21171 : NAND2_X1 port map( A1 => n15978, A2 => n13256, ZN => n28279);
   U21172 : XOR2_X1 port map( A1 => n21191, A2 => n20450, Z => n20485);
   U21177 : OAI22_X2 port map( A1 => n19971, A2 => n25431, B1 => n3802, B2 => 
                           n20125, ZN => n20450);
   U21182 : AOI21_X2 port map( A1 => n28280, A2 => n19988, B => n24037, ZN => 
                           n13330);
   U21184 : AND2_X1 port map( A1 => n19987, A2 => n809, Z => n28280);
   U21186 : INV_X2 port map( I => n21737, ZN => n1065);
   U21187 : NAND2_X2 port map( A1 => n21718, A2 => n9976, ZN => n21737);
   U21192 : XOR2_X1 port map( A1 => n19537, A2 => n28281, Z => n10201);
   U21193 : XOR2_X1 port map( A1 => n5560, A2 => n1359, Z => n28281);
   U21194 : AND2_X1 port map( A1 => n5445, A2 => n22554, Z => n9094);
   U21199 : NAND2_X2 port map( A1 => n14810, A2 => n7636, ZN => n20580);
   U21206 : OAI21_X2 port map( A1 => n28282, A2 => n26033, B => n3091, ZN => 
                           n9632);
   U21210 : NOR2_X2 port map( A1 => n17166, A2 => n24159, ZN => n28282);
   U21212 : XOR2_X1 port map( A1 => n3313, A2 => n28283, Z => n9070);
   U21217 : XOR2_X1 port map( A1 => n19194, A2 => n19560, Z => n19317);
   U21222 : OAI22_X1 port map( A1 => n23976, A2 => n13473, B1 => n13444, B2 => 
                           n11837, ZN => n4058);
   U21226 : OAI21_X2 port map( A1 => n28286, A2 => n11612, B => n22920, ZN => 
                           n11611);
   U21228 : NOR2_X2 port map( A1 => n19068, A2 => n21776, ZN => n28286);
   U21239 : INV_X4 port map( I => n13942, ZN => n19006);
   U21240 : NAND2_X2 port map( A1 => n13940, A2 => n13939, ZN => n13942);
   U21249 : XOR2_X1 port map( A1 => n28289, A2 => n10387, Z => n25120);
   U21259 : XOR2_X1 port map( A1 => n24077, A2 => n27104, Z => n28289);
   U21266 : NAND2_X2 port map( A1 => n28290, A2 => n6979, ZN => n5317);
   U21278 : NOR2_X2 port map( A1 => n22998, A2 => n13480, ZN => n28290);
   U21281 : XOR2_X1 port map( A1 => n21300, A2 => n28291, Z => n7638);
   U21282 : XOR2_X1 port map( A1 => n8581, A2 => n20725, Z => n28291);
   U21289 : BUF_X2 port map( I => n26058, Z => n28292);
   U21293 : NAND2_X2 port map( A1 => n5700, A2 => n5701, ZN => n5698);
   U21296 : XOR2_X1 port map( A1 => n18099, A2 => n18171, Z => n18336);
   U21311 : XOR2_X1 port map( A1 => n18270, A2 => n22886, Z => n28294);
   U21312 : NAND3_X1 port map( A1 => n26097, A2 => n10164, A3 => n27647, ZN => 
                           n6931);
   U21314 : XOR2_X1 port map( A1 => n7423, A2 => n15073, Z => n7422);
   U21327 : OR2_X2 port map( A1 => n16193, A2 => n14893, Z => n11660);
   U21332 : XOR2_X1 port map( A1 => n16627, A2 => n28296, Z => n22159);
   U21335 : XOR2_X1 port map( A1 => n16975, A2 => n16616, Z => n28296);
   U21344 : AOI22_X2 port map( A1 => n25406, A2 => n6332, B1 => n3286, B2 => 
                           n7656, ZN => n13235);
   U21363 : NAND3_X1 port map( A1 => n21473, A2 => n21483, A3 => n11622, ZN => 
                           n21470);
   U21366 : INV_X2 port map( I => n28301, ZN => n679);
   U21371 : XOR2_X1 port map( A1 => n26405, A2 => n26406, Z => n3417);
   U21384 : NAND3_X2 port map( A1 => n18389, A2 => n14207, A3 => n5192, ZN => 
                           n18390);
   U21386 : INV_X1 port map( I => n21695, ZN => n28304);
   U21400 : XOR2_X1 port map( A1 => Plaintext(191), A2 => Key(191), Z => n562);
   U21401 : INV_X1 port map( I => n16453, ZN => n28364);
   U21405 : NAND2_X2 port map( A1 => n6469, A2 => n28307, ZN => n6598);
   U21412 : XOR2_X1 port map( A1 => n18291, A2 => n6015, Z => n5823);
   U21420 : XOR2_X1 port map( A1 => n28310, A2 => n316, Z => n9411);
   U21421 : AOI21_X1 port map( A1 => n12517, A2 => n21608, B => n940, ZN => 
                           n21610);
   U21426 : NOR3_X2 port map( A1 => n2309, A2 => n8552, A3 => n8553, ZN => 
                           n19071);
   U21427 : NAND2_X2 port map( A1 => n7468, A2 => n2346, ZN => n8557);
   U21432 : OAI21_X2 port map( A1 => n24695, A2 => n9287, B => n2960, ZN => 
                           n9286);
   U21434 : XOR2_X1 port map( A1 => n20579, A2 => n13892, Z => n28312);
   U21435 : XOR2_X1 port map( A1 => n21198, A2 => n27418, Z => n20456);
   U21437 : XOR2_X1 port map( A1 => n9369, A2 => n18136, Z => n18140);
   U21441 : BUF_X2 port map( I => n20180, Z => n28314);
   U21447 : NAND3_X2 port map( A1 => n14889, A2 => n28317, A3 => n28316, ZN => 
                           n21371);
   U21449 : NAND2_X2 port map( A1 => n26459, A2 => n6470, ZN => n28317);
   U21452 : OAI21_X2 port map( A1 => n11834, A2 => n1780, B => n12899, ZN => 
                           n2772);
   U21453 : XOR2_X1 port map( A1 => n28318, A2 => n19419, Z => n5036);
   U21454 : OAI22_X2 port map( A1 => n5108, A2 => n5109, B1 => n5110, B2 => 
                           n9952, ZN => n19419);
   U21455 : NAND2_X2 port map( A1 => n13121, A2 => n19870, ZN => n19570);
   U21465 : OAI22_X2 port map( A1 => n25864, A2 => n2727, B1 => n18548, B2 => 
                           n24572, ZN => n9873);
   U21468 : NAND2_X2 port map( A1 => n20505, A2 => n28319, ZN => n20618);
   U21476 : AOI22_X2 port map( A1 => n78, A2 => n24327, B1 => n20733, B2 => 
                           n2536, ZN => n28319);
   U21482 : XOR2_X1 port map( A1 => n5742, A2 => n20381, Z => n28320);
   U21485 : XOR2_X1 port map( A1 => n28321, A2 => n539, Z => n17221);
   U21500 : XOR2_X1 port map( A1 => n12454, A2 => n17087, Z => n28321);
   U21510 : XOR2_X1 port map( A1 => n5127, A2 => n5129, Z => n22568);
   U21523 : XOR2_X1 port map( A1 => n5772, A2 => n28323, Z => n21253);
   U21525 : NOR2_X2 port map( A1 => n16063, A2 => n28152, ZN => n28324);
   U21528 : XOR2_X1 port map( A1 => n4631, A2 => n8964, Z => n8963);
   U21530 : BUF_X2 port map( I => n5921, Z => n28325);
   U21531 : NAND2_X2 port map( A1 => n28390, A2 => n11818, ZN => n28328);
   U21535 : NAND3_X1 port map( A1 => n6618, A2 => n28081, A3 => n6619, ZN => 
                           n28329);
   U21538 : XOR2_X1 port map( A1 => n23074, A2 => n28330, Z => n9332);
   U21542 : XOR2_X1 port map( A1 => n18120, A2 => n2604, Z => n28330);
   U21546 : AOI22_X2 port map( A1 => n28331, A2 => n19981, B1 => n3460, B2 => 
                           n3461, ZN => n25186);
   U21553 : NOR2_X2 port map( A1 => n4537, A2 => n4311, ZN => n28332);
   U21554 : XOR2_X1 port map( A1 => n28334, A2 => n20538, Z => n7077);
   U21559 : NAND2_X2 port map( A1 => n19984, A2 => n14258, ZN => n20538);
   U21563 : OAI21_X2 port map( A1 => n12676, A2 => n17844, B => n28335, ZN => 
                           n8782);
   U21565 : OAI21_X2 port map( A1 => n18543, A2 => n11873, B => n26321, ZN => 
                           n18376);
   U21569 : XOR2_X1 port map( A1 => n28336, A2 => n6751, Z => n8011);
   U21574 : XOR2_X1 port map( A1 => n7076, A2 => n15308, Z => n15624);
   U21577 : XOR2_X1 port map( A1 => n19288, A2 => n28337, Z => n9013);
   U21582 : XOR2_X1 port map( A1 => n25794, A2 => n22793, Z => n28337);
   U21583 : XOR2_X1 port map( A1 => n16768, A2 => n15256, Z => n16583);
   U21592 : XOR2_X1 port map( A1 => n20527, A2 => n27391, Z => n8259);
   U21595 : OAI21_X2 port map( A1 => n7094, A2 => n6005, B => n6004, ZN => 
                           n20527);
   U21597 : NAND2_X2 port map( A1 => n17644, A2 => n17643, ZN => n3701);
   U21598 : NAND2_X1 port map( A1 => n18654, A2 => n24568, ZN => n8357);
   U21605 : XOR2_X1 port map( A1 => n8361, A2 => n7285, Z => n24568);
   U21606 : NAND2_X2 port map( A1 => n5452, A2 => n28340, ZN => n13994);
   U21609 : NAND3_X1 port map( A1 => n21734, A2 => n26647, A3 => n9458, ZN => 
                           n4327);
   U21610 : XOR2_X1 port map( A1 => n20373, A2 => n25502, Z => n21547);
   U21619 : XOR2_X1 port map( A1 => n19463, A2 => n28341, Z => n9044);
   U21620 : XOR2_X1 port map( A1 => n11969, A2 => n19378, Z => n28341);
   U21624 : XNOR2_X1 port map( A1 => n12681, A2 => n12300, ZN => n28344);
   U21629 : XOR2_X1 port map( A1 => n26575, A2 => n28342, Z => n21895);
   U21632 : INV_X2 port map( I => n13048, ZN => n17185);
   U21634 : XOR2_X1 port map( A1 => n11275, A2 => n3372, Z => n10088);
   U21636 : NAND2_X2 port map( A1 => n25432, A2 => n12661, ZN => n11275);
   U21643 : AND2_X1 port map( A1 => n14855, A2 => n14854, Z => n3081);
   U21650 : NOR2_X2 port map( A1 => n24727, A2 => n3553, ZN => n16680);
   U21656 : NAND2_X1 port map( A1 => n21009, A2 => n12613, ZN => n28343);
   U21657 : NAND3_X2 port map( A1 => n3609, A2 => n1150, A3 => n5702, ZN => 
                           n25166);
   U21659 : INV_X4 port map( I => n26491, ZN => n11937);
   U21661 : NAND2_X2 port map( A1 => n22986, A2 => n28349, ZN => n26491);
   U21665 : INV_X2 port map( I => n421, ZN => n15227);
   U21666 : NAND2_X1 port map( A1 => n28345, A2 => n4706, ZN => n4704);
   U21667 : XOR2_X1 port map( A1 => n23502, A2 => n16993, Z => n11768);
   U21669 : AOI21_X2 port map( A1 => n14259, A2 => n16614, B => n145, ZN => 
                           n15013);
   U21670 : XOR2_X1 port map( A1 => n28348, A2 => n25227, Z => n1551);
   U21674 : XOR2_X1 port map( A1 => n18300, A2 => n594, Z => n28348);
   U21676 : NOR2_X2 port map( A1 => n24562, A2 => n802, ZN => n6037);
   U21680 : NAND2_X2 port map( A1 => n28469, A2 => n28351, ZN => n9047);
   U21683 : AOI22_X2 port map( A1 => n8217, A2 => n9057, B1 => n21671, B2 => 
                           n22747, ZN => n28351);
   U21693 : NOR2_X2 port map( A1 => n22506, A2 => n9987, ZN => n7405);
   U21694 : XOR2_X1 port map( A1 => n9791, A2 => n21218, Z => n5067);
   U21695 : AOI22_X2 port map( A1 => n18100, A2 => n1202, B1 => n25192, B2 => 
                           n11661, ZN => n5126);
   U21696 : NOR2_X2 port map( A1 => n27714, A2 => n22396, ZN => n18100);
   U21699 : NAND2_X2 port map( A1 => n28352, A2 => n16212, ZN => n8181);
   U21702 : NAND3_X2 port map( A1 => n23609, A2 => n23610, A3 => n12025, ZN => 
                           n28352);
   U21704 : XOR2_X1 port map( A1 => n16913, A2 => n24740, Z => n17081);
   U21707 : OAI21_X2 port map( A1 => n16463, A2 => n26594, B => n12608, ZN => 
                           n16913);
   U21708 : XOR2_X1 port map( A1 => n13906, A2 => n1975, Z => n19497);
   U21709 : NAND2_X2 port map( A1 => n28354, A2 => n15430, ZN => n15431);
   U21710 : NOR2_X1 port map( A1 => n13734, A2 => n13735, ZN => n28354);
   U21714 : XOR2_X1 port map( A1 => n24903, A2 => n17017, Z => n1998);
   U21718 : INV_X2 port map( I => n28357, ZN => n464);
   U21719 : INV_X2 port map( I => n19873, ZN => n28357);
   U21720 : NOR2_X2 port map( A1 => n14565, A2 => n8754, ZN => n19631);
   U21723 : NAND2_X2 port map( A1 => n159, A2 => n4409, ZN => n19392);
   U21726 : NAND3_X2 port map( A1 => n7939, A2 => n7938, A3 => n7937, ZN => 
                           n18793);
   U21727 : XOR2_X1 port map( A1 => n8503, A2 => n8504, Z => n24251);
   U21728 : NAND3_X2 port map( A1 => n7952, A2 => n28487, A3 => n18770, ZN => 
                           n18771);
   U21729 : XOR2_X1 port map( A1 => n12146, A2 => n28359, Z => n23279);
   U21736 : XOR2_X1 port map( A1 => n4618, A2 => n28360, Z => n28359);
   U21739 : INV_X1 port map( I => n20851, ZN => n28360);
   U21742 : NAND3_X2 port map( A1 => n28361, A2 => n4577, A3 => n24368, ZN => 
                           n25290);
   U21744 : NAND2_X2 port map( A1 => n13568, A2 => n27168, ZN => n28361);
   U21745 : INV_X2 port map( I => n792, ZN => n17078);
   U21754 : XOR2_X1 port map( A1 => n5499, A2 => n792, Z => n9399);
   U21757 : NOR2_X2 port map( A1 => n28364, A2 => n28363, ZN => n792);
   U21762 : OR2_X1 port map( A1 => n7839, A2 => n12729, Z => n28365);
   U21763 : NAND2_X2 port map( A1 => n23772, A2 => n5990, ZN => n6013);
   U21766 : BUF_X2 port map( I => n17436, Z => n28367);
   U21769 : OAI21_X2 port map( A1 => n9391, A2 => n16399, B => n9829, ZN => 
                           n28368);
   U21776 : BUF_X2 port map( I => n16483, Z => n28369);
   U21777 : XOR2_X1 port map( A1 => n26012, A2 => n4689, Z => n4688);
   U21778 : BUF_X2 port map( I => n12192, Z => n28373);
   U21781 : INV_X4 port map( I => n19720, ZN => n28378);
   U21782 : NAND2_X2 port map( A1 => n4006, A2 => n22052, ZN => n13119);
   U21784 : NAND2_X1 port map( A1 => n22016, A2 => n22017, ZN => n22015);
   U21795 : INV_X2 port map( I => n12947, ZN => n13422);
   U21796 : NAND3_X2 port map( A1 => n10019, A2 => n10023, A3 => n10024, ZN => 
                           n12947);
   U21803 : NAND2_X1 port map( A1 => n19845, A2 => n28375, ZN => n14660);
   U21804 : XOR2_X1 port map( A1 => n11277, A2 => n7301, Z => n15004);
   U21805 : AOI22_X2 port map( A1 => n11528, A2 => n11660, B1 => n11940, B2 => 
                           n16286, ZN => n16493);
   U21807 : XOR2_X1 port map( A1 => n23849, A2 => n3707, Z => n12142);
   U21811 : NOR2_X2 port map( A1 => n2717, A2 => n25860, ZN => n23849);
   U21817 : XOR2_X1 port map( A1 => n13370, A2 => n18266, Z => n5130);
   U21820 : NOR2_X2 port map( A1 => n24524, A2 => n2647, ZN => n28380);
   U21826 : NAND2_X1 port map( A1 => n28384, A2 => n28383, ZN => n28382);
   U21836 : INV_X1 port map( I => n11874, ZN => n28383);
   U21837 : NOR2_X1 port map( A1 => n13716, A2 => n20317, ZN => n28385);
   U21850 : OAI21_X1 port map( A1 => n8860, A2 => n10388, B => n28386, ZN => 
                           n2432);
   U21851 : XNOR2_X1 port map( A1 => n18319, A2 => n18318, ZN => n28445);
   U21855 : NAND2_X1 port map( A1 => n7960, A2 => n18776, ZN => n26482);
   U21856 : XOR2_X1 port map( A1 => n13714, A2 => n13710, Z => n26354);
   U21858 : NAND2_X2 port map( A1 => n26163, A2 => n12886, ZN => n12885);
   U21860 : AOI21_X2 port map( A1 => n10871, A2 => n17885, B => n23923, ZN => 
                           n17889);
   U21862 : XOR2_X1 port map( A1 => n28387, A2 => n14652, Z => Ciphertext(45));
   U21866 : NAND2_X1 port map( A1 => n22391, A2 => n6089, ZN => n9233);
   U21867 : XOR2_X1 port map( A1 => n1539, A2 => n19496, Z => n28388);
   U21869 : NAND2_X2 port map( A1 => n1780, A2 => n11579, ZN => n28390);
   U21870 : NAND2_X1 port map( A1 => n17270, A2 => n17271, ZN => n28392);
   U21871 : OAI21_X2 port map( A1 => n24980, A2 => n24981, B => n12438, ZN => 
                           n28394);
   U21875 : NOR2_X2 port map( A1 => n25701, A2 => n28395, ZN => n16538);
   U21879 : OAI22_X2 port map( A1 => n16291, A2 => n16292, B1 => n16290, B2 => 
                           n12678, ZN => n28395);
   U21883 : INV_X2 port map( I => n28396, ZN => n8223);
   U21885 : OR3_X1 port map( A1 => n7650, A2 => n15784, A3 => n7649, Z => 
                           n28396);
   U21888 : INV_X1 port map( I => n21228, ZN => n12430);
   U21889 : XOR2_X1 port map( A1 => n10075, A2 => n28397, Z => n7437);
   U21890 : XOR2_X1 port map( A1 => n16853, A2 => n16883, Z => n28397);
   U21892 : NAND2_X2 port map( A1 => n16314, A2 => n24872, ZN => n16242);
   U21893 : NAND2_X1 port map( A1 => n11961, A2 => n11048, ZN => n26229);
   U21896 : NAND2_X2 port map( A1 => n9731, A2 => n26653, ZN => n11961);
   U21897 : NAND2_X2 port map( A1 => n87, A2 => n9945, ZN => n4397);
   U21898 : NAND2_X2 port map( A1 => n18674, A2 => n18759, ZN => n5885);
   U21899 : NAND2_X2 port map( A1 => n25107, A2 => n12638, ZN => n17897);
   U21904 : XOR2_X1 port map( A1 => n21984, A2 => n21985, Z => n17983);
   U21907 : BUF_X2 port map( I => n15478, Z => n28402);
   U21908 : AND2_X2 port map( A1 => n13522, A2 => n3212, Z => n21759);
   U21914 : INV_X1 port map( I => n28496, ZN => n24640);
   U21915 : OR2_X1 port map( A1 => n28496, A2 => n6642, Z => n10510);
   U21917 : XOR2_X1 port map( A1 => n26726, A2 => n28403, Z => n2174);
   U21918 : XOR2_X1 port map( A1 => n981, A2 => n22804, Z => n28403);
   U21921 : NOR2_X1 port map( A1 => n20291, A2 => n20294, ZN => n7733);
   U21923 : AOI22_X2 port map( A1 => n28404, A2 => n25077, B1 => n1661, B2 => 
                           n24966, ZN => n2897);
   U21924 : NAND2_X2 port map( A1 => n22650, A2 => n17496, ZN => n28404);
   U21926 : NAND2_X2 port map( A1 => n13968, A2 => n14207, ZN => n11161);
   U21927 : OAI21_X1 port map( A1 => n625, A2 => n622, B => n17433, ZN => n4721
                           );
   U21931 : XOR2_X1 port map( A1 => n25317, A2 => n23849, Z => n13136);
   U21933 : NAND3_X2 port map( A1 => n2967, A2 => n24677, A3 => n1447, ZN => 
                           n25317);
   U21934 : OR2_X1 port map( A1 => n1458, A2 => n23420, Z => n12157);
   U21937 : XOR2_X1 port map( A1 => n12192, A2 => n16747, Z => n26183);
   U21939 : NAND2_X2 port map( A1 => n24792, A2 => n5732, ZN => n12192);
   U21944 : OAI21_X2 port map( A1 => n14829, A2 => n14828, B => n28406, ZN => 
                           n19088);
   U21946 : BUF_X2 port map( I => n18099, Z => n28407);
   U21952 : NAND2_X1 port map( A1 => n27871, A2 => n5115, ZN => n5294);
   U21961 : XOR2_X1 port map( A1 => n3662, A2 => n3664, Z => n26510);
   U21964 : NAND2_X2 port map( A1 => n24533, A2 => n27091, ZN => n20570);
   U21967 : AOI22_X2 port map( A1 => n11136, A2 => n22106, B1 => n11134, B2 => 
                           n21022, ZN => n25778);
   U21970 : XOR2_X1 port map( A1 => n6134, A2 => n19537, Z => n24926);
   U21971 : AOI21_X1 port map( A1 => n21612, A2 => n12517, B => n21608, ZN => 
                           n28409);
   U21972 : NOR2_X1 port map( A1 => n18793, A2 => n26831, ZN => n3867);
   U21974 : XOR2_X1 port map( A1 => n12081, A2 => n12080, Z => n20559);
   U21975 : NAND3_X2 port map( A1 => n5767, A2 => n5766, A3 => n17203, ZN => 
                           n12708);
   U21980 : NAND2_X2 port map( A1 => n25209, A2 => n6365, ZN => n15732);
   U21981 : NAND2_X1 port map( A1 => n14710, A2 => n5977, ZN => n28411);
   U21983 : NAND2_X2 port map( A1 => n12896, A2 => n25367, ZN => n28412);
   U21985 : NAND2_X1 port map( A1 => n28413, A2 => n13012, ZN => n25481);
   U21986 : NAND2_X1 port map( A1 => n5221, A2 => n22589, ZN => n28413);
   U21988 : NAND3_X2 port map( A1 => n28414, A2 => n5849, A3 => n1579, ZN => 
                           n9027);
   U21989 : NAND2_X2 port map( A1 => n5850, A2 => n16694, ZN => n28414);
   U21990 : XOR2_X1 port map( A1 => n2145, A2 => n28415, Z => n23440);
   U21991 : XOR2_X1 port map( A1 => n26823, A2 => n8880, Z => n28415);
   U21993 : OR2_X1 port map( A1 => n12524, A2 => n8135, Z => n12802);
   U21995 : INV_X2 port map( I => n21101, ZN => n11905);
   U21996 : XOR2_X1 port map( A1 => n19201, A2 => n19267, Z => n15662);
   U21997 : NOR2_X2 port map( A1 => n23147, A2 => n2908, ZN => n19267);
   U21999 : XOR2_X1 port map( A1 => n27449, A2 => n17016, Z => n28416);
   U22000 : XOR2_X1 port map( A1 => n28417, A2 => n10705, Z => n17018);
   U22001 : XOR2_X1 port map( A1 => n17016, A2 => n7231, Z => n28417);
   U22002 : XOR2_X1 port map( A1 => n28418, A2 => n2294, Z => n26193);
   U22003 : XOR2_X1 port map( A1 => n25751, A2 => n954, Z => n28418);
   U22007 : OAI21_X2 port map( A1 => n28419, A2 => n20313, B => n5664, ZN => 
                           n7094);
   U22011 : NAND2_X2 port map( A1 => n28420, A2 => n23438, ZN => n21487);
   U22012 : NOR2_X2 port map( A1 => n11737, A2 => n13625, ZN => n28420);
   U22014 : XOR2_X1 port map( A1 => n25813, A2 => n28421, Z => n7480);
   U22015 : XOR2_X1 port map( A1 => n18135, A2 => n3775, Z => n28421);
   U22017 : NAND3_X1 port map( A1 => n21685, A2 => n933, A3 => n721, ZN => 
                           n6035);
   U22018 : XOR2_X1 port map( A1 => n2743, A2 => n12261, Z => n2742);
   U22020 : NOR2_X1 port map( A1 => n14844, A2 => n1998, ZN => n24038);
   U22021 : NOR3_X2 port map( A1 => n7675, A2 => n28423, A3 => n28422, ZN => 
                           n7673);
   U22024 : NOR2_X1 port map( A1 => n2427, A2 => n3723, ZN => n28424);
   U22025 : XOR2_X1 port map( A1 => n4707, A2 => n16774, Z => n23865);
   U22026 : XOR2_X1 port map( A1 => n11103, A2 => n16941, Z => n16774);
   U22027 : XOR2_X1 port map( A1 => n7896, A2 => n3000, Z => n1420);
   U22028 : XOR2_X1 port map( A1 => n28531, A2 => n20304, Z => n3000);
   U22030 : OAI21_X2 port map( A1 => n23296, A2 => n22710, B => n21782, ZN => 
                           n28426);
   U22035 : BUF_X2 port map( I => n21389, Z => n28428);
   U22036 : XOR2_X1 port map( A1 => n28429, A2 => n14709, Z => n22889);
   U22039 : XOR2_X1 port map( A1 => n4420, A2 => n22363, Z => n28429);
   U22042 : NAND2_X1 port map( A1 => n8533, A2 => n8532, ZN => n25059);
   U22044 : NAND2_X1 port map( A1 => n1104, A2 => n2185, ZN => n24590);
   U22046 : XOR2_X1 port map( A1 => n1591, A2 => n1588, Z => n12396);
   U22048 : NAND3_X1 port map( A1 => n9829, A2 => n14254, A3 => n9830, ZN => 
                           n10228);
   U22049 : XOR2_X1 port map( A1 => n10378, A2 => n18180, Z => n18319);
   U22050 : INV_X2 port map( I => n28430, ZN => n10671);
   U22052 : XOR2_X1 port map( A1 => n19481, A2 => n12939, Z => n28430);
   U22054 : AOI21_X2 port map( A1 => n28433, A2 => n28431, B => n21669, ZN => 
                           n22695);
   U22055 : INV_X2 port map( I => n5673, ZN => n28433);
   U22058 : XOR2_X1 port map( A1 => n24843, A2 => n28435, Z => n22365);
   U22062 : XOR2_X1 port map( A1 => n25080, A2 => n15332, Z => n28435);
   U22064 : NAND2_X2 port map( A1 => n12346, A2 => n28436, ZN => n10474);
   U22065 : OR2_X2 port map( A1 => n2631, A2 => n24010, Z => n2057);
   U22071 : XOR2_X1 port map( A1 => n17127, A2 => n28438, Z => n9539);
   U22072 : NAND3_X1 port map( A1 => n13660, A2 => n26625, A3 => n24235, ZN => 
                           n9687);
   U22076 : XOR2_X1 port map( A1 => n28440, A2 => n7590, Z => n7586);
   U22080 : AND2_X1 port map( A1 => n15010, A2 => n25500, Z => n18371);
   U22083 : NAND2_X2 port map( A1 => n3861, A2 => n19839, ZN => n28441);
   U22084 : NOR2_X2 port map( A1 => n25283, A2 => n10650, ZN => n15547);
   U22085 : NAND2_X2 port map( A1 => n3866, A2 => n3865, ZN => n22768);
   U22086 : XOR2_X1 port map( A1 => n10998, A2 => n18328, Z => n10997);
   U22087 : NAND3_X2 port map( A1 => n26437, A2 => n6690, A3 => n17903, ZN => 
                           n6691);
   U22088 : INV_X2 port map( I => n22237, ZN => n28442);
   U22089 : INV_X4 port map( I => n9216, ZN => n1163);
   U22090 : NAND2_X2 port map( A1 => n13755, A2 => n14845, ZN => n28443);
   U22091 : XOR2_X1 port map( A1 => n17114, A2 => n5327, Z => n16411);
   U22092 : XOR2_X1 port map( A1 => n15675, A2 => n15694, Z => n7138);
   U22093 : XOR2_X1 port map( A1 => n18321, A2 => n28445, Z => n25806);
   U22094 : XOR2_X1 port map( A1 => n16922, A2 => n28447, Z => n3778);
   U22095 : XOR2_X1 port map( A1 => n62, A2 => n16819, Z => n28447);
   U22096 : NAND3_X2 port map( A1 => n2686, A2 => n26142, A3 => n28448, ZN => 
                           n14228);
   U22097 : NAND3_X2 port map( A1 => n914, A2 => n7226, A3 => n1268, ZN => 
                           n28448);
   U22098 : OAI22_X2 port map( A1 => n26009, A2 => n2599, B1 => n13422, B2 => 
                           n23401, ZN => n28449);
   U22099 : OAI22_X1 port map( A1 => n13307, A2 => n11223, B1 => n16063, B2 => 
                           n7053, ZN => n8409);
   U22100 : INV_X2 port map( I => n8407, ZN => n11223);
   U22101 : XOR2_X1 port map( A1 => n7748, A2 => Key(147), Z => n8407);
   U22102 : BUF_X4 port map( I => n6293, Z => n21793);
   U22103 : OAI21_X2 port map( A1 => n8978, A2 => n14592, B => n17061, ZN => 
                           n12610);
   U22104 : XOR2_X1 port map( A1 => n18167, A2 => n18348, Z => n24719);
   U22105 : NAND2_X2 port map( A1 => n9631, A2 => n9632, ZN => n6508);
   U22106 : OAI22_X2 port map( A1 => n4470, A2 => n6591, B1 => n6590, B2 => 
                           n6813, ZN => n14754);
   U22107 : NAND2_X2 port map( A1 => n24268, A2 => n26350, ZN => n24267);
   U22108 : XOR2_X1 port map( A1 => n14962, A2 => n15220, Z => n14538);
   U22109 : XOR2_X1 port map( A1 => n16825, A2 => n28450, Z => n5531);
   U22110 : XOR2_X1 port map( A1 => n16529, A2 => n27513, Z => n28450);
   U22111 : XOR2_X1 port map( A1 => n24944, A2 => n28451, Z => n17532);
   U22112 : XOR2_X1 port map( A1 => n17046, A2 => n25497, Z => n28451);
   U22113 : XOR2_X1 port map( A1 => n18140, A2 => n18139, Z => n18146);
   U22114 : OAI21_X1 port map( A1 => n23056, A2 => n15462, B => n17617, ZN => 
                           n2953);
   U22115 : NAND2_X1 port map( A1 => n8558, A2 => n8560, ZN => n28452);
   U22116 : NAND2_X2 port map( A1 => n28453, A2 => n14257, ZN => n25276);
   U22117 : XOR2_X1 port map( A1 => n28454, A2 => n6001, Z => n14795);
   U22118 : XOR2_X1 port map( A1 => n20420, A2 => n23585, Z => n28454);
   U22119 : XOR2_X1 port map( A1 => n26083, A2 => n22470, Z => n19684);
   U22120 : NOR2_X2 port map( A1 => n13770, A2 => n21447, ZN => n10844);
   U22121 : XOR2_X1 port map( A1 => n18217, A2 => n21651, Z => n6702);
   U22122 : NOR2_X1 port map( A1 => n15197, A2 => n24927, ZN => n25855);
   U22123 : AND2_X1 port map( A1 => n17460, A2 => n6293, Z => n17205);
   U22124 : XOR2_X1 port map( A1 => n19509, A2 => n19327, Z => n14940);
   U22125 : INV_X2 port map( I => n28455, ZN => n28551);
   U22126 : XOR2_X1 port map( A1 => n23565, A2 => n15356, Z => n28455);
   U22127 : NOR2_X2 port map( A1 => n12311, A2 => n28456, ZN => n12488);
   U22128 : NAND2_X2 port map( A1 => n28458, A2 => n5617, ZN => n16433);
   U22129 : NOR2_X2 port map( A1 => n841, A2 => n22991, ZN => n28461);
   U22130 : AOI21_X2 port map( A1 => n6690, A2 => n17904, B => n728, ZN => 
                           n26539);
   U22131 : XOR2_X1 port map( A1 => n9345, A2 => n19285, Z => n19528);
   U22132 : AOI21_X2 port map( A1 => n4171, A2 => n18961, B => n18960, ZN => 
                           n9345);
   U22133 : NAND2_X2 port map( A1 => n25898, A2 => n28462, ZN => n7308);
   U22134 : AOI21_X2 port map( A1 => n8868, A2 => n16106, B => n26488, ZN => 
                           n28462);
   U22135 : XOR2_X1 port map( A1 => n22757, A2 => n28463, Z => n19173);
   U22136 : NAND2_X1 port map( A1 => n13009, A2 => n11522, ZN => n13032);
   U22137 : NAND2_X2 port map( A1 => n24849, A2 => n3691, ZN => n13009);
   U22138 : OAI22_X2 port map( A1 => n9307, A2 => n12922, B1 => n9306, B2 => 
                           n9305, ZN => n13684);
   U22139 : BUF_X2 port map( I => n23480, Z => n28465);
   U22140 : XOR2_X1 port map( A1 => n7975, A2 => n8983, Z => n24096);
   U22141 : NAND3_X2 port map( A1 => n9138, A2 => n1429, A3 => n17684, ZN => 
                           n18071);
   U22142 : AND2_X1 port map( A1 => n1468, A2 => n1470, Z => n28478);
   U22143 : INV_X2 port map( I => n8546, ZN => n25216);
   U22144 : NAND2_X2 port map( A1 => n12950, A2 => n28467, ZN => n10894);
   U22145 : NOR2_X2 port map( A1 => n5211, A2 => n6075, ZN => n28467);
   U22146 : AND2_X1 port map( A1 => n14528, A2 => n17474, Z => n26472);
   U22147 : AOI21_X2 port map( A1 => n22942, A2 => n3530, B => n26554, ZN => 
                           n21274);
   U22148 : OR2_X1 port map( A1 => n14510, A2 => n18665, Z => n26030);
   U22149 : NAND3_X2 port map( A1 => n17768, A2 => n23115, A3 => n25493, ZN => 
                           n17769);
   U22150 : AOI22_X2 port map( A1 => n16346, A2 => n16348, B1 => n10186, B2 => 
                           n11, ZN => n6617);
   U22151 : XOR2_X1 port map( A1 => n25345, A2 => n5653, Z => n19319);
   U22152 : NAND2_X2 port map( A1 => n5433, A2 => n5652, ZN => n5653);
   U22153 : NAND2_X2 port map( A1 => n16447, A2 => n16446, ZN => n26578);
   U22154 : INV_X2 port map( I => n20626, ZN => n20623);
   U22155 : NAND3_X2 port map( A1 => n28471, A2 => n9119, A3 => n28470, ZN => 
                           n5578);
   U22156 : NAND2_X2 port map( A1 => n28472, A2 => n270, ZN => n819);
   U22157 : NAND2_X2 port map( A1 => n16597, A2 => n16640, ZN => n16403);
   U22158 : NOR2_X2 port map( A1 => n16023, A2 => n14881, ZN => n16597);
   U22159 : NOR2_X2 port map( A1 => n17728, A2 => n23245, ZN => n17656);
   U22160 : AOI21_X2 port map( A1 => n24687, A2 => n24686, B => n23815, ZN => 
                           n17728);
   U22161 : OAI21_X2 port map( A1 => n2739, A2 => n10272, B => n28473, ZN => 
                           n7749);
   U22162 : INV_X2 port map( I => n28474, ZN => n13695);
   U22163 : NAND2_X2 port map( A1 => n6982, A2 => n11409, ZN => n14203);
   U22164 : OAI21_X2 port map( A1 => n6538, A2 => n1048, B => n28475, ZN => 
                           n1968);
   U22165 : INV_X2 port map( I => n28476, ZN => n14843);
   U22166 : XOR2_X1 port map( A1 => Plaintext(138), A2 => Key(138), Z => n28476
                           );
   U22167 : XOR2_X1 port map( A1 => n28477, A2 => n682, Z => n22116);
   U22168 : XOR2_X1 port map( A1 => n23500, A2 => n24814, Z => n28477);
   U22169 : NAND2_X2 port map( A1 => n5099, A2 => n5100, ZN => n5080);
   U22170 : XOR2_X1 port map( A1 => n1534, A2 => n1535, Z => n3592);
   U22171 : NOR2_X1 port map( A1 => n7138, A2 => n8727, ZN => n2192);
   U22172 : NOR2_X2 port map( A1 => n24123, A2 => n28478, ZN => n632);
   U22173 : XOR2_X1 port map( A1 => n28479, A2 => n27365, Z => n5065);
   U22174 : XOR2_X1 port map( A1 => n5067, A2 => n27358, Z => n28479);
   U22175 : NOR2_X2 port map( A1 => n25167, A2 => n3102, ZN => n3101);
   U22176 : INV_X2 port map( I => n28480, ZN => n28554);
   U22177 : NAND2_X2 port map( A1 => n6568, A2 => n6567, ZN => n28480);
   U22178 : XOR2_X1 port map( A1 => n17013, A2 => n16943, Z => n8413);
   U22179 : NAND3_X2 port map( A1 => n25637, A2 => n10300, A3 => n9495, ZN => 
                           n6241);
   U22180 : NOR2_X2 port map( A1 => n22614, A2 => n15159, ZN => n16692);
   U22181 : NAND2_X2 port map( A1 => n3100, A2 => n23812, ZN => n12364);
   U22182 : INV_X2 port map( I => n28482, ZN => n18683);
   U22183 : NAND2_X2 port map( A1 => n19754, A2 => n2632, ZN => n28485);
   U22184 : NAND2_X1 port map( A1 => n5429, A2 => n10714, ZN => n28486);
   U22185 : NAND2_X1 port map( A1 => n18769, A2 => n1001, ZN => n28487);
   U22186 : BUF_X2 port map( I => n6699, Z => n28488);
   U22187 : NAND3_X2 port map( A1 => n11569, A2 => n217, A3 => n11572, ZN => 
                           n17694);
   U22188 : XOR2_X1 port map( A1 => n6202, A2 => n6201, Z => n20596);
   U22189 : XOR2_X1 port map( A1 => n11698, A2 => n28489, Z => n6144);
   U22190 : XOR2_X1 port map( A1 => n18283, A2 => n4560, Z => n28489);
   U22191 : AOI21_X2 port map( A1 => n24380, A2 => n5173, B => n6265, ZN => 
                           n14243);
   U22192 : INV_X2 port map( I => n14859, ZN => n28490);
   U22193 : OAI21_X2 port map( A1 => n28492, A2 => n28491, B => n4199, ZN => 
                           n18806);
   U22194 : INV_X1 port map( I => n25176, ZN => n28491);
   U22195 : XOR2_X1 port map( A1 => n4026, A2 => n14686, Z => n22591);
   U22196 : XOR2_X1 port map( A1 => n6445, A2 => n24189, Z => n14686);
   U22197 : NOR2_X1 port map( A1 => n14986, A2 => n23083, ZN => n11661);
   U22198 : NAND3_X2 port map( A1 => n24897, A2 => n4875, A3 => n9856, ZN => 
                           n23083);
   U22199 : NOR2_X2 port map( A1 => n288, A2 => n22973, ZN => n14784);
   U22200 : XOR2_X1 port map( A1 => n13001, A2 => n19368, Z => n19176);
   U22201 : NAND2_X2 port map( A1 => n24558, A2 => n7793, ZN => n7794);
   U22202 : NAND2_X2 port map( A1 => n13102, A2 => n28494, ZN => n14137);
   U22203 : AOI22_X2 port map( A1 => n15807, A2 => n6837, B1 => n16266, B2 => 
                           n15808, ZN => n28494);
   U22204 : XOR2_X1 port map( A1 => n7052, A2 => n16801, Z => n5624);
   U22205 : OAI22_X2 port map( A1 => n6269, A2 => n6268, B1 => n913, B2 => n833
                           , ZN => n7052);
   U22206 : BUF_X2 port map( I => n4802, Z => n28495);
   U22207 : NAND2_X2 port map( A1 => n17847, A2 => n17989, ZN => n28496);
   U22208 : XOR2_X1 port map( A1 => n8260, A2 => n28498, Z => n28497);
   U22209 : OAI21_X1 port map( A1 => n11194, A2 => n11195, B => n3979, ZN => 
                           n23362);
   U22210 : XOR2_X1 port map( A1 => n18317, A2 => n18182, Z => n11999);
   U22211 : OR2_X1 port map( A1 => n23538, A2 => n18740, Z => n18419);
   U22212 : XOR2_X1 port map( A1 => n8003, A2 => n8002, Z => n23538);
   U22213 : OR2_X2 port map( A1 => n24308, A2 => n14117, Z => n4415);
   U22214 : AOI22_X1 port map( A1 => n11841, A2 => n11840, B1 => n19090, B2 => 
                           n19092, ZN => n19524);
   U22215 : INV_X4 port map( I => n14879, ZN => n16587);
   U22216 : OAI22_X2 port map( A1 => n10503, A2 => n10504, B1 => n10505, B2 => 
                           n10507, ZN => n14879);
   U22217 : NAND2_X2 port map( A1 => n4255, A2 => n4256, ZN => n12360);
   U22218 : XOR2_X1 port map( A1 => n13856, A2 => n16874, Z => n7604);
   U22219 : XOR2_X1 port map( A1 => n22931, A2 => n15372, Z => n5450);
   U22220 : XOR2_X1 port map( A1 => n14701, A2 => n18015, Z => n3463);
   U22221 : XNOR2_X1 port map( A1 => n11780, A2 => n94, ZN => n17080);
   U22222 : NOR2_X2 port map( A1 => n10423, A2 => n22958, ZN => n11780);
   U22223 : XOR2_X1 port map( A1 => n22804, A2 => n28465, Z => n19455);
   U22224 : AOI21_X2 port map( A1 => n3239, A2 => n3238, B => n18577, ZN => 
                           n23480);
   U22225 : XOR2_X1 port map( A1 => n16965, A2 => n10294, Z => n14023);
   U22226 : AOI21_X2 port map( A1 => n11068, A2 => n13897, B => n11067, ZN => 
                           n16965);
   U22227 : XOR2_X1 port map( A1 => n19497, A2 => n12948, Z => n19253);
   U22228 : NAND2_X2 port map( A1 => n18963, A2 => n3833, ZN => n22001);
   U22229 : NAND2_X2 port map( A1 => n14188, A2 => n3312, ZN => n18963);
   U22230 : XOR2_X1 port map( A1 => n18292, A2 => n9736, Z => n10285);
   U22231 : XOR2_X1 port map( A1 => n18069, A2 => n18063, Z => n18292);
   U22232 : XOR2_X1 port map( A1 => n16809, A2 => n17053, Z => n16990);
   U22233 : NOR2_X2 port map( A1 => n1983, A2 => n10599, ZN => n16809);
   U22234 : NAND2_X2 port map( A1 => n23481, A2 => n24744, ZN => n28505);
   U22235 : NAND2_X1 port map( A1 => n3443, A2 => n12839, ZN => n14344);
   U22236 : NAND2_X2 port map( A1 => n18673, A2 => n24672, ZN => n3062);
   U22237 : XOR2_X1 port map( A1 => n1099, A2 => n4137, Z => n24095);
   U22238 : NAND2_X2 port map( A1 => n28506, A2 => n5539, ZN => n18733);
   U22239 : OAI21_X2 port map( A1 => n28509, A2 => n28508, B => n1080, ZN => 
                           n9807);
   U22240 : BUF_X2 port map( I => n25439, Z => n28510);
   U22241 : OAI21_X2 port map( A1 => n135, A2 => n28512, B => n28511, ZN => 
                           n20045);
   U22242 : INV_X2 port map( I => n24534, ZN => n28512);
   U22243 : AOI21_X1 port map( A1 => n21215, A2 => n21230, B => n21214, ZN => 
                           n14136);
   U22244 : AOI22_X2 port map( A1 => n10268, A2 => n6756, B1 => n9494, B2 => 
                           n26059, ZN => n21230);
   U22245 : NAND2_X2 port map( A1 => n3465, A2 => n15367, ZN => n24553);
   U22246 : NAND2_X2 port map( A1 => n19602, A2 => n28513, ZN => n6006);
   U22247 : OAI22_X2 port map( A1 => n15376, A2 => n19599, B1 => n977, B2 => 
                           n14423, ZN => n28513);
   U22248 : NOR3_X2 port map( A1 => n23700, A2 => n23558, A3 => n20186, ZN => 
                           n11051);
   U22249 : XOR2_X1 port map( A1 => n19419, A2 => n28514, Z => n26409);
   U22250 : INV_X2 port map( I => n4690, ZN => n28515);
   U22251 : NOR2_X2 port map( A1 => n737, A2 => n9508, ZN => n4690);
   U22252 : NAND3_X2 port map( A1 => n12876, A2 => n25590, A3 => n23804, ZN => 
                           n13524);
   U22253 : NAND2_X1 port map( A1 => n9236, A2 => n18426, ZN => n28516);
   U22254 : XOR2_X1 port map( A1 => n9102, A2 => n535, Z => n3338);
   U22255 : NAND2_X2 port map( A1 => n28520, A2 => n16237, ZN => n22572);
   U22256 : OAI21_X2 port map( A1 => n16232, A2 => n16233, B => n25816, ZN => 
                           n28520);
   U22257 : BUF_X2 port map( I => n21386, Z => n28521);
   U22258 : OAI21_X2 port map( A1 => n11088, A2 => n6593, B => n11087, ZN => 
                           n12195);
   U22259 : XOR2_X1 port map( A1 => n1912, A2 => n25356, Z => n20549);
   U22260 : NAND2_X2 port map( A1 => n1475, A2 => n1914, ZN => n25356);
   U22261 : BUF_X2 port map( I => n4709, Z => n28524);
   U22262 : NAND2_X2 port map( A1 => n28526, A2 => n2214, ZN => n2215);
   U22263 : NAND2_X1 port map( A1 => n7569, A2 => n11580, ZN => n8133);
   U22264 : BUF_X2 port map( I => n19264, Z => n28527);
   U22265 : AND2_X1 port map( A1 => n20431, A2 => n20200, Z => n24921);
   U22266 : XOR2_X1 port map( A1 => n9802, A2 => n18048, Z => n12742);
   U22267 : XOR2_X1 port map( A1 => n24938, A2 => n28528, Z => n21916);
   U22268 : XOR2_X1 port map( A1 => n19317, A2 => n6416, Z => n28528);
   U22269 : NAND2_X2 port map( A1 => n6987, A2 => n13194, ZN => n4088);
   U22270 : XOR2_X1 port map( A1 => n9477, A2 => n27623, Z => n28529);
   U22271 : XOR2_X1 port map( A1 => n1190, A2 => n24963, Z => n28530);
   U22272 : XOR2_X1 port map( A1 => n3869, A2 => n2998, Z => n24715);
   U22273 : NAND2_X2 port map( A1 => n13207, A2 => n28532, ZN => n12410);
   U22274 : AOI22_X2 port map( A1 => n24648, A2 => n3399, B1 => n16679, B2 => 
                           n16418, ZN => n28532);
   U22275 : NAND2_X2 port map( A1 => n28533, A2 => n6021, ZN => n13687);
   U22276 : NAND2_X2 port map( A1 => n4446, A2 => n8348, ZN => n28533);
   U22277 : XOR2_X1 port map( A1 => n19265, A2 => n19306, Z => n19237);
   U22278 : XOR2_X1 port map( A1 => n4128, A2 => n25507, Z => n4127);
   U22279 : OAI21_X1 port map( A1 => n10461, A2 => n28535, B => n28534, ZN => 
                           n5146);
   U22280 : OAI21_X1 port map( A1 => n8125, A2 => n24567, B => n10461, ZN => 
                           n28534);
   U22281 : NAND2_X2 port map( A1 => n2660, A2 => n2659, ZN => n8373);
   U22282 : INV_X2 port map( I => n19005, ZN => n3693);
   U22283 : OR2_X1 port map( A1 => n24235, A2 => n13660, Z => n148);
   U22284 : INV_X2 port map( I => n2631, ZN => n19796);
   U22285 : XNOR2_X1 port map( A1 => n13631, A2 => n7031, ZN => n28537);
   U22286 : INV_X2 port map( I => n17578, ZN => n25607);
   U22287 : INV_X2 port map( I => n9454, ZN => n25922);
   U22288 : AND2_X1 port map( A1 => n18694, A2 => n26880, Z => n28544);
   U22289 : NAND2_X2 port map( A1 => n999, A2 => n28019, ZN => n6834);
   U22290 : OAI21_X2 port map( A1 => n4090, A2 => n4089, B => n18429, ZN => 
                           n19148);
   U22291 : INV_X2 port map( I => n19889, ZN => n23782);
   U22292 : XNOR2_X1 port map( A1 => n4966, A2 => n14630, ZN => n28549);
   U22293 : XNOR2_X1 port map( A1 => n15130, A2 => n15242, ZN => n28550);
   U22294 : OAI21_X2 port map( A1 => n15180, A2 => n6321, B => n6318, ZN => 
                           n25370);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Top is

   port( clk : in std_logic;  Plaintext, Key : in std_logic_vector (191 downto 
         0);  Ciphertext : out std_logic_vector (191 downto 0));

end SPEEDY_Top;

architecture SYN_Behavioral of SPEEDY_Top is

   component DFFRNQ_X1
      port( D, CLK, RN : in std_logic;  Q : out std_logic);
   end component;
   
   component SPEEDY_Rounds5_0
      port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : 
            out std_logic_vector (191 downto 0));
   end component;
   
   component DFFSNQ_X1
      port( D, CLK, SN : in std_logic;  Q : out std_logic);
   end component;
   
   signal reg_in_191_port, reg_in_190_port, reg_in_189_port, reg_in_188_port, 
      reg_in_187_port, reg_in_186_port, reg_in_185_port, reg_in_184_port, 
      reg_in_183_port, reg_in_182_port, reg_in_181_port, reg_in_180_port, 
      reg_in_179_port, reg_in_178_port, reg_in_177_port, reg_in_176_port, 
      reg_in_175_port, reg_in_174_port, reg_in_173_port, reg_in_172_port, 
      reg_in_171_port, reg_in_170_port, reg_in_169_port, reg_in_168_port, 
      reg_in_167_port, reg_in_166_port, reg_in_165_port, reg_in_164_port, 
      reg_in_163_port, reg_in_162_port, reg_in_161_port, reg_in_160_port, 
      reg_in_159_port, reg_in_158_port, reg_in_157_port, reg_in_156_port, 
      reg_in_155_port, reg_in_154_port, reg_in_153_port, reg_in_152_port, 
      reg_in_151_port, reg_in_150_port, reg_in_149_port, reg_in_148_port, 
      reg_in_147_port, reg_in_146_port, reg_in_145_port, reg_in_144_port, 
      reg_in_143_port, reg_in_142_port, reg_in_141_port, reg_in_140_port, 
      reg_in_139_port, reg_in_138_port, reg_in_137_port, reg_in_136_port, 
      reg_in_135_port, reg_in_134_port, reg_in_133_port, reg_in_132_port, 
      reg_in_131_port, reg_in_130_port, reg_in_129_port, reg_in_128_port, 
      reg_in_127_port, reg_in_126_port, reg_in_125_port, reg_in_124_port, 
      reg_in_123_port, reg_in_122_port, reg_in_121_port, reg_in_120_port, 
      reg_in_119_port, reg_in_118_port, reg_in_117_port, reg_in_116_port, 
      reg_in_115_port, reg_in_114_port, reg_in_113_port, reg_in_112_port, 
      reg_in_111_port, reg_in_110_port, reg_in_109_port, reg_in_108_port, 
      reg_in_107_port, reg_in_106_port, reg_in_105_port, reg_in_104_port, 
      reg_in_103_port, reg_in_102_port, reg_in_101_port, reg_in_100_port, 
      reg_in_99_port, reg_in_98_port, reg_in_97_port, reg_in_96_port, 
      reg_in_95_port, reg_in_94_port, reg_in_93_port, reg_in_92_port, 
      reg_in_91_port, reg_in_90_port, reg_in_89_port, reg_in_88_port, 
      reg_in_87_port, reg_in_86_port, reg_in_85_port, reg_in_84_port, 
      reg_in_83_port, reg_in_82_port, reg_in_81_port, reg_in_80_port, 
      reg_in_79_port, reg_in_78_port, reg_in_77_port, reg_in_76_port, 
      reg_in_75_port, reg_in_74_port, reg_in_73_port, reg_in_72_port, 
      reg_in_71_port, reg_in_70_port, reg_in_69_port, reg_in_68_port, 
      reg_in_67_port, reg_in_66_port, reg_in_65_port, reg_in_64_port, 
      reg_in_63_port, reg_in_62_port, reg_in_61_port, reg_in_60_port, 
      reg_in_59_port, reg_in_58_port, reg_in_57_port, reg_in_56_port, 
      reg_in_55_port, reg_in_54_port, reg_in_53_port, reg_in_52_port, 
      reg_in_51_port, reg_in_50_port, reg_in_49_port, reg_in_48_port, 
      reg_in_47_port, reg_in_46_port, reg_in_45_port, reg_in_44_port, 
      reg_in_43_port, reg_in_42_port, reg_in_41_port, reg_in_40_port, 
      reg_in_39_port, reg_in_38_port, reg_in_37_port, reg_in_36_port, 
      reg_in_35_port, reg_in_34_port, reg_in_33_port, reg_in_32_port, 
      reg_in_31_port, reg_in_30_port, reg_in_29_port, reg_in_28_port, 
      reg_in_27_port, reg_in_26_port, reg_in_25_port, reg_in_24_port, 
      reg_in_23_port, reg_in_22_port, reg_in_21_port, reg_in_20_port, 
      reg_in_19_port, reg_in_18_port, reg_in_17_port, reg_in_16_port, 
      reg_in_15_port, reg_in_14_port, reg_in_13_port, reg_in_12_port, 
      reg_in_11_port, reg_in_10_port, reg_in_9_port, reg_in_8_port, 
      reg_in_7_port, reg_in_6_port, reg_in_5_port, reg_in_4_port, reg_in_3_port
      , reg_in_2_port, reg_in_1_port, reg_in_0_port, reg_key_191_port, 
      reg_key_190_port, reg_key_189_port, reg_key_188_port, reg_key_187_port, 
      reg_key_186_port, reg_key_185_port, reg_key_184_port, reg_key_183_port, 
      reg_key_182_port, reg_key_181_port, reg_key_180_port, reg_key_179_port, 
      reg_key_178_port, reg_key_177_port, reg_key_176_port, reg_key_175_port, 
      reg_key_174_port, reg_key_173_port, reg_key_172_port, reg_key_171_port, 
      reg_key_170_port, reg_key_169_port, reg_key_168_port, reg_key_167_port, 
      reg_key_166_port, reg_key_165_port, reg_key_164_port, reg_key_163_port, 
      reg_key_162_port, reg_key_161_port, reg_key_160_port, reg_key_159_port, 
      reg_key_158_port, reg_key_157_port, reg_key_156_port, reg_key_155_port, 
      reg_key_154_port, reg_key_153_port, reg_key_152_port, reg_key_151_port, 
      reg_key_150_port, reg_key_149_port, reg_key_148_port, reg_key_147_port, 
      reg_key_146_port, reg_key_145_port, reg_key_144_port, reg_key_143_port, 
      reg_key_142_port, reg_key_141_port, reg_key_140_port, reg_key_139_port, 
      reg_key_138_port, reg_key_137_port, reg_key_136_port, reg_key_135_port, 
      reg_key_134_port, reg_key_133_port, reg_key_132_port, reg_key_131_port, 
      reg_key_130_port, reg_key_129_port, reg_key_128_port, reg_key_127_port, 
      reg_key_126_port, reg_key_125_port, reg_key_124_port, reg_key_123_port, 
      reg_key_122_port, reg_key_121_port, reg_key_120_port, reg_key_119_port, 
      reg_key_118_port, reg_key_117_port, reg_key_116_port, reg_key_115_port, 
      reg_key_114_port, reg_key_113_port, reg_key_112_port, reg_key_111_port, 
      reg_key_110_port, reg_key_109_port, reg_key_108_port, reg_key_107_port, 
      reg_key_106_port, reg_key_105_port, reg_key_104_port, reg_key_103_port, 
      reg_key_102_port, reg_key_101_port, reg_key_100_port, reg_key_99_port, 
      reg_key_98_port, reg_key_97_port, reg_key_96_port, reg_key_95_port, 
      reg_key_94_port, reg_key_93_port, reg_key_92_port, reg_key_91_port, 
      reg_key_90_port, reg_key_89_port, reg_key_88_port, reg_key_87_port, 
      reg_key_86_port, reg_key_85_port, reg_key_84_port, reg_key_83_port, 
      reg_key_82_port, reg_key_81_port, reg_key_80_port, reg_key_79_port, 
      reg_key_78_port, reg_key_77_port, reg_key_76_port, reg_key_75_port, 
      reg_key_74_port, reg_key_73_port, reg_key_72_port, reg_key_71_port, 
      reg_key_70_port, reg_key_69_port, reg_key_68_port, reg_key_67_port, 
      reg_key_66_port, reg_key_65_port, reg_key_64_port, reg_key_63_port, 
      reg_key_62_port, reg_key_61_port, reg_key_60_port, reg_key_59_port, 
      reg_key_58_port, reg_key_57_port, reg_key_56_port, reg_key_55_port, 
      reg_key_54_port, reg_key_53_port, reg_key_52_port, reg_key_51_port, 
      reg_key_50_port, reg_key_49_port, reg_key_48_port, reg_key_47_port, 
      reg_key_46_port, reg_key_45_port, reg_key_44_port, reg_key_43_port, 
      reg_key_42_port, reg_key_41_port, reg_key_40_port, reg_key_39_port, 
      reg_key_38_port, reg_key_37_port, reg_key_36_port, reg_key_35_port, 
      reg_key_34_port, reg_key_33_port, reg_key_32_port, reg_key_31_port, 
      reg_key_30_port, reg_key_29_port, reg_key_28_port, reg_key_27_port, 
      reg_key_26_port, reg_key_25_port, reg_key_24_port, reg_key_23_port, 
      reg_key_22_port, reg_key_21_port, reg_key_20_port, reg_key_19_port, 
      reg_key_18_port, reg_key_17_port, reg_key_16_port, reg_key_15_port, 
      reg_key_14_port, reg_key_13_port, reg_key_12_port, reg_key_11_port, 
      reg_key_10_port, reg_key_9_port, reg_key_8_port, reg_key_7_port, 
      reg_key_6_port, reg_key_5_port, reg_key_4_port, reg_key_3_port, 
      reg_key_2_port, reg_key_1_port, reg_key_0_port, reg_out_191_port, 
      reg_out_190_port, reg_out_189_port, reg_out_188_port, reg_out_187_port, 
      reg_out_186_port, reg_out_185_port, reg_out_184_port, reg_out_183_port, 
      reg_out_182_port, reg_out_181_port, reg_out_180_port, reg_out_179_port, 
      reg_out_178_port, reg_out_177_port, reg_out_176_port, reg_out_175_port, 
      reg_out_174_port, reg_out_173_port, reg_out_172_port, reg_out_171_port, 
      reg_out_170_port, reg_out_169_port, reg_out_168_port, reg_out_167_port, 
      reg_out_166_port, reg_out_165_port, reg_out_164_port, reg_out_163_port, 
      reg_out_162_port, reg_out_161_port, reg_out_160_port, reg_out_159_port, 
      reg_out_158_port, reg_out_157_port, reg_out_156_port, reg_out_155_port, 
      reg_out_154_port, reg_out_153_port, reg_out_152_port, reg_out_151_port, 
      reg_out_150_port, reg_out_149_port, reg_out_148_port, reg_out_147_port, 
      reg_out_146_port, reg_out_145_port, reg_out_144_port, reg_out_143_port, 
      reg_out_142_port, reg_out_141_port, reg_out_140_port, reg_out_139_port, 
      reg_out_138_port, reg_out_137_port, reg_out_136_port, reg_out_135_port, 
      reg_out_134_port, reg_out_133_port, reg_out_132_port, reg_out_131_port, 
      reg_out_130_port, reg_out_129_port, reg_out_128_port, reg_out_127_port, 
      reg_out_126_port, reg_out_125_port, reg_out_124_port, reg_out_123_port, 
      reg_out_122_port, reg_out_121_port, reg_out_120_port, reg_out_119_port, 
      reg_out_118_port, reg_out_117_port, reg_out_116_port, reg_out_115_port, 
      reg_out_114_port, reg_out_113_port, reg_out_112_port, reg_out_111_port, 
      reg_out_110_port, reg_out_109_port, reg_out_108_port, reg_out_107_port, 
      reg_out_106_port, reg_out_105_port, reg_out_104_port, reg_out_103_port, 
      reg_out_102_port, reg_out_101_port, reg_out_100_port, reg_out_99_port, 
      reg_out_98_port, reg_out_97_port, reg_out_96_port, reg_out_95_port, 
      reg_out_94_port, reg_out_93_port, reg_out_92_port, reg_out_91_port, 
      reg_out_90_port, reg_out_89_port, reg_out_88_port, reg_out_87_port, 
      reg_out_86_port, reg_out_85_port, reg_out_84_port, reg_out_83_port, 
      reg_out_82_port, reg_out_81_port, reg_out_80_port, reg_out_79_port, 
      reg_out_78_port, reg_out_77_port, reg_out_76_port, reg_out_75_port, 
      reg_out_74_port, reg_out_73_port, reg_out_72_port, reg_out_71_port, 
      reg_out_70_port, reg_out_69_port, reg_out_68_port, reg_out_67_port, 
      reg_out_66_port, reg_out_65_port, reg_out_64_port, reg_out_63_port, 
      reg_out_62_port, reg_out_61_port, reg_out_60_port, reg_out_59_port, 
      reg_out_58_port, reg_out_57_port, reg_out_56_port, reg_out_55_port, 
      reg_out_54_port, reg_out_53_port, reg_out_52_port, reg_out_51_port, 
      reg_out_50_port, reg_out_49_port, reg_out_48_port, reg_out_47_port, 
      reg_out_46_port, reg_out_45_port, reg_out_44_port, reg_out_43_port, 
      reg_out_42_port, reg_out_41_port, reg_out_40_port, reg_out_39_port, 
      reg_out_38_port, reg_out_37_port, reg_out_36_port, reg_out_35_port, 
      reg_out_34_port, reg_out_33_port, reg_out_32_port, reg_out_31_port, 
      reg_out_30_port, reg_out_29_port, reg_out_28_port, reg_out_27_port, 
      reg_out_26_port, reg_out_25_port, reg_out_24_port, reg_out_23_port, 
      reg_out_22_port, reg_out_21_port, reg_out_20_port, reg_out_19_port, 
      reg_out_18_port, reg_out_17_port, reg_out_16_port, reg_out_15_port, 
      reg_out_14_port, reg_out_13_port, reg_out_12_port, reg_out_11_port, 
      reg_out_10_port, reg_out_9_port, reg_out_8_port, reg_out_7_port, 
      reg_out_6_port, reg_out_5_port, reg_out_4_port, reg_out_3_port, 
      reg_out_2_port, reg_out_1_port, reg_out_0_port, n2, n7, n8, n10, n15, n17
      , n19, n23, n24, n25, n26, n31, n32, n33, n36, n41, n43, n44, n45, n48, 
      n49, n50, n51, n55, n59, n62, n66, n69, n72, n73, n74, n75, n76, n78, n79
      , n80, n86, n87, n97, n98, n102, n103, n104, n107, n108, n109, n110, n114
      , n116, n117, n119, n122, n123, n124, n126, n131, n133, n136, n137, n138,
      n145, n146, n147, n148, n150, n151, n153, n154, n155, n157, n158, n161, 
      n162, n164, n165, n167, n168, n170, n172, n174, n176, n177, n180, n181, 
      n182, n183, n187, n191, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, 
      n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
      n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, 
      n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, 
      n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, 
      n579, n580, n581, n582, n583, n584, n585, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, 
      n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n654, 
      n655, n656, n657, n659, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692 : 
      std_logic;

begin
   
   reg_in_regx191x : DFFSNQ_X1 port map( D => Plaintext(191), CLK => clk, SN =>
                           n576, Q => reg_in_191_port);
   reg_in_regx190x : DFFSNQ_X1 port map( D => Plaintext(190), CLK => clk, SN =>
                           n575, Q => reg_in_190_port);
   reg_in_regx189x : DFFSNQ_X1 port map( D => Plaintext(189), CLK => clk, SN =>
                           n574, Q => reg_in_189_port);
   reg_in_regx188x : DFFSNQ_X1 port map( D => Plaintext(188), CLK => clk, SN =>
                           n573, Q => reg_in_188_port);
   reg_in_regx187x : DFFSNQ_X1 port map( D => Plaintext(187), CLK => clk, SN =>
                           n572, Q => reg_in_187_port);
   reg_in_regx186x : DFFSNQ_X1 port map( D => Plaintext(186), CLK => clk, SN =>
                           n571, Q => reg_in_186_port);
   reg_in_regx185x : DFFSNQ_X1 port map( D => Plaintext(185), CLK => clk, SN =>
                           n570, Q => reg_in_185_port);
   reg_in_regx184x : DFFSNQ_X1 port map( D => Plaintext(184), CLK => clk, SN =>
                           n569, Q => reg_in_184_port);
   reg_in_regx183x : DFFSNQ_X1 port map( D => Plaintext(183), CLK => clk, SN =>
                           n568, Q => reg_in_183_port);
   reg_in_regx182x : DFFSNQ_X1 port map( D => Plaintext(182), CLK => clk, SN =>
                           n567, Q => reg_in_182_port);
   reg_in_regx181x : DFFSNQ_X1 port map( D => Plaintext(181), CLK => clk, SN =>
                           n566, Q => reg_in_181_port);
   reg_in_regx180x : DFFSNQ_X1 port map( D => Plaintext(180), CLK => clk, SN =>
                           n565, Q => reg_in_180_port);
   reg_in_regx179x : DFFSNQ_X1 port map( D => Plaintext(179), CLK => clk, SN =>
                           n564, Q => reg_in_179_port);
   reg_in_regx178x : DFFSNQ_X1 port map( D => Plaintext(178), CLK => clk, SN =>
                           n563, Q => reg_in_178_port);
   reg_in_regx177x : DFFSNQ_X1 port map( D => Plaintext(177), CLK => clk, SN =>
                           n562, Q => reg_in_177_port);
   reg_in_regx176x : DFFSNQ_X1 port map( D => Plaintext(176), CLK => clk, SN =>
                           n561, Q => reg_in_176_port);
   reg_in_regx175x : DFFSNQ_X1 port map( D => Plaintext(175), CLK => clk, SN =>
                           n560, Q => reg_in_175_port);
   reg_in_regx174x : DFFSNQ_X1 port map( D => Plaintext(174), CLK => clk, SN =>
                           n559, Q => reg_in_174_port);
   reg_in_regx173x : DFFSNQ_X1 port map( D => Plaintext(173), CLK => clk, SN =>
                           n558, Q => reg_in_173_port);
   reg_in_regx172x : DFFSNQ_X1 port map( D => Plaintext(172), CLK => clk, SN =>
                           n557, Q => reg_in_172_port);
   reg_in_regx171x : DFFSNQ_X1 port map( D => Plaintext(171), CLK => clk, SN =>
                           n556, Q => reg_in_171_port);
   reg_in_regx170x : DFFSNQ_X1 port map( D => Plaintext(170), CLK => clk, SN =>
                           n555, Q => reg_in_170_port);
   reg_in_regx169x : DFFSNQ_X1 port map( D => Plaintext(169), CLK => clk, SN =>
                           n554, Q => reg_in_169_port);
   reg_in_regx168x : DFFSNQ_X1 port map( D => Plaintext(168), CLK => clk, SN =>
                           n553, Q => reg_in_168_port);
   reg_in_regx167x : DFFSNQ_X1 port map( D => Plaintext(167), CLK => clk, SN =>
                           n552, Q => reg_in_167_port);
   reg_in_regx166x : DFFSNQ_X1 port map( D => Plaintext(166), CLK => clk, SN =>
                           n551, Q => reg_in_166_port);
   reg_in_regx165x : DFFSNQ_X1 port map( D => Plaintext(165), CLK => clk, SN =>
                           n550, Q => reg_in_165_port);
   reg_in_regx164x : DFFSNQ_X1 port map( D => Plaintext(164), CLK => clk, SN =>
                           n549, Q => reg_in_164_port);
   reg_in_regx163x : DFFSNQ_X1 port map( D => Plaintext(163), CLK => clk, SN =>
                           n548, Q => reg_in_163_port);
   reg_in_regx162x : DFFSNQ_X1 port map( D => Plaintext(162), CLK => clk, SN =>
                           n547, Q => reg_in_162_port);
   reg_in_regx161x : DFFSNQ_X1 port map( D => Plaintext(161), CLK => clk, SN =>
                           n546, Q => reg_in_161_port);
   reg_in_regx160x : DFFSNQ_X1 port map( D => Plaintext(160), CLK => clk, SN =>
                           n545, Q => reg_in_160_port);
   reg_in_regx159x : DFFSNQ_X1 port map( D => Plaintext(159), CLK => clk, SN =>
                           n544, Q => reg_in_159_port);
   reg_in_regx158x : DFFSNQ_X1 port map( D => Plaintext(158), CLK => clk, SN =>
                           n543, Q => reg_in_158_port);
   reg_in_regx157x : DFFSNQ_X1 port map( D => Plaintext(157), CLK => clk, SN =>
                           n542, Q => reg_in_157_port);
   reg_in_regx156x : DFFSNQ_X1 port map( D => Plaintext(156), CLK => clk, SN =>
                           n541, Q => reg_in_156_port);
   reg_in_regx155x : DFFSNQ_X1 port map( D => Plaintext(155), CLK => clk, SN =>
                           n540, Q => reg_in_155_port);
   reg_in_regx154x : DFFSNQ_X1 port map( D => Plaintext(154), CLK => clk, SN =>
                           n539, Q => reg_in_154_port);
   reg_in_regx153x : DFFSNQ_X1 port map( D => Plaintext(153), CLK => clk, SN =>
                           n538, Q => reg_in_153_port);
   reg_in_regx152x : DFFSNQ_X1 port map( D => Plaintext(152), CLK => clk, SN =>
                           n537, Q => reg_in_152_port);
   reg_in_regx151x : DFFSNQ_X1 port map( D => Plaintext(151), CLK => clk, SN =>
                           n536, Q => reg_in_151_port);
   reg_in_regx150x : DFFSNQ_X1 port map( D => Plaintext(150), CLK => clk, SN =>
                           n535, Q => reg_in_150_port);
   reg_in_regx149x : DFFSNQ_X1 port map( D => Plaintext(149), CLK => clk, SN =>
                           n534, Q => reg_in_149_port);
   reg_in_regx148x : DFFSNQ_X1 port map( D => Plaintext(148), CLK => clk, SN =>
                           n533, Q => reg_in_148_port);
   reg_in_regx146x : DFFSNQ_X1 port map( D => Plaintext(146), CLK => clk, SN =>
                           n531, Q => reg_in_146_port);
   reg_in_regx145x : DFFSNQ_X1 port map( D => Plaintext(145), CLK => clk, SN =>
                           n530, Q => reg_in_145_port);
   reg_in_regx144x : DFFSNQ_X1 port map( D => Plaintext(144), CLK => clk, SN =>
                           n529, Q => reg_in_144_port);
   reg_in_regx143x : DFFSNQ_X1 port map( D => Plaintext(143), CLK => clk, SN =>
                           n528, Q => reg_in_143_port);
   reg_in_regx142x : DFFSNQ_X1 port map( D => Plaintext(142), CLK => clk, SN =>
                           n527, Q => reg_in_142_port);
   reg_in_regx141x : DFFSNQ_X1 port map( D => Plaintext(141), CLK => clk, SN =>
                           n526, Q => reg_in_141_port);
   reg_in_regx140x : DFFSNQ_X1 port map( D => Plaintext(140), CLK => clk, SN =>
                           n525, Q => reg_in_140_port);
   reg_in_regx139x : DFFSNQ_X1 port map( D => Plaintext(139), CLK => clk, SN =>
                           n524, Q => reg_in_139_port);
   reg_in_regx138x : DFFSNQ_X1 port map( D => Plaintext(138), CLK => clk, SN =>
                           n523, Q => reg_in_138_port);
   reg_in_regx137x : DFFSNQ_X1 port map( D => Plaintext(137), CLK => clk, SN =>
                           n522, Q => reg_in_137_port);
   reg_in_regx136x : DFFSNQ_X1 port map( D => Plaintext(136), CLK => clk, SN =>
                           n521, Q => reg_in_136_port);
   reg_in_regx135x : DFFSNQ_X1 port map( D => Plaintext(135), CLK => clk, SN =>
                           n520, Q => reg_in_135_port);
   reg_in_regx134x : DFFSNQ_X1 port map( D => Plaintext(134), CLK => clk, SN =>
                           n519, Q => reg_in_134_port);
   reg_in_regx133x : DFFSNQ_X1 port map( D => Plaintext(133), CLK => clk, SN =>
                           n518, Q => reg_in_133_port);
   reg_in_regx132x : DFFSNQ_X1 port map( D => Plaintext(132), CLK => clk, SN =>
                           n517, Q => reg_in_132_port);
   reg_in_regx130x : DFFSNQ_X1 port map( D => Plaintext(130), CLK => clk, SN =>
                           n515, Q => reg_in_130_port);
   reg_in_regx129x : DFFSNQ_X1 port map( D => Plaintext(129), CLK => clk, SN =>
                           n514, Q => reg_in_129_port);
   reg_in_regx128x : DFFSNQ_X1 port map( D => Plaintext(128), CLK => clk, SN =>
                           n513, Q => reg_in_128_port);
   reg_in_regx127x : DFFSNQ_X1 port map( D => Plaintext(127), CLK => clk, SN =>
                           n512, Q => reg_in_127_port);
   reg_in_regx126x : DFFSNQ_X1 port map( D => Plaintext(126), CLK => clk, SN =>
                           n511, Q => reg_in_126_port);
   reg_in_regx125x : DFFSNQ_X1 port map( D => Plaintext(125), CLK => clk, SN =>
                           n510, Q => reg_in_125_port);
   reg_in_regx124x : DFFSNQ_X1 port map( D => Plaintext(124), CLK => clk, SN =>
                           n509, Q => reg_in_124_port);
   reg_in_regx123x : DFFSNQ_X1 port map( D => Plaintext(123), CLK => clk, SN =>
                           n508, Q => reg_in_123_port);
   reg_in_regx122x : DFFSNQ_X1 port map( D => Plaintext(122), CLK => clk, SN =>
                           n507, Q => reg_in_122_port);
   reg_in_regx121x : DFFSNQ_X1 port map( D => Plaintext(121), CLK => clk, SN =>
                           n506, Q => reg_in_121_port);
   reg_in_regx120x : DFFSNQ_X1 port map( D => Plaintext(120), CLK => clk, SN =>
                           n505, Q => reg_in_120_port);
   reg_in_regx119x : DFFSNQ_X1 port map( D => Plaintext(119), CLK => clk, SN =>
                           n504, Q => reg_in_119_port);
   reg_in_regx118x : DFFSNQ_X1 port map( D => Plaintext(118), CLK => clk, SN =>
                           n503, Q => reg_in_118_port);
   reg_in_regx117x : DFFSNQ_X1 port map( D => Plaintext(117), CLK => clk, SN =>
                           n502, Q => reg_in_117_port);
   reg_in_regx116x : DFFSNQ_X1 port map( D => Plaintext(116), CLK => clk, SN =>
                           n501, Q => reg_in_116_port);
   reg_in_regx115x : DFFSNQ_X1 port map( D => Plaintext(115), CLK => clk, SN =>
                           n500, Q => reg_in_115_port);
   reg_in_regx114x : DFFSNQ_X1 port map( D => Plaintext(114), CLK => clk, SN =>
                           n499, Q => reg_in_114_port);
   reg_in_regx113x : DFFSNQ_X1 port map( D => Plaintext(113), CLK => clk, SN =>
                           n498, Q => reg_in_113_port);
   reg_in_regx112x : DFFSNQ_X1 port map( D => Plaintext(112), CLK => clk, SN =>
                           n497, Q => reg_in_112_port);
   reg_in_regx111x : DFFSNQ_X1 port map( D => Plaintext(111), CLK => clk, SN =>
                           n496, Q => reg_in_111_port);
   reg_in_regx110x : DFFSNQ_X1 port map( D => Plaintext(110), CLK => clk, SN =>
                           n495, Q => reg_in_110_port);
   reg_in_regx109x : DFFSNQ_X1 port map( D => Plaintext(109), CLK => clk, SN =>
                           n494, Q => reg_in_109_port);
   reg_in_regx108x : DFFSNQ_X1 port map( D => Plaintext(108), CLK => clk, SN =>
                           n493, Q => reg_in_108_port);
   reg_in_regx107x : DFFSNQ_X1 port map( D => Plaintext(107), CLK => clk, SN =>
                           n492, Q => reg_in_107_port);
   reg_in_regx106x : DFFSNQ_X1 port map( D => Plaintext(106), CLK => clk, SN =>
                           n491, Q => reg_in_106_port);
   reg_in_regx105x : DFFSNQ_X1 port map( D => Plaintext(105), CLK => clk, SN =>
                           n490, Q => reg_in_105_port);
   reg_in_regx104x : DFFSNQ_X1 port map( D => Plaintext(104), CLK => clk, SN =>
                           n489, Q => reg_in_104_port);
   reg_in_regx103x : DFFSNQ_X1 port map( D => Plaintext(103), CLK => clk, SN =>
                           n488, Q => reg_in_103_port);
   reg_in_regx102x : DFFSNQ_X1 port map( D => Plaintext(102), CLK => clk, SN =>
                           n487, Q => reg_in_102_port);
   reg_in_regx101x : DFFSNQ_X1 port map( D => Plaintext(101), CLK => clk, SN =>
                           n486, Q => reg_in_101_port);
   reg_in_regx100x : DFFSNQ_X1 port map( D => Plaintext(100), CLK => clk, SN =>
                           n485, Q => reg_in_100_port);
   reg_in_regx99x : DFFSNQ_X1 port map( D => Plaintext(99), CLK => clk, SN => 
                           n484, Q => reg_in_99_port);
   reg_in_regx98x : DFFSNQ_X1 port map( D => Plaintext(98), CLK => clk, SN => 
                           n483, Q => reg_in_98_port);
   reg_in_regx97x : DFFSNQ_X1 port map( D => Plaintext(97), CLK => clk, SN => 
                           n482, Q => reg_in_97_port);
   reg_in_regx96x : DFFSNQ_X1 port map( D => Plaintext(96), CLK => clk, SN => 
                           n481, Q => reg_in_96_port);
   reg_in_regx95x : DFFSNQ_X1 port map( D => Plaintext(95), CLK => clk, SN => 
                           n480, Q => reg_in_95_port);
   reg_in_regx94x : DFFSNQ_X1 port map( D => Plaintext(94), CLK => clk, SN => 
                           n479, Q => reg_in_94_port);
   reg_in_regx93x : DFFSNQ_X1 port map( D => Plaintext(93), CLK => clk, SN => 
                           n478, Q => reg_in_93_port);
   reg_in_regx92x : DFFSNQ_X1 port map( D => Plaintext(92), CLK => clk, SN => 
                           n477, Q => reg_in_92_port);
   reg_in_regx91x : DFFSNQ_X1 port map( D => Plaintext(91), CLK => clk, SN => 
                           n476, Q => reg_in_91_port);
   reg_in_regx90x : DFFSNQ_X1 port map( D => Plaintext(90), CLK => clk, SN => 
                           n475, Q => reg_in_90_port);
   reg_in_regx89x : DFFSNQ_X1 port map( D => Plaintext(89), CLK => clk, SN => 
                           n474, Q => reg_in_89_port);
   reg_in_regx88x : DFFSNQ_X1 port map( D => Plaintext(88), CLK => clk, SN => 
                           n473, Q => reg_in_88_port);
   reg_in_regx87x : DFFSNQ_X1 port map( D => Plaintext(87), CLK => clk, SN => 
                           n472, Q => reg_in_87_port);
   reg_in_regx86x : DFFSNQ_X1 port map( D => Plaintext(86), CLK => clk, SN => 
                           n471, Q => reg_in_86_port);
   reg_in_regx85x : DFFSNQ_X1 port map( D => Plaintext(85), CLK => clk, SN => 
                           n470, Q => reg_in_85_port);
   reg_in_regx84x : DFFSNQ_X1 port map( D => Plaintext(84), CLK => clk, SN => 
                           n469, Q => reg_in_84_port);
   reg_in_regx83x : DFFSNQ_X1 port map( D => Plaintext(83), CLK => clk, SN => 
                           n468, Q => reg_in_83_port);
   reg_in_regx82x : DFFSNQ_X1 port map( D => Plaintext(82), CLK => clk, SN => 
                           n467, Q => reg_in_82_port);
   reg_in_regx81x : DFFSNQ_X1 port map( D => Plaintext(81), CLK => clk, SN => 
                           n466, Q => reg_in_81_port);
   reg_in_regx80x : DFFSNQ_X1 port map( D => Plaintext(80), CLK => clk, SN => 
                           n465, Q => reg_in_80_port);
   reg_in_regx79x : DFFSNQ_X1 port map( D => Plaintext(79), CLK => clk, SN => 
                           n464, Q => reg_in_79_port);
   reg_in_regx78x : DFFSNQ_X1 port map( D => Plaintext(78), CLK => clk, SN => 
                           n463, Q => reg_in_78_port);
   reg_in_regx77x : DFFSNQ_X1 port map( D => Plaintext(77), CLK => clk, SN => 
                           n462, Q => reg_in_77_port);
   reg_in_regx76x : DFFSNQ_X1 port map( D => Plaintext(76), CLK => clk, SN => 
                           n461, Q => reg_in_76_port);
   reg_in_regx75x : DFFSNQ_X1 port map( D => Plaintext(75), CLK => clk, SN => 
                           n460, Q => reg_in_75_port);
   reg_in_regx74x : DFFSNQ_X1 port map( D => Plaintext(74), CLK => clk, SN => 
                           n459, Q => reg_in_74_port);
   reg_in_regx73x : DFFSNQ_X1 port map( D => Plaintext(73), CLK => clk, SN => 
                           n458, Q => reg_in_73_port);
   reg_in_regx72x : DFFSNQ_X1 port map( D => Plaintext(72), CLK => clk, SN => 
                           n457, Q => reg_in_72_port);
   reg_in_regx70x : DFFSNQ_X1 port map( D => Plaintext(70), CLK => clk, SN => 
                           n455, Q => reg_in_70_port);
   reg_in_regx69x : DFFSNQ_X1 port map( D => Plaintext(69), CLK => clk, SN => 
                           n454, Q => reg_in_69_port);
   reg_in_regx68x : DFFSNQ_X1 port map( D => Plaintext(68), CLK => clk, SN => 
                           n453, Q => reg_in_68_port);
   reg_in_regx67x : DFFSNQ_X1 port map( D => Plaintext(67), CLK => clk, SN => 
                           n452, Q => reg_in_67_port);
   reg_in_regx66x : DFFSNQ_X1 port map( D => Plaintext(66), CLK => clk, SN => 
                           n451, Q => reg_in_66_port);
   reg_in_regx65x : DFFSNQ_X1 port map( D => Plaintext(65), CLK => clk, SN => 
                           n450, Q => reg_in_65_port);
   reg_in_regx64x : DFFSNQ_X1 port map( D => Plaintext(64), CLK => clk, SN => 
                           n449, Q => reg_in_64_port);
   reg_in_regx63x : DFFSNQ_X1 port map( D => Plaintext(63), CLK => clk, SN => 
                           n448, Q => reg_in_63_port);
   reg_in_regx62x : DFFSNQ_X1 port map( D => Plaintext(62), CLK => clk, SN => 
                           n447, Q => reg_in_62_port);
   reg_in_regx61x : DFFSNQ_X1 port map( D => Plaintext(61), CLK => clk, SN => 
                           n446, Q => reg_in_61_port);
   reg_in_regx60x : DFFSNQ_X1 port map( D => Plaintext(60), CLK => clk, SN => 
                           n445, Q => reg_in_60_port);
   reg_in_regx59x : DFFSNQ_X1 port map( D => Plaintext(59), CLK => clk, SN => 
                           n444, Q => reg_in_59_port);
   reg_in_regx58x : DFFSNQ_X1 port map( D => Plaintext(58), CLK => clk, SN => 
                           n443, Q => reg_in_58_port);
   reg_in_regx57x : DFFSNQ_X1 port map( D => Plaintext(57), CLK => clk, SN => 
                           n442, Q => reg_in_57_port);
   reg_in_regx56x : DFFSNQ_X1 port map( D => Plaintext(56), CLK => clk, SN => 
                           n441, Q => reg_in_56_port);
   reg_in_regx55x : DFFSNQ_X1 port map( D => Plaintext(55), CLK => clk, SN => 
                           n440, Q => reg_in_55_port);
   reg_in_regx54x : DFFSNQ_X1 port map( D => Plaintext(54), CLK => clk, SN => 
                           n439, Q => reg_in_54_port);
   reg_in_regx53x : DFFSNQ_X1 port map( D => Plaintext(53), CLK => clk, SN => 
                           n438, Q => reg_in_53_port);
   reg_in_regx52x : DFFSNQ_X1 port map( D => Plaintext(52), CLK => clk, SN => 
                           n437, Q => reg_in_52_port);
   reg_in_regx50x : DFFSNQ_X1 port map( D => Plaintext(50), CLK => clk, SN => 
                           n435, Q => reg_in_50_port);
   reg_in_regx49x : DFFSNQ_X1 port map( D => Plaintext(49), CLK => clk, SN => 
                           n434, Q => reg_in_49_port);
   reg_in_regx48x : DFFSNQ_X1 port map( D => Plaintext(48), CLK => clk, SN => 
                           n433, Q => reg_in_48_port);
   reg_in_regx47x : DFFSNQ_X1 port map( D => Plaintext(47), CLK => clk, SN => 
                           n432, Q => reg_in_47_port);
   reg_in_regx46x : DFFSNQ_X1 port map( D => Plaintext(46), CLK => clk, SN => 
                           n431, Q => reg_in_46_port);
   reg_in_regx45x : DFFSNQ_X1 port map( D => Plaintext(45), CLK => clk, SN => 
                           n430, Q => reg_in_45_port);
   reg_in_regx44x : DFFSNQ_X1 port map( D => Plaintext(44), CLK => clk, SN => 
                           n429, Q => reg_in_44_port);
   reg_in_regx43x : DFFSNQ_X1 port map( D => Plaintext(43), CLK => clk, SN => 
                           n428, Q => reg_in_43_port);
   reg_in_regx42x : DFFSNQ_X1 port map( D => Plaintext(42), CLK => clk, SN => 
                           n427, Q => reg_in_42_port);
   reg_in_regx41x : DFFSNQ_X1 port map( D => Plaintext(41), CLK => clk, SN => 
                           n426, Q => reg_in_41_port);
   reg_in_regx40x : DFFSNQ_X1 port map( D => Plaintext(40), CLK => clk, SN => 
                           n425, Q => reg_in_40_port);
   reg_in_regx39x : DFFSNQ_X1 port map( D => Plaintext(39), CLK => clk, SN => 
                           n424, Q => reg_in_39_port);
   reg_in_regx38x : DFFSNQ_X1 port map( D => Plaintext(38), CLK => clk, SN => 
                           n423, Q => reg_in_38_port);
   reg_in_regx37x : DFFSNQ_X1 port map( D => Plaintext(37), CLK => clk, SN => 
                           n422, Q => reg_in_37_port);
   reg_in_regx36x : DFFSNQ_X1 port map( D => Plaintext(36), CLK => clk, SN => 
                           n421, Q => reg_in_36_port);
   reg_in_regx35x : DFFSNQ_X1 port map( D => Plaintext(35), CLK => clk, SN => 
                           n420, Q => reg_in_35_port);
   reg_in_regx34x : DFFSNQ_X1 port map( D => Plaintext(34), CLK => clk, SN => 
                           n419, Q => reg_in_34_port);
   reg_in_regx33x : DFFSNQ_X1 port map( D => Plaintext(33), CLK => clk, SN => 
                           n418, Q => reg_in_33_port);
   reg_in_regx32x : DFFSNQ_X1 port map( D => Plaintext(32), CLK => clk, SN => 
                           n417, Q => reg_in_32_port);
   reg_in_regx31x : DFFSNQ_X1 port map( D => Plaintext(31), CLK => clk, SN => 
                           n416, Q => reg_in_31_port);
   reg_in_regx30x : DFFSNQ_X1 port map( D => Plaintext(30), CLK => clk, SN => 
                           n415, Q => reg_in_30_port);
   reg_in_regx28x : DFFSNQ_X1 port map( D => Plaintext(28), CLK => clk, SN => 
                           n413, Q => reg_in_28_port);
   reg_in_regx27x : DFFSNQ_X1 port map( D => Plaintext(27), CLK => clk, SN => 
                           n412, Q => reg_in_27_port);
   reg_in_regx26x : DFFSNQ_X1 port map( D => Plaintext(26), CLK => clk, SN => 
                           n411, Q => reg_in_26_port);
   reg_in_regx25x : DFFSNQ_X1 port map( D => Plaintext(25), CLK => clk, SN => 
                           n410, Q => reg_in_25_port);
   reg_in_regx24x : DFFSNQ_X1 port map( D => Plaintext(24), CLK => clk, SN => 
                           n409, Q => reg_in_24_port);
   reg_in_regx23x : DFFSNQ_X1 port map( D => Plaintext(23), CLK => clk, SN => 
                           n408, Q => reg_in_23_port);
   reg_in_regx22x : DFFSNQ_X1 port map( D => Plaintext(22), CLK => clk, SN => 
                           n407, Q => reg_in_22_port);
   reg_in_regx21x : DFFSNQ_X1 port map( D => Plaintext(21), CLK => clk, SN => 
                           n406, Q => reg_in_21_port);
   reg_in_regx20x : DFFSNQ_X1 port map( D => Plaintext(20), CLK => clk, SN => 
                           n405, Q => reg_in_20_port);
   reg_in_regx19x : DFFSNQ_X1 port map( D => Plaintext(19), CLK => clk, SN => 
                           n404, Q => reg_in_19_port);
   reg_in_regx18x : DFFSNQ_X1 port map( D => Plaintext(18), CLK => clk, SN => 
                           n403, Q => reg_in_18_port);
   reg_in_regx17x : DFFSNQ_X1 port map( D => Plaintext(17), CLK => clk, SN => 
                           n402, Q => reg_in_17_port);
   reg_in_regx16x : DFFSNQ_X1 port map( D => Plaintext(16), CLK => clk, SN => 
                           n401, Q => reg_in_16_port);
   reg_in_regx15x : DFFSNQ_X1 port map( D => Plaintext(15), CLK => clk, SN => 
                           n400, Q => reg_in_15_port);
   reg_in_regx14x : DFFSNQ_X1 port map( D => Plaintext(14), CLK => clk, SN => 
                           n399, Q => reg_in_14_port);
   reg_in_regx13x : DFFSNQ_X1 port map( D => Plaintext(13), CLK => clk, SN => 
                           n398, Q => reg_in_13_port);
   reg_in_regx12x : DFFSNQ_X1 port map( D => Plaintext(12), CLK => clk, SN => 
                           n397, Q => reg_in_12_port);
   reg_in_regx11x : DFFSNQ_X1 port map( D => Plaintext(11), CLK => clk, SN => 
                           n396, Q => reg_in_11_port);
   reg_in_regx10x : DFFSNQ_X1 port map( D => Plaintext(10), CLK => clk, SN => 
                           n395, Q => reg_in_10_port);
   reg_in_regx9x : DFFSNQ_X1 port map( D => Plaintext(9), CLK => clk, SN => 
                           n394, Q => reg_in_9_port);
   reg_in_regx8x : DFFSNQ_X1 port map( D => Plaintext(8), CLK => clk, SN => 
                           n393, Q => reg_in_8_port);
   reg_in_regx7x : DFFSNQ_X1 port map( D => Plaintext(7), CLK => clk, SN => 
                           n392, Q => reg_in_7_port);
   reg_in_regx6x : DFFSNQ_X1 port map( D => Plaintext(6), CLK => clk, SN => 
                           n391, Q => reg_in_6_port);
   reg_in_regx5x : DFFSNQ_X1 port map( D => Plaintext(5), CLK => clk, SN => 
                           n390, Q => reg_in_5_port);
   reg_in_regx4x : DFFSNQ_X1 port map( D => Plaintext(4), CLK => clk, SN => 
                           n389, Q => reg_in_4_port);
   reg_in_regx3x : DFFSNQ_X1 port map( D => Plaintext(3), CLK => clk, SN => 
                           n388, Q => reg_in_3_port);
   reg_in_regx2x : DFFSNQ_X1 port map( D => Plaintext(2), CLK => clk, SN => 
                           n387, Q => reg_in_2_port);
   reg_in_regx1x : DFFSNQ_X1 port map( D => Plaintext(1), CLK => clk, SN => 
                           n386, Q => reg_in_1_port);
   reg_in_regx0x : DFFSNQ_X1 port map( D => Plaintext(0), CLK => clk, SN => 
                           n385, Q => reg_in_0_port);
   reg_key_regx191x : DFFSNQ_X1 port map( D => Key(191), CLK => clk, SN => n384
                           , Q => reg_key_191_port);
   reg_key_regx190x : DFFSNQ_X1 port map( D => Key(190), CLK => clk, SN => n383
                           , Q => reg_key_190_port);
   reg_key_regx189x : DFFSNQ_X1 port map( D => Key(189), CLK => clk, SN => n382
                           , Q => reg_key_189_port);
   reg_key_regx188x : DFFSNQ_X1 port map( D => Key(188), CLK => clk, SN => n381
                           , Q => reg_key_188_port);
   reg_key_regx187x : DFFSNQ_X1 port map( D => Key(187), CLK => clk, SN => n380
                           , Q => reg_key_187_port);
   reg_key_regx186x : DFFSNQ_X1 port map( D => Key(186), CLK => clk, SN => n379
                           , Q => reg_key_186_port);
   reg_key_regx185x : DFFSNQ_X1 port map( D => Key(185), CLK => clk, SN => n378
                           , Q => reg_key_185_port);
   reg_key_regx184x : DFFSNQ_X1 port map( D => Key(184), CLK => clk, SN => n377
                           , Q => reg_key_184_port);
   reg_key_regx183x : DFFSNQ_X1 port map( D => Key(183), CLK => clk, SN => n376
                           , Q => reg_key_183_port);
   reg_key_regx182x : DFFSNQ_X1 port map( D => Key(182), CLK => clk, SN => n375
                           , Q => reg_key_182_port);
   reg_key_regx181x : DFFSNQ_X1 port map( D => Key(181), CLK => clk, SN => n374
                           , Q => reg_key_181_port);
   reg_key_regx180x : DFFSNQ_X1 port map( D => Key(180), CLK => clk, SN => n373
                           , Q => reg_key_180_port);
   reg_key_regx179x : DFFSNQ_X1 port map( D => Key(179), CLK => clk, SN => n372
                           , Q => reg_key_179_port);
   reg_key_regx178x : DFFSNQ_X1 port map( D => Key(178), CLK => clk, SN => n371
                           , Q => reg_key_178_port);
   reg_key_regx177x : DFFSNQ_X1 port map( D => Key(177), CLK => clk, SN => n370
                           , Q => reg_key_177_port);
   reg_key_regx176x : DFFSNQ_X1 port map( D => Key(176), CLK => clk, SN => n369
                           , Q => reg_key_176_port);
   reg_key_regx175x : DFFSNQ_X1 port map( D => Key(175), CLK => clk, SN => n368
                           , Q => reg_key_175_port);
   reg_key_regx174x : DFFSNQ_X1 port map( D => Key(174), CLK => clk, SN => n367
                           , Q => reg_key_174_port);
   reg_key_regx173x : DFFSNQ_X1 port map( D => Key(173), CLK => clk, SN => n366
                           , Q => reg_key_173_port);
   reg_key_regx172x : DFFSNQ_X1 port map( D => Key(172), CLK => clk, SN => n365
                           , Q => reg_key_172_port);
   reg_key_regx171x : DFFSNQ_X1 port map( D => Key(171), CLK => clk, SN => n364
                           , Q => reg_key_171_port);
   reg_key_regx170x : DFFSNQ_X1 port map( D => Key(170), CLK => clk, SN => n363
                           , Q => reg_key_170_port);
   reg_key_regx169x : DFFSNQ_X1 port map( D => Key(169), CLK => clk, SN => n362
                           , Q => reg_key_169_port);
   reg_key_regx168x : DFFSNQ_X1 port map( D => Key(168), CLK => clk, SN => n361
                           , Q => reg_key_168_port);
   reg_key_regx167x : DFFSNQ_X1 port map( D => Key(167), CLK => clk, SN => n360
                           , Q => reg_key_167_port);
   reg_key_regx166x : DFFSNQ_X1 port map( D => Key(166), CLK => clk, SN => n359
                           , Q => reg_key_166_port);
   reg_key_regx165x : DFFSNQ_X1 port map( D => Key(165), CLK => clk, SN => n358
                           , Q => reg_key_165_port);
   reg_key_regx164x : DFFSNQ_X1 port map( D => Key(164), CLK => clk, SN => n357
                           , Q => reg_key_164_port);
   reg_key_regx163x : DFFSNQ_X1 port map( D => Key(163), CLK => clk, SN => n356
                           , Q => reg_key_163_port);
   reg_key_regx162x : DFFSNQ_X1 port map( D => Key(162), CLK => clk, SN => n355
                           , Q => reg_key_162_port);
   reg_key_regx161x : DFFSNQ_X1 port map( D => Key(161), CLK => clk, SN => n354
                           , Q => reg_key_161_port);
   reg_key_regx160x : DFFSNQ_X1 port map( D => Key(160), CLK => clk, SN => n353
                           , Q => reg_key_160_port);
   reg_key_regx159x : DFFSNQ_X1 port map( D => Key(159), CLK => clk, SN => n352
                           , Q => reg_key_159_port);
   reg_key_regx158x : DFFSNQ_X1 port map( D => Key(158), CLK => clk, SN => n351
                           , Q => reg_key_158_port);
   reg_key_regx157x : DFFSNQ_X1 port map( D => Key(157), CLK => clk, SN => n350
                           , Q => reg_key_157_port);
   reg_key_regx156x : DFFSNQ_X1 port map( D => Key(156), CLK => clk, SN => n349
                           , Q => reg_key_156_port);
   reg_key_regx155x : DFFSNQ_X1 port map( D => Key(155), CLK => clk, SN => n348
                           , Q => reg_key_155_port);
   reg_key_regx154x : DFFSNQ_X1 port map( D => Key(154), CLK => clk, SN => n347
                           , Q => reg_key_154_port);
   reg_key_regx153x : DFFSNQ_X1 port map( D => Key(153), CLK => clk, SN => n346
                           , Q => reg_key_153_port);
   reg_key_regx152x : DFFSNQ_X1 port map( D => Key(152), CLK => clk, SN => n345
                           , Q => reg_key_152_port);
   reg_key_regx151x : DFFSNQ_X1 port map( D => Key(151), CLK => clk, SN => n344
                           , Q => reg_key_151_port);
   reg_key_regx150x : DFFSNQ_X1 port map( D => Key(150), CLK => clk, SN => n343
                           , Q => reg_key_150_port);
   reg_key_regx149x : DFFSNQ_X1 port map( D => Key(149), CLK => clk, SN => n342
                           , Q => reg_key_149_port);
   reg_key_regx148x : DFFSNQ_X1 port map( D => Key(148), CLK => clk, SN => n341
                           , Q => reg_key_148_port);
   reg_key_regx147x : DFFSNQ_X1 port map( D => Key(147), CLK => clk, SN => n340
                           , Q => reg_key_147_port);
   reg_key_regx146x : DFFSNQ_X1 port map( D => Key(146), CLK => clk, SN => n339
                           , Q => reg_key_146_port);
   reg_key_regx145x : DFFSNQ_X1 port map( D => Key(145), CLK => clk, SN => n338
                           , Q => reg_key_145_port);
   reg_key_regx144x : DFFSNQ_X1 port map( D => Key(144), CLK => clk, SN => n337
                           , Q => reg_key_144_port);
   reg_key_regx143x : DFFSNQ_X1 port map( D => Key(143), CLK => clk, SN => n336
                           , Q => reg_key_143_port);
   reg_key_regx142x : DFFSNQ_X1 port map( D => Key(142), CLK => clk, SN => n335
                           , Q => reg_key_142_port);
   reg_key_regx141x : DFFSNQ_X1 port map( D => Key(141), CLK => clk, SN => n334
                           , Q => reg_key_141_port);
   reg_key_regx140x : DFFSNQ_X1 port map( D => Key(140), CLK => clk, SN => n333
                           , Q => reg_key_140_port);
   reg_key_regx139x : DFFSNQ_X1 port map( D => Key(139), CLK => clk, SN => n332
                           , Q => reg_key_139_port);
   reg_key_regx138x : DFFSNQ_X1 port map( D => Key(138), CLK => clk, SN => n331
                           , Q => reg_key_138_port);
   reg_key_regx137x : DFFSNQ_X1 port map( D => Key(137), CLK => clk, SN => n330
                           , Q => reg_key_137_port);
   reg_key_regx136x : DFFSNQ_X1 port map( D => Key(136), CLK => clk, SN => n329
                           , Q => reg_key_136_port);
   reg_key_regx135x : DFFSNQ_X1 port map( D => Key(135), CLK => clk, SN => n328
                           , Q => reg_key_135_port);
   reg_key_regx134x : DFFSNQ_X1 port map( D => Key(134), CLK => clk, SN => n327
                           , Q => reg_key_134_port);
   reg_key_regx133x : DFFSNQ_X1 port map( D => Key(133), CLK => clk, SN => n326
                           , Q => reg_key_133_port);
   reg_key_regx132x : DFFSNQ_X1 port map( D => Key(132), CLK => clk, SN => n325
                           , Q => reg_key_132_port);
   reg_key_regx131x : DFFSNQ_X1 port map( D => Key(131), CLK => clk, SN => n324
                           , Q => reg_key_131_port);
   reg_key_regx130x : DFFSNQ_X1 port map( D => Key(130), CLK => clk, SN => n323
                           , Q => reg_key_130_port);
   reg_key_regx129x : DFFSNQ_X1 port map( D => Key(129), CLK => clk, SN => n322
                           , Q => reg_key_129_port);
   reg_key_regx128x : DFFSNQ_X1 port map( D => Key(128), CLK => clk, SN => n321
                           , Q => reg_key_128_port);
   reg_key_regx127x : DFFSNQ_X1 port map( D => Key(127), CLK => clk, SN => n320
                           , Q => reg_key_127_port);
   reg_key_regx126x : DFFSNQ_X1 port map( D => Key(126), CLK => clk, SN => n319
                           , Q => reg_key_126_port);
   reg_key_regx125x : DFFSNQ_X1 port map( D => Key(125), CLK => clk, SN => n318
                           , Q => reg_key_125_port);
   reg_key_regx124x : DFFSNQ_X1 port map( D => Key(124), CLK => clk, SN => n317
                           , Q => reg_key_124_port);
   reg_key_regx123x : DFFSNQ_X1 port map( D => Key(123), CLK => clk, SN => n316
                           , Q => reg_key_123_port);
   reg_key_regx122x : DFFSNQ_X1 port map( D => Key(122), CLK => clk, SN => n315
                           , Q => reg_key_122_port);
   reg_key_regx121x : DFFSNQ_X1 port map( D => Key(121), CLK => clk, SN => n314
                           , Q => reg_key_121_port);
   reg_key_regx120x : DFFSNQ_X1 port map( D => Key(120), CLK => clk, SN => n313
                           , Q => reg_key_120_port);
   reg_key_regx119x : DFFSNQ_X1 port map( D => Key(119), CLK => clk, SN => n312
                           , Q => reg_key_119_port);
   reg_key_regx118x : DFFSNQ_X1 port map( D => Key(118), CLK => clk, SN => n311
                           , Q => reg_key_118_port);
   reg_key_regx117x : DFFSNQ_X1 port map( D => Key(117), CLK => clk, SN => n310
                           , Q => reg_key_117_port);
   reg_key_regx116x : DFFSNQ_X1 port map( D => Key(116), CLK => clk, SN => n309
                           , Q => reg_key_116_port);
   reg_key_regx115x : DFFSNQ_X1 port map( D => Key(115), CLK => clk, SN => n308
                           , Q => reg_key_115_port);
   reg_key_regx114x : DFFSNQ_X1 port map( D => Key(114), CLK => clk, SN => n307
                           , Q => reg_key_114_port);
   reg_key_regx113x : DFFSNQ_X1 port map( D => Key(113), CLK => clk, SN => n306
                           , Q => reg_key_113_port);
   reg_key_regx112x : DFFSNQ_X1 port map( D => Key(112), CLK => clk, SN => n305
                           , Q => reg_key_112_port);
   reg_key_regx111x : DFFSNQ_X1 port map( D => Key(111), CLK => clk, SN => n304
                           , Q => reg_key_111_port);
   reg_key_regx110x : DFFSNQ_X1 port map( D => Key(110), CLK => clk, SN => n303
                           , Q => reg_key_110_port);
   reg_key_regx109x : DFFSNQ_X1 port map( D => Key(109), CLK => clk, SN => n302
                           , Q => reg_key_109_port);
   reg_key_regx108x : DFFSNQ_X1 port map( D => Key(108), CLK => clk, SN => n301
                           , Q => reg_key_108_port);
   reg_key_regx107x : DFFSNQ_X1 port map( D => Key(107), CLK => clk, SN => n300
                           , Q => reg_key_107_port);
   reg_key_regx106x : DFFSNQ_X1 port map( D => Key(106), CLK => clk, SN => n299
                           , Q => reg_key_106_port);
   reg_key_regx105x : DFFSNQ_X1 port map( D => Key(105), CLK => clk, SN => n298
                           , Q => reg_key_105_port);
   reg_key_regx104x : DFFSNQ_X1 port map( D => Key(104), CLK => clk, SN => n297
                           , Q => reg_key_104_port);
   reg_key_regx103x : DFFSNQ_X1 port map( D => Key(103), CLK => clk, SN => n296
                           , Q => reg_key_103_port);
   reg_key_regx102x : DFFSNQ_X1 port map( D => Key(102), CLK => clk, SN => n295
                           , Q => reg_key_102_port);
   reg_key_regx101x : DFFSNQ_X1 port map( D => Key(101), CLK => clk, SN => n294
                           , Q => reg_key_101_port);
   reg_key_regx100x : DFFSNQ_X1 port map( D => Key(100), CLK => clk, SN => n293
                           , Q => reg_key_100_port);
   reg_key_regx99x : DFFSNQ_X1 port map( D => Key(99), CLK => clk, SN => n292, 
                           Q => reg_key_99_port);
   reg_key_regx98x : DFFSNQ_X1 port map( D => Key(98), CLK => clk, SN => n291, 
                           Q => reg_key_98_port);
   reg_key_regx97x : DFFSNQ_X1 port map( D => Key(97), CLK => clk, SN => n290, 
                           Q => reg_key_97_port);
   reg_key_regx96x : DFFSNQ_X1 port map( D => Key(96), CLK => clk, SN => n289, 
                           Q => reg_key_96_port);
   reg_key_regx95x : DFFSNQ_X1 port map( D => Key(95), CLK => clk, SN => n288, 
                           Q => reg_key_95_port);
   reg_key_regx94x : DFFSNQ_X1 port map( D => Key(94), CLK => clk, SN => n287, 
                           Q => reg_key_94_port);
   reg_key_regx93x : DFFSNQ_X1 port map( D => Key(93), CLK => clk, SN => n286, 
                           Q => reg_key_93_port);
   reg_key_regx92x : DFFSNQ_X1 port map( D => Key(92), CLK => clk, SN => n285, 
                           Q => reg_key_92_port);
   reg_key_regx91x : DFFSNQ_X1 port map( D => Key(91), CLK => clk, SN => n284, 
                           Q => reg_key_91_port);
   reg_key_regx90x : DFFSNQ_X1 port map( D => Key(90), CLK => clk, SN => n283, 
                           Q => reg_key_90_port);
   reg_key_regx89x : DFFSNQ_X1 port map( D => Key(89), CLK => clk, SN => n282, 
                           Q => reg_key_89_port);
   reg_key_regx88x : DFFSNQ_X1 port map( D => Key(88), CLK => clk, SN => n281, 
                           Q => reg_key_88_port);
   reg_key_regx87x : DFFSNQ_X1 port map( D => Key(87), CLK => clk, SN => n280, 
                           Q => reg_key_87_port);
   reg_key_regx86x : DFFSNQ_X1 port map( D => Key(86), CLK => clk, SN => n279, 
                           Q => reg_key_86_port);
   reg_key_regx85x : DFFSNQ_X1 port map( D => Key(85), CLK => clk, SN => n278, 
                           Q => reg_key_85_port);
   reg_key_regx84x : DFFSNQ_X1 port map( D => Key(84), CLK => clk, SN => n277, 
                           Q => reg_key_84_port);
   reg_key_regx83x : DFFSNQ_X1 port map( D => Key(83), CLK => clk, SN => n276, 
                           Q => reg_key_83_port);
   reg_key_regx82x : DFFSNQ_X1 port map( D => Key(82), CLK => clk, SN => n275, 
                           Q => reg_key_82_port);
   reg_key_regx81x : DFFSNQ_X1 port map( D => Key(81), CLK => clk, SN => n274, 
                           Q => reg_key_81_port);
   reg_key_regx80x : DFFSNQ_X1 port map( D => Key(80), CLK => clk, SN => n273, 
                           Q => reg_key_80_port);
   reg_key_regx79x : DFFSNQ_X1 port map( D => Key(79), CLK => clk, SN => n272, 
                           Q => reg_key_79_port);
   reg_key_regx78x : DFFSNQ_X1 port map( D => Key(78), CLK => clk, SN => n271, 
                           Q => reg_key_78_port);
   reg_key_regx77x : DFFSNQ_X1 port map( D => Key(77), CLK => clk, SN => n270, 
                           Q => reg_key_77_port);
   reg_key_regx76x : DFFSNQ_X1 port map( D => Key(76), CLK => clk, SN => n269, 
                           Q => reg_key_76_port);
   reg_key_regx75x : DFFSNQ_X1 port map( D => Key(75), CLK => clk, SN => n268, 
                           Q => reg_key_75_port);
   reg_key_regx74x : DFFSNQ_X1 port map( D => Key(74), CLK => clk, SN => n267, 
                           Q => reg_key_74_port);
   reg_key_regx73x : DFFSNQ_X1 port map( D => Key(73), CLK => clk, SN => n266, 
                           Q => reg_key_73_port);
   reg_key_regx72x : DFFSNQ_X1 port map( D => Key(72), CLK => clk, SN => n265, 
                           Q => reg_key_72_port);
   reg_key_regx71x : DFFSNQ_X1 port map( D => Key(71), CLK => clk, SN => n264, 
                           Q => reg_key_71_port);
   reg_key_regx70x : DFFSNQ_X1 port map( D => Key(70), CLK => clk, SN => n263, 
                           Q => reg_key_70_port);
   reg_key_regx69x : DFFSNQ_X1 port map( D => Key(69), CLK => clk, SN => n262, 
                           Q => reg_key_69_port);
   reg_key_regx68x : DFFSNQ_X1 port map( D => Key(68), CLK => clk, SN => n261, 
                           Q => reg_key_68_port);
   reg_key_regx67x : DFFSNQ_X1 port map( D => Key(67), CLK => clk, SN => n260, 
                           Q => reg_key_67_port);
   reg_key_regx66x : DFFSNQ_X1 port map( D => Key(66), CLK => clk, SN => n259, 
                           Q => reg_key_66_port);
   reg_key_regx65x : DFFSNQ_X1 port map( D => Key(65), CLK => clk, SN => n258, 
                           Q => reg_key_65_port);
   reg_key_regx64x : DFFSNQ_X1 port map( D => Key(64), CLK => clk, SN => n257, 
                           Q => reg_key_64_port);
   reg_key_regx63x : DFFSNQ_X1 port map( D => Key(63), CLK => clk, SN => n256, 
                           Q => reg_key_63_port);
   reg_key_regx62x : DFFSNQ_X1 port map( D => Key(62), CLK => clk, SN => n255, 
                           Q => reg_key_62_port);
   reg_key_regx61x : DFFSNQ_X1 port map( D => Key(61), CLK => clk, SN => n254, 
                           Q => reg_key_61_port);
   reg_key_regx60x : DFFSNQ_X1 port map( D => Key(60), CLK => clk, SN => n253, 
                           Q => reg_key_60_port);
   reg_key_regx59x : DFFSNQ_X1 port map( D => Key(59), CLK => clk, SN => n252, 
                           Q => reg_key_59_port);
   reg_key_regx58x : DFFSNQ_X1 port map( D => Key(58), CLK => clk, SN => n251, 
                           Q => reg_key_58_port);
   reg_key_regx57x : DFFSNQ_X1 port map( D => Key(57), CLK => clk, SN => n250, 
                           Q => reg_key_57_port);
   reg_key_regx56x : DFFSNQ_X1 port map( D => Key(56), CLK => clk, SN => n249, 
                           Q => reg_key_56_port);
   reg_key_regx55x : DFFSNQ_X1 port map( D => Key(55), CLK => clk, SN => n248, 
                           Q => reg_key_55_port);
   reg_key_regx54x : DFFSNQ_X1 port map( D => Key(54), CLK => clk, SN => n247, 
                           Q => reg_key_54_port);
   reg_key_regx53x : DFFSNQ_X1 port map( D => Key(53), CLK => clk, SN => n246, 
                           Q => reg_key_53_port);
   reg_key_regx52x : DFFSNQ_X1 port map( D => Key(52), CLK => clk, SN => n245, 
                           Q => reg_key_52_port);
   reg_key_regx51x : DFFSNQ_X1 port map( D => Key(51), CLK => clk, SN => n244, 
                           Q => reg_key_51_port);
   reg_key_regx50x : DFFSNQ_X1 port map( D => Key(50), CLK => clk, SN => n243, 
                           Q => reg_key_50_port);
   reg_key_regx49x : DFFSNQ_X1 port map( D => Key(49), CLK => clk, SN => n242, 
                           Q => reg_key_49_port);
   reg_key_regx48x : DFFSNQ_X1 port map( D => Key(48), CLK => clk, SN => n241, 
                           Q => reg_key_48_port);
   reg_key_regx47x : DFFSNQ_X1 port map( D => Key(47), CLK => clk, SN => n240, 
                           Q => reg_key_47_port);
   reg_key_regx46x : DFFSNQ_X1 port map( D => Key(46), CLK => clk, SN => n239, 
                           Q => reg_key_46_port);
   reg_key_regx45x : DFFSNQ_X1 port map( D => Key(45), CLK => clk, SN => n238, 
                           Q => reg_key_45_port);
   reg_key_regx44x : DFFSNQ_X1 port map( D => Key(44), CLK => clk, SN => n237, 
                           Q => reg_key_44_port);
   reg_key_regx43x : DFFSNQ_X1 port map( D => Key(43), CLK => clk, SN => n236, 
                           Q => reg_key_43_port);
   reg_key_regx42x : DFFSNQ_X1 port map( D => Key(42), CLK => clk, SN => n235, 
                           Q => reg_key_42_port);
   reg_key_regx41x : DFFSNQ_X1 port map( D => Key(41), CLK => clk, SN => n234, 
                           Q => reg_key_41_port);
   reg_key_regx40x : DFFSNQ_X1 port map( D => Key(40), CLK => clk, SN => n233, 
                           Q => reg_key_40_port);
   reg_key_regx39x : DFFSNQ_X1 port map( D => Key(39), CLK => clk, SN => n232, 
                           Q => reg_key_39_port);
   reg_key_regx38x : DFFSNQ_X1 port map( D => Key(38), CLK => clk, SN => n231, 
                           Q => reg_key_38_port);
   reg_key_regx37x : DFFSNQ_X1 port map( D => Key(37), CLK => clk, SN => n230, 
                           Q => reg_key_37_port);
   reg_key_regx36x : DFFSNQ_X1 port map( D => Key(36), CLK => clk, SN => n229, 
                           Q => reg_key_36_port);
   reg_key_regx35x : DFFSNQ_X1 port map( D => Key(35), CLK => clk, SN => n228, 
                           Q => reg_key_35_port);
   reg_key_regx34x : DFFSNQ_X1 port map( D => Key(34), CLK => clk, SN => n227, 
                           Q => reg_key_34_port);
   reg_key_regx33x : DFFSNQ_X1 port map( D => Key(33), CLK => clk, SN => n226, 
                           Q => reg_key_33_port);
   reg_key_regx32x : DFFSNQ_X1 port map( D => Key(32), CLK => clk, SN => n225, 
                           Q => reg_key_32_port);
   reg_key_regx31x : DFFSNQ_X1 port map( D => Key(31), CLK => clk, SN => n224, 
                           Q => reg_key_31_port);
   reg_key_regx30x : DFFSNQ_X1 port map( D => Key(30), CLK => clk, SN => n223, 
                           Q => reg_key_30_port);
   reg_key_regx29x : DFFSNQ_X1 port map( D => Key(29), CLK => clk, SN => n222, 
                           Q => reg_key_29_port);
   reg_key_regx28x : DFFSNQ_X1 port map( D => Key(28), CLK => clk, SN => n221, 
                           Q => reg_key_28_port);
   reg_key_regx27x : DFFSNQ_X1 port map( D => Key(27), CLK => clk, SN => n220, 
                           Q => reg_key_27_port);
   reg_key_regx26x : DFFSNQ_X1 port map( D => Key(26), CLK => clk, SN => n219, 
                           Q => reg_key_26_port);
   reg_key_regx25x : DFFSNQ_X1 port map( D => Key(25), CLK => clk, SN => n218, 
                           Q => reg_key_25_port);
   reg_key_regx24x : DFFSNQ_X1 port map( D => Key(24), CLK => clk, SN => n217, 
                           Q => reg_key_24_port);
   reg_key_regx23x : DFFSNQ_X1 port map( D => Key(23), CLK => clk, SN => n216, 
                           Q => reg_key_23_port);
   reg_key_regx22x : DFFSNQ_X1 port map( D => Key(22), CLK => clk, SN => n215, 
                           Q => reg_key_22_port);
   reg_key_regx21x : DFFSNQ_X1 port map( D => Key(21), CLK => clk, SN => n214, 
                           Q => reg_key_21_port);
   reg_key_regx20x : DFFSNQ_X1 port map( D => Key(20), CLK => clk, SN => n213, 
                           Q => reg_key_20_port);
   reg_key_regx19x : DFFSNQ_X1 port map( D => Key(19), CLK => clk, SN => n212, 
                           Q => reg_key_19_port);
   reg_key_regx18x : DFFSNQ_X1 port map( D => Key(18), CLK => clk, SN => n211, 
                           Q => reg_key_18_port);
   reg_key_regx17x : DFFSNQ_X1 port map( D => Key(17), CLK => clk, SN => n210, 
                           Q => reg_key_17_port);
   reg_key_regx16x : DFFSNQ_X1 port map( D => Key(16), CLK => clk, SN => n209, 
                           Q => reg_key_16_port);
   reg_key_regx15x : DFFSNQ_X1 port map( D => Key(15), CLK => clk, SN => n208, 
                           Q => reg_key_15_port);
   reg_key_regx14x : DFFSNQ_X1 port map( D => Key(14), CLK => clk, SN => n207, 
                           Q => reg_key_14_port);
   reg_key_regx13x : DFFSNQ_X1 port map( D => Key(13), CLK => clk, SN => n206, 
                           Q => reg_key_13_port);
   reg_key_regx12x : DFFSNQ_X1 port map( D => Key(12), CLK => clk, SN => n205, 
                           Q => reg_key_12_port);
   reg_key_regx10x : DFFSNQ_X1 port map( D => Key(10), CLK => clk, SN => n203, 
                           Q => reg_key_10_port);
   reg_key_regx9x : DFFSNQ_X1 port map( D => Key(9), CLK => clk, SN => n202, Q 
                           => reg_key_9_port);
   reg_key_regx8x : DFFSNQ_X1 port map( D => Key(8), CLK => clk, SN => n201, Q 
                           => reg_key_8_port);
   reg_key_regx7x : DFFSNQ_X1 port map( D => Key(7), CLK => clk, SN => n200, Q 
                           => reg_key_7_port);
   reg_key_regx6x : DFFSNQ_X1 port map( D => Key(6), CLK => clk, SN => n199, Q 
                           => reg_key_6_port);
   reg_key_regx5x : DFFSNQ_X1 port map( D => Key(5), CLK => clk, SN => n198, Q 
                           => reg_key_5_port);
   reg_key_regx4x : DFFSNQ_X1 port map( D => Key(4), CLK => clk, SN => n197, Q 
                           => reg_key_4_port);
   reg_key_regx3x : DFFSNQ_X1 port map( D => Key(3), CLK => clk, SN => n196, Q 
                           => reg_key_3_port);
   reg_key_regx2x : DFFSNQ_X1 port map( D => Key(2), CLK => clk, SN => n195, Q 
                           => reg_key_2_port);
   reg_key_regx1x : DFFSNQ_X1 port map( D => Key(1), CLK => clk, SN => n194, Q 
                           => reg_key_1_port);
   reg_key_regx0x : DFFSNQ_X1 port map( D => Key(0), CLK => clk, SN => n193, Q 
                           => reg_key_0_port);
   Ciphertext_regx190x : DFFSNQ_X1 port map( D => reg_out_190_port, CLK => clk,
                           SN => n191, Q => Ciphertext(190));
   Ciphertext_regx186x : DFFSNQ_X1 port map( D => reg_out_186_port, CLK => clk,
                           SN => n187, Q => Ciphertext(186));
   Ciphertext_regx182x : DFFSNQ_X1 port map( D => reg_out_182_port, CLK => clk,
                           SN => n183, Q => Ciphertext(182));
   Ciphertext_regx181x : DFFSNQ_X1 port map( D => reg_out_181_port, CLK => clk,
                           SN => n182, Q => Ciphertext(181));
   Ciphertext_regx180x : DFFSNQ_X1 port map( D => reg_out_180_port, CLK => clk,
                           SN => n181, Q => Ciphertext(180));
   Ciphertext_regx179x : DFFSNQ_X1 port map( D => reg_out_179_port, CLK => clk,
                           SN => n180, Q => Ciphertext(179));
   Ciphertext_regx176x : DFFSNQ_X1 port map( D => reg_out_176_port, CLK => clk,
                           SN => n177, Q => Ciphertext(176));
   Ciphertext_regx175x : DFFSNQ_X1 port map( D => reg_out_175_port, CLK => clk,
                           SN => n176, Q => Ciphertext(175));
   Ciphertext_regx173x : DFFSNQ_X1 port map( D => reg_out_173_port, CLK => clk,
                           SN => n174, Q => Ciphertext(173));
   Ciphertext_regx171x : DFFSNQ_X1 port map( D => reg_out_171_port, CLK => clk,
                           SN => n172, Q => Ciphertext(171));
   Ciphertext_regx169x : DFFSNQ_X1 port map( D => reg_out_169_port, CLK => clk,
                           SN => n170, Q => Ciphertext(169));
   Ciphertext_regx167x : DFFSNQ_X1 port map( D => reg_out_167_port, CLK => clk,
                           SN => n168, Q => Ciphertext(167));
   Ciphertext_regx166x : DFFSNQ_X1 port map( D => reg_out_166_port, CLK => clk,
                           SN => n167, Q => Ciphertext(166));
   Ciphertext_regx164x : DFFSNQ_X1 port map( D => reg_out_164_port, CLK => clk,
                           SN => n165, Q => Ciphertext(164));
   Ciphertext_regx163x : DFFSNQ_X1 port map( D => reg_out_163_port, CLK => clk,
                           SN => n164, Q => Ciphertext(163));
   Ciphertext_regx161x : DFFSNQ_X1 port map( D => reg_out_161_port, CLK => clk,
                           SN => n162, Q => Ciphertext(161));
   Ciphertext_regx160x : DFFSNQ_X1 port map( D => reg_out_160_port, CLK => clk,
                           SN => n161, Q => Ciphertext(160));
   Ciphertext_regx157x : DFFSNQ_X1 port map( D => reg_out_157_port, CLK => clk,
                           SN => n158, Q => Ciphertext(157));
   Ciphertext_regx156x : DFFSNQ_X1 port map( D => reg_out_156_port, CLK => clk,
                           SN => n157, Q => Ciphertext(156));
   Ciphertext_regx154x : DFFSNQ_X1 port map( D => reg_out_154_port, CLK => clk,
                           SN => n155, Q => Ciphertext(154));
   Ciphertext_regx153x : DFFSNQ_X1 port map( D => reg_out_153_port, CLK => clk,
                           SN => n154, Q => Ciphertext(153));
   Ciphertext_regx152x : DFFSNQ_X1 port map( D => reg_out_152_port, CLK => clk,
                           SN => n153, Q => Ciphertext(152));
   Ciphertext_regx150x : DFFSNQ_X1 port map( D => reg_out_150_port, CLK => clk,
                           SN => n151, Q => Ciphertext(150));
   Ciphertext_regx149x : DFFSNQ_X1 port map( D => reg_out_149_port, CLK => clk,
                           SN => n150, Q => Ciphertext(149));
   Ciphertext_regx147x : DFFSNQ_X1 port map( D => reg_out_147_port, CLK => clk,
                           SN => n148, Q => Ciphertext(147));
   Ciphertext_regx146x : DFFSNQ_X1 port map( D => reg_out_146_port, CLK => clk,
                           SN => n147, Q => Ciphertext(146));
   Ciphertext_regx145x : DFFSNQ_X1 port map( D => reg_out_145_port, CLK => clk,
                           SN => n146, Q => Ciphertext(145));
   Ciphertext_regx144x : DFFSNQ_X1 port map( D => reg_out_144_port, CLK => clk,
                           SN => n145, Q => Ciphertext(144));
   Ciphertext_regx137x : DFFSNQ_X1 port map( D => reg_out_137_port, CLK => clk,
                           SN => n138, Q => Ciphertext(137));
   Ciphertext_regx136x : DFFSNQ_X1 port map( D => reg_out_136_port, CLK => clk,
                           SN => n137, Q => Ciphertext(136));
   Ciphertext_regx135x : DFFSNQ_X1 port map( D => reg_out_135_port, CLK => clk,
                           SN => n136, Q => Ciphertext(135));
   Ciphertext_regx132x : DFFSNQ_X1 port map( D => reg_out_132_port, CLK => clk,
                           SN => n133, Q => Ciphertext(132));
   Ciphertext_regx130x : DFFSNQ_X1 port map( D => reg_out_130_port, CLK => clk,
                           SN => n131, Q => Ciphertext(130));
   Ciphertext_regx125x : DFFSNQ_X1 port map( D => reg_out_125_port, CLK => clk,
                           SN => n126, Q => Ciphertext(125));
   Ciphertext_regx123x : DFFSNQ_X1 port map( D => reg_out_123_port, CLK => clk,
                           SN => n124, Q => Ciphertext(123));
   Ciphertext_regx122x : DFFSNQ_X1 port map( D => reg_out_122_port, CLK => clk,
                           SN => n123, Q => Ciphertext(122));
   Ciphertext_regx121x : DFFSNQ_X1 port map( D => reg_out_121_port, CLK => clk,
                           SN => n122, Q => Ciphertext(121));
   Ciphertext_regx118x : DFFSNQ_X1 port map( D => reg_out_118_port, CLK => clk,
                           SN => n119, Q => Ciphertext(118));
   Ciphertext_regx116x : DFFSNQ_X1 port map( D => reg_out_116_port, CLK => clk,
                           SN => n117, Q => Ciphertext(116));
   Ciphertext_regx115x : DFFSNQ_X1 port map( D => reg_out_115_port, CLK => clk,
                           SN => n116, Q => Ciphertext(115));
   Ciphertext_regx113x : DFFSNQ_X1 port map( D => reg_out_113_port, CLK => clk,
                           SN => n114, Q => Ciphertext(113));
   Ciphertext_regx109x : DFFSNQ_X1 port map( D => reg_out_109_port, CLK => clk,
                           SN => n110, Q => Ciphertext(109));
   Ciphertext_regx108x : DFFSNQ_X1 port map( D => reg_out_108_port, CLK => clk,
                           SN => n109, Q => Ciphertext(108));
   Ciphertext_regx107x : DFFSNQ_X1 port map( D => reg_out_107_port, CLK => clk,
                           SN => n108, Q => Ciphertext(107));
   Ciphertext_regx106x : DFFSNQ_X1 port map( D => reg_out_106_port, CLK => clk,
                           SN => n107, Q => Ciphertext(106));
   Ciphertext_regx103x : DFFSNQ_X1 port map( D => reg_out_103_port, CLK => clk,
                           SN => n104, Q => Ciphertext(103));
   Ciphertext_regx102x : DFFSNQ_X1 port map( D => reg_out_102_port, CLK => clk,
                           SN => n103, Q => Ciphertext(102));
   Ciphertext_regx101x : DFFSNQ_X1 port map( D => reg_out_101_port, CLK => clk,
                           SN => n102, Q => Ciphertext(101));
   Ciphertext_regx97x : DFFSNQ_X1 port map( D => reg_out_97_port, CLK => clk, 
                           SN => n98, Q => Ciphertext(97));
   Ciphertext_regx96x : DFFSNQ_X1 port map( D => reg_out_96_port, CLK => clk, 
                           SN => n97, Q => Ciphertext(96));
   Ciphertext_regx86x : DFFSNQ_X1 port map( D => reg_out_86_port, CLK => clk, 
                           SN => n87, Q => Ciphertext(86));
   Ciphertext_regx85x : DFFSNQ_X1 port map( D => reg_out_85_port, CLK => clk, 
                           SN => n86, Q => Ciphertext(85));
   Ciphertext_regx79x : DFFSNQ_X1 port map( D => reg_out_79_port, CLK => clk, 
                           SN => n80, Q => Ciphertext(79));
   Ciphertext_regx78x : DFFSNQ_X1 port map( D => reg_out_78_port, CLK => clk, 
                           SN => n79, Q => Ciphertext(78));
   Ciphertext_regx77x : DFFSNQ_X1 port map( D => reg_out_77_port, CLK => clk, 
                           SN => n78, Q => Ciphertext(77));
   Ciphertext_regx75x : DFFSNQ_X1 port map( D => reg_out_75_port, CLK => clk, 
                           SN => n76, Q => Ciphertext(75));
   Ciphertext_regx74x : DFFSNQ_X1 port map( D => reg_out_74_port, CLK => clk, 
                           SN => n75, Q => Ciphertext(74));
   Ciphertext_regx73x : DFFSNQ_X1 port map( D => reg_out_73_port, CLK => clk, 
                           SN => n74, Q => Ciphertext(73));
   Ciphertext_regx72x : DFFSNQ_X1 port map( D => reg_out_72_port, CLK => clk, 
                           SN => n73, Q => Ciphertext(72));
   Ciphertext_regx71x : DFFSNQ_X1 port map( D => reg_out_71_port, CLK => clk, 
                           SN => n72, Q => Ciphertext(71));
   Ciphertext_regx68x : DFFSNQ_X1 port map( D => reg_out_68_port, CLK => clk, 
                           SN => n69, Q => Ciphertext(68));
   Ciphertext_regx65x : DFFSNQ_X1 port map( D => reg_out_65_port, CLK => clk, 
                           SN => n66, Q => Ciphertext(65));
   Ciphertext_regx61x : DFFSNQ_X1 port map( D => reg_out_61_port, CLK => clk, 
                           SN => n62, Q => Ciphertext(61));
   Ciphertext_regx58x : DFFSNQ_X1 port map( D => reg_out_58_port, CLK => clk, 
                           SN => n59, Q => Ciphertext(58));
   Ciphertext_regx54x : DFFSNQ_X1 port map( D => reg_out_54_port, CLK => clk, 
                           SN => n55, Q => Ciphertext(54));
   Ciphertext_regx50x : DFFSNQ_X1 port map( D => reg_out_50_port, CLK => clk, 
                           SN => n51, Q => Ciphertext(50));
   Ciphertext_regx49x : DFFSNQ_X1 port map( D => reg_out_49_port, CLK => clk, 
                           SN => n50, Q => Ciphertext(49));
   Ciphertext_regx48x : DFFSNQ_X1 port map( D => reg_out_48_port, CLK => clk, 
                           SN => n49, Q => Ciphertext(48));
   Ciphertext_regx47x : DFFSNQ_X1 port map( D => reg_out_47_port, CLK => clk, 
                           SN => n48, Q => Ciphertext(47));
   Ciphertext_regx44x : DFFSNQ_X1 port map( D => reg_out_44_port, CLK => clk, 
                           SN => n45, Q => Ciphertext(44));
   Ciphertext_regx43x : DFFSNQ_X1 port map( D => reg_out_43_port, CLK => clk, 
                           SN => n44, Q => Ciphertext(43));
   Ciphertext_regx42x : DFFSNQ_X1 port map( D => reg_out_42_port, CLK => clk, 
                           SN => n43, Q => Ciphertext(42));
   Ciphertext_regx40x : DFFSNQ_X1 port map( D => reg_out_40_port, CLK => clk, 
                           SN => n41, Q => Ciphertext(40));
   Ciphertext_regx35x : DFFSNQ_X1 port map( D => reg_out_35_port, CLK => clk, 
                           SN => n36, Q => Ciphertext(35));
   Ciphertext_regx32x : DFFSNQ_X1 port map( D => reg_out_32_port, CLK => clk, 
                           SN => n33, Q => Ciphertext(32));
   Ciphertext_regx31x : DFFSNQ_X1 port map( D => reg_out_31_port, CLK => clk, 
                           SN => n32, Q => Ciphertext(31));
   Ciphertext_regx30x : DFFSNQ_X1 port map( D => reg_out_30_port, CLK => clk, 
                           SN => n31, Q => Ciphertext(30));
   Ciphertext_regx25x : DFFSNQ_X1 port map( D => reg_out_25_port, CLK => clk, 
                           SN => n26, Q => Ciphertext(25));
   Ciphertext_regx24x : DFFSNQ_X1 port map( D => reg_out_24_port, CLK => clk, 
                           SN => n25, Q => Ciphertext(24));
   Ciphertext_regx23x : DFFSNQ_X1 port map( D => reg_out_23_port, CLK => clk, 
                           SN => n24, Q => Ciphertext(23));
   Ciphertext_regx22x : DFFSNQ_X1 port map( D => reg_out_22_port, CLK => clk, 
                           SN => n23, Q => Ciphertext(22));
   Ciphertext_regx18x : DFFSNQ_X1 port map( D => reg_out_18_port, CLK => clk, 
                           SN => n19, Q => Ciphertext(18));
   Ciphertext_regx16x : DFFSNQ_X1 port map( D => reg_out_16_port, CLK => clk, 
                           SN => n17, Q => Ciphertext(16));
   Ciphertext_regx14x : DFFSNQ_X1 port map( D => reg_out_14_port, CLK => clk, 
                           SN => n15, Q => Ciphertext(14));
   Ciphertext_regx9x : DFFSNQ_X1 port map( D => reg_out_9_port, CLK => clk, SN 
                           => n10, Q => Ciphertext(9));
   Ciphertext_regx7x : DFFSNQ_X1 port map( D => reg_out_7_port, CLK => clk, SN 
                           => n8, Q => Ciphertext(7));
   Ciphertext_regx6x : DFFSNQ_X1 port map( D => reg_out_6_port, CLK => clk, SN 
                           => n7, Q => Ciphertext(6));
   Ciphertext_regx1x : DFFSNQ_X1 port map( D => reg_out_1_port, CLK => clk, SN 
                           => n2, Q => Ciphertext(1));
   n2 <= '1';
   n7 <= '1';
   n8 <= '1';
   n10 <= '1';
   n15 <= '1';
   n17 <= '1';
   n19 <= '1';
   n23 <= '1';
   n24 <= '1';
   n25 <= '1';
   n26 <= '1';
   n31 <= '1';
   n32 <= '1';
   n33 <= '1';
   n36 <= '1';
   n41 <= '1';
   n43 <= '1';
   n44 <= '1';
   n45 <= '1';
   n48 <= '1';
   n49 <= '1';
   n50 <= '1';
   n51 <= '1';
   n55 <= '1';
   n59 <= '1';
   n62 <= '1';
   n66 <= '1';
   n69 <= '1';
   n72 <= '1';
   n73 <= '1';
   n74 <= '1';
   n75 <= '1';
   n76 <= '1';
   n78 <= '1';
   n79 <= '1';
   n80 <= '1';
   n86 <= '1';
   n87 <= '1';
   n97 <= '1';
   n98 <= '1';
   n102 <= '1';
   n103 <= '1';
   n104 <= '1';
   n107 <= '1';
   n108 <= '1';
   n109 <= '1';
   n110 <= '1';
   n114 <= '1';
   n116 <= '1';
   n117 <= '1';
   n119 <= '1';
   n122 <= '1';
   n123 <= '1';
   n124 <= '1';
   n126 <= '1';
   n131 <= '1';
   n133 <= '1';
   n136 <= '1';
   n137 <= '1';
   n138 <= '1';
   n145 <= '1';
   n146 <= '1';
   n147 <= '1';
   n148 <= '1';
   n150 <= '1';
   n151 <= '1';
   n153 <= '1';
   n154 <= '1';
   n155 <= '1';
   n157 <= '1';
   n158 <= '1';
   n161 <= '1';
   n162 <= '1';
   n164 <= '1';
   n165 <= '1';
   n167 <= '1';
   n168 <= '1';
   n170 <= '1';
   n172 <= '1';
   n174 <= '1';
   n176 <= '1';
   n177 <= '1';
   n180 <= '1';
   n181 <= '1';
   n182 <= '1';
   n183 <= '1';
   n187 <= '1';
   n191 <= '1';
   n193 <= '1';
   n194 <= '1';
   n195 <= '1';
   n196 <= '1';
   n197 <= '1';
   n198 <= '1';
   n199 <= '1';
   n200 <= '1';
   n201 <= '1';
   n202 <= '1';
   n203 <= '1';
   n205 <= '1';
   n206 <= '1';
   n207 <= '1';
   n208 <= '1';
   n209 <= '1';
   n210 <= '1';
   n211 <= '1';
   n212 <= '1';
   n213 <= '1';
   n214 <= '1';
   n215 <= '1';
   n216 <= '1';
   n217 <= '1';
   n218 <= '1';
   n219 <= '1';
   n220 <= '1';
   n221 <= '1';
   n222 <= '1';
   n223 <= '1';
   n224 <= '1';
   n225 <= '1';
   n226 <= '1';
   n227 <= '1';
   n228 <= '1';
   n229 <= '1';
   n230 <= '1';
   n231 <= '1';
   n232 <= '1';
   n233 <= '1';
   n234 <= '1';
   n235 <= '1';
   n236 <= '1';
   n237 <= '1';
   n238 <= '1';
   n239 <= '1';
   n240 <= '1';
   n241 <= '1';
   n242 <= '1';
   n243 <= '1';
   n244 <= '1';
   n245 <= '1';
   n246 <= '1';
   n247 <= '1';
   n248 <= '1';
   n249 <= '1';
   n250 <= '1';
   n251 <= '1';
   n252 <= '1';
   n253 <= '1';
   n254 <= '1';
   n255 <= '1';
   n256 <= '1';
   n257 <= '1';
   n258 <= '1';
   n259 <= '1';
   n260 <= '1';
   n261 <= '1';
   n262 <= '1';
   n263 <= '1';
   n264 <= '1';
   n265 <= '1';
   n266 <= '1';
   n267 <= '1';
   n268 <= '1';
   n269 <= '1';
   n270 <= '1';
   n271 <= '1';
   n272 <= '1';
   n273 <= '1';
   n274 <= '1';
   n275 <= '1';
   n276 <= '1';
   n277 <= '1';
   n278 <= '1';
   n279 <= '1';
   n280 <= '1';
   n281 <= '1';
   n282 <= '1';
   n283 <= '1';
   n284 <= '1';
   n285 <= '1';
   n286 <= '1';
   n287 <= '1';
   n288 <= '1';
   n289 <= '1';
   n290 <= '1';
   n291 <= '1';
   n292 <= '1';
   n293 <= '1';
   n294 <= '1';
   n295 <= '1';
   n296 <= '1';
   n297 <= '1';
   n298 <= '1';
   n299 <= '1';
   n300 <= '1';
   n301 <= '1';
   n302 <= '1';
   n303 <= '1';
   n304 <= '1';
   n305 <= '1';
   n306 <= '1';
   n307 <= '1';
   n308 <= '1';
   n309 <= '1';
   n310 <= '1';
   n311 <= '1';
   n312 <= '1';
   n313 <= '1';
   n314 <= '1';
   n315 <= '1';
   n316 <= '1';
   n317 <= '1';
   n318 <= '1';
   n319 <= '1';
   n320 <= '1';
   n321 <= '1';
   n322 <= '1';
   n323 <= '1';
   n324 <= '1';
   n325 <= '1';
   n326 <= '1';
   n327 <= '1';
   n328 <= '1';
   n329 <= '1';
   n330 <= '1';
   n331 <= '1';
   n332 <= '1';
   n333 <= '1';
   n334 <= '1';
   n335 <= '1';
   n336 <= '1';
   n337 <= '1';
   n338 <= '1';
   n339 <= '1';
   n340 <= '1';
   n341 <= '1';
   n342 <= '1';
   n343 <= '1';
   n344 <= '1';
   n345 <= '1';
   n346 <= '1';
   n347 <= '1';
   n348 <= '1';
   n349 <= '1';
   n350 <= '1';
   n351 <= '1';
   n352 <= '1';
   n353 <= '1';
   n354 <= '1';
   n355 <= '1';
   n356 <= '1';
   n357 <= '1';
   n358 <= '1';
   n359 <= '1';
   n360 <= '1';
   n361 <= '1';
   n362 <= '1';
   n363 <= '1';
   n364 <= '1';
   n365 <= '1';
   n366 <= '1';
   n367 <= '1';
   n368 <= '1';
   n369 <= '1';
   n370 <= '1';
   n371 <= '1';
   n372 <= '1';
   n373 <= '1';
   n374 <= '1';
   n375 <= '1';
   n376 <= '1';
   n377 <= '1';
   n378 <= '1';
   n379 <= '1';
   n380 <= '1';
   n381 <= '1';
   n382 <= '1';
   n383 <= '1';
   n384 <= '1';
   n385 <= '1';
   n386 <= '1';
   n387 <= '1';
   n388 <= '1';
   n389 <= '1';
   n390 <= '1';
   n391 <= '1';
   n392 <= '1';
   n393 <= '1';
   n394 <= '1';
   n395 <= '1';
   n396 <= '1';
   n397 <= '1';
   n398 <= '1';
   n399 <= '1';
   n400 <= '1';
   n401 <= '1';
   n402 <= '1';
   n403 <= '1';
   n404 <= '1';
   n405 <= '1';
   n406 <= '1';
   n407 <= '1';
   n408 <= '1';
   n409 <= '1';
   n410 <= '1';
   n411 <= '1';
   n412 <= '1';
   n413 <= '1';
   n415 <= '1';
   n416 <= '1';
   n417 <= '1';
   n418 <= '1';
   n419 <= '1';
   n420 <= '1';
   n421 <= '1';
   n422 <= '1';
   n423 <= '1';
   n424 <= '1';
   n425 <= '1';
   n426 <= '1';
   n427 <= '1';
   n428 <= '1';
   n429 <= '1';
   n430 <= '1';
   n431 <= '1';
   n432 <= '1';
   n433 <= '1';
   n434 <= '1';
   n435 <= '1';
   n437 <= '1';
   n438 <= '1';
   n439 <= '1';
   n440 <= '1';
   n441 <= '1';
   n442 <= '1';
   n443 <= '1';
   n444 <= '1';
   n445 <= '1';
   n446 <= '1';
   n447 <= '1';
   n448 <= '1';
   n449 <= '1';
   n450 <= '1';
   n451 <= '1';
   n452 <= '1';
   n453 <= '1';
   n454 <= '1';
   n455 <= '1';
   n457 <= '1';
   n458 <= '1';
   n459 <= '1';
   n460 <= '1';
   n461 <= '1';
   n462 <= '1';
   n463 <= '1';
   n464 <= '1';
   n465 <= '1';
   n466 <= '1';
   n467 <= '1';
   n468 <= '1';
   n469 <= '1';
   n470 <= '1';
   n471 <= '1';
   n472 <= '1';
   n473 <= '1';
   n474 <= '1';
   n475 <= '1';
   n476 <= '1';
   n477 <= '1';
   n478 <= '1';
   n479 <= '1';
   n480 <= '1';
   n481 <= '1';
   n482 <= '1';
   n483 <= '1';
   n484 <= '1';
   n485 <= '1';
   n486 <= '1';
   n487 <= '1';
   n488 <= '1';
   n489 <= '1';
   n490 <= '1';
   n491 <= '1';
   n492 <= '1';
   n493 <= '1';
   n494 <= '1';
   n495 <= '1';
   n496 <= '1';
   n497 <= '1';
   n498 <= '1';
   n499 <= '1';
   n500 <= '1';
   n501 <= '1';
   n502 <= '1';
   n503 <= '1';
   n504 <= '1';
   n505 <= '1';
   n506 <= '1';
   n507 <= '1';
   n508 <= '1';
   n509 <= '1';
   n510 <= '1';
   n511 <= '1';
   n512 <= '1';
   n513 <= '1';
   n514 <= '1';
   n515 <= '1';
   n517 <= '1';
   n518 <= '1';
   n519 <= '1';
   n520 <= '1';
   n521 <= '1';
   n522 <= '1';
   n523 <= '1';
   n524 <= '1';
   n525 <= '1';
   n526 <= '1';
   n527 <= '1';
   n528 <= '1';
   n529 <= '1';
   n530 <= '1';
   n531 <= '1';
   n533 <= '1';
   n534 <= '1';
   n535 <= '1';
   n536 <= '1';
   n537 <= '1';
   n538 <= '1';
   n539 <= '1';
   n540 <= '1';
   n541 <= '1';
   n542 <= '1';
   n543 <= '1';
   n544 <= '1';
   n545 <= '1';
   n546 <= '1';
   n547 <= '1';
   n548 <= '1';
   n549 <= '1';
   n550 <= '1';
   n551 <= '1';
   n552 <= '1';
   n553 <= '1';
   n554 <= '1';
   n555 <= '1';
   n556 <= '1';
   n557 <= '1';
   n558 <= '1';
   n559 <= '1';
   n560 <= '1';
   n561 <= '1';
   n562 <= '1';
   n563 <= '1';
   n564 <= '1';
   n565 <= '1';
   n566 <= '1';
   n567 <= '1';
   n568 <= '1';
   n569 <= '1';
   n570 <= '1';
   n571 <= '1';
   n572 <= '1';
   n573 <= '1';
   n574 <= '1';
   n575 <= '1';
   n576 <= '1';
   Ciphertext_regx36x : DFFRNQ_X1 port map( D => reg_out_36_port, CLK => clk, 
                           RN => n652, Q => Ciphertext(36));
   Ciphertext_regx178x : DFFRNQ_X1 port map( D => reg_out_178_port, CLK => clk,
                           RN => n651, Q => Ciphertext(178));
   Ciphertext_regx4x : DFFRNQ_X1 port map( D => reg_out_4_port, CLK => clk, RN 
                           => n650, Q => Ciphertext(4));
   Ciphertext_regx88x : DFFRNQ_X1 port map( D => reg_out_88_port, CLK => clk, 
                           RN => n649, Q => Ciphertext(88));
   Ciphertext_regx34x : DFFRNQ_X1 port map( D => reg_out_34_port, CLK => clk, 
                           RN => n648, Q => Ciphertext(34));
   Ciphertext_regx119x : DFFRNQ_X1 port map( D => reg_out_119_port, CLK => clk,
                           RN => n647, Q => Ciphertext(119));
   Ciphertext_regx39x : DFFRNQ_X1 port map( D => reg_out_39_port, CLK => clk, 
                           RN => n646, Q => Ciphertext(39));
   Ciphertext_regx37x : DFFRNQ_X1 port map( D => reg_out_37_port, CLK => clk, 
                           RN => n645, Q => Ciphertext(37));
   Ciphertext_regx174x : DFFRNQ_X1 port map( D => reg_out_174_port, CLK => clk,
                           RN => n644, Q => Ciphertext(174));
   Ciphertext_regx70x : DFFRNQ_X1 port map( D => reg_out_70_port, CLK => clk, 
                           RN => n643, Q => Ciphertext(70));
   Ciphertext_regx84x : DFFRNQ_X1 port map( D => reg_out_84_port, CLK => clk, 
                           RN => n642, Q => Ciphertext(84));
   Ciphertext_regx143x : DFFRNQ_X1 port map( D => reg_out_143_port, CLK => clk,
                           RN => n641, Q => Ciphertext(143));
   Ciphertext_regx57x : DFFRNQ_X1 port map( D => reg_out_57_port, CLK => clk, 
                           RN => n640, Q => Ciphertext(57));
   Ciphertext_regx46x : DFFRNQ_X1 port map( D => reg_out_46_port, CLK => clk, 
                           RN => n639, Q => Ciphertext(46));
   Ciphertext_regx3x : DFFRNQ_X1 port map( D => reg_out_3_port, CLK => clk, RN 
                           => n638, Q => Ciphertext(3));
   Ciphertext_regx66x : DFFRNQ_X1 port map( D => reg_out_66_port, CLK => clk, 
                           RN => n637, Q => Ciphertext(66));
   Ciphertext_regx170x : DFFRNQ_X1 port map( D => reg_out_170_port, CLK => clk,
                           RN => n636, Q => Ciphertext(170));
   Ciphertext_regx80x : DFFRNQ_X1 port map( D => reg_out_80_port, CLK => clk, 
                           RN => n635, Q => Ciphertext(80));
   Ciphertext_regx98x : DFFRNQ_X1 port map( D => reg_out_98_port, CLK => clk, 
                           RN => n634, Q => Ciphertext(98));
   Ciphertext_regx8x : DFFRNQ_X1 port map( D => reg_out_8_port, CLK => clk, RN 
                           => n633, Q => Ciphertext(8));
   Ciphertext_regx60x : DFFRNQ_X1 port map( D => reg_out_60_port, CLK => clk, 
                           RN => n632, Q => Ciphertext(60));
   Ciphertext_regx55x : DFFRNQ_X1 port map( D => reg_out_55_port, CLK => clk, 
                           RN => n630, Q => Ciphertext(55));
   Ciphertext_regx69x : DFFRNQ_X1 port map( D => reg_out_69_port, CLK => clk, 
                           RN => n629, Q => Ciphertext(69));
   Ciphertext_regx90x : DFFRNQ_X1 port map( D => reg_out_90_port, CLK => clk, 
                           RN => n628, Q => Ciphertext(90));
   Ciphertext_regx142x : DFFRNQ_X1 port map( D => reg_out_142_port, CLK => clk,
                           RN => n627, Q => Ciphertext(142));
   Ciphertext_regx159x : DFFRNQ_X1 port map( D => reg_out_159_port, CLK => clk,
                           RN => n626, Q => Ciphertext(159));
   Ciphertext_regx52x : DFFRNQ_X1 port map( D => reg_out_52_port, CLK => clk, 
                           RN => n625, Q => Ciphertext(52));
   Ciphertext_regx5x : DFFRNQ_X1 port map( D => reg_out_5_port, CLK => clk, RN 
                           => n624, Q => Ciphertext(5));
   Ciphertext_regx27x : DFFRNQ_X1 port map( D => reg_out_27_port, CLK => clk, 
                           RN => n623, Q => Ciphertext(27));
   Ciphertext_regx92x : DFFRNQ_X1 port map( D => reg_out_92_port, CLK => clk, 
                           RN => n622, Q => Ciphertext(92));
   Ciphertext_regx184x : DFFRNQ_X1 port map( D => reg_out_184_port, CLK => clk,
                           RN => n621, Q => Ciphertext(184));
   Ciphertext_regx138x : DFFRNQ_X1 port map( D => reg_out_138_port, CLK => clk,
                           RN => n620, Q => Ciphertext(138));
   Ciphertext_regx11x : DFFRNQ_X1 port map( D => reg_out_11_port, CLK => clk, 
                           RN => n619, Q => Ciphertext(11));
   Ciphertext_regx91x : DFFRNQ_X1 port map( D => reg_out_91_port, CLK => clk, 
                           RN => n618, Q => Ciphertext(91));
   Ciphertext_regx93x : DFFRNQ_X1 port map( D => reg_out_93_port, CLK => clk, 
                           RN => n617, Q => Ciphertext(93));
   Ciphertext_regx126x : DFFRNQ_X1 port map( D => reg_out_126_port, CLK => clk,
                           RN => n616, Q => Ciphertext(126));
   Ciphertext_regx29x : DFFRNQ_X1 port map( D => reg_out_29_port, CLK => clk, 
                           RN => n615, Q => Ciphertext(29));
   Ciphertext_regx38x : DFFRNQ_X1 port map( D => reg_out_38_port, CLK => clk, 
                           RN => n614, Q => Ciphertext(38));
   Ciphertext_regx133x : DFFRNQ_X1 port map( D => reg_out_133_port, CLK => clk,
                           RN => n613, Q => Ciphertext(133));
   Ciphertext_regx19x : DFFRNQ_X1 port map( D => reg_out_19_port, CLK => clk, 
                           RN => n612, Q => Ciphertext(19));
   Ciphertext_regx172x : DFFRNQ_X1 port map( D => reg_out_172_port, CLK => clk,
                           RN => n611, Q => Ciphertext(172));
   Ciphertext_regx177x : DFFRNQ_X1 port map( D => reg_out_177_port, CLK => clk,
                           RN => n610, Q => Ciphertext(177));
   Ciphertext_regx158x : DFFRNQ_X1 port map( D => reg_out_158_port, CLK => clk,
                           RN => n609, Q => Ciphertext(158));
   Ciphertext_regx162x : DFFRNQ_X1 port map( D => reg_out_162_port, CLK => clk,
                           RN => n608, Q => Ciphertext(162));
   Ciphertext_regx111x : DFFRNQ_X1 port map( D => reg_out_111_port, CLK => clk,
                           RN => n607, Q => Ciphertext(111));
   Ciphertext_regx165x : DFFRNQ_X1 port map( D => reg_out_165_port, CLK => clk,
                           RN => n606, Q => Ciphertext(165));
   Ciphertext_regx83x : DFFRNQ_X1 port map( D => reg_out_83_port, CLK => clk, 
                           RN => n605, Q => Ciphertext(83));
   Ciphertext_regx82x : DFFRNQ_X1 port map( D => reg_out_82_port, CLK => clk, 
                           RN => n604, Q => Ciphertext(82));
   Ciphertext_regx2x : DFFRNQ_X1 port map( D => reg_out_2_port, CLK => clk, RN 
                           => n603, Q => Ciphertext(2));
   Ciphertext_regx62x : DFFRNQ_X1 port map( D => reg_out_62_port, CLK => clk, 
                           RN => n602, Q => Ciphertext(62));
   Ciphertext_regx95x : DFFRNQ_X1 port map( D => reg_out_95_port, CLK => clk, 
                           RN => n601, Q => Ciphertext(95));
   Ciphertext_regx140x : DFFRNQ_X1 port map( D => reg_out_140_port, CLK => clk,
                           RN => n599, Q => Ciphertext(140));
   Ciphertext_regx183x : DFFRNQ_X1 port map( D => reg_out_183_port, CLK => clk,
                           RN => n598, Q => Ciphertext(183));
   Ciphertext_regx51x : DFFRNQ_X1 port map( D => reg_out_51_port, CLK => clk, 
                           RN => n597, Q => Ciphertext(51));
   Ciphertext_regx63x : DFFRNQ_X1 port map( D => reg_out_63_port, CLK => clk, 
                           RN => n596, Q => Ciphertext(63));
   Ciphertext_regx185x : DFFRNQ_X1 port map( D => reg_out_185_port, CLK => clk,
                           RN => n595, Q => Ciphertext(185));
   Ciphertext_regx81x : DFFRNQ_X1 port map( D => reg_out_81_port, CLK => clk, 
                           RN => n594, Q => Ciphertext(81));
   Ciphertext_regx26x : DFFRNQ_X1 port map( D => reg_out_26_port, CLK => clk, 
                           RN => n593, Q => Ciphertext(26));
   Ciphertext_regx94x : DFFRNQ_X1 port map( D => reg_out_94_port, CLK => clk, 
                           RN => n592, Q => Ciphertext(94));
   Ciphertext_regx10x : DFFRNQ_X1 port map( D => reg_out_10_port, CLK => clk, 
                           RN => n591, Q => Ciphertext(10));
   Ciphertext_regx87x : DFFRNQ_X1 port map( D => reg_out_87_port, CLK => clk, 
                           RN => n590, Q => Ciphertext(87));
   Ciphertext_regx59x : DFFRNQ_X1 port map( D => reg_out_59_port, CLK => clk, 
                           RN => n589, Q => Ciphertext(59));
   Ciphertext_regx117x : DFFRNQ_X1 port map( D => reg_out_117_port, CLK => clk,
                           RN => n588, Q => Ciphertext(117));
   Ciphertext_regx127x : DFFRNQ_X1 port map( D => reg_out_127_port, CLK => clk,
                           RN => n587, Q => Ciphertext(127));
   Ciphertext_regx15x : DFFRNQ_X1 port map( D => reg_out_15_port, CLK => clk, 
                           RN => n585, Q => Ciphertext(15));
   Ciphertext_regx105x : DFFRNQ_X1 port map( D => reg_out_105_port, CLK => clk,
                           RN => n584, Q => Ciphertext(105));
   Ciphertext_regx131x : DFFRNQ_X1 port map( D => reg_out_131_port, CLK => clk,
                           RN => n583, Q => Ciphertext(131));
   Ciphertext_regx20x : DFFRNQ_X1 port map( D => reg_out_20_port, CLK => clk, 
                           RN => n582, Q => Ciphertext(20));
   Ciphertext_regx21x : DFFRNQ_X1 port map( D => reg_out_21_port, CLK => clk, 
                           RN => n581, Q => Ciphertext(21));
   Ciphertext_regx13x : DFFRNQ_X1 port map( D => reg_out_13_port, CLK => clk, 
                           RN => n580, Q => Ciphertext(13));
   Ciphertext_regx129x : DFFRNQ_X1 port map( D => reg_out_129_port, CLK => clk,
                           RN => n579, Q => Ciphertext(129));
   Ciphertext_regx104x : DFFRNQ_X1 port map( D => reg_out_104_port, CLK => clk,
                           RN => n578, Q => Ciphertext(104));
   Ciphertext_regx33x : DFFRNQ_X1 port map( D => reg_out_33_port, CLK => clk, 
                           RN => n577, Q => Ciphertext(33));
   n577 <= '1';
   n578 <= '1';
   n579 <= '1';
   n580 <= '1';
   n581 <= '1';
   n582 <= '1';
   n583 <= '1';
   n584 <= '1';
   n585 <= '1';
   n587 <= '1';
   n588 <= '1';
   n589 <= '1';
   n590 <= '1';
   n591 <= '1';
   n592 <= '1';
   n593 <= '1';
   n594 <= '1';
   n595 <= '1';
   n596 <= '1';
   n597 <= '1';
   n598 <= '1';
   n599 <= '1';
   n601 <= '1';
   n602 <= '1';
   n603 <= '1';
   n604 <= '1';
   n605 <= '1';
   n606 <= '1';
   n607 <= '1';
   n608 <= '1';
   n609 <= '1';
   n610 <= '1';
   n611 <= '1';
   n612 <= '1';
   n613 <= '1';
   n614 <= '1';
   n615 <= '1';
   n616 <= '1';
   n617 <= '1';
   n618 <= '1';
   n619 <= '1';
   n620 <= '1';
   n621 <= '1';
   n622 <= '1';
   n623 <= '1';
   n624 <= '1';
   n625 <= '1';
   n626 <= '1';
   n627 <= '1';
   n628 <= '1';
   n629 <= '1';
   n630 <= '1';
   n632 <= '1';
   n633 <= '1';
   n634 <= '1';
   n635 <= '1';
   n636 <= '1';
   n637 <= '1';
   n638 <= '1';
   n639 <= '1';
   n640 <= '1';
   n641 <= '1';
   n642 <= '1';
   n643 <= '1';
   n644 <= '1';
   n645 <= '1';
   n646 <= '1';
   n647 <= '1';
   n648 <= '1';
   n649 <= '1';
   n650 <= '1';
   n651 <= '1';
   n652 <= '1';
   Ciphertext_regx110x : DFFRNQ_X1 port map( D => reg_out_110_port, CLK => clk,
                           RN => n671, Q => Ciphertext(110));
   Ciphertext_regx0x : DFFRNQ_X1 port map( D => reg_out_0_port, CLK => clk, RN 
                           => n670, Q => Ciphertext(0));
   Ciphertext_regx45x : DFFRNQ_X1 port map( D => reg_out_45_port, CLK => clk, 
                           RN => n669, Q => Ciphertext(45));
   Ciphertext_regx139x : DFFRNQ_X1 port map( D => reg_out_139_port, CLK => clk,
                           RN => n668, Q => Ciphertext(139));
   Ciphertext_regx188x : DFFRNQ_X1 port map( D => reg_out_188_port, CLK => clk,
                           RN => n667, Q => Ciphertext(188));
   Ciphertext_regx41x : DFFRNQ_X1 port map( D => reg_out_41_port, CLK => clk, 
                           RN => n666, Q => Ciphertext(41));
   Ciphertext_regx189x : DFFRNQ_X1 port map( D => reg_out_189_port, CLK => clk,
                           RN => n665, Q => Ciphertext(189));
   Ciphertext_regx151x : DFFRNQ_X1 port map( D => reg_out_151_port, CLK => clk,
                           RN => n664, Q => Ciphertext(151));
   Ciphertext_regx28x : DFFRNQ_X1 port map( D => reg_out_28_port, CLK => clk, 
                           RN => n663, Q => Ciphertext(28));
   Ciphertext_regx100x : DFFRNQ_X1 port map( D => reg_out_100_port, CLK => clk,
                           RN => n662, Q => Ciphertext(100));
   Ciphertext_regx64x : DFFRNQ_X1 port map( D => reg_out_64_port, CLK => clk, 
                           RN => n661, Q => Ciphertext(64));
   reg_in_regx51x : DFFRNQ_X1 port map( D => Plaintext(51), CLK => clk, RN => 
                           n659, Q => reg_in_51_port);
   Ciphertext_regx112x : DFFRNQ_X1 port map( D => reg_out_112_port, CLK => clk,
                           RN => n657, Q => Ciphertext(112));
   reg_in_regx29x : DFFRNQ_X1 port map( D => Plaintext(29), CLK => clk, RN => 
                           n656, Q => reg_in_29_port);
   Ciphertext_regx128x : DFFRNQ_X1 port map( D => reg_out_128_port, CLK => clk,
                           RN => n655, Q => Ciphertext(128));
   Ciphertext_regx89x : DFFRNQ_X1 port map( D => reg_out_89_port, CLK => clk, 
                           RN => n654, Q => Ciphertext(89));
   n654 <= '1';
   n655 <= '1';
   n656 <= '1';
   n657 <= '1';
   n659 <= '1';
   n661 <= '1';
   n662 <= '1';
   n663 <= '1';
   n664 <= '1';
   n665 <= '1';
   n666 <= '1';
   n667 <= '1';
   n668 <= '1';
   n669 <= '1';
   n670 <= '1';
   n671 <= '1';
   Ciphertext_regx12x : DFFRNQ_X1 port map( D => reg_out_12_port, CLK => clk, 
                           RN => n682, Q => Ciphertext(12));
   reg_in_regx71x : DFFRNQ_X1 port map( D => Plaintext(71), CLK => clk, RN => 
                           n681, Q => reg_in_71_port);
   reg_in_regx131x : DFFRNQ_X1 port map( D => Plaintext(131), CLK => clk, RN =>
                           n680, Q => reg_in_131_port);
   Ciphertext_regx124x : DFFRNQ_X1 port map( D => reg_out_124_port, CLK => clk,
                           RN => n679, Q => Ciphertext(124));
   Ciphertext_regx114x : DFFRNQ_X1 port map( D => reg_out_114_port, CLK => clk,
                           RN => n678, Q => Ciphertext(114));
   Ciphertext_regx120x : DFFRNQ_X1 port map( D => reg_out_120_port, CLK => clk,
                           RN => n677, Q => Ciphertext(120));
   reg_key_regx11x : DFFRNQ_X1 port map( D => Key(11), CLK => clk, RN => n676, 
                           Q => reg_key_11_port);
   Ciphertext_regx155x : DFFRNQ_X1 port map( D => reg_out_155_port, CLK => clk,
                           RN => n675, Q => Ciphertext(155));
   Ciphertext_regx17x : DFFRNQ_X1 port map( D => reg_out_17_port, CLK => clk, 
                           RN => n674, Q => Ciphertext(17));
   Ciphertext_regx99x : DFFRNQ_X1 port map( D => reg_out_99_port, CLK => clk, 
                           RN => n673, Q => Ciphertext(99));
   Ciphertext_regx56x : DFFSNQ_X1 port map( D => reg_out_56_port, CLK => clk, 
                           SN => n672, Q => Ciphertext(56));
   n672 <= '1';
   n673 <= '1';
   n674 <= '1';
   n675 <= '1';
   n676 <= '1';
   n677 <= '1';
   n678 <= '1';
   n679 <= '1';
   n680 <= '1';
   n681 <= '1';
   n682 <= '1';
   SPEEDY_instance : SPEEDY_Rounds5_0 port map( Plaintext(191) => 
                           reg_in_191_port, Plaintext(190) => reg_in_190_port, 
                           Plaintext(189) => reg_in_189_port, Plaintext(188) =>
                           reg_in_188_port, Plaintext(187) => reg_in_187_port, 
                           Plaintext(186) => reg_in_186_port, Plaintext(185) =>
                           reg_in_185_port, Plaintext(184) => reg_in_184_port, 
                           Plaintext(183) => reg_in_183_port, Plaintext(182) =>
                           reg_in_182_port, Plaintext(181) => reg_in_181_port, 
                           Plaintext(180) => reg_in_180_port, Plaintext(179) =>
                           reg_in_179_port, Plaintext(178) => reg_in_178_port, 
                           Plaintext(177) => reg_in_177_port, Plaintext(176) =>
                           reg_in_176_port, Plaintext(175) => reg_in_175_port, 
                           Plaintext(174) => reg_in_174_port, Plaintext(173) =>
                           reg_in_173_port, Plaintext(172) => reg_in_172_port, 
                           Plaintext(171) => reg_in_171_port, Plaintext(170) =>
                           reg_in_170_port, Plaintext(169) => reg_in_169_port, 
                           Plaintext(168) => reg_in_168_port, Plaintext(167) =>
                           reg_in_167_port, Plaintext(166) => reg_in_166_port, 
                           Plaintext(165) => reg_in_165_port, Plaintext(164) =>
                           reg_in_164_port, Plaintext(163) => reg_in_163_port, 
                           Plaintext(162) => reg_in_162_port, Plaintext(161) =>
                           reg_in_161_port, Plaintext(160) => reg_in_160_port, 
                           Plaintext(159) => reg_in_159_port, Plaintext(158) =>
                           reg_in_158_port, Plaintext(157) => reg_in_157_port, 
                           Plaintext(156) => reg_in_156_port, Plaintext(155) =>
                           reg_in_155_port, Plaintext(154) => reg_in_154_port, 
                           Plaintext(153) => reg_in_153_port, Plaintext(152) =>
                           reg_in_152_port, Plaintext(151) => reg_in_151_port, 
                           Plaintext(150) => reg_in_150_port, Plaintext(149) =>
                           reg_in_149_port, Plaintext(148) => reg_in_148_port, 
                           Plaintext(147) => reg_in_147_port, Plaintext(146) =>
                           reg_in_146_port, Plaintext(145) => reg_in_145_port, 
                           Plaintext(144) => reg_in_144_port, Plaintext(143) =>
                           reg_in_143_port, Plaintext(142) => reg_in_142_port, 
                           Plaintext(141) => reg_in_141_port, Plaintext(140) =>
                           reg_in_140_port, Plaintext(139) => reg_in_139_port, 
                           Plaintext(138) => reg_in_138_port, Plaintext(137) =>
                           reg_in_137_port, Plaintext(136) => reg_in_136_port, 
                           Plaintext(135) => reg_in_135_port, Plaintext(134) =>
                           reg_in_134_port, Plaintext(133) => reg_in_133_port, 
                           Plaintext(132) => reg_in_132_port, Plaintext(131) =>
                           reg_in_131_port, Plaintext(130) => reg_in_130_port, 
                           Plaintext(129) => reg_in_129_port, Plaintext(128) =>
                           reg_in_128_port, Plaintext(127) => reg_in_127_port, 
                           Plaintext(126) => reg_in_126_port, Plaintext(125) =>
                           reg_in_125_port, Plaintext(124) => reg_in_124_port, 
                           Plaintext(123) => reg_in_123_port, Plaintext(122) =>
                           reg_in_122_port, Plaintext(121) => reg_in_121_port, 
                           Plaintext(120) => reg_in_120_port, Plaintext(119) =>
                           reg_in_119_port, Plaintext(118) => reg_in_118_port, 
                           Plaintext(117) => reg_in_117_port, Plaintext(116) =>
                           reg_in_116_port, Plaintext(115) => reg_in_115_port, 
                           Plaintext(114) => reg_in_114_port, Plaintext(113) =>
                           reg_in_113_port, Plaintext(112) => reg_in_112_port, 
                           Plaintext(111) => reg_in_111_port, Plaintext(110) =>
                           reg_in_110_port, Plaintext(109) => reg_in_109_port, 
                           Plaintext(108) => reg_in_108_port, Plaintext(107) =>
                           reg_in_107_port, Plaintext(106) => reg_in_106_port, 
                           Plaintext(105) => reg_in_105_port, Plaintext(104) =>
                           reg_in_104_port, Plaintext(103) => reg_in_103_port, 
                           Plaintext(102) => reg_in_102_port, Plaintext(101) =>
                           reg_in_101_port, Plaintext(100) => reg_in_100_port, 
                           Plaintext(99) => reg_in_99_port, Plaintext(98) => 
                           reg_in_98_port, Plaintext(97) => reg_in_97_port, 
                           Plaintext(96) => reg_in_96_port, Plaintext(95) => 
                           reg_in_95_port, Plaintext(94) => reg_in_94_port, 
                           Plaintext(93) => reg_in_93_port, Plaintext(92) => 
                           reg_in_92_port, Plaintext(91) => reg_in_91_port, 
                           Plaintext(90) => reg_in_90_port, Plaintext(89) => 
                           reg_in_89_port, Plaintext(88) => reg_in_88_port, 
                           Plaintext(87) => reg_in_87_port, Plaintext(86) => 
                           reg_in_86_port, Plaintext(85) => reg_in_85_port, 
                           Plaintext(84) => reg_in_84_port, Plaintext(83) => 
                           reg_in_83_port, Plaintext(82) => reg_in_82_port, 
                           Plaintext(81) => reg_in_81_port, Plaintext(80) => 
                           reg_in_80_port, Plaintext(79) => reg_in_79_port, 
                           Plaintext(78) => reg_in_78_port, Plaintext(77) => 
                           reg_in_77_port, Plaintext(76) => reg_in_76_port, 
                           Plaintext(75) => reg_in_75_port, Plaintext(74) => 
                           reg_in_74_port, Plaintext(73) => reg_in_73_port, 
                           Plaintext(72) => reg_in_72_port, Plaintext(71) => 
                           reg_in_71_port, Plaintext(70) => reg_in_70_port, 
                           Plaintext(69) => reg_in_69_port, Plaintext(68) => 
                           reg_in_68_port, Plaintext(67) => reg_in_67_port, 
                           Plaintext(66) => reg_in_66_port, Plaintext(65) => 
                           reg_in_65_port, Plaintext(64) => reg_in_64_port, 
                           Plaintext(63) => reg_in_63_port, Plaintext(62) => 
                           reg_in_62_port, Plaintext(61) => reg_in_61_port, 
                           Plaintext(60) => reg_in_60_port, Plaintext(59) => 
                           reg_in_59_port, Plaintext(58) => reg_in_58_port, 
                           Plaintext(57) => reg_in_57_port, Plaintext(56) => 
                           reg_in_56_port, Plaintext(55) => reg_in_55_port, 
                           Plaintext(54) => reg_in_54_port, Plaintext(53) => 
                           reg_in_53_port, Plaintext(52) => reg_in_52_port, 
                           Plaintext(51) => reg_in_51_port, Plaintext(50) => 
                           reg_in_50_port, Plaintext(49) => reg_in_49_port, 
                           Plaintext(48) => reg_in_48_port, Plaintext(47) => 
                           reg_in_47_port, Plaintext(46) => reg_in_46_port, 
                           Plaintext(45) => reg_in_45_port, Plaintext(44) => 
                           reg_in_44_port, Plaintext(43) => reg_in_43_port, 
                           Plaintext(42) => reg_in_42_port, Plaintext(41) => 
                           reg_in_41_port, Plaintext(40) => reg_in_40_port, 
                           Plaintext(39) => reg_in_39_port, Plaintext(38) => 
                           reg_in_38_port, Plaintext(37) => reg_in_37_port, 
                           Plaintext(36) => reg_in_36_port, Plaintext(35) => 
                           reg_in_35_port, Plaintext(34) => reg_in_34_port, 
                           Plaintext(33) => reg_in_33_port, Plaintext(32) => 
                           reg_in_32_port, Plaintext(31) => reg_in_31_port, 
                           Plaintext(30) => reg_in_30_port, Plaintext(29) => 
                           reg_in_29_port, Plaintext(28) => reg_in_28_port, 
                           Plaintext(27) => reg_in_27_port, Plaintext(26) => 
                           reg_in_26_port, Plaintext(25) => reg_in_25_port, 
                           Plaintext(24) => reg_in_24_port, Plaintext(23) => 
                           reg_in_23_port, Plaintext(22) => reg_in_22_port, 
                           Plaintext(21) => reg_in_21_port, Plaintext(20) => 
                           reg_in_20_port, Plaintext(19) => reg_in_19_port, 
                           Plaintext(18) => reg_in_18_port, Plaintext(17) => 
                           reg_in_17_port, Plaintext(16) => reg_in_16_port, 
                           Plaintext(15) => reg_in_15_port, Plaintext(14) => 
                           reg_in_14_port, Plaintext(13) => reg_in_13_port, 
                           Plaintext(12) => reg_in_12_port, Plaintext(11) => 
                           reg_in_11_port, Plaintext(10) => reg_in_10_port, 
                           Plaintext(9) => reg_in_9_port, Plaintext(8) => 
                           reg_in_8_port, Plaintext(7) => reg_in_7_port, 
                           Plaintext(6) => reg_in_6_port, Plaintext(5) => 
                           reg_in_5_port, Plaintext(4) => reg_in_4_port, 
                           Plaintext(3) => reg_in_3_port, Plaintext(2) => 
                           reg_in_2_port, Plaintext(1) => reg_in_1_port, 
                           Plaintext(0) => reg_in_0_port, Key(191) => 
                           reg_key_191_port, Key(190) => reg_key_190_port, 
                           Key(189) => reg_key_189_port, Key(188) => 
                           reg_key_188_port, Key(187) => reg_key_187_port, 
                           Key(186) => reg_key_186_port, Key(185) => 
                           reg_key_185_port, Key(184) => reg_key_184_port, 
                           Key(183) => reg_key_183_port, Key(182) => 
                           reg_key_182_port, Key(181) => reg_key_181_port, 
                           Key(180) => reg_key_180_port, Key(179) => 
                           reg_key_179_port, Key(178) => reg_key_178_port, 
                           Key(177) => reg_key_177_port, Key(176) => 
                           reg_key_176_port, Key(175) => reg_key_175_port, 
                           Key(174) => reg_key_174_port, Key(173) => 
                           reg_key_173_port, Key(172) => reg_key_172_port, 
                           Key(171) => reg_key_171_port, Key(170) => 
                           reg_key_170_port, Key(169) => reg_key_169_port, 
                           Key(168) => reg_key_168_port, Key(167) => 
                           reg_key_167_port, Key(166) => reg_key_166_port, 
                           Key(165) => reg_key_165_port, Key(164) => 
                           reg_key_164_port, Key(163) => reg_key_163_port, 
                           Key(162) => reg_key_162_port, Key(161) => 
                           reg_key_161_port, Key(160) => reg_key_160_port, 
                           Key(159) => reg_key_159_port, Key(158) => 
                           reg_key_158_port, Key(157) => reg_key_157_port, 
                           Key(156) => reg_key_156_port, Key(155) => 
                           reg_key_155_port, Key(154) => reg_key_154_port, 
                           Key(153) => reg_key_153_port, Key(152) => 
                           reg_key_152_port, Key(151) => reg_key_151_port, 
                           Key(150) => reg_key_150_port, Key(149) => 
                           reg_key_149_port, Key(148) => reg_key_148_port, 
                           Key(147) => reg_key_147_port, Key(146) => 
                           reg_key_146_port, Key(145) => reg_key_145_port, 
                           Key(144) => reg_key_144_port, Key(143) => 
                           reg_key_143_port, Key(142) => reg_key_142_port, 
                           Key(141) => reg_key_141_port, Key(140) => 
                           reg_key_140_port, Key(139) => reg_key_139_port, 
                           Key(138) => reg_key_138_port, Key(137) => 
                           reg_key_137_port, Key(136) => reg_key_136_port, 
                           Key(135) => reg_key_135_port, Key(134) => 
                           reg_key_134_port, Key(133) => reg_key_133_port, 
                           Key(132) => reg_key_132_port, Key(131) => 
                           reg_key_131_port, Key(130) => reg_key_130_port, 
                           Key(129) => reg_key_129_port, Key(128) => 
                           reg_key_128_port, Key(127) => reg_key_127_port, 
                           Key(126) => reg_key_126_port, Key(125) => 
                           reg_key_125_port, Key(124) => reg_key_124_port, 
                           Key(123) => reg_key_123_port, Key(122) => 
                           reg_key_122_port, Key(121) => reg_key_121_port, 
                           Key(120) => reg_key_120_port, Key(119) => 
                           reg_key_119_port, Key(118) => reg_key_118_port, 
                           Key(117) => reg_key_117_port, Key(116) => 
                           reg_key_116_port, Key(115) => reg_key_115_port, 
                           Key(114) => reg_key_114_port, Key(113) => 
                           reg_key_113_port, Key(112) => reg_key_112_port, 
                           Key(111) => reg_key_111_port, Key(110) => 
                           reg_key_110_port, Key(109) => reg_key_109_port, 
                           Key(108) => reg_key_108_port, Key(107) => 
                           reg_key_107_port, Key(106) => reg_key_106_port, 
                           Key(105) => reg_key_105_port, Key(104) => 
                           reg_key_104_port, Key(103) => reg_key_103_port, 
                           Key(102) => reg_key_102_port, Key(101) => 
                           reg_key_101_port, Key(100) => reg_key_100_port, 
                           Key(99) => reg_key_99_port, Key(98) => 
                           reg_key_98_port, Key(97) => reg_key_97_port, Key(96)
                           => reg_key_96_port, Key(95) => reg_key_95_port, 
                           Key(94) => reg_key_94_port, Key(93) => 
                           reg_key_93_port, Key(92) => reg_key_92_port, Key(91)
                           => reg_key_91_port, Key(90) => reg_key_90_port, 
                           Key(89) => reg_key_89_port, Key(88) => 
                           reg_key_88_port, Key(87) => reg_key_87_port, Key(86)
                           => reg_key_86_port, Key(85) => reg_key_85_port, 
                           Key(84) => reg_key_84_port, Key(83) => 
                           reg_key_83_port, Key(82) => reg_key_82_port, Key(81)
                           => reg_key_81_port, Key(80) => reg_key_80_port, 
                           Key(79) => reg_key_79_port, Key(78) => 
                           reg_key_78_port, Key(77) => reg_key_77_port, Key(76)
                           => reg_key_76_port, Key(75) => reg_key_75_port, 
                           Key(74) => reg_key_74_port, Key(73) => 
                           reg_key_73_port, Key(72) => reg_key_72_port, Key(71)
                           => reg_key_71_port, Key(70) => reg_key_70_port, 
                           Key(69) => reg_key_69_port, Key(68) => 
                           reg_key_68_port, Key(67) => reg_key_67_port, Key(66)
                           => reg_key_66_port, Key(65) => reg_key_65_port, 
                           Key(64) => reg_key_64_port, Key(63) => 
                           reg_key_63_port, Key(62) => reg_key_62_port, Key(61)
                           => reg_key_61_port, Key(60) => reg_key_60_port, 
                           Key(59) => reg_key_59_port, Key(58) => 
                           reg_key_58_port, Key(57) => reg_key_57_port, Key(56)
                           => reg_key_56_port, Key(55) => reg_key_55_port, 
                           Key(54) => reg_key_54_port, Key(53) => 
                           reg_key_53_port, Key(52) => reg_key_52_port, Key(51)
                           => reg_key_51_port, Key(50) => reg_key_50_port, 
                           Key(49) => reg_key_49_port, Key(48) => 
                           reg_key_48_port, Key(47) => reg_key_47_port, Key(46)
                           => reg_key_46_port, Key(45) => reg_key_45_port, 
                           Key(44) => reg_key_44_port, Key(43) => 
                           reg_key_43_port, Key(42) => reg_key_42_port, Key(41)
                           => reg_key_41_port, Key(40) => reg_key_40_port, 
                           Key(39) => reg_key_39_port, Key(38) => 
                           reg_key_38_port, Key(37) => reg_key_37_port, Key(36)
                           => reg_key_36_port, Key(35) => reg_key_35_port, 
                           Key(34) => reg_key_34_port, Key(33) => 
                           reg_key_33_port, Key(32) => reg_key_32_port, Key(31)
                           => reg_key_31_port, Key(30) => reg_key_30_port, 
                           Key(29) => reg_key_29_port, Key(28) => 
                           reg_key_28_port, Key(27) => reg_key_27_port, Key(26)
                           => reg_key_26_port, Key(25) => reg_key_25_port, 
                           Key(24) => reg_key_24_port, Key(23) => 
                           reg_key_23_port, Key(22) => reg_key_22_port, Key(21)
                           => reg_key_21_port, Key(20) => reg_key_20_port, 
                           Key(19) => reg_key_19_port, Key(18) => 
                           reg_key_18_port, Key(17) => reg_key_17_port, Key(16)
                           => reg_key_16_port, Key(15) => reg_key_15_port, 
                           Key(14) => reg_key_14_port, Key(13) => 
                           reg_key_13_port, Key(12) => reg_key_12_port, Key(11)
                           => reg_key_11_port, Key(10) => reg_key_10_port, 
                           Key(9) => reg_key_9_port, Key(8) => reg_key_8_port, 
                           Key(7) => reg_key_7_port, Key(6) => reg_key_6_port, 
                           Key(5) => reg_key_5_port, Key(4) => reg_key_4_port, 
                           Key(3) => reg_key_3_port, Key(2) => reg_key_2_port, 
                           Key(1) => reg_key_1_port, Key(0) => reg_key_0_port, 
                           Ciphertext(191) => reg_out_191_port, Ciphertext(190)
                           => reg_out_190_port, Ciphertext(189) => 
                           reg_out_189_port, Ciphertext(188) => 
                           reg_out_188_port, Ciphertext(187) => 
                           reg_out_187_port, Ciphertext(186) => 
                           reg_out_186_port, Ciphertext(185) => 
                           reg_out_185_port, Ciphertext(184) => 
                           reg_out_184_port, Ciphertext(183) => 
                           reg_out_183_port, Ciphertext(182) => 
                           reg_out_182_port, Ciphertext(181) => 
                           reg_out_181_port, Ciphertext(180) => 
                           reg_out_180_port, Ciphertext(179) => 
                           reg_out_179_port, Ciphertext(178) => 
                           reg_out_178_port, Ciphertext(177) => 
                           reg_out_177_port, Ciphertext(176) => 
                           reg_out_176_port, Ciphertext(175) => 
                           reg_out_175_port, Ciphertext(174) => 
                           reg_out_174_port, Ciphertext(173) => 
                           reg_out_173_port, Ciphertext(172) => 
                           reg_out_172_port, Ciphertext(171) => 
                           reg_out_171_port, Ciphertext(170) => 
                           reg_out_170_port, Ciphertext(169) => 
                           reg_out_169_port, Ciphertext(168) => 
                           reg_out_168_port, Ciphertext(167) => 
                           reg_out_167_port, Ciphertext(166) => 
                           reg_out_166_port, Ciphertext(165) => 
                           reg_out_165_port, Ciphertext(164) => 
                           reg_out_164_port, Ciphertext(163) => 
                           reg_out_163_port, Ciphertext(162) => 
                           reg_out_162_port, Ciphertext(161) => 
                           reg_out_161_port, Ciphertext(160) => 
                           reg_out_160_port, Ciphertext(159) => 
                           reg_out_159_port, Ciphertext(158) => 
                           reg_out_158_port, Ciphertext(157) => 
                           reg_out_157_port, Ciphertext(156) => 
                           reg_out_156_port, Ciphertext(155) => 
                           reg_out_155_port, Ciphertext(154) => 
                           reg_out_154_port, Ciphertext(153) => 
                           reg_out_153_port, Ciphertext(152) => 
                           reg_out_152_port, Ciphertext(151) => 
                           reg_out_151_port, Ciphertext(150) => 
                           reg_out_150_port, Ciphertext(149) => 
                           reg_out_149_port, Ciphertext(148) => 
                           reg_out_148_port, Ciphertext(147) => 
                           reg_out_147_port, Ciphertext(146) => 
                           reg_out_146_port, Ciphertext(145) => 
                           reg_out_145_port, Ciphertext(144) => 
                           reg_out_144_port, Ciphertext(143) => 
                           reg_out_143_port, Ciphertext(142) => 
                           reg_out_142_port, Ciphertext(141) => 
                           reg_out_141_port, Ciphertext(140) => 
                           reg_out_140_port, Ciphertext(139) => 
                           reg_out_139_port, Ciphertext(138) => 
                           reg_out_138_port, Ciphertext(137) => 
                           reg_out_137_port, Ciphertext(136) => 
                           reg_out_136_port, Ciphertext(135) => 
                           reg_out_135_port, Ciphertext(134) => 
                           reg_out_134_port, Ciphertext(133) => 
                           reg_out_133_port, Ciphertext(132) => 
                           reg_out_132_port, Ciphertext(131) => 
                           reg_out_131_port, Ciphertext(130) => 
                           reg_out_130_port, Ciphertext(129) => 
                           reg_out_129_port, Ciphertext(128) => 
                           reg_out_128_port, Ciphertext(127) => 
                           reg_out_127_port, Ciphertext(126) => 
                           reg_out_126_port, Ciphertext(125) => 
                           reg_out_125_port, Ciphertext(124) => 
                           reg_out_124_port, Ciphertext(123) => 
                           reg_out_123_port, Ciphertext(122) => 
                           reg_out_122_port, Ciphertext(121) => 
                           reg_out_121_port, Ciphertext(120) => 
                           reg_out_120_port, Ciphertext(119) => 
                           reg_out_119_port, Ciphertext(118) => 
                           reg_out_118_port, Ciphertext(117) => 
                           reg_out_117_port, Ciphertext(116) => 
                           reg_out_116_port, Ciphertext(115) => 
                           reg_out_115_port, Ciphertext(114) => 
                           reg_out_114_port, Ciphertext(113) => 
                           reg_out_113_port, Ciphertext(112) => 
                           reg_out_112_port, Ciphertext(111) => 
                           reg_out_111_port, Ciphertext(110) => 
                           reg_out_110_port, Ciphertext(109) => 
                           reg_out_109_port, Ciphertext(108) => 
                           reg_out_108_port, Ciphertext(107) => 
                           reg_out_107_port, Ciphertext(106) => 
                           reg_out_106_port, Ciphertext(105) => 
                           reg_out_105_port, Ciphertext(104) => 
                           reg_out_104_port, Ciphertext(103) => 
                           reg_out_103_port, Ciphertext(102) => 
                           reg_out_102_port, Ciphertext(101) => 
                           reg_out_101_port, Ciphertext(100) => 
                           reg_out_100_port, Ciphertext(99) => reg_out_99_port,
                           Ciphertext(98) => reg_out_98_port, Ciphertext(97) =>
                           reg_out_97_port, Ciphertext(96) => reg_out_96_port, 
                           Ciphertext(95) => reg_out_95_port, Ciphertext(94) =>
                           reg_out_94_port, Ciphertext(93) => reg_out_93_port, 
                           Ciphertext(92) => reg_out_92_port, Ciphertext(91) =>
                           reg_out_91_port, Ciphertext(90) => reg_out_90_port, 
                           Ciphertext(89) => reg_out_89_port, Ciphertext(88) =>
                           reg_out_88_port, Ciphertext(87) => reg_out_87_port, 
                           Ciphertext(86) => reg_out_86_port, Ciphertext(85) =>
                           reg_out_85_port, Ciphertext(84) => reg_out_84_port, 
                           Ciphertext(83) => reg_out_83_port, Ciphertext(82) =>
                           reg_out_82_port, Ciphertext(81) => reg_out_81_port, 
                           Ciphertext(80) => reg_out_80_port, Ciphertext(79) =>
                           reg_out_79_port, Ciphertext(78) => reg_out_78_port, 
                           Ciphertext(77) => reg_out_77_port, Ciphertext(76) =>
                           reg_out_76_port, Ciphertext(75) => reg_out_75_port, 
                           Ciphertext(74) => reg_out_74_port, Ciphertext(73) =>
                           reg_out_73_port, Ciphertext(72) => reg_out_72_port, 
                           Ciphertext(71) => reg_out_71_port, Ciphertext(70) =>
                           reg_out_70_port, Ciphertext(69) => reg_out_69_port, 
                           Ciphertext(68) => reg_out_68_port, Ciphertext(67) =>
                           reg_out_67_port, Ciphertext(66) => reg_out_66_port, 
                           Ciphertext(65) => reg_out_65_port, Ciphertext(64) =>
                           reg_out_64_port, Ciphertext(63) => reg_out_63_port, 
                           Ciphertext(62) => reg_out_62_port, Ciphertext(61) =>
                           reg_out_61_port, Ciphertext(60) => reg_out_60_port, 
                           Ciphertext(59) => reg_out_59_port, Ciphertext(58) =>
                           reg_out_58_port, Ciphertext(57) => reg_out_57_port, 
                           Ciphertext(56) => reg_out_56_port, Ciphertext(55) =>
                           reg_out_55_port, Ciphertext(54) => reg_out_54_port, 
                           Ciphertext(53) => reg_out_53_port, Ciphertext(52) =>
                           reg_out_52_port, Ciphertext(51) => reg_out_51_port, 
                           Ciphertext(50) => reg_out_50_port, Ciphertext(49) =>
                           reg_out_49_port, Ciphertext(48) => reg_out_48_port, 
                           Ciphertext(47) => reg_out_47_port, Ciphertext(46) =>
                           reg_out_46_port, Ciphertext(45) => reg_out_45_port, 
                           Ciphertext(44) => reg_out_44_port, Ciphertext(43) =>
                           reg_out_43_port, Ciphertext(42) => reg_out_42_port, 
                           Ciphertext(41) => reg_out_41_port, Ciphertext(40) =>
                           reg_out_40_port, Ciphertext(39) => reg_out_39_port, 
                           Ciphertext(38) => reg_out_38_port, Ciphertext(37) =>
                           reg_out_37_port, Ciphertext(36) => reg_out_36_port, 
                           Ciphertext(35) => reg_out_35_port, Ciphertext(34) =>
                           reg_out_34_port, Ciphertext(33) => reg_out_33_port, 
                           Ciphertext(32) => reg_out_32_port, Ciphertext(31) =>
                           reg_out_31_port, Ciphertext(30) => reg_out_30_port, 
                           Ciphertext(29) => reg_out_29_port, Ciphertext(28) =>
                           reg_out_28_port, Ciphertext(27) => reg_out_27_port, 
                           Ciphertext(26) => reg_out_26_port, Ciphertext(25) =>
                           reg_out_25_port, Ciphertext(24) => reg_out_24_port, 
                           Ciphertext(23) => reg_out_23_port, Ciphertext(22) =>
                           reg_out_22_port, Ciphertext(21) => reg_out_21_port, 
                           Ciphertext(20) => reg_out_20_port, Ciphertext(19) =>
                           reg_out_19_port, Ciphertext(18) => reg_out_18_port, 
                           Ciphertext(17) => reg_out_17_port, Ciphertext(16) =>
                           reg_out_16_port, Ciphertext(15) => reg_out_15_port, 
                           Ciphertext(14) => reg_out_14_port, Ciphertext(13) =>
                           reg_out_13_port, Ciphertext(12) => reg_out_12_port, 
                           Ciphertext(11) => reg_out_11_port, Ciphertext(10) =>
                           reg_out_10_port, Ciphertext(9) => reg_out_9_port, 
                           Ciphertext(8) => reg_out_8_port, Ciphertext(7) => 
                           reg_out_7_port, Ciphertext(6) => reg_out_6_port, 
                           Ciphertext(5) => reg_out_5_port, Ciphertext(4) => 
                           reg_out_4_port, Ciphertext(3) => reg_out_3_port, 
                           Ciphertext(2) => reg_out_2_port, Ciphertext(1) => 
                           reg_out_1_port, Ciphertext(0) => reg_out_0_port);
   Ciphertext_regx187x : DFFRNQ_X1 port map( D => reg_out_187_port, CLK => clk,
                           RN => n692, Q => Ciphertext(187));
   Ciphertext_regx191x : DFFRNQ_X1 port map( D => reg_out_191_port, CLK => clk,
                           RN => n691, Q => Ciphertext(191));
   Ciphertext_regx76x : DFFRNQ_X1 port map( D => reg_out_76_port, CLK => clk, 
                           RN => n690, Q => Ciphertext(76));
   Ciphertext_regx53x : DFFRNQ_X1 port map( D => reg_out_53_port, CLK => clk, 
                           RN => n689, Q => Ciphertext(53));
   Ciphertext_regx134x : DFFRNQ_X1 port map( D => reg_out_134_port, CLK => clk,
                           RN => n688, Q => Ciphertext(134));
   reg_in_regx147x : DFFRNQ_X1 port map( D => Plaintext(147), CLK => clk, RN =>
                           n687, Q => reg_in_147_port);
   Ciphertext_regx168x : DFFRNQ_X1 port map( D => reg_out_168_port, CLK => clk,
                           RN => n686, Q => Ciphertext(168));
   Ciphertext_regx141x : DFFRNQ_X1 port map( D => reg_out_141_port, CLK => clk,
                           RN => n685, Q => Ciphertext(141));
   Ciphertext_regx67x : DFFRNQ_X1 port map( D => reg_out_67_port, CLK => clk, 
                           RN => n684, Q => Ciphertext(67));
   Ciphertext_regx148x : DFFRNQ_X1 port map( D => reg_out_148_port, CLK => clk,
                           RN => n683, Q => Ciphertext(148));
   n683 <= '1';
   n684 <= '1';
   n685 <= '1';
   n686 <= '1';
   n687 <= '1';
   n688 <= '1';
   n689 <= '1';
   n690 <= '1';
   n691 <= '1';
   n692 <= '1';

end SYN_Behavioral;
