
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_SPEEDY_Top is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_SPEEDY_Top;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Rounds6_0 is

   port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : out
         std_logic_vector (191 downto 0));

end SPEEDY_Rounds6_0;

architecture SYN_Behavioral of SPEEDY_Rounds6_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X4
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( I0, I1, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X12
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X4
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X8
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X8
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X8
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n21, n22, n24,
      n25, n27, n28, n29, n31, n32, n34, n36, n37, n38, n39, n42, n44, n46, n47
      , n50, n51, n52, n53, n54, n57, n60, n61, n62, n66, n67, n71, n72, n73, 
      n75, n78, n79, n81, n84, n85, n86, n87, n91, n92, n94, n97, n98, n100, 
      n101, n102, n107, n110, n111, n112, n115, n118, n119, n120, n123, n124, 
      n125, n128, n135, n136, n137, n138, n139, n144, n146, n149, n151, n152, 
      n153, n154, n155, n156, n161, n162, n164, n168, n169, n170, n171, n175, 
      n179, n180, n183, n184, n185, n187, n188, n193, n196, n204, n205, n206, 
      n207, n210, n214, n215, n219, n221, n224, n225, n227, n229, n230, n231, 
      n233, n236, n239, n242, n245, n250, n252, n253, n254, n258, n259, n261, 
      n262, n263, n265, n266, n268, n270, n273, n274, n275, n276, n277, n279, 
      n281, n283, n284, n285, n287, n292, n293, n294, n295, n297, n298, n299, 
      n300, n304, n305, n308, n313, n314, n315, n317, n319, n320, n321, n322, 
      n327, n328, n329, n330, n335, n337, n338, n339, n342, n343, n347, n348, 
      n349, n354, n355, n356, n358, n363, n365, n367, n371, n375, n376, n379, 
      n380, n384, n385, n386, n387, n388, n391, n392, n393, n396, n397, n398, 
      n400, n401, n402, n405, n406, n408, n410, n412, n413, n414, n415, n416, 
      n417, n419, n420, n421, n423, n424, n425, n431, n432, n433, n434, n436, 
      n437, n438, n439, n440, n442, n443, n444, n445, n446, n447, n448, n449, 
      n450, n452, n453, n454, n456, n457, n458, n460, n461, n462, n463, n465, 
      n467, n468, n469, n470, n471, n474, n475, n476, n477, n478, n479, n480, 
      n481, n485, n487, n488, n489, n490, n493, n494, n495, n496, n497, n498, 
      n499, n500, n502, n503, n505, n506, n507, n508, n509, n510, n511, n513, 
      n514, n515, n516, n517, n518, n519, n521, n522, n524, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n553, n554, 
      n556, n560, n561, n562, n563, n564, n565, n567, n568, n570, n571, n572, 
      n575, n576, n577, n578, n579, n580, n582, n583, n584, n586, n587, n589, 
      n590, n591, n595, n596, n598, n599, n600, n601, n602, n603, n606, n607, 
      n609, n610, n612, n613, n615, n616, n618, n620, n621, n622, n623, n624, 
      n625, n627, n628, n629, n630, n632, n634, n635, n636, n637, n639, n641, 
      n642, n643, n645, n646, n647, n651, n652, n654, n655, n657, n660, n661, 
      n662, n663, n664, n665, n666, n667, n668, n671, n673, n675, n676, n678, 
      n679, n680, n681, n686, n689, n690, n691, n692, n693, n694, n695, n696, 
      n698, n699, n700, n701, n702, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n721, n722, n723, n724, 
      n725, n727, n728, n729, n730, n732, n733, n734, n736, n737, n738, n739, 
      n741, n742, n743, n744, n745, n746, n747, n749, n750, n751, n752, n753, 
      n754, n755, n756, n757, n758, n760, n761, n763, n764, n765, n767, n769, 
      n770, n772, n773, n776, n777, n779, n780, n781, n782, n783, n784, n785, 
      n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, 
      n798, n801, n802, n803, n805, n806, n808, n809, n810, n812, n816, n817, 
      n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
      n830, n831, n832, n833, n834, n836, n837, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n855, n856, 
      n857, n858, n859, n861, n862, n864, n865, n867, n868, n870, n871, n873, 
      n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, 
      n887, n888, n889, n890, n891, n893, n895, n896, n897, n898, n899, n900, 
      n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, 
      n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n924, n925, 
      n926, n927, n929, n930, n931, n932, n933, n935, n936, n937, n938, n939, 
      n940, n941, n942, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n972, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n985, n986, n987, n989, n990, n992, n994, 
      n995, n996, n998, n1000, n1001, n1003, n1004, n1007, n1008, n1009, n1012,
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1022, n1023, 
      n1024, n1026, n1028, n1030, n1032, n1034, n1035, n1036, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1059, n1060, n1063, 
      n1064, n1065, n1067, n1069, n1070, n1071, n1074, n1075, n1076, n1077, 
      n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, 
      n1089, n1090, n1092, n1093, n1094, n1096, n1098, n1099, n1100, n1101, 
      n1102, n1104, n1106, n1107, n1108, n1109, n1112, n1113, n1116, n1117, 
      n1119, n1120, n1122, n1124, n1125, n1127, n1128, n1129, n1130, n1131, 
      n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, 
      n1142, n1143, n1145, n1146, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1163, n1164, 
      n1165, n1166, n1167, n1168, n1169, n1170, n1172, n1173, n1175, n1177, 
      n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1188, n1189, 
      n1190, n1191, n1192, n1193, n1194, n1196, n1197, n1198, n1200, n1201, 
      n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1218, n1219, n1221, n1223, n1224, n1225, 
      n1226, n1227, n1228, n1230, n1231, n1232, n1233, n1235, n1237, n1238, 
      n1239, n1240, n1241, n1243, n1244, n1245, n1246, n1247, n1249, n1250, 
      n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, 
      n1262, n1263, n1264, n1265, n1266, n1267, n1269, n1271, n1274, n1275, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1284, n1286, n1287, n1288, 
      n1289, n1290, n1291, n1292, n1294, n1296, n1297, n1298, n1299, n1300, 
      n1302, n1303, n1305, n1306, n1307, n1308, n1309, n1310, n1312, n1313, 
      n1315, n1316, n1317, n1318, n1319, n1321, n1322, n1323, n1325, n1326, 
      n1327, n1328, n1329, n1331, n1332, n1333, n1334, n1335, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1372, n1373, n1374, n1376, n1377, n1378, n1379, n1380, 
      n1382, n1384, n1385, n1386, n1387, n1389, n1390, n1391, n1392, n1393, 
      n1394, n1395, n1396, n1397, n1398, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1409, n1410, n1411, n1413, n1414, n1415, n1416, n1417, n1419, 
      n1420, n1421, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
      n1431, n1432, n1433, n1434, n1436, n1438, n1439, n1441, n1445, n1446, 
      n1449, n1450, n1451, n1452, n1453, n1454, n1456, n1457, n1458, n1462, 
      n1463, n1464, n1465, n1466, n1468, n1469, n1470, n1471, n1472, n1473, 
      n1474, n1475, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, 
      n1489, n1490, n1491, n1492, n1494, n1496, n1497, n1499, n1500, n1504, 
      n1506, n1507, n1508, n1511, n1513, n1516, n1519, n1521, n1522, n1523, 
      n1524, n1525, n1528, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
      n1538, n1540, n1541, n1543, n1544, n1545, n1546, n1547, n1549, n1550, 
      n1553, n1555, n1557, n1559, n1560, n1561, n1563, n1564, n1565, n1567, 
      n1571, n1572, n1573, n1577, n1579, n1580, n1581, n1587, n1588, n1589, 
      n1590, n1592, n1594, n1595, n1596, n1597, n1600, n1601, n1602, n1603, 
      n1604, n1607, n1609, n1610, n1612, n1613, n1615, n1616, n1617, n1619, 
      n1620, n1621, n1622, n1627, n1628, n1629, n1630, n1631, n1632, n1633, 
      n1634, n1635, n1636, n1640, n1641, n1642, n1644, n1645, n1646, n1647, 
      n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1658, n1659, 
      n1661, n1663, n1664, n1668, n1669, n1671, n1672, n1673, n1676, n1677, 
      n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, 
      n1688, n1690, n1694, n1695, n1696, n1698, n1699, n1700, n1702, n1703, 
      n1704, n1707, n1708, n1709, n1710, n1712, n1713, n1714, n1716, n1718, 
      n1719, n1720, n1726, n1727, n1728, n1730, n1731, n1732, n1733, n1734, 
      n1736, n1741, n1742, n1745, n1746, n1749, n1751, n1756, n1757, n1758, 
      n1760, n1761, n1762, n1763, n1764, n1766, n1767, n1768, n1769, n1770, 
      n1771, n1772, n1773, n1774, n1775, n1776, n1778, n1779, n1780, n1781, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1791, n1792, n1793, 
      n1794, n1795, n1796, n1799, n1800, n1801, n1803, n1805, n1807, n1808, 
      n1811, n1812, n1813, n1814, n1815, n1816, n1818, n1819, n1820, n1825, 
      n1826, n1828, n1830, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
      n1842, n1844, n1845, n1848, n1850, n1851, n1853, n1857, n1858, n1859, 
      n1861, n1862, n1863, n1864, n1865, n1867, n1868, n1869, n1870, n1871, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1881, n1882, n1883, n1884, 
      n1886, n1887, n1889, n1890, n1892, n1896, n1897, n1898, n1900, n1902, 
      n1903, n1905, n1908, n1909, n1910, n1911, n1913, n1914, n1915, n1916, 
      n1917, n1920, n1923, n1926, n1927, n1928, n1929, n1930, n1931, n1933, 
      n1934, n1935, n1936, n1937, n1938, n1940, n1941, n1942, n1944, n1945, 
      n1946, n1948, n1949, n1950, n1951, n1954, n1955, n1956, n1957, n1960, 
      n1961, n1962, n1963, n1964, n1965, n1967, n1968, n1970, n1971, n1973, 
      n1974, n1976, n1978, n1979, n1980, n1982, n1983, n1984, n1986, n1988, 
      n1990, n1991, n1992, n1993, n1994, n1995, n1997, n1998, n2000, n2001, 
      n2002, n2003, n2004, n2005, n2009, n2012, n2013, n2015, n2016, n2017, 
      n2018, n2019, n2021, n2022, n2023, n2024, n2028, n2029, n2031, n2032, 
      n2036, n2037, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2048, 
      n2049, n2052, n2053, n2054, n2055, n2060, n2061, n2064, n2066, n2069, 
      n2070, n2072, n2073, n2074, n2075, n2076, n2078, n2080, n2081, n2082, 
      n2084, n2085, n2086, n2088, n2089, n2092, n2095, n2097, n2098, n2099, 
      n2100, n2101, n2103, n2104, n2105, n2107, n2108, n2111, n2112, n2113, 
      n2114, n2117, n2118, n2122, n2123, n2124, n2125, n2126, n2128, n2129, 
      n2130, n2132, n2134, n2135, n2137, n2138, n2141, n2142, n2143, n2144, 
      n2145, n2146, n2147, n2148, n2149, n2150, n2152, n2153, n2154, n2155, 
      n2156, n2158, n2161, n2162, n2163, n2164, n2166, n2167, n2169, n2172, 
      n2173, n2174, n2176, n2177, n2178, n2180, n2182, n2186, n2190, n2191, 
      n2192, n2197, n2198, n2200, n2202, n2203, n2204, n2205, n2206, n2207, 
      n2208, n2209, n2210, n2211, n2212, n2214, n2215, n2217, n2219, n2221, 
      n2222, n2225, n2226, n2229, n2230, n2233, n2234, n2236, n2237, n2239, 
      n2241, n2242, n2245, n2247, n2250, n2251, n2252, n2253, n2256, n2257, 
      n2258, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2270, 
      n2271, n2272, n2275, n2277, n2278, n2279, n2280, n2281, n2282, n2283, 
      n2285, n2288, n2289, n2290, n2291, n2292, n2293, n2296, n2297, n2298, 
      n2299, n2300, n2301, n2302, n2304, n2305, n2306, n2308, n2309, n2311, 
      n2312, n2315, n2316, n2317, n2318, n2319, n2320, n2324, n2325, n2330, 
      n2331, n2333, n2334, n2335, n2337, n2338, n2339, n2342, n2345, n2347, 
      n2348, n2349, n2351, n2352, n2353, n2355, n2356, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2375, 
      n2378, n2380, n2381, n2383, n2384, n2386, n2387, n2388, n2389, n2390, 
      n2391, n2393, n2394, n2395, n2396, n2398, n2400, n2401, n2404, n2405, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2414, n2415, n2417, n2418, 
      n2420, n2421, n2423, n2424, n2427, n2430, n2432, n2435, n2436, n2440, 
      n2441, n2442, n2443, n2444, n2447, n2448, n2449, n2450, n2452, n2455, 
      n2456, n2458, n2460, n2463, n2464, n2466, n2468, n2469, n2470, n2471, 
      n2472, n2473, n2476, n2477, n2479, n2480, n2483, n2484, n2486, n2489, 
      n2490, n2491, n2492, n2495, n2497, n2498, n2499, n2500, n2501, n2502, 
      n2507, n2508, n2509, n2512, n2513, n2514, n2517, n2518, n2519, n2520, 
      n2522, n2523, n2524, n2525, n2526, n2529, n2534, n2535, n2536, n2537, 
      n2538, n2539, n2547, n2548, n2549, n2550, n2551, n2554, n2556, n2557, 
      n2558, n2560, n2561, n2563, n2564, n2565, n2566, n2568, n2569, n2570, 
      n2574, n2575, n2576, n2577, n2579, n2580, n2581, n2582, n2583, n2584, 
      n2585, n2587, n2589, n2590, n2591, n2592, n2593, n2595, n2596, n2598, 
      n2599, n2600, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, 
      n2610, n2611, n2612, n2613, n2614, n2616, n2618, n2619, n2620, n2621, 
      n2622, n2623, n2624, n2625, n2626, n2628, n2631, n2632, n2633, n2634, 
      n2635, n2636, n2637, n2638, n2639, n2640, n2642, n2643, n2646, n2647, 
      n2648, n2649, n2650, n2651, n2653, n2654, n2655, n2656, n2657, n2661, 
      n2664, n2665, n2666, n2667, n2668, n2671, n2672, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2682, n2683, n2684, n2686, n2687, n2689, 
      n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2703, 
      n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2712, n2713, n2715, 
      n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2731, n2732, n2733, n2734, n2738, n2739, n2741, 
      n2743, n2744, n2745, n2746, n2747, n2750, n2752, n2753, n2754, n2756, 
      n2757, n2758, n2759, n2761, n2763, n2764, n2766, n2767, n2770, n2771, 
      n2773, n2775, n2777, n2778, n2780, n2784, n2785, n2786, n2788, n2789, 
      n2790, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2801, n2802, 
      n2803, n2808, n2809, n2812, n2813, n2818, n2819, n2820, n2821, n2822, 
      n2824, n2825, n2826, n2831, n2833, n2834, n2838, n2839, n2840, n2841, 
      n2842, n2843, n2844, n2845, n2847, n2848, n2849, n2851, n2852, n2853, 
      n2854, n2855, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, 
      n2865, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2883, n2886, n2888, n2889, n2890, 
      n2891, n2894, n2896, n2898, n2899, n2900, n2901, n2902, n2903, n2904, 
      n2905, n2906, n2908, n2909, n2911, n2912, n2913, n2915, n2917, n2918, 
      n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
      n2930, n2933, n2934, n2935, n2936, n2937, n2939, n2940, n2941, n2943, 
      n2944, n2945, n2946, n2948, n2949, n2951, n2952, n2953, n2956, n2957, 
      n2958, n2959, n2960, n2961, n2962, n2964, n2965, n2967, n2968, n2969, 
      n2970, n2971, n2972, n2974, n2975, n2976, n2978, n2980, n2981, n2982, 
      n2983, n2986, n2987, n2989, n2990, n2992, n2993, n2996, n2997, n2998, 
      n2999, n3001, n3003, n3004, n3005, n3006, n3007, n3009, n3010, n3012, 
      n3013, n3014, n3016, n3018, n3019, n3021, n3022, n3023, n3024, n3026, 
      n3027, n3028, n3030, n3032, n3033, n3035, n3036, n3038, n3039, n3041, 
      n3042, n3043, n3045, n3047, n3048, n3049, n3050, n3051, n3052, n3055, 
      n3056, n3057, n3059, n3060, n3061, n3063, n3065, n3068, n3069, n3070, 
      n3071, n3072, n3073, n3074, n3076, n3077, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3090, n3091, n3092, n3093, n3094, 
      n3096, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3109, 
      n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, 
      n3122, n3123, n3124, n3126, n3128, n3131, n3132, n3133, n3134, n3135, 
      n3136, n3137, n3140, n3142, n3143, n3144, n3146, n3147, n3148, n3149, 
      n3152, n3155, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, 
      n3165, n3166, n3168, n3169, n3170, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3179, n3180, n3181, n3183, n3184, n3186, n3187, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3197, n3198, n3199, 
      n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
      n3211, n3212, n3213, n3214, n3216, n3217, n3218, n3219, n3220, n3221, 
      n3222, n3223, n3224, n3225, n3226, n3227, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3239, n3240, n3241, n3242, n3243, 
      n3244, n3245, n3247, n3248, n3250, n3251, n3253, n3255, n3256, n3257, 
      n3258, n3259, n3260, n3266, n3267, n3269, n3270, n3271, n3272, n3275, 
      n3280, n3281, n3282, n3283, n3285, n3286, n3288, n3289, n3292, n3293, 
      n3294, n3295, n3296, n3297, n3298, n3300, n3303, n3304, n3305, n3307, 
      n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, 
      n3318, n3319, n3322, n3324, n3325, n3327, n3328, n3329, n3332, n3334, 
      n3336, n3339, n3340, n3341, n3343, n3344, n3345, n3348, n3350, n3351, 
      n3352, n3353, n3354, n3355, n3357, n3358, n3360, n3361, n3364, n3365, 
      n3366, n3368, n3369, n3371, n3375, n3376, n3378, n3379, n3380, n3382, 
      n3384, n3385, n3388, n3389, n3390, n3391, n3392, n3393, n3395, n3396, 
      n3399, n3401, n3402, n3403, n3405, n3407, n3408, n3410, n3411, n3412, 
      n3415, n3416, n3417, n3418, n3420, n3421, n3424, n3425, n3428, n3429, 
      n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3439, n3440, 
      n3441, n3442, n3443, n3445, n3446, n3447, n3448, n3449, n3451, n3454, 
      n3455, n3461, n3462, n3463, n3465, n3467, n3468, n3469, n3472, n3475, 
      n3476, n3477, n3480, n3481, n3482, n3483, n3484, n3486, n3487, n3489, 
      n3491, n3493, n3494, n3495, n3497, n3499, n3501, n3502, n3503, n3504, 
      n3506, n3508, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3522, n3525, n3526, n3527, n3529, n3530, n3535, 
      n3536, n3539, n3540, n3541, n3544, n3545, n3546, n3547, n3548, n3549, 
      n3550, n3552, n3553, n3554, n3556, n3558, n3559, n3562, n3565, n3566, 
      n3567, n3568, n3569, n3570, n3571, n3574, n3575, n3576, n3578, n3579, 
      n3580, n3581, n3583, n3584, n3586, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3596, n3597, n3598, n3599, n3600, n3601, n3603, n3604, 
      n3605, n3606, n3614, n3617, n3618, n3619, n3620, n3621, n3622, n3624, 
      n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, 
      n3638, n3639, n3643, n3644, n3646, n3648, n3650, n3651, n3652, n3653, 
      n3654, n3656, n3657, n3658, n3659, n3663, n3665, n3667, n3668, n3669, 
      n3670, n3672, n3673, n3677, n3678, n3680, n3682, n3683, n3685, n3686, 
      n3687, n3689, n3692, n3694, n3695, n3696, n3698, n3702, n3703, n3704, 
      n3705, n3706, n3708, n3711, n3717, n3718, n3722, n3723, n3724, n3725, 
      n3727, n3728, n3729, n3730, n3731, n3732, n3735, n3736, n3737, n3739, 
      n3742, n3744, n3746, n3748, n3750, n3751, n3755, n3756, n3757, n3759, 
      n3760, n3767, n3769, n3770, n3771, n3772, n3773, n3774, n3777, n3778, 
      n3779, n3780, n3781, n3782, n3783, n3784, n3786, n3787, n3788, n3790, 
      n3791, n3792, n3793, n3794, n3796, n3797, n3798, n3799, n3800, n3801, 
      n3807, n3809, n3810, n3812, n3815, n3816, n3819, n3820, n3821, n3822, 
      n3824, n3825, n3826, n3827, n3828, n3830, n3835, n3836, n3840, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3851, n3852, n3854, n3856, n3860, 
      n3861, n3862, n3866, n3867, n3868, n3870, n3873, n3874, n3879, n3880, 
      n3883, n3884, n3885, n3888, n3889, n3891, n3893, n3894, n3896, n3898, 
      n3900, n3901, n3902, n3903, n3904, n3905, n3908, n3909, n3911, n3915, 
      n3916, n3918, n3919, n3920, n3922, n3923, n3924, n3925, n3926, n3927, 
      n3928, n3929, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, 
      n3940, n3941, n3944, n3945, n3946, n3947, n3950, n3951, n3954, n3955, 
      n3957, n3958, n3962, n3963, n3964, n3967, n3970, n3972, n3973, n3977, 
      n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, 
      n3989, n3990, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4003, 
      n4004, n4006, n4008, n4013, n4014, n4015, n4016, n4017, n4019, n4020, 
      n4021, n4024, n4025, n4026, n4028, n4029, n4034, n4035, n4036, n4040, 
      n4041, n4042, n4043, n4045, n4047, n4049, n4050, n4051, n4052, n4053, 
      n4054, n4055, n4056, n4057, n4059, n4060, n4061, n4062, n4063, n4065, 
      n4066, n4067, n4069, n4070, n4071, n4075, n4076, n4077, n4079, n4082, 
      n4084, n4086, n4087, n4088, n4089, n4091, n4095, n4097, n4098, n4099, 
      n4100, n4101, n4102, n4106, n4107, n4110, n4111, n4112, n4113, n4114, 
      n4117, n4118, n4119, n4123, n4124, n4130, n4131, n4133, n4134, n4135, 
      n4136, n4140, n4142, n4143, n4145, n4146, n4150, n4151, n4154, n4155, 
      n4156, n4157, n4158, n4161, n4162, n4163, n4164, n4167, n4168, n4169, 
      n4173, n4174, n4176, n4177, n4178, n4179, n4180, n4182, n4183, n4184, 
      n4186, n4187, n4188, n4191, n4192, n4193, n4194, n4196, n4197, n4200, 
      n4201, n4202, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, 
      n4212, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4224, 
      n4225, n4226, n4228, n4230, n4231, n4232, n4233, n4234, n4236, n4240, 
      n4241, n4243, n4244, n4245, n4246, n4248, n4251, n4253, n4254, n4255, 
      n4259, n4260, n4261, n4262, n4263, n4266, n4267, n4268, n4269, n4273, 
      n4274, n4279, n4280, n4281, n4283, n4284, n4285, n4286, n4287, n4289, 
      n4290, n4291, n4293, n4295, n4299, n4300, n4301, n4302, n4305, n4306, 
      n4308, n4310, n4311, n4312, n4314, n4315, n4318, n4319, n4321, n4324, 
      n4325, n4327, n4329, n4330, n4331, n4332, n4335, n4337, n4338, n4339, 
      n4340, n4341, n4342, n4349, n4350, n4352, n4353, n4354, n4355, n4356, 
      n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, 
      n4368, n4370, n4371, n4373, n4374, n4375, n4378, n4379, n4380, n4381, 
      n4382, n4384, n4385, n4386, n4387, n4390, n4391, n4392, n4393, n4395, 
      n4396, n4397, n4398, n4399, n4400, n4401, n4403, n4405, n4407, n4408, 
      n4409, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, 
      n4420, n4422, n4423, n4425, n4427, n4432, n4433, n4434, n4435, n4436, 
      n4437, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, 
      n4450, n4451, n4452, n4453, n4456, n4458, n4459, n4460, n4464, n4465, 
      n4466, n4467, n4468, n4469, n4471, n4472, n4474, n4476, n4477, n4481, 
      n4483, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4494, n4496, 
      n4497, n4498, n4500, n4502, n4503, n4504, n4505, n4506, n4507, n4508, 
      n4510, n4511, n4514, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
      n4524, n4525, n4529, n4530, n4531, n4533, n4534, n4535, n4536, n4538, 
      n4539, n4542, n4543, n4547, n4550, n4551, n4552, n4554, n4555, n4556, 
      n4557, n4559, n4560, n4562, n4563, n4564, n4565, n4566, n4567, n4568, 
      n4569, n4571, n4572, n4574, n4577, n4578, n4579, n4580, n4581, n4583, 
      n4585, n4586, n4587, n4589, n4590, n4591, n4592, n4594, n4595, n4596, 
      n4599, n4601, n4602, n4604, n4607, n4609, n4610, n4611, n4613, n4614, 
      n4616, n4617, n4618, n4619, n4622, n4624, n4626, n4627, n4628, n4629, 
      n4631, n4632, n4633, n4635, n4636, n4637, n4638, n4639, n4642, n4643, 
      n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4655, 
      n4656, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4668, 
      n4669, n4671, n4672, n4674, n4675, n4677, n4678, n4680, n4681, n4682, 
      n4683, n4685, n4686, n4687, n4688, n4689, n4693, n4699, n4700, n4701, 
      n4704, n4706, n4708, n4709, n4710, n4711, n4713, n4714, n4715, n4716, 
      n4717, n4718, n4719, n4720, n4723, n4724, n4725, n4726, n4727, n4728, 
      n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4739, n4740, n4741, 
      n4743, n4744, n4746, n4747, n4749, n4750, n4755, n4756, n4758, n4759, 
      n4760, n4761, n4762, n4763, n4765, n4767, n4768, n4769, n4770, n4771, 
      n4772, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4783, n4784, n4785, n4786, n4788, n4789, n4790, n4791, n4792, n4794, 
      n4797, n4798, n4800, n4801, n4803, n4804, n4805, n4806, n4807, n4808, 
      n4809, n4810, n4811, n4812, n4814, n4816, n4820, n4821, n4822, n4823, 
      n4824, n4831, n4833, n4834, n4835, n4840, n4841, n4842, n4843, n4845, 
      n4846, n4847, n4849, n4850, n4854, n4855, n4856, n4857, n4858, n4859, 
      n4861, n4862, n4863, n4865, n4867, n4868, n4869, n4871, n4872, n4873, 
      n4878, n4879, n4880, n4881, n4883, n4884, n4885, n4886, n4891, n4892, 
      n4893, n4894, n4895, n4897, n4898, n4899, n4900, n4903, n4906, n4908, 
      n4909, n4913, n4914, n4915, n4916, n4918, n4919, n4920, n4922, n4925, 
      n4926, n4927, n4928, n4930, n4931, n4932, n4935, n4936, n4937, n4938, 
      n4942, n4944, n4949, n4951, n4952, n4953, n4955, n4956, n4959, n4960, 
      n4961, n4964, n4965, n4967, n4968, n4971, n4972, n4975, n4976, n4980, 
      n4982, n4983, n4984, n4985, n4986, n4988, n4989, n4991, n4992, n4993, 
      n4994, n4996, n4997, n4999, n5000, n5002, n5003, n5004, n5009, n5011, 
      n5012, n5013, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5029, n5030, n5031, n5032, n5033, n5034, 
      n5035, n5038, n5039, n5040, n5041, n5043, n5045, n5047, n5048, n5049, 
      n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5058, n5059, n5061, 
      n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, 
      n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5086, n5089, n5090, 
      n5091, n5092, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5103, 
      n5104, n5105, n5106, n5107, n5109, n5111, n5112, n5113, n5115, n5116, 
      n5118, n5119, n5121, n5122, n5124, n5126, n5127, n5128, n5129, n5130, 
      n5132, n5133, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5145, 
      n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5154, n5155, n5157, 
      n5158, n5159, n5160, n5161, n5162, n5163, n5166, n5169, n5170, n5172, 
      n5173, n5174, n5177, n5178, n5182, n5184, n5185, n5186, n5187, n5188, 
      n5190, n5191, n5194, n5196, n5197, n5199, n5202, n5203, n5205, n5206, 
      n5207, n5209, n5210, n5211, n5212, n5215, n5216, n5217, n5218, n5219, 
      n5221, n5222, n5223, n5225, n5226, n5227, n5228, n5229, n5231, n5233, 
      n5236, n5237, n5238, n5239, n5240, n5241, n5243, n5244, n5248, n5250, 
      n5252, n5253, n5254, n5255, n5256, n5258, n5259, n5260, n5261, n5263, 
      n5264, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, 
      n5275, n5277, n5278, n5279, n5280, n5282, n5284, n5286, n5287, n5288, 
      n5289, n5292, n5296, n5297, n5300, n5301, n5303, n5304, n5305, n5306, 
      n5307, n5308, n5309, n5311, n5314, n5315, n5316, n5317, n5318, n5321, 
      n5322, n5324, n5327, n5328, n5329, n5332, n5333, n5335, n5336, n5337, 
      n5338, n5339, n5340, n5342, n5343, n5345, n5347, n5348, n5349, n5350, 
      n5351, n5352, n5353, n5356, n5357, n5358, n5361, n5366, n5367, n5371, 
      n5372, n5373, n5374, n5376, n5377, n5378, n5379, n5380, n5381, n5382, 
      n5383, n5384, n5385, n5387, n5389, n5392, n5394, n5395, n5396, n5399, 
      n5400, n5401, n5402, n5405, n5407, n5408, n5410, n5411, n5412, n5413, 
      n5414, n5415, n5416, n5417, n5418, n5421, n5422, n5424, n5425, n5428, 
      n5429, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5440, 
      n5441, n5445, n5448, n5449, n5451, n5452, n5453, n5454, n5455, n5456, 
      n5457, n5458, n5459, n5460, n5462, n5466, n5467, n5468, n5469, n5470, 
      n5471, n5472, n5473, n5474, n5476, n5477, n5478, n5480, n5481, n5482, 
      n5483, n5484, n5485, n5487, n5488, n5490, n5491, n5492, n5494, n5495, 
      n5496, n5497, n5498, n5500, n5501, n5503, n5504, n5505, n5508, n5509, 
      n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5520, n5522, 
      n5523, n5525, n5526, n5527, n5529, n5530, n5532, n5533, n5534, n5535, 
      n5539, n5543, n5544, n5545, n5546, n5548, n5549, n5550, n5553, n5555, 
      n5556, n5558, n5560, n5561, n5562, n5563, n5568, n5570, n5571, n5572, 
      n5573, n5575, n5577, n5578, n5581, n5582, n5583, n5586, n5587, n5588, 
      n5589, n5590, n5592, n5593, n5594, n5595, n5597, n5598, n5600, n5601, 
      n5602, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, 
      n5615, n5616, n5618, n5619, n5620, n5621, n5622, n5624, n5625, n5627, 
      n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, 
      n5638, n5640, n5641, n5642, n5644, n5645, n5646, n5647, n5648, n5653, 
      n5654, n5655, n5656, n5657, n5658, n5659, n5662, n5663, n5666, n5668, 
      n5669, n5670, n5671, n5672, n5673, n5675, n5676, n5677, n5678, n5679, 
      n5680, n5681, n5682, n5683, n5684, n5685, n5687, n5689, n5690, n5691, 
      n5692, n5693, n5694, n5696, n5697, n5698, n5699, n5700, n5702, n5703, 
      n5704, n5707, n5708, n5709, n5710, n5712, n5713, n5714, n5717, n5718, 
      n5722, n5724, n5725, n5726, n5730, n5732, n5733, n5734, n5735, n5736, 
      n5737, n5741, n5742, n5743, n5744, n5745, n5748, n5751, n5752, n5753, 
      n5754, n5755, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, 
      n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, 
      n5776, n5777, n5779, n5781, n5782, n5784, n5786, n5787, n5788, n5789, 
      n5790, n5791, n5792, n5793, n5795, n5796, n5801, n5804, n5805, n5810, 
      n5812, n5813, n5814, n5817, n5820, n5821, n5822, n5825, n5826, n5827, 
      n5828, n5830, n5832, n5834, n5835, n5836, n5837, n5838, n5839, n5842, 
      n5843, n5844, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5856, 
      n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, 
      n5867, n5869, n5870, n5871, n5872, n5874, n5875, n5876, n5877, n5878, 
      n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5888, n5889, 
      n5890, n5891, n5892, n5893, n5895, n5896, n5897, n5900, n5901, n5903, 
      n5904, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, 
      n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5925, n5926, n5929, 
      n5930, n5931, n5932, n5933, n5935, n5936, n5937, n5939, n5940, n5941, 
      n5942, n5944, n5945, n5946, n5948, n5949, n5950, n5951, n5952, n5953, 
      n5954, n5958, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5968, 
      n5969, n5970, n5971, n5972, n5973, n5975, n5976, n5978, n5979, n5980, 
      n5981, n5982, n5983, n5988, n5989, n5990, n5991, n5993, n5994, n5995, 
      n5996, n5997, n5999, n6001, n6003, n6005, n6006, n6007, n6008, n6009, 
      n6010, n6012, n6013, n6014, n6016, n6018, n6020, n6022, n6023, n6024, 
      n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, 
      n6035, n6037, n6039, n6041, n6042, n6043, n6047, n6050, n6051, n6052, 
      n6053, n6054, n6055, n6056, n6058, n6059, n6061, n6062, n6063, n6064, 
      n6067, n6068, n6069, n6071, n6072, n6073, n6074, n6075, n6076, n6078, 
      n6079, n6081, n6082, n6083, n6086, n6087, n6088, n6090, n6091, n6092, 
      n6093, n6094, n6095, n6097, n6098, n6099, n6101, n6102, n6103, n6104, 
      n6105, n6106, n6108, n6109, n6110, n6111, n6114, n6115, n6116, n6117, 
      n6118, n6119, n6121, n6123, n6127, n6129, n6131, n6132, n6133, n6134, 
      n6138, n6142, n6143, n6144, n6145, n6146, n6148, n6149, n6150, n6151, 
      n6152, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, 
      n6165, n6166, n6167, n6168, n6169, n6170, n6172, n6173, n6175, n6176, 
      n6177, n6178, n6179, n6181, n6182, n6183, n6185, n6186, n6187, n6188, 
      n6189, n6190, n6192, n6193, n6198, n6199, n6200, n6203, n6204, n6205, 
      n6206, n6207, n6209, n6211, n6212, n6213, n6215, n6216, n6218, n6219, 
      n6221, n6223, n6225, n6227, n6228, n6229, n6230, n6231, n6232, n6234, 
      n6235, n6236, n6237, n6238, n6242, n6244, n6245, n6247, n6248, n6249, 
      n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6259, n6262, 
      n6263, n6265, n6266, n6267, n6268, n6272, n6273, n6275, n6277, n6280, 
      n6281, n6282, n6283, n6285, n6286, n6287, n6288, n6290, n6293, n6294, 
      n6295, n6297, n6298, n6299, n6300, n6303, n6307, n6308, n6309, n6310, 
      n6311, n6312, n6313, n6316, n6318, n6319, n6320, n6321, n6322, n6324, 
      n6325, n6326, n6327, n6328, n6329, n6332, n6334, n6336, n6337, n6338, 
      n6341, n6342, n6343, n6344, n6345, n6346, n6348, n6350, n6351, n6354, 
      n6357, n6359, n6360, n6362, n6363, n6364, n6365, n6366, n6369, n6370, 
      n6371, n6373, n6376, n6377, n6380, n6382, n6384, n6386, n6387, n6388, 
      n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, 
      n6401, n6402, n6405, n6407, n6408, n6409, n6411, n6414, n6416, n6417, 
      n6420, n6421, n6424, n6425, n6426, n6427, n6428, n6429, n6431, n6432, 
      n6433, n6434, n6435, n6440, n6442, n6444, n6445, n6446, n6447, n6451, 
      n6452, n6453, n6454, n6455, n6457, n6458, n6461, n6462, n6464, n6465, 
      n6466, n6467, n6468, n6469, n6470, n6471, n6473, n6474, n6475, n6476, 
      n6477, n6478, n6479, n6482, n6483, n6484, n6485, n6488, n6489, n6490, 
      n6491, n6493, n6494, n6497, n6500, n6501, n6502, n6503, n6504, n6505, 
      n6507, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6519, n6520, 
      n6524, n6526, n6530, n6531, n6532, n6533, n6536, n6539, n6540, n6543, 
      n6544, n6545, n6547, n6548, n6549, n6551, n6552, n6553, n6555, n6556, 
      n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, 
      n6569, n6570, n6571, n6572, n6574, n6575, n6576, n6577, n6578, n6579, 
      n6580, n6581, n6584, n6587, n6590, n6591, n6592, n6593, n6595, n6597, 
      n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6607, n6608, n6609, 
      n6610, n6611, n6612, n6614, n6615, n6616, n6618, n6619, n6620, n6621, 
      n6624, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, 
      n6637, n6638, n6639, n6640, n6641, n6643, n6644, n6645, n6646, n6647, 
      n6649, n6650, n6651, n6654, n6656, n6657, n6658, n6659, n6660, n6661, 
      n6662, n6663, n6666, n6667, n6668, n6669, n6671, n6672, n6673, n6674, 
      n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, 
      n6685, n6686, n6687, n6688, n6689, n6691, n6693, n6694, n6696, n6698, 
      n6699, n6700, n6701, n6702, n6704, n6705, n6706, n6707, n6708, n6709, 
      n6710, n6711, n6712, n6713, n6716, n6718, n6719, n6720, n6721, n6722, 
      n6723, n6725, n6726, n6728, n6730, n6731, n6733, n6735, n6737, n6739, 
      n6741, n6743, n6745, n6746, n6748, n6749, n6750, n6751, n6753, n6754, 
      n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, 
      n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6775, 
      n6776, n6777, n6778, n6779, n6780, n6782, n6783, n6784, n6786, n6789, 
      n6790, n6791, n6792, n6793, n6794, n6795, n6797, n6798, n6799, n6800, 
      n6801, n6802, n6807, n6808, n6809, n6810, n6811, n6812, n6814, n6816, 
      n6817, n6818, n6819, n6820, n6822, n6824, n6825, n6826, n6827, n6828, 
      n6829, n6830, n6831, n6833, n6835, n6836, n6837, n6840, n6841, n6842, 
      n6843, n6846, n6848, n6849, n6850, n6851, n6852, n6854, n6855, n6856, 
      n6857, n6858, n6859, n6860, n6862, n6863, n6864, n6865, n6866, n6867, 
      n6869, n6872, n6873, n6874, n6876, n6877, n6878, n6879, n6880, n6881, 
      n6882, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6893, n6894, 
      n6895, n6897, n6898, n6899, n6901, n6903, n6904, n6905, n6906, n6907, 
      n6908, n6909, n6910, n6911, n6913, n6914, n6915, n6918, n6919, n6920, 
      n6921, n6923, n6924, n6925, n6926, n6929, n6930, n6931, n6932, n6935, 
      n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6945, n6948, n6950, 
      n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6960, n6961, 
      n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6973, 
      n6974, n6975, n6976, n6978, n6980, n6981, n6982, n6985, n6990, n6992, 
      n6994, n6995, n6996, n6997, n6999, n7001, n7003, n7004, n7005, n7007, 
      n7008, n7011, n7012, n7014, n7015, n7016, n7017, n7018, n7019, n7020, 
      n7022, n7023, n7024, n7025, n7027, n7029, n7030, n7031, n7032, n7033, 
      n7034, n7035, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, 
      n7045, n7046, n7047, n7049, n7050, n7051, n7052, n7053, n7054, n7055, 
      n7056, n7057, n7059, n7060, n7063, n7064, n7065, n7066, n7067, n7068, 
      n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, 
      n7080, n7081, n7083, n7084, n7085, n7086, n7087, n7088, n7090, n7091, 
      n7093, n7094, n7095, n7097, n7098, n7099, n7100, n7101, n7102, n7103, 
      n7105, n7107, n7108, n7109, n7110, n7113, n7114, n7115, n7116, n7118, 
      n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7129, n7131, 
      n7132, n7133, n7134, n7135, n7137, n7138, n7139, n7140, n7141, n7143, 
      n7144, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, 
      n7157, n7160, n7161, n7162, n7163, n7164, n7167, n7169, n7170, n7171, 
      n7173, n7176, n7178, n7179, n7181, n7182, n7183, n7184, n7185, n7186, 
      n7187, n7188, n7190, n7191, n7193, n7194, n7195, n7196, n7197, n7198, 
      n7199, n7200, n7201, n7203, n7204, n7205, n7206, n7207, n7211, n7212, 
      n7213, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7224, n7225, 
      n7226, n7228, n7229, n7232, n7233, n7234, n7235, n7236, n7237, n7238, 
      n7239, n7240, n7241, n7242, n7244, n7245, n7246, n7250, n7251, n7252, 
      n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7261, n7262, n7263, 
      n7265, n7266, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, 
      n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7285, n7286, 
      n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, 
      n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7307, 
      n7308, n7309, n7310, n7312, n7316, n7317, n7318, n7319, n7320, n7323, 
      n7324, n7325, n7326, n7327, n7328, n7330, n7331, n7332, n7334, n7335, 
      n7336, n7339, n7341, n7343, n7344, n7345, n7348, n7349, n7350, n7352, 
      n7356, n7357, n7358, n7360, n7361, n7363, n7365, n7366, n7368, n7369, 
      n7370, n7371, n7373, n7374, n7375, n7376, n7377, n7378, n7380, n7381, 
      n7382, n7383, n7384, n7386, n7387, n7388, n7392, n7394, n7395, n7396, 
      n7397, n7398, n7400, n7402, n7403, n7406, n7407, n7411, n7412, n7413, 
      n7415, n7417, n7418, n7419, n7420, n7425, n7426, n7427, n7429, n7430, 
      n7431, n7432, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7444, 
      n7446, n7447, n7450, n7452, n7453, n7454, n7457, n7458, n7460, n7461, 
      n7462, n7463, n7464, n7465, n7466, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7483, n7485, 
      n7486, n7488, n7490, n7492, n7493, n7495, n7496, n7497, n7501, n7502, 
      n7503, n7504, n7505, n7511, n7512, n7513, n7515, n7516, n7517, n7518, 
      n7520, n7524, n7525, n7526, n7528, n7529, n7530, n7532, n7535, n7537, 
      n7538, n7541, n7543, n7544, n7545, n7546, n7549, n7550, n7551, n7552, 
      n7553, n7554, n7555, n7557, n7559, n7560, n7561, n7562, n7565, n7566, 
      n7568, n7569, n7570, n7572, n7573, n7574, n7575, n7576, n7577, n7579, 
      n7580, n7581, n7582, n7584, n7586, n7589, n7590, n7591, n7592, n7594, 
      n7595, n7596, n7597, n7598, n7599, n7600, n7602, n7603, n7604, n7605, 
      n7606, n7607, n7609, n7610, n7611, n7613, n7614, n7615, n7616, n7619, 
      n7620, n7622, n7623, n7624, n7625, n7626, n7628, n7630, n7631, n7633, 
      n7634, n7635, n7636, n7638, n7639, n7640, n7641, n7643, n7644, n7645, 
      n7646, n7647, n7648, n7649, n7651, n7652, n7653, n7655, n7656, n7657, 
      n7658, n7659, n7660, n7662, n7663, n7664, n7665, n7666, n7667, n7668, 
      n7669, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, 
      n7681, n7682, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7693, 
      n7694, n7695, n7698, n7699, n7700, n7701, n7702, n7703, n7705, n7706, 
      n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7716, n7717, 
      n7719, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7729, n7730, 
      n7731, n7732, n7733, n7736, n7737, n7738, n7741, n7744, n7745, n7746, 
      n7747, n7748, n7749, n7751, n7753, n7754, n7756, n7757, n7759, n7761, 
      n7762, n7765, n7767, n7768, n7770, n7771, n7772, n7773, n7774, n7775, 
      n7776, n7777, n7778, n7779, n7780, n7781, n7785, n7786, n7787, n7789, 
      n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7802, 
      n7803, n7804, n7806, n7808, n7809, n7810, n7811, n7813, n7815, n7817, 
      n7819, n7820, n7822, n7823, n7825, n7826, n7828, n7829, n7830, n7831, 
      n7832, n7834, n7836, n7837, n7838, n7839, n7842, n7843, n7845, n7848, 
      n7850, n7851, n7852, n7853, n7854, n7855, n7857, n7859, n7860, n7861, 
      n7862, n7865, n7866, n7867, n7868, n7870, n7871, n7872, n7873, n7874, 
      n7875, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7887, n7888, 
      n7889, n7890, n7891, n7892, n7893, n7895, n7896, n7897, n7898, n7899, 
      n7900, n7901, n7904, n7905, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7915, n7916, n7917, n7918, n7920, n7921, n7922, n7923, n7924, n7925, 
      n7926, n7928, n7929, n7931, n7933, n7934, n7935, n7936, n7937, n7938, 
      n7939, n7940, n7941, n7942, n7943, n7945, n7946, n7947, n7949, n7951, 
      n7952, n7953, n7954, n7955, n7956, n7957, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7971, n7973, n7974, n7977, 
      n7978, n7984, n7986, n7987, n7988, n7989, n7990, n7991, n7993, n7994, 
      n7995, n7997, n7998, n7999, n8000, n8001, n8003, n8004, n8005, n8006, 
      n8007, n8010, n8011, n8012, n8013, n8015, n8016, n8018, n8020, n8021, 
      n8022, n8024, n8026, n8028, n8029, n8030, n8031, n8033, n8035, n8036, 
      n8037, n8038, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8049, 
      n8050, n8051, n8053, n8054, n8055, n8057, n8058, n8059, n8060, n8061, 
      n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, 
      n8073, n8074, n8076, n8077, n8078, n8079, n8081, n8082, n8083, n8084, 
      n8086, n8087, n8088, n8089, n8091, n8092, n8093, n8094, n8095, n8098, 
      n8099, n8100, n8105, n8106, n8107, n8108, n8109, n8110, n8112, n8113, 
      n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8125, 
      n8126, n8127, n8129, n8130, n8131, n8132, n8133, n8136, n8137, n8138, 
      n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, 
      n8149, n8150, n8152, n8154, n8156, n8160, n8164, n8165, n8166, n8167, 
      n8168, n8170, n8171, n8174, n8175, n8176, n8178, n8181, n8182, n8183, 
      n8184, n8186, n8189, n8190, n8192, n8193, n8194, n8195, n8196, n8197, 
      n8199, n8200, n8201, n8202, n8203, n8204, n8206, n8207, n8208, n8210, 
      n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8219, n8222, n8226, 
      n8227, n8228, n8230, n8232, n8233, n8235, n8236, n8237, n8238, n8241, 
      n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8251, n8252, 
      n8253, n8256, n8257, n8258, n8259, n8260, n8263, n8264, n8265, n8266, 
      n8267, n8268, n8269, n8270, n8271, n8273, n8274, n8275, n8276, n8277, 
      n8278, n8279, n8282, n8283, n8284, n8285, n8286, n8287, n8290, n8291, 
      n8292, n8293, n8294, n8295, n8298, n8299, n8301, n8302, n8303, n8304, 
      n8305, n8306, n8307, n8308, n8309, n8312, n8313, n8314, n8315, n8317, 
      n8318, n8320, n8323, n8324, n8325, n8327, n8328, n8330, n8331, n8332, 
      n8334, n8335, n8336, n8337, n8339, n8340, n8341, n8343, n8344, n8345, 
      n8347, n8348, n8349, n8352, n8353, n8354, n8356, n8358, n8359, n8360, 
      n8361, n8364, n8365, n8366, n8370, n8371, n8372, n8373, n8374, n8376, 
      n8378, n8379, n8380, n8381, n8382, n8383, n8386, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8405, n8406, n8408, n8409, n8411, n8412, n8413, n8415, n8416, n8418, 
      n8420, n8421, n8422, n8424, n8425, n8427, n8431, n8432, n8433, n8434, 
      n8435, n8437, n8438, n8440, n8442, n8443, n8444, n8450, n8452, n8453, 
      n8454, n8455, n8456, n8457, n8459, n8461, n8463, n8464, n8466, n8467, 
      n8468, n8469, n8470, n8471, n8472, n8473, n8475, n8478, n8479, n8480, 
      n8481, n8482, n8485, n8487, n8488, n8489, n8490, n8491, n8492, n8494, 
      n8496, n8497, n8499, n8500, n8502, n8504, n8505, n8506, n8507, n8515, 
      n8519, n8522, n8523, n8525, n8526, n8527, n8528, n8529, n8530, n8531, 
      n8532, n8533, n8535, n8536, n8537, n8539, n8541, n8542, n8543, n8544, 
      n8545, n8547, n8548, n8549, n8550, n8551, n8553, n8554, n8555, n8556, 
      n8557, n8558, n8560, n8561, n8562, n8567, n8568, n8569, n8570, n8571, 
      n8573, n8575, n8576, n8577, n8578, n8579, n8581, n8582, n8583, n8584, 
      n8587, n8589, n8591, n8592, n8593, n8594, n8595, n8596, n8601, n8602, 
      n8603, n8604, n8605, n8606, n8608, n8609, n8611, n8613, n8614, n8615, 
      n8616, n8617, n8618, n8619, n8622, n8625, n8627, n8628, n8629, n8630, 
      n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8639, n8645, n8648, 
      n8650, n8651, n8653, n8654, n8655, n8656, n8657, n8659, n8662, n8663, 
      n8664, n8665, n8666, n8667, n8671, n8672, n8674, n8675, n8676, n8678, 
      n8680, n8681, n8682, n8683, n8684, n8685, n8687, n8689, n8691, n8692, 
      n8694, n8695, n8700, n8701, n8702, n8703, n8705, n8706, n8707, n8708, 
      n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, 
      n8719, n8720, n8721, n8722, n8723, n8726, n8727, n8728, n8731, n8733, 
      n8734, n8735, n8736, n8737, n8739, n8740, n8741, n8742, n8743, n8745, 
      n8746, n8747, n8750, n8753, n8754, n8755, n8756, n8757, n8758, n8759, 
      n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8769, n8770, n8771, 
      n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8780, n8782, n8783, 
      n8784, n8785, n8786, n8787, n8788, n8790, n8791, n8792, n8794, n8795, 
      n8797, n8799, n8800, n8801, n8802, n8804, n8805, n8806, n8808, n8809, 
      n8810, n8811, n8812, n8813, n8816, n8817, n8819, n8820, n8821, n8822, 
      n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8831, n8832, n8834, 
      n8835, n8836, n8838, n8840, n8841, n8843, n8844, n8845, n8846, n8848, 
      n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8860, 
      n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, 
      n8875, n8876, n8882, n8883, n8885, n8886, n8892, n8893, n8894, n8895, 
      n8896, n8897, n8899, n8901, n8902, n8903, n8905, n8906, n8908, n8909, 
      n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, 
      n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, 
      n8930, n8931, n8932, n8933, n8934, n8937, n8939, n8940, n8941, n8942, 
      n8943, n8944, n8946, n8948, n8949, n8950, n8951, n8953, n8954, n8955, 
      n8957, n8958, n8959, n8960, n8962, n8963, n8964, n8965, n8966, n8967, 
      n8968, n8970, n8972, n8973, n8974, n8975, n8976, n8979, n8980, n8983, 
      n8984, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, 
      n8996, n8997, n8998, n9000, n9002, n9003, n9004, n9005, n9006, n9010, 
      n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9020, n9021, 
      n9022, n9025, n9026, n9027, n9028, n9030, n9031, n9032, n9033, n9037, 
      n9038, n9040, n9041, n9042, n9044, n9045, n9046, n9050, n9052, n9055, 
      n9057, n9058, n9059, n9062, n9064, n9065, n9066, n9068, n9071, n9073, 
      n9075, n9076, n9078, n9080, n9083, n9085, n9087, n9088, n9090, n9092, 
      n9093, n9095, n9097, n9098, n9099, n9101, n9102, n9103, n9105, n9106, 
      n9107, n9108, n9110, n9111, n9113, n9114, n9115, n9116, n9118, n9119, 
      n9120, n9121, n9123, n9125, n9126, n9127, n9129, n9131, n9133, n9134, 
      n9135, n9136, n9137, n9138, n9139, n9141, n9145, n9146, n9147, n9148, 
      n9149, n9151, n9152, n9153, n9154, n9155, n9156, n9158, n9159, n9160, 
      n9161, n9162, n9163, n9164, n9166, n9167, n9168, n9170, n9171, n9172, 
      n9173, n9174, n9176, n9177, n9178, n9180, n9181, n9182, n9183, n9184, 
      n9185, n9186, n9189, n9191, n9192, n9193, n9195, n9197, n9198, n9199, 
      n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, 
      n9211, n9212, n9213, n9214, n9215, n9217, n9218, n9219, n9220, n9221, 
      n9222, n9223, n9224, n9225, n9227, n9228, n9230, n9231, n9232, n9233, 
      n9234, n9235, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, 
      n9247, n9248, n9249, n9251, n9252, n9255, n9256, n9257, n9258, n9259, 
      n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9269, n9270, n9271, 
      n9272, n9273, n9274, n9275, n9277, n9278, n9280, n9281, n9282, n9283, 
      n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9292, n9293, n9294, 
      n9296, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9307, 
      n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, 
      n9318, n9319, n9320, n9322, n9323, n9324, n9325, n9326, n9327, n9328, 
      n9329, n9334, n9335, n9338, n9339, n9341, n9342, n9343, n9344, n9345, 
      n9346, n9347, n9349, n9350, n9351, n9352, n9353, n9356, n9361, n9362, 
      n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9373, n9374, 
      n9375, n9377, n9378, n9379, n9381, n9382, n9383, n9384, n9385, n9386, 
      n9387, n9388, n9390, n9391, n9392, n9393, n9395, n9396, n9397, n9398, 
      n9399, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9411, 
      n9412, n9413, n9414, n9418, n9419, n9420, n9422, n9423, n9424, n9425, 
      n9426, n9427, n9428, n9430, n9432, n9434, n9435, n9436, n9437, n9438, 
      n9439, n9440, n9441, n9442, n9443, n9444, n9446, n9447, n9448, n9449, 
      n9450, n9451, n9452, n9453, n9454, n9456, n9459, n9460, n9462, n9464, 
      n9467, n9468, n9469, n9472, n9473, n9474, n9475, n9476, n9478, n9479, 
      n9480, n9481, n9483, n9484, n9485, n9486, n9487, n9488, n9490, n9493, 
      n9495, n9496, n9500, n9502, n9503, n9504, n9505, n9506, n9507, n9508, 
      n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, 
      n9521, n9522, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, 
      n9535, n9536, n9538, n9539, n9540, n9542, n9544, n9545, n9546, n9547, 
      n9548, n9549, n9550, n9551, n9552, n9553, n9555, n9558, n9560, n9561, 
      n9563, n9564, n9567, n9568, n9569, n9571, n9573, n9574, n9575, n9577, 
      n9578, n9579, n9580, n9581, n9582, n9584, n9585, n9586, n9587, n9588, 
      n9589, n9590, n9591, n9592, n9593, n9597, n9599, n9601, n9603, n9604, 
      n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9615, n9616, 
      n9617, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, 
      n9629, n9630, n9631, n9634, n9635, n9636, n9637, n9640, n9641, n9644, 
      n9645, n9646, n9647, n9648, n9650, n9651, n9652, n9653, n9654, n9655, 
      n9658, n9659, n9660, n9661, n9663, n9664, n9665, n9666, n9667, n9668, 
      n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, 
      n9681, n9683, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, 
      n9694, n9695, n9696, n9697, n9698, n9699, n9701, n9703, n9704, n9705, 
      n9706, n9708, n9709, n9710, n9711, n9714, n9717, n9718, n9719, n9721, 
      n9724, n9725, n9728, n9729, n9731, n9732, n9733, n9734, n9736, n9737, 
      n9738, n9739, n9740, n9741, n9744, n9747, n9748, n9749, n9750, n9751, 
      n9752, n9753, n9754, n9757, n9758, n9759, n9760, n9761, n9762, n9764, 
      n9766, n9768, n9769, n9770, n9772, n9773, n9774, n9775, n9776, n9777, 
      n9778, n9780, n9781, n9782, n9783, n9785, n9786, n9787, n9788, n9789, 
      n9790, n9791, n9792, n9793, n9794, n9796, n9797, n9798, n9800, n9801, 
      n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, 
      n9812, n9813, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, 
      n9823, n9824, n9825, n9826, n9828, n9831, n9832, n9833, n9835, n9836, 
      n9837, n9838, n9839, n9840, n9842, n9843, n9844, n9846, n9847, n9848, 
      n9852, n9854, n9855, n9856, n9857, n9858, n9859, n9861, n9862, n9863, 
      n9865, n9866, n9867, n9868, n9870, n9871, n9874, n9875, n9876, n9877, 
      n9878, n9879, n9880, n9884, n9885, n9886, n9887, n9889, n9890, n9892, 
      n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, 
      n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9913, 
      n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9928, n9929, n9930, 
      n9931, n9932, n9933, n9934, n9936, n9937, n9939, n9941, n9943, n9945, 
      n9946, n9949, n9950, n9951, n9953, n9954, n9955, n9956, n9957, n9958, 
      n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, 
      n9969, n9973, n9975, n9976, n9977, n9978, n9980, n9981, n9982, n9983, 
      n9984, n9985, n9986, n9988, n9990, n9991, n9992, n9993, n9994, n9995, 
      n9998, n9999, n10000, n10001, n10003, n10004, n10005, n10006, n10007, 
      n10009, n10010, n10011, n10012, n10013, n10015, n10017, n10018, n10019, 
      n10020, n10024, n10026, n10028, n10030, n10031, n10033, n10035, n10038, 
      n10039, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10051, 
      n10052, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10062, 
      n10063, n10064, n10066, n10068, n10069, n10070, n10071, n10072, n10073, 
      n10074, n10075, n10076, n10077, n10079, n10080, n10081, n10082, n10084, 
      n10085, n10086, n10087, n10088, n10089, n10090, n10092, n10093, n10095, 
      n10096, n10097, n10098, n10099, n10100, n10103, n10104, n10105, n10106, 
      n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10116, 
      n10117, n10118, n10119, n10121, n10122, n10123, n10124, n10125, n10126, 
      n10127, n10128, n10129, n10130, n10132, n10133, n10134, n10135, n10136, 
      n10137, n10138, n10140, n10142, n10143, n10145, n10146, n10148, n10149, 
      n10150, n10152, n10154, n10155, n10157, n10159, n10160, n10163, n10164, 
      n10165, n10166, n10167, n10169, n10170, n10171, n10172, n10173, n10174, 
      n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, 
      n10184, n10186, n10187, n10188, n10192, n10193, n10194, n10195, n10196, 
      n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10205, n10206, 
      n10207, n10208, n10209, n10210, n10213, n10214, n10215, n10216, n10217, 
      n10218, n10219, n10220, n10221, n10224, n10226, n10227, n10228, n10229, 
      n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10241, n10243, 
      n10244, n10247, n10248, n10249, n10251, n10252, n10254, n10255, n10257, 
      n10258, n10259, n10260, n10261, n10262, n10264, n10265, n10266, n10268, 
      n10270, n10271, n10272, n10273, n10276, n10277, n10278, n10279, n10280, 
      n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, 
      n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10301, 
      n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10310, n10312, 
      n10313, n10314, n10315, n10316, n10317, n10320, n10321, n10322, n10323, 
      n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, 
      n10335, n10337, n10339, n10340, n10342, n10343, n10344, n10345, n10346, 
      n10347, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10357, 
      n10358, n10359, n10360, n10361, n10364, n10365, n10366, n10367, n10369, 
      n10370, n10371, n10372, n10373, n10374, n10376, n10379, n10380, n10381, 
      n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, 
      n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, 
      n10401, n10402, n10404, n10405, n10409, n10410, n10411, n10412, n10413, 
      n10414, n10416, n10419, n10420, n10421, n10422, n10423, n10424, n10426, 
      n10427, n10428, n10429, n10430, n10431, n10433, n10434, n10435, n10436, 
      n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10446, 
      n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10456, n10459, 
      n10460, n10461, n10462, n10463, n10465, n10466, n10467, n10468, n10469, 
      n10470, n10472, n10473, n10474, n10475, n10478, n10480, n10481, n10482, 
      n10483, n10484, n10485, n10486, n10488, n10489, n10490, n10491, n10492, 
      n10493, n10495, n10496, n10497, n10498, n10500, n10501, n10504, n10505, 
      n10507, n10508, n10510, n10511, n10513, n10514, n10515, n10516, n10519, 
      n10522, n10523, n10524, n10525, n10527, n10528, n10529, n10530, n10531, 
      n10532, n10533, n10535, n10536, n10537, n10539, n10542, n10546, n10547, 
      n10548, n10549, n10550, n10552, n10553, n10555, n10556, n10557, n10558, 
      n10560, n10561, n10564, n10565, n10566, n10567, n10568, n10569, n10570, 
      n10571, n10572, n10573, n10574, n10576, n10578, n10579, n10581, n10582, 
      n10583, n10584, n10585, n10587, n10588, n10589, n10598, n10599, n10600, 
      n10603, n10604, n10605, n10606, n10608, n10609, n10611, n10612, n10613, 
      n10614, n10615, n10616, n10617, n10619, n10620, n10621, n10622, n10623, 
      n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10637, 
      n10638, n10639, n10640, n10641, n10643, n10644, n10645, n10646, n10649, 
      n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, 
      n10659, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10669, 
      n10670, n10671, n10673, n10674, n10675, n10679, n10680, n10681, n10683, 
      n10685, n10686, n10687, n10689, n10693, n10694, n10695, n10696, n10697, 
      n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10707, n10708, 
      n10710, n10713, n10714, n10715, n10716, n10717, n10718, n10720, n10721, 
      n10722, n10723, n10724, n10725, n10727, n10728, n10729, n10730, n10731, 
      n10732, n10733, n10735, n10737, n10738, n10739, n10740, n10741, n10742, 
      n10743, n10744, n10745, n10747, n10748, n10749, n10750, n10752, n10753, 
      n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10762, n10763, 
      n10764, n10765, n10766, n10768, n10769, n10770, n10772, n10773, n10775, 
      n10776, n10777, n10778, n10780, n10783, n10784, n10785, n10786, n10787, 
      n10788, n10789, n10790, n10791, n10792, n10793, n10796, n10797, n10798, 
      n10799, n10800, n10804, n10805, n10806, n10808, n10809, n10810, n10811, 
      n10812, n10813, n10814, n10815, n10816, n10821, n10822, n10823, n10824, 
      n10825, n10827, n10828, n10829, n10831, n10832, n10833, n10834, n10835, 
      n10837, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, 
      n10849, n10850, n10853, n10854, n10855, n10856, n10857, n10858, n10859, 
      n10860, n10861, n10862, n10863, n10865, n10866, n10867, n10868, n10869, 
      n10870, n10871, n10872, n10873, n10874, n10875, n10877, n10878, n10883, 
      n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10895, 
      n10896, n10897, n10899, n10900, n10901, n10902, n10903, n10904, n10905, 
      n10907, n10908, n10909, n10910, n10914, n10915, n10916, n10917, n10921, 
      n10922, n10923, n10924, n10925, n10926, n10928, n10931, n10932, n10934, 
      n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, 
      n10944, n10945, n10946, n10947, n10948, n10949, n10951, n10953, n10954, 
      n10955, n10959, n10960, n10961, n10963, n10964, n10965, n10966, n10967, 
      n10968, n10970, n10971, n10972, n10973, n10974, n10975, n10977, n10978, 
      n10979, n10980, n10985, n10986, n10987, n10989, n10990, n10991, n10992, 
      n10993, n10999, n11000, n11003, n11004, n11005, n11006, n11008, n11010, 
      n11011, n11012, n11013, n11017, n11018, n11019, n11020, n11022, n11023, 
      n11027, n11028, n11031, n11033, n11034, n11035, n11036, n11037, n11038, 
      n11039, n11041, n11042, n11045, n11046, n11048, n11049, n11050, n11051, 
      n11052, n11053, n11055, n11057, n11058, n11059, n11061, n11062, n11063, 
      n11064, n11066, n11067, n11068, n11069, n11070, n11072, n11074, n11075, 
      n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, 
      n11086, n11089, n11090, n11091, n11092, n11093, n11095, n11096, n11097, 
      n11098, n11100, n11102, n11103, n11104, n11105, n11106, n11107, n11108, 
      n11109, n11110, n11111, n11112, n11113, n11118, n11119, n11120, n11121, 
      n11122, n11123, n11124, n11126, n11128, n11129, n11130, n11131, n11132, 
      n11133, n11134, n11135, n11136, n11138, n11139, n11140, n11141, n11142, 
      n11143, n11144, n11146, n11147, n11148, n11149, n11150, n11151, n11152, 
      n11153, n11155, n11156, n11157, n11158, n11159, n11161, n11162, n11164, 
      n11166, n11167, n11169, n11170, n11171, n11172, n11173, n11175, n11177, 
      n11178, n11179, n11180, n11181, n11182, n11185, n11186, n11187, n11192, 
      n11193, n11194, n11195, n11198, n11199, n11200, n11201, n11202, n11203, 
      n11204, n11205, n11206, n11208, n11210, n11211, n11212, n11213, n11214, 
      n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, 
      n11225, n11227, n11228, n11229, n11231, n11232, n11235, n11236, n11238, 
      n11240, n11241, n11243, n11244, n11245, n11246, n11247, n11248, n11249, 
      n11250, n11251, n11253, n11254, n11255, n11257, n11258, n11259, n11261, 
      n11262, n11263, n11264, n11265, n11266, n11268, n11269, n11270, n11271, 
      n11272, n11276, n11278, n11280, n11281, n11282, n11285, n11287, n11289, 
      n11290, n11291, n11292, n11294, n11295, n11297, n11298, n11299, n11300, 
      n11301, n11302, n11303, n11304, n11306, n11308, n11309, n11310, n11311, 
      n11312, n11315, n11317, n11318, n11319, n11320, n11321, n11322, n11323, 
      n11324, n11325, n11326, n11327, n11330, n11331, n11332, n11333, n11334, 
      n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11346, n11347, 
      n11348, n11349, n11350, n11351, n11353, n11354, n11355, n11356, n11357, 
      n11358, n11359, n11360, n11361, n11362, n11364, n11365, n11366, n11368, 
      n11370, n11372, n11374, n11376, n11378, n11379, n11380, n11381, n11382, 
      n11383, n11385, n11387, n11388, n11389, n11390, n11391, n11392, n11393, 
      n11394, n11396, n11397, n11398, n11399, n11401, n11402, n11405, n11406, 
      n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11416, n11418, 
      n11419, n11420, n11421, n11422, n11423, n11424, n11426, n11427, n11428, 
      n11429, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, 
      n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, 
      n11450, n11451, n11452, n11453, n11454, n11456, n11457, n11458, n11459, 
      n11460, n11461, n11463, n11464, n11465, n11466, n11467, n11468, n11469, 
      n11470, n11474, n11475, n11476, n11477, n11480, n11481, n11483, n11484, 
      n11485, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, 
      n11495, n11497, n11499, n11500, n11501, n11502, n11503, n11504, n11505, 
      n11507, n11508, n11510, n11511, n11512, n11513, n11514, n11515, n11516, 
      n11517, n11518, n11519, n11521, n11522, n11523, n11524, n11525, n11526, 
      n11527, n11528, n11529, n11530, n11531, n11532, n11534, n11535, n11536, 
      n11537, n11538, n11539, n11540, n11542, n11543, n11544, n11545, n11548, 
      n11551, n11552, n11555, n11556, n11557, n11558, n11559, n11560, n11562, 
      n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, 
      n11574, n11575, n11576, n11577, n11578, n11580, n11581, n11582, n11584, 
      n11585, n11586, n11587, n11589, n11590, n11591, n11593, n11595, n11596, 
      n11597, n11599, n11600, n11601, n11603, n11604, n11605, n11608, n11610, 
      n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, 
      n11620, n11621, n11622, n11623, n11624, n11626, n11627, n11628, n11629, 
      n11630, n11631, n11633, n11634, n11635, n11636, n11637, n11640, n11641, 
      n11643, n11644, n11645, n11646, n11651, n11652, n11653, n11654, n11655, 
      n11656, n11657, n11658, n11659, n11660, n11661, n11663, n11665, n11666, 
      n11667, n11668, n11669, n11670, n11673, n11675, n11676, n11677, n11678, 
      n11680, n11681, n11682, n11683, n11684, n11686, n11687, n11688, n11689, 
      n11690, n11691, n11693, n11694, n11695, n11696, n11697, n11698, n11699, 
      n11700, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, 
      n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, 
      n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, 
      n11730, n11732, n11733, n11734, n11735, n11736, n11737, n11740, n11741, 
      n11742, n11743, n11744, n11745, n11746, n11748, n11749, n11750, n11751, 
      n11752, n11754, n11755, n11756, n11757, n11759, n11760, n11761, n11762, 
      n11765, n11766, n11767, n11768, n11769, n11770, n11773, n11774, n11775, 
      n11776, n11777, n11778, n11780, n11781, n11782, n11783, n11784, n11785, 
      n11786, n11788, n11789, n11792, n11795, n11796, n11797, n11798, n11800, 
      n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, 
      n11812, n11814, n11815, n11816, n11817, n11819, n11820, n11821, n11822, 
      n11823, n11824, n11826, n11827, n11828, n11829, n11830, n11831, n11832, 
      n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, 
      n11842, n11843, n11844, n11845, n11847, n11848, n11850, n11852, n11853, 
      n11854, n11855, n11856, n11859, n11860, n11861, n11862, n11863, n11864, 
      n11865, n11866, n11867, n11868, n11869, n11871, n11872, n11873, n11874, 
      n11875, n11876, n11877, n11880, n11883, n11884, n11887, n11888, n11889, 
      n11890, n11891, n11892, n11893, n11895, n11897, n11898, n11899, n11900, 
      n11902, n11903, n11904, n11905, n11907, n11909, n11910, n11911, n11912, 
      n11913, n11915, n11916, n11917, n11918, n11919, n11920, n11922, n11923, 
      n11924, n11925, n11926, n11928, n11929, n11930, n11931, n11932, n11933, 
      n11934, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, 
      n11945, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, 
      n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, 
      n11964, n11966, n11967, n11968, n11969, n11970, n11971, n11973, n11974, 
      n11975, n11976, n11977, n11979, n11980, n11981, n11982, n11983, n11984, 
      n11985, n11986, n11987, n11988, n11990, n11991, n11992, n11994, n11995, 
      n11996, n11997, n11998, n11999, n12000, n12002, n12004, n12005, n12006, 
      n12008, n12010, n12011, n12013, n12014, n12016, n12017, n12018, n12019, 
      n12020, n12021, n12022, n12025, n12026, n12027, n12028, n12029, n12030, 
      n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, 
      n12040, n12041, n12042, n12043, n12044, n12045, n12048, n12049, n12051, 
      n12052, n12053, n12054, n12055, n12057, n12058, n12059, n12060, n12061, 
      n12062, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, 
      n12074, n12075, n12076, n12077, n12078, n12080, n12082, n12083, n12084, 
      n12085, n12086, n12088, n12089, n12090, n12091, n12093, n12094, n12095, 
      n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, 
      n12107, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12118, 
      n12119, n12120, n12121, n12122, n12123, n12124, n12127, n12128, n12130, 
      n12131, n12132, n12133, n12135, n12136, n12137, n12139, n12140, n12141, 
      n12142, n12143, n12144, n12145, n12147, n12148, n12149, n12150, n12151, 
      n12153, n12154, n12156, n12157, n12159, n12160, n12161, n12163, n12164, 
      n12165, n12166, n12168, n12169, n12170, n12171, n12172, n12173, n12174, 
      n12175, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, 
      n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, 
      n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, 
      n12208, n12209, n12211, n12212, n12213, n12214, n12215, n12217, n12218, 
      n12220, n12221, n12223, n12224, n12225, n12226, n12227, n12228, n12229, 
      n12230, n12231, n12232, n12235, n12236, n12237, n12238, n12239, n12240, 
      n12241, n12243, n12244, n12247, n12248, n12249, n12250, n12251, n12252, 
      n12253, n12254, n12256, n12257, n12258, n12259, n12260, n12262, n12263, 
      n12264, n12265, n12266, n12268, n12270, n12271, n12272, n12273, n12274, 
      n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, 
      n12284, n12285, n12286, n12287, n12288, n12290, n12291, n12293, n12295, 
      n12296, n12297, n12300, n12302, n12304, n12308, n12309, n12310, n12312, 
      n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12322, 
      n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, 
      n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12340, n12341, 
      n12342, n12343, n12344, n12345, n12347, n12348, n12351, n12353, n12354, 
      n12355, n12356, n12357, n12358, n12359, n12363, n12364, n12365, n12366, 
      n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, 
      n12376, n12377, n12379, n12380, n12381, n12382, n12383, n12384, n12386, 
      n12387, n12390, n12391, n12392, n12394, n12395, n12396, n12397, n12398, 
      n12399, n12402, n12403, n12407, n12408, n12409, n12410, n12411, n12413, 
      n12414, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, 
      n12424, n12429, n12430, n12431, n12432, n12433, n12434, n12439, n12440, 
      n12441, n12442, n12443, n12444, n12445, n12446, n12448, n12449, n12450, 
      n12452, n12453, n12454, n12456, n12457, n12458, n12459, n12461, n12462, 
      n12465, n12467, n12468, n12469, n12471, n12472, n12473, n12474, n12475, 
      n12476, n12478, n12479, n12482, n12485, n12486, n12487, n12488, n12490, 
      n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12500, 
      n12502, n12504, n12505, n12506, n12507, n12508, n12509, n12511, n12512, 
      n12513, n12514, n12515, n12516, n12517, n12519, n12520, n12521, n12522, 
      n12525, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, 
      n12535, n12536, n12538, n12539, n12540, n12541, n12542, n12545, n12546, 
      n12547, n12548, n12549, n12551, n12552, n12553, n12556, n12557, n12559, 
      n12561, n12562, n12563, n12564, n12565, n12567, n12568, n12570, n12572, 
      n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12582, 
      n12583, n12584, n12585, n12586, n12587, n12590, n12592, n12593, n12594, 
      n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, 
      n12604, n12605, n12609, n12610, n12611, n12613, n12614, n12615, n12616, 
      n12617, n12618, n12619, n12620, n12621, n12622, n12624, n12625, n12626, 
      n12627, n12628, n12629, n12632, n12634, n12636, n12637, n12640, n12641, 
      n12642, n12643, n12644, n12645, n12646, n12648, n12649, n12650, n12651, 
      n12652, n12653, n12654, n12657, n12658, n12659, n12662, n12663, n12665, 
      n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, 
      n12678, n12679, n12680, n12681, n12682, n12683, n12686, n12687, n12688, 
      n12689, n12690, n12691, n12692, n12693, n12695, n12696, n12697, n12698, 
      n12699, n12700, n12701, n12702, n12704, n12705, n12707, n12708, n12711, 
      n12712, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, 
      n12722, n12724, n12725, n12726, n12727, n12728, n12729, n12731, n12732, 
      n12733, n12735, n12736, n12738, n12742, n12743, n12744, n12746, n12747, 
      n12748, n12749, n12750, n12751, n12753, n12754, n12755, n12756, n12757, 
      n12758, n12759, n12760, n12762, n12763, n12764, n12765, n12768, n12770, 
      n12771, n12774, n12775, n12777, n12779, n12781, n12782, n12783, n12784, 
      n12785, n12786, n12787, n12788, n12789, n12790, n12792, n12793, n12794, 
      n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12803, n12804, 
      n12805, n12807, n12808, n12809, n12811, n12812, n12813, n12814, n12815, 
      n12816, n12817, n12821, n12823, n12824, n12826, n12827, n12828, n12830, 
      n12831, n12832, n12836, n12837, n12840, n12841, n12843, n12844, n12845, 
      n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12855, 
      n12856, n12858, n12861, n12862, n12863, n12864, n12865, n12866, n12868, 
      n12869, n12871, n12872, n12873, n12875, n12876, n12877, n12878, n12879, 
      n12880, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12891, 
      n12892, n12894, n12895, n12896, n12898, n12899, n12900, n12902, n12903, 
      n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, 
      n12913, n12915, n12916, n12917, n12918, n12919, n12921, n12922, n12923, 
      n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, 
      n12933, n12934, n12935, n12936, n12937, n12939, n12942, n12943, n12944, 
      n12945, n12947, n12948, n12950, n12951, n12952, n12954, n12955, n12956, 
      n12957, n12958, n12959, n12960, n12962, n12966, n12968, n12969, n12971, 
      n12972, n12973, n12974, n12975, n12976, n12977, n12980, n12981, n12982, 
      n12983, n12985, n12986, n12987, n12989, n12991, n12992, n12993, n12994, 
      n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, 
      n13004, n13006, n13008, n13009, n13011, n13012, n13013, n13014, n13015, 
      n13016, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13028, 
      n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, 
      n13040, n13041, n13042, n13043, n13045, n13046, n13047, n13048, n13049, 
      n13050, n13051, n13052, n13053, n13055, n13056, n13058, n13059, n13060, 
      n13061, n13063, n13065, n13066, n13067, n13068, n13070, n13071, n13072, 
      n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13082, 
      n13083, n13084, n13085, n13086, n13087, n13089, n13090, n13091, n13092, 
      n13093, n13095, n13099, n13100, n13101, n13102, n13103, n13104, n13105, 
      n13106, n13107, n13109, n13110, n13111, n13112, n13113, n13114, n13115, 
      n13116, n13120, n13121, n13122, n13123, n13124, n13125, n13127, n13129, 
      n13130, n13131, n13132, n13133, n13136, n13137, n13138, n13139, n13140, 
      n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, 
      n13151, n13152, n13154, n13157, n13159, n13160, n13161, n13162, n13163, 
      n13167, n13168, n13169, n13170, n13172, n13173, n13175, n13176, n13177, 
      n13178, n13179, n13180, n13181, n13185, n13186, n13187, n13188, n13189, 
      n13190, n13191, n13193, n13194, n13195, n13196, n13197, n13198, n13199, 
      n13200, n13201, n13202, n13204, n13205, n13208, n13209, n13210, n13212, 
      n13213, n13214, n13216, n13217, n13219, n13222, n13223, n13224, n13226, 
      n13227, n13230, n13231, n13232, n13234, n13235, n13236, n13237, n13238, 
      n13239, n13242, n13243, n13245, n13246, n13247, n13248, n13249, n13251, 
      n13252, n13253, n13254, n13255, n13258, n13260, n13261, n13262, n13263, 
      n13265, n13266, n13267, n13268, n13272, n13273, n13274, n13275, n13276, 
      n13279, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, 
      n13289, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, 
      n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13308, 
      n13309, n13310, n13312, n13313, n13314, n13315, n13316, n13318, n13319, 
      n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, 
      n13329, n13330, n13331, n13332, n13334, n13336, n13338, n13339, n13340, 
      n13341, n13342, n13343, n13345, n13346, n13347, n13348, n13349, n13353, 
      n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13363, 
      n13364, n13365, n13366, n13367, n13369, n13370, n13371, n13372, n13373, 
      n13374, n13375, n13377, n13378, n13379, n13380, n13381, n13382, n13384, 
      n13386, n13388, n13389, n13390, n13391, n13393, n13394, n13395, n13396, 
      n13397, n13401, n13402, n13403, n13404, n13405, n13407, n13408, n13409, 
      n13411, n13412, n13413, n13414, n13415, n13417, n13419, n13421, n13422, 
      n13423, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, 
      n13433, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, 
      n13444, n13445, n13448, n13449, n13450, n13451, n13452, n13453, n13454, 
      n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13464, 
      n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, 
      n13475, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13485, 
      n13488, n13489, n13490, n13491, n13494, n13495, n13496, n13497, n13498, 
      n13499, n13500, n13501, n13502, n13503, n13504, n13506, n13507, n13508, 
      n13509, n13510, n13511, n13513, n13514, n13517, n13519, n13520, n13521, 
      n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, 
      n13534, n13535, n13537, n13538, n13539, n13540, n13541, n13544, n13545, 
      n13546, n13547, n13548, n13549, n13551, n13552, n13553, n13554, n13555, 
      n13556, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, 
      n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, 
      n13575, n13576, n13578, n13579, n13580, n13581, n13582, n13583, n13585, 
      n13586, n13587, n13589, n13590, n13591, n13592, n13593, n13595, n13596, 
      n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13605, n13606, 
      n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, 
      n13617, n13618, n13619, n13621, n13622, n13623, n13624, n13627, n13628, 
      n13629, n13630, n13631, n13632, n13633, n13635, n13636, n13637, n13638, 
      n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, 
      n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, 
      n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, 
      n13667, n13668, n13669, n13670, n13673, n13677, n13678, n13679, n13680, 
      n13681, n13682, n13684, n13685, n13686, n13689, n13690, n13692, n13693, 
      n13694, n13695, n13696, n13698, n13700, n13702, n13703, n13704, n13705, 
      n13706, n13707, n13708, n13709, n13710, n13712, n13716, n13719, n13720, 
      n13721, n13723, n13724, n13725, n13727, n13730, n13732, n13733, n13735, 
      n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13745, 
      n13746, n13747, n13748, n13751, n13752, n13759, n13760, n13762, n13763, 
      n13764, n13765, n13766, n13767, n13768, n13770, n13771, n13772, n13773, 
      n13774, n13777, n13778, n13780, n13782, n13783, n13784, n13785, n13786, 
      n13787, n13788, n13791, n13792, n13793, n13794, n13796, n13800, n13802, 
      n13803, n13804, n13806, n13807, n13809, n13810, n13811, n13812, n13814, 
      n13815, n13816, n13817, n13819, n13822, n13824, n13825, n13826, n13828, 
      n13829, n13830, n13831, n13833, n13834, n13835, n13837, n13838, n13839, 
      n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13849, n13850, 
      n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, 
      n13860, n13861, n13862, n13863, n13864, n13865, n13867, n13869, n13872, 
      n13873, n13874, n13876, n13877, n13878, n13879, n13880, n13881, n13883, 
      n13884, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, 
      n13894, n13895, n13896, n13898, n13899, n13901, n13902, n13903, n13904, 
      n13905, n13906, n13907, n13908, n13909, n13911, n13912, n13913, n13914, 
      n13915, n13916, n13917, n13918, n13920, n13921, n13922, n13924, n13925, 
      n13927, n13928, n13930, n13931, n13932, n13933, n13934, n13935, n13936, 
      n13937, n13938, n13939, n13940, n13941, n13943, n13944, n13945, n13946, 
      n13947, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, 
      n13957, n13960, n13962, n13963, n13965, n13966, n13968, n13969, n13970, 
      n13971, n13972, n13973, n13974, n13975, n13977, n13978, n13979, n13981, 
      n13982, n13983, n13984, n13985, n13986, n13987, n13989, n13993, n13994, 
      n13995, n13996, n13998, n14000, n14001, n14002, n14004, n14005, n14008, 
      n14009, n14010, n14011, n14012, n14014, n14016, n14017, n14019, n14020, 
      n14021, n14022, n14023, n14024, n14027, n14029, n14030, n14031, n14032, 
      n14033, n14034, n14036, n14037, n14038, n14039, n14041, n14042, n14043, 
      n14044, n14045, n14047, n14049, n14050, n14051, n14052, n14053, n14054, 
      n14055, n14056, n14058, n14060, n14062, n14065, n14066, n14067, n14069, 
      n14070, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, 
      n14082, n14083, n14084, n14086, n14087, n14088, n14091, n14092, n14093, 
      n14094, n14095, n14098, n14099, n14100, n14101, n14102, n14103, n14104, 
      n14106, n14107, n14108, n14110, n14111, n14112, n14113, n14114, n14117, 
      n14118, n14119, n14120, n14122, n14123, n14124, n14125, n14126, n14129, 
      n14130, n14131, n14132, n14133, n14134, n14136, n14137, n14138, n14139, 
      n14142, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14153, 
      n14154, n14155, n14156, n14157, n14159, n14160, n14161, n14162, n14163, 
      n14164, n14166, n14168, n14170, n14171, n14172, n14173, n14174, n14176, 
      n14177, n14178, n14179, n14181, n14183, n14184, n14187, n14188, n14189, 
      n14190, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, 
      n14201, n14202, n14203, n14206, n14207, n14208, n14209, n14210, n14211, 
      n14212, n14213, n14214, n14215, n14216, n14217, n14219, n14220, n14221, 
      n14222, n14223, n14227, n14228, n14230, n14231, n14232, n14233, n14234, 
      n14236, n14237, n14238, n14239, n14242, n14243, n14244, n14245, n14246, 
      n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14255, n14257, 
      n14258, n14259, n14261, n14262, n14263, n14264, n14265, n14266, n14267, 
      n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14276, n14277, 
      n14279, n14280, n14281, n14282, n14283, n14284, n14288, n14289, n14290, 
      n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, 
      n14301, n14305, n14306, n14307, n14308, n14309, n14311, n14312, n14314, 
      n14315, n14316, n14318, n14320, n14321, n14322, n14325, n14326, n14327, 
      n14328, n14329, n14331, n14332, n14334, n14335, n14336, n14337, n14339, 
      n14340, n14342, n14344, n14346, n14348, n14349, n14350, n14352, n14354, 
      n14355, n14359, n14361, n14362, n14363, n14364, n14365, n14366, n14367, 
      n14368, n14369, n14370, n14371, n14373, n14375, n14376, n14381, n14382, 
      n14383, n14384, n14385, n14386, n14387, n14388, n14391, n14392, n14393, 
      n14394, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14404, 
      n14407, n14409, n14410, n14411, n14412, n14415, n14416, n14417, n14418, 
      n14419, n14420, n14422, n14423, n14424, n14425, n14426, n14428, n14429, 
      n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, 
      n14442, n14443, n14444, n14445, n14447, n14449, n14450, n14451, n14453, 
      n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14463, 
      n14464, n14465, n14466, n14470, n14471, n14472, n14473, n14478, n14479, 
      n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, 
      n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, 
      n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, 
      n14509, n14510, n14511, n14513, n14514, n14516, n14517, n14518, n14519, 
      n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14529, n14530, 
      n14531, n14532, n14533, n14534, n14536, n14537, n14539, n14540, n14541, 
      n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14550, n14551, 
      n14552, n14555, n14556, n14557, n14559, n14560, n14561, n14562, n14563, 
      n14564, n14565, n14566, n14567, n14568, n14571, n14572, n14573, n14574, 
      n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, 
      n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, 
      n14593, n14594, n14595, n14597, n14598, n14600, n14601, n14602, n14603, 
      n14605, n14606, n14607, n14609, n14610, n14611, n14612, n14613, n14614, 
      n14615, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, 
      n14625, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, 
      n14635, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, 
      n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, 
      n14654, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, 
      n14664, n14665, n14666, n14667, n14668, n14671, n14673, n14674, n14676, 
      n14677, n14678, n14680, n14681, n14682, n14683, n14684, n14685, n14686, 
      n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, 
      n14698, n14699, n14701, n14702, n14703, n14704, n14705, n14706, n14708, 
      n14709, n14710, n14711, n14712, n14713, n14716, n14717, n14719, n14720, 
      n14721, n14722, n14724, n14725, n14726, n14727, n14728, n14729, n14730, 
      n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, 
      n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, 
      n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, 
      n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, 
      n14770, n14772, n14773, n14774, n14775, n14776, n14778, n14779, n14780, 
      n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, 
      n14791, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14801, 
      n14802, n14803, n14805, n14806, n14809, n14810, n14811, n14812, n14813, 
      n14814, n14815, n14817, n14818, n14819, n14820, n14821, n14822, n14828, 
      n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, 
      n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, 
      n14847, n14848, n14849, n14851, n14853, n14854, n14855, n14856, n14858, 
      n14859, n14860, n14861, n14863, n14864, n14865, n14866, n14867, n14868, 
      n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14878, 
      n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, 
      n14890, n14891, n14892, n14893, n14895, n14896, n14897, n14898, n14899, 
      n14901, n14902, n14903, n14905, n14906, n14907, n14908, n14911, n14912, 
      n14913, n14914, n14915, n14916, n14917, n14918, n14920, n14922, n14924, 
      n14925, n14926, n14927, n14930, n14931, n14932, n14933, n14934, n14935, 
      n14937, n14938, n14939, n14940, n14942, n14943, n14944, n14945, n14948, 
      n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14957, n14959, 
      n14960, n14964, n14965, n14966, n14967, n14968, n14969, n14971, n14972, 
      n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14983, 
      n14985, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, 
      n14996, n14997, n14998, n14999, n15000, n15002, n15004, n15005, n15006, 
      n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15015, n15016, 
      n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, 
      n15026, n15027, n15028, n15029, n15031, n15032, n15033, n15035, n15036, 
      n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, 
      n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, 
      n15055, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, 
      n15065, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15077, 
      n15078, n15079, n15083, n15084, n15085, n15086, n15089, n15091, n15092, 
      n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15101, n15103, 
      n15106, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, 
      n15116, n15117, n15119, n15120, n15121, n15123, n15124, n15126, n15127, 
      n15129, n15130, n15132, n15133, n15134, n15135, n15136, n15137, n15139, 
      n15140, n15141, n15142, n15143, n15144, n15146, n15147, n15148, n15149, 
      n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, 
      n15160, n15161, n15162, n15165, n15166, n15167, n15168, n15169, n15171, 
      n15172, n15173, n15174, n15175, n15176, n15177, n15179, n15183, n15184, 
      n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, 
      n15194, n15195, n15196, n15198, n15204, n15205, n15206, n15207, n15208, 
      n15211, n15212, n15213, n15215, n15216, n15217, n15219, n15220, n15223, 
      n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, 
      n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, 
      n15243, n15245, n15246, n15247, n15249, n15250, n15253, n15254, n15255, 
      n15256, n15257, n15258, n15259, n15260, n15261, n15264, n15265, n15266, 
      n15267, n15268, n15270, n15271, n15272, n15274, n15275, n15276, n15277, 
      n15278, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, 
      n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, 
      n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, 
      n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, 
      n15319, n15321, n15322, n15323, n15324, n15326, n15327, n15328, n15329, 
      n15330, n15331, n15332, n15334, n15335, n15337, n15338, n15339, n15340, 
      n15341, n15343, n15344, n15346, n15347, n15348, n15349, n15350, n15351, 
      n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, 
      n15362, n15364, n15365, n15366, n15367, n15368, n15370, n15371, n15372, 
      n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15381, n15382, 
      n15383, n15384, n15385, n15386, n15389, n15390, n15391, n15393, n15394, 
      n15395, n15396, n15397, n15399, n15400, n15401, n15402, n15404, n15405, 
      n15406, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, 
      n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, 
      n15425, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, 
      n15435, n15436, n15437, n15438, n15441, n15442, n15443, n15444, n15446, 
      n15448, n15449, n15450, n15451, n15452, n15455, n15456, n15457, n15458, 
      n15459, n15460, n15462, n15464, n15465, n15466, n15467, n15468, n15470, 
      n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, 
      n15480, n15481, n15483, n15484, n15485, n15486, n15487, n15489, n15490, 
      n15494, n15495, n15496, n15497, n15498, n15500, n15501, n15502, n15505, 
      n15506, n15507, n15508, n15514, n15515, n15516, n15517, n15518, n15519, 
      n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, 
      n15529, n15530, n15531, n15534, n15536, n15537, n15538, n15539, n15540, 
      n15543, n15544, n15546, n15548, n15550, n15551, n15553, n15555, n15556, 
      n15557, n15559, n15560, n15561, n15562, n15564, n15565, n15566, n15569, 
      n15570, n15571, n15573, n15574, n15575, n15576, n15577, n15578, n15579, 
      n15580, n15581, n15583, n15584, n15585, n15588, n15589, n15590, n15591, 
      n15592, n15593, n15594, n15595, n15597, n15598, n15599, n15600, n15601, 
      n15602, n15606, n15607, n15608, n15609, n15611, n15612, n15613, n15614, 
      n15615, n15616, n15617, n15618, n15621, n15622, n15623, n15624, n15627, 
      n15628, n15629, n15630, n15631, n15632, n15633, n15635, n15636, n15638, 
      n15639, n15640, n15641, n15642, n15643, n15644, n15646, n15650, n15652, 
      n15653, n15655, n15658, n15659, n15660, n15661, n15662, n15663, n15665, 
      n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, 
      n15675, n15676, n15677, n15679, n15680, n15681, n15682, n15683, n15685, 
      n15686, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, 
      n15698, n15699, n15701, n15702, n15704, n15705, n15707, n15708, n15709, 
      n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, 
      n15719, n15720, n15721, n15722, n15725, n15726, n15727, n15728, n15729, 
      n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, 
      n15740, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, 
      n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15759, n15761, 
      n15763, n15765, n15768, n15769, n15770, n15771, n15772, n15774, n15775, 
      n15776, n15777, n15778, n15779, n15780, n15781, n15783, n15785, n15786, 
      n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15795, n15796, 
      n15797, n15798, n15799, n15801, n15802, n15803, n15804, n15805, n15806, 
      n15807, n15808, n15811, n15812, n15813, n15814, n15815, n15816, n15817, 
      n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15827, 
      n15828, n15829, n15830, n15831, n15832, n15833, n15835, n15836, n15837, 
      n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, 
      n15847, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15857, 
      n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15867, 
      n15869, n15870, n15872, n15873, n15874, n15875, n15876, n15877, n15880, 
      n15882, n15883, n15885, n15886, n15887, n15888, n15889, n15890, n15891, 
      n15893, n15894, n15896, n15897, n15898, n15899, n15900, n15902, n15904, 
      n15905, n15906, n15907, n15909, n15910, n15911, n15912, n15913, n15914, 
      n15915, n15917, n15919, n15920, n15923, n15925, n15927, n15928, n15929, 
      n15930, n15931, n15932, n15934, n15935, n15936, n15939, n15941, n15942, 
      n15943, n15944, n15946, n15947, n15948, n15949, n15950, n15951, n15953, 
      n15954, n15955, n15956, n15957, n15959, n15960, n15961, n15963, n15964, 
      n15965, n15966, n15967, n15968, n15969, n15971, n15973, n15974, n15976, 
      n15977, n15978, n15979, n15982, n15983, n15984, n15985, n15986, n15987, 
      n15988, n15990, n15991, n15992, n15993, n15994, n15996, n15997, n15998, 
      n15999, n16000, n16001, n16002, n16004, n16005, n16007, n16008, n16009, 
      n16010, n16011, n16012, n16013, n16014, n16016, n16017, n16018, n16021, 
      n16022, n16023, n16024, n16025, n16027, n16028, n16029, n16030, n16033, 
      n16034, n16035, n16036, n16038, n16039, n16041, n16042, n16045, n16046, 
      n16047, n16048, n16050, n16051, n16052, n16053, n16054, n16058, n16059, 
      n16060, n16062, n16065, n16066, n16068, n16070, n16072, n16073, n16076, 
      n16077, n16078, n16080, n16081, n16083, n16084, n16085, n16086, n16088, 
      n16090, n16091, n16092, n16093, n16094, n16096, n16097, n16098, n16099, 
      n16100, n16104, n16105, n16106, n16108, n16109, n16110, n16111, n16112, 
      n16113, n16115, n16117, n16118, n16120, n16121, n16122, n16123, n16124, 
      n16125, n16127, n16128, n16129, n16132, n16133, n16134, n16136, n16137, 
      n16138, n16139, n16140, n16141, n16142, n16144, n16146, n16147, n16148, 
      n16149, n16150, n16152, n16154, n16155, n16156, n16157, n16158, n16159, 
      n16160, n16162, n16163, n16164, n16165, n16166, n16167, n16169, n16170, 
      n16173, n16174, n16175, n16176, n16178, n16180, n16181, n16182, n16184, 
      n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, 
      n16194, n16195, n16196, n16197, n16198, n16200, n16202, n16203, n16204, 
      n16205, n16207, n16209, n16210, n16211, n16212, n16215, n16216, n16217, 
      n16218, n16220, n16221, n16222, n16224, n16225, n16226, n16228, n16229, 
      n16231, n16232, n16235, n16236, n16237, n16238, n16239, n16240, n16241, 
      n16242, n16243, n16246, n16247, n16248, n16249, n16251, n16253, n16254, 
      n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16265, n16266, 
      n16267, n16269, n16271, n16272, n16273, n16274, n16275, n16276, n16277, 
      n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16286, n16287, 
      n16288, n16290, n16291, n16292, n16293, n16295, n16297, n16298, n16300, 
      n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, 
      n16310, n16311, n16313, n16315, n16317, n16318, n16319, n16320, n16321, 
      n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16331, n16332, 
      n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16343, n16344, 
      n16345, n16346, n16347, n16348, n16349, n16351, n16352, n16353, n16354, 
      n16355, n16356, n16357, n16358, n16359, n16361, n16363, n16364, n16366, 
      n16367, n16370, n16371, n16372, n16373, n16374, n16375, n16377, n16378, 
      n16380, n16381, n16382, n16383, n16384, n16386, n16387, n16388, n16389, 
      n16390, n16392, n16393, n16394, n16395, n16397, n16398, n16400, n16401, 
      n16402, n16403, n16406, n16408, n16409, n16410, n16411, n16412, n16413, 
      n16414, n16416, n16417, n16418, n16420, n16421, n16422, n16423, n16424, 
      n16425, n16426, n16429, n16430, n16431, n16432, n16434, n16435, n16437, 
      n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16447, 
      n16448, n16450, n16451, n16452, n16453, n16454, n16457, n16458, n16459, 
      n16461, n16462, n16463, n16464, n16466, n16467, n16468, n16469, n16472, 
      n16473, n16474, n16477, n16479, n16481, n16482, n16483, n16484, n16485, 
      n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, 
      n16496, n16497, n16501, n16502, n16503, n16504, n16505, n16506, n16507, 
      n16509, n16510, n16512, n16513, n16514, n16515, n16516, n16518, n16519, 
      n16520, n16522, n16523, n16525, n16526, n16527, n16528, n16529, n16530, 
      n16531, n16532, n16533, n16534, n16535, n16536, n16538, n16539, n16540, 
      n16541, n16543, n16544, n16545, n16546, n16548, n16549, n16550, n16551, 
      n16552, n16553, n16554, n16555, n16556, n16558, n16559, n16560, n16561, 
      n16562, n16563, n16564, n16566, n16567, n16568, n16569, n16570, n16572, 
      n16573, n16574, n16575, n16577, n16578, n16579, n16581, n16582, n16583, 
      n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, 
      n16595, n16596, n16597, n16598, n16600, n16601, n16602, n16603, n16604, 
      n16605, n16606, n16607, n16608, n16609, n16611, n16612, n16613, n16614, 
      n16615, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, 
      n16625, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, 
      n16635, n16636, n16637, n16639, n16640, n16641, n16642, n16643, n16646, 
      n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, 
      n16657, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, 
      n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, 
      n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, 
      n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, 
      n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16703, n16704, 
      n16705, n16708, n16710, n16711, n16712, n16713, n16716, n16717, n16718, 
      n16719, n16722, n16723, n16724, n16725, n16727, n16728, n16729, n16730, 
      n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, 
      n16741, n16743, n16745, n16747, n16748, n16749, n16750, n16751, n16752, 
      n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16762, n16763, 
      n16766, n16767, n16768, n16769, n16770, n16773, n16774, n16775, n16776, 
      n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, 
      n16786, n16787, n16788, n16789, n16790, n16792, n16793, n16795, n16796, 
      n16797, n16798, n16799, n16800, n16801, n16803, n16804, n16805, n16806, 
      n16807, n16809, n16810, n16811, n16812, n16815, n16816, n16817, n16818, 
      n16819, n16820, n16823, n16824, n16826, n16827, n16828, n16829, n16831, 
      n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16841, n16842, 
      n16844, n16845, n16847, n16848, n16849, n16850, n16851, n16852, n16853, 
      n16854, n16855, n16857, n16858, n16859, n16861, n16862, n16863, n16864, 
      n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, 
      n16875, n16876, n16877, n16879, n16881, n16882, n16883, n16884, n16885, 
      n16886, n16887, n16888, n16889, n16891, n16893, n16896, n16897, n16898, 
      n16899, n16901, n16904, n16905, n16906, n16907, n16908, n16909, n16910, 
      n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, 
      n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, 
      n16930, n16933, n16934, n16937, n16938, n16939, n16940, n16943, n16945, 
      n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, 
      n16955, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, 
      n16966, n16969, n16971, n16972, n16973, n16974, n16975, n16976, n16977, 
      n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, 
      n16987, n16989, n16992, n16993, n16995, n16996, n16997, n16998, n17001, 
      n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, 
      n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, 
      n17021, n17022, n17023, n17026, n17028, n17029, n17030, n17035, n17036, 
      n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17046, 
      n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, 
      n17056, n17058, n17060, n17061, n17062, n17063, n17064, n17065, n17066, 
      n17067, n17068, n17069, n17072, n17073, n17074, n17076, n17077, n17078, 
      n17079, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, 
      n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, 
      n17100, n17101, n17102, n17104, n17105, n17106, n17108, n17109, n17110, 
      n17112, n17113, n17114, n17115, n17117, n17118, n17119, n17120, n17122, 
      n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, 
      n17132, n17133, n17134, n17135, n17136, n17139, n17140, n17141, n17143, 
      n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17153, 
      n17155, n17156, n17157, n17159, n17161, n17162, n17163, n17164, n17165, 
      n17166, n17167, n17168, n17169, n17171, n17172, n17174, n17175, n17177, 
      n17178, n17180, n17181, n17183, n17184, n17185, n17186, n17187, n17188, 
      n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17199, 
      n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17211, 
      n17212, n17213, n17214, n17215, n17217, n17218, n17219, n17220, n17222, 
      n17223, n17224, n17225, n17226, n17227, n17228, n17231, n17232, n17233, 
      n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, 
      n17243, n17244, n17245, n17247, n17248, n17249, n17251, n17253, n17254, 
      n17255, n17257, n17258, n17259, n17260, n17261, n17263, n17266, n17268, 
      n17269, n17270, n17271, n17272, n17273, n17274, n17277, n17278, n17280, 
      n17281, n17282, n17284, n17285, n17286, n17287, n17288, n17289, n17290, 
      n17291, n17293, n17295, n17296, n17297, n17298, n17299, n17300, n17301, 
      n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, 
      n17311, n17313, n17316, n17317, n17318, n17319, n17320, n17321, n17322, 
      n17323, n17324, n17325, n17327, n17328, n17329, n17330, n17331, n17333, 
      n17334, n17335, n17336, n17338, n17339, n17341, n17342, n17346, n17347, 
      n17348, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, 
      n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17367, n17368, 
      n17369, n17370, n17371, n17373, n17374, n17375, n17377, n17378, n17379, 
      n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17389, 
      n17392, n17393, n17394, n17395, n17396, n17398, n17399, n17400, n17401, 
      n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17411, 
      n17414, n17415, n17416, n17418, n17419, n17420, n17422, n17423, n17424, 
      n17425, n17426, n17428, n17429, n17430, n17431, n17432, n17434, n17435, 
      n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, 
      n17445, n17446, n17448, n17450, n17452, n17453, n17455, n17456, n17457, 
      n17458, n17460, n17462, n17463, n17464, n17465, n17466, n17467, n17472, 
      n17473, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, 
      n17483, n17485, n17486, n17487, n17488, n17489, n17490, n17492, n17493, 
      n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, 
      n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, 
      n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, 
      n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17531, 
      n17532, n17535, n17537, n17538, n17540, n17541, n17542, n17543, n17544, 
      n17546, n17547, n17548, n17549, n17551, n17552, n17553, n17554, n17555, 
      n17556, n17557, n17558, n17559, n17561, n17562, n17563, n17564, n17565, 
      n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, 
      n17575, n17576, n17578, n17579, n17580, n17581, n17582, n17584, n17585, 
      n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, 
      n17595, n17597, n17598, n17599, n17600, n17601, n17602, n17604, n17605, 
      n17606, n17608, n17609, n17612, n17613, n17616, n17617, n17618, n17621, 
      n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17630, n17631, 
      n17633, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, 
      n17643, n17644, n17647, n17649, n17650, n17651, n17652, n17653, n17655, 
      n17658, n17659, n17661, n17662, n17663, n17664, n17665, n17666, n17668, 
      n17669, n17670, n17672, n17673, n17675, n17676, n17677, n17678, n17679, 
      n17680, n17681, n17682, n17683, n17684, n17685, n17687, n17688, n17689, 
      n17691, n17692, n17693, n17694, n17696, n17697, n17698, n17699, n17701, 
      n17703, n17704, n17705, n17707, n17708, n17709, n17711, n17712, n17713, 
      n17714, n17715, n17716, n17717, n17718, n17720, n17721, n17722, n17723, 
      n17725, n17726, n17728, n17729, n17730, n17731, n17732, n17734, n17735, 
      n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, 
      n17745, n17746, n17747, n17748, n17750, n17752, n17753, n17754, n17755, 
      n17756, n17758, n17759, n17760, n17762, n17764, n17765, n17766, n17767, 
      n17768, n17770, n17771, n17773, n17774, n17775, n17777, n17778, n17779, 
      n17781, n17782, n17784, n17785, n17786, n17787, n17790, n17791, n17792, 
      n17793, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, 
      n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, 
      n17814, n17815, n17816, n17817, n17819, n17820, n17821, n17822, n17824, 
      n17826, n17828, n17829, n17830, n17832, n17833, n17834, n17835, n17837, 
      n17838, n17839, n17840, n17841, n17843, n17844, n17845, n17849, n17850, 
      n17853, n17855, n17857, n17858, n17859, n17860, n17861, n17863, n17865, 
      n17866, n17867, n17869, n17871, n17872, n17873, n17874, n17875, n17876, 
      n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17886, 
      n17887, n17888, n17889, n17890, n17891, n17893, n17894, n17895, n17896, 
      n17897, n17898, n17899, n17900, n17903, n17904, n17905, n17906, n17907, 
      n17910, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, 
      n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, 
      n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, 
      n17940, n17941, n17943, n17944, n17945, n17947, n17948, n17949, n17950, 
      n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17963, 
      n17964, n17967, n17968, n17970, n17971, n17973, n17974, n17975, n17977, 
      n17978, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, 
      n17991, n17992, n17993, n17995, n17996, n17997, n17998, n17999, n18001, 
      n18002, n18003, n18005, n18006, n18007, n18010, n18011, n18012, n18013, 
      n18015, n18017, n18018, n18019, n18020, n18021, n18022, n18024, n18025, 
      n18026, n18028, n18029, n18031, n18032, n18033, n18034, n18035, n18036, 
      n18037, n18038, n18039, n18041, n18042, n18043, n18044, n18047, n18048, 
      n18049, n18050, n18051, n18054, n18055, n18056, n18058, n18059, n18062, 
      n18064, n18065, n18068, n18071, n18072, n18073, n18074, n18075, n18076, 
      n18077, n18078, n18079, n18080, n18082, n18083, n18084, n18085, n18088, 
      n18089, n18090, n18091, n18094, n18095, n18096, n18098, n18099, n18100, 
      n18101, n18102, n18103, n18105, n18106, n18107, n18108, n18109, n18110, 
      n18112, n18113, n18114, n18117, n18118, n18119, n18120, n18121, n18122, 
      n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, 
      n18132, n18133, n18135, n18136, n18137, n18138, n18139, n18141, n18142, 
      n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, 
      n18152, n18154, n18155, n18156, n18159, n18160, n18161, n18162, n18163, 
      n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, 
      n18174, n18175, n18177, n18179, n18180, n18181, n18182, n18184, n18185, 
      n18186, n18187, n18188, n18189, n18190, n18192, n18194, n18195, n18196, 
      n18197, n18198, n18199, n18200, n18204, n18205, n18206, n18207, n18208, 
      n18209, n18210, n18213, n18215, n18216, n18217, n18218, n18219, n18220, 
      n18221, n18224, n18225, n18226, n18227, n18228, n18230, n18231, n18235, 
      n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18246, n18251, 
      n18254, n18256, n18257, n18259, n18260, n18261, n18264, n18265, n18266, 
      n18267, n18268, n18269, n18270, n18274, n18275, n18276, n18277, n18278, 
      n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, 
      n18288, n18289, n18290, n18292, n18293, n18294, n18295, n18297, n18298, 
      n18299, n18300, n18301, n18302, n18303, n18304, n18307, n18308, n18309, 
      n18310, n18311, n18313, n18314, n18315, n18316, n18317, n18318, n18320, 
      n18321, n18322, n18323, n18324, n18326, n18327, n18328, n18329, n18330, 
      n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, 
      n18340, n18341, n18344, n18345, n18346, n18347, n18348, n18349, n18350, 
      n18352, n18354, n18356, n18357, n18359, n18360, n18361, n18362, n18363, 
      n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, 
      n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18381, n18382, 
      n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, 
      n18392, n18393, n18395, n18396, n18397, n18398, n18399, n18400, n18401, 
      n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, 
      n18411, n18412, n18413, n18415, n18416, n18417, n18418, n18419, n18420, 
      n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, 
      n18431, n18432, n18433, n18434, n18435, n18437, n18438, n18439, n18440, 
      n18441, n18443, n18444, n18445, n18446, n18447, n18449, n18450, n18452, 
      n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18462, 
      n18463, n18464, n18467, n18468, n18469, n18470, n18471, n18472, n18473, 
      n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, 
      n18483, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, 
      n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, 
      n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, 
      n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, 
      n18520, n18521, n18522, n18524, n18525, n18526, n18527, n18528, n18530, 
      n18531, n18532, n18534, n18535, n18536, n18537, n18538, n18539, n18540, 
      n18541, n18543, n18546, n18548, n18549, n18550, n18551, n18553, n18554, 
      n18555, n18556, n18557, n18559, n18560, n18561, n18563, n18565, n18566, 
      n18567, n18569, n18571, n18572, n18573, n18574, n18575, n18576, n18577, 
      n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, 
      n18587, n18588, n18590, n18591, n18593, n18594, n18595, n18596, n18598, 
      n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, 
      n18608, n18609, n18613, n18615, n18616, n18617, n18618, n18619, n18621, 
      n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18631, 
      n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, 
      n18641, n18642, n18643, n18647, n18648, n18649, n18650, n18651, n18653, 
      n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18662, n18663, 
      n18664, n18665, n18666, n18667, n18668, n18669, n18671, n18672, n18674, 
      n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18686, 
      n18687, n18688, n18691, n18692, n18693, n18694, n18695, n18696, n18697, 
      n18698, n18699, n18700, n18701, n18702, n18704, n18705, n18706, n18707, 
      n18708, n18709, n18710, n18711, n18714, n18715, n18716, n18717, n18718, 
      n18719, n18720, n18721, n18722, n18723, n18724, n18726, n18727, n18729, 
      n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, 
      n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, 
      n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, 
      n18757, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, 
      n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, 
      n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18784, n18785, 
      n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, 
      n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, 
      n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, 
      n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, 
      n18822, n18823, n18824, n18825, n18827, n18828, n18829, n18830, n18831, 
      n18832, n18833, n18835, n18836, n18838, n18839, n18840, n18841, n18842, 
      n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, 
      n18853, n18854, n18855, n18856, n18858, n18859, n18860, n18861, n18862, 
      n18863, n18864, n18865, n18866, n18867, n18869, n18870, n18871, n18873, 
      n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, 
      n18884, n18885, n18886, n18887, n18888, n18889, n18891, n18892, n18893, 
      n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, 
      n18903, n18904, n18905, n18907, n18908, n18909, n18910, n18911, n18912, 
      n18913, n18914, n18915, n18916, n18917, n18919, n18920, n18921, n18922, 
      n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, 
      n18932, n18935, n18937, n18938, n18939, n18940, n18941, n18942, n18943, 
      n18944, n18945, n18946, n18947, n18948, n18949, n18952, n18953, n18955, 
      n18956, n18957, n18958, n18959, n18960, n18962, n18963, n18964, n18965, 
      n18966, n18967, n18969, n18970, n18971, n18973, n18974, n18975, n18976, 
      n18977, n18978, n18979, n18980, n18982, n18983, n18984, n18985, n18986, 
      n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, 
      n18996, n18997, n18999, n19000, n19002, n19003, n19004, n19006, n19007, 
      n19008, n19009, n19010, n19011, n19013, n19014, n19016, n19017, n19020, 
      n19021, n19022, n19023, n19024, n19026, n19027, n19028, n19029, n19030, 
      n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, 
      n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, 
      n19049, n19050, n19051, n19052, n19053, n19056, n19057, n19058, n19059, 
      n19060, n19061, n19062, n19063, n19064, n19065, n19067, n19068, n19069, 
      n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, 
      n19079, n19080, n19084, n19085, n19087, n19088, n19089, n19090, n19091, 
      n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19100, n19101, 
      n19102, n19103, n19104, n19105, n19107, n19108, n19109, n19110, n19111, 
      n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, 
      n19121, n19122, n19123, n19124, n19125, n19126, n19128, n19130, n19131, 
      n19132, n19133, n19134, n19135, n19136, n19137, n19139, n19140, n19141, 
      n19142, n19143, n19144, n19146, n19147, n19148, n19149, n19150, n19151, 
      n19152, n19153, n19154, n19155, n19156, n19158, n19160, n19161, n19162, 
      n19163, n19164, n19165, n19167, n19168, n19170, n19171, n19172, n19173, 
      n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, 
      n19183, n19185, n19186, n19188, n19189, n19190, n19193, n19195, n19196, 
      n19197, n19198, n19199, n19200, n19202, n19203, n19204, n19205, n19206, 
      n19209, n19210, n19211, n19212, n19214, n19215, n19216, n19217, n19218, 
      n19219, n19220, n19222, n19224, n19225, n19226, n19227, n19228, n19229, 
      n19230, n19232, n19233, n19234, n19235, n19236, n19238, n19239, n19240, 
      n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, 
      n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, 
      n19259, n19260, n19261, n19262, n19263, n19265, n19267, n19268, n19269, 
      n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, 
      n19280, n19281, n19282, n19283, n19284, n19285, n19287, n19288, n19289, 
      n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, 
      n19300, n19301, n19302, n19303, n19305, n19307, n19308, n19309, n19310, 
      n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, 
      n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19328, n19329, 
      n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, 
      n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, 
      n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, 
      n19357, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, 
      n19367, n19368, n19370, n19371, n19372, n19373, n19374, n19375, n19376, 
      n19377, n19378, n19379, n19380, n19381, n19382, n19384, n19385, n19386, 
      n19387, n19388, n19389, n19390, n19391, n19394, n19395, n19397, n19398, 
      n19399, n19400, n19401, n19402, n19403, n19405, n19406, n19407, n19408, 
      n19409, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, 
      n19419, n19420, n19421, n19422, n19423, n19424, n19426, n19427, n19428, 
      n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19438, 
      n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, 
      n19448, n19449, n19450, n19451, n19453, n19454, n19455, n19456, n19457, 
      n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, 
      n19468, n19469, n19470, n19471, n19473, n19474, n19475, n19476, n19479, 
      n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19490, 
      n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19500, 
      n19501, n19502, n19503, n19504, n19505, n19507, n19508, n19509, n19510, 
      n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, 
      n19520, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, 
      n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, 
      n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, 
      n19549, n19550, n19551, n19552, n19554, n19555, n19556, n19557, n19558, 
      n19559, n19561, n19562, n19564, n19565, n19566, n19567, n19568, n19570, 
      n19571, n19573, n19574, n19575, n19577, n19578, n19579, n19580, n19582, 
      n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, 
      n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19601, 
      n19602, n19603, n19604, n19605, n19606, n19607, n19609, n19610, n19611, 
      n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, 
      n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, 
      n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, 
      n19639, n19640, n19641, n19642, n19644, n19647, n19648, n19649, n19651, 
      n19653, n19654, n19655, n19657, n19658, n19659, n19660, n19661, n19662, 
      n19663, n19664, n19666, n19667, n19668, n19669, n19671, n19672, n19673, 
      n19675, n19676, n19677, n19679, n19680, n19681, n19682, n19683, n19684, 
      n19685, n19686, n19687, n19689, n19690, n19691, n19693, n19694, n19695, 
      n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19705, 
      n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19716, 
      n19717, n19718, n19719, n19721, n19722, n19723, n19724, n19726, n19727, 
      n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, 
      n19737, n19739, n19740, n19741, n19742, n19743, n19744, n19746, n19748, 
      n19749, n19750, n19751, n19752, n19754, n19755, n19757, n19759, n19761, 
      n19763, n19764, n19766, n19767, n19768, n19769, n19770, n19771, n19772, 
      n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19782, 
      n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, 
      n19792, n19794, n19796, n19798, n19799, n19800, n19801, n19803, n19804, 
      n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19814, 
      n19816, n19817, n19818, n19819, n19820, n19822, n19823, n19824, n19825, 
      n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, 
      n19835, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, 
      n19845, n19846, n19847, n19849, n19850, n19851, n19853, n19854, n19855, 
      n19856, n19857, n19861, n19862, n19863, n19864, n19865, n19866, n19867, 
      n19868, n19869, n19871, n19872, n19874, n19875, n19876, n19878, n19879, 
      n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19888, n19889, 
      n19891, n19892, n19893, n19894, n19896, n19897, n19898, n19899, n19900, 
      n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, 
      n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, 
      n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, 
      n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19938, 
      n19939, n19940, n19941, n19942, n19943, n19944, n19947, n19948, n19949, 
      n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, 
      n19959, n19960, n19961, n19962, n19964, n19965, n19966, n19967, n19968, 
      n19969, n19970, n19971, n19972, n19974, n19975, n19976, n19977, n19979, 
      n19984, n19986, n19987, n19990, n19991, n19992, n19993, n19994, n19995, 
      n19996, n19997, n19998, n20000, n20001, n20002, n20003, n20004, n20005, 
      n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, 
      n20015, n20017, n20018, n20019, n20020, n20021, n20022, n20024, n20025, 
      n20026, n20028, n20029, n20032, n20033, n20034, n20035, n20036, n20037, 
      n20038, n20039, n20040, n20042, n20043, n20044, n20045, n20047, n20048, 
      n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, 
      n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, 
      n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20075, n20076, 
      n20077, n20078, n20079, n20080, n20081, n20083, n20084, n20085, n20086, 
      n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, 
      n20096, n20097, n20098, n20099, n20100, n20102, n20103, n20104, n20105, 
      n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20116, 
      n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, 
      n20126, n20127, n20128, n20130, n20132, n20133, n20134, n20135, n20136, 
      n20137, n20138, n20139, n20141, n20142, n20143, n20144, n20147, n20148, 
      n20149, n20150, n20152, n20153, n20154, n20155, n20156, n20157, n20158, 
      n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, 
      n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, 
      n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20186, n20187, 
      n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20196, n20197, 
      n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, 
      n20208, n20209, n20210, n20213, n20216, n20217, n20218, n20219, n20220, 
      n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, 
      n20230, n20231, n20233, n20234, n20235, n20236, n20237, n20238, n20239, 
      n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, 
      n20249, n20251, n20252, n20254, n20255, n20256, n20257, n20258, n20259, 
      n20261, n20263, n20266, n20267, n20268, n20269, n20270, n20271, n20272, 
      n20273, n20274, n20275, n20276, n20277, n20278, n20280, n20281, n20282, 
      n20283, n20284, n20285, n20287, n20288, n20289, n20290, n20291, n20292, 
      n20293, n20294, n20296, n20297, n20298, n20299, n20300, n20301, n20302, 
      n20304, n20305, n20306, n20308, n20309, n20310, n20311, n20312, n20313, 
      n20314, n20315, n20316, n20317, n20318, n20319, n20321, n20322, n20323, 
      n20324, n20325, n20327, n20328, n20329, n20330, n20332, n20333, n20334, 
      n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20344, 
      n20345, n20347, n20349, n20350, n20351, n20352, n20353, n20354, n20356, 
      n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20366, 
      n20367, n20368, n20371, n20373, n20374, n20375, n20376, n20377, n20378, 
      n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, 
      n20389, n20390, n20392, n20393, n20395, n20396, n20397, n20399, n20400, 
      n20401, n20403, n20404, n20405, n20406, n20407, n20408, n20410, n20411, 
      n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, 
      n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, 
      n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, 
      n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, 
      n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, 
      n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20466, n20467, 
      n20468, n20471, n20472, n20475, n20476, n20479, n20480, n20481, n20482, 
      n20483, n20484, n20485, n20486, n20487, n20489, n20490, n20492, n20493, 
      n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, 
      n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, 
      n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, 
      n20521, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20531, 
      n20533, n20534, n20535, n20536, n20537, n20538, n20540, n20541, n20542, 
      n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, 
      n20554, n20555, n20556, n20557, n20558, n20560, n20561, n20562, n20563, 
      n20564, n20565, n20566, n20568, n20569, n20570, n20571, n20572, n20573, 
      n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, 
      n20583, n20584, n20585, n20586, n20588, n20589, n20590, n20591, n20592, 
      n20593, n20594, n20595, n20598, n20599, n20600, n20601, n20602, n20603, 
      n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20612, n20613, 
      n20614, n20615, n20616, n20617, n20619, n20620, n20621, n20622, n20623, 
      n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, 
      n20633, n20634, n20635, n20636, n20639, n20640, n20641, n20642, n20644, 
      n20645, n20647, n20648, n20649, n20650, n20651, n20652, n20654, n20657, 
      n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20667, n20668, 
      n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, 
      n20678, n20679, n20680, n20682, n20684, n20686, n20687, n20688, n20690, 
      n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, 
      n20700, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, 
      n20710, n20711, n20712, n20713, n20715, n20716, n20717, n20718, n20719, 
      n20720, n20721, n20722, n20723, n20724, n20726, n20727, n20729, n20730, 
      n20731, n20732, n20733, n20736, n20737, n20738, n20739, n20740, n20742, 
      n20743, n20744, n20746, n20747, n20748, n20749, n20751, n20752, n20753, 
      n20754, n20755, n20756, n20757, n20758, n20759, n20762, n20764, n20765, 
      n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, 
      n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, 
      n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, 
      n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20801, n20802, 
      n20803, n20804, n20806, n20807, n20808, n20809, n20810, n20813, n20815, 
      n20816, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, 
      n20827, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, 
      n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20848, n20849, 
      n20850, n20851, n20852, n20853, n20855, n20856, n20857, n20858, n20859, 
      n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, 
      n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20877, n20879, 
      n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, 
      n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, 
      n20899, n20900, n20902, n20904, n20905, n20906, n20907, n20908, n20909, 
      n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, 
      n20919, n20920, n20921, n20922, n20924, n20925, n20926, n20927, n20928, 
      n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20938, 
      n20939, n20940, n20941, n20944, n20945, n20946, n20947, n20949, n20950, 
      n20951, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, 
      n20961, n20962, n20963, n20964, n20966, n20967, n20968, n20970, n20971, 
      n20972, n20974, n20975, n20976, n20977, n20978, n20979, n20982, n20983, 
      n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20992, n20993, 
      n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, 
      n21003, n21004, n21005, n21006, n21007, n21009, n21010, n21011, n21012, 
      n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21022, n21023, 
      n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, 
      n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, 
      n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, 
      n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, 
      n21060, n21061, n21064, n21065, n21066, n21067, n21068, n21069, n21070, 
      n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, 
      n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, 
      n21089, n21090, n21091, n21093, n21095, n21096, n21097, n21098, n21099, 
      n21100, n21101, n21104, n21107, n21109, n21110, n21112, n21113, n21114, 
      n21115, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21125, 
      n21126, n21127, n21129, n21131, n21132, n21134, n21136, n21137, n21138, 
      n21139, n21140, n21141, n21143, n21145, n21146, n21147, n21148, n21149, 
      n21151, n21152, n21153, n21154, n21155, n21156, n21158, n21159, n21160, 
      n21161, n21162, n21163, n21164, n21165, n21167, n21168, n21169, n21170, 
      n21171, n21172, n21173, n21175, n21176, n21178, n21179, n21180, n21181, 
      n21182, n21183, n21184, n21187, n21188, n21189, n21190, n21191, n21192, 
      n21193, n21195, n21196, n21198, n21199, n21200, n21202, n21203, n21204, 
      n21206, n21207, n21209, n21210, n21211, n21212, n21213, n21214, n21215, 
      n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, 
      n21225, n21226, n21228, n21230, n21232, n21233, n21234, n21235, n21237, 
      n21239, n21240, n21241, n21243, n21244, n21247, n21248, n21249, n21251, 
      n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, 
      n21261, n21263, n21264, n21265, n21266, n21267, n21269, n21270, n21272, 
      n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, 
      n21282, n21283, n21284, n21285, n21286, n21289, n21291, n21292, n21295, 
      n21297, n21298, n21299, n21300, n21302, n21303, n21304, n21305, n21306, 
      n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, 
      n21316, n21317, n21320, n21321, n21322, n21323, n21324, n21325, n21326, 
      n21328, n21330, n21331, n21332, n21334, n21335, n21336, n21337, n21338, 
      n21339, n21340, n21341, n21343, n21345, n21346, n21347, n21348, n21349, 
      n21350, n21351, n21353, n21354, n21356, n21357, n21358, n21359, n21361, 
      n21362, n21363, n21365, n21366, n21367, n21368, n21369, n21370, n21372, 
      n21373, n21374, n21375, n21377, n21378, n21379, n21381, n21382, n21383, 
      n21385, n21386, n21387, n21389, n21390, n21391, n21392, n21393, n21394, 
      n21395, n21396, n21398, n21399, n21400, n21401, n21402, n21403, n21404, 
      n21405, n21406, n21407, n21408, n21410, n21411, n21412, n21413, n21414, 
      n21415, n21416, n21418, n21419, n21420, n21421, n21423, n21424, n21426, 
      n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21437, 
      n21438, n21439, n21440, n21441, n21442, n21443, n21445, n21447, n21448, 
      n21449, n21451, n21452, n21453, n21454, n21455, n21457, n21458, n21459, 
      n21460, n21461, n21462, n21463, n21465, n21466, n21467, n21468, n21469, 
      n21470, n21471, n21472, n21473, n21475, n21477, n21478, n21479, n21480, 
      n21481, n21482, n21483, n21484, n21485, n21487, n21488, n21489, n21490, 
      n21491, n21492, n21494, n21495, n21496, n21497, n21498, n21499, n21500, 
      n21501, n21502, n21503, n21504, n21505, n21506, n21509, n21510, n21512, 
      n21514, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, 
      n21525, n21527, n21529, n21530, n21531, n21532, n21534, n21535, n21536, 
      n21537, n21538, n21539, n21540, n21542, n21544, n21545, n21546, n21548, 
      n21549, n21550, n21551, n21553, n21554, n21555, n21556, n21558, n21559, 
      n21560, n21561, n21562, n21564, n21566, n21568, n21569, n21570, n21571, 
      n21572, n21573, n21574, n21576, n21577, n21579, n21580, n21581, n21582, 
      n21583, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, 
      n21594, n21595, n21596, n21597, n21599, n21600, n21601, n21602, n21603, 
      n21604, n21606, n21607, n21608, n21609, n21610, n21612, n21613, n21614, 
      n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, 
      n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21632, n21633, 
      n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, 
      n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, 
      n21652, n21653, n21655, n21656, n21657, n21658, n21659, n21660, n21661, 
      n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21671, 
      n21672, n21673, n21674, n21676, n21678, n21680, n21681, n21682, n21683, 
      n21684, n21685, n21686, n21687, n21688, n21690, n21691, n21692, n21693, 
      n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21704, n21705, 
      n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21715, 
      n21716, n21717, n21719, n21720, n21721, n21722, n21723, n21724, n21725, 
      n21726, n21727, n21728, n21730, n21731, n21732, n21733, n21736, n21737, 
      n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21746, n21747, 
      n21748, n21749, n21750, n21752, n21753, n21754, n21755, n21756, n21757, 
      n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, 
      n21768, n21769, n21771, n21772, n21775, n21776, n21777, n21778, n21779, 
      n21780, n21781, n21785, n21786, n21789, n21790, n21791, n21792, n21793, 
      n21794, n21795, n21796, n21797, n21799, n21800, n21801, n21804, n21805, 
      n21806, n21808, n21809, n21811, n21812, n21813, n21814, n21815, n21816, 
      n21817, n21818, n21819, n21820, n21821, n21823, n21824, n21825, n21826, 
      n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, 
      n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, 
      n21846, n21847, n21848, n21849, n21850, n21852, n21853, n21854, n21855, 
      n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, 
      n21865, n21866, n21867, n21869, n21870, n21871, n21872, n21873, n21874, 
      n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, 
      n21884, n21885, n21886, n21887, n21888, n21889, n21891, n21892, n21893, 
      n21894, n21896, n21898, n21899, n21900, n21901, n21902, n21903, n21905, 
      n21906, n21907, n21909, n21910, n21911, n21912, n21913, n21915, n21916, 
      n21918, n21919, n21920, n21921, n21923, n21924, n21925, n21926, n21927, 
      n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, 
      n21938, n21939, n21940, n21941, n21944, n21945, n21946, n21947, n21948, 
      n21949, n21950, n21951, n21952, n21953, n21956, n21957, n21958, n21959, 
      n21960, n21961, n21962, n21963, n21964, n21965, n21967, n21968, n21970, 
      n21971, n21972, n21974, n21975, n21979, n21980, n21981, n21983, n21984, 
      n21985, n21986, n21988, n21990, n21992, n21993, n21994, n21995, n21996, 
      n21997, n21998, n21999, n22000, n22002, n22003, n22004, n22005, n22006, 
      n22008, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, 
      n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, 
      n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, 
      n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, 
      n22046, n22047, n22048, n22049, n22051, n22053, n22054, n22055, n22056, 
      n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22066, 
      n22067, n22070, n22071, n22072, n22075, n22076, n22078, n22079, n22080, 
      n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, 
      n22090, n22091, n22092, n22093, n22094, n22096, n22098, n22099, n22100, 
      n22102, n22103, n22104, n22105, n22107, n22108, n22109, n22110, n22111, 
      n22112, n22113, n22114, n22115, n22118, n22119, n22120, n22121, n22123, 
      n22125, n22126, n22127, n22128, n22130, n22131, n22132, n22133, n22134, 
      n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, 
      n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, 
      n22154, n22155, n22156, n22157, n22158, n22160, n22161, n22162, n22163, 
      n22164, n22165, n22166, n22167, n22168, n22169, n22171, n22172, n22173, 
      n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, 
      n22183, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, 
      n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, 
      n22202, n22203, n22205, n22206, n22208, n22210, n22211, n22213, n22214, 
      n22216, n22217, n22218, n22220, n22221, n22222, n22223, n22224, n22225, 
      n22226, n22227, n22229, n22230, n22231, n22232, n22233, n22235, n22237, 
      n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22246, n22247, 
      n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, 
      n22258, n22259, n22260, n22261, n22264, n22265, n22266, n22267, n22268, 
      n22269, n22271, n22273, n22274, n22275, n22276, n22277, n22280, n22282, 
      n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22291, n22292, 
      n22293, n22294, n22295, n22296, n22297, n22299, n22300, n22301, n22302, 
      n22303, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, 
      n22313, n22314, n22315, n22317, n22318, n22319, n22320, n22322, n22324, 
      n22325, n22326, n22327, n22328, n22329, n22330, n22332, n22333, n22335, 
      n22336, n22337, n22338, n22339, n22340, n22342, n22343, n22344, n22348, 
      n22350, n22351, n22353, n22356, n22357, n22358, n22359, n22360, n22361, 
      n22362, n22363, n22364, n22366, n22367, n22368, n22369, n22372, n22375, 
      n22377, n22379, n22380, n22382, n22383, n22384, n22385, n22386, n22387, 
      n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22396, n22397, 
      n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22406, n22407, 
      n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, 
      n22418, n22420, n22421, n22422, n22424, n22425, n22426, n22427, n22428, 
      n22429, n22430, n22431, n22433, n22434, n22435, n22436, n22437, n22438, 
      n22439, n22441, n22442, n22443, n22444, n22446, n22448, n22449, n22450, 
      n22452, n22454, n22455, n22457, n22458, n22459, n22460, n22461, n22462, 
      n22463, n22464, n22466, n22467, n22468, n22470, n22471, n22472, n22473, 
      n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22482, n22483, 
      n22484, n22486, n22487, n22488, n22489, n22490, n22491, n22495, n22496, 
      n22497, n22498, n22499, n22500, n22502, n22503, n22504, n22505, n22508, 
      n22509, n22510, n22511, n22512, n22513, n22515, n22516, n22517, n22518, 
      n22521, n22522, n22523, n22524, n22526, n22527, n22529, n22530, n22531, 
      n22534, n22535, n22536, n22537, n22539, n22540, n22542, n22543, n22544, 
      n22546, n22547, n22549, n22550, n22551, n22552, n22553, n22555, n22556, 
      n22557, n22558, n22560, n22561, n22562, n22563, n22564, n22565, n22566, 
      n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, 
      n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, 
      n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22594, 
      n22595, n22596, n22597, n22598, n22599, n22600, n22602, n22603, n22604, 
      n22605, n22606, n22607, n22608, n22610, n22612, n22613, n22614, n22615, 
      n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, 
      n22625, n22626, n22627, n22628, n22629, n22631, n22633, n22634, n22635, 
      n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, 
      n22645, n22646, n22647, n22648, n22650, n22651, n22652, n22653, n22654, 
      n22655, n22656, n22657, n22658, n22659, n22660, n22662, n22663, n22664, 
      n22665, n22666, n22667, n22669, n22670, n22671, n22672, n22673, n22674, 
      n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22685, n22686, 
      n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22697, n22698, 
      n22699, n22701, n22704, n22705, n22706, n22707, n22709, n22710, n22711, 
      n22712, n22714, n22715, n22716, n22717, n22719, n22720, n22721, n22722, 
      n22723, n22724, n22725, n22726, n22728, n22729, n22730, n22731, n22732, 
      n22737, n22738, n22739, n22740, n22741, n22743, n22744, n22745, n22747, 
      n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, 
      n22757, n22758, n22759, n22760, n22761, n22762, n22765, n22766, n22767, 
      n22768, n22769, n22770, n22772, n22773, n22774, n22775, n22776, n22777, 
      n22778, n22779, n22780, n22781, n22783, n22784, n22785, n22786, n22789, 
      n22790, n22791, n22792, n22795, n22798, n22799, n22800, n22801, n22803, 
      n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22813, 
      n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22822, n22823, 
      n22824, n22825, n22826, n22827, n22828, n22830, n22831, n22832, n22833, 
      n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, 
      n22843, n22845, n22848, n22849, n22851, n22852, n22853, n22855, n22856, 
      n22857, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, 
      n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, 
      n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, 
      n22885, n22886, n22888, n22889, n22890, n22892, n22893, n22894, n22895, 
      n22896, n22897, n22899, n22900, n22901, n22904, n22905, n22906, n22907, 
      n22908, n22909, n22910, n22913, n22914, n22915, n22916, n22919, n22920, 
      n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, 
      n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22940, 
      n22942, n22943, n22944, n22945, n22946, n22948, n22949, n22950, n22951, 
      n22952, n22953, n22954, n22955, n22956, n22957, n22959, n22960, n22961, 
      n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, 
      n22971, n22972, n22973, n22974, n22977, n22978, n22979, n22981, n22982, 
      n22983, n22984, n22985, n22986, n22988, n22990, n22992, n22993, n22996, 
      n22997, n22999, n23000, n23002, n23003, n23004, n23005, n23006, n23007, 
      n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, 
      n23017, n23018, n23021, n23022, n23023, n23024, n23025, n23026, n23027, 
      n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23037, 
      n23038, n23039, n23040, n23041, n23042, n23043, n23045, n23046, n23047, 
      n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, 
      n23057, n23058, n23060, n23062, n23064, n23065, n23066, n23067, n23068, 
      n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, 
      n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, 
      n23088, n23089, n23090, n23092, n23093, n23094, n23096, n23100, n23101, 
      n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, 
      n23112, n23113, n23115, n23116, n23117, n23118, n23119, n23120, n23121, 
      n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23130, n23131, 
      n23132, n23136, n23137, n23138, n23139, n23140, n23143, n23144, n23145, 
      n23146, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, 
      n23158, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, 
      n23170, n23171, n23173, n23174, n23176, n23177, n23178, n23179, n23180, 
      n23181, n23182, n23183, n23184, n23185, n23186, n23188, n23189, n23190, 
      n23191, n23192, n23194, n23196, n23197, n23198, n23199, n23200, n23201, 
      n23202, n23203, n23205, n23206, n23207, n23209, n23210, n23211, n23212, 
      n23213, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, 
      n23224, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, 
      n23234, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, 
      n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23253, 
      n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, 
      n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, 
      n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, 
      n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, 
      n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, 
      n23300, n23301, n23302, n23303, n23304, n23306, n23307, n23308, n23310, 
      n23311, n23312, n23313, n23314, n23315, n23316, n23318, n23319, n23320, 
      n23321, n23322, n23324, n23326, n23328, n23329, n23330, n23331, n23332, 
      n23333, n23334, n23335, n23336, n23337, n23338, n23340, n23341, n23342, 
      n23343, n23344, n23346, n23347, n23348, n23349, n23350, n23351, n23352, 
      n23353, n23354, n23355, n23356, n23358, n23359, n23361, n23362, n23363, 
      n23364, n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, 
      n23374, n23375, n23376, n23377, n23382, n23383, n23384, n23385, n23386, 
      n23387, n23388, n23389, n23390, n23391, n23393, n23395, n23396, n23397, 
      n23398, n23399, n23400, n23402, n23403, n23404, n23405, n23406, n23407, 
      n23408, n23411, n23412, n23413, n23414, n23415, n23417, n23419, n23420, 
      n23421, n23422, n23424, n23425, n23426, n23427, n23429, n23430, n23431, 
      n23432, n23433, n23435, n23436, n23437, n23438, n23439, n23440, n23441, 
      n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, 
      n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, 
      n23460, n23461, n23462, n23463, n23464, n23465, n23467, n23468, n23469, 
      n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23478, n23479, 
      n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, 
      n23489, n23490, n23491, n23493, n23494, n23495, n23496, n23497, n23498, 
      n23499, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, 
      n23509, n23510, n23511, n23512, n23513, n23514, n23516, n23517, n23518, 
      n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, 
      n23528, n23529, n23530, n23532, n23533, n23534, n23535, n23536, n23537, 
      n23538, n23539, n23540, n23542, n23543, n23544, n23547, n23548, n23549, 
      n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23558, n23559, 
      n23560, n23561, n23562, n23564, n23565, n23566, n23567, n23569, n23570, 
      n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, 
      n23581, n23582, n23583, n23584, n23586, n23587, n23588, n23590, n23593, 
      n23594, n23595, n23597, n23598, n23600, n23601, n23602, n23603, n23604, 
      n23605, n23606, n23608, n23609, n23610, n23611, n23612, n23613, n23616, 
      n23618, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, 
      n23628, n23629, n23631, n23632, n23633, n23634, n23635, n23636, n23637, 
      n23638, n23639, n23640, n23642, n23643, n23644, n23646, n23647, n23649, 
      n23650, n23651, n23653, n23654, n23655, n23656, n23657, n23658, n23659, 
      n23660, n23663, n23664, n23665, n23666, n23668, n23669, n23670, n23671, 
      n23672, n23675, n23676, n23677, n23679, n23680, n23681, n23682, n23683, 
      n23684, n23685, n23688, n23689, n23690, n23691, n23692, n23694, n23695, 
      n23696, n23697, n23698, n23699, n23701, n23702, n23703, n23704, n23705, 
      n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, 
      n23715, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, 
      n23726, n23727, n23728, n23729, n23730, n23731, n23735, n23736, n23737, 
      n23738, n23739, n23740, n23741, n23742, n23745, n23746, n23747, n23748, 
      n23749, n23750, n23752, n23753, n23754, n23755, n23756, n23757, n23758, 
      n23759, n23760, n23763, n23764, n23765, n23766, n23767, n23768, n23769, 
      n23770, n23771, n23772, n23773, n23775, n23776, n23777, n23778, n23780, 
      n23781, n23782, n23784, n23785, n23786, n23787, n23788, n23790, n23791, 
      n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, 
      n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, 
      n23811, n23812, n23813, n23815, n23816, n23817, n23818, n23819, n23821, 
      n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23832, n23833, 
      n23834, n23835, n23840, n23841, n23842, n23843, n23847, n23848, n23849, 
      n23850, n23851, n23852, n23853, n23855, n23856, n23857, n23858, n23859, 
      n23860, n23862, n23864, n23866, n23867, n23868, n23869, n23870, n23871, 
      n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23880, n23881, 
      n23882, n23884, n23885, n23886, n23887, n23888, n23889, n23891, n23892, 
      n23894, n23895, n23896, n23897, n23899, n23901, n23902, n23903, n23904, 
      n23905, n23906, n23910, n23912, n23914, n23915, n23916, n23917, n23918, 
      n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23927, n23928, 
      n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23938, 
      n23939, n23940, n23942, n23943, n23944, n23945, n23946, n23947, n23949, 
      n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, 
      n23959, n23960, n23961, n23962, n23964, n23965, n23966, n23967, n23968, 
      n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23978, 
      n23981, n23982, n23984, n23987, n23988, n23989, n23990, n23991, n23992, 
      n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, 
      n24004, n24005, n24007, n24008, n24009, n24010, n24011, n24012, n24013, 
      n24014, n24015, n24016, n24017, n24018, n24020, n24021, n24024, n24025, 
      n24027, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, 
      n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24046, n24047, 
      n24048, n24049, n24050, n24051, n24052, n24053, n24056, n24057, n24059, 
      n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24069, 
      n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, 
      n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24089, 
      n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, 
      n24099, n24101, n24102, n24103, n24104, n24106, n24107, n24108, n24109, 
      n24110, n24111, n24112, n24114, n24115, n24116, n24117, n24118, n24119, 
      n24120, n24121, n24123, n24124, n24125, n24126, n24127, n24128, n24129, 
      n24130, n24131, n24132, n24133, n24134, n24135, n24137, n24138, n24139, 
      n24140, n24141, n24142, n24143, n24144, n24147, n24148, n24149, n24150, 
      n24152, n24153, n24154, n24156, n24157, n24158, n24159, n24161, n24162, 
      n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24171, n24172, 
      n24173, n24174, n24176, n24177, n24178, n24179, n24180, n24181, n24182, 
      n24183, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24193, 
      n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, 
      n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, 
      n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, 
      n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, 
      n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, 
      n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24248, n24249, 
      n24250, n24251, n24253, n24254, n24255, n24256, n24257, n24259, n24260, 
      n24262, n24263, n24265, n24266, n24267, n24268, n24269, n24270, n24271, 
      n24272, n24273, n24275, n24276, n24277, n24278, n24279, n24280, n24281, 
      n24283, n24284, n24285, n24286, n24288, n24289, n24290, n24292, n24293, 
      n24294, n24295, n24296, n24297, n24299, n24300, n24301, n24302, n24304, 
      n24305, n24306, n24308, n24309, n24310, n24311, n24312, n24313, n24314, 
      n24315, n24316, n24317, n24318, n24319, n24321, n24322, n24324, n24325, 
      n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, 
      n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, 
      n24344, n24346, n24347, n24348, n24349, n24350, n24351, n24353, n24354, 
      n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24364, 
      n24365, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, 
      n24376, n24377, n24378, n24379, n24382, n24383, n24384, n24385, n24386, 
      n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, 
      n24398, n24399, n24401, n24402, n24403, n24404, n24405, n24407, n24408, 
      n24409, n24410, n24411, n24412, n24413, n24415, n24416, n24417, n24418, 
      n24419, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, 
      n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, 
      n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, 
      n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, 
      n24456, n24457, n24459, n24460, n24461, n24462, n24463, n24466, n24467, 
      n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, 
      n24478, n24479, n24481, n24482, n24484, n24485, n24486, n24487, n24488, 
      n24489, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, 
      n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, 
      n24508, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, 
      n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, 
      n24528, n24529, n24531, n24532, n24533, n24536, n24537, n24538, n24539, 
      n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, 
      n24549, n24551, n24552, n24553, n24554, n24556, n24557, n24559, n24560, 
      n24561, n24562, n24563, n24564, n24565, n24567, n24568, n24569, n24570, 
      n24572, n24573, n24574, n24575, n24576, n24578, n24579, n24580, n24581, 
      n24582, n24583, n24584, n24585, n24587, n24588, n24590, n24591, n24592, 
      n24593, n24595, n24596, n24597, n24598, n24600, n24602, n24603, n24604, 
      n24605, n24606, n24607, n24609, n24610, n24611, n24613, n24615, n24616, 
      n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, 
      n24626, n24628, n24629, n24631, n24632, n24633, n24634, n24635, n24636, 
      n24637, n24638, n24639, n24642, n24643, n24644, n24645, n24646, n24647, 
      n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, 
      n24657, n24658, n24659, n24660, n24662, n24664, n24665, n24666, n24667, 
      n24668, n24671, n24672, n24673, n24674, n24675, n24676, n24678, n24679, 
      n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, 
      n24689, n24691, n24692, n24693, n24695, n24696, n24697, n24698, n24699, 
      n24701, n24702, n24703, n24704, n24705, n24707, n24708, n24709, n24710, 
      n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, 
      n24720, n24721, n24723, n24724, n24725, n24726, n24728, n24729, n24730, 
      n24732, n24733, n24734, n24735, n24737, n24738, n24740, n24741, n24742, 
      n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, 
      n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760, 
      n24761, n24762, n24763, n24764, n24766, n24768, n24769, n24770, n24771, 
      n24773, n24774, n24776, n24777, n24778, n24779, n24780, n24781, n24782, 
      n24783, n24785, n24786, n24787, n24788, n24789, n24790, n24792, n24793, 
      n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, 
      n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, 
      n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, 
      n24821, n24822, n24823, n24824, n24825, n24826, n24828, n24829, n24830, 
      n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, 
      n24840, n24841, n24842, n24843, n24845, n24846, n24847, n24848, n24849, 
      n24852, n24853, n24854, n24855, n24856, n24857, n24860, n24861, n24862, 
      n24863, n24864, n24865, n24866, n24867, n24869, n24870, n24873, n24874, 
      n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, 
      n24884, n24885, n24886, n24888, n24889, n24892, n24893, n24894, n24895, 
      n24896, n24897, n24899, n24901, n24902, n24903, n24904, n24905, n24906, 
      n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, 
      n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, 
      n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, 
      n24934, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, 
      n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24953, n24954, 
      n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24964, 
      n24965, n24966, n24967, n24968, n24969, n24970, n24972, n24973, n24974, 
      n24975, n24976, n24977, n24981, n24983, n24984, n24985, n24988, n24989, 
      n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, 
      n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, 
      n25009, n25010, n25012, n25013, n25014, n25015, n25017, n25019, n25020, 
      n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, 
      n25031, n25033, n25034, n25035, n25036, n25037, n25038, n25040, n25041, 
      n25042, n25043, n25044, n25045, n25046, n25048, n25049, n25050, n25051, 
      n25052, n25053, n25054, n25055, n25057, n25058, n25059, n25060, n25062, 
      n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, 
      n25072, n25074, n25076, n25078, n25079, n25081, n25082, n25083, n25084, 
      n25086, n25087, n25088, n25089, n25090, n25091, n25093, n25094, n25095, 
      n25097, n25098, n25100, n25102, n25104, n25105, n25106, n25107, n25108, 
      n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, 
      n25118, n25119, n25120, n25121, n25123, n25124, n25125, n25126, n25127, 
      n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, 
      n25138, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, 
      n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, 
      n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25165, n25166, 
      n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, 
      n25176, n25177, n25179, n25180, n25181, n25182, n25183, n25184, n25185, 
      n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, 
      n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, 
      n25204, n25205, n25206, n25207, n25208, n25210, n25211, n25213, n25214, 
      n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, 
      n25224, n25225, n25227, n25228, n25229, n25231, n25232, n25233, n25234, 
      n25235, n25236, n25237, n25238, n25239, n25242, n25243, n25245, n25246, 
      n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, 
      n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, 
      n25265, n25266, n25267, n25268, n25271, n25272, n25273, n25274, n25276, 
      n25277, n25278, n25279, n25280, n25281, n25282, n25284, n25285, n25286, 
      n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, 
      n25297, n25299, n25302, n25303, n25306, n25308, n25309, n25311, n25312, 
      n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25322, 
      n25323, n25324, n25325, n25326, n25328, n25329, n25330, n25331, n25332, 
      n25334, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, 
      n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25352, n25353, 
      n25354, n25355, n25356, n25357, n25358, n25360, n25361, n25362, n25364, 
      n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, 
      n25375, n25376, n25377, n25378, n25379, n25380, n25382, n25383, n25385, 
      n25387, n25388, n25390, n25391, n25392, n25394, n25396, n25397, n25398, 
      n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25409, 
      n25410, n25411, n25412, n25415, n25416, n25417, n25418, n25419, n25420, 
      n25424, n25425, n25427, n25428, n25429, n25430, n25432, n25433, n25434, 
      n25436, n25437, n25439, n25440, n25441, n25442, n25443, n25444, n25445, 
      n25446, n25447, n25449, n25450, n25452, n25453, n25454, n25455, n25456, 
      n25457, n25458, n25459, n25460, n25462, n25463, n25464, n25465, n25466, 
      n25467, n25468, n25470, n25471, n25472, n25473, n25474, n25475, n25476, 
      n25477, n25478, n25479, n25480, n25481, n25482, n25485, n25486, n25487, 
      n25488, n25490, n25492, n25493, n25494, n25495, n25496, n25497, n25498, 
      n25499, n25500, n25501, n25504, n25506, n25507, n25509, n25510, n25511, 
      n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, 
      n25522, n25523, n25526, n25527, n25529, n25530, n25531, n25534, n25535, 
      n25536, n25537, n25539, n25541, n25542, n25543, n25544, n25545, n25546, 
      n25547, n25548, n25549, n25550, n25552, n25554, n25555, n25556, n25557, 
      n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, 
      n25568, n25569, n25570, n25571, n25572, n25573, n25575, n25577, n25578, 
      n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, 
      n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25598, n25600, 
      n25602, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, 
      n25612, n25613, n25615, n25617, n25618, n25619, n25620, n25621, n25624, 
      n25627, n25628, n25630, n25632, n25633, n25634, n25636, n25637, n25638, 
      n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25648, 
      n25650, n25651, n25653, n25654, n25657, n25658, n25659, n25660, n25664, 
      n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, 
      n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, 
      n25684, n25685, n25686, n25687, n25689, n25691, n25692, n25693, n25694, 
      n25695, n25696, n25697, n25699, n25700, n25701, n25702, n25703, n25704, 
      n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, 
      n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, 
      n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, 
      n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, 
      n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, 
      n25750, n25751, n25752, n25753, n25755, n25756, n25757, n25760, n25761, 
      n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, 
      n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, 
      n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, 
      n25790, n25791, n25792, n25793, n25795, n25796, n25797, n25798, n25799, 
      n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, 
      n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, 
      n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, 
      n25828, n25829, n25830, n25832, n25833, n25834, n25835, n25836, n25837, 
      n25838, n25839, n25840, n25841, n25843, n25844, n25845, n25846, n25847, 
      n25848, n25849, n25851, n25852, n25853, n25854, n25855, n25856, n25857, 
      n25858, n25859, n25860, n25861, n25863, n25864, n25865, n25866, n25867, 
      n25868, n25870, n25871, n25872, n25874, n25875, n25876, n25877, n25878, 
      n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, 
      n25889, n25890, n25891, n25892, n25893, n25894, n25896, n25897, n25899, 
      n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, 
      n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, 
      n25918, n25919, n25920, n25922, n25923, n25924, n25925, n25926, n25927, 
      n25929, n25941, n25942, n25943, n25944, n25945, n25947, n25951, n25954, 
      n25959, n25960, n25961, n25962, n25963, n25966, n25967, n25968, n25969, 
      n25971, n25973, n25974, n25975, n25977, n25979, n25980, n25981, n25985, 
      n25987, n25988, n25990, n25991, n25993, n25994, n25995, n25996, n25997, 
      n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, 
      n26007, n26008, n26012, n26013, n26014, n26015, n26016, n26018, n26020, 
      n26021, n26022, n26023, n26025, n26026, n26027, n26028, n26029, n26030, 
      n26031, n26032, n26033, n26035, n26036, n26037, n26038, n26040, n26041, 
      n26043, n26045, n26046, n26047, n26049, n26051, n26053, n26054, n26055, 
      n26056, n26057, n26058, n26059, n26060, n26061, n26065, n26067, n26068, 
      n26069, n26070, n26072, n26073, n26074, n26075, n26076, n26078, n26079, 
      n26081, n26082, n26083, n26084, n26085, n26087, n26088, n26089, n26093, 
      n26094, n26096, n26097, n26098, n26100, n26101, n26102, n26103, n26104, 
      n26106, n26108, n26109, n26111, n26113, n26114, n26115, n26116, n26118, 
      n26120, n26121, n26123, n26124, n26125, n26126, n26127, n26130, n26133, 
      n26140, n26142, n26144, n26145, n26150, n26152, n26153, n26154, n26155, 
      n26156, n26157, n26158, n26160, n26161, n26162, n26163, n26164, n26165, 
      n26166, n26167, n26168, n26169, n26170, n26172, n26173, n26175, n26176, 
      n26178, n26181, n26182, n26185, n26193, n26194, n26195, n26197, n26198, 
      n26199, n26202, n26203, n26204, n26206, n26207, n26208, n26211, n26212, 
      n26214, n26215, n26216, n26217, n26220, n26221, n26222, n26224, n26228, 
      n26230, n26231, n26232, n26233, n26236, n26237, n26238, n26239, n26241, 
      n26242, n26243, n26244, n26247, n26249, n26250, n26251, n26253, n26255, 
      n26256, n26257, n26261, n26262, n26265, n26268, n26270, n26272, n26274, 
      n26275, n26276, n26277, n26278, n26279, n26281, n26282, n26283, n26284, 
      n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, 
      n26298, n26300, n26301, n26302, n26304, n26305, n26307, n26311, n26312, 
      n26314, n26317, n26318, n26320, n26322, n26324, n26325, n26326, n26328, 
      n26330, n26333, n26334, n26336, n26337, n26338, n26340, n26341, n26343, 
      n26345, n26347, n26350, n26351, n26355, n26357, n26358, n26362, n26363, 
      n26365, n26367, n26368, n26369, n26370, n26371, n26373, n26374, n26375, 
      n26376, n26378, n26380, n26383, n26384, n26385, n26386, n26387, n26388, 
      n26389, n26390, n26391, n26392, n26393, n26394, n26397, n26398, n26399, 
      n26400, n26401, n26404, n26406, n26407, n26408, n26409, n26410, n26411, 
      n26412, n26413, n26415, n26416, n26417, n26418, n26422, n26423, n26424, 
      n26426, n26429, n26431, n26432, n26433, n26435, n26436, n26438, n26439, 
      n26440, n26442, n26443, n26444, n26445, n26447, n26448, n26451, n26452, 
      n26453, n26455, n26456, n26458, n26459, n26462, n26464, n26465, n26466, 
      n26468, n26469, n26471, n26472, n26474, n26478, n26479, n26484, n26485, 
      n26487, n26488, n26490, n26492, n26493, n26494, n26497, n26499, n26501, 
      n26502, n26503, n26504, n26505, n26506, n26507, n26511, n26513, n26515, 
      n26516, n26518, n26520, n26521, n26522, n26524, n26525, n26526, n26527, 
      n26528, n26529, n26530, n26533, n26534, n26537, n26540, n26542, n26543, 
      n26544, n26545, n26547, n26550, n26551, n26552, n26553, n26554, n26555, 
      n26556, n26557, n26562, n26563, n26566, n26567, n26568, n26569, n26570, 
      n26571, n26572, n26573, n26575, n26576, n26579, n26580, n26581, n26582, 
      n26583, n26585, n26587, n26588, n26589, n26590, n26591, n26593, n26594, 
      n26595, n26597, n26600, n26603, n26606, n26607, n26608, n26609, n26611, 
      n26612, n26614, n26615, n26617, n26622, n26623, n26625, n26627, n26628, 
      n26630, n26631, n26632, n26633, n26635, n26637, n26640, n26641, n26642, 
      n26643, n26644, n26646, n26647, n26648, n26655, n26656, n26660, n26663, 
      n26665, n26666, n26667, n26671, n26674, n26677, n26679, n26680, n26682, 
      n26683, n26688, n26690, n26691, n26692, n26693, n26696, n26699, n26701, 
      n26702, n26705, n26708, n26709, n26710, n26711, n26712, n26713, n26715, 
      n26716, n26717, n26720, n26722, n26724, n26725, n26726, n26727, n26728, 
      n26730, n26731, n26732, n26733, n26735, n26736, n26738, n26739, n26740, 
      n26741, n26742, n26744, n26745, n26747, n26750, n26751, n26753, n26754, 
      n26755, n26756, n26758, n26761, n26762, n26765, n26766, n26767, n26768, 
      n26769, n26772, n26774, n26775, n26777, n26778, n26780, n26782, n26784, 
      n26785, n26787, n26790, n26791, n26793, n26794, n26795, n26796, n26798, 
      n26799, n26800, n26801, n26803, n26806, n26807, n26808, n26810, n26812, 
      n26813, n26814, n26815, n26817, n26818, n26821, n26822, n26823, n26825, 
      n26827, n26829, n26830, n26834, n26835, n26836, n26837, n26842, n26844, 
      n26845, n26846, n26848, n26851, n26854, n26855, n26856, n26858, n26861, 
      n26862, n26863, n26865, n26867, n26868, n26869, n26872, n26873, n26874, 
      n26875, n26877, n26878, n26881, n26882, n26883, n26884, n26885, n26886, 
      n26887, n26888, n26889, n26890, n26891, n26892, n26896, n26897, n26898, 
      n26899, n26900, n26903, n26904, n26907, n26909, n26912, n26913, n26914, 
      n26915, n26916, n26917, n26918, n26920, n26921, n26922, n26923, n26924, 
      n26925, n26927, n26929, n26930, n26931, n26933, n26934, n26936, n26937, 
      n26938, n26941, n26942, n26945, n26947, n26948, n26949, n26950, n26953, 
      n26954, n26955, n26956, n26957, n26958, n26960, n26961, n26962, n26965, 
      n26966, n26967, n26969, n26971, n26974, n26976, n26977, n26978, n26979, 
      n26980, n26983, n26986, n26987, n26988, n26990, n26991, n26992, n26993, 
      n26994, n26995, n26996, n26997, n26998, n27000, n27004, n27005, n27007, 
      n27008, n27010, n27011, n27012, n27014, n27015, n27016, n27018, n27019, 
      n27020, n27021, n27023, n27024, n27026, n27028, n27033, n27034, n27038, 
      n27041, n27042, n27044, n27046, n27047, n27049, n27050, n27052, n27053, 
      n27054, n27055, n27057, n27058, n27060, n27062, n27063, n27064, n27065, 
      n27066, n27067, n27070, n27072, n27073, n27075, n27076, n27077, n27078, 
      n27079, n27080, n27081, n27082, n27088, n27090, n27091, n27092, n27094, 
      n27097, n27098, n27099, n27100, n27101, n27103, n27104, n27105, n27106, 
      n27110, n27111, n27113, n27114, n27115, n27117, n27118, n27119, n27120, 
      n27121, n27122, n27123, n27125, n27126, n27127, n27128, n27129, n27130, 
      n27131, n27132, n27134, n27135, n27136, n27137, n27138, n27139, n27142, 
      n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, 
      n27152, n27153, n27154, n27155, n27156, n27157, n27159, n27160, n27162, 
      n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, 
      n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, 
      n27182, n27183, n27184, n27185, n27186, n27188, n27189, n27190, n27191, 
      n27192, n27193, n27196, n27198, n27200, n27201, n27202, n27203, n27207, 
      n27208, n27211, n27212, n27214, n27215, n27217, n27218, n27219, n27220, 
      n27225, n27226, n27227, n27228, n27230, n27232, n27233, n27234, n27236, 
      n27237, n27238, n27240, n27242, n27243, n27244, n27245, n27246, n27248, 
      n27249, n27252, n27253, n27257, n27259, n27261, n27262, n27263, n27265, 
      n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, 
      n27275, n27276, n27277, n27279, n27281, n27282, n27283, n27284, n27285, 
      n27289, n27290, n27294, n27296, n27297, n27298, n27299, n27300, n27301, 
      n27302, n27303, n27305, n27307, n27308, n27309, n27311, n27312, n27314, 
      n27315, n27316, n27317, n27318, n27320, n27321, n27324, n27326, n27329, 
      n27330, n27332, n27334, n27336, n27337, n27338, n27340, n27341, n27342, 
      n27343, n27344, n27345, n27349, n27352, n27353, n27354, n27357, n27358, 
      n27359, n27360, n27361, n27362, n27363, n27365, n27367, n27368, n27369, 
      n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27381, 
      n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390, 
      n27391, n27392, n27395, n27396, n27397, n27398, n27401, n27402, n27403, 
      n27406, n27408, n27409, n27410, n27411, n27412, n27413, n27415, n27416, 
      n27419, n27420, n27423, n27424, n27426, n27428, n27429, n27430, n27431, 
      n27432, n27435, n27436, n27437, n27439, n27440, n27441, n27442, n27443, 
      n27444, n27445, n27446, n27450, n27451, n27453, n27454, n27455, n27456, 
      n27457, n27458, n27459, n27460, n27461, n27462, n27466, n27471, n27472, 
      n27474, n27475, n27478, n27479, n27480, n27481, n27482, n27485, n27486, 
      n27487, n27490, n27491, n27495, n27500, n27501, n27503, n27504, n27505, 
      n27506, n27509, n27514, n27515, n27516, n27517, n27518, n27520, n27523, 
      n27525, n27526, n27528, n27529, n27531, n27532, n27534, n27535, n27537, 
      n27538, n27539, n27541, n27542, n27543, n27544, n27545, n27548, n27550, 
      n27551, n27552, n27553, n27555, n27556, n27560, n27561, n27563, n27565, 
      n27566, n27567, n27569, n27570, n27571, n27573, n27574, n27575, n27577, 
      n27580, n27582, n27583, n27585, n27586, n27587, n27588, n27589, n27590, 
      n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27599, n27600, 
      n27601, n27604, n27605, n27607, n27608, n27609, n27610, n27611, n27612, 
      n27613, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622, 
      n27624, n27625, n27627, n27628, n27629, n27630, n27631, n27633, n27635, 
      n27637, n27638, n27639, n27641, n27642, n27643, n27645, n27646, n27648, 
      n27649, n27650, n27651, n27652, n27654, n27655, n27658, n27659, n27660, 
      n27661, n27662, n27664, n27667, n27668, n27669, n27670, n27672, n27673, 
      n27676, n27678, n27679, n27680, n27683, n27684, n27685, n27686, n27687, 
      n27688, n27689, n27690, n27691, n27693, n27694, n27695, n27696, n27697, 
      n27698, n27699, n27701, n27703, n27704, n27706, n27707, n27708, n27709, 
      n27711, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721, 
      n27724, n27726, n27728, n27729, n27731, n27732, n27733, n27734, n27735, 
      n27736, n27737, n27738, n27739, n27741, n27743, n27745, n27747, n27748, 
      n27750, n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, 
      n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, 
      n27769, n27771, n27773, n27775, n27776, n27778, n27779, n27781, n27785, 
      n27786, n27787, n27788, n27790, n27791, n27792, n27793, n27797, n27798, 
      n27799, n27801, n27802, n27804, n27805, n27806, n27807, n27808, n27811, 
      n27812, n27814, n27816, n27818, n27819, n27823, n27824, n27825, n27826, 
      n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836, 
      n27837, n27838, n27840, n27841, n27842, n27845, n27846, n27850, n27851, 
      n27852, n27854, n27856, n27857, n27860, n27861, n27862, n27863, n27864, 
      n27865, n27866, n27867, n27868, n27872, n27873, n27875, n27876, n27877, 
      n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27886, n27887, 
      n27889, n27893, n27894, n27895, n27896, n27897, n27899, n27900, n27901, 
      n27902, n27904, n27907, n27908, n27909, n27910, n27911, n27912, n27914, 
      n27916, n27919, n27920, n27921, n27922, n27923, n27925, n27926, n27929, 
      n27930, n27931, n27933, n27934, n27936, n27937, n27938, n27939, n27940, 
      n27941, n27942, n27943, n27946, n27947, n27950, n27951, n27952, n27953, 
      n27954, n27955, n27957, n27958, n27959, n27960, n27961, n27962, n27963, 
      n27965, n27968, n27969, n27970, n27971, n27972, n27973, n27975, n27976, 
      n27977, n27980, n27981, n27982, n27984, n27987, n27988, n27990, n27991, 
      n27992, n27993, n27994, n27995, n27996, n27998, n28000, n28001, n28002, 
      n28003, n28004, n28005, n28009, n28010, n28011, n28012, n28014, n28016, 
      n28017, n28018, n28019, n28020, n28021, n28022, n28025, n28027, n28028, 
      n28029, n28030, n28031, n28034, n28035, n28037, n28038, n28039, n28040, 
      n28043, n28052, n28056, n28057, n28058, n28059, n28061, n28062, n28064, 
      n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28077, 
      n28078, n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28091, 
      n28093, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28104, 
      n28105, n28107, n28108, n28109, n28110, n28111, n28113, n28114, n28116, 
      n28117, n28118, n28119, n28120, n28121, n28123, n28124, n28126, n28128, 
      n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138, 
      n28139, n28141, n28142, n28144, n28147, n28150, n28151, n28152, n28153, 
      n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28162, n28163, 
      n28166, n28167, n28170, n28171, n28172, n28174, n28175, n28177, n28178, 
      n28179, n28181, n28183, n28186, n28188, n28190, n28194, n28196, n28197, 
      n28199, n28200, n28202, n28203, n28205, n28206, n28208, n28209, n28210, 
      n28211, n28214, n28216, n28217, n28218, n28219, n28220, n28222, n28223, 
      n28225, n28226, n28227, n28228, n28231, n28232, n28234, n28235, n28236, 
      n28237, n28238, n28239, n28240, n28242, n28243, n28244, n28245, n28246, 
      n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28260, 
      n28261, n28262, n28263, n28265, n28266, n28268, n28269, n28270, n28273, 
      n28275, n28276, n28277, n28278, n28279, n28281, n28283, n28285, n28286, 
      n28287, n28288, n28289, n28293, n28295, n28296, n28297, n28298, n28299, 
      n28300, n28302, n28303, n28304, n28306, n28307, n28308, n28309, n28311, 
      n28312, n28313, n28314, n28315, n28316, n28318, n28320, n28321, n28323, 
      n28324, n28327, n28328, n28329, n28330, n28331, n28332, n28338, n28340, 
      n28342, n28343, n28344, n28345, n28347, n28348, n28349, n28350, n28351, 
      n28353, n28354, n28355, n28356, n28357, n28358, n28361, n28364, n28365, 
      n28366, n28367, n28371, n28372, n28373, n28374, n28375, n28376, n28378, 
      n28379, n28380, n28381, n28382, n28383, n28385, n28386, n28387, n28388, 
      n28390, n28391, n28393, n28395, n28396, n28397, n28399, n28400, n28401, 
      n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, 
      n28411, n28413, n28414, n28415, n28416, n28418, n28419, n28420, n28421, 
      n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430, 
      n28431, n28432, n28435, n28436, n28437, n28438, n28439, n28441, n28442, 
      n28443, n28444, n28446, n28447, n28448, n28449, n28450, n28451, n28452, 
      n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461, 
      n28462, n28463, n28465, n28466, n28467, n28469, n28470, n28471, n28472, 
      n28473, n28474, n28475, n28478, n28479, n28480, n28482, n28483, n28484, 
      n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493, 
      n28494, n28495, n28496, n28497, n28498, n28501, n28502, n28503, n28504, 
      n28505, n28506, n28507, n28509, n28510, n28513, n28514, n28516, n28517, 
      n28519, n28520, n28522, n28523, n28524, n28525, n28526, n28527, n28528, 
      n28530, n28531, n28532, n28534, n28536, n28538, n28539, n28540, n28541, 
      n28542, n28543, n28544, n28545, n28548, n28549, n28552, n28553, n28554, 
      n28555, n28557, n28560, n28562, n28564, n28565, n28566, n28567, n28568, 
      n28571, n28573, n28574, n28575, n28578, n28579, n28580, n28581, n28584, 
      n28585, n28586, n28587, n28589, n28590, n28591, n28592, n28593, n28594, 
      n28595, n28600, n28601, n28602, n28603, n28605, n28606, n28607, n28608, 
      n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28621, 
      n28622, n28623, n28624, n28625, n28626, n28627, n28631, n28632, n28633, 
      n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, 
      n28644, n28645, n28647, n28648, n28649, n28651, n28652, n28654, n28655, 
      n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665, 
      n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676, 
      n28680, n28681, n28683, n28684, n28685, n28686, n28687, n28688, n28689, 
      n28691, n28692, n28694, n28696, n28697, n28698, n28699, n28700, n28701, 
      n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710, 
      n28711, n28712, n28714, n28715, n28721, n28722, n28723, n28724, n28725, 
      n28726, n28728, n28729, n28730, n28731, n28733, n28734, n28735, n28736, 
      n28737, n28738, n28740, n28743, n28744, n28745, n28746, n28747, n28748, 
      n28750, n28751, n28752, n28753, n28754, n28755, n28757, n28758, n28759, 
      n28760, n28761, n28762, n28763, n28765, n28767, n28769, n28770, n28771, 
      n28773, n28775, n28776, n28777, n28778, n28779, n28781, n28782, n28783, 
      n28784, n28786, n28788, n28789, n28791, n28796, n28797, n28799, n28800, 
      n28801, n28802, n28803, n28806, n28807, n28811, n28812, n28813, n28814, 
      n28815, n28816, n28817, n28818, n28819, n28821, n28822, n28823, n28824, 
      n28825, n28826, n28827, n28829, n28830, n28831, n28833, n28835, n28836, 
      n28837, n28838, n28839, n28840, n28844, n28846, n28847, n28848, n28849, 
      n28850, n28852, n28853, n28854, n28855, n28856, n28857, n28859, n28860, 
      n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869, 
      n28870, n28872, n28873, n28875, n28876, n28877, n28878, n28880, n28882, 
      n28883, n28885, n28886, n28887, n28888, n28889, n28891, n28893, n28894, 
      n28895, n28896, n28897, n28898, n28899, n28900, n28902, n28903, n28904, 
      n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, 
      n28917, n28918, n28921, n28922, n28923, n28924, n28926, n28927, n28929, 
      n28931, n28932, n28933, n28934, n28935, n28937, n28938, n28939, n28940, 
      n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949, 
      n28950, n28951, n28952, n28953, n28954, n28956, n28957, n28958, n28964, 
      n28967, n28968, n28970, n28972, n28973, n28974, n28975, n28977, n28978, 
      n28979, n28981, n28982, n28983, n28987, n28989, n28990, n28992, n28993, 
      n28995, n28996, n28998, n28999, n29000, n29001, n29002, n29003, n29004, 
      n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29018, n29020, 
      n29021, n29022, n29026, n29027, n29028, n29029, n29030, n29032, n29033, 
      n29034, n29035, n29037, n29039, n29040, n29042, n29043, n29044, n29046, 
      n29047, n29048, n29049, n29050, n29051, n29052, n29054, n29056, n29057, 
      n29060, n29061, n29062, n29063, n29064, n29068, n29069, n29070, n29071, 
      n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, 
      n29081, n29082, n29084, n29085, n29087, n29088, n29089, n29090, n29093, 
      n29094, n29095, n29098, n29099, n29101, n29102, n29106, n29107, n29108, 
      n29110, n29111, n29114, n29115, n29116, n29118, n29119, n29120, n29121, 
      n29122, n29123, n29124, n29127, n29130, n29131, n29133, n29134, n29135, 
      n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29146, n29147, 
      n29148, n29149, n29152, n29153, n29155, n29156, n29157, n29158, n29159, 
      n29160, n29162, n29167, n29168, n29169, n29170, n29172, n29173, n29174, 
      n29175, n29176, n29178, n29180, n29182, n29184, n29185, n29187, n29189, 
      n29190, n29194, n29196, n29198, n29200, n29201, n29202, n29203, n29205, 
      n29206, n29207, n29208, n29209, n29211, n29212, n29213, n29214, n29215, 
      n29216, n29217, n29218, n29220, n29221, n29222, n29223, n29224, n29225, 
      n29227, n29228, n29230, n29231, n29232, n29233, n29234, n29235, n29236, 
      n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29250, 
      n29252, n29253, n29254, n29255, n29256, n29258, n29259, n29260, n29261, 
      n29262, n29263, n29266, n29268, n29269, n29270, n29271, n29272, n29273, 
      n29274, n29275, n29277, n29278, n29279, n29280, n29281, n29282, n29283, 
      n29284, n29285, n29286, n29287, n29288, n29291, n29292, n29293, n29294, 
      n29296, n29299, n29302, n29303, n29304, n29305, n29306, n29307, n29308, 
      n29309, n29312, n29313, n29314, n29315, n29317, n29318, n29320, n29321, 
      n29322, n29323, n29325, n29328, n29329, n29330, n29331, n29334, n29335, 
      n29336, n29337, n29338, n29339, n29341, n29342, n29343, n29344, n29345, 
      n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354, 
      n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363, 
      n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372, 
      n29373, n29375, n29376, n29378, n29379, n29380, n29382, n29383, n29384, 
      n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, 
      n29394, n29395, n29396, n29397, n29398, n29400, n29401, n29402, n29404, 
      n29405, n29406, n29407, n29408, n29409, n29412, n29413, n29415, n29416, 
      n29417, n29418, n29420, n29421, n29422, n29423, n29424, n29426, n29427, 
      n29428, n29430, n29431, n29432, n29433, n29434, n29435, n29437, n29438, 
      n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, 
      n29450, n29451, n29453, n29454, n29455, n29457, n29458, n29460, n29461, 
      n29462, n29463, n29464, n29467, n29469, n29470, n29471, n29472, n29473, 
      n29474, n29475, n29476, n29477, n29480, n29481, n29482, n29483, n29485, 
      n29486, n29487, n29488, n29489, n29492, n29494, n29495, n29497, n29498, 
      n29499, n29501, n29502, n29503, n29507, n29508, n29509, n29510, n29512, 
      n29514, n29515, n29517, n29518, n29520, n29521, n29522, n29523, n29525, 
      n29526, n29527, n29528, n29531, n29532, n29534, n29536, n29537, n29538, 
      n29539, n29540, n29541, n29543, n29545, n29547, n29548, n29550, n29551, 
      n29552, n29553, n29554, n29555, n29557, n29559, n29560, n29561, n29562, 
      n29563, n29566, n29567, n29568, n29570, n29572, n29573, n29574, n29575, 
      n29576, n29577, n29578, n29580, n29581, n29582, n29583, n29584, n29586, 
      n29588, n29589, n29590, n29593, n29594, n29595, n29597, n29598, n29600, 
      n29602, n29603, n29605, n29606, n29607, n29608, n29609, n29610, n29614, 
      n29615, n29618, n29620, n29621, n29623, n29624, n29626, n29628, n29629, 
      n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29638, n29639, 
      n29642, n29643, n29644, n29645, n29646, n29648, n29650, n29651, n29652, 
      n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661, 
      n29662, n29663, n29664, n29666, n29667, n29668, n29670, n29671, n29672, 
      n29673, n29674, n29675, n29676, n29678, n29679, n29680, n29681, n29682, 
      n29683, n29684, n29687, n29688, n29689, n29690, n29692, n29693, n29695, 
      n29696, n29699, n29702, n29704, n29705, n29706, n29707, n29708, n29709, 
      n29711, n29712, n29714, n29715, n29717, n29718, n29719, n29720, n29721, 
      n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730, 
      n29731, n29732, n29733, n29734, n29736, n29737, n29738, n29739, n29740, 
      n29741, n29742, n29743, n29748, n29750, n29751, n29753, n29754, n29755, 
      n29757, n29758, n29759, n29761, n29762, n29763, n29765, n29767, n29768, 
      n29769, n29771, n29772, n29773, n29774, n29776, n29777, n29778, n29780, 
      n29781, n29784, n29785, n29787, n29788, n29789, n29790, n29791, n29792, 
      n29795, n29796, n29799, n29800, n29801, n29802, n29803, n29804, n29806, 
      n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, 
      n29817, n29818, n29819, n29820, n29821, n29823, n29825, n29827, n29828, 
      n29829, n29830, n29832, n29833, n29834, n29835, n29836, n29837, n29838, 
      n29839, n29840, n29841, n29843, n29844, n29845, n29846, n29847, n29848, 
      n29849, n29850, n29851, n29853, n29854, n29855, n29856, n29858, n29863, 
      n29864, n29865, n29866, n29867, n29868, n29870, n29872, n29873, n29875, 
      n29876, n29877, n29878, n29879, n29880, n29882, n29883, n29885, n29888, 
      n29890, n29895, n29896, n29898, n29899, n29900, n29901, n29903, n29904, 
      n29905, n29906, n29907, n29908, n29909, n29911, n29912, n29913, n29914, 
      n29915, n29916, n29918, n29919, n29920, n29921, n29922, n29924, n29927, 
      n29928, n29930, n29931, n29932, n29933, n29934, n29936, n29937, n29938, 
      n29943, n29944, n29946, n29947, n29949, n29951, n29952, n29953, n29954, 
      n29955, n29957, n29958, n29960, n29962, n29963, n29964, n29965, n29967, 
      n29969, n29970, n29972, n29973, n29975, n29976, n29977, n29978, n29980, 
      n29981, n29982, n29983, n29985, n29986, n29987, n29988, n29989, n29993, 
      n29994, n29995, n29997, n30000, n30001, n30003, n30004, n30005, n30006, 
      n30007, n30008, n30010, n30011, n30012, n30013, n30014, n30015, n30016, 
      n30017, n30018, n30019, n30020, n30021, n30022, n30025, n30028, n30029, 
      n30031, n30032, n30033, n30036, n30038, n30039, n30041, n30042, n30044, 
      n30045, n30047, n30048, n30049, n30050, n30054, n30057, n30058, n30059, 
      n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30069, 
      n30070, n30071, n30072, n30074, n30075, n30076, n30078, n30079, n30080, 
      n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, 
      n30090, n30091, n30093, n30094, n30096, n30097, n30098, n30099, n30102, 
      n30104, n30105, n30106, n30107, n30109, n30110, n30111, n30112, n30114, 
      n30115, n30116, n30117, n30118, n30119, n30121, n30122, n30123, n30124, 
      n30125, n30126, n30127, n30129, n30130, n30131, n30134, n30135, n30136, 
      n30137, n30138, n30139, n30140, n30142, n30143, n30144, n30145, n30146, 
      n30148, n30149, n30151, n30152, n30154, n30155, n30156, n30157, n30159, 
      n30163, n30165, n30167, n30168, n30169, n30171, n30172, n30173, n30174, 
      n30175, n30176, n30177, n30180, n30181, n30182, n30183, n30185, n30186, 
      n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30195, n30197, 
      n30198, n30199, n30200, n30202, n30203, n30204, n30205, n30207, n30209, 
      n30212, n30214, n30215, n30216, n30218, n30219, n30220, n30221, n30222, 
      n30223, n30224, n30225, n30226, n30227, n30229, n30230, n30231, n30232, 
      n30233, n30234, n30235, n30236, n30237, n30240, n30241, n30243, n30246, 
      n30247, n30248, n30250, n30251, n30252, n30255, n30257, n30258, n30259, 
      n30262, n30265, n30267, n30269, n30270, n30271, n30272, n30273, n30274, 
      n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283, 
      n30284, n30285, n30288, n30289, n30290, n30291, n30293, n30294, n30295, 
      n30296, n30297, n30301, n30302, n30303, n30304, n30305, n30306, n30307, 
      n30308, n30309, n30311, n30313, n30314, n30315, n30316, n30317, n30318, 
      n30319, n30320, n30321, n30322, n30323, n30326, n30327, n30328, n30329, 
      n30330, n30331, n30332, n30333, n30334, n30336, n30338, n30339, n30340, 
      n30341, n30342, n30344, n30345, n30346, n30348, n30349, n30353, n30354, 
      n30355, n30356, n30357, n30358, n30359, n30360, n30362, n30364, n30365, 
      n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30374, n30375, 
      n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387, 
      n30388, n30389, n30390, n30391, n30393, n30394, n30396, n30398, n30400, 
      n30401, n30402, n30403, n30404, n30405, n30407, n30408, n30409, n30410, 
      n30411, n30412, n30413, n30414, n30417, n30418, n30420, n30421, n30423, 
      n30425, n30426, n30427, n30428, n30429, n30430, n30433, n30435, n30436, 
      n30437, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446, 
      n30447, n30448, n30449, n30450, n30453, n30454, n30455, n30458, n30459, 
      n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30469, n30470, 
      n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30479, n30480, 
      n30482, n30483, n30486, n30487, n30488, n30489, n30492, n30493, n30494, 
      n30495, n30496, n30497, n30498, n30501, n30502, n30503, n30504, n30505, 
      n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, 
      n30515, n30517, n30521, n30522, n30523, n30524, n30526, n30527, n30528, 
      n30529, n30530, n30532, n30535, n30536, n30537, n30538, n30539, n30540, 
      n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549, 
      n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558, 
      n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30568, n30569, 
      n30570, n30571, n30572, n30573, n30574, n30575, n30578, n30579, n30583, 
      n30584, n30586, n30587, n30592, n30593, n30594, n30595, n30596, n30597, 
      n30598, n30600, n30601, n30602, n30603, n30607, n30608, n30610, n30612, 
      n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, 
      n30623, n30624, n30625, n30626, n30627, n30628, n30631, n30632, n30633, 
      n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30643, 
      n30644, n30645, n30646, n30648, n30649, n30651, n30652, n30653, n30654, 
      n30656, n30658, n30660, n30661, n30663, n30664, n30666, n30668, n30669, 
      n30670, n30671, n30673, n30676, n30677, n30678, n30679, n30681, n30682, 
      n30685, n30686, n30687, n30688, n30690, n30691, n30692, n30693, n30694, 
      n30695, n30696, n30697, n30698, n30699, n30700, n30702, n30703, n30705, 
      n30706, n30707, n30708, n30710, n30711, n30712, n30713, n30714, n30715, 
      n30716, n30717, n30718, n30720, n30721, n30722, n30723, n30724, n30725, 
      n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734, 
      n30736, n30737, n30740, n30741, n30742, n30743, n30744, n30745, n30746, 
      n30747, n30748, n30749, n30753, n30754, n30755, n30757, n30758, n30760, 
      n30762, n30763, n30765, n30766, n30767, n30768, n30769, n30770, n30771, 
      n30774, n30776, n30777, n30778, n30779, n30780, n30781, n30783, n30784, 
      n30789, n30790, n30792, n30793, n30794, n30795, n30798, n30800, n30802, 
      n30803, n30805, n30806, n30807, n30808, n30810, n30811, n30813, n30815, 
      n30816, n30817, n30818, n30819, n30820, n30822, n30824, n30825, n30826, 
      n30828, n30830, n30831, n30832, n30833, n30837, n30838, n30840, n30843, 
      n30844, n30845, n30846, n30849, n30850, n30852, n30853, n30854, n30855, 
      n30856, n30857, n30858, n30861, n30862, n30863, n30865, n30866, n30867, 
      n30868, n30869, n30870, n30871, n30872, n30873, n30875, n30876, n30877, 
      n30878, n30879, n30880, n30881, n30882, n30883, n30885, n30886, n30887, 
      n30888, n30889, n30892, n30894, n30895, n30898, n30899, n30900, n30901, 
      n30902, n30904, n30905, n30906, n30907, n30908, n30909, n30912, n30913, 
      n30914, n30915, n30917, n30919, n30922, n30923, n30924, n30925, n30926, 
      n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936, 
      n30937, n30938, n30940, n30942, n30943, n30945, n30946, n30948, n30949, 
      n30951, n30952, n30953, n30954, n30955, n30957, n30958, n30959, n30960, 
      n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, 
      n30970, n30971, n30972, n30973, n30976, n30978, n30979, n30980, n30981, 
      n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990, 
      n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999, 
      n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31009, n31012, 
      n31015, n31016, n31017, n31019, n31021, n31022, n31025, n31026, n31028, 
      n31029, n31030, n31032, n31033, n31034, n31036, n31037, n31039, n31040, 
      n31041, n31042, n31043, n31044, n31046, n31047, n31048, n31051, n31052, 
      n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31062, n31063, 
      n31065, n31066, n31070, n31071, n31072, n31073, n31074, n31075, n31077, 
      n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, 
      n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, 
      n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, 
      n31105, n31106, n31108, n31109, n31110, n31111, n31112, n31113, n31114, 
      n31115, n31116, n31117, n31118, n31120, n31121, n31122, n31123, n31124, 
      n31126, n31127, n31128, n31129, n31132, n31133, n31135, n31136, n31137, 
      n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, 
      n31147, n31148, n31149, n31150, n31151, n31152, n31155, n31156, n31157, 
      n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31167, 
      n31168, n31169, n31170, n31171, n31173, n31174, n31175, n31177, n31178, 
      n31179, n31180, n31181, n31182, n31184, n31185, n31186, n31188, n31189, 
      n31190, n31191, n31194, n31195, n31197, n31200, n31201, n31202, n31203, 
      n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31213, n31214, 
      n31215, n31216, n31217, n31218, n31220, n31221, n31223, n31225, n31226, 
      n31228, n31229, n31231, n31232, n31233, n31234, n31235, n31236, n31237, 
      n31238, n31239, n31241, n31242, n31243, n31244, n31245, n31246, n31247, 
      n31248, n31250, n31251, n31252, n31253, n31254, n31258, n31259, n31260, 
      n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31271, 
      n31272, n31273, n31274, n31275, n31277, n31279, n31280, n31281, n31282, 
      n31284, n31285, n31286, n31287, n31288, n31290, n31291, n31292, n31293, 
      n31294, n31295, n31296, n31297, n31301, n31303, n31306, n31308, n31309, 
      n31311, n31312, n31314, n31315, n31316, n31317, n31318, n31319, n31320, 
      n31321, n31323, n31324, n31325, n31327, n31329, n31330, n31331, n31333, 
      n31334, n31335, n31336, n31338, n31339, n31340, n31341, n31342, n31344, 
      n31345, n31346, n31348, n31349, n31350, n31351, n31352, n31354, n31355, 
      n31356, n31357, n31358, n31359, n31360, n31361, n31363, n31365, n31366, 
      n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31377, 
      n31378, n31379, n31380, n31381, n31385, n31387, n31389, n31390, n31393, 
      n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402, 
      n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411, 
      n31414, n31415, n31416, n31417, n31418, n31419, n31421, n31422, n31423, 
      n31424, n31426, n31427, n31428, n31429, n31432, n31434, n31435, n31437, 
      n31438, n31440, n31442, n31443, n31444, n31445, n31448, n31450, n31451, 
      n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31461, n31463, 
      n31464, n31467, n31468, n31469, n31470, n31471, n31473, n31474, n31475, 
      n31476, n31477, n31478, n31479, n31483, n31484, n31485, n31486, n31487, 
      n31488, n31489, n31490, n31491, n31492, n31493, n31495, n31496, n31497, 
      n31498, n31499, n31500, n31503, n31504, n31505, n31506, n31507, n31508, 
      n31509, n31510, n31511, n31512, n31513, n31514, n31516, n31519, n31521, 
      n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31531, 
      n31532, n31533, n31534, n31538, n31539, n31542, n31543, n31544, n31545, 
      n31547, n31548, n31549, n31551, n31552, n31553, n31554, n31557, n31559, 
      n31560, n31561, n31562, n31563, n31564, n31566, n31567, n31568, n31569, 
      n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31579, n31583, 
      n31584, n31585, n31588, n31590, n31591, n31593, n31594, n31596, n31597, 
      n31598, n31599, n31601, n31602, n31603, n31604, n31606, n31607, n31608, 
      n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619, 
      n31622, n31623, n31626, n31627, n31629, n31630, n31634, n31635, n31636, 
      n31637, n31638, n31639, n31640, n31642, n31643, n31644, n31645, n31646, 
      n31647, n31649, n31650, n31653, n31654, n31655, n31656, n31657, n31658, 
      n31660, n31661, n31662, n31663, n31664, n31666, n31667, n31668, n31669, 
      n31670, n31671, n31673, n31674, n31675, n31676, n31677, n31678, n31679, 
      n31682, n31683, n31684, n31686, n31687, n31689, n31690, n31691, n31692, 
      n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31701, n31702, 
      n31703, n31704, n31706, n31707, n31709, n31710, n31711, n31712, n31713, 
      n31714, n31715, n31716, n31718, n31719, n31720, n31721, n31722, n31724, 
      n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31734, 
      n31736, n31737, n31738, n31739, n31742, n31745, n31746, n31747, n31748, 
      n31749, n31750, n31751, n31753, n31754, n31755, n31756, n31757, n31758, 
      n31759, n31760, n31761, n31762, n31763, n31765, n31766, n31767, n31768, 
      n31769, n31770, n31771, n31772, n31773, n31776, n31777, n31778, n31779, 
      n31780, n31781, n31783, n31784, n31785, n31786, n31787, n31788, n31790, 
      n31793, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31803, 
      n31804, n31805, n31807, n31810, n31811, n31813, n31814, n31815, n31819, 
      n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, 
      n31830, n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31841, 
      n31843, n31844, n31848, n31849, n31850, n31852, n31853, n31854, n31856, 
      n31857, n31859, n31860, n31861, n31862, n31863, n31866, n31867, n31868, 
      n31869, n31871, n31872, n31873, n31874, n31875, n31876, n31878, n31880, 
      n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890, 
      n31891, n31892, n31893, n31894, n31895, n31898, n31899, n31900, n31901, 
      n31902, n31903, n31904, n31906, n31907, n31908, n31909, n31910, n31911, 
      n31912, n31913, n31914, n31915, n31916, n31918, n31919, n31920, n31921, 
      n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, 
      n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, 
      n31940, n31941, n31942, n31943, n31945, n31946, n31947, n31948, n31949, 
      n31950, n31951, n31953, n31954, n31956, n31957, n31958, n31959, n31960, 
      n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969, 
      n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978, 
      n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987, 
      n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996, 
      n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005, 
      n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014, 
      n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023, 
      n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032, 
      n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041, 
      n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050, 
      n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059, 
      n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068, 
      n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077, 
      n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, 
      n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, 
      n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, 
      n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, 
      n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122, 
      n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131, 
      n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140, 
      n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149, 
      n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158, 
      n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167, 
      n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176, 
      n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185, 
      n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194, 
      n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203, 
      n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212, 
      n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221, 
      n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230, 
      n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239, 
      n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248, 
      n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257, 
      n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266, 
      n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275, 
      n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284, 
      n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293, 
      n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302, 
      n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311, 
      n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320, 
      n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329, 
      n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338, 
      n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347, 
      n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356, 
      n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365, 
      n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374, 
      n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383, 
      n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392, 
      n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401, 
      n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410, 
      n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419, 
      n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428, 
      n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437, 
      n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446, 
      n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455, 
      n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, 
      n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, 
      n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, 
      n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, 
      n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500, 
      n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509, 
      n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518, 
      n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527, 
      n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536, 
      n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545, 
      n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554, 
      n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563, 
      n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572, 
      n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581, 
      n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590, 
      n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599, 
      n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608, 
      n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617, 
      n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626, 
      n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635, 
      n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644, 
      n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653, 
      n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662, 
      n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671, 
      n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680, 
      n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689, 
      n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698, 
      n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707, 
      n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716, 
      n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725, 
      n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734, 
      n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743, 
      n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752, 
      n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761, 
      n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770, 
      n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779, 
      n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788, 
      n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797, 
      n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806, 
      n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815, 
      n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824, 
      n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833, 
      n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842, 
      n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851, 
      n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860, 
      n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869, 
      n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878, 
      n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887, 
      n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896, 
      n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905, 
      n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914, 
      n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923, 
      n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932, 
      n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941, 
      n32942, n32943, n32945, n32946, n32947, n32948, n32949, n32950, n32951, 
      n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960, 
      n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969, 
      n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978, 
      n32979, n32980, n32981, n32983, n32984, n32985, n32986, n32987, n32988, 
      n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997, 
      n32998, n32999, n33001, n33002, n33003, n33004, n33005, n33006, n33007, 
      n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016, 
      n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025, 
      n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034, 
      n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043, 
      n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052, 
      n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061, 
      n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070, 
      n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079, 
      n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088, 
      n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097, 
      n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, 
      n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115, 
      n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124, 
      n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133, 
      n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142, 
      n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151, 
      n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160, 
      n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169, 
      n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178, 
      n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187, 
      n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196, 
      n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205, 
      n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214, 
      n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223, 
      n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232, 
      n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241, 
      n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250, 
      n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259, 
      n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268, 
      n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277, 
      n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286, 
      n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295, 
      n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304, 
      n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313, 
      n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322, 
      n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331, 
      n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340, 
      n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349, 
      n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358, 
      n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367, 
      n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376, 
      n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385, 
      n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, 
      n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403, 
      n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412, 
      n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, 
      n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430, 
      n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439, 
      n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448, 
      n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457, 
      n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466, 
      n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475, 
      n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484, 
      n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493, 
      n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502, 
      n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511, 
      n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520, 
      n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529, 
      n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, 
      n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547, 
      n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556, 
      n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565, 
      n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574, 
      n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583, 
      n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33593, 
      n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602, 
      n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611, 
      n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620, 
      n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629, 
      n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638, 
      n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647, 
      n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656, 
      n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665, 
      n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674, 
      n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683, 
      n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692, 
      n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701, 
      n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710, 
      n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719, 
      n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728, 
      n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737, 
      n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746, 
      n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755, 
      n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764, 
      n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773, 
      n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782, 
      n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791, 
      n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800, 
      n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809, 
      n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818, 
      n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827, 
      n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836, 
      n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845, 
      n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854, 
      n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863, 
      n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872, 
      n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881, 
      n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890, 
      n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899, 
      n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908, 
      n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917, 
      n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926, 
      n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935, 
      n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944, 
      n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953, 
      n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962, 
      n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971, 
      n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980, 
      n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989, 
      n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998, 
      n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007, 
      n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016, 
      n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025, 
      n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034, 
      n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043, 
      n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052, 
      n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061, 
      n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070, 
      n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079, 
      n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088, 
      n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097, 
      n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106, 
      n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115, 
      n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124, 
      n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132, n34133, 
      n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142, 
      n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151, 
      n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160, 
      n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169, 
      n34170 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n5901, A2 => n964, ZN => n433);
   U10 : NOR2_X1 port map( A1 => n17637, A2 => n25517, ZN => n25509);
   U35 : NAND3_X1 port map( A1 => n24584, A2 => n24583, A3 => n24582, ZN => 
                           n10608);
   U39 : NAND2_X1 port map( A1 => n10174, A2 => n32856, ZN => n10173);
   U130 : INV_X1 port map( I => n13236, ZN => n24592);
   U138 : INV_X1 port map( I => n5284, ZN => n24782);
   U145 : NAND2_X1 port map( A1 => n2444, A2 => n23618, ZN => n214);
   U192 : NOR2_X1 port map( A1 => n24271, A2 => n29307, ZN => n2923);
   U251 : NAND2_X1 port map( A1 => n16676, A2 => n13549, ZN => n7504);
   U278 : INV_X2 port map( I => n33722, ZN => n16786);
   U313 : INV_X1 port map( I => n23450, ZN => n169);
   U317 : INV_X1 port map( I => n24386, ZN => n12797);
   U320 : INV_X1 port map( I => n23534, ZN => n23227);
   U325 : INV_X1 port map( I => n16703, ZN => n18122);
   U330 : INV_X1 port map( I => n29885, ZN => n8883);
   U371 : INV_X1 port map( I => n13679, ZN => n13751);
   U390 : INV_X1 port map( I => n12729, ZN => n11308);
   U429 : INV_X2 port map( I => n2860, ZN => n1106);
   U438 : NAND2_X1 port map( A1 => n11250, A2 => n29287, ZN => n22685);
   U442 : AOI21_X1 port map( A1 => n22672, A2 => n29304, B => n9753, ZN => 
                           n22673);
   U447 : INV_X1 port map( I => n17151, ZN => n22577);
   U452 : OR2_X1 port map( A1 => n639, A2 => n9953, Z => n22682);
   U487 : NAND2_X1 port map( A1 => n22562, A2 => n22403, ZN => n6384);
   U489 : INV_X1 port map( I => n22679, ZN => n22562);
   U512 : INV_X1 port map( I => n21958, ZN => n1306);
   U554 : OR2_X1 port map( A1 => n31511, A2 => n21651, Z => n21641);
   U577 : INV_X1 port map( I => n21708, ZN => n9119);
   U586 : NAND2_X1 port map( A1 => n21491, A2 => n21568, ZN => n21492);
   U680 : NOR2_X1 port map( A1 => n21374, A2 => n4145, ZN => n15814);
   U695 : INV_X2 port map( I => n21203, ZN => n21400);
   U738 : OAI21_X1 port map( A1 => n27177, A2 => n1034, B => n3787, ZN => n3558
                           );
   U752 : NAND3_X1 port map( A1 => n20591, A2 => n20589, A3 => n384, ZN => 
                           n20173);
   U760 : CLKBUF_X2 port map( I => n15230, Z => n8353);
   U780 : INV_X2 port map( I => n17544, ZN => n20486);
   U802 : OAI21_X1 port map( A1 => n11909, A2 => n16065, B => n6644, ZN => 
                           n10056);
   U804 : NAND2_X1 port map( A1 => n1826, A2 => n402, ZN => n9015);
   U815 : NOR2_X1 port map( A1 => n10086, A2 => n6200, ZN => n402);
   U818 : NAND3_X1 port map( A1 => n25997, A2 => n16, A3 => n13747, ZN => 
                           n15435);
   U876 : INV_X2 port map( I => n28951, ZN => n1044);
   U882 : INV_X1 port map( I => n25208, ZN => n293);
   U884 : INV_X1 port map( I => n15960, ZN => n876);
   U891 : INV_X1 port map( I => n2581, ZN => n18840);
   U954 : INV_X2 port map( I => n9319, ZN => n7687);
   U958 : INV_X1 port map( I => n6846, ZN => n18913);
   U963 : NAND2_X1 port map( A1 => n7900, A2 => n30744, ZN => n436);
   U970 : INV_X1 port map( I => n31971, ZN => n952);
   U994 : NAND2_X1 port map( A1 => n18515, A2 => n13663, ZN => n16086);
   U1011 : INV_X1 port map( I => n18700, ZN => n18007);
   U1014 : INV_X2 port map( I => n494, ZN => n1188);
   U1027 : NAND2_X2 port map( A1 => n34037, A2 => n1333, ZN => n1915);
   U1061 : NOR2_X2 port map( A1 => n21715, A2 => n21601, ZN => n21710);
   U1070 : NAND2_X2 port map( A1 => n29185, A2 => n23721, ZN => n13342);
   U1088 : INV_X2 port map( I => n18018, ZN => n18616);
   U1102 : NAND2_X2 port map( A1 => n14246, A2 => n27182, ZN => n25404);
   U1162 : INV_X2 port map( I => n13442, ZN => n13816);
   U1167 : NOR2_X2 port map( A1 => n20361, A2 => n27887, ZN => n20451);
   U1178 : NOR2_X2 port map( A1 => n25891, A2 => n25890, ZN => n9941);
   U1299 : INV_X2 port map( I => n10335, ZN => n17456);
   U1317 : NOR2_X2 port map( A1 => n3455, A2 => n9800, ZN => n3124);
   U1353 : OAI22_X2 port map( A1 => n1143, A2 => n21237, B1 => n424, B2 => n780
                           , ZN => n12836);
   U1384 : INV_X2 port map( I => n16748, ZN => n14198);
   U1415 : INV_X4 port map( I => n4656, ZN => n19301);
   U1424 : AOI22_X2 port map( A1 => n3189, A2 => n1720, B1 => n3188, B2 => 
                           n1120, ZN => n3187);
   U1440 : NAND2_X2 port map( A1 => n1384, A2 => n18990, ZN => n19091);
   U1452 : NAND2_X2 port map( A1 => n7600, A2 => n19255, ZN => n2177);
   U1465 : INV_X2 port map( I => n17352, ZN => n23904);
   U1470 : INV_X2 port map( I => n18674, ZN => n18881);
   U1482 : BUF_X2 port map( I => n22535, Z => n16434);
   U1517 : INV_X2 port map( I => n18990, ZN => n878);
   U1528 : BUF_X4 port map( I => n16801, Z => n10828);
   U1536 : NAND2_X2 port map( A1 => n8787, A2 => n19115, ZN => n19186);
   U1543 : BUF_X2 port map( I => n29781, Z => n2582);
   U1548 : AOI21_X2 port map( A1 => n18347, A2 => n18346, B => n18345, ZN => 
                           n2331);
   U1557 : NOR2_X1 port map( A1 => n25971, A2 => n16740, ZN => n16876);
   U1559 : NAND3_X1 port map( A1 => n1358, A2 => n13327, A3 => n19949, ZN => 
                           n20191);
   U1569 : OAI21_X1 port map( A1 => n31407, A2 => n1074, B => n694, ZN => n66);
   U1571 : NAND2_X1 port map( A1 => n14764, A2 => n712, ZN => n14763);
   U1616 : INV_X1 port map( I => n5492, ZN => n5113);
   U1624 : NOR2_X1 port map( A1 => n33563, A2 => n268, ZN => n17336);
   U1625 : INV_X2 port map( I => n11984, ZN => n13499);
   U1630 : NAND2_X2 port map( A1 => n14311, A2 => n11831, ZN => n24548);
   U1648 : NAND2_X1 port map( A1 => n16800, A2 => n29866, ZN => n363);
   U1651 : NAND3_X1 port map( A1 => n4770, A2 => n786, A3 => n4782, ZN => n3433
                           );
   U1678 : AOI21_X1 port map( A1 => n21669, A2 => n21672, B => n16345, ZN => 
                           n21278);
   U1685 : NAND2_X1 port map( A1 => n22919, A2 => n8365, ZN => n268);
   U1727 : INV_X2 port map( I => n19641, ZN => n1045);
   U1736 : NAND2_X1 port map( A1 => n3722, A2 => n3723, ZN => n15796);
   U1749 : OR2_X2 port map( A1 => n5392, A2 => n11847, Z => n21202);
   U1766 : INV_X1 port map( I => n18310, ZN => n1184);
   U1771 : NAND2_X2 port map( A1 => n17334, A2 => n17335, ZN => n23346);
   U1779 : OAI21_X2 port map( A1 => n827, A2 => n29, B => n19050, ZN => n13448)
                           ;
   U1788 : XOR2_X1 port map( A1 => n2278, A2 => n31259, Z => n12011);
   U1806 : NOR2_X2 port map( A1 => n12074, A2 => n16766, ZN => n14284);
   U1807 : NAND2_X1 port map( A1 => n24138, A2 => n16286, ZN => n6980);
   U1810 : INV_X2 port map( I => n9436, ZN => n11372);
   U1820 : NAND2_X1 port map( A1 => n9695, A2 => n9697, ZN => n13065);
   U1821 : NOR2_X1 port map( A1 => n27123, A2 => n10858, ZN => n9696);
   U1830 : INV_X2 port map( I => n12241, ZN => n13852);
   U1836 : NAND2_X2 port map( A1 => n11, A2 => n4209, ZN => n20468);
   U1844 : BUF_X2 port map( I => n24117, Z => n13);
   U1849 : INV_X2 port map( I => n5837, ZN => n17495);
   U1876 : AOI21_X2 port map( A1 => n17371, A2 => n28219, B => n15366, ZN => 
                           n9099);
   U1877 : INV_X1 port map( I => n25985, ZN => n8450);
   U1890 : XOR2_X1 port map( A1 => n18948, A2 => n17613, Z => n367);
   U1898 : BUF_X2 port map( I => n18700, Z => n22);
   U1901 : XOR2_X1 port map( A1 => n24837, A2 => n16504, Z => n13849);
   U1908 : AOI21_X2 port map( A1 => n15585, A2 => n17234, B => n14778, ZN => 
                           n15584);
   U1913 : AOI21_X2 port map( A1 => n6069, A2 => n761, B => n4162, ZN => n6068)
                           ;
   U1920 : NAND2_X2 port map( A1 => n6074, A2 => n21581, ZN => n21666);
   U1923 : XOR2_X1 port map( A1 => n8861, A2 => n10328, Z => n3304);
   U1936 : AOI21_X2 port map( A1 => n22607, A2 => n9155, B => n5958, ZN => 
                           n23110);
   U1943 : AND2_X1 port map( A1 => n28338, A2 => n29279, Z => n696);
   U1954 : XOR2_X1 port map( A1 => n29277, A2 => n31, Z => n4951);
   U1955 : XOR2_X1 port map( A1 => n24538, A2 => n14079, Z => n31);
   U1957 : XOR2_X1 port map( A1 => n23473, A2 => n11667, Z => n4661);
   U1960 : XOR2_X1 port map( A1 => n7566, A2 => n34, Z => n606);
   U1961 : XOR2_X1 port map( A1 => n7565, A2 => n29413, Z => n34);
   U1982 : BUF_X2 port map( I => Key(54), Z => n16690);
   U1987 : INV_X4 port map( I => n18683, ZN => n1659);
   U1996 : XOR2_X1 port map( A1 => n29275, A2 => n44, Z => n5965);
   U1997 : XOR2_X1 port map( A1 => n24773, A2 => n24476, Z => n44);
   U2014 : NAND2_X2 port map( A1 => n18400, A2 => n46, ZN => n19294);
   U2024 : XOR2_X1 port map( A1 => n4986, A2 => n702, Z => n4984);
   U2034 : XOR2_X1 port map( A1 => n52, A2 => n14809, Z => n15733);
   U2041 : XOR2_X1 port map( A1 => n23463, A2 => n54, Z => n14783);
   U2042 : XOR2_X1 port map( A1 => n23299, A2 => n23489, Z => n54);
   U2070 : XOR2_X1 port map( A1 => n23136, A2 => n62, Z => n17591);
   U2071 : XOR2_X1 port map( A1 => n26101, A2 => n14818, Z => n62);
   U2076 : NAND2_X2 port map( A1 => n2677, A2 => n16084, ZN => n20529);
   U2082 : NAND2_X2 port map( A1 => n16669, A2 => n31324, ZN => n17239);
   U2101 : NAND2_X1 port map( A1 => n18462, A2 => n18463, ZN => n94);
   U2102 : AOI21_X2 port map( A1 => n4879, A2 => n4643, B => n8091, ZN => n4878
                           );
   U2116 : INV_X2 port map( I => n11562, ZN => n22139);
   U2150 : NAND2_X2 port map( A1 => n28904, A2 => n3157, ZN => n20334);
   U2151 : XOR2_X1 port map( A1 => n81, A2 => n23132, Z => n23263);
   U2157 : NAND2_X2 port map( A1 => n21559, A2 => n6489, ZN => n21821);
   U2162 : XOR2_X1 port map( A1 => n10399, A2 => n6571, Z => n86);
   U2165 : INV_X2 port map( I => n87, ZN => n563);
   U2168 : INV_X2 port map( I => n14980, ZN => n13759);
   U2179 : OR2_X1 port map( A1 => n14212, A2 => n28891, Z => n4611);
   U2185 : NAND2_X1 port map( A1 => n11419, A2 => n15835, ZN => n92);
   U2211 : NAND2_X1 port map( A1 => n33583, A2 => n31807, ZN => n97);
   U2243 : OAI21_X1 port map( A1 => n25278, A2 => n12431, B => n25284, ZN => 
                           n16290);
   U2247 : INV_X4 port map( I => n4746, ZN => n15179);
   U2251 : INV_X2 port map( I => n11833, ZN => n22926);
   U2252 : NAND2_X1 port map( A1 => n107, A2 => n16347, ZN => n25255);
   U2265 : OAI21_X2 port map( A1 => n21298, A2 => n15807, B => n21299, ZN => 
                           n21721);
   U2292 : BUF_X4 port map( I => n9125, Z => n9127);
   U2294 : NAND2_X2 port map( A1 => n7144, A2 => n17888, ZN => n21877);
   U2302 : XOR2_X1 port map( A1 => n20746, A2 => n3209, Z => n11689);
   U2308 : XOR2_X1 port map( A1 => n16917, A2 => n6973, Z => n119);
   U2330 : AOI21_X2 port map( A1 => n11709, A2 => n9854, B => n124, ZN => 
                           n20727);
   U2341 : XOR2_X1 port map( A1 => n34160, A2 => n22072, Z => n22307);
   U2343 : XOR2_X1 port map( A1 => n19554, A2 => n26032, Z => n128);
   U2348 : NOR2_X1 port map( A1 => n4953, A2 => n17927, ZN => n4952);
   U2367 : OAI21_X1 port map( A1 => n25526, A2 => n15295, B => n15155, ZN => 
                           n25527);
   U2377 : INV_X2 port map( I => n10371, ZN => n8778);
   U2379 : NOR2_X2 port map( A1 => n1352, A2 => n14545, ZN => n10323);
   U2381 : XOR2_X1 port map( A1 => n15353, A2 => n136, Z => n10558);
   U2382 : XOR2_X1 port map( A1 => n15352, A2 => n20962, Z => n136);
   U2386 : OAI21_X1 port map( A1 => n25488, A2 => n25487, B => n25486, ZN => 
                           n138);
   U2388 : XOR2_X1 port map( A1 => n16693, A2 => n25190, Z => n139);
   U2390 : NAND2_X2 port map( A1 => n7278, A2 => n7277, ZN => n12491);
   U2394 : INV_X2 port map( I => n23949, ZN => n23947);
   U2407 : INV_X2 port map( I => n3340, ZN => n19236);
   U2419 : INV_X2 port map( I => n4113, ZN => n18241);
   U2426 : OAI22_X1 port map( A1 => n25668, A2 => n9365, B1 => n25645, B2 => 
                           n25651, ZN => n25642);
   U2432 : INV_X2 port map( I => n18884, ZN => n18662);
   U2436 : BUF_X4 port map( I => n14702, Z => n1337);
   U2438 : INV_X2 port map( I => n10146, ZN => n24811);
   U2449 : NOR2_X2 port map( A1 => n11759, A2 => n152, ZN => n17927);
   U2456 : XOR2_X1 port map( A1 => n153, A2 => n25195, Z => Ciphertext(71));
   U2457 : NAND3_X1 port map( A1 => n4767, A2 => n4768, A3 => n4769, ZN => n153
                           );
   U2459 : INV_X2 port map( I => n12811, ZN => n12992);
   U2462 : NAND2_X2 port map( A1 => n7492, A2 => n5455, ZN => n11074);
   U2488 : NAND2_X2 port map( A1 => n4337, A2 => n28701, ZN => n20940);
   U2491 : OAI21_X2 port map( A1 => n16712, A2 => n10778, B => n28240, ZN => 
                           n10777);
   U2497 : XOR2_X1 port map( A1 => n21035, A2 => n1993, Z => n11424);
   U2498 : NAND2_X2 port map( A1 => n11617, A2 => n11618, ZN => n21035);
   U2503 : NAND2_X2 port map( A1 => n21812, A2 => n18184, ZN => n11848);
   U2511 : OR2_X2 port map( A1 => n1850, A2 => n28591, Z => n12247);
   U2523 : XOR2_X1 port map( A1 => n1454, A2 => n168, Z => n652);
   U2524 : XOR2_X1 port map( A1 => n23199, A2 => n169, Z => n168);
   U2528 : XOR2_X1 port map( A1 => n170, A2 => n29108, Z => n17535);
   U2529 : XOR2_X1 port map( A1 => n6417, A2 => n15334, Z => n170);
   U2538 : XOR2_X1 port map( A1 => n175, A2 => n12062, Z => n18037);
   U2540 : NAND2_X2 port map( A1 => n15166, A2 => n15165, ZN => n18997);
   U2553 : XOR2_X1 port map( A1 => n3504, A2 => n5051, Z => n24549);
   U2558 : XOR2_X1 port map( A1 => n5231, A2 => n5229, Z => n25112);
   U2564 : AOI22_X2 port map( A1 => n11815, A2 => n18556, B1 => n16564, B2 => 
                           n18328, ZN => n5892);
   U2565 : NAND3_X2 port map( A1 => n5890, A2 => n5892, A3 => n5891, ZN => 
                           n5545);
   U2575 : OR2_X1 port map( A1 => n21733, A2 => n13872, Z => n187);
   U2579 : INV_X2 port map( I => n10327, ZN => n17814);
   U2594 : INV_X2 port map( I => n193, ZN => n502);
   U2595 : XOR2_X1 port map( A1 => n5151, A2 => n5152, Z => n193);
   U2596 : INV_X2 port map( I => n29814, ZN => n1353);
   U2627 : INV_X2 port map( I => n3967, ZN => n19907);
   U2631 : XOR2_X1 port map( A1 => n21990, A2 => n29259, Z => n13704);
   U2632 : OAI21_X2 port map( A1 => n6117, A2 => n15697, B => n6116, ZN => 
                           n7134);
   U2634 : XOR2_X1 port map( A1 => n7674, A2 => n26085, Z => n15309);
   U2651 : XOR2_X1 port map( A1 => n2330, A2 => n19467, Z => n2335);
   U2653 : NAND3_X1 port map( A1 => n20361, A2 => n27887, A3 => n10939, ZN => 
                           n5349);
   U2659 : INV_X4 port map( I => n17408, ZN => n22705);
   U2661 : OR2_X1 port map( A1 => n9719, A2 => n20375, Z => n204);
   U2672 : NAND2_X1 port map( A1 => n2209, A2 => n6288, ZN => n13023);
   U2674 : INV_X2 port map( I => n625, ZN => n5440);
   U2709 : OAI21_X2 port map( A1 => n18956, A2 => n784, B => n13009, ZN => 
                           n13482);
   U2717 : XOR2_X1 port map( A1 => n23254, A2 => n22841, Z => n225);
   U2726 : XOR2_X1 port map( A1 => n29194, A2 => n6923, Z => n227);
   U2734 : XOR2_X1 port map( A1 => n22230, A2 => n233, Z => n17284);
   U2735 : XOR2_X1 port map( A1 => n32084, A2 => n22092, Z => n233);
   U2751 : NAND2_X2 port map( A1 => n19283, A2 => n19285, ZN => n19080);
   U2756 : NOR2_X2 port map( A1 => n1864, A2 => n6073, ZN => n10717);
   U2786 : INV_X4 port map( I => n5610, ZN => n1378);
   U2827 : INV_X2 port map( I => n23143, ZN => n23211);
   U2856 : NAND2_X1 port map( A1 => n20573, A2 => n20572, ZN => n258);
   U2859 : AOI21_X1 port map( A1 => n7680, A2 => n16274, B => n259, ZN => 
                           n19250);
   U2868 : XOR2_X1 port map( A1 => n30443, A2 => n19494, Z => n19431);
   U2869 : OAI21_X2 port map( A1 => n1451, A2 => n1453, B => n1450, ZN => 
                           n19494);
   U2872 : NAND2_X2 port map( A1 => n9967, A2 => n11452, ZN => n21651);
   U2885 : NAND2_X1 port map( A1 => n5948, A2 => n12654, ZN => n262);
   U2896 : OAI21_X2 port map( A1 => n22774, A2 => n15718, B => n22759, ZN => 
                           n7625);
   U2901 : XOR2_X1 port map( A1 => Plaintext(70), A2 => Key(70), Z => n270);
   U2917 : XOR2_X1 port map( A1 => n12011, A2 => n24441, Z => n16877);
   U2918 : XOR2_X1 port map( A1 => n24475, A2 => n9386, Z => n24441);
   U2924 : NAND3_X2 port map( A1 => n273, A2 => n2922, A3 => n23991, ZN => 
                           n24664);
   U2926 : INV_X2 port map( I => n2236, ZN => n694);
   U2929 : XOR2_X1 port map( A1 => n24596, A2 => n24576, Z => n17097);
   U2936 : INV_X2 port map( I => n23904, ZN => n11050);
   U2958 : XOR2_X1 port map( A1 => n6706, A2 => n15761, Z => n281);
   U2970 : XOR2_X1 port map( A1 => n9644, A2 => n13888, Z => n16030);
   U2983 : INV_X2 port map( I => n292, ZN => n547);
   U2986 : XOR2_X1 port map( A1 => n16429, A2 => n293, Z => n476);
   U2992 : NAND2_X2 port map( A1 => n11961, A2 => n294, ZN => n19951);
   U2993 : INV_X4 port map( I => n16681, ZN => n2694);
   U3004 : NOR2_X2 port map( A1 => n14659, A2 => n14658, ZN => n14657);
   U3008 : XOR2_X1 port map( A1 => n7387, A2 => n13863, Z => n17126);
   U3009 : NAND2_X2 port map( A1 => n13478, A2 => n13479, ZN => n7387);
   U3029 : INV_X2 port map( I => n15057, ZN => n16009);
   U3032 : INV_X4 port map( I => n17598, ZN => n18761);
   U3044 : AND2_X1 port map( A1 => n24138, A2 => n24141, Z => n11832);
   U3050 : XOR2_X1 port map( A1 => n5381, A2 => n30319, Z => n23313);
   U3052 : XOR2_X1 port map( A1 => n308, A2 => n19539, Z => n7193);
   U3053 : XOR2_X1 port map( A1 => n31568, A2 => n16301, Z => n308);
   U3065 : INV_X4 port map( I => n21056, ZN => n9191);
   U3079 : NAND2_X2 port map( A1 => n5969, A2 => n5968, ZN => n5970);
   U3082 : NAND2_X2 port map( A1 => n10513, A2 => n24207, ZN => n24062);
   U3100 : BUF_X2 port map( I => n24852, Z => n322);
   U3105 : NOR2_X2 port map( A1 => n14951, A2 => n16844, ZN => n13800);
   U3117 : XOR2_X1 port map( A1 => n15093, A2 => n15934, Z => n16778);
   U3118 : XOR2_X1 port map( A1 => n22114, A2 => n29851, Z => n3101);
   U3127 : BUF_X4 port map( I => n13531, Z => n13548);
   U3135 : NAND2_X1 port map( A1 => n8305, A2 => n5595, ZN => n329);
   U3138 : NAND2_X2 port map( A1 => n10615, A2 => n10614, ZN => n20412);
   U3141 : INV_X2 port map( I => n25228, ZN => n25306);
   U3144 : NOR2_X2 port map( A1 => n24036, A2 => n24035, ZN => n24796);
   U3161 : OR2_X1 port map( A1 => n11827, A2 => n11826, Z => n337);
   U3178 : INV_X2 port map( I => n25711, ZN => n1077);
   U3183 : XOR2_X1 port map( A1 => n19626, A2 => n4942, Z => n19577);
   U3189 : XOR2_X1 port map( A1 => n22235, A2 => n22152, Z => n2696);
   U3190 : XOR2_X1 port map( A1 => n16210, A2 => n22017, Z => n22235);
   U3192 : OAI22_X1 port map( A1 => n18777, A2 => n28686, B1 => n954, B2 => 
                           n16585, ZN => n12877);
   U3200 : INV_X1 port map( I => n8243, ZN => n13730);
   U3210 : NAND2_X2 port map( A1 => n2905, A2 => n15285, ZN => n20632);
   U3215 : INV_X2 port map( I => n18048, ZN => n349);
   U3233 : XOR2_X1 port map( A1 => n15630, A2 => n26075, Z => n5133);
   U3235 : NOR2_X2 port map( A1 => n6943, A2 => n642, ZN => n6874);
   U3237 : OR2_X1 port map( A1 => n28338, A2 => n11899, Z => n13819);
   U3257 : INV_X2 port map( I => n18654, ZN => n18798);
   U3264 : INV_X2 port map( I => n5441, ZN => n22585);
   U3265 : OAI21_X2 port map( A1 => n18327, A2 => n180, B => n9840, ZN => n2581
                           );
   U3274 : NAND3_X2 port map( A1 => n365, A2 => n5990, A3 => n5989, ZN => n5988
                           );
   U3280 : OAI21_X2 port map( A1 => n7330, A2 => n10460, B => n7332, ZN => 
                           n14522);
   U3283 : XOR2_X1 port map( A1 => n10809, A2 => n367, Z => n11969);
   U3294 : INV_X2 port map( I => n24204, ZN => n24061);
   U3297 : INV_X4 port map( I => n8832, ZN => n18515);
   U3304 : NOR2_X2 port map( A1 => n5121, A2 => n5122, ZN => n6846);
   U3315 : XOR2_X1 port map( A1 => n1941, A2 => n1942, Z => n7573);
   U3321 : NAND2_X2 port map( A1 => n4130, A2 => n8144, ZN => n3929);
   U3345 : XOR2_X1 port map( A1 => n15367, A2 => n26057, Z => n380);
   U3351 : INV_X2 port map( I => n627, ZN => n1284);
   U3361 : XOR2_X1 port map( A1 => n19611, A2 => n9599, Z => n2672);
   U3369 : XOR2_X1 port map( A1 => n16877, A2 => n385, Z => n2315);
   U3370 : XOR2_X1 port map( A1 => n18174, A2 => n18173, Z => n385);
   U3400 : INV_X2 port map( I => n18037, ZN => n17147);
   U3405 : NAND2_X2 port map( A1 => n25402, A2 => n25401, ZN => n25440);
   U3423 : AOI21_X2 port map( A1 => n12026, A2 => n27455, B => n6363, ZN => 
                           n12434);
   U3442 : OR2_X1 port map( A1 => n22439, A2 => n8409, Z => n17008);
   U3446 : NAND2_X2 port map( A1 => n25391, A2 => n17717, ZN => n25346);
   U3450 : NAND2_X2 port map( A1 => n3554, A2 => n3552, ZN => n4746);
   U3455 : NAND3_X1 port map( A1 => n12682, A2 => n20040, A3 => n20138, ZN => 
                           n410);
   U3463 : NAND3_X1 port map( A1 => n6072, A2 => n8409, A3 => n1125, ZN => n413
                           );
   U3467 : BUF_X2 port map( I => n26049, Z => n414);
   U3474 : XOR2_X1 port map( A1 => n10205, A2 => n10979, Z => n5847);
   U3477 : INV_X4 port map( I => n18720, ZN => n18855);
   U3481 : OR2_X1 port map( A1 => n25366, A2 => n30400, Z => n25371);
   U3483 : XOR2_X1 port map( A1 => n3493, A2 => n416, Z => n17932);
   U3508 : INV_X2 port map( I => n4798, ZN => n424);
   U3509 : XOR2_X1 port map( A1 => n17384, A2 => n425, Z => n5340);
   U3510 : XOR2_X1 port map( A1 => n30327, A2 => n24516, Z => n425);
   U3514 : XOR2_X1 port map( A1 => n22311, A2 => n22233, Z => n9432);
   U3515 : XOR2_X1 port map( A1 => n27130, A2 => n2863, Z => n22311);
   U3518 : XOR2_X1 port map( A1 => n19585, A2 => n10434, Z => n2064);
   U3526 : XOR2_X1 port map( A1 => n5244, A2 => n30311, Z => n3584);
   U3551 : AOI21_X2 port map( A1 => n19889, A2 => n11475, B => n19949, ZN => 
                           n7245);
   U3563 : XOR2_X1 port map( A1 => n439, A2 => n16381, Z => Ciphertext(7));
   U3569 : INV_X2 port map( I => n12906, ZN => n17373);
   U3570 : XOR2_X1 port map( A1 => n12962, A2 => n440, Z => n12960);
   U3571 : XOR2_X1 port map( A1 => n11784, A2 => n26100, Z => n440);
   U3583 : OR2_X1 port map( A1 => n20376, A2 => n20361, Z => n5351);
   U3593 : INV_X1 port map( I => n22677, ZN => n22403);
   U3624 : XNOR2_X1 port map( A1 => n19540, A2 => n1364, ZN => n444);
   U3625 : XNOR2_X1 port map( A1 => n19539, A2 => n16578, ZN => n445);
   U3628 : XNOR2_X1 port map( A1 => n20730, A2 => n25735, ZN => n447);
   U3633 : XNOR2_X1 port map( A1 => n30532, A2 => n16696, ZN => n452);
   U3635 : XNOR2_X1 port map( A1 => n34150, A2 => n16698, ZN => n454);
   U3637 : XNOR2_X1 port map( A1 => n19473, A2 => n25195, ZN => n456);
   U3638 : XNOR2_X1 port map( A1 => n31229, A2 => n1403, ZN => n457);
   U3639 : XNOR2_X1 port map( A1 => n283, A2 => n1409, ZN => n458);
   U3642 : XNOR2_X1 port map( A1 => n19691, A2 => n25108, ZN => n461);
   U3644 : XNOR2_X1 port map( A1 => n19463, A2 => n25182, ZN => n463);
   U3646 : XNOR2_X1 port map( A1 => n23475, A2 => n23474, ZN => n465);
   U3652 : XNOR2_X1 port map( A1 => n19651, A2 => n25465, ZN => n467);
   U3660 : XNOR2_X1 port map( A1 => n14132, A2 => n16674, ZN => n474);
   U3661 : XNOR2_X1 port map( A1 => n23535, A2 => n16679, ZN => n475);
   U3662 : XNOR2_X1 port map( A1 => n15517, A2 => n25098, ZN => n477);
   U3663 : XNOR2_X1 port map( A1 => n30212, A2 => n24386, ZN => n478);
   U3665 : XNOR2_X1 port map( A1 => n10294, A2 => n1197, ZN => n480);
   U3666 : XNOR2_X1 port map( A1 => n34100, A2 => n16619, ZN => n481);
   U3670 : AND2_X2 port map( A1 => n17558, A2 => n4869, Z => n485);
   U3672 : XNOR2_X1 port map( A1 => n15236, A2 => n25319, ZN => n487);
   U3673 : XOR2_X1 port map( A1 => Plaintext(34), A2 => Key(34), Z => n488);
   U3678 : XOR2_X1 port map( A1 => Plaintext(97), A2 => Key(97), Z => n493);
   U3679 : XNOR2_X1 port map( A1 => Plaintext(115), A2 => Key(115), ZN => n494)
                           ;
   U3680 : XOR2_X1 port map( A1 => Plaintext(190), A2 => Key(190), Z => n495);
   U3681 : XNOR2_X1 port map( A1 => n10180, A2 => n8685, ZN => n496);
   U3683 : XOR2_X1 port map( A1 => Plaintext(96), A2 => Key(96), Z => n498);
   U3685 : XNOR2_X1 port map( A1 => n20963, A2 => n24065, ZN => n500);
   U3689 : XNOR2_X1 port map( A1 => n17010, A2 => n17009, ZN => n503);
   U3692 : XNOR2_X1 port map( A1 => n20813, A2 => n25693, ZN => n506);
   U3693 : XNOR2_X1 port map( A1 => n20921, A2 => n29707, ZN => n507);
   U3694 : XNOR2_X1 port map( A1 => n5414, A2 => n16654, ZN => n508);
   U3697 : XNOR2_X1 port map( A1 => n16634, A2 => n16448, ZN => n511);
   U3699 : XNOR2_X1 port map( A1 => n28762, A2 => n25001, ZN => n513);
   U3700 : XNOR2_X1 port map( A1 => n8269, A2 => n1427, ZN => n514);
   U3704 : XNOR2_X1 port map( A1 => n4285, A2 => n32130, ZN => n518);
   U3707 : XNOR2_X1 port map( A1 => n30309, A2 => n25506, ZN => n521);
   U3710 : XNOR2_X1 port map( A1 => n23475, A2 => n17400, ZN => n524);
   U3713 : XNOR2_X1 port map( A1 => n32050, A2 => n27176, ZN => n528);
   U3714 : XNOR2_X1 port map( A1 => n23196, A2 => n25648, ZN => n529);
   U3715 : XNOR2_X1 port map( A1 => n23200, A2 => n23291, ZN => n530);
   U3716 : XNOR2_X1 port map( A1 => n10535, A2 => n16504, ZN => n531);
   U3717 : XNOR2_X1 port map( A1 => n29217, A2 => n25716, ZN => n532);
   U3718 : XNOR2_X1 port map( A1 => n7046, A2 => n18019, ZN => n533);
   U3720 : XOR2_X1 port map( A1 => n10659, A2 => n11148, Z => n535);
   U3721 : XNOR2_X1 port map( A1 => n22056, A2 => n25457, ZN => n536);
   U3722 : XNOR2_X1 port map( A1 => n13844, A2 => n16381, ZN => n537);
   U3723 : XNOR2_X1 port map( A1 => n16160, A2 => n25001, ZN => n538);
   U3725 : INV_X1 port map( I => n23931, ZN => n23527);
   U3726 : XNOR2_X1 port map( A1 => n6262, A2 => n23295, ZN => n540);
   U3727 : XNOR2_X1 port map( A1 => n22113, A2 => n3704, ZN => n541);
   U3728 : XNOR2_X1 port map( A1 => n22113, A2 => n22173, ZN => n542);
   U3729 : XNOR2_X1 port map( A1 => n25751, A2 => n27801, ZN => n543);
   U3730 : XNOR2_X1 port map( A1 => n24738, A2 => n24632, ZN => n544);
   U3731 : XNOR2_X1 port map( A1 => n24790, A2 => n25040, ZN => n545);
   U3732 : XNOR2_X1 port map( A1 => n24787, A2 => n25493, ZN => n546);
   U3734 : XNOR2_X1 port map( A1 => n14789, A2 => n25879, ZN => n549);
   U3735 : XNOR2_X1 port map( A1 => n24816, A2 => n24895, ZN => n550);
   U3736 : XNOR2_X1 port map( A1 => n23467, A2 => n13033, ZN => n551);
   U3738 : XNOR2_X1 port map( A1 => n24545, A2 => n25104, ZN => n553);
   U3739 : XNOR2_X1 port map( A1 => n25428, A2 => n24512, ZN => n554);
   U3742 : XNOR2_X1 port map( A1 => n12821, A2 => n25578, ZN => n556);
   U3755 : XNOR2_X1 port map( A1 => n9044, A2 => n6254, ZN => n567);
   U3759 : XNOR2_X1 port map( A1 => n10663, A2 => n10661, ZN => n571);
   U3764 : XOR2_X1 port map( A1 => n7636, A2 => n7634, Z => n576);
   U3769 : BUF_X2 port map( I => n11910, Z => n11350);
   U3775 : INV_X2 port map( I => n20117, ZN => n20045);
   U3782 : XOR2_X1 port map( A1 => n32478, A2 => n16705, Z => n586);
   U3789 : XNOR2_X1 port map( A1 => n20242, A2 => n20241, ZN => n590);
   U3790 : XNOR2_X1 port map( A1 => n20873, A2 => n25878, ZN => n591);
   U3795 : XNOR2_X1 port map( A1 => n18095, A2 => n16820, ZN => n595);
   U3800 : XNOR2_X1 port map( A1 => n8827, A2 => n8826, ZN => n598);
   U3803 : INV_X2 port map( I => n8632, ZN => n21149);
   U3804 : XNOR2_X1 port map( A1 => n20699, A2 => n20698, ZN => n600);
   U3805 : XOR2_X1 port map( A1 => n1487, A2 => n2009, Z => n601);
   U3807 : XNOR2_X1 port map( A1 => n10164, A2 => n20390, ZN => n603);
   U3810 : INV_X2 port map( I => n20468, ZN => n3462);
   U3817 : NAND2_X2 port map( A1 => n4785, A2 => n4784, ZN => n21466);
   U3819 : XNOR2_X1 port map( A1 => n15268, A2 => n20644, ZN => n609);
   U3826 : NAND3_X2 port map( A1 => n1651, A2 => n1649, A3 => n1648, ZN => 
                           n22012);
   U3827 : XNOR2_X1 port map( A1 => n22145, A2 => n25167, ZN => n612);
   U3828 : XNOR2_X1 port map( A1 => n18189, A2 => n24999, ZN => n613);
   U3834 : XNOR2_X1 port map( A1 => n22047, A2 => n22013, ZN => n618);
   U3837 : XNOR2_X1 port map( A1 => n22140, A2 => n22142, ZN => n620);
   U3840 : XNOR2_X1 port map( A1 => n22029, A2 => n22021, ZN => n623);
   U3841 : XNOR2_X1 port map( A1 => n5476, A2 => n31094, ZN => n624);
   U3852 : NAND2_X2 port map( A1 => n12845, A2 => n14878, ZN => n12594);
   U3858 : NOR2_X2 port map( A1 => n14044, A2 => n14765, ZN => n22957);
   U3867 : NAND2_X2 port map( A1 => n15608, A2 => n15607, ZN => n12729);
   U3874 : XNOR2_X1 port map( A1 => n14036, A2 => n9228, ZN => n647);
   U3884 : XOR2_X1 port map( A1 => n23304, A2 => n10129, Z => n657);
   U3890 : XNOR2_X1 port map( A1 => n11551, A2 => n23468, ZN => n660);
   U3891 : XOR2_X1 port map( A1 => n11039, A2 => n23077, Z => n661);
   U3900 : NAND2_X2 port map( A1 => n9343, A2 => n23671, ZN => n9342);
   U3904 : OAI21_X2 port map( A1 => n17730, A2 => n11975, B => n13603, ZN => 
                           n24275);
   U3919 : INV_X2 port map( I => n4951, ZN => n17861);
   U3923 : INV_X4 port map( I => n25871, ZN => n883);
   U3942 : INV_X2 port map( I => n17476, ZN => n25903);
   U3944 : INV_X2 port map( I => n8044, ZN => n25892);
   U3947 : OR2_X1 port map( A1 => n25067, A2 => n1951, Z => n693);
   U3949 : OR2_X1 port map( A1 => n24922, A2 => n15799, Z => n698);
   U3965 : NAND2_X2 port map( A1 => n4420, A2 => n15350, ZN => n20450);
   U3970 : AOI21_X2 port map( A1 => n28395, A2 => n28838, B => n2551, ZN => 
                           n1771);
   U3978 : INV_X1 port map( I => n19583, ZN => n16110);
   U3988 : NAND3_X2 port map( A1 => n17511, A2 => n20490, A3 => n17513, ZN => 
                           n20726);
   U3997 : OAI21_X2 port map( A1 => n10167, A2 => n17269, B => n10166, ZN => 
                           n23053);
   U4012 : INV_X1 port map( I => n22390, ZN => n22549);
   U4021 : AOI21_X2 port map( A1 => n5473, A2 => n5053, B => n5052, ZN => 
                           n16047);
   U4034 : AOI21_X2 port map( A1 => n12634, A2 => n20135, B => n19964, ZN => 
                           n2905);
   U4039 : NAND2_X1 port map( A1 => n6288, A2 => n7842, ZN => n25679);
   U4043 : OR2_X1 port map( A1 => n24910, A2 => n10755, Z => n8304);
   U4050 : NAND2_X2 port map( A1 => n25765, A2 => n25704, ZN => n9804);
   U4051 : AOI21_X2 port map( A1 => n17475, A2 => n25904, B => n8299, ZN => 
                           n10285);
   U4074 : INV_X2 port map( I => n14142, ZN => n25563);
   U4101 : INV_X2 port map( I => n7825, ZN => n15423);
   U4109 : INV_X2 port map( I => n2200, ZN => n23201);
   U4144 : INV_X2 port map( I => n9753, ZN => n10622);
   U4146 : INV_X2 port map( I => n9750, ZN => n10568);
   U4154 : INV_X2 port map( I => n8964, ZN => n8965);
   U4179 : INV_X1 port map( I => n28429, ZN => n12278);
   U4213 : NAND2_X2 port map( A1 => n11141, A2 => n5910, ZN => n17544);
   U4214 : NAND2_X2 port map( A1 => n9099, A2 => n9098, ZN => n12563);
   U4221 : INV_X2 port map( I => n29252, ZN => n821);
   U4226 : BUF_X4 port map( I => n19455, Z => n16694);
   U4229 : INV_X2 port map( I => n12467, ZN => n20067);
   U4237 : AND2_X1 port map( A1 => n13252, A2 => n1452, Z => n1451);
   U4255 : AND2_X1 port map( A1 => n15873, A2 => n5834, Z => n15870);
   U4262 : INV_X2 port map( I => n3954, ZN => n5225);
   U4270 : CLKBUF_X2 port map( I => n18823, Z => n4868);
   U4272 : BUF_X1 port map( I => Key(133), Z => n25156);
   U4275 : BUF_X1 port map( I => Key(105), Z => n16506);
   U4286 : BUF_X1 port map( I => Key(189), Z => n24527);
   U4291 : BUF_X1 port map( I => Key(168), Z => n25086);
   U4293 : BUF_X1 port map( I => Key(161), Z => n25288);
   U4299 : BUF_X1 port map( I => Key(59), Z => n24231);
   U4304 : BUF_X1 port map( I => Key(135), Z => n24417);
   U4308 : BUF_X1 port map( I => Key(9), Z => n25570);
   U4312 : BUF_X1 port map( I => Key(165), Z => n16597);
   U4314 : BUF_X1 port map( I => Key(125), Z => n25108);
   U4315 : BUF_X1 port map( I => Key(104), Z => n24514);
   U4320 : BUF_X1 port map( I => Key(131), Z => n24426);
   U4333 : NAND3_X1 port map( A1 => n25575, A2 => n25571, A3 => n30285, ZN => 
                           n6730);
   U4339 : NAND3_X1 port map( A1 => n25916, A2 => n25915, A3 => n25925, ZN => 
                           n25917);
   U4341 : NAND2_X1 port map( A1 => n25851, A2 => n13049, ZN => n13953);
   U4344 : NAND2_X1 port map( A1 => n24904, A2 => n24915, ZN => n3820);
   U4347 : AOI21_X1 port map( A1 => n15054, A2 => n25258, B => n2191, ZN => 
                           n25246);
   U4359 : INV_X1 port map( I => n25687, ZN => n7843);
   U4361 : INV_X1 port map( I => n3229, ZN => n3230);
   U4363 : NAND3_X1 port map( A1 => n27113, A2 => n5926, A3 => n25571, ZN => 
                           n25573);
   U4366 : NAND2_X1 port map( A1 => n31178, A2 => n25313, ZN => n25314);
   U4384 : AOI22_X1 port map( A1 => n700, A2 => n14104, B1 => n10136, B2 => 
                           n25900, ZN => n17195);
   U4398 : NAND2_X1 port map( A1 => n12856, A2 => n25591, ZN => n1751);
   U4404 : NAND2_X1 port map( A1 => n24725, A2 => n25871, ZN => n9110);
   U4408 : OAI21_X1 port map( A1 => n12359, A2 => n12358, B => n3828, ZN => 
                           n5763);
   U4411 : AND2_X1 port map( A1 => n18219, A2 => n10062, Z => n10221);
   U4431 : NAND2_X1 port map( A1 => n28096, A2 => n15295, ZN => n9718);
   U4445 : INV_X1 port map( I => n25111, ZN => n9506);
   U4463 : NAND4_X1 port map( A1 => n1816, A2 => n1818, A3 => n1819, A4 => 
                           n23594, ZN => n7962);
   U4486 : NAND2_X1 port map( A1 => n23581, A2 => n29068, ZN => n23582);
   U4499 : NAND3_X2 port map( A1 => n22410, A2 => n9747, A3 => n17481, ZN => 
                           n6386);
   U4532 : NAND2_X1 port map( A1 => n22550, A2 => n22551, ZN => n6366);
   U4536 : NAND2_X1 port map( A1 => n22025, A2 => n628, ZN => n11378);
   U4538 : INV_X2 port map( I => n8167, ZN => n9737);
   U4542 : INV_X2 port map( I => n16136, ZN => n996);
   U4551 : NOR3_X1 port map( A1 => n14949, A2 => n11755, A3 => n11229, ZN => 
                           n11228);
   U4552 : AND2_X1 port map( A1 => n11755, A2 => n6442, Z => n21676);
   U4562 : NAND2_X2 port map( A1 => n6014, A2 => n6013, ZN => n16077);
   U4572 : NOR2_X1 port map( A1 => n5822, A2 => n16633, ZN => n21311);
   U4578 : NAND3_X1 port map( A1 => n14682, A2 => n10523, A3 => n20173, ZN => 
                           n2647);
   U4580 : NOR2_X1 port map( A1 => n20547, A2 => n30130, ZN => n1961);
   U4585 : NOR2_X1 port map( A1 => n20548, A2 => n710, ZN => n6134);
   U4591 : NAND2_X1 port map( A1 => n1964, A2 => n26182, ZN => n1963);
   U4595 : INV_X1 port map( I => n20503, ZN => n16146);
   U4611 : INV_X2 port map( I => n8373, ZN => n8857);
   U4612 : INV_X2 port map( I => n11507, ZN => n14761);
   U4615 : INV_X1 port map( I => n7575, ZN => n7008);
   U4643 : INV_X2 port map( I => n15216, ZN => n18307);
   U4646 : INV_X2 port map( I => n6265, ZN => n15216);
   U4648 : BUF_X1 port map( I => Key(103), Z => n16701);
   U4659 : NAND3_X1 port map( A1 => n1208, A2 => n24969, A3 => n24970, ZN => 
                           n1934);
   U4664 : NAND2_X1 port map( A1 => n10755, A2 => n24910, ZN => n9991);
   U4670 : INV_X1 port map( I => n3843, ZN => n12783);
   U4677 : INV_X1 port map( I => n32855, ZN => n25613);
   U4681 : INV_X1 port map( I => n27173, ZN => n2049);
   U4700 : NAND2_X1 port map( A1 => n14267, A2 => n25890, ZN => n12678);
   U4704 : NAND2_X1 port map( A1 => n25233, A2 => n25232, ZN => n17925);
   U4720 : NOR2_X1 port map( A1 => n17535, A2 => n31920, ZN => n4491);
   U4726 : AOI21_X1 port map( A1 => n25229, A2 => n25306, B => n18059, ZN => 
                           n9428);
   U4732 : INV_X1 port map( I => n2378, ZN => n25526);
   U4736 : INV_X2 port map( I => n686, ZN => n13763);
   U4741 : INV_X2 port map( I => n30277, ZN => n837);
   U4749 : INV_X1 port map( I => n10048, ZN => n7602);
   U4760 : NAND2_X1 port map( A1 => n9178, A2 => n10687, ZN => n11788);
   U4766 : AOI21_X1 port map( A1 => n27159, A2 => n26750, B => n24106, ZN => 
                           n13237);
   U4769 : NAND2_X1 port map( A1 => n10687, A2 => n32737, ZN => n15158);
   U4787 : NOR2_X1 port map( A1 => n6474, A2 => n14078, ZN => n9812);
   U4803 : INV_X1 port map( I => n17285, ZN => n23708);
   U4811 : INV_X1 port map( I => n17857, ZN => n23857);
   U4812 : INV_X1 port map( I => n23287, ZN => n23242);
   U4815 : INV_X1 port map( I => n3600, ZN => n4777);
   U4819 : NAND2_X1 port map( A1 => n3773, A2 => n22977, ZN => n2624);
   U4833 : INV_X1 port map( I => n9335, ZN => n9334);
   U4865 : INV_X1 port map( I => n19894, ZN => n20417);
   U4867 : INV_X1 port map( I => n20595, ZN => n20499);
   U4879 : INV_X2 port map( I => n571, ZN => n14559);
   U4894 : AOI21_X1 port map( A1 => n18835, A2 => n13846, B => n18832, ZN => 
                           n14393);
   U4917 : AOI22_X1 port map( A1 => n12783, A2 => n24969, B1 => n8622, B2 => 
                           n27134, ZN => n3136);
   U4953 : AOI21_X1 port map( A1 => n25637, A2 => n9718, B => n27188, ZN => 
                           n9717);
   U4954 : OR2_X1 port map( A1 => n25876, A2 => n1211, Z => n3955);
   U4959 : NAND3_X1 port map( A1 => n14630, A2 => n17595, A3 => n14629, ZN => 
                           n14628);
   U4963 : AOI21_X1 port map( A1 => n17169, A2 => n24606, B => n9941, ZN => 
                           n24025);
   U4977 : NOR2_X1 port map( A1 => n1083, A2 => n34115, ZN => n8840);
   U4995 : AOI21_X1 port map( A1 => n9202, A2 => n970, B => n9275, ZN => n9366)
                           ;
   U5022 : NAND2_X1 port map( A1 => n23715, A2 => n707, ZN => n6248);
   U5045 : INV_X1 port map( I => n11621, ZN => n4111);
   U5076 : NAND2_X1 port map( A1 => n2418, A2 => n22567, ZN => n22444);
   U5095 : NAND2_X1 port map( A1 => n12794, A2 => n34046, ZN => n21576);
   U5102 : INV_X1 port map( I => n7753, ZN => n21752);
   U5122 : INV_X1 port map( I => n20650, ZN => n20270);
   U5161 : NOR2_X1 port map( A1 => n12316, A2 => n18993, ZN => n1453);
   U5175 : NAND2_X1 port map( A1 => n5328, A2 => n5327, ZN => n4053);
   U5180 : NAND3_X1 port map( A1 => n17073, A2 => n10786, A3 => n29659, ZN => 
                           n10785);
   U5181 : INV_X1 port map( I => n5328, ZN => n4178);
   U5186 : NOR2_X1 port map( A1 => n493, A2 => n16450, ZN => n5753);
   U5194 : NAND4_X1 port map( A1 => n5622, A2 => n25206, A3 => n5621, A4 => 
                           n7304, ZN => n7302);
   U5195 : NAND3_X1 port map( A1 => n4770, A2 => n4781, A3 => n10858, ZN => 
                           n4769);
   U5200 : NOR2_X1 port map( A1 => n4781, A2 => n9247, ZN => n3988);
   U5221 : NOR2_X1 port map( A1 => n24484, A2 => n17684, ZN => n6365);
   U5230 : INV_X1 port map( I => n11409, ZN => n25263);
   U5234 : NAND2_X1 port map( A1 => n15555, A2 => n25870, ZN => n15670);
   U5236 : INV_X2 port map( I => n17861, ZN => n25292);
   U5240 : INV_X2 port map( I => n15295, ZN => n13032);
   U5241 : INV_X1 port map( I => n1786, ZN => n25203);
   U5242 : INV_X1 port map( I => n17092, ZN => n15355);
   U5249 : NOR2_X1 port map( A1 => n25564, A2 => n25582, ZN => n25634);
   U5290 : NAND2_X1 port map( A1 => n707, A2 => n8370, ZN => n7190);
   U5295 : NAND2_X1 port map( A1 => n23816, A2 => n17616, ZN => n17816);
   U5301 : NAND2_X1 port map( A1 => n23949, A2 => n11621, ZN => n9894);
   U5303 : NAND2_X1 port map( A1 => n15865, A2 => n27136, ZN => n23555);
   U5304 : OAI21_X1 port map( A1 => n3553, A2 => n11621, B => n30360, ZN => 
                           n3552);
   U5309 : INV_X1 port map( I => n16536, ZN => n23713);
   U5311 : AND2_X1 port map( A1 => n34009, A2 => n28914, Z => n8850);
   U5315 : OAI21_X1 port map( A1 => n847, A2 => n8760, B => n23721, ZN => 
                           n23115);
   U5324 : INV_X1 port map( I => n11887, ZN => n7088);
   U5328 : INV_X2 port map( I => n17591, ZN => n23888);
   U5329 : INV_X1 port map( I => n26114, ZN => n16097);
   U5331 : INV_X2 port map( I => n9798, ZN => n11943);
   U5335 : INV_X2 port map( I => n23286, ZN => n770);
   U5337 : NAND3_X1 port map( A1 => n10528, A2 => n28891, A3 => n1271, ZN => 
                           n17774);
   U5375 : NOR2_X1 port map( A1 => n22608, A2 => n32512, ZN => n7426);
   U5378 : NAND2_X1 port map( A1 => n22535, A2 => n22428, ZN => n22540);
   U5433 : INV_X1 port map( I => n17746, ZN => n15468);
   U5443 : NAND3_X1 port map( A1 => n6405, A2 => n13451, A3 => n32746, ZN => 
                           n13301);
   U5471 : INV_X1 port map( I => n13450, ZN => n19051);
   U5476 : OAI21_X1 port map( A1 => n12707, A2 => n19048, B => n28705, ZN => 
                           n12600);
   U5482 : NAND2_X1 port map( A1 => n5545, A2 => n5889, ZN => n5907);
   U5508 : NAND2_X1 port map( A1 => n13360, A2 => n8208, ZN => n17073);
   U5509 : INV_X1 port map( I => n3344, ZN => n18311);
   U5516 : INV_X1 port map( I => n13531, ZN => n1063);
   U5536 : NAND2_X1 port map( A1 => n830, A2 => n27123, ZN => n3706);
   U5542 : NAND3_X1 port map( A1 => n715, A2 => n25220, A3 => n25210, ZN => 
                           n7304);
   U5545 : INV_X1 port map( I => n31236, ZN => n25550);
   U5555 : INV_X1 port map( I => n25746, ZN => n832);
   U5559 : AOI22_X1 port map( A1 => n4492, A2 => n31920, B1 => n4407, B2 => 
                           n4491, ZN => n5886);
   U5566 : AND2_X1 port map( A1 => n833, A2 => n24667, Z => n25537);
   U5573 : NAND2_X1 port map( A1 => n13985, A2 => n25261, ZN => n24581);
   U5576 : AND2_X1 port map( A1 => n25334, A2 => n25536, Z => n12088);
   U5578 : NOR2_X1 port map( A1 => n317, A2 => n6551, ZN => n6640);
   U5580 : AOI21_X1 port map( A1 => n15235, A2 => n33393, B => n765, ZN => 
                           n5929);
   U5581 : NAND3_X1 port map( A1 => n10497, A2 => n15295, A3 => n2378, ZN => 
                           n25715);
   U5582 : AOI22_X1 port map( A1 => n15235, A2 => n25561, B1 => n765, B2 => 
                           n16704, ZN => n5930);
   U5591 : AND2_X1 port map( A1 => n25586, A2 => n25590, Z => n12423);
   U5592 : NAND2_X1 port map( A1 => n678, A2 => n25409, ZN => n25326);
   U5599 : INV_X1 port map( I => n25115, ZN => n16025);
   U5613 : INV_X1 port map( I => n24763, ZN => n1225);
   U5625 : NAND2_X1 port map( A1 => n24156, A2 => n10513, ZN => n9283);
   U5627 : NAND3_X1 port map( A1 => n7150, A2 => n16868, A3 => n24253, ZN => 
                           n3546);
   U5640 : AND2_X1 port map( A1 => n24061, A2 => n24156, Z => n2463);
   U5641 : NAND3_X1 port map( A1 => n767, A2 => n29566, A3 => n2847, ZN => 
                           n7094);
   U5700 : NAND3_X1 port map( A1 => n23867, A2 => n17895, A3 => n23868, ZN => 
                           n23821);
   U5701 : NAND3_X1 port map( A1 => n8408, A2 => n23868, A3 => n1257, ZN => 
                           n10132);
   U5717 : NAND2_X1 port map( A1 => n23947, A2 => n4111, ZN => n1525);
   U5735 : INV_X1 port map( I => n23346, ZN => n23132);
   U5746 : AND3_X1 port map( A1 => n4067, A2 => n22826, A3 => n30437, Z => 
                           n22652);
   U5766 : OAI21_X1 port map( A1 => n6593, A2 => n17720, B => n22955, ZN => 
                           n2002);
   U5777 : INV_X1 port map( I => n17890, ZN => n22389);
   U5788 : NAND3_X1 port map( A1 => n902, A2 => n22330, A3 => n14376, ZN => 
                           n11008);
   U5795 : INV_X1 port map( I => n29451, ZN => n14008);
   U5801 : INV_X1 port map( I => n22576, ZN => n16148);
   U5815 : OAI21_X1 port map( A1 => n21123, A2 => n31910, B => n31260, ZN => 
                           n21126);
   U5838 : INV_X2 port map( I => n21432, ZN => n5049);
   U5840 : AOI21_X1 port map( A1 => n21453, A2 => n9186, B => n780, ZN => n9393
                           );
   U5841 : NOR2_X1 port map( A1 => n11966, A2 => n21367, ZN => n2605);
   U5847 : INV_X1 port map( I => n8398, ZN => n3931);
   U5862 : OAI21_X1 port map( A1 => n26182, A2 => n20545, B => n3157, ZN => 
                           n13631);
   U5870 : OAI21_X1 port map( A1 => n2566, A2 => n17497, B => n8293, ZN => 
                           n19955);
   U5875 : NAND4_X1 port map( A1 => n1678, A2 => n1680, A3 => n1677, A4 => 
                           n1679, ZN => n20306);
   U5886 : OAI21_X1 port map( A1 => n10286, A2 => n18142, B => n14306, ZN => 
                           n3945);
   U5901 : NOR2_X1 port map( A1 => n13605, A2 => n20088, ZN => n11501);
   U5907 : INV_X2 port map( I => n4881, ZN => n6275);
   U5908 : AND2_X1 port map( A1 => n16489, A2 => n20052, Z => n16675);
   U5916 : INV_X1 port map( I => n11910, ZN => n19863);
   U5944 : NAND2_X1 port map( A1 => n27726, A2 => n3388, ZN => n3390);
   U5959 : OAI21_X1 port map( A1 => n15495, A2 => n9937, B => n16538, ZN => 
                           n15576);
   U5962 : OR2_X2 port map( A1 => n18709, A2 => n17625, Z => n10700);
   U5964 : NOR2_X1 port map( A1 => n15902, A2 => n1709, ZN => n9937);
   U5974 : NOR2_X1 port map( A1 => n13548, A2 => n15146, ZN => n13526);
   U5997 : INV_X1 port map( I => n17189, ZN => n881);
   U5999 : INV_X2 port map( I => n18559, ZN => n828);
   U6002 : CLKBUF_X2 port map( I => Key(58), Z => n16691);
   U6004 : CLKBUF_X2 port map( I => Key(187), Z => n16655);
   U6006 : CLKBUF_X2 port map( I => Key(91), Z => n24869);
   U6007 : CLKBUF_X2 port map( I => Key(79), Z => n16555);
   U6010 : CLKBUF_X2 port map( I => Key(151), Z => n16654);
   U6015 : NOR2_X1 port map( A1 => n17927, A2 => n27123, ZN => n9703);
   U6020 : AOI21_X1 port map( A1 => n714, A2 => n25007, B => n3232, ZN => n3231
                           );
   U6021 : OAI21_X1 port map( A1 => n1076, A2 => n10376, B => n25724, ZN => 
                           n4253);
   U6022 : AND2_X1 port map( A1 => n27123, A2 => n786, Z => n12060);
   U6023 : NOR2_X1 port map( A1 => n27123, A2 => n9247, ZN => n3435);
   U6025 : OR2_X1 port map( A1 => n4415, A2 => n25744, Z => n24432);
   U6027 : INV_X1 port map( I => n32859, ZN => n25105);
   U6029 : NAND2_X1 port map( A1 => n28358, A2 => n16509, ZN => n25216);
   U6030 : NOR2_X1 port map( A1 => n5926, A2 => n5942, ZN => n5918);
   U6042 : INV_X2 port map( I => n16509, ZN => n15340);
   U6053 : INV_X1 port map( I => n25200, ZN => n17005);
   U6055 : NOR2_X1 port map( A1 => n27651, A2 => n16025, ZN => n12165);
   U6056 : OAI21_X1 port map( A1 => n25134, A2 => n5611, B => n16589, ZN => 
                           n25135);
   U6057 : NOR2_X1 port map( A1 => n25117, A2 => n14495, ZN => n9956);
   U6058 : INV_X1 port map( I => n24724, ZN => n7963);
   U6059 : NOR2_X1 port map( A1 => n14495, A2 => n27651, ZN => n8608);
   U6065 : AND2_X1 port map( A1 => n25884, A2 => n15152, Z => n25886);
   U6068 : NOR2_X1 port map( A1 => n25229, A2 => n13985, ZN => n9427);
   U6080 : INV_X1 port map( I => n25977, ZN => n1224);
   U6104 : NAND2_X1 port map( A1 => n7361, A2 => n8399, ZN => n13632);
   U6112 : AND2_X1 port map( A1 => n7060, A2 => n16643, Z => n7059);
   U6128 : NOR2_X1 port map( A1 => n17178, A2 => n17180, ZN => n16663);
   U6129 : NAND2_X1 port map( A1 => n24177, A2 => n4897, ZN => n5041);
   U6153 : NOR2_X1 port map( A1 => n28222, A2 => n23754, ZN => n23347);
   U6160 : OAI21_X1 port map( A1 => n6869, A2 => n23917, B => n8372, ZN => 
                           n23116);
   U6181 : AND2_X1 port map( A1 => n29272, A2 => n756, Z => n7710);
   U6198 : NAND2_X1 port map( A1 => n17895, A2 => n657, ZN => n3650);
   U6207 : NOR2_X1 port map( A1 => n16431, A2 => n29270, ZN => n23643);
   U6209 : NAND2_X1 port map( A1 => n1099, A2 => n29323, ZN => n12817);
   U6216 : INV_X2 port map( I => n17506, ZN => n843);
   U6238 : OR2_X1 port map( A1 => n22868, A2 => n25994, Z => n7103);
   U6253 : NAND2_X1 port map( A1 => n12729, A2 => n16458, ZN => n12726);
   U6256 : INV_X1 port map( I => n27719, ZN => n11565);
   U6263 : NAND3_X1 port map( A1 => n23066, A2 => n4734, A3 => n13807, ZN => 
                           n10411);
   U6265 : NAND3_X1 port map( A1 => n805, A2 => n2479, A3 => n31795, ZN => 
                           n7582);
   U6266 : NAND3_X1 port map( A1 => n1109, A2 => n31129, A3 => n22798, ZN => 
                           n17481);
   U6308 : AND2_X1 port map( A1 => n22430, A2 => n2538, Z => n2537);
   U6309 : AND2_X1 port map( A1 => n16529, A2 => n9515, Z => n9516);
   U6310 : NAND3_X1 port map( A1 => n14008, A2 => n809, A3 => n16483, ZN => 
                           n14066);
   U6324 : NAND2_X1 port map( A1 => n22575, A2 => n5743, ZN => n5744);
   U6330 : OAI21_X1 port map( A1 => n14251, A2 => n32830, B => n14253, ZN => 
                           n1663);
   U6351 : NAND2_X1 port map( A1 => n11629, A2 => n22486, ZN => n8318);
   U6354 : INV_X1 port map( I => n29868, ZN => n22359);
   U6370 : NOR2_X1 port map( A1 => n13167, A2 => n2801, ZN => n7017);
   U6428 : NOR2_X1 port map( A1 => n21074, A2 => n21434, ZN => n14951);
   U6438 : OR2_X1 port map( A1 => n12441, A2 => n21353, Z => n12465);
   U6441 : NOR2_X1 port map( A1 => n11272, A2 => n21095, ZN => n7512);
   U6455 : AND3_X1 port map( A1 => n10599, A2 => n21239, A3 => n5822, Z => 
                           n13100);
   U6470 : INV_X1 port map( I => n20730, ZN => n20824);
   U6501 : OR3_X1 port map( A1 => n6679, A2 => n1357, A3 => n20635, Z => n6616)
                           ;
   U6506 : OR2_X1 port map( A1 => n13282, A2 => n28836, Z => n12115);
   U6513 : INV_X1 port map( I => n20605, ZN => n20130);
   U6517 : OAI21_X1 port map( A1 => n8100, A2 => n29253, B => n19850, ZN => 
                           n19234);
   U6520 : NAND3_X1 port map( A1 => n12253, A2 => n18119, A3 => n1168, ZN => 
                           n4854);
   U6533 : NOR2_X1 port map( A1 => n1172, A2 => n31161, ZN => n3311);
   U6535 : NAND2_X1 port map( A1 => n16848, A2 => n29153, ZN => n6960);
   U6537 : NAND3_X1 port map( A1 => n15665, A2 => n4180, A3 => n20056, ZN => 
                           n15313);
   U6539 : OR2_X1 port map( A1 => n19456, A2 => n28293, Z => n19994);
   U6543 : NAND3_X1 port map( A1 => n4215, A2 => n33419, A3 => n20156, ZN => 
                           n8589);
   U6548 : INV_X1 port map( I => n19936, ZN => n14172);
   U6551 : INV_X2 port map( I => n29254, ZN => n1168);
   U6570 : INV_X1 port map( I => n15786, ZN => n19524);
   U6580 : NAND3_X1 port map( A1 => n3822, A2 => n19016, A3 => n19017, ZN => 
                           n4985);
   U6585 : AOI21_X1 port map( A1 => n16669, A2 => n18838, B => n13925, ZN => 
                           n18839);
   U6589 : AND2_X1 port map( A1 => n19183, A2 => n2612, Z => n7568);
   U6598 : NAND3_X1 port map( A1 => n28379, A2 => n16740, A3 => n19140, ZN => 
                           n5333);
   U6611 : AND2_X1 port map( A1 => n10423, A2 => n29781, Z => n2149);
   U6633 : OAI21_X1 port map( A1 => n15018, A2 => n8376, B => n9886, ZN => 
                           n3023);
   U6637 : NAND3_X1 port map( A1 => n952, A2 => n711, A3 => n29315, ZN => 
                           n10306);
   U6647 : NAND2_X1 port map( A1 => n15902, A2 => n11459, ZN => n10133);
   U6653 : NAND2_X1 port map( A1 => n18480, A2 => n18605, ZN => n16763);
   U6657 : NOR2_X1 port map( A1 => n6783, A2 => n11389, ZN => n14843);
   U6661 : NOR2_X1 port map( A1 => n18682, A2 => n1659, ZN => n12051);
   U6677 : NAND2_X1 port map( A1 => n4677, A2 => n33621, ZN => n6777);
   U6680 : NAND2_X1 port map( A1 => n4808, A2 => n962, ZN => n11389);
   U6697 : OR2_X2 port map( A1 => n16855, A2 => n7216, Z => n3779);
   U6699 : NAND2_X1 port map( A1 => n6783, A2 => n14926, ZN => n6887);
   U6702 : NAND2_X1 port map( A1 => n493, A2 => n498, ZN => n17557);
   U6704 : NOR2_X1 port map( A1 => n9766, A2 => n16420, ZN => n15697);
   U6708 : NAND2_X1 port map( A1 => n16855, A2 => n7216, ZN => n14906);
   U6714 : AND2_X1 port map( A1 => n17223, A2 => n16948, Z => n8948);
   U6719 : BUF_X2 port map( I => n16450, Z => n5473);
   U6720 : INV_X1 port map( I => n25578, ZN => n960);
   U6723 : CLKBUF_X2 port map( I => Key(82), Z => n16642);
   U6725 : CLKBUF_X2 port map( I => Key(87), Z => n25465);
   U6726 : CLKBUF_X2 port map( I => Key(80), Z => n25720);
   U6728 : INV_X2 port map( I => n18085, ZN => n882);
   U6729 : CLKBUF_X2 port map( I => Key(14), Z => n25880);
   U6736 : NOR2_X1 port map( A1 => n12431, A2 => n25271, ZN => n10605);
   U6737 : NAND2_X1 port map( A1 => n25571, A2 => n5942, ZN => n3638);
   U6739 : AND2_X1 port map( A1 => n5043, A2 => n15340, Z => n4613);
   U6740 : NAND2_X1 port map( A1 => n3646, A2 => n2191, ZN => n25256);
   U6743 : NOR2_X1 port map( A1 => n28736, A2 => n25128, ZN => n6828);
   U6745 : NOR2_X1 port map( A1 => n31456, A2 => n30241, ZN => n14873);
   U6758 : NOR2_X1 port map( A1 => n10097, A2 => n967, ZN => n8247);
   U6763 : OAI21_X1 port map( A1 => n25202, A2 => n16632, B => n25203, ZN => 
                           n3385);
   U6770 : INV_X1 port map( I => n16783, ZN => n6641);
   U6772 : OR2_X1 port map( A1 => n15425, A2 => n29063, Z => n14925);
   U6775 : AND2_X1 port map( A1 => n12039, A2 => n6034, Z => n6825);
   U6783 : NAND2_X1 port map( A1 => n11049, A2 => n16066, ZN => n3212);
   U6790 : NAND2_X1 port map( A1 => n8058, A2 => n24094, ZN => n23382);
   U6794 : NOR2_X1 port map( A1 => n7097, A2 => n7361, ZN => n7100);
   U6801 : OAI21_X1 port map( A1 => n32520, A2 => n23995, B => n15175, ZN => 
                           n9659);
   U6804 : AOI21_X1 port map( A1 => n10987, A2 => n24328, B => n24245, ZN => 
                           n7097);
   U6811 : OAI21_X1 port map( A1 => n24210, A2 => n24212, B => n24211, ZN => 
                           n6840);
   U6815 : NAND2_X1 port map( A1 => n24132, A2 => n32102, ZN => n8336);
   U6816 : NOR2_X1 port map( A1 => n4024, A2 => n7503, ZN => n24202);
   U6817 : NAND3_X1 port map( A1 => n24097, A2 => n840, A3 => n26516, ZN => 
                           n24038);
   U6820 : NAND2_X1 port map( A1 => n24092, A2 => n17261, ZN => n5914);
   U6833 : NAND2_X1 port map( A1 => n23347, A2 => n28297, ZN => n14118);
   U6841 : INV_X1 port map( I => n31096, ZN => n14891);
   U6871 : NOR2_X1 port map( A1 => n23848, A2 => n15423, ZN => n6132);
   U6885 : NOR2_X1 port map( A1 => n23872, A2 => n23695, ZN => n23577);
   U6892 : NOR2_X1 port map( A1 => n13308, A2 => n23949, ZN => n3553);
   U6910 : NAND2_X1 port map( A1 => n2623, A2 => n30573, ZN => n11669);
   U6931 : NOR2_X1 port map( A1 => n8954, A2 => n13751, ZN => n8953);
   U6934 : INV_X1 port map( I => n22862, ZN => n9435);
   U6935 : OAI21_X1 port map( A1 => n10644, A2 => n849, B => n10411, ZN => 
                           n10410);
   U6938 : OR2_X1 port map( A1 => n28314, A2 => n22810, Z => n15730);
   U6953 : NOR2_X1 port map( A1 => n12727, A2 => n851, ZN => n5982);
   U6954 : AND2_X1 port map( A1 => n23096, A2 => n25979, Z => n3173);
   U6966 : NAND2_X1 port map( A1 => n13694, A2 => n5915, ZN => n4182);
   U6967 : INV_X1 port map( I => n23111, ZN => n17099);
   U6969 : OAI21_X1 port map( A1 => n13008, A2 => n29335, B => n12688, ZN => 
                           n12687);
   U6977 : NAND2_X1 port map( A1 => n10388, A2 => n22681, ZN => n10387);
   U6986 : NOR2_X1 port map( A1 => n15260, A2 => n30668, ZN => n7659);
   U7001 : INV_X1 port map( I => n22393, ZN => n7490);
   U7007 : NOR2_X1 port map( A1 => n27402, A2 => n22550, ZN => n8098);
   U7009 : NOR2_X1 port map( A1 => n26878, A2 => n29078, ZN => n1519);
   U7014 : AOI21_X1 port map( A1 => n628, A2 => n9234, B => n9757, ZN => n15643
                           );
   U7036 : NOR2_X1 port map( A1 => n22595, A2 => n22599, ZN => n4055);
   U7037 : INV_X1 port map( I => n1289, ZN => n11244);
   U7046 : INV_X2 port map( I => n17899, ZN => n907);
   U7047 : INV_X1 port map( I => n22078, ZN => n11859);
   U7064 : AOI22_X1 port map( A1 => n534, A2 => n31765, B1 => n28450, B2 => 
                           n3821, ZN => n10874);
   U7081 : NOR2_X1 port map( A1 => n21856, A2 => n21, ZN => n1595);
   U7082 : NOR2_X1 port map( A1 => n30885, A2 => n1013, ZN => n4435);
   U7085 : NOR2_X1 port map( A1 => n27178, A2 => n21719, ZN => n21720);
   U7106 : AND2_X1 port map( A1 => n16386, A2 => n21842, Z => n1535);
   U7115 : OAI22_X1 port map( A1 => n17078, A2 => n14640, B1 => n1652, B2 => 
                           n14577, ZN => n1769);
   U7118 : INV_X1 port map( I => n21350, ZN => n1012);
   U7119 : NOR2_X1 port map( A1 => n10720, A2 => n12561, ZN => n15747);
   U7124 : NAND2_X1 port map( A1 => n14577, A2 => n1652, ZN => n21723);
   U7128 : INV_X2 port map( I => n8313, ZN => n915);
   U7135 : INV_X1 port map( I => n8140, ZN => n1139);
   U7142 : INV_X1 port map( I => n18213, ZN => n6471);
   U7157 : AOI21_X1 port map( A1 => n28642, A2 => n1017, B => n20676, ZN => 
                           n20677);
   U7172 : NAND2_X1 port map( A1 => n6451, A2 => n26167, ZN => n1784);
   U7204 : INV_X1 port map( I => n20657, ZN => n21249);
   U7207 : AOI21_X1 port map( A1 => n9405, A2 => n21452, B => n21237, ZN => 
                           n9406);
   U7210 : INV_X1 port map( I => n30727, ZN => n8393);
   U7240 : INV_X1 port map( I => n20836, ZN => n1592);
   U7259 : NOR2_X1 port map( A1 => n16146, A2 => n14719, ZN => n4857);
   U7263 : NOR2_X1 port map( A1 => n28390, A2 => n20549, ZN => n10834);
   U7264 : NAND3_X1 port map( A1 => n20575, A2 => n420, A3 => n20571, ZN => 
                           n4816);
   U7273 : INV_X1 port map( I => n20430, ZN => n11017);
   U7287 : NAND2_X1 port map( A1 => n13631, A2 => n28261, ZN => n13630);
   U7301 : NOR2_X1 port map( A1 => n20267, A2 => n26585, ZN => n8293);
   U7304 : INV_X1 port map( I => n10939, ZN => n20452);
   U7313 : NAND3_X1 port map( A1 => n20256, A2 => n13380, A3 => n20404, ZN => 
                           n13379);
   U7321 : BUF_X2 port map( I => n16452, Z => n10057);
   U7332 : NAND2_X1 port map( A1 => n13611, A2 => n12078, ZN => n13608);
   U7339 : NAND2_X1 port map( A1 => n5642, A2 => n17456, ZN => n5641);
   U7346 : AOI21_X1 port map( A1 => n29357, A2 => n29013, B => n10340, ZN => 
                           n19822);
   U7347 : NAND2_X1 port map( A1 => n19876, A2 => n31103, ZN => n20289);
   U7380 : INV_X1 port map( I => n11593, ZN => n13841);
   U7386 : NAND2_X1 port map( A1 => n1039, A2 => n14281, ZN => n2291);
   U7389 : NAND2_X1 port map( A1 => n13912, A2 => n5073, ZN => n4051);
   U7394 : AND2_X1 port map( A1 => n9748, A2 => n3526, Z => n3525);
   U7401 : AND2_X1 port map( A1 => n8301, A2 => n20008, Z => n9875);
   U7418 : INV_X1 port map( I => n10696, ZN => n20157);
   U7429 : INV_X1 port map( I => n8808, ZN => n12100);
   U7432 : INV_X1 port map( I => n20088, ZN => n16493);
   U7439 : NOR3_X1 port map( A1 => n19174, A2 => n19134, A3 => n3535, ZN => 
                           n19135);
   U7455 : NAND2_X1 port map( A1 => n17370, A2 => n16699, ZN => n1450);
   U7458 : NOR2_X1 port map( A1 => n19313, A2 => n19152, ZN => n11075);
   U7468 : NAND2_X1 port map( A1 => n19604, A2 => n2799, ZN => n3391);
   U7474 : NAND2_X1 port map( A1 => n19176, A2 => n19253, ZN => n2123);
   U7476 : NOR2_X1 port map( A1 => n18994, A2 => n14892, ZN => n5655);
   U7478 : AOI22_X1 port map( A1 => n19287, A2 => n3388, B1 => n6059, B2 => 
                           n27726, ZN => n1869);
   U7479 : NOR2_X1 port map( A1 => n16916, A2 => n18979, ZN => n2390);
   U7486 : NOR2_X1 port map( A1 => n8606, A2 => n19229, ZN => n9424);
   U7504 : AND2_X1 port map( A1 => n19313, A2 => n763, Z => n18969);
   U7508 : AND2_X1 port map( A1 => n12707, A2 => n30682, Z => n12131);
   U7510 : NOR2_X1 port map( A1 => n16274, A2 => n9553, ZN => n3244);
   U7511 : OR2_X1 port map( A1 => n27726, A2 => n17817, Z => n3365);
   U7512 : NOR2_X1 port map( A1 => n19107, A2 => n19108, ZN => n10054);
   U7524 : INV_X2 port map( I => n19123, ZN => n8233);
   U7526 : AND2_X1 port map( A1 => n25985, A2 => n1056, Z => n9710);
   U7537 : OR2_X2 port map( A1 => n10365, A2 => n4659, Z => n4656);
   U7565 : OAI21_X1 port map( A1 => n31579, A2 => n4259, B => n18768, ZN => 
                           n18765);
   U7581 : AOI21_X1 port map( A1 => n13514, A2 => n8376, B => n7454, ZN => 
                           n11555);
   U7584 : NAND2_X1 port map( A1 => n18795, A2 => n6119, ZN => n7682);
   U7585 : AOI21_X1 port map( A1 => n3601, A2 => n11941, B => n26717, ZN => 
                           n3111);
   U7586 : NAND2_X1 port map( A1 => n17359, A2 => n18737, ZN => n7733);
   U7590 : NOR2_X1 port map( A1 => n17687, A2 => n18863, ZN => n4506);
   U7595 : NAND2_X1 port map( A1 => n18511, A2 => n16855, ZN => n14453);
   U7596 : OAI21_X1 port map( A1 => n13254, A2 => n34141, B => n4677, ZN => 
                           n12173);
   U7598 : NOR2_X1 port map( A1 => n17477, A2 => n1060, ZN => n6890);
   U7599 : OAI21_X1 port map( A1 => n18785, A2 => n18801, B => n8395, ZN => 
                           n18628);
   U7600 : NAND3_X1 port map( A1 => n3601, A2 => n10095, A3 => n732, ZN => 
                           n3149);
   U7603 : NAND2_X1 port map( A1 => n9766, A2 => n31724, ZN => n11693);
   U7607 : NOR2_X1 port map( A1 => n18815, A2 => n11918, ZN => n8043);
   U7611 : NAND2_X1 port map( A1 => n18797, A2 => n16420, ZN => n7713);
   U7613 : NOR2_X1 port map( A1 => n18706, A2 => n18707, ZN => n18745);
   U7621 : INV_X1 port map( I => n10182, ZN => n1189);
   U7626 : AND2_X1 port map( A1 => n9909, A2 => n11459, Z => n15495);
   U7628 : NAND2_X1 port map( A1 => n16766, A2 => n31579, ZN => n18764);
   U7630 : INV_X1 port map( I => n25832, ZN => n1064);
   U7631 : INV_X1 port map( I => n25493, ZN => n1065);
   U7636 : INV_X1 port map( I => n18335, ZN => n18481);
   U7638 : INV_X2 port map( I => n32034, ZN => n13254);
   U7642 : INV_X1 port map( I => n16464, ZN => n1070);
   U7643 : BUF_X2 port map( I => n9909, Z => n1709);
   U7644 : INV_X1 port map( I => n11905, ZN => n8208);
   U7646 : INV_X1 port map( I => n16548, ZN => n1419);
   U7647 : INV_X1 port map( I => n25108, ZN => n1067);
   U7653 : INV_X1 port map( I => n16701, ZN => n1069);
   U7654 : CLKBUF_X2 port map( I => Key(102), Z => n16548);
   U7656 : CLKBUF_X2 port map( I => Key(93), Z => n24968);
   U7657 : CLKBUF_X2 port map( I => Key(65), Z => n24386);
   U7664 : CLKBUF_X2 port map( I => Key(132), Z => n24943);
   U7665 : INV_X2 port map( I => n16914, ZN => n962);
   U7667 : CLKBUF_X2 port map( I => Key(101), Z => n16423);
   U7676 : OAI21_X1 port map( A1 => n25746, A2 => n27189, B => n1979, ZN => 
                           n4417);
   U7679 : NAND3_X1 port map( A1 => n11003, A2 => n25816, A3 => n25804, ZN => 
                           n11004);
   U7683 : NAND2_X1 port map( A1 => n6111, A2 => n13624, ZN => n5917);
   U7684 : NAND2_X1 port map( A1 => n7929, A2 => n14511, ZN => n11133);
   U7685 : INV_X1 port map( I => n25223, ZN => n4188);
   U7688 : NAND2_X1 port map( A1 => n25247, A2 => n2191, ZN => n11135);
   U7690 : NAND2_X1 port map( A1 => n25743, A2 => n32863, ZN => n9414);
   U7692 : NAND2_X1 port map( A1 => n25006, A2 => n3232, ZN => n3155);
   U7693 : NAND2_X1 port map( A1 => n715, A2 => n25214, ZN => n4614);
   U7697 : AND2_X1 port map( A1 => n7273, A2 => n1395, Z => n7270);
   U7699 : INV_X1 port map( I => n11571, ZN => n8035);
   U7701 : NAND2_X1 port map( A1 => n25220, A2 => n7515, ZN => n25222);
   U7706 : INV_X4 port map( I => n24896, ZN => n965);
   U7707 : INV_X1 port map( I => n2983, ZN => n2876);
   U7710 : NAND2_X1 port map( A1 => n885, A2 => n17684, ZN => n4101);
   U7712 : NAND2_X1 port map( A1 => n10570, A2 => n25289, ZN => n5535);
   U7717 : NOR2_X1 port map( A1 => n24884, A2 => n25020, ZN => n6473);
   U7721 : INV_X1 port map( I => n7081, ZN => n10748);
   U7725 : NOR3_X1 port map( A1 => n14454, A2 => n24780, A3 => n15719, ZN => 
                           n2996);
   U7730 : OAI21_X1 port map( A1 => n13042, A2 => n25885, B => n25871, ZN => 
                           n8541);
   U7731 : NAND2_X1 port map( A1 => n15318, A2 => n4885, ZN => n5659);
   U7740 : NOR2_X1 port map( A1 => n5202, A2 => n25119, ZN => n5203);
   U7741 : INV_X4 port map( I => n25382, ZN => n16783);
   U7743 : OAI21_X1 port map( A1 => n2158, A2 => n2156, B => n10924, ZN => 
                           n1645);
   U7760 : NAND2_X1 port map( A1 => n24051, A2 => n15720, ZN => n15790);
   U7767 : NOR2_X1 port map( A1 => n9202, A2 => n796, ZN => n17601);
   U7786 : AOI21_X1 port map( A1 => n9323, A2 => n6286, B => n16651, ZN => 
                           n3548);
   U7791 : NAND2_X1 port map( A1 => n2558, A2 => n14399, ZN => n14995);
   U7792 : OAI21_X1 port map( A1 => n13175, A2 => n24110, B => n10530, ZN => 
                           n10529);
   U7793 : OAI21_X1 port map( A1 => n28945, A2 => n11200, B => n13356, ZN => 
                           n24178);
   U7796 : OR3_X1 port map( A1 => n1087, A2 => n13343, A3 => n17068, Z => 
                           n24115);
   U7803 : INV_X2 port map( I => n14123, ZN => n1088);
   U7805 : OAI21_X1 port map( A1 => n26158, A2 => n1775, B => n27931, ZN => 
                           n5045);
   U7811 : OR2_X1 port map( A1 => n16643, A2 => n3718, Z => n2686);
   U7812 : INV_X1 port map( I => n7581, ZN => n24236);
   U7831 : NOR2_X1 port map( A1 => n15660, A2 => n4408, ZN => n3995);
   U7832 : NAND2_X1 port map( A1 => n17980, A2 => n14664, ZN => n14166);
   U7849 : NOR2_X1 port map( A1 => n13521, A2 => n895, ZN => n5954);
   U7851 : NAND2_X1 port map( A1 => n15623, A2 => n23910, ZN => n3449);
   U7861 : NAND3_X1 port map( A1 => n4177, A2 => n28347, A3 => n23857, ZN => 
                           n23801);
   U7869 : OR2_X1 port map( A1 => n23778, A2 => n11392, Z => n11391);
   U7882 : NAND2_X1 port map( A1 => n29294, A2 => n11676, ZN => n9893);
   U7890 : NOR2_X1 port map( A1 => n10193, A2 => n34008, ZN => n12070);
   U7914 : NOR2_X1 port map( A1 => n22400, A2 => n33007, ZN => n11411);
   U7934 : NAND2_X1 port map( A1 => n1104, A2 => n10528, ZN => n2342);
   U7935 : OAI21_X1 port map( A1 => n1106, A2 => n7463, B => n3668, ZN => n3783
                           );
   U7944 : NAND2_X1 port map( A1 => n22944, A2 => n3657, ZN => n9259);
   U7948 : NAND2_X1 port map( A1 => n1484, A2 => n23104, ZN => n10790);
   U7950 : NAND3_X1 port map( A1 => n31531, A2 => n22981, A3 => n32935, ZN => 
                           n17411);
   U7951 : NOR2_X1 port map( A1 => n23109, A2 => n853, ZN => n5895);
   U7957 : NOR2_X1 port map( A1 => n6453, A2 => n16022, ZN => n4937);
   U7960 : OAI21_X1 port map( A1 => n29242, A2 => n31798, B => n22828, ZN => 
                           n8200);
   U7982 : INV_X1 port map( I => n32531, ZN => n23032);
   U7994 : NAND2_X1 port map( A1 => n1286, A2 => n8801, ZN => n6712);
   U7996 : NOR2_X1 port map( A1 => n31561, A2 => n22637, ZN => n4511);
   U8001 : NAND2_X1 port map( A1 => n1842, A2 => n7659, ZN => n7658);
   U8006 : NOR2_X1 port map( A1 => n22025, A2 => n8131, ZN => n8349);
   U8025 : NAND2_X1 port map( A1 => n21957, A2 => n10724, ZN => n9547);
   U8033 : NAND2_X1 port map( A1 => n12488, A2 => n639, ZN => n10216);
   U8038 : NOR2_X1 port map( A1 => n3063, A2 => n22503, ZN => n3328);
   U8041 : AND2_X1 port map( A1 => n14251, A2 => n1294, Z => n1664);
   U8048 : NOR2_X1 port map( A1 => n22690, A2 => n22689, ZN => n3454);
   U8055 : OAI21_X1 port map( A1 => n26878, A2 => n27378, B => n12213, ZN => 
                           n7541);
   U8057 : INV_X1 port map( I => n16375, ZN => n22604);
   U8059 : NAND2_X1 port map( A1 => n901, A2 => n22524, ZN => n1727);
   U8067 : NOR2_X1 port map( A1 => n22645, A2 => n16166, ZN => n8595);
   U8069 : NAND2_X1 port map( A1 => n10282, A2 => n10354, ZN => n10355);
   U8073 : NOR2_X1 port map( A1 => n22625, A2 => n634, ZN => n7559);
   U8076 : INV_X1 port map( I => n11986, ZN => n9155);
   U8078 : BUF_X2 port map( I => n22504, Z => n3063);
   U8104 : INV_X1 port map( I => n22231, ZN => n10429);
   U8110 : INV_X2 port map( I => n21910, ZN => n1003);
   U8128 : AOI21_X1 port map( A1 => n32073, A2 => n1134, B => n13133, ZN => 
                           n21599);
   U8130 : NAND3_X1 port map( A1 => n1650, A2 => n21723, A3 => n28838, ZN => 
                           n1649);
   U8151 : NOR2_X1 port map( A1 => n727, A2 => n16441, ZN => n2443);
   U8158 : NOR2_X1 port map( A1 => n3043, A2 => n31197, ZN => n3042);
   U8161 : NOR2_X1 port map( A1 => n28581, A2 => n15302, ZN => n21657);
   U8168 : NOR2_X1 port map( A1 => n21489, A2 => n6718, ZN => n3418);
   U8175 : NOR2_X1 port map( A1 => n21738, A2 => n21866, ZN => n2625);
   U8178 : NAND2_X1 port map( A1 => n21235, A2 => n8029, ZN => n11381);
   U8182 : NOR2_X1 port map( A1 => n1136, A2 => n21581, ZN => n21164);
   U8186 : NAND2_X1 port map( A1 => n21461, A2 => n14640, ZN => n1650);
   U8227 : INV_X1 port map( I => n15022, ZN => n12587);
   U8255 : OAI22_X1 port map( A1 => n1784, A2 => n1632, B1 => n925, B2 => n1783
                           , ZN => n1457);
   U8262 : NOR2_X1 port map( A1 => n21451, A2 => n33498, ZN => n1968);
   U8267 : OR2_X1 port map( A1 => n21080, A2 => n17467, Z => n13968);
   U8268 : NAND2_X1 port map( A1 => n34131, A2 => n3236, ZN => n20941);
   U8274 : NAND2_X1 port map( A1 => n21393, A2 => n21367, ZN => n16311);
   U8280 : AOI22_X1 port map( A1 => n16505, A2 => n16473, B1 => n21152, B2 => 
                           n31835, ZN => n12689);
   U8292 : NOR2_X1 port map( A1 => n921, A2 => n21259, ZN => n3867);
   U8308 : NOR2_X1 port map( A1 => n21085, A2 => n26861, ZN => n1867);
   U8321 : NOR2_X1 port map( A1 => n1335, A2 => n14290, ZN => n20790);
   U8328 : OR3_X1 port map( A1 => n151, A2 => n21200, A3 => n17455, Z => n9794)
                           ;
   U8329 : INV_X1 port map( I => n7007, ZN => n2277);
   U8365 : INV_X1 port map( I => n20885, ZN => n5558);
   U8367 : OR2_X1 port map( A1 => n20954, A2 => n6158, Z => n6157);
   U8385 : NAND3_X1 port map( A1 => n20601, A2 => n28288, A3 => n12583, ZN => 
                           n2753);
   U8416 : OAI21_X1 port map( A1 => n28390, A2 => n20549, B => n12563, ZN => 
                           n11827);
   U8418 : OR2_X1 port map( A1 => n20487, A2 => n9808, Z => n11139);
   U8431 : NOR2_X1 port map( A1 => n31390, A2 => n13693, ZN => n11826);
   U8449 : NOR2_X1 port map( A1 => n1155, A2 => n30637, ZN => n11055);
   U8456 : NOR2_X1 port map( A1 => n32240, A2 => n20534, ZN => n11839);
   U8465 : OR2_X1 port map( A1 => n17947, A2 => n20485, Z => n5878);
   U8470 : AND2_X1 port map( A1 => n9688, A2 => n26881, Z => n9689);
   U8471 : NAND2_X1 port map( A1 => n8454, A2 => n4807, ZN => n20572);
   U8472 : NOR2_X1 port map( A1 => n15230, A2 => n28288, ZN => n5030);
   U8476 : AND2_X1 port map( A1 => n20570, A2 => n17236, Z => n12999);
   U8480 : NAND2_X1 port map( A1 => n1156, A2 => n20635, ZN => n2904);
   U8495 : NOR2_X1 port map( A1 => n33117, A2 => n30763, ZN => n3442);
   U8496 : INV_X1 port map( I => n11557, ZN => n12142);
   U8497 : NAND2_X1 port map( A1 => n5641, A2 => n32296, ZN => n5910);
   U8498 : NOR2_X1 port map( A1 => n17237, A2 => n17236, ZN => n5592);
   U8505 : NOR2_X1 port map( A1 => n937, A2 => n13077, ZN => n15849);
   U8506 : AND2_X1 port map( A1 => n19952, A2 => n14927, Z => n19953);
   U8510 : NAND2_X1 port map( A1 => n3197, A2 => n729, ZN => n1679);
   U8523 : NAND2_X1 port map( A1 => n2291, A2 => n2289, ZN => n2292);
   U8536 : NAND3_X1 port map( A1 => n13771, A2 => n12100, A3 => n9876, ZN => 
                           n1815);
   U8539 : NAND2_X1 port map( A1 => n821, A2 => n19884, ZN => n8382);
   U8540 : AOI21_X1 port map( A1 => n13605, A2 => n16493, B => n1161, ZN => 
                           n5693);
   U8542 : NAND2_X1 port map( A1 => n6263, A2 => n4674, ZN => n14011);
   U8545 : NOR2_X1 port map( A1 => n12179, A2 => n20156, ZN => n12178);
   U8553 : NAND2_X1 port map( A1 => n1438, A2 => n3790, ZN => n12351);
   U8555 : INV_X1 port map( I => n19935, ZN => n14171);
   U8556 : OAI21_X1 port map( A1 => n20128, A2 => n875, B => n431, ZN => n7893)
                           ;
   U8570 : NAND2_X1 port map( A1 => n26551, A2 => n19456, ZN => n5827);
   U8571 : NOR2_X1 port map( A1 => n12075, A2 => n20052, ZN => n7244);
   U8585 : NOR2_X1 port map( A1 => n11959, A2 => n9724, ZN => n9027);
   U8587 : NOR3_X1 port map( A1 => n20052, A2 => n584, A3 => n17495, ZN => 
                           n3769);
   U8588 : AND2_X1 port map( A1 => n17243, A2 => n4215, Z => n16029);
   U8593 : NOR2_X1 port map( A1 => n15189, A2 => n9724, ZN => n14793);
   U8609 : INV_X1 port map( I => n11219, ZN => n9263);
   U8610 : INV_X1 port map( I => n7108, ZN => n5606);
   U8613 : INV_X1 port map( I => n19589, ZN => n13095);
   U8614 : NAND2_X1 port map( A1 => n4592, A2 => n7810, ZN => n10073);
   U8617 : NAND2_X1 port map( A1 => n4405, A2 => n7680, ZN => n4592);
   U8635 : NAND2_X1 port map( A1 => n10943, A2 => n19284, ZN => n9383);
   U8656 : AND2_X1 port map( A1 => n14597, A2 => n8742, Z => n19336);
   U8657 : INV_X1 port map( I => n26600, ZN => n19202);
   U8659 : NOR2_X1 port map( A1 => n1386, A2 => n2935, ZN => n7201);
   U8663 : NOR2_X1 port map( A1 => n13806, A2 => n947, ZN => n6009);
   U8665 : NAND2_X1 port map( A1 => n2612, A2 => n19325, ZN => n16872);
   U8669 : NOR2_X1 port map( A1 => n877, A2 => n4202, ZN => n4218);
   U8671 : NAND2_X1 port map( A1 => n2101, A2 => n19269, ZN => n2100);
   U8678 : AND2_X1 port map( A1 => n34018, A2 => n3340, Z => n18935);
   U8686 : NOR2_X1 port map( A1 => n31108, A2 => n10017, ZN => n18908);
   U8687 : NAND2_X1 port map( A1 => n19252, A2 => n29757, ZN => n19176);
   U8689 : NOR2_X1 port map( A1 => n18983, A2 => n8233, ZN => n5636);
   U8693 : INV_X1 port map( I => n4436, ZN => n19175);
   U8695 : NOR2_X1 port map( A1 => n950, A2 => n19116, ZN => n19117);
   U8699 : INV_X1 port map( I => n19020, ZN => n13426);
   U8702 : NAND2_X1 port map( A1 => n4053, A2 => n5646, ZN => n5645);
   U8703 : INV_X1 port map( I => n25960, ZN => n19121);
   U8707 : INV_X1 port map( I => n13796, ZN => n19036);
   U8709 : NAND2_X1 port map( A1 => n30958, A2 => n31949, ZN => n4364);
   U8715 : INV_X1 port map( I => n19143, ZN => n19253);
   U8718 : AND2_X1 port map( A1 => n11203, A2 => n4016, Z => n10453);
   U8721 : NAND2_X1 port map( A1 => n8395, A2 => n6399, ZN => n12174);
   U8738 : NOR2_X1 port map( A1 => n11555, A2 => n18892, ZN => n6794);
   U8739 : NOR2_X1 port map( A1 => n28548, A2 => n12290, ZN => n15695);
   U8742 : INV_X1 port map( I => n18653, ZN => n9264);
   U8745 : OAI21_X1 port map( A1 => n18737, A2 => n6429, B => n6428, ZN => 
                           n18740);
   U8761 : OAI22_X1 port map( A1 => n6597, A2 => n18511, B1 => n956, B2 => 
                           n11380, ZN => n18513);
   U8762 : NOR2_X1 port map( A1 => n2733, A2 => n18893, ZN => n2732);
   U8765 : NAND2_X1 port map( A1 => n13548, A2 => n13514, ZN => n7518);
   U8766 : NAND2_X1 port map( A1 => n16403, A2 => n8395, ZN => n18366);
   U8768 : OAI21_X1 port map( A1 => n16435, A2 => n18602, B => n15115, ZN => 
                           n18292);
   U8771 : NAND2_X1 port map( A1 => n15406, A2 => n1184, ZN => n6173);
   U8780 : NAND2_X1 port map( A1 => n18739, A2 => n18863, ZN => n6428);
   U8783 : NOR2_X1 port map( A1 => n29315, A2 => n31971, ZN => n2596);
   U8784 : NAND2_X1 port map( A1 => n18101, A2 => n1189, ZN => n1571);
   U8785 : NOR2_X1 port map( A1 => n16181, A2 => n8208, ZN => n13243);
   U8789 : AOI21_X1 port map( A1 => n28344, A2 => n18808, B => n16474, ZN => 
                           n2432);
   U8790 : INV_X1 port map( I => n18812, ZN => n3180);
   U8794 : NOR2_X1 port map( A1 => n7899, A2 => n18797, ZN => n7681);
   U8796 : INV_X1 port map( I => n18569, ZN => n15070);
   U8797 : INV_X2 port map( I => n16766, ZN => n18642);
   U8799 : NAND2_X1 port map( A1 => n16487, A2 => n497, ZN => n6037);
   U8808 : OAI21_X1 port map( A1 => n29087, A2 => n171, B => n5473, ZN => 
                           n17737);
   U8810 : INV_X1 port map( I => n493, ZN => n1190);
   U8814 : NOR2_X1 port map( A1 => n12290, A2 => n962, ZN => n2964);
   U8818 : INV_X1 port map( I => n18548, ZN => n18808);
   U8826 : AND2_X1 port map( A1 => n1709, A2 => n961, Z => n8184);
   U8827 : CLKBUF_X2 port map( I => n18707, Z => n16487);
   U8828 : INV_X2 port map( I => n18888, ZN => n1060);
   U8831 : INV_X1 port map( I => n18823, ZN => n4869);
   U8832 : BUF_X2 port map( I => n18402, Z => n18849);
   U8833 : INV_X2 port map( I => n15240, ZN => n16855);
   U8834 : INV_X1 port map( I => n14926, ZN => n16370);
   U8836 : INV_X1 port map( I => n16355, ZN => n1191);
   U8839 : INV_X1 port map( I => n25190, ZN => n1197);
   U8840 : INV_X1 port map( I => n16575, ZN => n1196);
   U8841 : INV_X1 port map( I => n16685, ZN => n1194);
   U8842 : INV_X1 port map( I => n16612, ZN => n1192);
   U8843 : INV_X1 port map( I => n25373, ZN => n1193);
   U8846 : CLKBUF_X2 port map( I => Key(140), Z => n24966);
   U8847 : CLKBUF_X2 port map( I => Key(41), Z => n25751);
   U8848 : CLKBUF_X2 port map( I => Key(68), Z => n25648);
   U8849 : CLKBUF_X2 port map( I => Key(77), Z => n24917);
   U8851 : CLKBUF_X2 port map( I => Key(127), Z => n16685);
   U8854 : CLKBUF_X2 port map( I => Key(38), Z => n24953);
   U8856 : CLKBUF_X2 port map( I => Key(188), Z => n25191);
   U8865 : CLKBUF_X2 port map( I => Key(176), Z => n25126);
   U8868 : CLKBUF_X2 port map( I => Key(86), Z => n25161);
   U8870 : CLKBUF_X2 port map( I => Key(95), Z => n25519);
   U8872 : NOR2_X1 port map( A1 => n13624, A2 => n30557, ZN => n10012);
   U8873 : NAND3_X1 port map( A1 => n11005, A2 => n25819, A3 => n11004, ZN => 
                           n15959);
   U8876 : AOI22_X1 port map( A1 => n7270, A2 => n7271, B1 => n7274, B2 => 
                           n1395, ZN => n7266);
   U8881 : OAI21_X1 port map( A1 => n25510, A2 => n749, B => n1946, ZN => n1945
                           );
   U8885 : OAI21_X1 port map( A1 => n16833, A2 => n16973, B => n963, ZN => 
                           n6047);
   U8889 : OAI21_X1 port map( A1 => n25812, A2 => n25803, B => n25826, ZN => 
                           n11005);
   U8891 : AOI22_X1 port map( A1 => n10959, A2 => n25569, B1 => n5918, B2 => 
                           n5917, ZN => n5916);
   U8892 : NAND2_X1 port map( A1 => n7271, A2 => n7273, ZN => n7269);
   U8893 : NOR2_X1 port map( A1 => n3435, A2 => n786, ZN => n3434);
   U8899 : AOI22_X1 port map( A1 => n30318, A2 => n30288, B1 => n14737, B2 => 
                           n32059, ZN => n5303);
   U8900 : NAND2_X1 port map( A1 => n25193, A2 => n786, ZN => n13245);
   U8902 : NOR2_X1 port map( A1 => n32059, A2 => n2536, ZN => n7339);
   U8905 : NAND2_X1 port map( A1 => n25100, A2 => n1203, ZN => n7335);
   U8906 : OAI21_X1 port map( A1 => n9495, A2 => n13640, B => n6915, ZN => 
                           n9552);
   U8907 : OAI21_X1 port map( A1 => n6092, A2 => n25575, B => n25571, ZN => 
                           n3639);
   U8909 : NAND2_X1 port map( A1 => n11571, A2 => n25247, ZN => n11569);
   U8911 : NAND2_X1 port map( A1 => n25906, A2 => n1206, ZN => n7716);
   U8914 : NAND2_X1 port map( A1 => n10941, A2 => n15359, ZN => n10940);
   U8915 : NAND2_X1 port map( A1 => n27149, A2 => n4781, ZN => n25189);
   U8918 : INV_X1 port map( I => n17637, ZN => n8902);
   U8919 : NOR2_X1 port map( A1 => n25665, A2 => n25657, ZN => n6299);
   U8935 : NAND2_X1 port map( A1 => n25391, A2 => n11556, ZN => n6909);
   U8944 : NAND2_X1 port map( A1 => n13323, A2 => n11306, ZN => n5989);
   U8945 : NAND2_X1 port map( A1 => n24734, A2 => n24733, ZN => n24735);
   U8951 : AOI21_X1 port map( A1 => n16442, A2 => n9127, B => n11718, ZN => 
                           n24364);
   U8954 : NOR2_X1 port map( A1 => n25872, A2 => n25884, ZN => n9111);
   U8958 : NOR2_X1 port map( A1 => n9195, A2 => n24713, ZN => n24714);
   U8959 : NAND2_X1 port map( A1 => n5203, A2 => n25116, ZN => n3794);
   U8961 : NOR2_X1 port map( A1 => n3033, A2 => n17787, ZN => n2998);
   U8962 : NAND2_X1 port map( A1 => n24875, A2 => n14959, ZN => n5624);
   U8965 : NOR2_X1 port map( A1 => n5468, A2 => n25232, ZN => n5467);
   U8966 : INV_X1 port map( I => n11752, ZN => n25868);
   U8969 : NOR2_X1 port map( A1 => n18219, A2 => n25900, ZN => n14104);
   U8973 : NOR2_X1 port map( A1 => n25388, A2 => n25590, ZN => n10042);
   U8976 : NOR2_X1 port map( A1 => n790, A2 => n1223, ZN => n10548);
   U8979 : NAND2_X1 port map( A1 => n24729, A2 => n754, ZN => n8195);
   U8980 : NOR2_X1 port map( A1 => n25566, A2 => n16648, ZN => n10396);
   U8983 : OAI21_X1 port map( A1 => n16025, A2 => n25116, B => n25119, ZN => 
                           n24981);
   U8989 : NAND2_X1 port map( A1 => n25867, A2 => n1223, ZN => n17489);
   U8990 : INV_X1 port map( I => n25117, ZN => n12164);
   U8993 : NAND2_X1 port map( A1 => n6034, A2 => n12039, ZN => n25204);
   U8994 : AOI21_X1 port map( A1 => n4407, A2 => n17120, B => n25760, ZN => 
                           n2872);
   U8996 : AOI21_X1 port map( A1 => n25114, A2 => n560, B => n18154, ZN => 
                           n9957);
   U8998 : AND2_X1 port map( A1 => n25760, A2 => n754, Z => n13258);
   U9002 : AND2_X1 port map( A1 => n5254, A2 => n28455, Z => n12113);
   U9004 : NAND2_X1 port map( A1 => n837, A2 => n12042, ZN => n9859);
   U9008 : INV_X2 port map( I => n17867, ZN => n25382);
   U9012 : INV_X1 port map( I => n24770, ZN => n6862);
   U9013 : INV_X1 port map( I => n9681, ZN => n8215);
   U9016 : INV_X1 port map( I => n18028, ZN => n4244);
   U9017 : INV_X1 port map( I => n24622, ZN => n3294);
   U9018 : INV_X1 port map( I => n12313, ZN => n3305);
   U9021 : INV_X2 port map( I => n24548, ZN => n1084);
   U9039 : NAND2_X1 port map( A1 => n24140, A2 => n7203, ZN => n6166);
   U9047 : NOR2_X1 port map( A1 => n31862, A2 => n3181, ZN => n24129);
   U9052 : NAND2_X1 port map( A1 => n33680, A2 => n24242, ZN => n2325);
   U9054 : OAI21_X1 port map( A1 => n1237, A2 => n30061, B => n3548, ZN => 
                           n3547);
   U9058 : NAND3_X1 port map( A1 => n14530, A2 => n24223, A3 => n24042, ZN => 
                           n9965);
   U9061 : NOR2_X1 port map( A1 => n24236, A2 => n32102, ZN => n15271);
   U9067 : NOR2_X1 port map( A1 => n24159, A2 => n29748, ZN => n11435);
   U9071 : OR2_X1 port map( A1 => n719, A2 => n24073, Z => n11387);
   U9073 : NAND2_X1 port map( A1 => n1240, A2 => n13412, ZN => n7019);
   U9084 : OAI21_X1 port map( A1 => n24237, A2 => n14542, B => n32862, ZN => 
                           n15270);
   U9085 : AOI21_X1 port map( A1 => n2686, A2 => n13458, B => n24209, ZN => 
                           n6819);
   U9090 : OAI21_X1 port map( A1 => n26750, A2 => n8058, B => n23665, ZN => 
                           n23666);
   U9093 : INV_X1 port map( I => n24228, ZN => n13733);
   U9103 : NOR2_X1 port map( A1 => n15065, A2 => n24177, ZN => n13356);
   U9106 : NOR2_X1 port map( A1 => n24251, A2 => n28553, ZN => n3221);
   U9112 : NOR2_X1 port map( A1 => n14399, A2 => n16868, ZN => n3632);
   U9118 : AOI22_X1 port map( A1 => n23895, A2 => n23894, B1 => n28265, B2 => 
                           n707, ZN => n5754);
   U9127 : NAND2_X1 port map( A1 => n15207, A2 => n13720, ZN => n15206);
   U9153 : NAND2_X1 port map( A1 => n23632, A2 => n33337, ZN => n6467);
   U9157 : NOR2_X1 port map( A1 => n8145, A2 => n23912, ZN => n3446);
   U9159 : NAND2_X1 port map( A1 => n16271, A2 => n8547, ZN => n14038);
   U9167 : NAND2_X1 port map( A1 => n31435, A2 => n23847, ZN => n9329);
   U9168 : NAND2_X1 port map( A1 => n7077, A2 => n1253, ZN => n7076);
   U9183 : NOR2_X1 port map( A1 => n23860, A2 => n17661, ZN => n8865);
   U9184 : NAND2_X1 port map( A1 => n4891, A2 => n8525, ZN => n23952);
   U9200 : NOR2_X1 port map( A1 => n23857, A2 => n4177, ZN => n15186);
   U9201 : NOR2_X1 port map( A1 => n31890, A2 => n13521, ZN => n14496);
   U9204 : NOR2_X1 port map( A1 => n17694, A2 => n29246, ZN => n12031);
   U9207 : NAND2_X1 port map( A1 => n10955, A2 => n29246, ZN => n9740);
   U9226 : NAND3_X1 port map( A1 => n12823, A2 => n16587, A3 => n22874, ZN => 
                           n1671);
   U9227 : AOI21_X1 port map( A1 => n12823, A2 => n22874, B => n16587, ZN => 
                           n1673);
   U9234 : AOI21_X1 port map( A1 => n22893, A2 => n22894, B => n23034, ZN => 
                           n8150);
   U9248 : AOI21_X1 port map( A1 => n31861, A2 => n4113, B => n22915, ZN => 
                           n15717);
   U9259 : NAND2_X1 port map( A1 => n22972, A2 => n14420, ZN => n2639);
   U9263 : NOR2_X1 port map( A1 => n22862, A2 => n6800, ZN => n4609);
   U9264 : INV_X1 port map( I => n11018, ZN => n3348);
   U9270 : NAND2_X1 port map( A1 => n1112, A2 => n1267, ZN => n15831);
   U9272 : AOI21_X1 port map( A1 => n897, A2 => n15704, B => n15301, ZN => 
                           n2029);
   U9274 : OAI21_X1 port map( A1 => n11268, A2 => n641, B => n10031, ZN => 
                           n2032);
   U9276 : INV_X1 port map( I => n1267, ZN => n2773);
   U9278 : NAND3_X1 port map( A1 => n724, A2 => n13751, A3 => n23073, ZN => 
                           n3162);
   U9279 : NAND2_X1 port map( A1 => n10884, A2 => n723, ZN => n10883);
   U9280 : OAI21_X1 port map( A1 => n22962, A2 => n13592, B => n8334, ZN => 
                           n8127);
   U9297 : AND2_X1 port map( A1 => n15718, A2 => n27090, Z => n1719);
   U9300 : NAND2_X1 port map( A1 => n27798, A2 => n31867, ZN => n8201);
   U9302 : NOR2_X1 port map( A1 => n27719, A2 => n31325, ZN => n11828);
   U9312 : AND2_X1 port map( A1 => n22834, A2 => n10360, Z => n9384);
   U9314 : INV_X1 port map( I => n12687, ZN => n12686);
   U9315 : INV_X1 port map( I => n22871, ZN => n15389);
   U9326 : INV_X2 port map( I => n15243, ZN => n1109);
   U9328 : OAI21_X1 port map( A1 => n3502, A2 => n8260, B => n16483, ZN => 
                           n3501);
   U9331 : NAND3_X1 port map( A1 => n15204, A2 => n12530, A3 => n13710, ZN => 
                           n21883);
   U9335 : OAI21_X1 port map( A1 => n3329, A2 => n3328, B => n1287, ZN => n3327
                           );
   U9348 : AOI21_X1 port map( A1 => n22449, A2 => n2381, B => n22557, ZN => 
                           n2380);
   U9349 : OAI21_X1 port map( A1 => n11895, A2 => n28473, B => n14591, ZN => 
                           n14590);
   U9358 : NAND2_X1 port map( A1 => n16367, A2 => n22461, ZN => n16366);
   U9360 : AOI21_X1 port map( A1 => n22404, A2 => n12496, B => n3325, ZN => 
                           n3324);
   U9363 : NAND2_X1 port map( A1 => n11866, A2 => n29232, ZN => n11865);
   U9366 : NAND2_X1 port map( A1 => n22434, A2 => n28472, ZN => n13008);
   U9371 : INV_X1 port map( I => n22430, ZN => n22431);
   U9373 : NOR2_X1 port map( A1 => n22329, A2 => n10354, ZN => n9653);
   U9374 : NOR2_X1 port map( A1 => n31701, A2 => n10355, ZN => n6401);
   U9376 : NAND2_X1 port map( A1 => n8594, A2 => n4315, ZN => n8593);
   U9387 : NOR2_X1 port map( A1 => n907, A2 => n10206, ZN => n1820);
   U9394 : NOR2_X1 port map( A1 => n22544, A2 => n10288, ZN => n7237);
   U9401 : NAND2_X1 port map( A1 => n13485, A2 => n8318, ZN => n1658);
   U9403 : AOI21_X1 port map( A1 => n15195, A2 => n1296, B => n13169, ZN => 
                           n13168);
   U9404 : NOR2_X1 port map( A1 => n14376, A2 => n22672, ZN => n4810);
   U9407 : NAND2_X1 port map( A1 => n14307, A2 => n22576, ZN => n4547);
   U9422 : NOR2_X1 port map( A1 => n3063, A2 => n9370, ZN => n3332);
   U9425 : AND2_X1 port map( A1 => n17916, A2 => n1291, Z => n15740);
   U9427 : NAND3_X1 port map( A1 => n11244, A2 => n11629, A3 => n1296, ZN => 
                           n11243);
   U9431 : NAND2_X1 port map( A1 => n22540, A2 => n12844, ZN => n4504);
   U9439 : AND2_X1 port map( A1 => n12496, A2 => n3063, Z => n3329);
   U9443 : NOR2_X1 port map( A1 => n8318, A2 => n11244, ZN => n2137);
   U9450 : AND2_X1 port map( A1 => n16166, A2 => n22642, Z => n22643);
   U9452 : AOI21_X1 port map( A1 => n16166, A2 => n30641, B => n22645, ZN => 
                           n17191);
   U9453 : AND2_X1 port map( A1 => n16432, A2 => n8527, Z => n8529);
   U9458 : AND3_X1 port map( A1 => n22452, A2 => n16567, A3 => n22576, Z => 
                           n14219);
   U9476 : INV_X1 port map( I => n34160, ZN => n1970);
   U9490 : NOR2_X1 port map( A1 => n11796, A2 => n1647, ZN => n7326);
   U9495 : NAND3_X1 port map( A1 => n2551, A2 => n1647, A3 => n32282, ZN => 
                           n1651);
   U9504 : NAND2_X1 port map( A1 => n31910, A2 => n913, ZN => n7323);
   U9525 : NAND2_X1 port map( A1 => n21653, A2 => n21592, ZN => n21154);
   U9529 : NAND2_X1 port map( A1 => n11890, A2 => n21832, ZN => n2300);
   U9532 : NOR2_X1 port map( A1 => n21840, A2 => n4234, ZN => n21610);
   U9533 : INV_X1 port map( I => n21823, ZN => n8006);
   U9546 : NAND3_X1 port map( A1 => n21663, A2 => n777, A3 => n31197, ZN => 
                           n7949);
   U9549 : NAND2_X1 port map( A1 => n21664, A2 => n21662, ZN => n3049);
   U9551 : OR2_X1 port map( A1 => n27619, A2 => n15026, Z => n12448);
   U9559 : AND2_X1 port map( A1 => n21737, A2 => n30152, Z => n16371);
   U9560 : NAND2_X1 port map( A1 => n11683, A2 => n11215, ZN => n11682);
   U9564 : OAI21_X1 port map( A1 => n1328, A2 => n28181, B => n21460, ZN => 
                           n9284);
   U9567 : NAND2_X1 port map( A1 => n32642, A2 => n6489, ZN => n16735);
   U9570 : INV_X1 port map( I => n21697, ZN => n21656);
   U9573 : NAND2_X1 port map( A1 => n432, A2 => n16194, ZN => n6935);
   U9588 : NAND2_X1 port map( A1 => n11684, A2 => n29460, ZN => n11683);
   U9591 : NAND2_X1 port map( A1 => n26407, A2 => n28642, ZN => n11684);
   U9610 : NAND2_X1 port map( A1 => n29256, A2 => n16933, ZN => n17984);
   U9625 : INV_X1 port map( I => n21387, ZN => n6182);
   U9626 : NAND2_X1 port map( A1 => n12195, A2 => n20677, ZN => n1559);
   U9635 : AND2_X1 port map( A1 => n15506, A2 => n151, Z => n2724);
   U9636 : NOR2_X1 port map( A1 => n8657, A2 => n33454, ZN => n5730);
   U9645 : NAND2_X1 port map( A1 => n28257, A2 => n1022, ZN => n4088);
   U9656 : NOR2_X1 port map( A1 => n21269, A2 => n1017, ZN => n12865);
   U9659 : AND2_X1 port map( A1 => n21259, A2 => n21257, Z => n10096);
   U9667 : NAND2_X1 port map( A1 => n21149, A2 => n2738, ZN => n2716);
   U9668 : NAND2_X1 port map( A1 => n21389, A2 => n29901, ZN => n6181);
   U9675 : NAND2_X1 port map( A1 => n1332, A2 => n14483, ZN => n14482);
   U9679 : INV_X1 port map( I => n349, ZN => n21217);
   U9683 : OAI21_X1 port map( A1 => n11272, A2 => n510, B => n17455, ZN => 
                           n12091);
   U9684 : NAND2_X1 port map( A1 => n28737, A2 => n398, ZN => n5683);
   U9687 : NAND3_X1 port map( A1 => n927, A2 => n21441, A3 => n926, ZN => n2664
                           );
   U9692 : NAND2_X1 port map( A1 => n8605, A2 => n10558, ZN => n8604);
   U9695 : NAND2_X1 port map( A1 => n21215, A2 => n12525, ZN => n21216);
   U9696 : INV_X1 port map( I => n21263, ZN => n21057);
   U9706 : NAND2_X1 port map( A1 => n21448, A2 => n5822, ZN => n21449);
   U9709 : INV_X1 port map( I => n30313, ZN => n21084);
   U9722 : AOI22_X1 port map( A1 => n4618, A2 => n1398, B1 => n4617, B2 => 
                           n4616, ZN => n10110);
   U9725 : INV_X1 port map( I => n20711, ZN => n8343);
   U9726 : NOR2_X1 port map( A1 => n18265, A2 => n1398, ZN => n4617);
   U9737 : NOR2_X1 port map( A1 => n13572, A2 => n11634, ZN => n8579);
   U9752 : NOR2_X1 port map( A1 => n20338, A2 => n20590, ZN => n20592);
   U9755 : INV_X1 port map( I => n14858, ZN => n1828);
   U9756 : NAND2_X1 port map( A1 => n5496, A2 => n8268, ZN => n5350);
   U9760 : NAND2_X1 port map( A1 => n4807, A2 => n816, ZN => n8820);
   U9783 : AND2_X1 port map( A1 => n9783, A2 => n31873, Z => n10488);
   U9787 : NAND2_X1 port map( A1 => n26041, A2 => n20523, ZN => n15257);
   U9789 : NOR2_X1 port map( A1 => n3443, A2 => n3442, ZN => n3441);
   U9790 : NAND3_X1 port map( A1 => n20313, A2 => n20314, A3 => n20481, ZN => 
                           n20315);
   U9795 : NAND2_X1 port map( A1 => n20525, A2 => n12169, ZN => n9485);
   U9799 : NAND2_X1 port map( A1 => n16190, A2 => n16144, ZN => n2621);
   U9801 : NAND2_X1 port map( A1 => n20377, A2 => n14179, ZN => n5497);
   U9808 : NAND2_X1 port map( A1 => n1350, A2 => n14545, ZN => n3425);
   U9809 : OAI21_X1 port map( A1 => n16518, A2 => n20533, B => n15027, ZN => 
                           n11038);
   U9817 : NOR2_X1 port map( A1 => n20570, A2 => n31968, ZN => n12793);
   U9832 : NOR2_X1 port map( A1 => n819, A2 => n11988, ZN => n5026);
   U9848 : NOR2_X1 port map( A1 => n6864, A2 => n10752, ZN => n7308);
   U9849 : NAND2_X1 port map( A1 => n8382, A2 => n11593, ZN => n2147);
   U9850 : NOR2_X1 port map( A1 => n19921, A2 => n33525, ZN => n7631);
   U9853 : OAI21_X1 port map( A1 => n29003, A2 => n31742, B => n15135, ZN => 
                           n7551);
   U9868 : OR2_X1 port map( A1 => n19883, A2 => n19794, Z => n17944);
   U9869 : NOR2_X1 port map( A1 => n28600, A2 => n19975, ZN => n1898);
   U9879 : NOR2_X1 port map( A1 => n10752, A2 => n19921, ZN => n19922);
   U9888 : NOR2_X1 port map( A1 => n19459, A2 => n7609, ZN => n7607);
   U9893 : INV_X1 port map( I => n13859, ZN => n9221);
   U9895 : NOR2_X1 port map( A1 => n12168, A2 => n16848, ZN => n5718);
   U9901 : NAND2_X1 port map( A1 => n20120, A2 => n14815, ZN => n6221);
   U9909 : AOI21_X1 port map( A1 => n9563, A2 => n8100, B => n17967, ZN => 
                           n3270);
   U9917 : OR3_X1 port map( A1 => n17260, A2 => n28600, A3 => n873, Z => n15176
                           );
   U9923 : INV_X1 port map( I => n13605, ZN => n11119);
   U9924 : NAND2_X1 port map( A1 => n34154, A2 => n29153, ZN => n15602);
   U9927 : NOR2_X1 port map( A1 => n12038, A2 => n11913, ZN => n10804);
   U9929 : AND2_X1 port map( A1 => n942, A2 => n15110, Z => n9302);
   U9931 : INV_X1 port map( I => n15237, ZN => n20138);
   U9935 : OR2_X1 port map( A1 => n397, A2 => n14210, Z => n6409);
   U9939 : INV_X1 port map( I => n20119, ZN => n20018);
   U9947 : INV_X1 port map( I => n20098, ZN => n19891);
   U9956 : INV_X1 port map( I => n15236, ZN => n4976);
   U9958 : INV_X1 port map( I => n3652, ZN => n3194);
   U9963 : INV_X1 port map( I => n11102, ZN => n1365);
   U9964 : INV_X1 port map( I => n17430, ZN => n5484);
   U9974 : NAND2_X1 port map( A1 => n9383, A2 => n1376, ZN => n3206);
   U9979 : OAI21_X1 port map( A1 => n18935, A2 => n1386, B => n7133, ZN => 
                           n1655);
   U9981 : NAND2_X1 port map( A1 => n8437, A2 => n33672, ZN => n5222);
   U9983 : NOR2_X1 port map( A1 => n2100, A2 => n2098, ZN => n19073);
   U9996 : NAND2_X1 port map( A1 => n14331, A2 => n4436, ZN => n2587);
   U10004 : AOI21_X1 port map( A1 => n19334, A2 => n8212, B => n12815, ZN => 
                           n6440);
   U10007 : NAND2_X1 port map( A1 => n12502, A2 => n7557, ZN => n6577);
   U10008 : NOR2_X1 port map( A1 => n25999, A2 => n5636, ZN => n5635);
   U10011 : AOI22_X1 port map( A1 => n19182, A2 => n19181, B1 => n33078, B2 => 
                           n29769, ZN => n2125);
   U10013 : NOR2_X1 port map( A1 => n2283, A2 => n3340, ZN => n6779);
   U10016 : AND2_X1 port map( A1 => n19186, A2 => n947, Z => n15675);
   U10018 : OAI22_X1 port map( A1 => n17386, A2 => n19096, B1 => n29093, B2 => 
                           n10203, ZN => n3115);
   U10019 : NAND2_X1 port map( A1 => n31451, A2 => n5889, ZN => n7187);
   U10020 : OR2_X1 port map( A1 => n33845, A2 => n10260, Z => n14113);
   U10021 : AND2_X1 port map( A1 => n1386, A2 => n31139, Z => n7200);
   U10022 : NAND2_X1 port map( A1 => n15021, A2 => n1384, ZN => n7901);
   U10024 : NAND2_X1 port map( A1 => n13568, A2 => n824, ZN => n9177);
   U10026 : NAND2_X1 port map( A1 => n19110, A2 => n17725, ZN => n6563);
   U10028 : OAI21_X1 port map( A1 => n19334, A2 => n9538, B => n8742, ZN => 
                           n6282);
   U10030 : INV_X1 port map( I => n18454, ZN => n18285);
   U10032 : NAND2_X1 port map( A1 => n17817, A2 => n10124, ZN => n3360);
   U10034 : INV_X1 port map( I => n16790, ZN => n2871);
   U10039 : NAND2_X1 port map( A1 => n27807, A2 => n6290, ZN => n11262);
   U10042 : OAI21_X1 port map( A1 => n9423, A2 => n19229, B => n34107, ZN => 
                           n18440);
   U10046 : OAI22_X1 port map( A1 => n5877, A2 => n19199, B1 => n29047, B2 => 
                           n5876, ZN => n18789);
   U10047 : INV_X1 port map( I => n5789, ZN => n19209);
   U10048 : NOR2_X1 port map( A1 => n9423, A2 => n19357, ZN => n16769);
   U10049 : AND2_X1 port map( A1 => n19262, A2 => n25971, Z => n18751);
   U10051 : AOI21_X1 port map( A1 => n25985, A2 => n33822, B => n19146, ZN => 
                           n10259);
   U10054 : NAND2_X1 port map( A1 => n7134, A2 => n19002, ZN => n5033);
   U10060 : NAND3_X1 port map( A1 => n4365, A2 => n4364, A3 => n5789, ZN => 
                           n4363);
   U10064 : NAND2_X1 port map( A1 => n5545, A2 => n19360, ZN => n18931);
   U10067 : AOI21_X1 port map( A1 => n1053, A2 => n19109, B => n19107, ZN => 
                           n19111);
   U10068 : NAND2_X1 port map( A1 => n19088, A2 => n19087, ZN => n7435);
   U10069 : AND3_X1 port map( A1 => n19216, A2 => n32805, A3 => n827, Z => 
                           n6575);
   U10072 : AOI21_X1 port map( A1 => n1054, A2 => n13796, B => n11940, ZN => 
                           n1836);
   U10073 : INV_X1 port map( I => n32788, ZN => n18474);
   U10074 : NAND2_X1 port map( A1 => n2901, A2 => n2902, ZN => n19214);
   U10081 : NOR2_X1 port map( A1 => n19257, A2 => n25971, ZN => n4596);
   U10082 : INV_X1 port map( I => n4835, ZN => n14806);
   U10097 : NAND2_X1 port map( A1 => n8376, A2 => n7454, ZN => n3364);
   U10099 : NAND2_X1 port map( A1 => n18682, A2 => n746, ZN => n7275);
   U10100 : NOR2_X1 port map( A1 => n14614, A2 => n18407, ZN => n10207);
   U10101 : NAND2_X1 port map( A1 => n18653, A2 => n9266, ZN => n9265);
   U10105 : NAND2_X1 port map( A1 => n16854, A2 => n16855, ZN => n3437);
   U10108 : NOR2_X1 port map( A1 => n7163, A2 => n7216, ZN => n7162);
   U10109 : NAND2_X1 port map( A1 => n18311, A2 => n6173, ZN => n6172);
   U10115 : NAND2_X1 port map( A1 => n15211, A2 => n18854, ZN => n3928);
   U10118 : NOR2_X1 port map( A1 => n1571, A2 => n16538, ZN => n14659);
   U10124 : NAND2_X1 port map( A1 => n9437, A2 => n2936, ZN => n14654);
   U10134 : NOR2_X1 port map( A1 => n14695, A2 => n18875, ZN => n14694);
   U10135 : NAND2_X1 port map( A1 => n18881, A2 => n18880, ZN => n9266);
   U10136 : NAND2_X1 port map( A1 => n16995, A2 => n18539, ZN => n14326);
   U10146 : OAI21_X1 port map( A1 => n1709, A2 => n10181, B => n11460, ZN => 
                           n18686);
   U10148 : NOR2_X1 port map( A1 => n14093, A2 => n18761, ZN => n18336);
   U10149 : OR2_X1 port map( A1 => n14906, A2 => n18511, Z => n6918);
   U10150 : OR2_X1 port map( A1 => n18566, A2 => n18492, Z => n14678);
   U10152 : NAND2_X1 port map( A1 => n18406, A2 => n18875, ZN => n9401);
   U10155 : NAND3_X1 port map( A1 => n3251, A2 => n18822, A3 => n29514, ZN => 
                           n15957);
   U10156 : OR2_X1 port map( A1 => n18463, A2 => n16915, Z => n11954);
   U10157 : AOI21_X1 port map( A1 => n18708, A2 => n18742, B => n10665, ZN => 
                           n17625);
   U10159 : NAND2_X1 port map( A1 => n18854, A2 => n18307, ZN => n18718);
   U10160 : NAND2_X1 port map( A1 => n18856, A2 => n18853, ZN => n3927);
   U10161 : NOR2_X1 port map( A1 => n11097, A2 => n18085, ZN => n11098);
   U10163 : NAND2_X1 port map( A1 => n8739, A2 => n30371, ZN => n6587);
   U10164 : AND2_X1 port map( A1 => n34139, A2 => n18492, Z => n18460);
   U10167 : OR2_X1 port map( A1 => n18539, A2 => n14651, Z => n2936);
   U10174 : BUF_X2 port map( I => n15265, Z => n7454);
   U10175 : AND2_X1 port map( A1 => n18770, A2 => n18774, Z => n18274);
   U10181 : NOR2_X1 port map( A1 => n18637, A2 => n18537, ZN => n13381);
   U10186 : INV_X1 port map( I => n17419, ZN => n11122);
   U10188 : INV_X1 port map( I => n16462, ZN => n9729);
   U10191 : INV_X1 port map( I => n25879, ZN => n1395);
   U10193 : INV_X1 port map( I => n16657, ZN => n1427);
   U10196 : INV_X2 port map( I => n12166, ZN => n18588);
   U10197 : INV_X1 port map( I => n25036, ZN => n1398);
   U10199 : INV_X1 port map( I => n24999, ZN => n1415);
   U10200 : INV_X1 port map( I => n25252, ZN => n1424);
   U10201 : CLKBUF_X2 port map( I => n32034, Z => n1446);
   U10206 : INV_X1 port map( I => n25156, ZN => n1393);
   U10207 : INV_X1 port map( I => n16497, ZN => n1396);
   U10209 : INV_X1 port map( I => n24707, ZN => n1407);
   U10210 : INV_X1 port map( I => n25167, ZN => n1413);
   U10211 : INV_X1 port map( I => n25772, ZN => n1431);
   U10212 : INV_X1 port map( I => n24992, ZN => n1406);
   U10217 : CLKBUF_X2 port map( I => Key(155), Z => n24738);
   U10219 : CLKBUF_X2 port map( I => Key(153), Z => n16666);
   U10220 : CLKBUF_X2 port map( I => Key(171), Z => n16622);
   U10221 : CLKBUF_X2 port map( I => Key(146), Z => n25549);
   U10224 : CLKBUF_X2 port map( I => Key(118), Z => n25319);
   U10225 : CLKBUF_X2 port map( I => Key(150), Z => n16520);
   U10226 : CLKBUF_X2 port map( I => Key(119), Z => n25669);
   U10227 : CLKBUF_X2 port map( I => Key(83), Z => n25457);
   U10228 : CLKBUF_X2 port map( I => Key(56), Z => n24374);
   U10230 : CLKBUF_X2 port map( I => Key(152), Z => n25001);
   U10233 : CLKBUF_X2 port map( I => Key(5), Z => n25560);
   U10234 : CLKBUF_X2 port map( I => Key(117), Z => n25079);
   U10236 : CLKBUF_X2 port map( I => Key(44), Z => n25506);
   U10237 : CLKBUF_X2 port map( I => Key(23), Z => n24895);
   U10238 : CLKBUF_X2 port map( I => Key(128), Z => n24923);
   U10239 : CLKBUF_X2 port map( I => Key(53), Z => n25827);
   U10241 : CLKBUF_X2 port map( I => Key(74), Z => n25098);
   U10242 : CLKBUF_X2 port map( I => Key(50), Z => n24992);
   U10243 : CLKBUF_X2 port map( I => Key(25), Z => n16687);
   U10245 : CLKBUF_X2 port map( I => Key(8), Z => n25252);
   U10246 : INV_X1 port map( I => n25641, ZN => n1198);
   U10249 : CLKBUF_X2 port map( I => Key(71), Z => n25324);
   U10250 : CLKBUF_X2 port map( I => Key(62), Z => n25040);
   U10255 : CLKBUF_X2 port map( I => Key(149), Z => n25224);
   U10267 : AOI21_X1 port map( A1 => n3706, A2 => n3434, B => n3432, ZN => 
                           n3431);
   U10268 : INV_X1 port map( I => n7303, ZN => n5622);
   U10278 : OAI22_X1 port map( A1 => n4642, A2 => n832, B1 => n25743, B2 => 
                           n1979, ZN => n24434);
   U10279 : NAND2_X1 port map( A1 => n25173, A2 => n25174, ZN => n8339);
   U10281 : OAI21_X1 port map( A1 => n5113, A2 => n7831, B => n14321, ZN => 
                           n14320);
   U10285 : NAND2_X1 port map( A1 => n2129, A2 => n13935, ZN => n2128);
   U10287 : NAND2_X1 port map( A1 => n24934, A2 => n24925, ZN => n5773);
   U10292 : OAI21_X1 port map( A1 => n24967, A2 => n24970, B => n3843, ZN => 
                           n3135);
   U10294 : NAND2_X1 port map( A1 => n25681, A2 => n26447, ZN => n1757);
   U10296 : NAND2_X1 port map( A1 => n25691, A2 => n25689, ZN => n1758);
   U10298 : INV_X1 port map( I => n24972, ZN => n2103);
   U10299 : NAND2_X1 port map( A1 => n3376, A2 => n14208, ZN => n5900);
   U10301 : NAND2_X1 port map( A1 => n25650, A2 => n6299, ZN => n7084);
   U10302 : NAND2_X1 port map( A1 => n11428, A2 => n965, ZN => n15250);
   U10304 : NAND2_X1 port map( A1 => n24967, A2 => n33434, ZN => n3846);
   U10310 : INV_X1 port map( I => n24913, ZN => n10214);
   U10312 : NAND2_X1 port map( A1 => n32859, A2 => n5712, ZN => n5520);
   U10318 : INV_X1 port map( I => n25067, ZN => n5865);
   U10324 : OAI21_X1 port map( A1 => n3123, A2 => n3122, B => n31640, ZN => 
                           n6424);
   U10325 : OR3_X1 port map( A1 => n25670, A2 => n25687, A3 => n25686, Z => 
                           n24860);
   U10328 : NAND2_X1 port map( A1 => n25222, A2 => n28651, ZN => n5638);
   U10332 : NOR2_X1 port map( A1 => n27183, A2 => n1074, ZN => n9732);
   U10335 : NAND2_X1 port map( A1 => n13023, A2 => n29243, ZN => n12217);
   U10336 : INV_X1 port map( I => n25851, ZN => n25860);
   U10338 : NOR2_X1 port map( A1 => n25171, A2 => n18227, ZN => n8930);
   U10340 : NOR2_X1 port map( A1 => n2049, A2 => n25686, ZN => n8156);
   U10341 : NOR2_X1 port map( A1 => n25059, A2 => n25060, ZN => n8257);
   U10342 : INV_X1 port map( I => n14732, ZN => n2017);
   U10349 : INV_X1 port map( I => n27162, ZN => n18022);
   U10352 : NAND2_X1 port map( A1 => n2536, A2 => n10469, ZN => n5408);
   U10355 : INV_X2 port map( I => n3019, ZN => n3232);
   U10358 : INV_X1 port map( I => n17488, ZN => n11247);
   U10359 : INV_X1 port map( I => n2191, ZN => n25257);
   U10361 : OAI21_X1 port map( A1 => n28136, A2 => n25391, B => n6909, ZN => 
                           n24587);
   U10363 : INV_X1 port map( I => n25172, ZN => n18227);
   U10370 : INV_X1 port map( I => n28736, ZN => n8073);
   U10373 : NAND2_X1 port map( A1 => n15894, A2 => n11703, ZN => n15771);
   U10393 : AND2_X1 port map( A1 => n15964, A2 => n25590, Z => n12025);
   U10399 : NAND2_X1 port map( A1 => n29476, A2 => n13322, ZN => n5990);
   U10400 : NAND2_X1 port map( A1 => n5467, A2 => n17110, ZN => n2214);
   U10402 : NOR2_X1 port map( A1 => n25839, A2 => n7143, ZN => n25840);
   U10403 : NOR2_X1 port map( A1 => n10396, A2 => n10395, ZN => n13422);
   U10404 : NAND2_X1 port map( A1 => n15770, A2 => n32798, ZN => n15894);
   U10408 : INV_X1 port map( I => n24718, ZN => n12369);
   U10417 : NOR2_X1 port map( A1 => n25761, A2 => n4407, ZN => n4531);
   U10420 : NAND2_X1 port map( A1 => n24448, A2 => n27127, ZN => n11697);
   U10423 : OAI21_X1 port map( A1 => n7064, A2 => n24714, B => n25763, ZN => 
                           n24717);
   U10430 : NAND2_X1 port map( A1 => n1081, A2 => n13429, ZN => n25010);
   U10432 : OR2_X1 port map( A1 => n1786, A2 => n13709, Z => n7855);
   U10434 : NOR2_X1 port map( A1 => n752, A2 => n25299, ZN => n10251);
   U10441 : NAND2_X1 port map( A1 => n24981, A2 => n25114, ZN => n3378);
   U10442 : NAND2_X1 port map( A1 => n25326, A2 => n15528, ZN => n6144);
   U10447 : INV_X1 port map( I => n4491, ZN => n25761);
   U10455 : NAND2_X1 port map( A1 => n24732, A2 => n13349, ZN => n12968);
   U10462 : OAI21_X1 port map( A1 => n17120, A2 => n25712, B => n2872, ZN => 
                           n2961);
   U10469 : AND2_X1 port map( A1 => n13709, A2 => n25201, Z => n25202);
   U10471 : OR2_X1 port map( A1 => n25891, A2 => n25892, Z => n12359);
   U10472 : OR2_X1 port map( A1 => n25584, A2 => n718, Z => n25585);
   U10473 : NOR2_X1 port map( A1 => n886, A2 => n15528, ZN => n10252);
   U10475 : NAND2_X1 port map( A1 => n31945, A2 => n25590, ZN => n11992);
   U10480 : NAND2_X1 port map( A1 => n754, A2 => n24729, ZN => n4452);
   U10481 : AND2_X1 port map( A1 => n13050, A2 => n13042, Z => n11976);
   U10486 : INV_X1 port map( I => n11973, ZN => n25709);
   U10488 : INV_X2 port map( I => n675, ZN => n1218);
   U10492 : INV_X4 port map( I => n24466, ZN => n1221);
   U10498 : INV_X1 port map( I => n24575, ZN => n17153);
   U10499 : INV_X1 port map( I => n17448, ZN => n24845);
   U10500 : INV_X1 port map( I => n24518, ZN => n13145);
   U10507 : INV_X1 port map( I => n24544, ZN => n4566);
   U10511 : INV_X1 port map( I => n24773, ZN => n17865);
   U10512 : INV_X1 port map( I => n24813, ZN => n11537);
   U10516 : INV_X1 port map( I => n15508, ZN => n8507);
   U10518 : INV_X1 port map( I => n24545, ZN => n10257);
   U10524 : AND2_X1 port map( A1 => n24166, A2 => n24165, Z => n6051);
   U10528 : NAND2_X1 port map( A1 => n3767, A2 => n3506, ZN => n6268);
   U10533 : INV_X1 port map( I => n4728, ZN => n8895);
   U10534 : NAND2_X1 port map( A1 => n23994, A2 => n28691, ZN => n11440);
   U10541 : INV_X2 port map( I => n283, ZN => n1228);
   U10549 : NAND2_X1 port map( A1 => n12068, A2 => n16090, ZN => n18128);
   U10569 : NOR2_X1 port map( A1 => n13047, A2 => n15253, ZN => n7101);
   U10573 : NAND2_X1 port map( A1 => n24336, A2 => n33680, ZN => n2400);
   U10577 : OR2_X1 port map( A1 => n24005, A2 => n1089, Z => n5424);
   U10578 : INV_X1 port map( I => n17112, ZN => n12353);
   U10581 : INV_X1 port map( I => n14530, ZN => n13082);
   U10583 : NAND2_X1 port map( A1 => n13748, A2 => n11346, ZN => n10450);
   U10594 : NAND2_X1 port map( A1 => n23666, A2 => n32459, ZN => n7883);
   U10601 : NAND2_X1 port map( A1 => n16574, A2 => n9323, ZN => n3549);
   U10607 : NOR2_X1 port map( A1 => n15271, A2 => n15270, ZN => n24238);
   U10608 : NOR2_X1 port map( A1 => n1096, A2 => n1800, ZN => n14411);
   U10610 : INV_X1 port map( I => n6819, ZN => n6818);
   U10613 : AND2_X1 port map( A1 => n24138, A2 => n3880, Z => n24140);
   U10614 : NOR2_X1 port map( A1 => n10342, A2 => n1093, ZN => n8399);
   U10619 : NAND2_X1 port map( A1 => n2944, A2 => n13268, ZN => n2943);
   U10620 : AND3_X1 port map( A1 => n24305, A2 => n12903, A3 => n24304, Z => 
                           n24306);
   U10623 : INV_X1 port map( I => n2686, ZN => n2945);
   U10636 : NAND2_X1 port map( A1 => n32041, A2 => n795, ZN => n11725);
   U10639 : NAND2_X1 port map( A1 => n24321, A2 => n8, ZN => n6841);
   U10645 : NAND3_X1 port map( A1 => n793, A2 => n27168, A3 => n13334, ZN => 
                           n1838);
   U10646 : NAND2_X1 port map( A1 => n15011, A2 => n24084, ZN => n24085);
   U10654 : OR2_X1 port map( A1 => n24210, A2 => n13530, Z => n11963);
   U10658 : INV_X1 port map( I => n1090, ZN => n1238);
   U10659 : INV_X1 port map( I => n24148, ZN => n24121);
   U10662 : NAND4_X1 port map( A1 => n4822, A2 => n4824, A3 => n4823, A4 => 
                           n4821, ZN => n24256);
   U10663 : AND2_X1 port map( A1 => n12997, A2 => n14907, Z => n4775);
   U10687 : NAND2_X1 port map( A1 => n5116, A2 => n13666, ZN => n11079);
   U10691 : NAND2_X1 port map( A1 => n13906, A2 => n13904, ZN => n12237);
   U10700 : INV_X1 port map( I => n15474, ZN => n5633);
   U10705 : AND2_X1 port map( A1 => n16786, A2 => n23692, Z => n8613);
   U10708 : NAND2_X1 port map( A1 => n23875, A2 => n26882, ZN => n16326);
   U10710 : NAND2_X1 port map( A1 => n662, A2 => n23938, ZN => n12080);
   U10712 : INV_X1 port map( I => n10069, ZN => n2447);
   U10715 : NAND2_X1 port map( A1 => n14164, A2 => n11095, ZN => n12884);
   U10729 : NAND2_X1 port map( A1 => n3873, A2 => n29839, ZN => n3744);
   U10733 : NAND2_X1 port map( A1 => n14088, A2 => n842, ZN => n8344);
   U10734 : NAND2_X1 port map( A1 => n12069, A2 => n14207, ZN => n11310);
   U10737 : NAND2_X1 port map( A1 => n23642, A2 => n4891, ZN => n3757);
   U10738 : NAND2_X1 port map( A1 => n12031, A2 => n548, ZN => n3708);
   U10740 : NOR2_X1 port map( A1 => n13103, A2 => n15446, ZN => n8064);
   U10765 : NAND2_X1 port map( A1 => n8865, A2 => n11904, ZN => n2003);
   U10767 : NAND2_X1 port map( A1 => n10140, A2 => n844, ZN => n9931);
   U10770 : NAND2_X1 port map( A1 => n33345, A2 => n844, ZN => n8655);
   U10771 : NOR2_X1 port map( A1 => n23637, A2 => n3650, ZN => n11653);
   U10776 : NOR2_X1 port map( A1 => n23868, A2 => n17895, ZN => n13137);
   U10781 : OR2_X1 port map( A1 => n23862, A2 => n23527, Z => n4079);
   U10783 : INV_X1 port map( I => n16033, ZN => n11157);
   U10785 : AND2_X1 port map( A1 => n16320, A2 => n977, Z => n12069);
   U10794 : INV_X1 port map( I => n23738, ZN => n14155);
   U10798 : AND2_X1 port map( A1 => n15682, A2 => n14325, Z => n11975);
   U10800 : NAND3_X1 port map( A1 => n1489, A2 => n23763, A3 => n23736, ZN => 
                           n23737);
   U10806 : NOR2_X1 port map( A1 => n757, A2 => n11887, ZN => n10068);
   U10808 : INV_X1 port map( I => n13342, ZN => n9444);
   U10811 : NAND2_X1 port map( A1 => n23902, A2 => n27474, ZN => n23176);
   U10814 : AND2_X1 port map( A1 => n23848, A2 => n23807, Z => n13544);
   U10821 : INV_X1 port map( I => n9391, ZN => n3375);
   U10830 : NAND2_X1 port map( A1 => n14585, A2 => n23763, ZN => n23723);
   U10837 : CLKBUF_X2 port map( I => n23435, Z => n8298);
   U10842 : INV_X1 port map( I => n12538, ZN => n23298);
   U10843 : INV_X1 port map( I => n23386, ZN => n9671);
   U10848 : INV_X1 port map( I => n10535, ZN => n4409);
   U10850 : INV_X1 port map( I => n1673, ZN => n1672);
   U10856 : INV_X1 port map( I => n23294, ZN => n7520);
   U10858 : INV_X1 port map( I => n30321, ZN => n23320);
   U10861 : INV_X1 port map( I => n23387, ZN => n5514);
   U10863 : INV_X1 port map( I => n12491, ZN => n11426);
   U10868 : INV_X1 port map( I => n4399, ZN => n22811);
   U10894 : NAND2_X1 port map( A1 => n12135, A2 => n4731, ZN => n4730);
   U10900 : NAND2_X1 port map( A1 => n2639, A2 => n2638, ZN => n2637);
   U10909 : INV_X1 port map( I => n5971, ZN => n2633);
   U10912 : NAND2_X1 port map( A1 => n23030, A2 => n13066, ZN => n14617);
   U10915 : NAND2_X1 port map( A1 => n2624, A2 => n23103, ZN => n2623);
   U10921 : NAND2_X1 port map( A1 => n22399, A2 => n12375, ZN => n3770);
   U10929 : AND2_X1 port map( A1 => n12417, A2 => n12418, Z => n12099);
   U10931 : OAI21_X1 port map( A1 => n12016, A2 => n14114, B => n31784, ZN => 
                           n3513);
   U10932 : NOR2_X1 port map( A1 => n23015, A2 => n27652, ZN => n13288);
   U10944 : NAND2_X1 port map( A1 => n11829, A2 => n11828, ZN => n11837);
   U10947 : NOR2_X1 port map( A1 => n22897, A2 => n27984, ZN => n16142);
   U10958 : NAND2_X1 port map( A1 => n13838, A2 => n4833, ZN => n13837);
   U10965 : INV_X1 port map( I => n22961, ZN => n5260);
   U10976 : AND2_X1 port map( A1 => n23003, A2 => n23000, Z => n12135);
   U10982 : AND2_X1 port map( A1 => n32119, A2 => n33675, Z => n23090);
   U10984 : NAND2_X1 port map( A1 => n12218, A2 => n990, ZN => n12180);
   U10989 : AND2_X1 port map( A1 => n3891, A2 => n22836, Z => n12033);
   U10990 : INV_X1 port map( I => n3614, ZN => n5981);
   U10992 : INV_X1 port map( I => n22800, ZN => n22801);
   U10994 : NAND2_X1 port map( A1 => n852, A2 => n8967, ZN => n8966);
   U10998 : INV_X1 port map( I => n9184, ZN => n6098);
   U11004 : AOI21_X1 port map( A1 => n17503, A2 => n31943, B => n22753, ZN => 
                           n17502);
   U11012 : NAND2_X1 port map( A1 => n22592, A2 => n22705, ZN => n11829);
   U11013 : NOR2_X1 port map( A1 => n990, A2 => n30297, ZN => n7747);
   U11015 : NAND3_X1 port map( A1 => n23079, A2 => n23082, A3 => n22885, ZN => 
                           n12646);
   U11024 : INV_X1 port map( I => n11330, ZN => n7745);
   U11029 : INV_X1 port map( I => n3566, ZN => n10166);
   U11030 : INV_X2 port map( I => n3668, ZN => n23026);
   U11031 : AND2_X1 port map( A1 => n23009, A2 => n23008, Z => n23010);
   U11033 : NAND2_X1 port map( A1 => n22900, A2 => n17211, ZN => n11048);
   U11037 : AND4_X1 port map( A1 => n22358, A2 => n17627, A3 => n12697, A4 => 
                           n22357, Z => n9584);
   U11038 : NAND2_X1 port map( A1 => n1274, A2 => n33591, ZN => n13977);
   U11049 : INV_X1 port map( I => n17631, ZN => n13746);
   U11057 : NAND2_X1 port map( A1 => n1113, A2 => n10121, ZN => n11853);
   U11067 : INV_X1 port map( I => n17569, ZN => n11615);
   U11070 : AOI21_X1 port map( A1 => n6384, A2 => n22678, B => n32172, ZN => 
                           n9738);
   U11076 : NOR2_X1 port map( A1 => n30066, A2 => n22600, ZN => n7649);
   U11084 : NAND2_X1 port map( A1 => n22498, A2 => n5769, ZN => n22499);
   U11085 : INV_X1 port map( I => n22409, ZN => n1749);
   U11089 : NAND2_X1 port map( A1 => n14830, A2 => n22639, ZN => n15607);
   U11091 : NAND2_X1 port map( A1 => n8529, A2 => n30066, ZN => n7648);
   U11092 : NAND2_X1 port map( A1 => n14830, A2 => n16240, ZN => n11746);
   U11097 : OAI21_X1 port map( A1 => n14221, A2 => n14220, B => n22666, ZN => 
                           n4628);
   U11099 : NAND2_X1 port map( A1 => n1728, A2 => n1727, ZN => n1726);
   U11109 : NAND2_X1 port map( A1 => n9789, A2 => n1124, ZN => n22254);
   U11111 : NOR2_X1 port map( A1 => n22402, A2 => n16556, ZN => n16232);
   U11114 : OR2_X1 port map( A1 => n22544, A2 => n252, Z => n10137);
   U11116 : INV_X1 port map( I => n22369, ZN => n3522);
   U11118 : NAND2_X1 port map( A1 => n14713, A2 => n701, ZN => n3382);
   U11120 : NAND2_X1 port map( A1 => n11575, A2 => n9603, ZN => n3594);
   U11121 : INV_X1 port map( I => n22437, ZN => n16414);
   U11123 : NAND2_X1 port map( A1 => n4810, A2 => n905, ZN => n4809);
   U11137 : NAND2_X1 port map( A1 => n11011, A2 => n22673, ZN => n11010);
   U11139 : INV_X2 port map( I => n12488, ZN => n3567);
   U11140 : NOR2_X1 port map( A1 => n22510, A2 => n8527, ZN => n14765);
   U11146 : INV_X1 port map( I => n11378, ZN => n3325);
   U11149 : NOR2_X1 port map( A1 => n22536, A2 => n17626, ZN => n17146);
   U11156 : NAND2_X1 port map( A1 => n29158, A2 => n9737, ZN => n8287);
   U11158 : INV_X1 port map( I => n22522, ZN => n9654);
   U11164 : NOR2_X1 port map( A1 => n7964, A2 => n22558, ZN => n2844);
   U11174 : INV_X1 port map( I => n22455, ZN => n13665);
   U11175 : NAND2_X1 port map( A1 => n28865, A2 => n10622, ZN => n11147);
   U11178 : NAND2_X1 port map( A1 => n22639, A2 => n22640, ZN => n13881);
   U11180 : AND2_X1 port map( A1 => n1116, A2 => n28865, Z => n22112);
   U11183 : NOR2_X1 port map( A1 => n22537, A2 => n909, ZN => n3188);
   U11186 : NOR2_X1 port map( A1 => n22491, A2 => n26305, ZN => n12931);
   U11187 : INV_X1 port map( I => n22669, ZN => n15650);
   U11199 : NAND2_X1 port map( A1 => n17394, A2 => n907, ZN => n7897);
   U11208 : INV_X1 port map( I => n22504, ZN => n22025);
   U11210 : INV_X2 port map( I => n22414, ZN => n2066);
   U11213 : CLKBUF_X2 port map( I => n22677, Z => n16556);
   U11217 : INV_X1 port map( I => n22289, ZN => n16027);
   U11225 : INV_X1 port map( I => n10186, ZN => n21874);
   U11230 : NOR2_X1 port map( A1 => n14151, A2 => n14150, ZN => n15698);
   U11233 : NAND2_X1 port map( A1 => n15798, A2 => n22126, ZN => n15797);
   U11240 : INV_X1 port map( I => n15606, ZN => n4789);
   U11242 : INV_X1 port map( I => n13651, ZN => n4187);
   U11244 : INV_X1 port map( I => n17362, ZN => n4788);
   U11250 : NAND2_X1 port map( A1 => n15840, A2 => n6176, ZN => n10671);
   U11251 : OAI21_X1 port map( A1 => n21562, A2 => n21561, B => n22220, ZN => 
                           n13370);
   U11252 : OR2_X1 port map( A1 => n31930, A2 => n29180, Z => n9961);
   U11257 : INV_X1 port map( I => n22196, ZN => n9531);
   U11260 : NAND2_X1 port map( A1 => n21756, A2 => n33403, ZN => n15410);
   U11268 : INV_X1 port map( I => n21126, ZN => n9312);
   U11273 : NAND2_X1 port map( A1 => n21521, A2 => n21520, ZN => n11590);
   U11284 : NAND2_X1 port map( A1 => n21542, A2 => n30677, ZN => n15129);
   U11288 : NAND2_X1 port map( A1 => n5788, A2 => n5787, ZN => n7792);
   U11295 : INV_X1 port map( I => n21754, ZN => n21756);
   U11299 : OAI21_X1 port map( A1 => n12041, A2 => n21610, B => n27937, ZN => 
                           n3050);
   U11301 : INV_X1 port map( I => n26113, ZN => n2949);
   U11303 : OR2_X1 port map( A1 => n2441, A2 => n7592, Z => n2440);
   U11313 : INV_X1 port map( I => n21527, ZN => n8459);
   U11319 : NAND2_X1 port map( A1 => n21641, A2 => n21640, ZN => n4688);
   U11327 : NAND2_X1 port map( A1 => n21766, A2 => n28395, ZN => n5997);
   U11328 : NOR2_X1 port map( A1 => n21647, A2 => n26573, ZN => n11633);
   U11329 : INV_X1 port map( I => n21818, ZN => n21819);
   U11340 : AOI21_X1 port map( A1 => n10357, A2 => n21864, B => n15465, ZN => 
                           n21527);
   U11343 : AND2_X1 port map( A1 => n14738, A2 => n14739, Z => n9299);
   U11346 : INV_X1 port map( I => n21491, ZN => n11582);
   U11347 : NOR2_X1 port map( A1 => n33325, A2 => n15302, ZN => n9811);
   U11348 : NAND2_X1 port map( A1 => n777, A2 => n3497, ZN => n10346);
   U11349 : NOR2_X1 port map( A1 => n16441, A2 => n25975, ZN => n21479);
   U11352 : NOR2_X1 port map( A1 => n1138, A2 => n16735, ZN => n17164);
   U11356 : NAND2_X1 port map( A1 => n21496, A2 => n21601, ZN => n6237);
   U11358 : INV_X1 port map( I => n21797, ZN => n21800);
   U11371 : INV_X1 port map( I => n21842, ZN => n21750);
   U11373 : INV_X1 port map( I => n21643, ZN => n8733);
   U11375 : INV_X1 port map( I => n21740, ZN => n18055);
   U11377 : AND2_X1 port map( A1 => n29864, A2 => n21460, Z => n7388);
   U11378 : NOR2_X1 port map( A1 => n1139, A2 => n9205, ZN => n9204);
   U11381 : AND2_X1 port map( A1 => n29980, A2 => n15302, Z => n2202);
   U11382 : NAND2_X1 port map( A1 => n13213, A2 => n28099, ZN => n7947);
   U11386 : NOR2_X1 port map( A1 => n14397, A2 => n7182, ZN => n13869);
   U11387 : NAND2_X1 port map( A1 => n6181, A2 => n21387, ZN => n6179);
   U11388 : NOR2_X1 port map( A1 => n31197, A2 => n28099, ZN => n4098);
   U11392 : INV_X1 port map( I => n21510, ZN => n9059);
   U11397 : INV_X1 port map( I => n10357, ZN => n21587);
   U11398 : AND2_X1 port map( A1 => n2575, A2 => n2576, Z => n11362);
   U11399 : INV_X1 port map( I => n21723, ZN => n13187);
   U11401 : NAND2_X1 port map( A1 => n31042, A2 => n12827, ZN => n7365);
   U11407 : NOR2_X1 port map( A1 => n7182, A2 => n196, ZN => n15827);
   U11410 : INV_X1 port map( I => n13800, ZN => n11229);
   U11412 : INV_X1 port map( I => n21559, ZN => n12229);
   U11413 : INV_X1 port map( I => n12792, ZN => n1323);
   U11414 : NAND2_X1 port map( A1 => n8267, A2 => n6182, ZN => n6178);
   U11416 : INV_X1 port map( I => n12587, ZN => n6751);
   U11421 : INV_X1 port map( I => n11266, ZN => n21616);
   U11429 : NOR2_X1 port map( A1 => n21084, A2 => n10573, ZN => n10572);
   U11430 : OR2_X1 port map( A1 => n26635, A2 => n20940, Z => n12133);
   U11433 : INV_X1 port map( I => n13130, ZN => n21107);
   U11437 : NAND2_X1 port map( A1 => n7673, A2 => n17341, ZN => n11315);
   U11438 : NAND2_X1 port map( A1 => n21110, A2 => n21222, ZN => n8468);
   U11445 : NOR2_X1 port map( A1 => n21423, A2 => n32347, ZN => n6881);
   U11450 : INV_X1 port map( I => n6199, ZN => n6198);
   U11452 : NAND2_X1 port map( A1 => n21413, A2 => n8657, ZN => n3916);
   U11456 : OAI21_X1 port map( A1 => n28257, A2 => n921, B => n4088, ZN => 
                           n21051);
   U11460 : NAND2_X1 port map( A1 => n21115, A2 => n21114, ZN => n6743);
   U11463 : NAND2_X1 port map( A1 => n3105, A2 => n505, ZN => n3104);
   U11469 : AND2_X1 port map( A1 => n21209, A2 => n20874, Z => n9095);
   U11472 : NAND2_X1 port map( A1 => n11285, A2 => n21163, ZN => n12536);
   U11479 : NAND2_X1 port map( A1 => n21260, A2 => n921, ZN => n10655);
   U11481 : NAND2_X1 port map( A1 => n12492, A2 => n21270, ZN => n10339);
   U11482 : INV_X1 port map( I => n21074, ZN => n7147);
   U11485 : INV_X1 port map( I => n3937, ZN => n3936);
   U11492 : INV_X1 port map( I => n6303, ZN => n21361);
   U11494 : OAI21_X1 port map( A1 => n5684, A2 => n17341, B => n5683, ZN => 
                           n3937);
   U11495 : INV_X1 port map( I => n1783, ZN => n21127);
   U11501 : NAND2_X1 port map( A1 => n32242, A2 => n27382, ZN => n12340);
   U11502 : NAND2_X1 port map( A1 => n21357, A2 => n6307, ZN => n9462);
   U11509 : NOR2_X1 port map( A1 => n398, A2 => n7673, ZN => n1911);
   U11512 : INV_X1 port map( I => n21302, ZN => n21447);
   U11513 : NAND2_X1 port map( A1 => n21096, A2 => n15024, ZN => n15023);
   U11516 : OAI21_X1 port map( A1 => n4683, A2 => n320, B => n29255, ZN => 
                           n16545);
   U11517 : NAND2_X1 port map( A1 => n1146, A2 => n320, ZN => n21073);
   U11518 : NAND3_X1 port map( A1 => n11292, A2 => n9186, A3 => n1143, ZN => 
                           n11291);
   U11522 : NAND2_X1 port map( A1 => n13101, A2 => n21311, ZN => n11452);
   U11524 : NOR2_X1 port map( A1 => n12091, A2 => n15506, ZN => n2725);
   U11525 : OAI21_X1 port map( A1 => n21131, A2 => n21307, B => n31729, ZN => 
                           n6199);
   U11534 : NOR2_X1 port map( A1 => n8792, A2 => n8924, ZN => n7343);
   U11535 : NOR2_X1 port map( A1 => n599, A2 => n15015, ZN => n21415);
   U11536 : NOR2_X1 port map( A1 => n11513, A2 => n13367, ZN => n14489);
   U11539 : AND2_X1 port map( A1 => n21139, A2 => n21374, Z => n11979);
   U11541 : INV_X1 port map( I => n21081, ZN => n1868);
   U11544 : AND2_X1 port map( A1 => n21295, A2 => n9721, Z => n12111);
   U11552 : OAI21_X1 port map( A1 => n15874, A2 => n21398, B => n32625, ZN => 
                           n15112);
   U11561 : INV_X1 port map( I => n21053, ZN => n21054);
   U11564 : CLKBUF_X2 port map( I => n21053, Z => n16308);
   U11565 : INV_X2 port map( I => n7738, ZN => n21259);
   U11566 : INV_X1 port map( I => n20931, ZN => n21182);
   U11570 : AND2_X1 port map( A1 => n10533, A2 => n33566, Z => n3032);
   U11571 : INV_X1 port map( I => n21184, ZN => n21363);
   U11573 : INV_X1 port map( I => n27711, ZN => n16905);
   U11574 : INV_X1 port map( I => n21136, ZN => n21269);
   U11578 : INV_X2 port map( I => n9744, ZN => n17985);
   U11583 : INV_X1 port map( I => n10110, ZN => n9908);
   U11585 : INV_X1 port map( I => n8581, ZN => n11512);
   U11594 : NAND2_X1 port map( A1 => n7253, A2 => n7252, ZN => n6158);
   U11603 : INV_X1 port map( I => n18266, ZN => n4616);
   U11612 : INV_X1 port map( I => n20769, ZN => n17592);
   U11614 : NAND2_X1 port map( A1 => n20380, A2 => n20442, ZN => n4913);
   U11615 : NOR2_X1 port map( A1 => n20270, A2 => n28575, ZN => n20271);
   U11618 : INV_X1 port map( I => n20861, ZN => n7888);
   U11625 : NAND2_X1 port map( A1 => n3441, A2 => n3462, ZN => n3440);
   U11628 : NAND2_X1 port map( A1 => n33902, A2 => n12224, ZN => n6083);
   U11629 : NOR2_X1 port map( A1 => n12757, A2 => n12759, ZN => n5804);
   U11630 : INV_X1 port map( I => n20736, ZN => n20816);
   U11640 : INV_X1 port map( I => n15168, ZN => n3308);
   U11641 : INV_X1 port map( I => n20219, ZN => n17003);
   U11649 : NAND2_X1 port map( A1 => n20194, A2 => n32941, ZN => n11216);
   U11662 : NOR2_X1 port map( A1 => n5878, A2 => n20221, ZN => n7478);
   U11673 : NAND2_X1 port map( A1 => n9693, A2 => n1151, ZN => n4130);
   U11674 : NOR2_X1 port map( A1 => n20400, A2 => n819, ZN => n8354);
   U11675 : NAND2_X1 port map( A1 => n5498, A2 => n5497, ZN => n5496);
   U11676 : INV_X1 port map( I => n26424, ZN => n8868);
   U11680 : NAND2_X1 port map( A1 => n34013, A2 => n1863, ZN => n9419);
   U11681 : NAND2_X1 port map( A1 => n5275, A2 => n20345, ZN => n10716);
   U11684 : INV_X1 port map( I => n26041, ZN => n17791);
   U11689 : NAND2_X1 port map( A1 => n6925, A2 => n27771, ZN => n5835);
   U11692 : NAND2_X1 port map( A1 => n11038, A2 => n1153, ZN => n11037);
   U11693 : INV_X1 port map( I => n20197, ZN => n3069);
   U11694 : NAND2_X1 port map( A1 => n10351, A2 => n20515, ZN => n7254);
   U11697 : NAND2_X1 port map( A1 => n12583, A2 => n5415, ZN => n12582);
   U11704 : INV_X1 port map( I => n20405, ZN => n11445);
   U11712 : NAND2_X1 port map( A1 => n32940, A2 => n16190, ZN => n10623);
   U11713 : OAI21_X1 port map( A1 => n15553, A2 => n9774, B => n20563, ZN => 
                           n9773);
   U11715 : NAND3_X1 port map( A1 => n14719, A2 => n12966, A3 => n28376, ZN => 
                           n20501);
   U11724 : AND2_X1 port map( A1 => n20284, A2 => n20527, Z => n8582);
   U11730 : INV_X1 port map( I => n15225, ZN => n20319);
   U11731 : NAND2_X1 port map( A1 => n20227, A2 => n29938, ZN => n11666);
   U11733 : NAND2_X1 port map( A1 => n20304, A2 => n1028, ZN => n7698);
   U11740 : INV_X1 port map( I => n9719, ZN => n20199);
   U11741 : NOR2_X1 port map( A1 => n1811, A2 => n1032, ZN => n7033);
   U11743 : INV_X1 port map( I => n20304, ZN => n5217);
   U11744 : INV_X1 port map( I => n20306, ZN => n2134);
   U11748 : INV_X1 port map( I => n27600, ZN => n20300);
   U11749 : OR2_X1 port map( A1 => n5879, A2 => n5909, Z => n5908);
   U11752 : AND2_X1 port map( A1 => n16132, A2 => n933, Z => n20230);
   U11753 : NAND2_X1 port map( A1 => n819, A2 => n11988, ZN => n10431);
   U11754 : AND2_X1 port map( A1 => n20460, A2 => n20395, Z => n20366);
   U11755 : NAND2_X1 port map( A1 => n16606, A2 => n6531, ZN => n17393);
   U11768 : NAND2_X1 port map( A1 => n13538, A2 => n26881, ZN => n20181);
   U11769 : NAND2_X1 port map( A1 => n16146, A2 => n12421, ZN => n20502);
   U11770 : NAND2_X1 port map( A1 => n9688, A2 => n20310, ZN => n20179);
   U11778 : OAI21_X1 port map( A1 => n11502, A2 => n11501, B => n11500, ZN => 
                           n19816);
   U11783 : AND2_X1 port map( A1 => n20290, A2 => n20289, Z => n20291);
   U11788 : NAND2_X1 port map( A1 => n19534, A2 => n20037, ZN => n19535);
   U11796 : NAND2_X1 port map( A1 => n11501, A2 => n28644, ZN => n11500);
   U11800 : NAND2_X1 port map( A1 => n11350, A2 => n568, ZN => n19861);
   U11805 : NAND2_X1 port map( A1 => n14989, A2 => n4841, ZN => n5888);
   U11810 : INV_X1 port map( I => n6963, ZN => n7001);
   U11811 : NAND2_X1 port map( A1 => n14033, A2 => n31683, ZN => n14032);
   U11815 : INV_X1 port map( I => n13058, ZN => n19913);
   U11818 : NAND2_X1 port map( A1 => n3271, A2 => n3270, ZN => n3269);
   U11819 : NAND2_X1 port map( A1 => n8148, A2 => n20061, ZN => n19892);
   U11822 : NAND2_X1 port map( A1 => n19869, A2 => n8137, ZN => n19872);
   U11825 : OAI21_X1 port map( A1 => n16193, A2 => n20088, B => n1161, ZN => 
                           n6963);
   U11827 : INV_X1 port map( I => n14801, ZN => n3096);
   U11828 : NAND2_X1 port map( A1 => n1955, A2 => n10750, ZN => n1954);
   U11833 : OR2_X1 port map( A1 => n13425, A2 => n19991, Z => n13423);
   U11836 : NAND2_X1 port map( A1 => n10683, A2 => n16346, ZN => n8592);
   U11837 : NAND2_X1 port map( A1 => n7153, A2 => n20045, ZN => n6663);
   U11841 : NAND2_X1 port map( A1 => n20055, A2 => n9379, ZN => n11871);
   U11846 : AOI21_X1 port map( A1 => n579, A2 => n16491, B => n7460, ZN => 
                           n15906);
   U11847 : AND2_X1 port map( A1 => n1165, A2 => n5433, Z => n6951);
   U11853 : NAND2_X1 port map( A1 => n19818, A2 => n6961, ZN => n14107);
   U11855 : INV_X1 port map( I => n10484, ZN => n14173);
   U11856 : NAND2_X1 port map( A1 => n5718, A2 => n13583, ZN => n5717);
   U11870 : NAND2_X1 port map( A1 => n29187, A2 => n25980, ZN => n1799);
   U11875 : AND2_X1 port map( A1 => n28183, A2 => n33848, Z => n4308);
   U11878 : INV_X1 port map( I => n7525, ZN => n1974);
   U11880 : INV_X1 port map( I => n13346, ZN => n20077);
   U11881 : INV_X1 port map( I => n20118, ZN => n7153);
   U11884 : INV_X1 port map( I => n34153, ZN => n13425);
   U11889 : NOR2_X1 port map( A1 => n17711, A2 => n20068, ZN => n16516);
   U11891 : NOR2_X1 port map( A1 => n19965, A2 => n8371, ZN => n9105);
   U11899 : OAI21_X1 port map( A1 => n19891, A2 => n20096, B => n30692, ZN => 
                           n8148);
   U11904 : NAND2_X1 port map( A1 => n1040, A2 => n19456, ZN => n5828);
   U11909 : NOR2_X1 port map( A1 => n17060, A2 => n16694, ZN => n8216);
   U11910 : NAND2_X1 port map( A1 => n27097, A2 => n20152, ZN => n19979);
   U11911 : INV_X1 port map( I => n12085, ZN => n2290);
   U11915 : NAND2_X1 port map( A1 => n1043, A2 => n16579, ZN => n7737);
   U11916 : AND2_X1 port map( A1 => n13852, A2 => n19942, Z => n12061);
   U11917 : INV_X1 port map( I => n17060, ZN => n11142);
   U11921 : INV_X1 port map( I => n20106, ZN => n17696);
   U11923 : NAND3_X1 port map( A1 => n20106, A2 => n20107, A3 => n16243, ZN => 
                           n7579);
   U11924 : AND2_X1 port map( A1 => n19874, A2 => n149, Z => n11909);
   U11932 : INV_X2 port map( I => n5287, ZN => n13605);
   U11934 : NAND2_X1 port map( A1 => n577, A2 => n20096, ZN => n17441);
   U11940 : INV_X1 port map( I => n19469, ZN => n7191);
   U11942 : INV_X1 port map( I => n19433, ZN => n4894);
   U11945 : INV_X1 port map( I => n19462, ZN => n5190);
   U11948 : OAI21_X1 port map( A1 => n17293, A2 => n17291, B => n17290, ZN => 
                           n19633);
   U11949 : INV_X1 port map( I => n19682, ZN => n2469);
   U11950 : INV_X1 port map( I => n19545, ZN => n6680);
   U11953 : INV_X1 port map( I => n18125, ZN => n8266);
   U11954 : INV_X1 port map( I => n15188, ZN => n19757);
   U11962 : INV_X1 port map( I => n19461, ZN => n19696);
   U11963 : INV_X1 port map( I => n2282, ZN => n2281);
   U11965 : INV_X1 port map( I => n26683, ZN => n19570);
   U11967 : INV_X1 port map( I => n19352, ZN => n3073);
   U11969 : INV_X1 port map( I => n32697, ZN => n19448);
   U11972 : INV_X1 port map( I => n19445, ZN => n19587);
   U11975 : INV_X1 port map( I => n7109, ZN => n5608);
   U11988 : NAND2_X1 port map( A1 => n15930, A2 => n11262, ZN => n11261);
   U11993 : NOR2_X1 port map( A1 => n7575, A2 => n32802, ZN => n5332);
   U11995 : NAND2_X1 port map( A1 => n10828, A2 => n19164, ZN => n11278);
   U11997 : NAND2_X1 port map( A1 => n6282, A2 => n13252, ZN => n12894);
   U12000 : NAND2_X1 port map( A1 => n10856, A2 => n10855, ZN => n10854);
   U12004 : OAI21_X1 port map( A1 => n8233, A2 => n19128, B => n5635, ZN => 
                           n5637);
   U12007 : INV_X1 port map( I => n6440, ZN => n6029);
   U12010 : NAND2_X1 port map( A1 => n11263, A2 => n30817, ZN => n2518);
   U12019 : NAND2_X1 port map( A1 => n3115, A2 => n15910, ZN => n3114);
   U12021 : AND2_X1 port map( A1 => n18987, A2 => n19033, Z => n3116);
   U12024 : INV_X1 port map( I => n8092, ZN => n4879);
   U12027 : INV_X2 port map( I => n19370, ZN => n1372);
   U12029 : NAND2_X1 port map( A1 => n1766, A2 => n19219, ZN => n6795);
   U12034 : AOI21_X1 port map( A1 => n19093, A2 => n5813, B => n17386, ZN => 
                           n5946);
   U12035 : OAI22_X1 port map( A1 => n12034, A2 => n17725, B1 => n19107, B2 => 
                           n5907, ZN => n18457);
   U12036 : NAND2_X1 port map( A1 => n19209, A2 => n31948, ZN => n9318);
   U12038 : NOR2_X1 port map( A1 => n16444, A2 => n31451, ZN => n18455);
   U12042 : NAND2_X1 port map( A1 => n4363, A2 => n4202, ZN => n4360);
   U12043 : INV_X1 port map( I => n19243, ZN => n4217);
   U12050 : NAND2_X1 port map( A1 => n3022, A2 => n14597, ZN => n5221);
   U12057 : NAND2_X1 port map( A1 => n19128, A2 => n7967, ZN => n7966);
   U12059 : NOR2_X1 port map( A1 => n14806, A2 => n10828, ZN => n17527);
   U12060 : NAND2_X1 port map( A1 => n19215, A2 => n1836, ZN => n6603);
   U12064 : OAI21_X1 port map( A1 => n13389, A2 => n11807, B => n13390, ZN => 
                           n13391);
   U12075 : INV_X1 port map( I => n9508, ZN => n8671);
   U12086 : INV_X1 port map( I => n9887, ZN => n3024);
   U12087 : INV_X1 port map( I => n3516, ZN => n3499);
   U12089 : NOR2_X1 port map( A1 => n19293, A2 => n7275, ZN => n19297);
   U12090 : NAND2_X1 port map( A1 => n15928, A2 => n15927, ZN => n10910);
   U12093 : NOR2_X1 port map( A1 => n7517, A2 => n13526, ZN => n7516);
   U12097 : NAND2_X1 port map( A1 => n14327, A2 => n14328, ZN => n8489);
   U12111 : OAI21_X1 port map( A1 => n18659, A2 => n12199, B => n12198, ZN => 
                           n10693);
   U12117 : NOR2_X1 port map( A1 => n7454, A2 => n7518, ZN => n7517);
   U12120 : INV_X1 port map( I => n18896, ZN => n7714);
   U12121 : NOR2_X1 port map( A1 => n12799, A2 => n18339, ZN => n18996);
   U12122 : NAND2_X1 port map( A1 => n18686, A2 => n15575, ZN => n15574);
   U12123 : NAND2_X1 port map( A1 => n5587, A2 => n1060, ZN => n5561);
   U12125 : NAND2_X1 port map( A1 => n5586, A2 => n18680, ZN => n4717);
   U12128 : NAND2_X1 port map( A1 => n18803, A2 => n18785, ZN => n6399);
   U12135 : AOI21_X1 port map( A1 => n10367, A2 => n10366, B => n18678, ZN => 
                           n10365);
   U12136 : NAND2_X1 port map( A1 => n18336, A2 => n18755, ZN => n9835);
   U12138 : NOR2_X1 port map( A1 => n18499, A2 => n18605, ZN => n16328);
   U12140 : NAND2_X1 port map( A1 => n4868, A2 => n1190, ZN => n8570);
   U12143 : OAI21_X1 port map( A1 => n17926, A2 => n18894, B => n18795, ZN => 
                           n12814);
   U12150 : NOR2_X1 port map( A1 => n18870, A2 => n18871, ZN => n10305);
   U12153 : NOR2_X1 port map( A1 => n3218, A2 => n18891, ZN => n14544);
   U12158 : NAND3_X1 port map( A1 => n15348, A2 => n18579, A3 => n18856, ZN => 
                           n5124);
   U12159 : NAND2_X1 port map( A1 => n11410, A2 => n6891, ZN => n6889);
   U12162 : INV_X1 port map( I => n18410, ZN => n18522);
   U12163 : NAND2_X1 port map( A1 => n6612, A2 => n16614, ZN => n18309);
   U12166 : AND2_X1 port map( A1 => n18702, A2 => n16352, Z => n12132);
   U12169 : NOR2_X1 port map( A1 => n18130, A2 => n13738, ZN => n18333);
   U12172 : NAND2_X1 port map( A1 => n33205, A2 => n16287, ZN => n6429);
   U12174 : INV_X1 port map( I => n18659, ZN => n11517);
   U12175 : NAND2_X1 port map( A1 => n18881, A2 => n28578, ZN => n10639);
   U12177 : AND2_X1 port map( A1 => n16474, A2 => n18349, Z => n16120);
   U12180 : INV_X1 port map( I => n18576, ZN => n10565);
   U12182 : INV_X1 port map( I => n15265, ZN => n18792);
   U12186 : CLKBUF_X2 port map( I => n18654, Z => n18446);
   U12189 : CLKBUF_X2 port map( I => n18756, Z => n14093);
   U12191 : INV_X1 port map( I => n25693, ZN => n25694);
   U12192 : INV_X1 port map( I => n25126, ZN => n11034);
   U12193 : AND2_X1 port map( A1 => n12006, A2 => n22, Z => n12130);
   U12194 : INV_X1 port map( I => n25319, ZN => n24507);
   U12196 : INV_X1 port map( I => n16479, ZN => n3259);
   U12197 : INV_X1 port map( I => n16654, ZN => n10308);
   U12198 : INV_X1 port map( I => n25815, ZN => n10584);
   U12199 : INV_X1 port map( I => n25751, ZN => n13033);
   U12203 : INV_X1 port map( I => n16502, ZN => n15409);
   U12204 : INV_X1 port map( I => n24426, ZN => n12754);
   U12206 : INV_X1 port map( I => n16423, ZN => n9874);
   U12208 : INV_X1 port map( I => n25598, ZN => n1546);
   U12212 : INV_X1 port map( I => n24943, ZN => n24944);
   U12218 : INV_X1 port map( I => n25131, ZN => n1653);
   U12219 : INV_X1 port map( I => n25288, ZN => n14526);
   U12220 : INV_X1 port map( I => n25191, ZN => n25192);
   U12222 : INV_X1 port map( I => n24738, ZN => n5101);
   U12223 : INV_X1 port map( I => n16679, ZN => n14300);
   U12224 : INV_X1 port map( I => n25465, ZN => n25466);
   U12225 : INV_X1 port map( I => n25074, ZN => n15742);
   U12226 : INV_X1 port map( I => n25506, ZN => n25507);
   U12227 : INV_X1 port map( I => n24917, ZN => n24918);
   U12230 : INV_X1 port map( I => n16454, ZN => n15779);
   U12232 : INV_X1 port map( I => n24748, ZN => n9527);
   U12233 : INV_X1 port map( I => n24907, ZN => n13438);
   U12237 : INV_X1 port map( I => n25457, ZN => n3027);
   U12238 : CLKBUF_X2 port map( I => n18335, Z => n18755);
   U12240 : INV_X1 port map( I => n25560, ZN => n8500);
   U12241 : INV_X1 port map( I => n16613, ZN => n14885);
   U12243 : INV_X1 port map( I => n16671, ZN => n17063);
   U12244 : INV_X1 port map( I => n16482, ZN => n8139);
   U12245 : INV_X1 port map( I => n16602, ZN => n10553);
   U12246 : INV_X1 port map( I => n16696, ZN => n12719);
   U12248 : INV_X1 port map( I => n25001, ZN => n12695);
   U12249 : INV_X1 port map( I => n16680, ZN => n15147);
   U12250 : INV_X1 port map( I => n16642, ZN => n1390);
   U12254 : CLKBUF_X2 port map( I => Key(89), Z => n24962);
   U12255 : INV_X1 port map( I => n16322, ZN => n1397);
   U12257 : INV_X1 port map( I => n25722, ZN => n1402);
   U12259 : INV_X1 port map( I => n16690, ZN => n1403);
   U12260 : INV_X1 port map( I => n16631, ZN => n1405);
   U12262 : INV_X1 port map( I => n25554, ZN => n1409);
   U12263 : INV_X1 port map( I => n16390, ZN => n1411);
   U12266 : CLKBUF_X2 port map( I => Key(137), Z => n25182);
   U12268 : INV_X1 port map( I => n25218, ZN => n1414);
   U12270 : INV_X1 port map( I => n25049, ZN => n1416);
   U12271 : INV_X1 port map( I => n25908, ZN => n1417);
   U12273 : INV_X1 port map( I => n16578, ZN => n1420);
   U12274 : INV_X1 port map( I => n25716, ZN => n1421);
   U12276 : INV_X1 port map( I => n25038, ZN => n1423);
   U12277 : CLKBUF_X2 port map( I => Key(21), Z => n16698);
   U12278 : CLKBUF_X2 port map( I => Key(63), Z => n25282);
   U12280 : INV_X1 port map( I => n16584, ZN => n1425);
   U12282 : INV_X1 port map( I => n16506, ZN => n1426);
   U12283 : INV_X1 port map( I => n16301, ZN => n1429);
   U12284 : CLKBUF_X2 port map( I => Key(164), Z => n25074);
   U12285 : INV_X1 port map( I => n16666, ZN => n1432);
   U12286 : INV_X1 port map( I => n25009, ZN => n1433);
   U12287 : INV_X1 port map( I => n16622, ZN => n1434);
   U12289 : XOR2_X1 port map( A1 => n31491, A2 => n10776, Z => n1436);
   U12293 : NAND3_X1 port map( A1 => n1438, A2 => n3790, A3 => n1163, ZN => 
                           n19934);
   U12294 : XOR2_X1 port map( A1 => Plaintext(129), A2 => Key(129), Z => n17189
                           );
   U12304 : XOR2_X1 port map( A1 => n22235, A2 => n13740, Z => n1445);
   U12305 : NOR2_X1 port map( A1 => n32787, A2 => n12317, ZN => n18802);
   U12306 : INV_X2 port map( I => n6776, ZN => n12317);
   U12320 : INV_X1 port map( I => n1464, ZN => n19485);
   U12321 : XOR2_X1 port map( A1 => n1464, A2 => n16654, Z => n2980);
   U12323 : XOR2_X1 port map( A1 => n1464, A2 => n3568, Z => n19648);
   U12324 : XOR2_X1 port map( A1 => n1464, A2 => n2469, Z => n1541);
   U12326 : NOR2_X1 port map( A1 => n1465, A2 => n31907, ZN => n3746);
   U12332 : XOR2_X1 port map( A1 => n24758, A2 => n24757, Z => n1468);
   U12337 : XOR2_X1 port map( A1 => n23277, A2 => n1470, Z => n2164);
   U12338 : XOR2_X1 port map( A1 => n23299, A2 => n25500, Z => n1470);
   U12339 : OAI21_X2 port map( A1 => n23080, A2 => n18129, B => n3786, ZN => 
                           n23299);
   U12343 : NAND2_X2 port map( A1 => n1474, A2 => n1473, ZN => n16798);
   U12346 : XOR2_X1 port map( A1 => n17385, A2 => n3550, Z => n2436);
   U12348 : XOR2_X1 port map( A1 => n17385, A2 => n25554, Z => n17564);
   U12349 : XOR2_X1 port map( A1 => n22120, A2 => n17385, Z => n4397);
   U12350 : XOR2_X1 port map( A1 => n1481, A2 => n1483, Z => n10287);
   U12352 : XOR2_X1 port map( A1 => n27174, A2 => n24968, Z => n1482);
   U12355 : XOR2_X1 port map( A1 => n21014, A2 => n21015, Z => n1483);
   U12356 : XOR2_X1 port map( A1 => n20818, A2 => n20801, Z => n21015);
   U12359 : XOR2_X1 port map( A1 => n20819, A2 => n20717, Z => n21014);
   U12362 : NOR2_X2 port map( A1 => n10905, A2 => n10904, ZN => n1485);
   U12368 : NOR2_X1 port map( A1 => n23763, A2 => n1489, ZN => n17537);
   U12379 : NAND2_X2 port map( A1 => n1497, A2 => n1496, ZN => n5268);
   U12383 : AOI22_X2 port map( A1 => n1506, A2 => n23869, B1 => n13224, B2 => 
                           n23867, ZN => n13223);
   U12398 : OAI21_X2 port map( A1 => n1524, A2 => n1523, B => n17357, ZN => 
                           n22909);
   U12405 : XOR2_X1 port map( A1 => n23166, A2 => n1537, Z => n1536);
   U12406 : XOR2_X1 port map( A1 => n23183, A2 => n23218, Z => n23166);
   U12407 : XOR2_X1 port map( A1 => n51, A2 => n1391, Z => n1537);
   U12412 : NAND3_X2 port map( A1 => n9950, A2 => n23054, A3 => n9949, ZN => 
                           n23267);
   U12417 : NAND2_X2 port map( A1 => n2281, A2 => n2279, ZN => n3568);
   U12418 : XOR2_X1 port map( A1 => n2470, A2 => n1541, Z => n1540);
   U12424 : XOR2_X1 port map( A1 => n32861, A2 => n27252, Z => n4467);
   U12427 : XOR2_X1 port map( A1 => n20670, A2 => n1546, Z => n1545);
   U12436 : XOR2_X1 port map( A1 => n24356, A2 => n1560, Z => n18091);
   U12438 : XOR2_X1 port map( A1 => n1560, A2 => n16655, Z => n24391);
   U12439 : XOR2_X1 port map( A1 => n14789, A2 => n1560, Z => n7259);
   U12440 : XOR2_X1 port map( A1 => n1560, A2 => n1230, Z => n10089);
   U12448 : NAND2_X2 port map( A1 => n1565, A2 => n1564, ZN => n23293);
   U12455 : NOR2_X2 port map( A1 => n32878, A2 => n4885, ZN => n1573);
   U12467 : XOR2_X1 port map( A1 => n3550, A2 => n21952, Z => n1590);
   U12468 : XOR2_X1 port map( A1 => n5482, A2 => n14289, Z => n1587);
   U12470 : XOR2_X1 port map( A1 => n22217, A2 => n454, Z => n1588);
   U12471 : XOR2_X1 port map( A1 => n11736, A2 => n22098, Z => n22217);
   U12481 : NOR2_X1 port map( A1 => n15110, A2 => n823, ZN => n1596);
   U12482 : XOR2_X1 port map( A1 => n31843, A2 => n16551, Z => n17858);
   U12497 : XOR2_X1 port map( A1 => n20443, A2 => n20669, Z => n1612);
   U12498 : XOR2_X1 port map( A1 => n8568, A2 => n20917, Z => n20669);
   U12504 : XOR2_X1 port map( A1 => n12121, A2 => n19519, Z => n1616);
   U12513 : XOR2_X1 port map( A1 => n4554, A2 => n23440, Z => n1621);
   U12517 : XOR2_X1 port map( A1 => n23334, A2 => n452, Z => n1622);
   U12522 : XOR2_X1 port map( A1 => n27114, A2 => n13545, Z => n24538);
   U12523 : XOR2_X1 port map( A1 => n27114, A2 => n7574, Z => n18174);
   U12528 : OAI21_X1 port map( A1 => n4150, A2 => n5872, B => n25693, ZN => 
                           n1627);
   U12529 : OR2_X1 port map( A1 => n5872, A2 => n25693, Z => n1628);
   U12530 : XOR2_X1 port map( A1 => n19746, A2 => n9880, Z => n19766);
   U12532 : AOI21_X2 port map( A1 => n1631, A2 => n19254, B => n1629, ZN => 
                           n19746);
   U12535 : OAI21_X1 port map( A1 => n20523, A2 => n1150, B => n1635, ZN => 
                           n20231);
   U12537 : NAND2_X2 port map( A1 => n17786, A2 => n17784, ZN => n1636);
   U12543 : XOR2_X1 port map( A1 => n17384, A2 => n2155, Z => n1644);
   U12544 : NAND2_X2 port map( A1 => n1646, A2 => n1645, ZN => n17384);
   U12545 : XOR2_X1 port map( A1 => n22012, A2 => n25908, Z => n21889);
   U12549 : INV_X2 port map( I => n11238, ZN => n22487);
   U12552 : NAND2_X2 port map( A1 => n12823, A2 => n22874, ZN => n23331);
   U12554 : XOR2_X1 port map( A1 => n10201, A2 => n23507, Z => n1676);
   U12555 : NAND2_X2 port map( A1 => n2112, A2 => n2111, ZN => n23507);
   U12559 : AOI22_X2 port map( A1 => n4255, A2 => n18784, B1 => n18787, B2 => 
                           n18786, ZN => n4392);
   U12560 : NAND2_X1 port map( A1 => n4392, A2 => n2150, ZN => n5876);
   U12561 : XOR2_X1 port map( A1 => n1686, A2 => n1682, Z => n17271);
   U12562 : XOR2_X1 port map( A1 => n1685, A2 => n1683, Z => n1682);
   U12563 : XOR2_X1 port map( A1 => n20970, A2 => n25001, Z => n1683);
   U12565 : XOR2_X1 port map( A1 => n20891, A2 => n20892, Z => n1685);
   U12567 : NAND2_X2 port map( A1 => n20385, A2 => n20386, ZN => n20891);
   U12569 : XOR2_X1 port map( A1 => n3705, A2 => n20839, Z => n20890);
   U12571 : NAND2_X2 port map( A1 => n20351, A2 => n20350, ZN => n20982);
   U12572 : INV_X2 port map( I => n20727, ZN => n20822);
   U12578 : XOR2_X1 port map( A1 => n14789, A2 => n24403, Z => n24556);
   U12584 : XOR2_X1 port map( A1 => n9577, A2 => n2122, Z => n1695);
   U12592 : XOR2_X1 port map( A1 => n24567, A2 => n10163, Z => n5530);
   U12598 : XOR2_X1 port map( A1 => n20782, A2 => n3119, Z => n1704);
   U12599 : INV_X2 port map( I => n15865, ZN => n17661);
   U12605 : XOR2_X1 port map( A1 => Plaintext(179), A2 => Key(179), Z => n18874
                           );
   U12606 : INV_X2 port map( I => n10181, ZN => n18101);
   U12607 : XOR2_X1 port map( A1 => Plaintext(178), A2 => Key(178), Z => n9909)
                           ;
   U12609 : XOR2_X1 port map( A1 => n13477, A2 => n29312, Z => n3178);
   U12610 : NAND2_X2 port map( A1 => n2037, A2 => n12368, ZN => n2041);
   U12613 : XOR2_X1 port map( A1 => n28239, A2 => n24804, Z => n1712);
   U12618 : NAND2_X2 port map( A1 => n7325, A2 => n11590, ZN => n10979);
   U12623 : INV_X1 port map( I => n23858, ZN => n1732);
   U12628 : XOR2_X1 port map( A1 => n11349, A2 => n25969, Z => n1741);
   U12634 : XOR2_X1 port map( A1 => n12124, A2 => n541, Z => n1742);
   U12639 : INV_X2 port map( I => n6288, ZN => n25687);
   U12645 : NOR2_X1 port map( A1 => n25675, A2 => n14732, ZN => n1756);
   U12648 : XOR2_X1 port map( A1 => n9189, A2 => n1760, Z => n1761);
   U12649 : XOR2_X1 port map( A1 => n16693, A2 => n1069, Z => n1760);
   U12658 : INV_X2 port map( I => n11628, ZN => n6474);
   U12679 : XOR2_X1 port map( A1 => n1780, A2 => n1779, Z => n1778);
   U12680 : XOR2_X1 port map( A1 => n14789, A2 => n13419, Z => n1779);
   U12681 : XOR2_X1 port map( A1 => n24761, A2 => n8306, Z => n1780);
   U12682 : XOR2_X1 port map( A1 => n24472, A2 => n14967, Z => n1781);
   U12683 : NAND2_X2 port map( A1 => n7660, A2 => n7658, ZN => n4124);
   U12685 : XOR2_X1 port map( A1 => n1791, A2 => n1794, Z => n15365);
   U12686 : XOR2_X1 port map( A1 => n1793, A2 => n1792, Z => n1791);
   U12687 : XOR2_X1 port map( A1 => n23336, A2 => n24374, Z => n1792);
   U12689 : XOR2_X1 port map( A1 => n1796, A2 => n1795, Z => n1794);
   U12693 : OAI21_X1 port map( A1 => n25980, A2 => n1362, B => n1799, ZN => 
                           n3925);
   U12694 : NAND2_X2 port map( A1 => n1818, A2 => n23594, ZN => n9964);
   U12696 : NAND4_X1 port map( A1 => n14548, A2 => n1818, A3 => n14550, A4 => 
                           n23594, ZN => n1800);
   U12697 : NAND2_X1 port map( A1 => n3779, A2 => n32005, ZN => n3856);
   U12700 : XOR2_X1 port map( A1 => n20886, A2 => n5024, Z => n1801);
   U12704 : NAND2_X1 port map( A1 => n1803, A2 => n16041, ZN => n17089);
   U12706 : OAI21_X1 port map( A1 => n9732, A2 => n31178, B => n32867, ZN => 
                           n9731);
   U12714 : XOR2_X1 port map( A1 => n1825, A2 => n23425, Z => n23426);
   U12716 : XOR2_X1 port map( A1 => n17775, A2 => n1825, Z => n23062);
   U12717 : XOR2_X1 port map( A1 => n23529, A2 => n1825, Z => n23182);
   U12721 : XOR2_X1 port map( A1 => n20593, A2 => n20997, Z => n2009);
   U12723 : NOR3_X2 port map( A1 => n7478, A2 => n19957, A3 => n7479, ZN => 
                           n20699);
   U12725 : OAI21_X1 port map( A1 => n7555, A2 => n28736, B => n15323, ZN => 
                           n1832);
   U12726 : NAND2_X1 port map( A1 => n1834, A2 => n25124, ZN => n1833);
   U12727 : NAND2_X1 port map( A1 => n7554, A2 => n15323, ZN => n1834);
   U12729 : NOR2_X1 port map( A1 => n881, A2 => n32337, ZN => n15429);
   U12738 : OAI21_X1 port map( A1 => n5628, A2 => n30033, B => n17644, ZN => 
                           n20877);
   U12741 : XOR2_X1 port map( A1 => n3929, A2 => n24748, Z => n1844);
   U12742 : XOR2_X1 port map( A1 => n20776, A2 => n7294, Z => n1845);
   U12762 : NAND2_X2 port map( A1 => n1862, A2 => n3385, ZN => n25221);
   U12767 : XOR2_X1 port map( A1 => n32822, A2 => n2388, Z => n3357);
   U12775 : NAND2_X2 port map( A1 => n9195, A2 => n25701, ZN => n1874);
   U12780 : XOR2_X1 port map( A1 => n1881, A2 => n3176, Z => n3816);
   U12781 : XOR2_X1 port map( A1 => n12413, A2 => n19441, Z => n1881);
   U12788 : INV_X1 port map( I => n33621, ZN => n18803);
   U12790 : XOR2_X1 port map( A1 => n28730, A2 => n24923, Z => n1884);
   U12794 : XOR2_X1 port map( A1 => n20838, A2 => n20748, Z => n1886);
   U12795 : XOR2_X1 port map( A1 => n20747, A2 => n21043, Z => n20838);
   U12798 : NAND2_X1 port map( A1 => n19837, A2 => n20037, ZN => n19838);
   U12808 : OR2_X1 port map( A1 => n19976, A2 => n32746, Z => n1900);
   U12811 : XOR2_X1 port map( A1 => n859, A2 => n1903, Z => n1902);
   U12814 : XOR2_X1 port map( A1 => n10824, A2 => n1970, Z => n1905);
   U12817 : INV_X1 port map( I => n11617, ZN => n1909);
   U12824 : AOI21_X1 port map( A1 => n28737, A2 => n17341, B => n16184, ZN => 
                           n1914);
   U12827 : XOR2_X1 port map( A1 => n31616, A2 => n24962, Z => n5012);
   U12828 : XOR2_X1 port map( A1 => n31616, A2 => n25182, Z => n21947);
   U12829 : XOR2_X1 port map( A1 => n22055, A2 => n31616, Z => n16912);
   U12835 : AOI21_X1 port map( A1 => n25234, A2 => n16589, B => n8219, ZN => 
                           n8121);
   U12837 : XOR2_X1 port map( A1 => n1928, A2 => n1927, Z => n10436);
   U12838 : XOR2_X1 port map( A1 => n20679, A2 => n25476, Z => n1927);
   U12839 : XOR2_X1 port map( A1 => n3929, A2 => n21016, Z => n1928);
   U12842 : XOR2_X1 port map( A1 => n14897, A2 => n11170, Z => n11169);
   U12844 : XOR2_X1 port map( A1 => n2362, A2 => n12141, Z => n12260);
   U12849 : XOR2_X1 port map( A1 => n4295, A2 => n32981, Z => n1936);
   U12864 : XOR2_X1 port map( A1 => n27167, A2 => n1191, Z => n1948);
   U12865 : XOR2_X1 port map( A1 => n13470, A2 => n14665, Z => n24774);
   U12868 : NAND2_X1 port map( A1 => n30330, A2 => n1951, ZN => n25069);
   U12869 : NOR2_X1 port map( A1 => n25076, A2 => n1951, ZN => n12304);
   U12870 : NAND3_X1 port map( A1 => n25076, A2 => n25066, A3 => n1951, ZN => 
                           n25068);
   U12874 : OAI21_X1 port map( A1 => n12329, A2 => n25066, B => n1951, ZN => 
                           n1950);
   U12879 : MUX2_X1 port map( I0 => n10086, I1 => n19921, S => n10752, Z => 
                           n1955);
   U12889 : INV_X1 port map( I => n1982, ZN => n13149);
   U12891 : XOR2_X1 port map( A1 => n19672, A2 => n1984, Z => n11627);
   U12892 : XOR2_X1 port map( A1 => n1984, A2 => n16598, Z => n17538);
   U12894 : NAND2_X1 port map( A1 => n24076, A2 => n1233, ZN => n24077);
   U12899 : XOR2_X1 port map( A1 => n4134, A2 => n6966, Z => n1988);
   U12903 : XOR2_X1 port map( A1 => n34078, A2 => n22198, Z => n1990);
   U12905 : XOR2_X1 port map( A1 => n14851, A2 => n22240, Z => n1992);
   U12908 : INV_X2 port map( I => n6462, ZN => n13612);
   U12913 : XOR2_X1 port map( A1 => n20852, A2 => n1993, Z => n14668);
   U12918 : NAND2_X1 port map( A1 => n219, A2 => n1040, ZN => n19995);
   U12929 : XOR2_X1 port map( A1 => n24812, A2 => n24554, Z => n2012);
   U12934 : XOR2_X1 port map( A1 => n24664, A2 => n25071, Z => n2015);
   U12937 : AOI22_X2 port map( A1 => n2018, A2 => n11497, B1 => n27947, B2 => 
                           n24460, ZN => n25686);
   U12947 : XOR2_X1 port map( A1 => n24486, A2 => n2048, Z => n2043);
   U12948 : XOR2_X1 port map( A1 => n24770, A2 => n2864, Z => n24486);
   U12949 : XOR2_X1 port map( A1 => n16917, A2 => n13810, Z => n2044);
   U12951 : XOR2_X1 port map( A1 => n1228, A2 => n14762, Z => n13810);
   U12955 : NAND2_X1 port map( A1 => n26447, A2 => n2049, ZN => n25673);
   U12959 : XOR2_X1 port map( A1 => n16608, A2 => n19767, Z => n2053);
   U12960 : XOR2_X1 port map( A1 => n3357, A2 => n3358, Z => n2054);
   U12968 : XOR2_X1 port map( A1 => n23233, A2 => n23536, Z => n15497);
   U12969 : XOR2_X1 port map( A1 => n1258, A2 => n721, Z => n14122);
   U12976 : NOR2_X1 port map( A1 => n22487, A2 => n2066, ZN => n13169);
   U12977 : NAND2_X1 port map( A1 => n31964, A2 => n2066, ZN => n16963);
   U12978 : MUX2_X1 port map( I0 => n2066, I1 => n31964, S => n33046, Z => 
                           n11246);
   U12981 : AOI22_X2 port map( A1 => n13364, A2 => n17398, B1 => n8145, B2 => 
                           n13936, ZN => n24240);
   U12990 : NAND2_X1 port map( A1 => n1098, A2 => n34009, ZN => n8852);
   U12991 : NAND3_X1 port map( A1 => n763, A2 => n7197, A3 => n2081, ZN => 
                           n18905);
   U12992 : OAI21_X1 port map( A1 => n825, A2 => n31970, B => n2081, ZN => 
                           n16908);
   U12996 : XOR2_X1 port map( A1 => n2082, A2 => n22155, Z => n8341);
   U12999 : NOR2_X1 port map( A1 => n23046, A2 => n808, ZN => n2084);
   U13000 : NOR2_X1 port map( A1 => n13121, A2 => n13120, ZN => n2085);
   U13018 : XOR2_X1 port map( A1 => n2095, A2 => n2097, Z => n8099);
   U13021 : XOR2_X1 port map( A1 => n22309, A2 => n22310, Z => n2097);
   U13022 : XOR2_X1 port map( A1 => n11736, A2 => n13564, Z => n22310);
   U13023 : AOI21_X2 port map( A1 => n4688, A2 => n21643, B => n4687, ZN => 
                           n13564);
   U13029 : NAND2_X2 port map( A1 => n11396, A2 => n14844, ZN => n15502);
   U13040 : INV_X2 port map( I => n2108, ZN => n5897);
   U13042 : XOR2_X1 port map( A1 => n3599, A2 => n19632, Z => n19636);
   U13043 : XOR2_X1 port map( A1 => n3599, A2 => n19072, Z => n10224);
   U13051 : NAND2_X1 port map( A1 => n11153, A2 => n2118, ZN => n11152);
   U13054 : XOR2_X1 port map( A1 => n2331, A2 => n25669, Z => n2122);
   U13068 : XOR2_X1 port map( A1 => n30749, A2 => n20729, Z => n15936);
   U13073 : XOR2_X1 port map( A1 => n22150, A2 => n5352, Z => n2144);
   U13079 : NOR2_X1 port map( A1 => n10203, A2 => n26417, ZN => n19092);
   U13080 : NAND3_X1 port map( A1 => n10203, A2 => n31658, A3 => n26417, ZN => 
                           n18987);
   U13081 : AOI21_X1 port map( A1 => n31658, A2 => n8141, B => n26417, ZN => 
                           n18790);
   U13082 : OAI21_X1 port map( A1 => n5813, A2 => n8141, B => n26417, ZN => 
                           n5812);
   U13087 : NAND2_X1 port map( A1 => n9521, A2 => n4019, ZN => n2154);
   U13089 : XOR2_X1 port map( A1 => n33700, A2 => n15000, Z => n2155);
   U13092 : XOR2_X1 port map( A1 => n13020, A2 => n5031, Z => n2161);
   U13093 : INV_X2 port map( I => n2163, ZN => n13297);
   U13095 : AND2_X1 port map( A1 => n31916, A2 => n13297, Z => n23562);
   U13099 : XOR2_X1 port map( A1 => n582, A2 => n16678, Z => n9201);
   U13101 : XOR2_X1 port map( A1 => Plaintext(191), A2 => Key(191), Z => n10891
                           );
   U13108 : AOI21_X1 port map( A1 => n24924, A2 => n2180, B => n15799, ZN => 
                           n24931);
   U13115 : XOR2_X1 port map( A1 => n23454, A2 => n27243, Z => n2190);
   U13116 : NOR2_X1 port map( A1 => n5568, A2 => n2191, ZN => n16348);
   U13117 : NAND3_X1 port map( A1 => n3646, A2 => n7929, A3 => n2191, ZN => 
                           n16583);
   U13118 : OAI21_X1 port map( A1 => n25247, A2 => n34109, B => n2191, ZN => 
                           n8036);
   U13119 : NAND2_X2 port map( A1 => n4552, A2 => n25245, ZN => n2191);
   U13123 : NAND3_X2 port map( A1 => n2197, A2 => n13563, A3 => n13562, ZN => 
                           n16331);
   U13128 : NAND2_X1 port map( A1 => n20379, A2 => n2205, ZN => n2204);
   U13129 : NOR2_X1 port map( A1 => n6679, A2 => n20635, ZN => n2205);
   U13132 : NAND2_X1 port map( A1 => n2209, A2 => n25687, ZN => n25680);
   U13134 : OAI22_X1 port map( A1 => n26447, A2 => n27173, B1 => n25687, B2 => 
                           n2209, ZN => n2208);
   U13136 : XOR2_X1 port map( A1 => n24370, A2 => n16733, Z => n9681);
   U13140 : XOR2_X1 port map( A1 => n2212, A2 => n24541, Z => n2211);
   U13141 : XOR2_X1 port map( A1 => n705, A2 => n26002, Z => n2212);
   U13143 : OAI21_X2 port map( A1 => n12919, A2 => n2219, B => n2215, ZN => 
                           n21910);
   U13149 : NAND2_X1 port map( A1 => n3007, A2 => n1274, ZN => n2226);
   U13151 : XOR2_X1 port map( A1 => n11641, A2 => n620, Z => n2547);
   U13154 : NOR2_X1 port map( A1 => n31046, A2 => n2229, ZN => n19817);
   U13158 : NAND3_X1 port map( A1 => n28734, A2 => n25322, A3 => n16041, ZN => 
                           n25323);
   U13161 : NAND2_X1 port map( A1 => n25320, A2 => n28734, ZN => n9733);
   U13162 : NOR2_X1 port map( A1 => n8770, A2 => n2237, ZN => n12917);
   U13164 : NAND3_X1 port map( A1 => n1028, A2 => n1151, A3 => n2237, ZN => 
                           n7252);
   U13181 : XOR2_X1 port map( A1 => n22036, A2 => n16523, Z => n2261);
   U13182 : XOR2_X1 port map( A1 => n2262, A2 => n12695, Z => Ciphertext(32));
   U13186 : OAI21_X1 port map( A1 => n3019, A2 => n30279, B => n2266, ZN => 
                           n2265);
   U13189 : XOR2_X1 port map( A1 => n21023, A2 => n2268, Z => n2267);
   U13190 : XOR2_X1 port map( A1 => n7717, A2 => n25545, Z => n2268);
   U13195 : XOR2_X1 port map( A1 => n19701, A2 => n19697, Z => n18166);
   U13196 : XNOR2_X1 port map( A1 => n16349, A2 => n19661, ZN => n19701);
   U13198 : NAND2_X1 port map( A1 => n2271, A2 => n7001, ZN => n6995);
   U13199 : NAND2_X1 port map( A1 => n26088, A2 => n2271, ZN => n6994);
   U13202 : XOR2_X1 port map( A1 => Plaintext(54), A2 => Key(54), Z => n16849);
   U13207 : XOR2_X1 port map( A1 => n24747, A2 => n2278, Z => n2699);
   U13209 : OAI21_X2 port map( A1 => n11042, A2 => n24199, B => n24020, ZN => 
                           n2278);
   U13210 : AOI21_X1 port map( A1 => n19038, A2 => n19039, B => n28157, ZN => 
                           n2282);
   U13214 : NAND2_X1 port map( A1 => n2290, A2 => n10845, ZN => n2289);
   U13220 : NAND2_X1 port map( A1 => n12147, A2 => n12148, ZN => n2302);
   U13225 : XOR2_X1 port map( A1 => n21020, A2 => n2306, Z => n2305);
   U13226 : XOR2_X1 port map( A1 => n21019, A2 => n1923, Z => n2306);
   U13235 : INV_X2 port map( I => n2312, ZN => n2450);
   U13236 : INV_X2 port map( I => n2315, ZN => n2378);
   U13237 : MUX2_X1 port map( I0 => n15295, I1 => n18151, S => n2378, Z => 
                           n9198);
   U13240 : OAI21_X2 port map( A1 => n20360, A2 => n2320, B => n2319, ZN => 
                           n20813);
   U13243 : INV_X2 port map( I => n14934, ZN => n21438);
   U13247 : XOR2_X1 port map( A1 => n19772, A2 => n24426, Z => n2333);
   U13248 : XOR2_X1 port map( A1 => n13106, A2 => n31731, Z => n2334);
   U13264 : XOR2_X1 port map( A1 => n7256, A2 => n24763, Z => n24472);
   U13268 : XOR2_X1 port map( A1 => n26623, A2 => n358, Z => n2365);
   U13270 : XOR2_X1 port map( A1 => n2367, A2 => n23151, Z => n2968);
   U13271 : XOR2_X1 port map( A1 => n2367, A2 => n23236, Z => n15374);
   U13279 : OAI21_X1 port map( A1 => n3032, A2 => n6520, B => n2369, ZN => 
                           n2371);
   U13281 : NOR2_X1 port map( A1 => n33566, A2 => n30813, ZN => n12027);
   U13288 : XNOR2_X1 port map( A1 => n10979, A2 => n22028, ZN => n22070);
   U13290 : OR2_X1 port map( A1 => n6798, A2 => n22949, Z => n6675);
   U13298 : XOR2_X1 port map( A1 => n31950, A2 => n1413, Z => n2384);
   U13305 : XOR2_X1 port map( A1 => n19168, A2 => n2389, Z => n5402);
   U13306 : XOR2_X1 port map( A1 => n19484, A2 => n2388, Z => n2389);
   U13317 : NOR2_X1 port map( A1 => n2479, A2 => n22949, ZN => n2405);
   U13324 : XOR2_X1 port map( A1 => n11869, A2 => n14784, Z => n2414);
   U13325 : XOR2_X1 port map( A1 => n20958, A2 => n14785, Z => n2415);
   U13330 : NAND3_X1 port map( A1 => n10046, A2 => n24675, A3 => n23964, ZN => 
                           n2420);
   U13340 : XOR2_X1 port map( A1 => n5875, A2 => n2436, Z => n2435);
   U13344 : NAND2_X2 port map( A1 => n2442, A2 => n2440, ZN => n17385);
   U13345 : AOI21_X1 port map( A1 => n21715, A2 => n21601, B => n21496, ZN => 
                           n2441);
   U13351 : NAND2_X1 port map( A1 => n2449, A2 => n28942, ZN => n10496);
   U13352 : NOR2_X1 port map( A1 => n9224, A2 => n2449, ZN => n9003);
   U13358 : XOR2_X1 port map( A1 => n2045, A2 => n16253, Z => n2452);
   U13359 : XNOR2_X1 port map( A1 => n24810, A2 => n91, ZN => n16002);
   U13370 : INV_X2 port map( I => n2455, ZN => n6976);
   U13371 : NAND2_X2 port map( A1 => n1083, A2 => n18080, ZN => n2456);
   U13375 : XOR2_X1 port map( A1 => n2221, A2 => n6386, Z => n2458);
   U13376 : INV_X2 port map( I => n12617, ZN => n24308);
   U13379 : NAND2_X2 port map( A1 => n2466, A2 => n2464, ZN => n15716);
   U13381 : XOR2_X1 port map( A1 => n4321, A2 => n1069, Z => n2470);
   U13382 : XOR2_X1 port map( A1 => n17830, A2 => n2472, Z => n2473);
   U13383 : XOR2_X1 port map( A1 => n20905, A2 => n25815, Z => n2472);
   U13388 : XOR2_X1 port map( A1 => n20928, A2 => n15, Z => n2476);
   U13389 : INV_X1 port map( I => n22274, ZN => n18058);
   U13394 : NAND2_X1 port map( A1 => n1204, A2 => n6595, ZN => n18215);
   U13401 : NAND2_X1 port map( A1 => n25146, A2 => n5020, ZN => n17525);
   U13402 : XOR2_X1 port map( A1 => n24829, A2 => n5021, Z => n2489);
   U13403 : OAI21_X2 port map( A1 => n17385, A2 => n22099, B => n2490, ZN => 
                           n16971);
   U13404 : NAND2_X2 port map( A1 => n2491, A2 => n21126, ZN => n22099);
   U13408 : NOR2_X2 port map( A1 => n23565, A2 => n23564, ZN => n24150);
   U13409 : NAND2_X1 port map( A1 => n4065, A2 => n25119, ZN => n2498);
   U13410 : NAND2_X1 port map( A1 => n1205, A2 => n254, ZN => n15016);
   U13411 : NAND2_X2 port map( A1 => n2498, A2 => n2497, ZN => n25007);
   U13412 : AND2_X1 port map( A1 => n24885, A2 => n24886, Z => n2497);
   U13415 : XOR2_X1 port map( A1 => n4028, A2 => n19681, Z => n2500);
   U13417 : XOR2_X1 port map( A1 => n19726, A2 => n5081, Z => n2501);
   U13419 : NAND3_X1 port map( A1 => n31074, A2 => n19252, A3 => n1180, ZN => 
                           n2867);
   U13420 : AOI21_X2 port map( A1 => n2794, A2 => n22071, B => n2502, ZN => 
                           n15123);
   U13432 : OAI21_X2 port map( A1 => n911, A2 => n21602, B => n2513, ZN => 
                           n8533);
   U13438 : NAND3_X2 port map( A1 => n11261, A2 => n2519, A3 => n2518, ZN => 
                           n15786);
   U13441 : NAND2_X1 port map( A1 => n8756, A2 => n29309, ZN => n2523);
   U13445 : XOR2_X1 port map( A1 => n1024, A2 => n28864, Z => n2525);
   U13446 : XOR2_X1 port map( A1 => n3351, A2 => n507, Z => n2526);
   U13456 : NAND2_X2 port map( A1 => n2535, A2 => n16951, ZN => n9320);
   U13457 : NOR2_X1 port map( A1 => n10752, A2 => n1826, ZN => n2534);
   U13460 : INV_X2 port map( I => n2978, ZN => n6200);
   U13461 : NAND2_X2 port map( A1 => n5270, A2 => n5271, ZN => n2536);
   U13468 : NAND2_X2 port map( A1 => n29258, A2 => n21462, ZN => n6599);
   U13470 : XOR2_X1 port map( A1 => n2556, A2 => n26124, Z => n3782);
   U13471 : XOR2_X1 port map( A1 => n2557, A2 => n11681, Z => n2556);
   U13474 : XOR2_X1 port map( A1 => n23293, A2 => n1194, Z => n2564);
   U13477 : NOR2_X1 port map( A1 => n7287, A2 => n23057, ZN => n2580);
   U13479 : XOR2_X1 port map( A1 => n15960, A2 => n16657, Z => n11726);
   U13480 : OAI21_X2 port map( A1 => n18841, A2 => n12052, B => n2583, ZN => 
                           n15960);
   U13488 : XOR2_X1 port map( A1 => n20786, A2 => n5414, Z => n2590);
   U13489 : XOR2_X1 port map( A1 => n4681, A2 => n13491, Z => n2591);
   U13495 : NOR2_X1 port map( A1 => n29330, A2 => n13684, ZN => n2960);
   U13496 : NOR2_X1 port map( A1 => n29331, A2 => n13640, ZN => n12885);
   U13499 : OAI22_X1 port map( A1 => n25717, A2 => n29331, B1 => n1076, B2 => 
                           n6915, ZN => n5784);
   U13504 : XOR2_X1 port map( A1 => n17931, A2 => n19719, Z => n2607);
   U13506 : XOR2_X1 port map( A1 => n17430, A2 => n1370, Z => n19719);
   U13507 : XOR2_X1 port map( A1 => n19701, A2 => n467, Z => n2608);
   U13508 : XOR2_X1 port map( A1 => n28822, A2 => n2616, Z => n12673);
   U13511 : OR2_X1 port map( A1 => n31156, A2 => n7394, Z => n2610);
   U13519 : XOR2_X1 port map( A1 => n14588, A2 => n2611, Z => n19519);
   U13521 : NAND2_X1 port map( A1 => n18648, A2 => n18373, ZN => n2613);
   U13522 : NAND2_X1 port map( A1 => n18650, A2 => n2614, ZN => n18549);
   U13530 : XOR2_X1 port map( A1 => n31477, A2 => n16698, Z => n13725);
   U13531 : XOR2_X1 port map( A1 => n31477, A2 => n1416, Z => n9762);
   U13535 : XOR2_X1 port map( A1 => n31908, A2 => n478, Z => n2626);
   U13544 : NAND4_X1 port map( A1 => n5973, A2 => n5971, A3 => n22654, A4 => 
                           n11669, ZN => n2632);
   U13545 : INV_X1 port map( I => n11669, ZN => n2634);
   U13556 : OAI21_X2 port map( A1 => n2646, A2 => n730, B => n26600, ZN => 
                           n3051);
   U13558 : XOR2_X1 port map( A1 => n10522, A2 => n21017, Z => n10437);
   U13559 : NAND2_X2 port map( A1 => n2648, A2 => n2647, ZN => n10522);
   U13564 : XOR2_X1 port map( A1 => n23231, A2 => n540, Z => n2651);
   U13571 : XOR2_X1 port map( A1 => n11636, A2 => n7717, Z => n2661);
   U13581 : XOR2_X1 port map( A1 => n3694, A2 => n7603, Z => n2666);
   U13583 : XOR2_X1 port map( A1 => n7562, A2 => n24769, Z => n2668);
   U13585 : XOR2_X1 port map( A1 => n19712, A2 => n876, Z => n2671);
   U13589 : OAI21_X2 port map( A1 => n19339, A2 => n20000, B => n7327, ZN => 
                           n15005);
   U13590 : NAND2_X1 port map( A1 => n20196, A2 => n2675, ZN => n5103);
   U13598 : OAI21_X1 port map( A1 => n31753, A2 => n18893, B => n11941, ZN => 
                           n2682);
   U13607 : OAI21_X1 port map( A1 => n4045, A2 => n2694, B => n2693, ZN => 
                           n19847);
   U13609 : XOR2_X1 port map( A1 => n2696, A2 => n2695, Z => n8396);
   U13610 : XOR2_X1 port map( A1 => n22268, A2 => n22057, Z => n2695);
   U13612 : XOR2_X1 port map( A1 => n24790, A2 => n1391, Z => n2698);
   U13620 : XOR2_X1 port map( A1 => n22289, A2 => n2707, Z => n2917);
   U13621 : XOR2_X1 port map( A1 => n343, A2 => n1390, Z => n2707);
   U13625 : XOR2_X1 port map( A1 => n2483, A2 => n12719, Z => n12718);
   U13626 : XOR2_X1 port map( A1 => n32822, A2 => n1415, Z => n19427);
   U13648 : OAI21_X2 port map( A1 => n18555, A2 => n3429, B => n2731, ZN => 
                           n9553);
   U13657 : XOR2_X1 port map( A1 => Plaintext(28), A2 => Key(28), Z => n11605);
   U13659 : XOR2_X1 port map( A1 => n4134, A2 => n14668, Z => n2739);
   U13666 : NAND2_X2 port map( A1 => n10710, A2 => n13173, ZN => n13232);
   U13669 : XOR2_X1 port map( A1 => n31755, A2 => n19763, Z => n2747);
   U13675 : NAND2_X2 port map( A1 => n2754, A2 => n2753, ZN => n20921);
   U13683 : XOR2_X1 port map( A1 => n2759, A2 => n2757, Z => n20054);
   U13684 : XOR2_X1 port map( A1 => n19742, A2 => n2758, Z => n2757);
   U13685 : XOR2_X1 port map( A1 => n19768, A2 => n16525, Z => n2758);
   U13701 : XOR2_X1 port map( A1 => n15560, A2 => n624, Z => n10076);
   U13710 : XOR2_X1 port map( A1 => n2786, A2 => n2784, Z => n20882);
   U13716 : XOR2_X1 port map( A1 => n17837, A2 => n24527, Z => n2788);
   U13717 : NAND2_X2 port map( A1 => n2790, A2 => n12536, ZN => n12535);
   U13721 : XOR2_X1 port map( A1 => n19431, A2 => n17104, Z => n19687);
   U13722 : XOR2_X1 port map( A1 => n17835, A2 => n17834, Z => n2796);
   U13723 : XOR2_X1 port map( A1 => n28460, A2 => n16701, Z => n23113);
   U13726 : AOI21_X2 port map( A1 => n24385, A2 => n24384, B => n24383, ZN => 
                           n6484);
   U13729 : NAND2_X1 port map( A1 => n31228, A2 => n27104, ZN => n24384);
   U13739 : XOR2_X1 port map( A1 => n9018, A2 => n23470, Z => n2808);
   U13748 : NOR2_X2 port map( A1 => n2813, A2 => n2844, ZN => n23057);
   U13754 : XOR2_X1 port map( A1 => n9629, A2 => n16551, Z => n2818);
   U13755 : XOR2_X1 port map( A1 => n4134, A2 => n20989, Z => n2819);
   U13760 : NAND3_X2 port map( A1 => n3461, A2 => n3465, A3 => n6536, ZN => 
                           n2989);
   U13764 : AOI21_X1 port map( A1 => n12966, A2 => n28376, B => n2821, ZN => 
                           n20505);
   U13765 : NOR2_X1 port map( A1 => n2822, A2 => n1145, ZN => n21418);
   U13767 : NAND2_X1 port map( A1 => n28017, A2 => n2822, ZN => n7121);
   U13773 : XOR2_X1 port map( A1 => n22126, A2 => n25274, Z => n2825);
   U13784 : XOR2_X1 port map( A1 => n32467, A2 => n25274, Z => n2838);
   U13786 : XOR2_X1 port map( A1 => n2842, A2 => n2840, Z => n16563);
   U13787 : XOR2_X1 port map( A1 => n15055, A2 => n2841, Z => n2840);
   U13791 : NAND3_X1 port map( A1 => n14054, A2 => n15005, A3 => n2843, ZN => 
                           n14546);
   U13794 : XOR2_X1 port map( A1 => n2331, A2 => n34082, Z => n3654);
   U13796 : XOR2_X1 port map( A1 => n34082, A2 => n25619, Z => n19391);
   U13797 : XOR2_X1 port map( A1 => n3653, A2 => n3651, Z => n9469);
   U13815 : NAND2_X1 port map( A1 => n19143, A2 => n2869, ZN => n2868);
   U13819 : NAND3_X1 port map( A1 => n2876, A2 => n25007, A3 => n254, ZN => 
                           n25004);
   U13823 : NAND2_X2 port map( A1 => n3293, A2 => n3292, ZN => n8374);
   U13824 : XOR2_X1 port map( A1 => n2881, A2 => n2880, Z => n2946);
   U13825 : XOR2_X1 port map( A1 => n9569, A2 => n20837, Z => n2880);
   U13826 : XOR2_X1 port map( A1 => n21007, A2 => n21043, Z => n9569);
   U13831 : XOR2_X1 port map( A1 => n20813, A2 => n1193, Z => n2883);
   U13837 : XOR2_X1 port map( A1 => n2891, A2 => n2890, Z => n2889);
   U13838 : XOR2_X1 port map( A1 => n29652, A2 => n24964, Z => n2890);
   U13839 : XOR2_X1 port map( A1 => n9303, A2 => n20926, Z => n2891);
   U13848 : XOR2_X1 port map( A1 => n22158, A2 => n1067, Z => n2898);
   U13849 : XOR2_X1 port map( A1 => n2894, A2 => n4285, Z => n2899);
   U13858 : NOR2_X1 port map( A1 => n2901, A2 => n2902, ZN => n10808);
   U13859 : OAI22_X1 port map( A1 => n26640, A2 => n32253, B1 => n11940, B2 => 
                           n2902, ZN => n19037);
   U13863 : INV_X1 port map( I => n2909, ZN => n25026);
   U13868 : INV_X2 port map( I => n2915, ZN => n13998);
   U13871 : XOR2_X1 port map( A1 => n22118, A2 => n22115, Z => n2918);
   U13874 : XOR2_X1 port map( A1 => n2920, A2 => n16697, Z => n19442);
   U13879 : XOR2_X1 port map( A1 => n20974, A2 => n2925, Z => n2924);
   U13882 : XOR2_X1 port map( A1 => n20743, A2 => n8774, Z => n2926);
   U13891 : INV_X2 port map( I => n2946, ZN => n21237);
   U13898 : XOR2_X1 port map( A1 => n13908, A2 => n13909, Z => n2952);
   U13907 : NAND2_X1 port map( A1 => n868, A2 => n2958, ZN => n15951);
   U13911 : AOI21_X1 port map( A1 => n25732, A2 => n6915, B => n2959, ZN => 
                           n5838);
   U13912 : NOR2_X1 port map( A1 => n13124, A2 => n2960, ZN => n2959);
   U13915 : NOR2_X2 port map( A1 => n13637, A2 => n13636, ZN => n13640);
   U13926 : XOR2_X1 port map( A1 => n2972, A2 => n2975, Z => n8634);
   U13930 : XOR2_X1 port map( A1 => n30041, A2 => n23387, Z => n23522);
   U13931 : XOR2_X1 port map( A1 => n13190, A2 => n17704, Z => n2975);
   U13933 : NAND2_X2 port map( A1 => n3658, A2 => n4982, ZN => n23441);
   U13939 : OAI21_X2 port map( A1 => n8867, A2 => n8864, B => n8863, ZN => 
                           n19484);
   U13941 : NAND2_X2 port map( A1 => n18717, A2 => n17617, ZN => n19470);
   U13943 : OAI22_X1 port map( A1 => n25006, A2 => n3019, B1 => n2983, B2 => 
                           n14865, ZN => n25008);
   U13952 : NOR2_X1 port map( A1 => n9090, A2 => n27142, ZN => n2986);
   U13953 : XOR2_X1 port map( A1 => n2989, A2 => n25722, Z => n20644);
   U13956 : INV_X2 port map( I => n11599, ZN => n11941);
   U13968 : NAND2_X1 port map( A1 => n11680, A2 => n1331, ZN => n3003);
   U13978 : XOR2_X1 port map( A1 => n6484, A2 => n7256, Z => n17571);
   U13979 : INV_X2 port map( I => n3012, ZN => n8370);
   U13980 : NAND4_X1 port map( A1 => n24333, A2 => n24334, A3 => n24332, A4 => 
                           n3014, ZN => n24336);
   U13984 : NAND2_X2 port map( A1 => n24880, A2 => n24879, ZN => n3019);
   U13990 : NOR2_X2 port map( A1 => n24083, A2 => n24082, ZN => n24753);
   U13993 : NOR2_X2 port map( A1 => n3024, A2 => n3023, ZN => n9885);
   U13995 : XOR2_X1 port map( A1 => n33293, A2 => n3027, Z => n3026);
   U13996 : XOR2_X1 port map( A1 => n7229, A2 => n30320, Z => n3028);
   U13999 : INV_X1 port map( I => n3033, ZN => n15013);
   U14008 : NAND2_X1 port map( A1 => n3049, A2 => n3048, ZN => n3047);
   U14018 : NOR2_X1 port map( A1 => n20196, A2 => n295, ZN => n3068);
   U14020 : XOR2_X1 port map( A1 => n19549, A2 => n3071, Z => n3070);
   U14021 : XOR2_X1 port map( A1 => n19550, A2 => n25049, Z => n3071);
   U14023 : XOR2_X1 port map( A1 => n19699, A2 => n7971, Z => n19549);
   U14028 : NAND2_X2 port map( A1 => n16363, A2 => n19131, ZN => n16727);
   U14029 : XOR2_X1 port map( A1 => n19661, A2 => n19580, Z => n19551);
   U14038 : XOR2_X1 port map( A1 => n3081, A2 => n3082, Z => n23586);
   U14043 : XOR2_X1 port map( A1 => n1262, A2 => n27186, Z => n3083);
   U14050 : XOR2_X1 port map( A1 => n20984, A2 => n20986, Z => n3099);
   U14051 : XOR2_X1 port map( A1 => n17377, A2 => n3101, Z => n3100);
   U14052 : XOR2_X1 port map( A1 => n12495, A2 => n21985, Z => n3102);
   U14059 : OAI21_X1 port map( A1 => n17640, A2 => n26677, B => n4971, ZN => 
                           n3105);
   U14068 : XOR2_X1 port map( A1 => n10443, A2 => n32880, Z => n3109);
   U14074 : INV_X1 port map( I => n20781, ZN => n20867);
   U14078 : XOR2_X1 port map( A1 => n17517, A2 => n16390, Z => n3118);
   U14079 : XOR2_X1 port map( A1 => n21019, A2 => n15275, Z => n3119);
   U14081 : XOR2_X1 port map( A1 => n22203, A2 => n10165, Z => n3120);
   U14091 : XNOR2_X1 port map( A1 => n23200, A2 => n7772, ZN => n23165);
   U14092 : XOR2_X1 port map( A1 => n33465, A2 => n14435, Z => n3126);
   U14096 : INV_X2 port map( I => n19222, ZN => n15137);
   U14102 : XOR2_X1 port map( A1 => n3134, A2 => n24964, Z => Ciphertext(18));
   U14107 : XOR2_X1 port map( A1 => n22030, A2 => n22031, Z => n3142);
   U14108 : XOR2_X1 port map( A1 => n16321, A2 => n16472, Z => n24595);
   U14109 : XOR2_X1 port map( A1 => n16321, A2 => n1417, Z => n24357);
   U14111 : XOR2_X1 port map( A1 => n15308, A2 => n17384, Z => n3143);
   U14116 : NAND3_X1 port map( A1 => n3148, A2 => n24268, A3 => n31228, ZN => 
                           n23996);
   U14119 : XOR2_X1 port map( A1 => n20772, A2 => n3158, Z => n4246);
   U14120 : XOR2_X1 port map( A1 => n32399, A2 => n20992, Z => n3158);
   U14126 : XOR2_X1 port map( A1 => n17519, A2 => n3164, Z => n14494);
   U14127 : XOR2_X1 port map( A1 => n29011, A2 => n8356, Z => n3164);
   U14128 : NAND2_X1 port map( A1 => n29043, A2 => n3165, ZN => n17588);
   U14137 : XOR2_X1 port map( A1 => n7987, A2 => n6464, Z => n10791);
   U14140 : NAND2_X1 port map( A1 => n24780, A2 => n24874, ZN => n24604);
   U14141 : XOR2_X1 port map( A1 => n32467, A2 => n21037, Z => n12171);
   U14143 : XOR2_X1 port map( A1 => n22143, A2 => n21984, Z => n3175);
   U14145 : XOR2_X1 port map( A1 => n27240, A2 => n13091, Z => n3177);
   U14147 : NAND2_X1 port map( A1 => n8125, A2 => n3181, ZN => n17589);
   U14149 : AND2_X1 port map( A1 => n22537, A2 => n28170, Z => n3189);
   U14151 : XOR2_X1 port map( A1 => n21038, A2 => n6872, Z => n3190);
   U14152 : XOR2_X1 port map( A1 => n21039, A2 => n586, Z => n3191);
   U14155 : XOR2_X1 port map( A1 => n3194, A2 => n19413, Z => n19414);
   U14157 : XOR2_X1 port map( A1 => n11422, A2 => n22194, Z => n11421);
   U14161 : NOR2_X1 port map( A1 => n10831, A2 => n19856, ZN => n3197);
   U14162 : XOR2_X1 port map( A1 => n3199, A2 => n3198, Z => n13298);
   U14163 : XOR2_X1 port map( A1 => n13236, A2 => n1420, Z => n3198);
   U14164 : XOR2_X1 port map( A1 => n28579, A2 => n28939, Z => n3199);
   U14168 : NAND2_X1 port map( A1 => n30678, A2 => n3203, ZN => n21536);
   U14172 : NAND2_X1 port map( A1 => n24260, A2 => n30280, ZN => n16573);
   U14188 : AOI21_X1 port map( A1 => n18891, A2 => n18676, B => n3218, ZN => 
                           n12198);
   U14189 : NOR2_X1 port map( A1 => n11398, A2 => n3218, ZN => n11397);
   U14190 : AOI21_X1 port map( A1 => n3586, A2 => n14874, B => n3218, ZN => 
                           n3516);
   U14194 : NOR2_X1 port map( A1 => n9162, A2 => n9164, ZN => n3224);
   U14200 : OAI21_X2 port map( A1 => n17906, A2 => n3240, B => n3239, ZN => 
                           n24242);
   U14202 : NAND2_X2 port map( A1 => n5083, A2 => n3242, ZN => n6387);
   U14203 : NAND3_X2 port map( A1 => n3245, A2 => n19173, A3 => n19172, ZN => 
                           n19473);
   U14208 : NAND2_X1 port map( A1 => n12508, A2 => n6111, ZN => n25572);
   U14213 : XOR2_X1 port map( A1 => n1363, A2 => n3258, Z => n3358);
   U14214 : XOR2_X1 port map( A1 => n3260, A2 => n3259, Z => n3258);
   U14217 : XOR2_X1 port map( A1 => n23399, A2 => n23398, Z => n3267);
   U14220 : NAND2_X1 port map( A1 => n4663, A2 => n31742, ZN => n3271);
   U14238 : XOR2_X1 port map( A1 => n11604, A2 => n34082, Z => n19591);
   U14242 : XOR2_X1 port map( A1 => n17912, A2 => n1084, Z => n24401);
   U14247 : INV_X2 port map( I => n23853, ZN => n8614);
   U14251 : OAI21_X2 port map( A1 => n2537, A2 => n1300, B => n6685, ZN => 
                           n22856);
   U14254 : NAND3_X2 port map( A1 => n25342, A2 => n25341, A3 => n25340, ZN => 
                           n3300);
   U14255 : NOR2_X1 port map( A1 => n3300, A2 => n25367, ZN => n25362);
   U14256 : AOI21_X1 port map( A1 => n25367, A2 => n25368, B => n3300, ZN => 
                           n25350);
   U14257 : NOR2_X1 port map( A1 => n18711, A2 => n27142, ZN => n11269);
   U14262 : XOR2_X1 port map( A1 => n3350, A2 => n1407, Z => n20621);
   U14263 : XOR2_X1 port map( A1 => n3350, A2 => n7705, Z => n20798);
   U14264 : XOR2_X1 port map( A1 => n3350, A2 => n30543, Z => n13093);
   U14266 : INV_X2 port map( I => n13189, ZN => n15522);
   U14272 : XOR2_X1 port map( A1 => n438, A2 => n32796, Z => n3319);
   U14276 : OAI21_X2 port map( A1 => n3324, A2 => n29232, B => n11865, ZN => 
                           n15243);
   U14279 : XOR2_X1 port map( A1 => n30041, A2 => n14613, Z => n13777);
   U14288 : NAND2_X1 port map( A1 => n18538, A2 => n3344, ZN => n14327);
   U14291 : XOR2_X1 port map( A1 => n3345, A2 => n31416, Z => n24552);
   U14292 : XOR2_X1 port map( A1 => n33700, A2 => n24804, Z => n14532);
   U14296 : NAND2_X2 port map( A1 => n4234, A2 => n13113, ZN => n21839);
   U14298 : XOR2_X1 port map( A1 => n3355, A2 => n3354, Z => n3353);
   U14299 : XOR2_X1 port map( A1 => n29121, A2 => n1421, Z => n3354);
   U14300 : XOR2_X1 port map( A1 => n12789, A2 => n7808, Z => n3355);
   U14302 : OAI21_X2 port map( A1 => n7516, A2 => n10125, B => n3361, ZN => 
                           n10124);
   U14305 : XOR2_X1 port map( A1 => n22187, A2 => n3369, Z => n3368);
   U14306 : XOR2_X1 port map( A1 => n16060, A2 => n25910, Z => n3369);
   U14309 : NAND3_X2 port map( A1 => n3384, A2 => n32031, A3 => n3382, ZN => 
                           n6798);
   U14314 : INV_X2 port map( I => n3392, ZN => n4396);
   U14316 : XOR2_X1 port map( A1 => n30571, A2 => n27920, Z => n3396);
   U14319 : XOR2_X1 port map( A1 => n19716, A2 => n10123, Z => n3399);
   U14324 : XOR2_X1 port map( A1 => n21045, A2 => n20967, Z => n4260);
   U14327 : NOR2_X1 port map( A1 => n3405, A2 => n25564, ZN => n24460);
   U14332 : OAI21_X2 port map( A1 => n1260, A2 => n9843, B => n3408, ZN => 
                           n4955);
   U14336 : XOR2_X1 port map( A1 => n4955, A2 => n23386, Z => n3410);
   U14337 : XOR2_X1 port map( A1 => n3412, A2 => n537, Z => n3411);
   U14338 : XOR2_X1 port map( A1 => n27220, A2 => n5514, Z => n3412);
   U14342 : XOR2_X1 port map( A1 => n26623, A2 => n25218, Z => n3415);
   U14346 : XOR2_X1 port map( A1 => n13477, A2 => n3417, Z => n19705);
   U14348 : XOR2_X1 port map( A1 => n22119, A2 => n30993, Z => n22120);
   U14355 : AND2_X1 port map( A1 => n20419, A2 => n15005, Z => n3428);
   U14356 : INV_X1 port map( I => n3430, ZN => n10745);
   U14357 : XOR2_X1 port map( A1 => n3431, A2 => n25192, Z => Ciphertext(68));
   U14358 : OAI21_X1 port map( A1 => n10574, A2 => n27149, B => n3433, ZN => 
                           n3432);
   U14372 : NOR2_X1 port map( A1 => n632, A2 => n14339, ZN => n3502);
   U14374 : MUX2_X1 port map( I0 => n809, I1 => n30065, S => n14227, Z => 
                           n22448);
   U14376 : XOR2_X1 port map( A1 => n24749, A2 => n3477, Z => n3476);
   U14377 : XOR2_X1 port map( A1 => n24839, A2 => n25864, Z => n3477);
   U14389 : NOR2_X1 port map( A1 => n30318, A2 => n3489, ZN => n5301);
   U14390 : NAND2_X1 port map( A1 => n5408, A2 => n3489, ZN => n5407);
   U14394 : XOR2_X1 port map( A1 => n16998, A2 => n18015, Z => n3493);
   U14396 : NAND2_X1 port map( A1 => n26292, A2 => n3495, ZN => n11420);
   U14399 : NAND2_X1 port map( A1 => n31197, A2 => n32898, ZN => n3497);
   U14404 : XOR2_X1 port map( A1 => n10422, A2 => n10421, Z => n16710);
   U14410 : XOR2_X1 port map( A1 => n3514, A2 => n23535, Z => n9983);
   U14418 : XOR2_X1 port map( A1 => n23183, A2 => n26656, Z => n23494);
   U14435 : NAND3_X1 port map( A1 => n21781, A2 => n31220, A3 => n3539, ZN => 
                           n21746);
   U14439 : XOR2_X1 port map( A1 => n11217, A2 => n3541, Z => n3540);
   U14440 : XOR2_X1 port map( A1 => n17301, A2 => n8139, Z => n3541);
   U14442 : XOR2_X1 port map( A1 => n5932, A2 => n24652, Z => n24824);
   U14449 : XOR2_X1 port map( A1 => n20747, A2 => n1191, Z => n3559);
   U14454 : NAND2_X1 port map( A1 => n3567, A2 => n31019, ZN => n17631);
   U14456 : NOR2_X1 port map( A1 => n22406, A2 => n3567, ZN => n3566);
   U14457 : INV_X1 port map( I => n3569, ZN => n12159);
   U14458 : NAND3_X1 port map( A1 => n3570, A2 => n22982, A3 => n22983, ZN => 
                           n22984);
   U14460 : NOR2_X1 port map( A1 => n22800, A2 => n3570, ZN => n13045);
   U14465 : XOR2_X1 port map( A1 => n23375, A2 => n23294, Z => n23240);
   U14466 : NAND2_X2 port map( A1 => n16993, A2 => n11837, ZN => n23294);
   U14468 : NAND2_X2 port map( A1 => n15208, A2 => n17175, ZN => n16373);
   U14470 : XOR2_X1 port map( A1 => n23343, A2 => n3575, Z => n3574);
   U14471 : XOR2_X1 port map( A1 => n15183, A2 => n16602, Z => n3575);
   U14483 : XOR2_X1 port map( A1 => n22139, A2 => n16390, Z => n3583);
   U14487 : XOR2_X1 port map( A1 => n27186, A2 => n12797, Z => n10776);
   U14488 : XOR2_X1 port map( A1 => n27186, A2 => n9223, Z => n7131);
   U14491 : AOI21_X2 port map( A1 => n19074, A2 => n29398, B => n19073, ZN => 
                           n3599);
   U14497 : XOR2_X1 port map( A1 => n17918, A2 => n3606, Z => n3605);
   U14498 : XOR2_X1 port map( A1 => n8617, A2 => n16525, Z => n3606);
   U14500 : XOR2_X1 port map( A1 => n33468, A2 => n16598, Z => n12624);
   U14508 : INV_X2 port map( I => n20788, ZN => n20907);
   U14511 : XOR2_X1 port map( A1 => n3621, A2 => n3622, Z => n3618);
   U14514 : XOR2_X1 port map( A1 => n23461, A2 => n23321, Z => n3620);
   U14516 : XOR2_X1 port map( A1 => n30322, A2 => n15114, Z => n3622);
   U14520 : XOR2_X1 port map( A1 => n3628, A2 => n20894, Z => n3627);
   U14521 : XOR2_X1 port map( A1 => n20992, A2 => n1069, Z => n3628);
   U14527 : XOR2_X1 port map( A1 => n3634, A2 => n25541, Z => n9269);
   U14543 : XOR2_X1 port map( A1 => n11762, A2 => n10278, Z => n3648);
   U14544 : XOR2_X1 port map( A1 => n3652, A2 => n18031, Z => n3651);
   U14545 : XOR2_X1 port map( A1 => n3815, A2 => n3654, Z => n3653);
   U14546 : AOI21_X1 port map( A1 => n17055, A2 => n15475, B => n25996, ZN => 
                           n15474);
   U14549 : MUX2_X1 port map( I0 => n30769, I1 => n30885, S => n21697, Z => 
                           n3656);
   U14550 : NAND2_X2 port map( A1 => n18136, A2 => n12133, ZN => n21697);
   U14553 : AND2_X1 port map( A1 => n33627, A2 => n29446, Z => n4301);
   U14555 : XOR2_X1 port map( A1 => n19620, A2 => n5919, Z => n3665);
   U14561 : NAND2_X1 port map( A1 => n5821, A2 => n3668, ZN => n22750);
   U14571 : XOR2_X1 port map( A1 => n24552, A2 => n3677, Z => n4302);
   U14572 : XOR2_X1 port map( A1 => n8949, A2 => n5268, Z => n3677);
   U14576 : XOR2_X1 port map( A1 => n21945, A2 => n3682, Z => n3683);
   U14577 : INV_X2 port map( I => n3686, ZN => n9172);
   U14578 : NOR2_X1 port map( A1 => n17694, A2 => n3687, ZN => n13879);
   U14579 : NAND2_X2 port map( A1 => n22496, A2 => n22495, ZN => n14686);
   U14585 : XOR2_X1 port map( A1 => n3694, A2 => n2864, Z => n9093);
   U14591 : XOR2_X1 port map( A1 => n3704, A2 => n17555, Z => n22300);
   U14594 : XOR2_X1 port map( A1 => n9536, A2 => n3704, Z => n9532);
   U14597 : XOR2_X1 port map( A1 => n12342, A2 => n3705, Z => n20242);
   U14598 : XOR2_X1 port map( A1 => n20726, A2 => n3705, Z => n21027);
   U14599 : NAND2_X2 port map( A1 => n15142, A2 => n20237, ZN => n3705);
   U14609 : OAI21_X2 port map( A1 => n11991, A2 => n918, B => n11856, ZN => 
                           n3723);
   U14617 : XOR2_X1 port map( A1 => n3727, A2 => n19679, Z => n9819);
   U14618 : NAND2_X1 port map( A1 => n5433, A2 => n502, ZN => n4841);
   U14620 : NAND2_X2 port map( A1 => n3730, A2 => n3728, ZN => n6402);
   U14621 : INV_X2 port map( I => n18080, ZN => n25236);
   U14623 : XOR2_X1 port map( A1 => n30219, A2 => n24231, Z => n3735);
   U14624 : XOR2_X1 port map( A1 => n14858, A2 => n16173, Z => n12618);
   U14625 : XOR2_X1 port map( A1 => n20870, A2 => n3737, Z => n3736);
   U14626 : XOR2_X1 port map( A1 => n21040, A2 => n5772, Z => n3737);
   U14634 : XOR2_X1 port map( A1 => n24469, A2 => n17753, Z => n17752);
   U14639 : AOI22_X2 port map( A1 => n24378, A2 => n14547, B1 => n25753, B2 => 
                           n25581, ZN => n25746);
   U14643 : NOR2_X1 port map( A1 => n12906, A2 => n12948, ZN => n9391);
   U14647 : NAND2_X2 port map( A1 => n23792, A2 => n23791, ZN => n12493);
   U14654 : INV_X2 port map( I => n3755, ZN => n10182);
   U14655 : XOR2_X1 port map( A1 => Plaintext(174), A2 => Key(174), Z => n3755)
                           ;
   U14657 : XOR2_X1 port map( A1 => n4240, A2 => n16642, Z => n24794);
   U14663 : NOR3_X2 port map( A1 => n26025, A2 => n15466, A3 => n14098, ZN => 
                           n8530);
   U14667 : XOR2_X1 port map( A1 => n17524, A2 => n20514, Z => n21442);
   U14673 : NAND2_X2 port map( A1 => n20651, A2 => n20650, ZN => n20769);
   U14674 : AOI21_X2 port map( A1 => n2565, A2 => n20438, B => n17424, ZN => 
                           n20651);
   U14679 : NAND2_X1 port map( A1 => n20501, A2 => n20502, ZN => n16758);
   U14682 : OAI21_X1 port map( A1 => n25349, A2 => n25360, B => n25379, ZN => 
                           n3771);
   U14683 : OR2_X1 port map( A1 => n25350, A2 => n25361, Z => n3772);
   U14686 : XOR2_X1 port map( A1 => n24848, A2 => n17448, Z => n5022);
   U14693 : XOR2_X1 port map( A1 => n4915, A2 => n23245, Z => n3777);
   U14694 : NAND2_X1 port map( A1 => n4066, A2 => n14811, ZN => n16007);
   U14695 : OAI21_X2 port map( A1 => n4178, A2 => n5752, B => n5751, ZN => 
                           n4066);
   U14696 : XNOR2_X1 port map( A1 => n13309, A2 => n11803, ZN => n4004);
   U14705 : INV_X2 port map( I => n3782, ZN => n11820);
   U14707 : AND2_X1 port map( A1 => n25174, A2 => n25175, Z => n8931);
   U14708 : NAND2_X2 port map( A1 => n25172, A2 => n25169, ZN => n25174);
   U14718 : NAND2_X1 port map( A1 => n3788, A2 => n1425, ZN => n14295);
   U14730 : XOR2_X1 port map( A1 => Plaintext(116), A2 => Key(116), Z => n18131
                           );
   U14731 : XOR2_X1 port map( A1 => n23220, A2 => n23198, Z => n11144);
   U14736 : OAI21_X1 port map( A1 => n14830, A2 => n22636, B => n12043, ZN => 
                           n22495);
   U14748 : XOR2_X1 port map( A1 => n8656, A2 => n24050, Z => n9968);
   U14757 : XOR2_X1 port map( A1 => n9200, A2 => n660, Z => n9199);
   U14759 : XOR2_X1 port map( A1 => n23189, A2 => n4409, Z => n23465);
   U14761 : XOR2_X1 port map( A1 => n24533, A2 => n27950, Z => n16891);
   U14762 : AND2_X1 port map( A1 => n23660, A2 => n30252, Z => n4350);
   U14766 : NAND2_X1 port map( A1 => n32884, A2 => n32798, ZN => n15867);
   U14771 : XOR2_X1 port map( A1 => n24439, A2 => n3809, Z => n11527);
   U14772 : XOR2_X1 port map( A1 => n24592, A2 => n25364, Z => n3809);
   U14780 : INV_X2 port map( I => n3816, ZN => n11333);
   U14783 : NAND2_X1 port map( A1 => n9469, A2 => n563, ZN => n12119);
   U14784 : XOR2_X1 port map( A1 => n3819, A2 => n12672, Z => n8545);
   U14785 : XOR2_X1 port map( A1 => n20796, A2 => n20797, Z => n3819);
   U14786 : XOR2_X1 port map( A1 => n21025, A2 => n6561, Z => n6560);
   U14789 : NAND2_X2 port map( A1 => n9237, A2 => n9238, ZN => n14293);
   U14794 : AOI21_X1 port map( A1 => n832, A2 => n27189, B => n7038, ZN => 
                           n7037);
   U14797 : OAI21_X2 port map( A1 => n14693, A2 => n19889, B => n3827, ZN => 
                           n20485);
   U14801 : XNOR2_X1 port map( A1 => n11481, A2 => n5848, ZN => n9673);
   U14803 : XOR2_X1 port map( A1 => n15708, A2 => n19552, Z => n19555);
   U14823 : XOR2_X1 port map( A1 => n23370, A2 => n16300, Z => n6152);
   U14824 : XOR2_X1 port map( A1 => n8630, A2 => n22301, Z => n12828);
   U14825 : XOR2_X1 port map( A1 => n4723, A2 => n15825, Z => n22301);
   U14826 : NAND2_X1 port map( A1 => n21594, A2 => n21145, ZN => n21156);
   U14828 : NOR2_X1 port map( A1 => n6778, A2 => n33621, ZN => n6579);
   U14837 : OAI21_X2 port map( A1 => n15675, A2 => n6009, B => n3920, ZN => 
                           n19778);
   U14863 : NOR2_X1 port map( A1 => n13733, A2 => n24229, ZN => n13732);
   U14864 : XOR2_X1 port map( A1 => n23315, A2 => n13812, Z => n11416);
   U14866 : XOR2_X1 port map( A1 => n20600, A2 => n5209, Z => n16239);
   U14869 : NAND2_X2 port map( A1 => n414, A2 => n5834, ZN => n18682);
   U14887 : XOR2_X1 port map( A1 => n23385, A2 => n17188, Z => n23284);
   U14893 : NAND2_X2 port map( A1 => n6206, A2 => n6570, ZN => n6571);
   U14897 : XOR2_X1 port map( A1 => n14908, A2 => n26623, Z => n3870);
   U14900 : OR2_X1 port map( A1 => n24712, A2 => n4490, Z => n4451);
   U14904 : XOR2_X1 port map( A1 => n11221, A2 => n11220, Z => n19958);
   U14905 : NAND2_X2 port map( A1 => n21827, A2 => n21824, ZN => n5170);
   U14912 : XNOR2_X1 port map( A1 => n23203, A2 => n24917, ZN => n4466);
   U14913 : NAND2_X1 port map( A1 => n23690, A2 => n23856, ZN => n17056);
   U14921 : XOR2_X1 port map( A1 => n3884, A2 => n14206, Z => n14296);
   U14922 : NAND2_X1 port map( A1 => n14295, A2 => n14294, ZN => n3884);
   U14924 : XOR2_X1 port map( A1 => n12491, A2 => n30320, Z => n9012);
   U14928 : INV_X1 port map( I => n4342, ZN => n22188);
   U14932 : AOI21_X2 port map( A1 => n18334, A2 => n3893, B => n18333, ZN => 
                           n16847);
   U14933 : XOR2_X1 port map( A1 => n7184, A2 => n446, Z => n16105);
   U14943 : XOR2_X1 port map( A1 => n17565, A2 => n23320, Z => n23194);
   U14946 : XOR2_X1 port map( A1 => n10200, A2 => n3896, Z => n17779);
   U14947 : XOR2_X1 port map( A1 => n14779, A2 => n24098, Z => n3896);
   U14948 : NAND2_X2 port map( A1 => n7770, A2 => n7768, ZN => n25107);
   U14955 : NAND3_X2 port map( A1 => n3900, A2 => n5333, A3 => n19136, ZN => 
                           n19773);
   U14956 : INV_X1 port map( I => n23446, ZN => n17350);
   U14959 : AND2_X1 port map( A1 => n4405, A2 => n7810, Z => n19174);
   U14961 : XOR2_X1 port map( A1 => n3905, A2 => n17457, Z => n8834);
   U14963 : AND2_X1 port map( A1 => n6483, A2 => n3467, Z => n8970);
   U14971 : NAND2_X2 port map( A1 => n3908, A2 => n12939, ZN => n22291);
   U14973 : NAND2_X1 port map( A1 => n19863, A2 => n10335, ZN => n7922);
   U14974 : XOR2_X1 port map( A1 => n9326, A2 => n9325, Z => n10335);
   U14979 : INV_X1 port map( I => n25882, ZN => n7274);
   U14980 : AND2_X1 port map( A1 => n25882, A2 => n25879, Z => n7268);
   U14985 : XNOR2_X1 port map( A1 => n21281, A2 => n21280, ZN => n9593);
   U14992 : NOR2_X1 port map( A1 => n19799, A2 => n16625, ZN => n19800);
   U14995 : INV_X2 port map( I => n9992, ZN => n11887);
   U14998 : NAND2_X2 port map( A1 => n13461, A2 => n13462, ZN => n23066);
   U15004 : XOR2_X1 port map( A1 => n23220, A2 => n3923, Z => n8488);
   U15005 : XOR2_X1 port map( A1 => n27252, A2 => n31354, Z => n3923);
   U15006 : XNOR2_X1 port map( A1 => n15341, A2 => n27763, ZN => n14733);
   U15010 : NOR2_X1 port map( A1 => n21066, A2 => n31965, ZN => n6213);
   U15012 : XNOR2_X1 port map( A1 => n28262, A2 => n16551, ZN => n10878);
   U15018 : NAND2_X1 port map( A1 => n8966, A2 => n3926, ZN => n14465);
   U15019 : AOI21_X1 port map( A1 => n5035, A2 => n6593, B => n22957, ZN => 
                           n3926);
   U15021 : NAND2_X2 port map( A1 => n23989, A2 => n13144, ZN => n7511);
   U15025 : NOR2_X1 port map( A1 => n5842, A2 => n18945, ZN => n18946);
   U15027 : NAND2_X2 port map( A1 => n24217, A2 => n29010, ZN => n23964);
   U15028 : NAND2_X2 port map( A1 => n14966, A2 => n14965, ZN => n6906);
   U15035 : XOR2_X1 port map( A1 => n5881, A2 => n3938, Z => n5880);
   U15036 : XOR2_X1 port map( A1 => n5882, A2 => n524, Z => n3938);
   U15067 : NAND2_X1 port map( A1 => n6234, A2 => n694, ZN => n16661);
   U15071 : XOR2_X1 port map( A1 => Plaintext(9), A2 => Key(9), Z => n3954);
   U15072 : AOI21_X1 port map( A1 => n5113, A2 => n24994, B => n9901, ZN => 
                           n9903);
   U15074 : INV_X2 port map( I => n10725, ZN => n16166);
   U15078 : XOR2_X1 port map( A1 => n24846, A2 => n7256, Z => n24849);
   U15082 : XOR2_X1 port map( A1 => n20757, A2 => n20712, Z => n20713);
   U15085 : XOR2_X1 port map( A1 => n10109, A2 => n15562, Z => n3957);
   U15086 : XOR2_X1 port map( A1 => n3958, A2 => n9487, Z => n9486);
   U15087 : XOR2_X1 port map( A1 => n24778, A2 => n550, Z => n3958);
   U15088 : XOR2_X1 port map( A1 => n20852, A2 => n10159, Z => n15630);
   U15090 : OAI22_X2 port map( A1 => n21602, A2 => n21716, B1 => n21710, B2 => 
                           n21712, ZN => n6462);
   U15093 : XOR2_X1 port map( A1 => n6169, A2 => n15653, Z => n16300);
   U15104 : OAI22_X2 port map( A1 => n3963, A2 => n21298, B1 => n4989, B2 => 
                           n21199, ZN => n21870);
   U15106 : XOR2_X1 port map( A1 => n24634, A2 => n24494, Z => n10945);
   U15108 : XOR2_X1 port map( A1 => n20899, A2 => n9706, Z => n10951);
   U15114 : NAND2_X2 port map( A1 => n964, A2 => n5072, ZN => n9481);
   U15124 : OAI22_X2 port map( A1 => n19060, A2 => n1179, B1 => n4366, B2 => 
                           n16185, ZN => n4150);
   U15137 : NAND2_X1 port map( A1 => n22832, A2 => n13635, ZN => n12156);
   U15140 : XOR2_X1 port map( A1 => n16259, A2 => n23433, Z => n17285);
   U15146 : XOR2_X1 port map( A1 => n9528, A2 => n3980, Z => n10934);
   U15148 : XOR2_X1 port map( A1 => n3981, A2 => n444, Z => n5074);
   U15149 : XOR2_X1 port map( A1 => n4984, A2 => n15788, Z => n3981);
   U15150 : INV_X1 port map( I => n19523, ZN => n20141);
   U15151 : NAND2_X1 port map( A1 => n27110, A2 => n15237, ZN => n19523);
   U15157 : AND2_X1 port map( A1 => n10182, A2 => n11460, Z => n18877);
   U15159 : OR2_X1 port map( A1 => n7465, A2 => n13334, Z => n5490);
   U15165 : NAND2_X2 port map( A1 => n3985, A2 => n12814, ZN => n16699);
   U15169 : XOR2_X1 port map( A1 => n20752, A2 => n3990, Z => n18050);
   U15170 : XOR2_X1 port map( A1 => n4618, A2 => n24804, Z => n3990);
   U15180 : OAI21_X2 port map( A1 => n3996, A2 => n3995, B => n4675, ZN => 
                           n24002);
   U15181 : OR2_X1 port map( A1 => n4734, A2 => n23065, Z => n3997);
   U15186 : XOR2_X1 port map( A1 => n20759, A2 => n16191, Z => n4000);
   U15197 : AND2_X1 port map( A1 => n1278, A2 => n15633, Z => n12218);
   U15209 : OR2_X1 port map( A1 => n1430, A2 => n10080, Z => n4008);
   U15212 : XOR2_X1 port map( A1 => n4013, A2 => n13067, Z => n10186);
   U15216 : INV_X1 port map( I => n24870, ZN => n16607);
   U15217 : XOR2_X1 port map( A1 => n4015, A2 => n9607, Z => n9606);
   U15218 : XOR2_X1 port map( A1 => n9608, A2 => n21007, Z => n4015);
   U15229 : XOR2_X1 port map( A1 => n5939, A2 => n14122, Z => n4020);
   U15238 : XOR2_X1 port map( A1 => n30327, A2 => n5539, Z => n14779);
   U15240 : NAND2_X2 port map( A1 => n4628, A2 => n4629, ZN => n4599);
   U15249 : XOR2_X1 port map( A1 => n4035, A2 => n16423, Z => Ciphertext(29));
   U15259 : AOI22_X1 port map( A1 => n17165, A2 => n17687, B1 => n17166, B2 => 
                           n18863, ZN => n12193);
   U15261 : NOR2_X2 port map( A1 => n19816, A2 => n19817, ZN => n20595);
   U15262 : OR2_X1 port map( A1 => n10413, A2 => n19891, Z => n17443);
   U15268 : XOR2_X1 port map( A1 => n19695, A2 => n4042, Z => n20088);
   U15269 : XOR2_X1 port map( A1 => n19693, A2 => n19694, Z => n4042);
   U15286 : XOR2_X1 port map( A1 => n4052, A2 => n496, Z => n8684);
   U15294 : XOR2_X1 port map( A1 => n21035, A2 => n1409, Z => n20929);
   U15299 : XOR2_X1 port map( A1 => n23124, A2 => n481, Z => n4059);
   U15303 : OR2_X1 port map( A1 => n21707, A2 => n230, Z => n14461);
   U15309 : NAND2_X2 port map( A1 => n5801, A2 => n4062, ZN => n4646);
   U15311 : XOR2_X1 port map( A1 => n4063, A2 => n27126, Z => n7381);
   U15315 : NAND2_X1 port map( A1 => n24882, A2 => n25117, ZN => n4065);
   U15337 : NOR2_X1 port map( A1 => n14544, A2 => n14543, ZN => n10128);
   U15339 : NAND2_X1 port map( A1 => n4177, A2 => n23855, ZN => n23800);
   U15340 : OAI21_X2 port map( A1 => n8800, A2 => n18925, B => n18924, ZN => 
                           n19632);
   U15342 : AND2_X1 port map( A1 => n23949, A2 => n11676, Z => n9002);
   U15343 : NAND2_X1 port map( A1 => n11623, A2 => n2635, ZN => n5233);
   U15347 : XOR2_X1 port map( A1 => n15308, A2 => n24387, Z => n4419);
   U15351 : AND2_X1 port map( A1 => n25867, A2 => n25897, Z => n8780);
   U15354 : XOR2_X1 port map( A1 => Plaintext(189), A2 => Key(189), Z => n5594)
                           ;
   U15356 : INV_X1 port map( I => n23705, ZN => n4086);
   U15360 : OAI21_X1 port map( A1 => n25375, A2 => n30276, B => n4089, ZN => 
                           n25357);
   U15363 : XOR2_X1 port map( A1 => n11836, A2 => n11835, Z => n11834);
   U15365 : XOR2_X1 port map( A1 => n24593, A2 => n4091, Z => n5429);
   U15366 : XOR2_X1 port map( A1 => n24645, A2 => n28898, Z => n4091);
   U15375 : NAND2_X1 port map( A1 => n28825, A2 => n8846, ZN => n5814);
   U15379 : INV_X1 port map( I => n16596, ZN => n18779);
   U15395 : NAND2_X2 port map( A1 => n1337, A2 => n9678, ZN => n8041);
   U15396 : XOR2_X1 port map( A1 => n1227, A2 => n4112, Z => n15484);
   U15397 : XOR2_X1 port map( A1 => n27151, A2 => n25856, Z => n4112);
   U15407 : XOR2_X1 port map( A1 => n24424, A2 => n24425, Z => n6726);
   U15408 : XOR2_X1 port map( A1 => n24416, A2 => n24796, Z => n24425);
   U15410 : BUF_X2 port map( I => n8190, Z => n4119);
   U15420 : OAI21_X1 port map( A1 => n27619, A2 => n27336, B => n12028, ZN => 
                           n21549);
   U15436 : XOR2_X1 port map( A1 => n23441, A2 => n17871, Z => n4559);
   U15440 : INV_X2 port map( I => n4133, ZN => n20156);
   U15451 : INV_X1 port map( I => n6259, ZN => n12570);
   U15452 : NAND2_X1 port map( A1 => n12570, A2 => n25197, ZN => n4533);
   U15457 : XOR2_X1 port map( A1 => n7731, A2 => n30540, Z => n24629);
   U15461 : AOI22_X2 port map( A1 => n8461, A2 => n18422, B1 => n18616, B2 => 
                           n17224, ZN => n14811);
   U15478 : XOR2_X1 port map( A1 => n22799, A2 => n4154, Z => n14381);
   U15479 : XOR2_X1 port map( A1 => n13347, A2 => n15941, Z => n4154);
   U15485 : NOR2_X1 port map( A1 => n12930, A2 => n12931, ZN => n9502);
   U15486 : OAI21_X1 port map( A1 => n917, A2 => n916, B => n9898, ZN => n9897)
                           ;
   U15487 : NAND2_X1 port map( A1 => n9897, A2 => n9896, ZN => n9895);
   U15488 : OAI22_X2 port map( A1 => n18647, A2 => n5456, B1 => n10125, B2 => 
                           n17792, ZN => n5455);
   U15490 : XOR2_X1 port map( A1 => n11860, A2 => n11859, Z => n4158);
   U15491 : XNOR2_X1 port map( A1 => n22273, A2 => n21931, ZN => n6543);
   U15493 : INV_X1 port map( I => n10404, ZN => n4456);
   U15512 : NAND2_X1 port map( A1 => n15043, A2 => n15169, ZN => n20341);
   U15515 : INV_X1 port map( I => n18002, ZN => n4168);
   U15525 : NOR2_X1 port map( A1 => n8207, A2 => n25179, ZN => n8932);
   U15528 : NAND2_X2 port map( A1 => n21867, A2 => n13652, ZN => n21863);
   U15530 : INV_X1 port map( I => n20015, ZN => n4893);
   U15532 : XOR2_X1 port map( A1 => n8921, A2 => n19702, Z => n7184);
   U15533 : XOR2_X1 port map( A1 => n18911, A2 => n19743, Z => n19702);
   U15534 : XOR2_X1 port map( A1 => n14743, A2 => n14744, Z => n17821);
   U15536 : XOR2_X1 port map( A1 => n5702, A2 => n533, Z => n4173);
   U15539 : AOI21_X2 port map( A1 => n23818, A2 => n23819, B => n23817, ZN => 
                           n24327);
   U15547 : XOR2_X1 port map( A1 => n4176, A2 => n19512, Z => n16646);
   U15548 : XOR2_X1 port map( A1 => n12801, A2 => n12683, Z => n4176);
   U15553 : INV_X2 port map( I => n4180, ZN => n11958);
   U15554 : XNOR2_X1 port map( A1 => n17356, A2 => n17355, ZN => n4180);
   U15557 : XOR2_X1 port map( A1 => n6316, A2 => n10901, Z => n10900);
   U15559 : XOR2_X1 port map( A1 => n14833, A2 => n4187, Z => n4186);
   U15573 : XOR2_X1 port map( A1 => n8682, A2 => n4196, Z => n8681);
   U15574 : XOR2_X1 port map( A1 => n11783, A2 => n15936, Z => n4196);
   U15578 : NAND3_X2 port map( A1 => n24856, A2 => n7853, A3 => n7854, ZN => 
                           n25082);
   U15583 : INV_X2 port map( I => n4200, ZN => n18349);
   U15587 : XOR2_X1 port map( A1 => n20723, A2 => n20859, Z => n16803);
   U15590 : NAND2_X1 port map( A1 => n4447, A2 => n9181, ZN => n25814);
   U15604 : NAND2_X2 port map( A1 => n6010, A2 => n8667, ZN => n23111);
   U15609 : XOR2_X1 port map( A1 => n19594, A2 => n463, Z => n5138);
   U15613 : XNOR2_X1 port map( A1 => n23249, A2 => n23450, ZN => n5263);
   U15614 : INV_X2 port map( I => n4224, ZN => n4373);
   U15616 : XOR2_X1 port map( A1 => n21044, A2 => n27169, Z => n9607);
   U15619 : NOR2_X1 port map( A1 => n16440, A2 => n21338, ZN => n7115);
   U15633 : AOI21_X2 port map( A1 => n18084, A2 => n4232, B => n24364, ZN => 
                           n24910);
   U15636 : INV_X1 port map( I => n21146, ZN => n4865);
   U15639 : NAND2_X1 port map( A1 => n22645, A2 => n10724, ZN => n13973);
   U15641 : INV_X2 port map( I => n4243, ZN => n11045);
   U15645 : AOI21_X2 port map( A1 => n24301, A2 => n24302, B => n24306, ZN => 
                           n24645);
   U15649 : OR2_X1 port map( A1 => n18800, A2 => n8395, Z => n4255);
   U15650 : XOR2_X1 port map( A1 => n24281, A2 => n24280, Z => n11717);
   U15663 : NAND3_X1 port map( A1 => n7855, A2 => n16632, A3 => n15254, ZN => 
                           n7853);
   U15664 : AOI21_X1 port map( A1 => n5908, A2 => n12194, B => n1346, ZN => 
                           n4261);
   U15668 : XOR2_X1 port map( A1 => n20762, A2 => n26058, Z => n4263);
   U15678 : XOR2_X1 port map( A1 => n8488, A2 => n9993, Z => n9992);
   U15685 : XOR2_X1 port map( A1 => n23441, A2 => n23368, Z => n4273);
   U15687 : XOR2_X1 port map( A1 => n24416, A2 => n30540, Z => n12067);
   U15694 : OR2_X1 port map( A1 => n10335, A2 => n568, Z => n17060);
   U15696 : XOR2_X1 port map( A1 => n8214, A2 => n4280, Z => n9239);
   U15697 : XOR2_X1 port map( A1 => n24371, A2 => n9241, Z => n4280);
   U15704 : XOR2_X1 port map( A1 => n32860, A2 => n12491, Z => n11551);
   U15705 : XOR2_X1 port map( A1 => n24847, A2 => n10084, Z => n24541);
   U15712 : OR2_X1 port map( A1 => n20575, A2 => n20574, Z => n4290);
   U15721 : OAI21_X2 port map( A1 => n4370, A2 => n4368, B => n4367, ZN => 
                           n20627);
   U15722 : NAND2_X2 port map( A1 => n8332, A2 => n4299, ZN => n17408);
   U15725 : XOR2_X1 port map( A1 => Plaintext(102), A2 => Key(102), Z => n6634)
                           ;
   U15727 : OR2_X1 port map( A1 => n5753, A2 => n5327, Z => n5752);
   U15730 : AND2_X1 port map( A1 => n7161, A2 => n27021, Z => n7967);
   U15734 : AND2_X1 port map( A1 => n21621, A2 => n21620, Z => n4310);
   U15745 : XOR2_X1 port map( A1 => n24549, A2 => n9694, Z => n5231);
   U15747 : INV_X2 port map( I => n4330, ZN => n8420);
   U15749 : XOR2_X1 port map( A1 => n4332, A2 => n24646, Z => n6417);
   U15752 : NAND2_X1 port map( A1 => n8156, A2 => n7843, ZN => n25671);
   U15756 : OAI21_X2 port map( A1 => n5804, A2 => n26778, B => n4335, ZN => 
                           n17793);
   U15758 : XOR2_X1 port map( A1 => n4338, A2 => n23377, Z => n10936);
   U15759 : XOR2_X1 port map( A1 => n3723, A2 => n25040, Z => n7999);
   U15760 : XOR2_X1 port map( A1 => n32881, A2 => n3723, Z => n21900);
   U15769 : XOR2_X1 port map( A1 => n24764, A2 => n24620, Z => n4352);
   U15770 : XOR2_X1 port map( A1 => n5268, A2 => n13060, Z => n4353);
   U15771 : OAI21_X2 port map( A1 => n12985, A2 => n14913, B => n12983, ZN => 
                           n13060);
   U15772 : XOR2_X1 port map( A1 => n4355, A2 => n24354, Z => n4354);
   U15773 : XOR2_X1 port map( A1 => n5539, A2 => n1231, Z => n4355);
   U15777 : INV_X2 port map( I => n4362, ZN => n19630);
   U15778 : NAND2_X1 port map( A1 => n18876, A2 => n31948, ZN => n4365);
   U15788 : XOR2_X1 port map( A1 => n28823, A2 => n25224, Z => n15025);
   U15789 : XOR2_X1 port map( A1 => n28823, A2 => n21018, Z => n5068);
   U15793 : XOR2_X1 port map( A1 => n22043, A2 => n22266, Z => n4379);
   U15794 : XOR2_X1 port map( A1 => n12627, A2 => n22045, Z => n4380);
   U15797 : NOR2_X2 port map( A1 => n4387, A2 => n4386, ZN => n15028);
   U15804 : XOR2_X1 port map( A1 => n7363, A2 => n29299, Z => n7107);
   U15807 : XOR2_X1 port map( A1 => n19537, A2 => n4403, Z => n4401);
   U15809 : XOR2_X1 port map( A1 => n19597, A2 => n25001, Z => n4403);
   U15814 : XOR2_X1 port map( A1 => n4413, A2 => n4412, Z => n4411);
   U15815 : XOR2_X1 port map( A1 => n29235, A2 => n26000, Z => n4412);
   U15816 : XOR2_X1 port map( A1 => n23383, A2 => n23465, Z => n4414);
   U15826 : XOR2_X1 port map( A1 => n21993, A2 => n514, Z => n4427);
   U15832 : NAND3_X1 port map( A1 => n23031, A2 => n22945, A3 => n773, ZN => 
                           n7277);
   U15834 : INV_X2 port map( I => n16272, ZN => n22681);
   U15836 : XOR2_X1 port map( A1 => n22182, A2 => n22148, Z => n4437);
   U15840 : XOR2_X1 port map( A1 => n4446, A2 => n4444, Z => n17150);
   U15841 : XOR2_X1 port map( A1 => n4955, A2 => n4445, Z => n4444);
   U15842 : XOR2_X1 port map( A1 => n30321, A2 => n15147, Z => n4445);
   U15845 : MUX2_X1 port map( I0 => n25820, I1 => n25804, S => n4450, Z => 
                           n4447);
   U15847 : XOR2_X1 port map( A1 => n20907, A2 => n28864, Z => n4448);
   U15848 : INV_X2 port map( I => n4449, ZN => n4490);
   U15849 : INV_X2 port map( I => n4450, ZN => n25823);
   U15850 : XOR2_X1 port map( A1 => n3682, A2 => n24374, Z => n22081);
   U15851 : XOR2_X1 port map( A1 => n3682, A2 => n25126, Z => n21899);
   U15854 : XOR2_X1 port map( A1 => n12419, A2 => n3682, Z => n10815);
   U15868 : XOR2_X1 port map( A1 => n6156, A2 => n5964, Z => n4464);
   U15870 : XOR2_X1 port map( A1 => n4792, A2 => n4466, Z => n13932);
   U15875 : NOR2_X2 port map( A1 => n6672, A2 => n6377, ZN => n14564);
   U15877 : OAI21_X2 port map( A1 => n24338, A2 => n767, B => n2847, ZN => 
                           n24165);
   U15878 : NAND2_X2 port map( A1 => n16859, A2 => n33990, ZN => n24166);
   U15883 : NAND2_X1 port map( A1 => n15243, A2 => n31129, ZN => n4486);
   U15885 : INV_X2 port map( I => n31920, ZN => n25712);
   U15890 : OR2_X1 port map( A1 => n10858, A2 => n4770, Z => n9248);
   U15891 : OAI21_X2 port map( A1 => n5532, A2 => n9428, B => n9426, ZN => 
                           n10858);
   U15898 : XOR2_X1 port map( A1 => n4236, A2 => n1424, Z => n6376);
   U15903 : NAND2_X1 port map( A1 => n17767, A2 => n17971, ZN => n16266);
   U15909 : MUX2_X1 port map( I0 => n21536, I1 => n17274, S => n21569, Z => 
                           n21537);
   U15910 : NOR2_X1 port map( A1 => n3376, A2 => n4525, ZN => n14322);
   U15911 : NOR2_X1 port map( A1 => n5113, A2 => n4525, ZN => n17838);
   U15912 : OAI21_X1 port map( A1 => n9481, A2 => n4525, B => n4524, ZN => 
                           n9480);
   U15920 : XOR2_X1 port map( A1 => n28926, A2 => n1395, Z => n4530);
   U15921 : XOR2_X1 port map( A1 => n29918, A2 => n17723, Z => n17722);
   U15925 : OR2_X1 port map( A1 => n17662, A2 => n397, Z => n12077);
   U15928 : XOR2_X1 port map( A1 => n4557, A2 => n4556, Z => n4555);
   U15929 : XOR2_X1 port map( A1 => n26915, A2 => n16555, Z => n4556);
   U15930 : XOR2_X1 port map( A1 => n32899, A2 => n6905, Z => n4557);
   U15942 : XOR2_X1 port map( A1 => n13596, A2 => n4565, Z => n9164);
   U15943 : XOR2_X1 port map( A1 => n7173, A2 => n13595, Z => n4565);
   U15944 : XOR2_X1 port map( A1 => n5970, A2 => n24475, Z => n7173);
   U15946 : XOR2_X1 port map( A1 => n30314, A2 => n30329, Z => n5600);
   U15955 : XOR2_X1 port map( A1 => n26084, A2 => n5169, Z => n4579);
   U15959 : XOR2_X1 port map( A1 => n22153, A2 => n17187, Z => n4583);
   U15960 : NAND2_X1 port map( A1 => n20447, A2 => n31454, ZN => n4585);
   U15965 : XOR2_X1 port map( A1 => n6650, A2 => n22151, Z => n4590);
   U15966 : NAND2_X1 port map( A1 => n1271, A2 => n4599, ZN => n23015);
   U15967 : NAND2_X1 port map( A1 => n14540, A2 => n4599, ZN => n17399);
   U15969 : INV_X2 port map( I => n29061, ZN => n18891);
   U15970 : NOR2_X1 port map( A1 => n29061, A2 => n14926, ZN => n11410);
   U15971 : INV_X1 port map( I => Plaintext(16), ZN => n4601);
   U15978 : XOR2_X1 port map( A1 => n15183, A2 => n27126, Z => n4610);
   U15980 : OR2_X1 port map( A1 => n18266, A2 => n18265, Z => n4618);
   U15983 : XOR2_X1 port map( A1 => n14382, A2 => n14381, Z => n8523);
   U15984 : NOR2_X1 port map( A1 => n32127, A2 => n18643, ZN => n4624);
   U15986 : AOI21_X1 port map( A1 => n17266, A2 => n4626, B => n28238, ZN => 
                           n18378);
   U16000 : AOI21_X1 port map( A1 => n11893, A2 => n565, B => n16317, ZN => 
                           n4636);
   U16002 : AOI21_X1 port map( A1 => n7039, A2 => n4642, B => n7037, ZN => 
                           n10157);
   U16003 : XOR2_X1 port map( A1 => n2045, A2 => n25167, Z => n10163);
   U16011 : OAI21_X1 port map( A1 => n19301, A2 => n1052, B => n4658, ZN => 
                           n14736);
   U16012 : XOR2_X1 port map( A1 => n23182, A2 => n538, Z => n4660);
   U16014 : XOR2_X1 port map( A1 => n23138, A2 => n529, Z => n4662);
   U16015 : XOR2_X1 port map( A1 => n23267, A2 => n31727, Z => n23138);
   U16016 : INV_X1 port map( I => n31161, ZN => n4663);
   U16025 : XNOR2_X1 port map( A1 => Plaintext(182), A2 => Key(182), ZN => 
                           n4669);
   U16028 : XOR2_X1 port map( A1 => n32648, A2 => n16506, Z => n4671);
   U16035 : NAND2_X1 port map( A1 => n7802, A2 => n4834, ZN => n4678);
   U16039 : XOR2_X1 port map( A1 => n29918, A2 => n16525, Z => n4681);
   U16041 : AOI21_X1 port map( A1 => n25265, A2 => n25264, B => n4685, ZN => 
                           n25267);
   U16042 : OAI22_X1 port map( A1 => n1207, A2 => n4686, B1 => n12431, B2 => 
                           n25284, ZN => n4685);
   U16044 : OR2_X1 port map( A1 => n25285, A2 => n25277, Z => n4686);
   U16048 : AOI21_X1 port map( A1 => n20635, A2 => n4693, B => n26278, ZN => 
                           n20322);
   U16054 : NOR2_X1 port map( A1 => n21721, A2 => n3467, ZN => n4699);
   U16059 : XOR2_X1 port map( A1 => n4704, A2 => n16705, Z => n8718);
   U16060 : XOR2_X1 port map( A1 => n4704, A2 => n19570, Z => n11354);
   U16065 : NAND2_X2 port map( A1 => n18694, A2 => n18693, ZN => n10714);
   U16066 : NAND2_X1 port map( A1 => n7687, A2 => n11477, ZN => n4716);
   U16067 : NAND2_X2 port map( A1 => n15576, A2 => n15574, ZN => n11477);
   U16073 : XOR2_X1 port map( A1 => n8306, A2 => n16555, Z => n4720);
   U16080 : XOR2_X1 port map( A1 => n4727, A2 => n4724, Z => n10337);
   U16081 : XOR2_X1 port map( A1 => n4726, A2 => n4725, Z => n4724);
   U16082 : XOR2_X1 port map( A1 => n1923, A2 => n25669, Z => n4725);
   U16083 : XOR2_X1 port map( A1 => n20783, A2 => n20955, Z => n4726);
   U16088 : XOR2_X1 port map( A1 => n4783, A2 => n15707, Z => n17498);
   U16089 : XOR2_X1 port map( A1 => n4729, A2 => n13825, Z => n4783);
   U16091 : NAND3_X2 port map( A1 => n5130, A2 => n5129, A3 => n668, ZN => 
                           n14855);
   U16092 : NAND2_X2 port map( A1 => n10313, A2 => n9462, ZN => n5016);
   U16104 : XOR2_X1 port map( A1 => n22017, A2 => n22033, Z => n4739);
   U16106 : XOR2_X1 port map( A1 => n12376, A2 => n22108, Z => n22016);
   U16112 : NOR2_X1 port map( A1 => n8270, A2 => n9172, ZN => n4743);
   U16124 : XOR2_X1 port map( A1 => n20897, A2 => n11066, Z => n4759);
   U16125 : NOR2_X1 port map( A1 => n21604, A2 => n17098, ZN => n11081);
   U16126 : XOR2_X1 port map( A1 => n4763, A2 => n4762, Z => n4761);
   U16127 : XOR2_X1 port map( A1 => n10292, A2 => n25086, Z => n4762);
   U16128 : NOR2_X2 port map( A1 => n6266, A2 => n4765, ZN => n10953);
   U16129 : NAND3_X2 port map( A1 => n4772, A2 => n14546, A3 => n13933, ZN => 
                           n6857);
   U16132 : XOR2_X1 port map( A1 => Plaintext(15), A2 => Key(15), Z => n4808);
   U16133 : XOR2_X1 port map( A1 => n4783, A2 => n13824, Z => n10617);
   U16134 : XOR2_X1 port map( A1 => n15606, A2 => n25190, Z => n5031);
   U16135 : XOR2_X1 port map( A1 => n31597, A2 => n3977, Z => n22320);
   U16136 : XOR2_X1 port map( A1 => n3977, A2 => n4788, Z => n22002);
   U16137 : XOR2_X1 port map( A1 => n11750, A2 => n4789, Z => n11748);
   U16142 : XOR2_X1 port map( A1 => n23358, A2 => n25801, Z => n4794);
   U16149 : XOR2_X1 port map( A1 => n13970, A2 => n32310, Z => n10799);
   U16154 : XOR2_X1 port map( A1 => n27130, A2 => n30495, Z => n22111);
   U16159 : INV_X2 port map( I => n4808, ZN => n11390);
   U16160 : NAND2_X2 port map( A1 => n4811, A2 => n4809, ZN => n23056);
   U16163 : NAND2_X2 port map( A1 => n7253, A2 => n7252, ZN => n20899);
   U16165 : AOI21_X2 port map( A1 => n23952, A2 => n16281, B => n17664, ZN => 
                           n4821);
   U16174 : XOR2_X1 port map( A1 => n22264, A2 => n27120, Z => n15367);
   U16176 : XOR2_X1 port map( A1 => n22214, A2 => n16530, Z => n4831);
   U16181 : NAND2_X2 port map( A1 => n10693, A2 => n10694, ZN => n4835);
   U16183 : NOR2_X1 port map( A1 => n4835, A2 => n11444, ZN => n11263);
   U16186 : NOR2_X1 port map( A1 => n11085, A2 => n4835, ZN => n11688);
   U16191 : XOR2_X1 port map( A1 => n15674, A2 => n24267, Z => n4840);
   U16194 : NAND2_X2 port map( A1 => n24259, A2 => n17800, ZN => n6547);
   U16195 : XOR2_X1 port map( A1 => n4849, A2 => n598, Z => n11733);
   U16197 : NOR2_X1 port map( A1 => n29495, A2 => n4396, ZN => n11195);
   U16198 : NOR2_X1 port map( A1 => n22558, A2 => n22671, ZN => n4850);
   U16207 : XOR2_X1 port map( A1 => n21926, A2 => n8979, Z => n4861);
   U16208 : NAND2_X1 port map( A1 => n8079, A2 => n27543, ZN => n21790);
   U16209 : AOI21_X2 port map( A1 => n4865, A2 => n27842, B => n4863, ZN => 
                           n21789);
   U16211 : NAND2_X1 port map( A1 => n171, A2 => n4869, ZN => n18384);
   U16212 : NOR2_X1 port map( A1 => n18571, A2 => n4869, ZN => n18385);
   U16213 : OAI21_X1 port map( A1 => n1190, A2 => n4869, B => n29087, ZN => 
                           n5053);
   U16214 : XOR2_X1 port map( A1 => Plaintext(99), A2 => Key(99), Z => n18823);
   U16218 : XOR2_X1 port map( A1 => n19584, A2 => n8089, Z => n4884);
   U16219 : XOR2_X1 port map( A1 => n27733, A2 => n25911, Z => n14407);
   U16221 : XOR2_X1 port map( A1 => n27733, A2 => n24968, Z => n24404);
   U16222 : XOR2_X1 port map( A1 => n1604, A2 => n1394, Z => n17041);
   U16223 : XOR2_X1 port map( A1 => n10006, A2 => n27185, Z => n10005);
   U16224 : INV_X2 port map( I => n11888, ZN => n4891);
   U16225 : NAND2_X1 port map( A1 => n23919, A2 => n4892, ZN => n15095);
   U16226 : NAND2_X1 port map( A1 => n16620, A2 => n33221, ZN => n23349);
   U16234 : NAND3_X1 port map( A1 => n24903, A2 => n27248, A3 => n10099, ZN => 
                           n4899);
   U16235 : NAND2_X2 port map( A1 => n4903, A2 => n4900, ZN => n24915);
   U16236 : INV_X1 port map( I => n5763, ZN => n4903);
   U16242 : XOR2_X1 port map( A1 => n34047, A2 => n25319, Z => n4915);
   U16243 : XOR2_X1 port map( A1 => n18180, A2 => n20816, Z => n20956);
   U16247 : NAND2_X2 port map( A1 => n4919, A2 => n6501, ZN => n16023);
   U16248 : OR2_X1 port map( A1 => n1335, A2 => n11915, Z => n4922);
   U16263 : NAND2_X2 port map( A1 => n5534, A2 => n5533, ZN => n5128);
   U16266 : OR2_X1 port map( A1 => n13601, A2 => n30191, Z => n4960);
   U16269 : XOR2_X1 port map( A1 => n31229, A2 => n29121, Z => n17042);
   U16272 : NAND2_X1 port map( A1 => n3657, A2 => n32531, ZN => n4982);
   U16276 : NOR2_X1 port map( A1 => n19855, A2 => n3989, ZN => n5909);
   U16280 : MUX2_X1 port map( I0 => n5073, I1 => n20155, S => n9724, Z => 
                           n12322);
   U16284 : XOR2_X1 port map( A1 => n4992, A2 => n26076, Z => n11351);
   U16296 : XOR2_X1 port map( A1 => n5013, A2 => n5011, Z => n9757);
   U16297 : XOR2_X1 port map( A1 => n5012, A2 => n9758, Z => n5011);
   U16301 : XOR2_X1 port map( A1 => n24830, A2 => n11297, Z => n5021);
   U16304 : XNOR2_X1 port map( A1 => n5022, A2 => n5023, ZN => n5019);
   U16306 : NAND2_X2 port map( A1 => n5027, A2 => n5025, ZN => n20968);
   U16307 : XOR2_X1 port map( A1 => n20968, A2 => n16612, Z => n5431);
   U16308 : NOR2_X1 port map( A1 => n16789, A2 => n20096, ZN => n18041);
   U16309 : XOR2_X1 port map( A1 => n7375, A2 => n7374, Z => n10414);
   U16311 : XOR2_X1 port map( A1 => n22012, A2 => n13067, Z => n22168);
   U16314 : NAND2_X1 port map( A1 => n15601, A2 => n5035, ZN => n22959);
   U16316 : XOR2_X1 port map( A1 => n23261, A2 => n556, Z => n5038);
   U16322 : INV_X1 port map( I => n24132, ZN => n5066);
   U16324 : XOR2_X1 port map( A1 => n5070, A2 => n5069, Z => n11515);
   U16325 : XOR2_X1 port map( A1 => n20721, A2 => n5071, Z => n5069);
   U16326 : XOR2_X1 port map( A1 => n5772, A2 => n1067, Z => n5071);
   U16327 : INV_X2 port map( I => n7940, ZN => n7941);
   U16331 : INV_X2 port map( I => n5074, ZN => n9724);
   U16336 : XOR2_X1 port map( A1 => n2073, A2 => n16613, Z => n5081);
   U16337 : OAI22_X2 port map( A1 => n7438, A2 => n12532, B1 => n7437, B2 => 
                           n7436, ZN => n19426);
   U16343 : INV_X1 port map( I => n5089, ZN => n24656);
   U16344 : XOR2_X1 port map( A1 => n5090, A2 => n16402, Z => n9694);
   U16345 : XOR2_X1 port map( A1 => n5090, A2 => n16605, Z => n24379);
   U16347 : NAND2_X1 port map( A1 => n979, A2 => n5097, ZN => n6694);
   U16350 : XOR2_X1 port map( A1 => n28709, A2 => n22248, Z => n5099);
   U16353 : XOR2_X1 port map( A1 => n5106, A2 => n5104, Z => n22579);
   U16354 : XOR2_X1 port map( A1 => n5105, A2 => n13371, Z => n5104);
   U16357 : XOR2_X1 port map( A1 => n22296, A2 => n22147, Z => n5107);
   U16359 : XOR2_X1 port map( A1 => n22149, A2 => n16613, Z => n5109);
   U16368 : XOR2_X1 port map( A1 => n22004, A2 => n21658, Z => n5126);
   U16372 : XOR2_X1 port map( A1 => n5133, A2 => n20661, Z => n9980);
   U16374 : NOR2_X2 port map( A1 => n12181, A2 => n15317, ZN => n5380);
   U16381 : INV_X1 port map( I => n5140, ZN => n9800);
   U16385 : XOR2_X1 port map( A1 => n5146, A2 => n5147, Z => n5145);
   U16386 : XOR2_X1 port map( A1 => n16733, A2 => n29954, Z => n5147);
   U16388 : NAND2_X2 port map( A1 => n9314, A2 => n9317, ZN => n17430);
   U16389 : XOR2_X1 port map( A1 => n19551, A2 => n19465, Z => n5152);
   U16395 : XOR2_X1 port map( A1 => n23502, A2 => n7994, Z => n5159);
   U16409 : XOR2_X1 port map( A1 => n32255, A2 => n13438, Z => n13437);
   U16410 : XOR2_X1 port map( A1 => n32255, A2 => n25208, Z => n13453);
   U16411 : XOR2_X1 port map( A1 => n16429, A2 => n24907, Z => n5169);
   U16421 : XOR2_X1 port map( A1 => n30303, A2 => n20784, Z => n21011);
   U16422 : INV_X2 port map( I => n5188, ZN => n8443);
   U16433 : XOR2_X1 port map( A1 => n5197, A2 => n10004, Z => n16392);
   U16434 : XOR2_X1 port map( A1 => n7288, A2 => n21457, Z => n5197);
   U16440 : XOR2_X1 port map( A1 => n13198, A2 => n26103, Z => n5207);
   U16442 : XOR2_X1 port map( A1 => n5462, A2 => n25450, Z => n18902);
   U16443 : XOR2_X1 port map( A1 => n24785, A2 => n25832, Z => n24537);
   U16444 : XOR2_X1 port map( A1 => n24785, A2 => n16520, Z => n6053);
   U16446 : XOR2_X1 port map( A1 => n20899, A2 => n24937, Z => n5210);
   U16451 : XOR2_X1 port map( A1 => n23502, A2 => n23406, Z => n5215);
   U16454 : NAND2_X2 port map( A1 => n5218, A2 => n5216, ZN => n20885);
   U16457 : NOR2_X1 port map( A1 => n21801, A2 => n5228, ZN => n15639);
   U16460 : NAND2_X2 port map( A1 => n10811, A2 => n24119, ZN => n24573);
   U16461 : XNOR2_X1 port map( A1 => n10631, A2 => n5790, ZN => n10729);
   U16465 : XOR2_X1 port map( A1 => n5237, A2 => n1045, Z => n5236);
   U16466 : XOR2_X1 port map( A1 => n19772, A2 => n1065, Z => n5237);
   U16467 : NAND2_X1 port map( A1 => n17640, A2 => n5239, ZN => n9558);
   U16472 : XOR2_X1 port map( A1 => n5724, A2 => n9908, Z => n5240);
   U16475 : XOR2_X1 port map( A1 => n20873, A2 => n20872, Z => n20902);
   U16477 : XOR2_X1 port map( A1 => n5243, A2 => n25225, Z => Ciphertext(77));
   U16480 : XOR2_X1 port map( A1 => n5256, A2 => n5255, Z => n6552);
   U16481 : XOR2_X1 port map( A1 => n24415, A2 => n554, Z => n5255);
   U16487 : XOR2_X1 port map( A1 => Plaintext(140), A2 => Key(140), Z => n10664
                           );
   U16488 : INV_X1 port map( I => n5273, ZN => n5272);
   U16492 : XOR2_X1 port map( A1 => n23209, A2 => n16464, Z => n5277);
   U16495 : XOR2_X1 port map( A1 => n6156, A2 => n19707, Z => n5279);
   U16496 : XOR2_X1 port map( A1 => n14337, A2 => n11219, Z => n19707);
   U16497 : XOR2_X1 port map( A1 => n19709, A2 => n18082, Z => n5280);
   U16504 : MUX2_X1 port map( I0 => n16493, I1 => n20012, S => n13605, Z => 
                           n19880);
   U16507 : XOR2_X1 port map( A1 => n29885, A2 => n26915, Z => n15690);
   U16515 : XOR2_X1 port map( A1 => n12414, A2 => n1070, Z => n5297);
   U16516 : AOI22_X2 port map( A1 => n21748, A2 => n21750, B1 => n13815, B2 => 
                           n30346, ZN => n11458);
   U16518 : NOR2_X1 port map( A1 => n23081, A2 => n1577, ZN => n8126);
   U16519 : MUX2_X1 port map( I0 => n6985, I1 => n23082, S => n1577, Z => 
                           n23080);
   U16520 : NOR2_X1 port map( A1 => n12869, A2 => n1124, ZN => n5305);
   U16526 : XOR2_X1 port map( A1 => n5316, A2 => n29344, Z => n5315);
   U16531 : XOR2_X1 port map( A1 => n15527, A2 => n12998, Z => n5322);
   U16534 : NAND3_X1 port map( A1 => n25410, A2 => n752, A3 => n25405, ZN => 
                           n24702);
   U16536 : XOR2_X1 port map( A1 => n17548, A2 => Key(101), Z => n17558);
   U16541 : XOR2_X1 port map( A1 => n20710, A2 => n5337, Z => n5336);
   U16545 : XOR2_X1 port map( A1 => n5340, A2 => n5338, Z => n6143);
   U16546 : XOR2_X1 port map( A1 => n24568, A2 => n5339, Z => n5338);
   U16547 : XOR2_X1 port map( A1 => n12454, A2 => n24943, Z => n5339);
   U16550 : XOR2_X1 port map( A1 => n15114, A2 => n17871, Z => n12659);
   U16555 : XOR2_X1 port map( A1 => n4295, A2 => n25358, Z => n5352);
   U16570 : INV_X2 port map( I => n5361, ZN => n6855);
   U16571 : NAND2_X1 port map( A1 => n22462, A2 => n22343, ZN => n23011);
   U16580 : MUX2_X1 port map( I0 => n23902, I1 => n23629, S => n1254, Z => 
                           n23631);
   U16583 : INV_X2 port map( I => n11988, ZN => n7116);
   U16588 : INV_X2 port map( I => n5392, ZN => n11915);
   U16589 : XOR2_X1 port map( A1 => Plaintext(133), A2 => Key(133), Z => n14156
                           );
   U16590 : INV_X2 port map( I => n5401, ZN => n17967);
   U16599 : XOR2_X1 port map( A1 => n11762, A2 => n5422, Z => n5421);
   U16600 : XOR2_X1 port map( A1 => n14125, A2 => n25598, Z => n5422);
   U16603 : XOR2_X1 port map( A1 => n29318, A2 => n24750, Z => n5425);
   U16609 : NAND2_X1 port map( A1 => n886, A2 => n752, ZN => n24701);
   U16614 : INV_X2 port map( I => n5432, ZN => n24975);
   U16616 : XOR2_X1 port map( A1 => n19742, A2 => n5435, Z => n5434);
   U16617 : XOR2_X1 port map( A1 => n19466, A2 => n27995, Z => n5435);
   U16622 : XOR2_X1 port map( A1 => Key(136), A2 => Plaintext(136), Z => n16995
                           );
   U16625 : XOR2_X1 port map( A1 => n23402, A2 => n23226, Z => n5445);
   U16636 : XOR2_X1 port map( A1 => n15844, A2 => n19641, Z => n19467);
   U16641 : NAND2_X2 port map( A1 => n5460, A2 => n9352, ZN => n20554);
   U16642 : NAND2_X1 port map( A1 => n20169, A2 => n5460, ZN => n20172);
   U16643 : INV_X2 port map( I => n20521, ZN => n5460);
   U16644 : XOR2_X1 port map( A1 => n5472, A2 => n3929, Z => n9605);
   U16645 : XOR2_X1 port map( A1 => n5472, A2 => n16530, Z => n10424);
   U16646 : XOR2_X1 port map( A1 => Plaintext(98), A2 => Key(98), Z => n16450);
   U16649 : INV_X2 port map( I => n7348, ZN => n5476);
   U16651 : OAI21_X2 port map( A1 => n18824, A2 => n17735, B => n5478, ZN => 
                           n19128);
   U16653 : NOR2_X1 port map( A1 => n16093, A2 => n26600, ZN => n13957);
   U16654 : NOR2_X1 port map( A1 => n4656, A2 => n26600, ZN => n19084);
   U16656 : INV_X2 port map( I => n6854, ZN => n5480);
   U16657 : XOR2_X1 port map( A1 => n5483, A2 => n19481, Z => n19482);
   U16658 : XOR2_X1 port map( A1 => n7971, A2 => n5484, Z => n5483);
   U16668 : XOR2_X1 port map( A1 => n5513, A2 => n21650, Z => n5501);
   U16670 : XOR2_X1 port map( A1 => n859, A2 => n22099, Z => n5503);
   U16671 : INV_X2 port map( I => n5504, ZN => n15746);
   U16672 : AOI21_X2 port map( A1 => n23404, A2 => n5742, B => n5505, ZN => 
                           n11326);
   U16675 : XOR2_X1 port map( A1 => n26582, A2 => n27179, Z => n5508);
   U16680 : XOR2_X1 port map( A1 => n14289, A2 => n4057, Z => n5513);
   U16681 : XOR2_X1 port map( A1 => n27148, A2 => n5399, Z => n23386);
   U16682 : XOR2_X1 port map( A1 => n5518, A2 => n5515, Z => n21168);
   U16683 : XOR2_X1 port map( A1 => n5517, A2 => n5516, Z => n5515);
   U16684 : XOR2_X1 port map( A1 => n20860, A2 => n16502, Z => n5516);
   U16685 : XOR2_X1 port map( A1 => n17554, A2 => n21016, Z => n5517);
   U16693 : XOR2_X1 port map( A1 => n31508, A2 => n24748, Z => n5522);
   U16696 : XOR2_X1 port map( A1 => n6156, A2 => n19343, Z => n5526);
   U16697 : INV_X2 port map( I => n5527, ZN => n23765);
   U16701 : NOR2_X1 port map( A1 => n33714, A2 => n820, ZN => n5582);
   U16709 : AOI21_X1 port map( A1 => n17725, A2 => n19063, B => n1053, ZN => 
                           n7186);
   U16711 : NOR3_X1 port map( A1 => n21560, A2 => n14236, A3 => n5546, ZN => 
                           n15319);
   U16713 : NOR2_X1 port map( A1 => n3657, A2 => n850, ZN => n6696);
   U16714 : INV_X1 port map( I => n21636, ZN => n21638);
   U16715 : NOR2_X2 port map( A1 => n9186, A2 => n780, ZN => n5575);
   U16720 : XOR2_X1 port map( A1 => n19564, A2 => n456, Z => n5562);
   U16723 : NAND2_X1 port map( A1 => n5575, A2 => n21453, ZN => n20436);
   U16724 : AOI21_X1 port map( A1 => n25217, A2 => n5043, B => n5577, ZN => 
                           n25219);
   U16732 : INV_X2 port map( I => n22535, ZN => n22537);
   U16739 : OAI21_X2 port map( A1 => n31923, A2 => n12610, B => n5602, ZN => 
                           n19556);
   U16742 : NOR2_X2 port map( A1 => n17556, A2 => n12744, ZN => n19424);
   U16744 : XOR2_X1 port map( A1 => n9955, A2 => n16824, Z => n5609);
   U16751 : OAI21_X2 port map( A1 => n5656, A2 => n5655, B => n4643, ZN => 
                           n15073);
   U16756 : XOR2_X1 port map( A1 => n16708, A2 => n25355, Z => n5629);
   U16760 : NAND2_X2 port map( A1 => n18986, A2 => n5637, ZN => n19589);
   U16770 : XNOR2_X1 port map( A1 => n22144, A2 => n21920, ZN => n5658);
   U16771 : XOR2_X1 port map( A1 => n21726, A2 => n22100, Z => n21920);
   U16775 : XOR2_X1 port map( A1 => n9848, A2 => n5666, Z => n5663);
   U16779 : XOR2_X1 port map( A1 => n24532, A2 => n16301, Z => n5666);
   U16788 : INV_X2 port map( I => n5675, ZN => n16625);
   U16790 : NOR2_X1 port map( A1 => n5677, A2 => n18493, ZN => n18424);
   U16791 : NOR2_X1 port map( A1 => n18326, A2 => n5677, ZN => n5676);
   U16792 : NAND2_X2 port map( A1 => n5682, A2 => n8786, ZN => n23485);
   U16795 : NAND4_X2 port map( A1 => n11725, A2 => n11724, A3 => n15781, A4 => 
                           n5690, ZN => n11722);
   U16797 : XOR2_X1 port map( A1 => n5692, A2 => n5691, Z => n17812);
   U16798 : XOR2_X1 port map( A1 => n23249, A2 => n23251, Z => n5691);
   U16804 : OAI22_X1 port map( A1 => n32868, A2 => n803, B1 => n724, B2 => 
                           n3163, ZN => n22693);
   U16805 : XOR2_X1 port map( A1 => n5699, A2 => n5697, Z => n15009);
   U16806 : XOR2_X1 port map( A1 => n5698, A2 => n14415, Z => n5697);
   U16807 : XOR2_X1 port map( A1 => n4400, A2 => n25098, Z => n5698);
   U16813 : XOR2_X1 port map( A1 => n34056, A2 => n23224, Z => n5702);
   U16818 : NOR2_X1 port map( A1 => n5707, A2 => n31017, ZN => n13649);
   U16822 : NAND2_X1 port map( A1 => n7334, A2 => n5713, ZN => n25083);
   U16823 : NAND2_X1 port map( A1 => n5713, A2 => n25106, ZN => n5712);
   U16827 : XOR2_X1 port map( A1 => n546, A2 => n24817, Z => n5714);
   U16832 : XOR2_X1 port map( A1 => n511, A2 => n13901, Z => n5722);
   U16834 : INV_X2 port map( I => n6894, ZN => n16668);
   U16837 : XOR2_X1 port map( A1 => n26084, A2 => n18011, Z => n5726);
   U16842 : XOR2_X1 port map( A1 => n20977, A2 => n5733, Z => n5732);
   U16843 : XOR2_X1 port map( A1 => n16708, A2 => n16381, Z => n5733);
   U16851 : NOR2_X1 port map( A1 => n978, A2 => n28222, ZN => n5745);
   U16853 : NAND2_X2 port map( A1 => n7538, A2 => n5754, ZN => n14147);
   U16855 : XOR2_X1 port map( A1 => n22021, A2 => n21886, Z => n21903);
   U16857 : XOR2_X1 port map( A1 => n30069, A2 => n31308, Z => n10923);
   U16859 : NAND2_X1 port map( A1 => n1384, A2 => n5760, ZN => n7434);
   U16862 : XOR2_X1 port map( A1 => n24643, A2 => n30104, Z => n24376);
   U16866 : XOR2_X1 port map( A1 => n7135, A2 => n7606, Z => n5767);
   U16868 : NAND2_X1 port map( A1 => n16205, A2 => n1122, ZN => n5771);
   U16869 : NAND3_X1 port map( A1 => n30328, A2 => n24922, A3 => n15569, ZN => 
                           n5774);
   U16870 : MUX2_X1 port map( I0 => n32571, I1 => n1211, S => n33585, Z => 
                           n25786);
   U16872 : XOR2_X1 port map( A1 => n5775, A2 => n6324, Z => n15994);
   U16879 : INV_X1 port map( I => n5792, ZN => n5791);
   U16883 : XOR2_X1 port map( A1 => n8232, A2 => n17793, Z => n13899);
   U16884 : NAND2_X1 port map( A1 => n5805, A2 => n28987, ZN => n5890);
   U16893 : NOR2_X2 port map( A1 => n7464, A2 => n21929, ZN => n7463);
   U16896 : XOR2_X1 port map( A1 => n24785, A2 => n1421, Z => n13793);
   U16899 : XOR2_X1 port map( A1 => n22085, A2 => n22096, Z => n21921);
   U16903 : XOR2_X1 port map( A1 => n5838, A2 => n1194, Z => Ciphertext(151));
   U16905 : NAND3_X1 port map( A1 => n30346, A2 => n13816, A3 => n21840, ZN => 
                           n14739);
   U16906 : NAND2_X1 port map( A1 => n16987, A2 => n5843, ZN => n21685);
   U16907 : NAND2_X1 port map( A1 => n16386, A2 => n30346, ZN => n21841);
   U16909 : XOR2_X1 port map( A1 => n5844, A2 => n11766, Z => n11765);
   U16912 : XOR2_X1 port map( A1 => n23474, A2 => n16597, Z => n5846);
   U16915 : AOI21_X1 port map( A1 => n18492, A2 => n17813, B => n17316, ZN => 
                           n5852);
   U16922 : NAND2_X1 port map( A1 => n6493, A2 => n780, ZN => n9273);
   U16923 : NAND2_X1 port map( A1 => n17437, A2 => n1337, ZN => n5857);
   U16924 : XOR2_X1 port map( A1 => n5862, A2 => n5859, Z => n5870);
   U16925 : XOR2_X1 port map( A1 => n5861, A2 => n5860, Z => n5859);
   U16926 : XOR2_X1 port map( A1 => n14588, A2 => n16655, Z => n5860);
   U16933 : INV_X1 port map( I => n22336, ZN => n22413);
   U16944 : INV_X2 port map( I => n5870, ZN => n16154);
   U16946 : XOR2_X1 port map( A1 => n9160, A2 => n16734, Z => n15077);
   U16947 : XOR2_X1 port map( A1 => n23324, A2 => n12200, Z => n5881);
   U16948 : INV_X1 port map( I => n23213, ZN => n5882);
   U16950 : XOR2_X1 port map( A1 => n21911, A2 => n6183, Z => n5885);
   U16952 : NAND2_X1 port map( A1 => n18274, A2 => n27129, ZN => n5891);
   U16960 : XOR2_X1 port map( A1 => n5904, A2 => n26701, Z => n14036);
   U16963 : NOR2_X1 port map( A1 => n6899, A2 => n17947, ZN => n5911);
   U16966 : XOR2_X1 port map( A1 => n5916, A2 => n1069, Z => Ciphertext(127));
   U16968 : XOR2_X1 port map( A1 => n19649, A2 => n16506, Z => n5919);
   U16970 : XOR2_X1 port map( A1 => n19721, A2 => n5921, Z => n5920);
   U16981 : NAND3_X2 port map( A1 => n19904, A2 => n19905, A3 => n5931, ZN => 
                           n20561);
   U16983 : XOR2_X1 port map( A1 => n5940, A2 => n23535, Z => n5939);
   U16984 : XOR2_X1 port map( A1 => n23534, A2 => n16634, Z => n5940);
   U16985 : XOR2_X1 port map( A1 => n7933, A2 => n5941, Z => n8167);
   U16986 : XOR2_X1 port map( A1 => n22293, A2 => n610, Z => n5941);
   U16989 : NAND2_X1 port map( A1 => n19033, A2 => n5946, ZN => n5945);
   U16990 : NAND2_X1 port map( A1 => n21404, A2 => n596, ZN => n5948);
   U16992 : INV_X2 port map( I => n5962, ZN => n10871);
   U16994 : NAND2_X1 port map( A1 => n2858, A2 => n5991, ZN => n5963);
   U16995 : INV_X2 port map( I => n19230, ZN => n19783);
   U16996 : XOR2_X1 port map( A1 => n19230, A2 => n1406, Z => n5964);
   U16997 : INV_X2 port map( I => n5965, ZN => n17240);
   U16998 : NAND2_X1 port map( A1 => n885, A2 => n25012, ZN => n24477);
   U17003 : XOR2_X1 port map( A1 => n22130, A2 => n22192, Z => n22293);
   U17008 : NAND2_X2 port map( A1 => n13707, A2 => n13708, ZN => n19384);
   U17010 : INV_X2 port map( I => n9203, ZN => n11912);
   U17013 : OAI21_X1 port map( A1 => n15456, A2 => n5981, B => n15457, ZN => 
                           n5983);
   U17016 : XOR2_X1 port map( A1 => n11332, A2 => n24442, Z => n24795);
   U17018 : NAND2_X1 port map( A1 => n22606, A2 => n5991, ZN => n6186);
   U17019 : NAND2_X1 port map( A1 => n4066, A2 => n19156, ZN => n15120);
   U17020 : NOR2_X1 port map( A1 => n18426, A2 => n4066, ZN => n18979);
   U17021 : XOR2_X1 port map( A1 => n3799, A2 => n25801, Z => n20647);
   U17022 : XOR2_X1 port map( A1 => n5994, A2 => n22005, Z => n21916);
   U17024 : XOR2_X1 port map( A1 => n28082, A2 => n31308, Z => n8755);
   U17027 : NAND2_X1 port map( A1 => n6003, A2 => n30146, ZN => n12692);
   U17031 : XOR2_X1 port map( A1 => n6008, A2 => n6005, Z => n24459);
   U17032 : XOR2_X1 port map( A1 => n6007, A2 => n6006, Z => n6005);
   U17033 : XOR2_X1 port map( A1 => n24526, A2 => n25722, Z => n6006);
   U17034 : XOR2_X1 port map( A1 => n24799, A2 => n24809, Z => n6007);
   U17039 : NAND2_X2 port map( A1 => n6322, A2 => n7648, ZN => n23109);
   U17044 : XOR2_X1 port map( A1 => n22130, A2 => n25545, Z => n6018);
   U17046 : XOR2_X1 port map( A1 => n13020, A2 => n22049, Z => n6020);
   U17048 : INV_X1 port map( I => n6673, ZN => n10011);
   U17054 : XOR2_X1 port map( A1 => n24478, A2 => n25206, Z => n12032);
   U17057 : XOR2_X1 port map( A1 => n19763, A2 => n19649, Z => n6028);
   U17058 : OAI21_X2 port map( A1 => n6030, A2 => n6029, B => n9134, ZN => 
                           n19763);
   U17059 : XOR2_X1 port map( A1 => n6033, A2 => n6032, Z => n6031);
   U17060 : XOR2_X1 port map( A1 => n19764, A2 => n25783, Z => n6032);
   U17066 : XOR2_X1 port map( A1 => n31229, A2 => n24833, Z => n14217);
   U17067 : XOR2_X1 port map( A1 => n7046, A2 => n25728, Z => n7994);
   U17068 : XOR2_X1 port map( A1 => n7046, A2 => n15409, Z => n15408);
   U17075 : XOR2_X1 port map( A1 => n13471, A2 => n6053, Z => n6052);
   U17080 : XOR2_X1 port map( A1 => n22213, A2 => n6056, Z => n6055);
   U17081 : XOR2_X1 port map( A1 => n15825, A2 => n16527, Z => n6056);
   U17089 : XOR2_X1 port map( A1 => n26683, A2 => n27101, Z => n16824);
   U17090 : XOR2_X1 port map( A1 => n26683, A2 => n16671, Z => n7875);
   U17091 : XOR2_X1 port map( A1 => n26683, A2 => n25506, Z => n14315);
   U17092 : XOR2_X1 port map( A1 => n26530, A2 => n20747, Z => n6078);
   U17101 : XOR2_X1 port map( A1 => n6088, A2 => n6087, Z => n6086);
   U17102 : XOR2_X1 port map( A1 => n20825, A2 => n25880, Z => n6087);
   U17103 : XOR2_X1 port map( A1 => n23181, A2 => n10218, Z => n10219);
   U17112 : XOR2_X1 port map( A1 => n6095, A2 => n25466, Z => Ciphertext(111));
   U17114 : MUX2_X1 port map( I0 => n25462, I1 => n25473, S => n6310, Z => 
                           n6097);
   U17115 : AOI21_X2 port map( A1 => n13249, A2 => n16490, B => n9738, ZN => 
                           n23051);
   U17116 : XOR2_X1 port map( A1 => n6103, A2 => n24643, Z => n9943);
   U17119 : NAND3_X1 port map( A1 => n9625, A2 => n33597, A3 => n5308, ZN => 
                           n6104);
   U17122 : XOR2_X1 port map( A1 => n19385, A2 => n6115, Z => n19387);
   U17127 : XOR2_X1 port map( A1 => n2896, A2 => n13579, Z => n6318);
   U17132 : XOR2_X1 port map( A1 => n27922, A2 => n1192, Z => n6127);
   U17134 : NAND2_X1 port map( A1 => n14652, A2 => n6138, ZN => n13686);
   U17137 : XOR2_X1 port map( A1 => n16897, A2 => n22242, Z => n9790);
   U17141 : NOR2_X1 port map( A1 => n22963, A2 => n6149, ZN => n6150);
   U17144 : XOR2_X1 port map( A1 => n23449, A2 => n23288, Z => n6151);
   U17147 : NAND2_X1 port map( A1 => n8304, A2 => n24908, ZN => n6155);
   U17148 : XOR2_X1 port map( A1 => n6159, A2 => n6160, Z => n13304);
   U17152 : NAND2_X2 port map( A1 => n7255, A2 => n7254, ZN => n20954);
   U17153 : INV_X2 port map( I => n9627, ZN => n9706);
   U17154 : XOR2_X1 port map( A1 => n20833, A2 => n6161, Z => n6160);
   U17155 : XOR2_X1 port map( A1 => n9627, A2 => n6162, Z => n6161);
   U17156 : INV_X1 port map( I => n25324, ZN => n6162);
   U17157 : XNOR2_X1 port map( A1 => n17517, A2 => n6906, ZN => n20833);
   U17162 : XOR2_X1 port map( A1 => n11206, A2 => n16597, Z => n6183);
   U17163 : XOR2_X1 port map( A1 => n9809, A2 => n27837, Z => n22042);
   U17165 : XOR2_X1 port map( A1 => n24809, A2 => n25465, Z => n6185);
   U17167 : NAND2_X1 port map( A1 => n21256, A2 => n6192, ZN => n21261);
   U17170 : OAI21_X1 port map( A1 => n18979, A2 => n18425, B => n18978, ZN => 
                           n6193);
   U17172 : NOR2_X1 port map( A1 => n14810, A2 => n6402, ZN => n9227);
   U17173 : AND2_X1 port map( A1 => n25312, A2 => n694, Z => n17709);
   U17175 : NOR2_X1 port map( A1 => n24121, A2 => n1775, ZN => n13748);
   U17176 : NAND2_X1 port map( A1 => n8932, A2 => n16273, ZN => n8340);
   U17179 : XOR2_X1 port map( A1 => Plaintext(22), A2 => Key(22), Z => n8317);
   U17192 : OR2_X1 port map( A1 => n19967, A2 => n14576, Z => n20022);
   U17193 : XOR2_X1 port map( A1 => n20669, A2 => n20667, Z => n6205);
   U17196 : AND2_X1 port map( A1 => n15528, A2 => n16528, Z => n15530);
   U17197 : XOR2_X1 port map( A1 => n18903, A2 => n6209, Z => n6281);
   U17200 : XOR2_X1 port map( A1 => n24768, A2 => n6211, Z => n7042);
   U17201 : XOR2_X1 port map( A1 => n13060, A2 => n16561, Z => n6211);
   U17204 : NAND2_X1 port map( A1 => n24084, A2 => n24087, ZN => n14912);
   U17207 : OAI21_X2 port map( A1 => n11788, A2 => n10119, B => n10116, ZN => 
                           n24819);
   U17213 : XOR2_X1 port map( A1 => Plaintext(60), A2 => Key(60), Z => n6215);
   U17228 : XOR2_X1 port map( A1 => n31450, A2 => n11889, Z => n6229);
   U17229 : NAND3_X1 port map( A1 => n11517, A2 => n12197, A3 => n12196, ZN => 
                           n10694);
   U17237 : XNOR2_X1 port map( A1 => n24537, A2 => n24835, ZN => n6341);
   U17243 : XOR2_X1 port map( A1 => n22044, A2 => n9129, Z => n6245);
   U17245 : XNOR2_X1 port map( A1 => n19620, A2 => n15621, ZN => n6867);
   U17246 : CLKBUF_X2 port map( I => Key(29), Z => n24861);
   U17251 : NAND2_X2 port map( A1 => n6252, A2 => n16763, ZN => n19348);
   U17253 : XOR2_X1 port map( A1 => n10902, A2 => n19721, Z => n6254);
   U17254 : NAND2_X1 port map( A1 => n22156, A2 => n17151, ZN => n22665);
   U17264 : XOR2_X1 port map( A1 => Plaintext(158), A2 => Key(158), Z => n6265)
                           ;
   U17268 : XOR2_X1 port map( A1 => n24654, A2 => n1226, Z => n6267);
   U17269 : XOR2_X1 port map( A1 => n21912, A2 => n6318, Z => n6811);
   U17271 : NAND3_X2 port map( A1 => n6268, A2 => n9542, A3 => n11534, ZN => 
                           n10146);
   U17277 : XOR2_X1 port map( A1 => n20957, A2 => n474, Z => n6273);
   U17279 : AND2_X1 port map( A1 => n25628, A2 => n4146, Z => n16096);
   U17286 : NOR2_X2 port map( A1 => n8064, A2 => n8063, ZN => n24177);
   U17289 : INV_X1 port map( I => n16828, ZN => n16827);
   U17297 : NOR2_X2 port map( A1 => n13295, A2 => n34107, ZN => n19356);
   U17298 : AND2_X1 port map( A1 => n9692, A2 => n20576, Z => n8144);
   U17299 : OR2_X1 port map( A1 => n12042, A2 => n32875, Z => n7974);
   U17300 : INV_X2 port map( I => n6281, ZN => n11913);
   U17303 : OAI21_X2 port map( A1 => n4245, A2 => n6283, B => n24893, ZN => 
                           n14954);
   U17306 : XOR2_X1 port map( A1 => n14239, A2 => n8575, Z => n14238);
   U17309 : XNOR2_X1 port map( A1 => n12785, A2 => n13553, ZN => n22256);
   U17313 : XOR2_X1 port map( A1 => n24823, A2 => n24548, Z => n18042);
   U17314 : NAND3_X2 port map( A1 => n11830, A2 => n16950, A3 => n29292, ZN => 
                           n24823);
   U17323 : XOR2_X1 port map( A1 => n10869, A2 => n24574, Z => n8747);
   U17334 : NOR2_X1 port map( A1 => n15302, A2 => n21530, ZN => n12095);
   U17341 : XOR2_X1 port map( A1 => n18315, A2 => Key(130), Z => n16462);
   U17347 : XOR2_X1 port map( A1 => n20977, A2 => n14522, Z => n9635);
   U17353 : XOR2_X1 port map( A1 => n10277, A2 => n10276, Z => n9301);
   U17354 : XOR2_X1 port map( A1 => n12971, A2 => n543, Z => n6316);
   U17362 : NAND2_X1 port map( A1 => n14258, A2 => n14257, ZN => n10783);
   U17367 : XOR2_X1 port map( A1 => n14428, A2 => n20871, Z => n6324);
   U17372 : XOR2_X1 port map( A1 => n17004, A2 => n22091, Z => n6327);
   U17373 : XOR2_X1 port map( A1 => n10813, A2 => n10816, Z => n14514);
   U17376 : XNOR2_X1 port map( A1 => n24814, A2 => n11537, ZN => n8537);
   U17387 : XOR2_X1 port map( A1 => n13163, A2 => n6341, Z => n7080);
   U17392 : XOR2_X1 port map( A1 => n15743, A2 => n17938, Z => n15754);
   U17394 : NOR2_X1 port map( A1 => n16534, A2 => n10937, ZN => n11067);
   U17398 : NAND2_X1 port map( A1 => n30308, A2 => n25345, ZN => n6345);
   U17399 : INV_X2 port map( I => n6346, ZN => n7216);
   U17400 : XOR2_X1 port map( A1 => Plaintext(104), A2 => Key(104), Z => n6346)
                           ;
   U17403 : XOR2_X1 port map( A1 => n18109, A2 => n11604, Z => n19690);
   U17410 : XNOR2_X1 port map( A1 => n23200, A2 => n16527, ZN => n9228);
   U17417 : XOR2_X1 port map( A1 => n16080, A2 => n19673, Z => n6721);
   U17421 : NAND2_X2 port map( A1 => n12547, A2 => n12546, ZN => n23540);
   U17424 : NOR2_X1 port map( A1 => n23067, A2 => n29070, ZN => n6677);
   U17426 : XOR2_X1 port map( A1 => n23152, A2 => n23240, Z => n22518);
   U17427 : XOR2_X1 port map( A1 => n20757, A2 => n15025, Z => n7908);
   U17433 : XOR2_X1 port map( A1 => n7452, A2 => n600, Z => n7234);
   U17434 : XOR2_X1 port map( A1 => n33380, A2 => n13638, Z => n9131);
   U17447 : NAND2_X1 port map( A1 => n7897, A2 => n13318, ZN => n6710);
   U17449 : INV_X1 port map( I => n8951, ZN => n8950);
   U17452 : XNOR2_X1 port map( A1 => n19468, A2 => n19394, ZN => n8401);
   U17455 : XOR2_X1 port map( A1 => n24116, A2 => n24375, Z => n6397);
   U17459 : NAND2_X2 port map( A1 => n1356, A2 => n7577, ZN => n20604);
   U17460 : XOR2_X1 port map( A1 => n19731, A2 => n19732, Z => n10576);
   U17463 : NAND2_X1 port map( A1 => n2471, A2 => n10310, ZN => n22806);
   U17465 : XOR2_X1 port map( A1 => n20887, A2 => n10557, Z => n7126);
   U17468 : XOR2_X1 port map( A1 => n28983, A2 => n26530, Z => n7565);
   U17470 : OR2_X1 port map( A1 => n19899, A2 => n17688, Z => n20106);
   U17489 : AND2_X1 port map( A1 => n1786, A2 => n11987, Z => n7656);
   U17491 : INV_X1 port map( I => n25020, ZN => n9052);
   U17493 : NOR2_X1 port map( A1 => n884, A2 => n14832, ZN => n6425);
   U17498 : OR2_X1 port map( A1 => n20755, A2 => n6431, Z => n7952);
   U17501 : INV_X2 port map( I => n6434, ZN => n17306);
   U17509 : INV_X1 port map( I => n15581, ZN => n15195);
   U17510 : OR2_X1 port map( A1 => n15581, A2 => n22487, Z => n11245);
   U17513 : XOR2_X1 port map( A1 => n7772, A2 => n1404, Z => n17546);
   U17516 : XOR2_X1 port map( A1 => n5381, A2 => n31491, Z => n6445);
   U17519 : XOR2_X1 port map( A1 => Plaintext(19), A2 => Key(19), Z => n7712);
   U17526 : XOR2_X1 port map( A1 => n16717, A2 => n16718, Z => n6452);
   U17527 : OR2_X1 port map( A1 => n10435, A2 => n579, Z => n7525);
   U17531 : XOR2_X1 port map( A1 => n22132, A2 => n31105, Z => n22134);
   U17535 : OR2_X1 port map( A1 => n21374, A2 => n4145, Z => n12110);
   U17547 : XOR2_X1 port map( A1 => n16949, A2 => n6465, Z => n6464);
   U17549 : INV_X2 port map( I => n15721, ZN => n16568);
   U17551 : XOR2_X1 port map( A1 => n24474, A2 => n24421, Z => n24373);
   U17552 : XOR2_X1 port map( A1 => n17682, A2 => n458, Z => n24678);
   U17554 : XOR2_X1 port map( A1 => n6469, A2 => n1410, Z => Ciphertext(144));
   U17556 : NAND3_X1 port map( A1 => n28767, A2 => n16154, A3 => n29840, ZN => 
                           n18147);
   U17563 : OR2_X1 port map( A1 => n11255, A2 => n24327, Z => n7099);
   U17569 : NOR2_X1 port map( A1 => n12937, A2 => n18842, ZN => n10451);
   U17570 : OAI21_X1 port map( A1 => n24432, A2 => n27164, B => n6477, ZN => 
                           n24433);
   U17571 : NAND2_X1 port map( A1 => n24431, A2 => n27164, ZN => n6477);
   U17572 : NAND2_X1 port map( A1 => n22588, A2 => n16562, ZN => n22590);
   U17573 : XOR2_X1 port map( A1 => n22173, A2 => n28490, Z => n22175);
   U17576 : XOR2_X1 port map( A1 => n1345, A2 => n13970, Z => n7030);
   U17579 : XOR2_X1 port map( A1 => n17549, A2 => n9764, Z => n6485);
   U17584 : OR2_X1 port map( A1 => n13059, A2 => n16916, Z => n16788);
   U17596 : NOR2_X1 port map( A1 => n18609, A2 => n18485, ZN => n18276);
   U17598 : XOR2_X1 port map( A1 => n6720, A2 => n6885, Z => n6719);
   U17605 : NOR2_X2 port map( A1 => n6504, A2 => n10128, ZN => n17820);
   U17606 : XOR2_X1 port map( A1 => n6507, A2 => n348, Z => n8485);
   U17609 : NOR2_X2 port map( A1 => n18502, A2 => n18503, ZN => n19089);
   U17612 : XOR2_X1 port map( A1 => n24389, A2 => n24600, Z => n6513);
   U17613 : XOR2_X1 port map( A1 => n21965, A2 => n6515, Z => n15229);
   U17617 : XOR2_X1 port map( A1 => n23258, A2 => n23476, Z => n23520);
   U17622 : AND2_X1 port map( A1 => n24063, A2 => n9946, Z => n9945);
   U17629 : XOR2_X1 port map( A1 => n21037, A2 => n20389, Z => n20390);
   U17633 : AOI21_X1 port map( A1 => n25742, A2 => n25741, B => n6524, ZN => 
                           n10082);
   U17637 : AND2_X1 port map( A1 => n33078, A2 => n13200, Z => n8662);
   U17640 : OR2_X1 port map( A1 => n21666, A2 => n28618, Z => n11584);
   U17643 : XOR2_X1 port map( A1 => n6526, A2 => n16454, Z => Ciphertext(184));
   U17653 : XOR2_X1 port map( A1 => n19574, A2 => n10866, Z => n10865);
   U17663 : NAND3_X2 port map( A1 => n22356, A2 => n22511, A3 => n13078, ZN => 
                           n22357);
   U17669 : XOR2_X1 port map( A1 => n24796, A2 => n16525, Z => n14689);
   U17675 : NAND3_X1 port map( A1 => n9148, A2 => n32186, A3 => n31862, ZN => 
                           n9147);
   U17676 : XOR2_X1 port map( A1 => n2142, A2 => n12580, Z => n12579);
   U17683 : XOR2_X1 port map( A1 => n31277, A2 => n14206, Z => n6561);
   U17684 : XOR2_X1 port map( A1 => n20863, A2 => n508, Z => n6562);
   U17687 : OR2_X1 port map( A1 => n18931, A2 => n17725, Z => n6567);
   U17688 : XOR2_X1 port map( A1 => n9018, A2 => n11586, Z => n6572);
   U17690 : XOR2_X1 port map( A1 => n7861, A2 => n7860, Z => n6574);
   U17691 : OAI21_X1 port map( A1 => n12175, A2 => n6579, B => n13254, ZN => 
                           n7027);
   U17692 : XOR2_X1 port map( A1 => Plaintext(51), A2 => Key(51), Z => n6776);
   U17701 : XOR2_X1 port map( A1 => n14401, A2 => n6601, Z => n20049);
   U17702 : XOR2_X1 port map( A1 => n28822, A2 => n20836, Z => n6601);
   U17703 : XOR2_X1 port map( A1 => n14132, A2 => n2616, Z => n14401);
   U17704 : XOR2_X1 port map( A1 => Plaintext(73), A2 => Key(73), Z => n18557);
   U17707 : NAND2_X1 port map( A1 => n15119, A2 => n29626, ZN => n15326);
   U17714 : NAND2_X1 port map( A1 => n23033, A2 => n6605, ZN => n22893);
   U17719 : XOR2_X1 port map( A1 => n51, A2 => n25161, Z => n6607);
   U17722 : XOR2_X1 port map( A1 => n2330, A2 => n6680, Z => n6609);
   U17727 : OAI22_X1 port map( A1 => n18853, A2 => n6860, B1 => n15216, B2 => 
                           n15211, ZN => n6612);
   U17728 : INV_X2 port map( I => n8400, ZN => n15211);
   U17731 : XOR2_X1 port map( A1 => n11691, A2 => n28687, Z => n6614);
   U17737 : XOR2_X1 port map( A1 => n20987, A2 => n6618, Z => n8160);
   U17738 : XOR2_X1 port map( A1 => n20754, A2 => n16666, Z => n6618);
   U17740 : XOR2_X1 port map( A1 => n24783, A2 => n6621, Z => n6620);
   U17741 : XOR2_X1 port map( A1 => n30307, A2 => n16657, Z => n6621);
   U17746 : XOR2_X1 port map( A1 => n6627, A2 => n6628, Z => n8632);
   U17747 : XOR2_X1 port map( A1 => n587, A2 => n9984, Z => n6628);
   U17748 : NAND2_X1 port map( A1 => n33702, A2 => n7555, ZN => n12251);
   U17750 : INV_X2 port map( I => n6634, ZN => n16854);
   U17753 : NAND2_X2 port map( A1 => n6919, A2 => n6918, ZN => n19156);
   U17755 : INV_X2 port map( I => n33393, ZN => n25562);
   U17758 : XOR2_X1 port map( A1 => n24683, A2 => n6647, Z => n6646);
   U17759 : XOR2_X1 port map( A1 => n24474, A2 => n24789, Z => n24683);
   U17762 : XOR2_X1 port map( A1 => n25191, A2 => n27385, Z => n6647);
   U17765 : XOR2_X1 port map( A1 => n1129, A2 => n28005, Z => n6650);
   U17767 : OAI21_X2 port map( A1 => n22770, A2 => n32960, B => n15914, ZN => 
                           n23183);
   U17774 : NOR2_X1 port map( A1 => n16418, A2 => n15108, ZN => n6668);
   U17777 : MUX2_X1 port map( I0 => n14729, I1 => n19959, S => n20112, Z => 
                           n6672);
   U17778 : NAND3_X1 port map( A1 => n6673, A2 => n13624, A3 => n30557, ZN => 
                           n10007);
   U17781 : NAND2_X2 port map( A1 => n16085, A2 => n13580, ZN => n21665);
   U17782 : XNOR2_X1 port map( A1 => n15539, A2 => n6682, ZN => n6681);
   U17783 : XOR2_X1 port map( A1 => n6683, A2 => n15538, Z => n6682);
   U17786 : XOR2_X1 port map( A1 => n6687, A2 => n6688, Z => n6686);
   U17792 : XOR2_X1 port map( A1 => n6701, A2 => n6700, Z => n21228);
   U17796 : XOR2_X1 port map( A1 => n31950, A2 => n17600, Z => n6702);
   U17798 : INV_X2 port map( I => n14834, ZN => n19874);
   U17799 : INV_X2 port map( I => n6705, ZN => n11922);
   U17800 : XOR2_X1 port map( A1 => n6706, A2 => n6708, Z => n6707);
   U17801 : XOR2_X1 port map( A1 => n23300, A2 => n23535, Z => n6708);
   U17802 : XOR2_X1 port map( A1 => n23301, A2 => n10201, Z => n23124);
   U17807 : NOR2_X1 port map( A1 => n29757, A2 => n19143, ZN => n7882);
   U17810 : INV_X2 port map( I => n6725, ZN => n25697);
   U17811 : AOI21_X2 port map( A1 => n13662, A2 => n1327, B => n6728, ZN => 
                           n8291);
   U17813 : NAND3_X2 port map( A1 => n15023, A2 => n21097, A3 => n21098, ZN => 
                           n15022);
   U17819 : XOR2_X1 port map( A1 => n20926, A2 => n25832, Z => n6737);
   U17822 : XOR2_X1 port map( A1 => n16958, A2 => n20715, Z => n6739);
   U17825 : XOR2_X1 port map( A1 => n23256, A2 => n475, Z => n6746);
   U17830 : XOR2_X1 port map( A1 => n6756, A2 => n6755, Z => n6893);
   U17831 : XOR2_X1 port map( A1 => n21033, A2 => n31950, Z => n6755);
   U17834 : XOR2_X1 port map( A1 => n6757, A2 => n4771, Z => n6756);
   U17837 : XOR2_X1 port map( A1 => n6761, A2 => n23524, Z => n6760);
   U17838 : XOR2_X1 port map( A1 => n32899, A2 => n10773, Z => n6761);
   U17839 : XOR2_X1 port map( A1 => n23367, A2 => n2520, Z => n23524);
   U17840 : XOR2_X1 port map( A1 => n8882, A2 => n23248, Z => n6762);
   U17844 : NAND2_X1 port map( A1 => n3909, A2 => n31402, ZN => n22654);
   U17846 : AOI21_X1 port map( A1 => n747, A2 => n14737, B => n32059, ZN => 
                           n7373);
   U17847 : XOR2_X1 port map( A1 => n22285, A2 => n16344, Z => n10422);
   U17848 : XOR2_X1 port map( A1 => n24492, A2 => n7132, Z => n15427);
   U17849 : NAND3_X2 port map( A1 => n6773, A2 => n7729, A3 => n7727, ZN => 
                           n15671);
   U17854 : INV_X1 port map( I => n12317, ZN => n6778);
   U17858 : OAI21_X2 port map( A1 => n6786, A2 => n16473, B => n6784, ZN => 
                           n9472);
   U17862 : XOR2_X1 port map( A1 => n20978, A2 => n10424, Z => n6790);
   U17863 : INV_X1 port map( I => Plaintext(32), ZN => n6791);
   U17864 : XOR2_X1 port map( A1 => n6791, A2 => Key(32), Z => n7194);
   U17865 : INV_X2 port map( I => n7368, ZN => n7195);
   U17866 : OR2_X1 port map( A1 => n22950, A2 => n6798, Z => n6801);
   U17872 : XOR2_X1 port map( A1 => n6808, A2 => n7138, Z => n7137);
   U17875 : XOR2_X1 port map( A1 => n12614, A2 => n6810, Z => n6809);
   U17876 : XOR2_X1 port map( A1 => n9412, A2 => n24386, Z => n6810);
   U17879 : INV_X2 port map( I => n6820, ZN => n9162);
   U17884 : XOR2_X1 port map( A1 => n6827, A2 => n16584, Z => Ciphertext(55));
   U17885 : NAND3_X1 port map( A1 => n1075, A2 => n28736, A3 => n7555, ZN => 
                           n6829);
   U17895 : XOR2_X1 port map( A1 => n11869, A2 => n13393, Z => n6843);
   U17901 : NOR2_X1 port map( A1 => n1214, A2 => n25889, ZN => n24718);
   U17902 : INV_X1 port map( I => n13622, ZN => n12231);
   U17903 : NOR2_X2 port map( A1 => n22326, A2 => n22325, ZN => n16267);
   U17906 : XNOR2_X1 port map( A1 => n15309, A2 => n6856, ZN => n6854);
   U17907 : XOR2_X1 port map( A1 => n29285, A2 => n20998, Z => n6856);
   U17908 : XOR2_X1 port map( A1 => n15, A2 => n25436, Z => n11374);
   U17915 : NAND3_X1 port map( A1 => n6200, A2 => n6263, A3 => n4674, ZN => 
                           n6866);
   U17920 : XOR2_X1 port map( A1 => n21036, A2 => n21037, Z => n6872);
   U17921 : NOR2_X1 port map( A1 => n580, A2 => n1158, ZN => n20616);
   U17923 : NAND2_X1 port map( A1 => n14559, A2 => n16489, ZN => n6930);
   U17924 : XOR2_X1 port map( A1 => n19741, A2 => n25880, Z => n6885);
   U17925 : XOR2_X1 port map( A1 => n27156, A2 => n19424, Z => n19673);
   U17929 : INV_X2 port map( I => n6893, ZN => n12044);
   U17935 : XOR2_X1 port map( A1 => n24638, A2 => n16581, Z => n6897);
   U17936 : XOR2_X1 port map( A1 => n9145, A2 => n24394, Z => n24505);
   U17938 : XOR2_X1 port map( A1 => n15886, A2 => n11194, Z => n6903);
   U17939 : XOR2_X1 port map( A1 => n21019, A2 => n6906, Z => n20700);
   U17942 : NAND2_X1 port map( A1 => n27501, A2 => n30586, ZN => n9846);
   U17943 : NAND2_X1 port map( A1 => n27501, A2 => n24158, ZN => n24313);
   U17945 : XOR2_X1 port map( A1 => n19705, A2 => n487, Z => n6914);
   U17946 : AOI21_X1 port map( A1 => n16854, A2 => n18459, B => n7216, ZN => 
                           n6921);
   U17949 : XOR2_X1 port map( A1 => n32880, A2 => n23474, Z => n6923);
   U17952 : XOR2_X1 port map( A1 => n3322, A2 => n12059, Z => n6924);
   U17955 : NAND2_X1 port map( A1 => n21612, A2 => n17472, ZN => n6937);
   U17956 : INV_X2 port map( I => n6938, ZN => n6939);
   U17958 : XOR2_X1 port map( A1 => n24377, A2 => n6941, Z => n6940);
   U17959 : XOR2_X1 port map( A1 => n24559, A2 => n1411, Z => n6941);
   U17964 : INV_X2 port map( I => n6955, ZN => n12076);
   U17966 : INV_X2 port map( I => n6957, ZN => n21165);
   U17970 : XOR2_X1 port map( A1 => n10159, A2 => n16301, Z => n6966);
   U17972 : AOI21_X1 port map( A1 => n19915, A2 => n19914, B => n6970, ZN => 
                           n19916);
   U17974 : XOR2_X1 port map( A1 => n24771, A2 => n25610, Z => n6973);
   U17977 : NAND2_X1 port map( A1 => n18041, A2 => n2606, ZN => n6999);
   U17988 : INV_X2 port map( I => n7020, ZN => n16650);
   U17990 : INV_X2 port map( I => n7022, ZN => n13905);
   U17992 : INV_X2 port map( I => n21970, ZN => n7023);
   U17994 : XOR2_X1 port map( A1 => n22167, A2 => n11027, Z => n7025);
   U17995 : XOR2_X1 port map( A1 => n7030, A2 => n7031, Z => n7029);
   U18000 : NAND2_X1 port map( A1 => n8820, A2 => n31968, ZN => n8819);
   U18003 : NOR2_X1 port map( A1 => n9985, A2 => n27901, ZN => n11635);
   U18004 : XOR2_X1 port map( A1 => n9467, A2 => n7042, Z => n7043);
   U18005 : INV_X2 port map( I => n7043, ZN => n25700);
   U18010 : OAI21_X1 port map( A1 => n468, A2 => n2417, B => n11250, ZN => 
                           n7052);
   U18013 : AOI22_X2 port map( A1 => n7055, A2 => n7116, B1 => n8353, B2 => 
                           n7054, ZN => n20776);
   U18014 : XOR2_X1 port map( A1 => n7057, A2 => n30305, Z => n14415);
   U18017 : XOR2_X1 port map( A1 => n29137, A2 => n25560, Z => n13435);
   U18024 : XOR2_X1 port map( A1 => n23362, A2 => n7823, Z => n7071);
   U18028 : NOR2_X1 port map( A1 => n7073, A2 => n12906, ZN => n7077);
   U18029 : XOR2_X1 port map( A1 => n3739, A2 => n24895, Z => n9867);
   U18030 : XOR2_X1 port map( A1 => n7078, A2 => n24836, Z => n18138);
   U18031 : INV_X2 port map( I => n7080, ZN => n25232);
   U18032 : INV_X2 port map( I => n17214, ZN => n7081);
   U18038 : NOR2_X1 port map( A1 => n10018, A2 => n7088, ZN => n23221);
   U18042 : NAND2_X1 port map( A1 => n11255, A2 => n24245, ZN => n24128);
   U18046 : NOR2_X1 port map( A1 => n22868, A2 => n28555, ZN => n22869);
   U18047 : NAND2_X1 port map( A1 => n23050, A2 => n28555, ZN => n9950);
   U18048 : XOR2_X1 port map( A1 => n23224, A2 => n1414, Z => n11586);
   U18049 : XOR2_X1 port map( A1 => n17929, A2 => n23224, Z => n12387);
   U18053 : XOR2_X1 port map( A1 => n20839, A2 => n20892, Z => n7113);
   U18056 : INV_X2 port map( I => n21971, ZN => n22411);
   U18057 : XOR2_X1 port map( A1 => n7114, A2 => n21901, Z => n21971);
   U18061 : INV_X2 port map( I => n7250, ZN => n10205);
   U18062 : INV_X2 port map( I => n7124, ZN => n8490);
   U18063 : XNOR2_X1 port map( A1 => n7126, A2 => n7125, ZN => n7124);
   U18064 : XOR2_X1 port map( A1 => n15823, A2 => n20671, Z => n7125);
   U18066 : XOR2_X1 port map( A1 => n9222, A2 => n13739, Z => n7129);
   U18069 : XOR2_X1 port map( A1 => n10331, A2 => n16703, Z => n7132);
   U18072 : XOR2_X1 port map( A1 => n20837, A2 => n20860, Z => n20978);
   U18073 : NAND2_X2 port map( A1 => n20425, A2 => n20424, ZN => n20837);
   U18075 : NAND2_X1 port map( A1 => n7140, A2 => n13281, ZN => n7139);
   U18076 : XOR2_X1 port map( A1 => n22105, A2 => n12127, Z => n7152);
   U18079 : XOR2_X1 port map( A1 => n22318, A2 => n22295, Z => n22273);
   U18080 : NAND2_X1 port map( A1 => n16811, A2 => n19907, ZN => n20118);
   U18084 : AOI21_X2 port map( A1 => n18577, A2 => n33941, B => n7162, ZN => 
                           n7161);
   U18085 : OR2_X1 port map( A1 => n16854, A2 => n11379, Z => n7164);
   U18090 : NAND3_X1 port map( A1 => n26232, A2 => n6230, A3 => n26471, ZN => 
                           n20583);
   U18102 : XOR2_X1 port map( A1 => n16005, A2 => n19763, Z => n19469);
   U18104 : INV_X2 port map( I => n7194, ZN => n15146);
   U18108 : NOR2_X1 port map( A1 => n14940, A2 => n25995, ZN => n7369);
   U18115 : NAND3_X1 port map( A1 => n10511, A2 => n24991, A3 => n10510, ZN => 
                           n7212);
   U18117 : NAND3_X1 port map( A1 => n9320, A2 => n14436, A3 => n7218, ZN => 
                           n9692);
   U18120 : XOR2_X1 port map( A1 => n4157, A2 => n16527, Z => n7222);
   U18121 : NOR2_X1 port map( A1 => n17640, A2 => n4971, ZN => n7224);
   U18122 : INV_X2 port map( I => n18197, ZN => n21170);
   U18125 : XOR2_X1 port map( A1 => n19699, A2 => n5150, Z => n7938);
   U18129 : XOR2_X1 port map( A1 => n16053, A2 => n7229, Z => n23342);
   U18133 : NOR3_X1 port map( A1 => n7776, A2 => n7775, A3 => n7232, ZN => 
                           n7774);
   U18135 : XOR2_X1 port map( A1 => n21041, A2 => n18010, Z => n7235);
   U18138 : NAND2_X1 port map( A1 => n21517, A2 => n21847, ZN => n7241);
   U18144 : XOR2_X1 port map( A1 => n7259, A2 => n7258, Z => n7257);
   U18145 : XOR2_X1 port map( A1 => n24796, A2 => n16696, Z => n7258);
   U18153 : XOR2_X1 port map( A1 => n31523, A2 => n24065, Z => n23452);
   U18160 : XOR2_X1 port map( A1 => n7294, A2 => n1405, Z => n9608);
   U18161 : XOR2_X1 port map( A1 => n21044, A2 => n28983, Z => n14785);
   U18163 : NAND2_X2 port map( A1 => n20368, A2 => n20367, ZN => n7294);
   U18165 : XOR2_X1 port map( A1 => n19733, A2 => n7296, Z => n7295);
   U18166 : XOR2_X1 port map( A1 => n15117, A2 => n16703, Z => n7296);
   U18168 : NAND2_X1 port map( A1 => n7303, A2 => n27920, ZN => n7298);
   U18169 : NOR2_X1 port map( A1 => n7301, A2 => n7300, ZN => n7299);
   U18170 : NOR3_X1 port map( A1 => n7305, A2 => n15359, A3 => n25206, ZN => 
                           n7300);
   U18171 : NOR2_X1 port map( A1 => n7304, A2 => n25206, ZN => n7301);
   U18173 : NOR2_X1 port map( A1 => n10750, A2 => n7308, ZN => n7307);
   U18179 : NAND3_X1 port map( A1 => n5834, A2 => n18683, A3 => n30116, ZN => 
                           n7318);
   U18180 : NOR2_X1 port map( A1 => n26049, A2 => n18683, ZN => n9476);
   U18182 : XOR2_X1 port map( A1 => n20688, A2 => n7331, Z => n7328);
   U18184 : XOR2_X1 port map( A1 => n32749, A2 => n16687, Z => n7331);
   U18186 : XOR2_X1 port map( A1 => n7336, A2 => n25881, Z => Ciphertext(183));
   U18191 : XOR2_X1 port map( A1 => n16693, A2 => n7352, Z => n24798);
   U18192 : XOR2_X1 port map( A1 => n16128, A2 => n24741, Z => n7352);
   U18204 : XOR2_X1 port map( A1 => n7381, A2 => n14748, Z => n7380);
   U18205 : XOR2_X1 port map( A1 => n23511, A2 => n16482, Z => n7382);
   U18207 : XOR2_X1 port map( A1 => n24603, A2 => n15573, Z => n12935);
   U18208 : XOR2_X1 port map( A1 => n7387, A2 => n2363, Z => n14391);
   U18214 : OR2_X1 port map( A1 => n20387, A2 => n53, Z => n7395);
   U18215 : OR2_X1 port map( A1 => n18899, A2 => n878, Z => n7402);
   U18221 : XOR2_X1 port map( A1 => n23230, A2 => n12252, Z => n15055);
   U18223 : AND2_X1 port map( A1 => n22716, A2 => n22808, Z => n7412);
   U18225 : INV_X1 port map( I => n7413, ZN => n10567);
   U18226 : NAND2_X1 port map( A1 => n16274, A2 => n9553, ZN => n7417);
   U18227 : NOR2_X1 port map( A1 => n28707, A2 => n7496, ZN => n17368);
   U18229 : XOR2_X1 port map( A1 => n7431, A2 => n7432, Z => n11942);
   U18230 : XOR2_X1 port map( A1 => n21045, A2 => n8526, Z => n7432);
   U18235 : XOR2_X1 port map( A1 => n25991, A2 => n1405, Z => n7450);
   U18237 : NOR2_X1 port map( A1 => n1063, A2 => n18792, ZN => n18794);
   U18238 : XOR2_X1 port map( A1 => n18350, A2 => Key(30), Z => n15265);
   U18248 : XOR2_X1 port map( A1 => n7471, A2 => n7470, Z => n7469);
   U18249 : XOR2_X1 port map( A1 => n4997, A2 => n16604, Z => n7470);
   U18251 : XOR2_X1 port map( A1 => n10869, A2 => n24774, Z => n7472);
   U18252 : NAND2_X1 port map( A1 => n9025, A2 => n11312, ZN => n11311);
   U18258 : OAI21_X2 port map( A1 => n20299, A2 => n14835, B => n20554, ZN => 
                           n20698);
   U18262 : NOR2_X1 port map( A1 => n4024, A2 => n24201, ZN => n7485);
   U18269 : NAND2_X1 port map( A1 => n470, A2 => n7496, ZN => n7495);
   U18270 : NOR2_X1 port map( A1 => n31407, A2 => n25317, ZN => n11998);
   U18281 : NAND2_X1 port map( A1 => n15906, A2 => n7525, ZN => n9381);
   U18283 : XOR2_X1 port map( A1 => n28953, A2 => n5024, Z => n13209);
   U18284 : XOR2_X1 port map( A1 => n400, A2 => n7530, Z => n9373);
   U18285 : XOR2_X1 port map( A1 => n27275, A2 => n7530, Z => n8053);
   U18291 : INV_X2 port map( I => n10770, ZN => n24780);
   U18292 : XOR2_X1 port map( A1 => n4240, A2 => n1404, Z => n7537);
   U18303 : INV_X1 port map( I => n12609, ZN => n21042);
   U18306 : XOR2_X1 port map( A1 => n31277, A2 => n33693, Z => n7569);
   U18308 : INV_X2 port map( I => n7573, ZN => n18089);
   U18309 : OAI21_X1 port map( A1 => n24657, A2 => n24656, B => n7576, ZN => 
                           n24659);
   U18310 : NAND2_X1 port map( A1 => n31428, A2 => n10325, ZN => n18889);
   U18317 : XOR2_X1 port map( A1 => n8785, A2 => n1365, Z => n7589);
   U18318 : XOR2_X1 port map( A1 => n33749, A2 => n19675, Z => n7590);
   U18320 : NAND2_X1 port map( A1 => n25115, A2 => n18156, ZN => n25020);
   U18324 : XOR2_X1 port map( A1 => n7595, A2 => n5024, Z => n7594);
   U18328 : XOR2_X1 port map( A1 => n17395, A2 => n7598, Z => n7597);
   U18329 : XOR2_X1 port map( A1 => n30331, A2 => n30906, Z => n7598);
   U18330 : XOR2_X1 port map( A1 => n12760, A2 => n16974, Z => n7599);
   U18331 : NOR2_X1 port map( A1 => n7600, A2 => n19255, ZN => n15040);
   U18332 : AOI21_X2 port map( A1 => n24676, A2 => n24799, B => n7604, ZN => 
                           n17811);
   U18333 : XOR2_X1 port map( A1 => n17811, A2 => n16972, Z => n7605);
   U18334 : XOR2_X1 port map( A1 => n13236, A2 => n1432, Z => n7606);
   U18335 : NOR2_X1 port map( A1 => n7609, A2 => n12038, ZN => n19997);
   U18337 : XOR2_X1 port map( A1 => n7611, A2 => n9641, Z => n9640);
   U18338 : XOR2_X1 port map( A1 => n9006, A2 => n10210, Z => n7611);
   U18340 : XOR2_X1 port map( A1 => n23245, A2 => n7615, Z => n7614);
   U18341 : XOR2_X1 port map( A1 => n23186, A2 => n16605, Z => n7615);
   U18343 : XOR2_X1 port map( A1 => n32930, A2 => n19582, Z => n7619);
   U18346 : XOR2_X1 port map( A1 => n20904, A2 => n25610, Z => n7622);
   U18347 : XOR2_X1 port map( A1 => n8795, A2 => n20905, Z => n7623);
   U18348 : INV_X1 port map( I => n32051, ZN => n18518);
   U18350 : INV_X2 port map( I => n7624, ZN => n25889);
   U18352 : XOR2_X1 port map( A1 => n20736, A2 => n1923, Z => n7628);
   U18353 : AOI22_X2 port map( A1 => n9852, A2 => n16050, B1 => n7631, B2 => 
                           n14011, ZN => n20614);
   U18354 : XOR2_X1 port map( A1 => n19588, A2 => n7635, Z => n7634);
   U18355 : XOR2_X1 port map( A1 => n29890, A2 => n207, Z => n7635);
   U18360 : XOR2_X1 port map( A1 => n29011, A2 => n16464, Z => n7638);
   U18363 : XOR2_X1 port map( A1 => n21910, A2 => n21958, Z => n22046);
   U18368 : XOR2_X1 port map( A1 => n20648, A2 => n7645, Z => n7644);
   U18369 : XOR2_X1 port map( A1 => n20996, A2 => n12957, Z => n7645);
   U18370 : XOR2_X1 port map( A1 => n20698, A2 => n20954, Z => n20648);
   U18371 : XOR2_X1 port map( A1 => n19703, A2 => n27281, Z => n7652);
   U18372 : XOR2_X1 port map( A1 => n32581, A2 => n25465, Z => n20858);
   U18378 : INV_X2 port map( I => n7657, ZN => n21070);
   U18379 : NOR2_X1 port map( A1 => n4202, A2 => n30010, ZN => n9315);
   U18381 : NOR2_X1 port map( A1 => n8408, A2 => n23867, ZN => n7663);
   U18382 : INV_X2 port map( I => n15356, ZN => n19938);
   U18384 : XOR2_X1 port map( A1 => n2894, A2 => n24917, Z => n7664);
   U18386 : XOR2_X1 port map( A1 => n8997, A2 => n25131, Z => n7675);
   U18388 : XOR2_X1 port map( A1 => n19632, A2 => n1196, Z => n7676);
   U18394 : XOR2_X1 port map( A1 => n22076, A2 => n22158, Z => n21919);
   U18396 : NAND2_X1 port map( A1 => n12358, A2 => n7689, ZN => n7688);
   U18399 : XOR2_X1 port map( A1 => n29318, A2 => n1397, Z => n7693);
   U18400 : XOR2_X1 port map( A1 => n356, A2 => n25990, Z => n7694);
   U18404 : INV_X2 port map( I => n7700, ZN => n8408);
   U18406 : NAND2_X2 port map( A1 => n17022, A2 => n17023, ZN => n7702);
   U18407 : NOR2_X1 port map( A1 => n25916, A2 => n7701, ZN => n25907);
   U18409 : NOR2_X1 port map( A1 => n31476, A2 => n1018, ZN => n21272);
   U18413 : INV_X2 port map( I => n7712, ZN => n16420);
   U18414 : NAND2_X1 port map( A1 => n9272, A2 => n1287, ZN => n11866);
   U18418 : MUX2_X1 port map( I0 => n26950, I1 => n9323, S => n7809, Z => n7730
                           );
   U18420 : XOR2_X1 port map( A1 => n7731, A2 => n16687, Z => n11484);
   U18421 : NOR2_X1 port map( A1 => n8862, A2 => n7732, ZN => n8867);
   U18425 : NAND2_X1 port map( A1 => n2444, A2 => n1244, ZN => n23621);
   U18426 : NAND2_X1 port map( A1 => n24111, A2 => n1244, ZN => n24112);
   U18427 : NOR2_X1 port map( A1 => n15977, A2 => n1244, ZN => n10177);
   U18431 : INV_X2 port map( I => n7912, ZN => n10187);
   U18435 : XOR2_X1 port map( A1 => n9904, A2 => n33749, Z => n7741);
   U18440 : AOI22_X2 port map( A1 => n7745, A2 => n22864, B1 => n7744, B2 => 
                           n14978, ZN => n23262);
   U18442 : NAND2_X1 port map( A1 => n31019, A2 => n12488, ZN => n17268);
   U18447 : XOR2_X1 port map( A1 => n7838, A2 => n17296, Z => n7761);
   U18449 : OAI21_X1 port map( A1 => n25154, A2 => n7765, B => n25175, ZN => 
                           n16098);
   U18452 : XOR2_X1 port map( A1 => n7772, A2 => n16355, Z => n23472);
   U18457 : AOI21_X1 port map( A1 => n3994, A2 => n24936, B => n15799, ZN => 
                           n7785);
   U18462 : XOR2_X1 port map( A1 => n7794, A2 => n7793, Z => n24870);
   U18463 : XOR2_X1 port map( A1 => n28258, A2 => n7795, Z => n7793);
   U18465 : XOR2_X1 port map( A1 => n30301, A2 => n7511, Z => n7795);
   U18467 : INV_X1 port map( I => n14201, ZN => n22855);
   U18470 : NAND2_X1 port map( A1 => n29253, A2 => n27345, ZN => n7803);
   U18473 : XOR2_X1 port map( A1 => n7808, A2 => n14300, Z => n14299);
   U18477 : XOR2_X1 port map( A1 => n31950, A2 => n16038, Z => n16754);
   U18478 : XOR2_X1 port map( A1 => n27708, A2 => n25036, Z => n7823);
   U18484 : XOR2_X1 port map( A1 => n7828, A2 => n16530, Z => n7829);
   U18487 : NOR2_X1 port map( A1 => n24995, A2 => n7831, ZN => n14450);
   U18492 : OR2_X1 port map( A1 => n25677, A2 => n25678, Z => n7842);
   U18494 : XOR2_X1 port map( A1 => n22139, A2 => n30332, Z => n16837);
   U18498 : XOR2_X1 port map( A1 => n7859, A2 => n18231, Z => n11220);
   U18499 : XOR2_X1 port map( A1 => n24826, A2 => n1426, Z => n7860);
   U18500 : XOR2_X1 port map( A1 => n28579, A2 => n12313, Z => n7861);
   U18503 : INV_X2 port map( I => n7865, ZN => n13969);
   U18504 : XOR2_X1 port map( A1 => n15357, A2 => n15819, Z => n7866);
   U18505 : XOR2_X1 port map( A1 => n1341, A2 => n7960, Z => n7870);
   U18508 : XOR2_X1 port map( A1 => n16080, A2 => n7875, Z => n7874);
   U18519 : XOR2_X1 port map( A1 => n13457, A2 => n7888, Z => n13491);
   U18521 : XOR2_X1 port map( A1 => n20906, A2 => n447, Z => n7890);
   U18524 : NAND2_X1 port map( A1 => n7895, A2 => n1099, ZN => n23649);
   U18525 : NAND2_X1 port map( A1 => n7895, A2 => n27455, ZN => n23348);
   U18529 : NOR2_X1 port map( A1 => n6215, A2 => n1430, ZN => n7900);
   U18530 : XOR2_X1 port map( A1 => Plaintext(65), A2 => Key(65), Z => n18186);
   U18533 : XOR2_X1 port map( A1 => n24686, A2 => n10924, Z => n24524);
   U18534 : AOI21_X2 port map( A1 => n11121, A2 => n28120, B => n24169, ZN => 
                           n24686);
   U18537 : XOR2_X1 port map( A1 => n7910, A2 => n7909, Z => n14307);
   U18538 : XOR2_X1 port map( A1 => n16896, A2 => n15778, Z => n7909);
   U18539 : XOR2_X1 port map( A1 => n12495, A2 => n7911, Z => n7910);
   U18543 : XOR2_X1 port map( A1 => n23121, A2 => n22948, Z => n7916);
   U18544 : XOR2_X1 port map( A1 => n23184, A2 => n22954, Z => n7917);
   U18545 : NAND2_X1 port map( A1 => n8467, A2 => n17439, ZN => n8466);
   U18546 : INV_X2 port map( I => n7918, ZN => n17439);
   U18548 : XOR2_X1 port map( A1 => n17766, A2 => n15121, Z => n7931);
   U18550 : NAND2_X2 port map( A1 => n21742, A2 => n14041, ZN => n9960);
   U18551 : XOR2_X1 port map( A1 => n11784, A2 => n7934, Z => n7933);
   U18552 : XOR2_X1 port map( A1 => n22294, A2 => n22295, Z => n7934);
   U18555 : XOR2_X1 port map( A1 => n7939, A2 => n7936, Z => n12241);
   U18556 : XOR2_X1 port map( A1 => n7937, A2 => n7938, Z => n7936);
   U18559 : NAND2_X1 port map( A1 => n713, A2 => n7941, ZN => n14451);
   U18560 : NAND2_X2 port map( A1 => n13940, A2 => n9422, ZN => n19230);
   U18561 : OAI21_X2 port map( A1 => n21310, A2 => n21447, B => n21309, ZN => 
                           n21662);
   U18566 : XOR2_X1 port map( A1 => n22168, A2 => n28926, Z => n22247);
   U18571 : AND2_X1 port map( A1 => n19130, A2 => n7966, Z => n16363);
   U18572 : INV_X2 port map( I => n11379, ZN => n18459);
   U18579 : XOR2_X1 port map( A1 => n19546, A2 => n19690, Z => n7988);
   U18581 : XOR2_X1 port map( A1 => n19734, A2 => n19401, Z => n7989);
   U18583 : INV_X2 port map( I => n7993, ZN => n23795);
   U18585 : XOR2_X1 port map( A1 => n7999, A2 => n22250, Z => n7998);
   U18590 : XOR2_X1 port map( A1 => n8701, A2 => n17999, Z => n8700);
   U18593 : XOR2_X1 port map( A1 => n23393, A2 => n16454, Z => n8018);
   U18595 : XOR2_X1 port map( A1 => n8021, A2 => n23403, Z => n8020);
   U18596 : XOR2_X1 port map( A1 => n11193, A2 => n27613, Z => n8021);
   U18601 : NAND2_X1 port map( A1 => n12827, A2 => n8029, ZN => n8030);
   U18602 : XOR2_X1 port map( A1 => n27169, A2 => n3929, Z => n20695);
   U18604 : INV_X2 port map( I => n14788, ZN => n17110);
   U18605 : XOR2_X1 port map( A1 => n10617, A2 => n10616, Z => n14788);
   U18607 : NAND2_X2 port map( A1 => n17959, A2 => n22527, ZN => n22983);
   U18609 : INV_X2 port map( I => n8042, ZN => n23742);
   U18619 : XOR2_X1 port map( A1 => n8050, A2 => n24646, Z => n24411);
   U18622 : XOR2_X1 port map( A1 => n13339, A2 => n1024, Z => n13338);
   U18624 : INV_X1 port map( I => n9481, ZN => n9479);
   U18631 : NAND2_X2 port map( A1 => n19241, A2 => n19240, ZN => n19676);
   U18632 : NOR2_X2 port map( A1 => n19239, A2 => n19238, ZN => n19779);
   U18633 : NOR2_X1 port map( A1 => n8058, A2 => n24106, ZN => n14375);
   U18634 : NOR2_X1 port map( A1 => n17310, A2 => n8058, ZN => n12098);
   U18636 : XOR2_X1 port map( A1 => n8060, A2 => n8059, Z => n8721);
   U18638 : XOR2_X1 port map( A1 => n27130, A2 => n16060, Z => n8061);
   U18641 : NOR2_X1 port map( A1 => n13102, A2 => n23930, ZN => n8063);
   U18643 : XOR2_X1 port map( A1 => n32895, A2 => n8066, Z => n8065);
   U18644 : XOR2_X1 port map( A1 => n23519, A2 => n25465, Z => n8066);
   U18645 : XOR2_X1 port map( A1 => n23518, A2 => n23520, Z => n8067);
   U18648 : XOR2_X1 port map( A1 => n23125, A2 => n15049, Z => n8070);
   U18651 : AOI21_X1 port map( A1 => n712, A2 => n14810, B => n6402, ZN => 
                           n25125);
   U18655 : XOR2_X1 port map( A1 => n22296, A2 => n16381, Z => n21878);
   U18657 : XOR2_X1 port map( A1 => n16138, A2 => n16110, Z => n8089);
   U18667 : NOR2_X2 port map( A1 => n21306, A2 => n21305, ZN => n8106);
   U18673 : XOR2_X1 port map( A1 => n13695, A2 => n25009, Z => n8112);
   U18674 : XOR2_X1 port map( A1 => n14899, A2 => n20318, Z => n8116);
   U18676 : XOR2_X1 port map( A1 => n23387, A2 => n25772, Z => n8129);
   U18677 : XOR2_X1 port map( A1 => n10205, A2 => n1064, Z => n22194);
   U18678 : XOR2_X1 port map( A1 => n8133, A2 => n8132, Z => n9871);
   U18679 : XOR2_X1 port map( A1 => n21927, A2 => n10429, Z => n8132);
   U18683 : XOR2_X1 port map( A1 => n30729, A2 => n8139, Z => n12103);
   U18684 : XOR2_X1 port map( A1 => n30729, A2 => n16631, Z => n19316);
   U18686 : NAND2_X2 port map( A1 => n18769, A2 => n17905, ZN => n8141);
   U18694 : NAND2_X2 port map( A1 => n12371, A2 => n12373, ZN => n8313);
   U18697 : NAND2_X2 port map( A1 => n21609, A2 => n21608, ZN => n22021);
   U18702 : NAND2_X1 port map( A1 => n32605, A2 => n22608, ZN => n12112);
   U18706 : OAI21_X1 port map( A1 => n18583, A2 => n12190, B => n18582, ZN => 
                           n12191);
   U18715 : NOR2_X1 port map( A1 => n22690, A2 => n16205, ZN => n9603);
   U18716 : OAI21_X1 port map( A1 => n17709, A2 => n17708, B => n8629, ZN => 
                           n11558);
   U18718 : OAI21_X1 port map( A1 => n15858, A2 => n32867, B => n25312, ZN => 
                           n15857);
   U18725 : XOR2_X1 port map( A1 => n11434, A2 => n11432, Z => n16904);
   U18727 : NAND2_X2 port map( A1 => n8481, A2 => n11347, ZN => n9247);
   U18730 : INV_X1 port map( I => n12498, ZN => n12497);
   U18736 : XOR2_X1 port map( A1 => Plaintext(170), A2 => Key(170), Z => n18411
                           );
   U18738 : XOR2_X1 port map( A1 => n19587, A2 => n32844, Z => n15044);
   U18748 : NAND2_X1 port map( A1 => n21653, A2 => n21595, ZN => n21596);
   U18749 : OR2_X1 port map( A1 => n29658, A2 => n8208, Z => n10786);
   U18756 : NOR2_X1 port map( A1 => n24328, A2 => n10987, ZN => n10342);
   U18757 : INV_X2 port map( I => n18182, ZN => n10213);
   U18760 : INV_X2 port map( I => n8213, ZN => n18880);
   U18762 : XOR2_X1 port map( A1 => n24845, A2 => n8215, Z => n8214);
   U18764 : NAND2_X1 port map( A1 => n23105, A2 => n22971, ZN => n11623);
   U18772 : OAI22_X1 port map( A1 => n19022, A2 => n19023, B1 => n19021, B2 => 
                           n19290, ZN => n8227);
   U18773 : AOI21_X1 port map( A1 => n17850, A2 => n25463, B => n25470, ZN => 
                           n17849);
   U18774 : INV_X2 port map( I => n8228, ZN => n9133);
   U18778 : XOR2_X1 port map( A1 => n1341, A2 => n11636, Z => n8232);
   U18785 : XOR2_X1 port map( A1 => n8236, A2 => n31094, Z => Ciphertext(122));
   U18786 : NAND3_X1 port map( A1 => n25548, A2 => n17401, A3 => n25547, ZN => 
                           n8236);
   U18787 : XOR2_X1 port map( A1 => n24578, A2 => n14250, Z => n17504);
   U18792 : XOR2_X1 port map( A1 => n8241, A2 => n30275, Z => n11271);
   U18793 : INV_X1 port map( I => n9536, ZN => n8241);
   U18803 : NAND2_X1 port map( A1 => n7144, A2 => n21876, ZN => n8253);
   U18806 : XNOR2_X1 port map( A1 => n32255, A2 => n22078, ZN => n9208);
   U18812 : NOR2_X1 port map( A1 => n881, A2 => n6295, ZN => n18318);
   U18813 : OR2_X1 port map( A1 => n15397, A2 => n19330, Z => n19155);
   U18814 : XOR2_X1 port map( A1 => n8556, A2 => n14429, Z => n14534);
   U18821 : XOR2_X1 port map( A1 => n11574, A2 => n8266, Z => n8265);
   U18824 : NOR2_X1 port map( A1 => n4373, A2 => n16848, ZN => n19818);
   U18825 : NAND2_X1 port map( A1 => n17670, A2 => n33561, ZN => n12253);
   U18830 : AOI21_X1 port map( A1 => n23108, A2 => n6453, B => n23111, ZN => 
                           n9042);
   U18837 : XOR2_X1 port map( A1 => n22099, A2 => n22031, Z => n8282);
   U18844 : OAI21_X1 port map( A1 => n17877, A2 => n298, B => n11257, ZN => 
                           n17876);
   U18849 : INV_X1 port map( I => n21160, ZN => n21139);
   U18855 : XOR2_X1 port map( A1 => n20710, A2 => n20709, Z => n11542);
   U18859 : OR2_X1 port map( A1 => n17403, A2 => n13483, Z => n25548);
   U18860 : NAND2_X1 port map( A1 => n11646, A2 => n28203, ZN => n11645);
   U18864 : AND2_X1 port map( A1 => n1099, A2 => n29323, Z => n12026);
   U18869 : OR3_X1 port map( A1 => n17156, A2 => n17155, A3 => n4587, Z => 
                           n10850);
   U18870 : XOR2_X1 port map( A1 => n12342, A2 => n20921, Z => n20758);
   U18872 : INV_X1 port map( I => n9612, ZN => n9611);
   U18885 : AND2_X1 port map( A1 => n10574, A2 => n27149, Z => n9676);
   U18890 : NOR2_X1 port map( A1 => n10549, A2 => n18219, ZN => n8470);
   U18893 : NOR2_X1 port map( A1 => n23670, A2 => n29198, ZN => n9344);
   U18895 : XOR2_X1 port map( A1 => n12681, A2 => n22221, Z => n8324);
   U18900 : XOR2_X1 port map( A1 => n8557, A2 => n8987, Z => n10372);
   U18907 : NOR2_X2 port map( A1 => n11983, A2 => n31854, ZN => n22781);
   U18910 : AND2_X1 port map( A1 => n21676, A2 => n15595, Z => n8331);
   U18911 : OR2_X1 port map( A1 => n18955, A2 => n18983, Z => n18964);
   U18915 : AND3_X1 port map( A1 => n14321, A2 => n24995, A3 => n24996, Z => 
                           n9901);
   U18919 : XOR2_X1 port map( A1 => n21892, A2 => n30332, Z => n10963);
   U18928 : XOR2_X1 port map( A1 => n8341, A2 => n14216, Z => n22156);
   U18929 : NAND2_X1 port map( A1 => n9273, A2 => n6908, ZN => n8958);
   U18934 : XOR2_X1 port map( A1 => n8345, A2 => n16402, Z => Ciphertext(172));
   U18941 : XOR2_X1 port map( A1 => n22018, A2 => n521, Z => n8352);
   U18946 : XOR2_X1 port map( A1 => n8361, A2 => n11600, Z => n9753);
   U18948 : XOR2_X1 port map( A1 => n21885, A2 => n16439, Z => n17109);
   U18953 : XOR2_X1 port map( A1 => n14400, A2 => n8364, Z => n12670);
   U18954 : XOR2_X1 port map( A1 => n14647, A2 => n14646, Z => n8364);
   U18956 : XOR2_X1 port map( A1 => n11282, A2 => n8366, Z => n11281);
   U18965 : NAND3_X1 port map( A1 => n10897, A2 => n27162, A3 => n25851, ZN => 
                           n18021);
   U18968 : XOR2_X1 port map( A1 => n19406, A2 => n445, Z => n8383);
   U18977 : AND2_X1 port map( A1 => n11987, A2 => n28591, Z => n14895);
   U18984 : XOR2_X1 port map( A1 => n8394, A2 => n25910, Z => Ciphertext(188));
   U18986 : NAND2_X2 port map( A1 => n12690, A2 => n12689, ZN => n8457);
   U18987 : XOR2_X1 port map( A1 => n10916, A2 => n10914, Z => n14834);
   U18988 : NOR2_X1 port map( A1 => n8397, A2 => n25416, ZN => n25417);
   U18989 : AOI21_X1 port map( A1 => n25415, A2 => n25418, B => n25452, ZN => 
                           n8397);
   U18994 : XOR2_X1 port map( A1 => Key(159), A2 => Plaintext(159), Z => n8400)
                           ;
   U18995 : INV_X4 port map( I => n9162, ZN => n14922);
   U18997 : INV_X2 port map( I => n20091, ZN => n19936);
   U18998 : XOR2_X1 port map( A1 => n14222, A2 => n8401, Z => n20091);
   U18999 : INV_X1 port map( I => n16007, ZN => n14611);
   U19000 : AND2_X1 port map( A1 => n16275, A2 => n599, Z => n12743);
   U19001 : NOR2_X1 port map( A1 => n21590, A2 => n7144, ZN => n8402);
   U19003 : XOR2_X1 port map( A1 => n10076, A2 => n8405, Z => n22390);
   U19008 : XOR2_X1 port map( A1 => n27852, A2 => n322, Z => n8413);
   U19012 : NAND2_X2 port map( A1 => n985, A2 => n9280, ZN => n8786);
   U19014 : INV_X2 port map( I => n10860, ZN => n11198);
   U19015 : XOR2_X1 port map( A1 => n10861, A2 => n8416, Z => n10860);
   U19021 : XOR2_X1 port map( A1 => Plaintext(94), A2 => Key(94), Z => n16782);
   U19023 : INV_X2 port map( I => n8422, ZN => n10080);
   U19026 : XOR2_X1 port map( A1 => n11320, A2 => n15565, Z => n8424);
   U19029 : XNOR2_X1 port map( A1 => n22014, A2 => n16587, ZN => n8979);
   U19038 : INV_X2 port map( I => n8435, ZN => n19947);
   U19043 : XOR2_X1 port map( A1 => n8440, A2 => n1426, Z => Ciphertext(33));
   U19045 : INV_X1 port map( I => n17578, ZN => n23870);
   U19047 : NOR2_X1 port map( A1 => n29294, A2 => n10187, ZN => n10753);
   U19050 : INV_X2 port map( I => n8444, ZN => n11945);
   U19051 : XOR2_X1 port map( A1 => n14886, A2 => n14883, Z => n8444);
   U19065 : XNOR2_X1 port map( A1 => n19773, A2 => n13826, ZN => n15188);
   U19072 : OR2_X1 port map( A1 => n21490, A2 => n21489, Z => n8463);
   U19077 : NAND2_X1 port map( A1 => n34097, A2 => n15976, ZN => n11740);
   U19078 : INV_X2 port map( I => n8469, ZN => n21109);
   U19080 : INV_X2 port map( I => n10372, ZN => n25867);
   U19082 : XOR2_X1 port map( A1 => n6569, A2 => n16701, Z => n8475);
   U19084 : OR2_X1 port map( A1 => n17879, A2 => n22580, Z => n22348);
   U19099 : NAND2_X1 port map( A1 => n31549, A2 => n23103, ZN => n8494);
   U19101 : XOR2_X1 port map( A1 => n10391, A2 => n8496, Z => n10390);
   U19103 : XOR2_X1 port map( A1 => n3722, A2 => n22078, Z => n8497);
   U19108 : XOR2_X1 port map( A1 => n8997, A2 => n8500, Z => n11066);
   U19111 : INV_X1 port map( I => n9839, ZN => n10886);
   U19114 : INV_X2 port map( I => n8505, ZN => n11920);
   U19115 : XOR2_X1 port map( A1 => n14298, A2 => n14301, Z => n8505);
   U19116 : XOR2_X1 port map( A1 => n24777, A2 => n24778, Z => n16719);
   U19117 : XOR2_X1 port map( A1 => n8507, A2 => n24643, Z => n24777);
   U19120 : NAND2_X1 port map( A1 => n25804, A2 => n25818, ZN => n25819);
   U19123 : NOR2_X2 port map( A1 => n8515, A2 => n9956, ZN => n25072);
   U19125 : XNOR2_X1 port map( A1 => n19544, A2 => n19446, ZN => n16678);
   U19128 : XOR2_X1 port map( A1 => n24679, A2 => n24678, Z => n24680);
   U19132 : XOR2_X1 port map( A1 => n8949, A2 => n25878, Z => n8531);
   U19133 : XOR2_X1 port map( A1 => n19742, A2 => n13222, Z => n8532);
   U19134 : NAND2_X1 port map( A1 => n23822, A2 => n11887, ZN => n18152);
   U19135 : XOR2_X1 port map( A1 => n8536, A2 => n16587, Z => Ciphertext(60));
   U19137 : NAND2_X1 port map( A1 => n14531, A2 => n25140, ZN => n15228);
   U19142 : XOR2_X1 port map( A1 => n23196, A2 => n16160, Z => n23373);
   U19145 : NAND2_X1 port map( A1 => n8542, A2 => n8541, ZN => n10100);
   U19148 : NOR2_X1 port map( A1 => n21478, A2 => n32904, ZN => n9590);
   U19150 : AND2_X1 port map( A1 => n23882, A2 => n8544, Z => n10621);
   U19153 : INV_X2 port map( I => n8545, ZN => n11966);
   U19157 : AOI22_X1 port map( A1 => n25153, A2 => n25179, B1 => n14531, B2 => 
                           n25174, ZN => n17635);
   U19161 : NAND2_X2 port map( A1 => n8551, A2 => n8550, ZN => n19104);
   U19162 : XOR2_X1 port map( A1 => n24762, A2 => n24541, Z => n14886);
   U19166 : OAI21_X2 port map( A1 => n11318, A2 => n11319, B => n8554, ZN => 
                           n18257);
   U19169 : XOR2_X1 port map( A1 => n24793, A2 => n17858, Z => n8557);
   U19172 : XOR2_X1 port map( A1 => n19698, A2 => n23239, Z => n8561);
   U19174 : XOR2_X1 port map( A1 => n19527, A2 => n19526, Z => n20137);
   U19176 : NAND2_X1 port map( A1 => n8664, A2 => n24276, ZN => n8663);
   U19186 : NAND2_X1 port map( A1 => n19233, A2 => n19274, ZN => n9407);
   U19190 : OAI21_X2 port map( A1 => n8581, A2 => n11636, B => n8578, ZN => 
                           n12539);
   U19192 : XOR2_X1 port map( A1 => n1340, A2 => n11349, Z => n8583);
   U19194 : NAND2_X1 port map( A1 => n32857, A2 => n28228, ZN => n25089);
   U19200 : XOR2_X1 port map( A1 => n19503, A2 => n13829, Z => n10060);
   U19211 : NOR2_X1 port map( A1 => n19229, A2 => n8606, ZN => n11807);
   U19218 : INV_X2 port map( I => n18541, ZN => n13279);
   U19222 : XOR2_X1 port map( A1 => n8633, A2 => n16679, Z => n13951);
   U19223 : XOR2_X1 port map( A1 => n8633, A2 => n12998, Z => n12519);
   U19224 : INV_X2 port map( I => n8634, ZN => n17895);
   U19226 : XOR2_X1 port map( A1 => n8480, A2 => n25827, Z => n8635);
   U19228 : INV_X2 port map( I => n24947, ZN => n24958);
   U19232 : XOR2_X1 port map( A1 => n32243, A2 => n8659, Z => n23390);
   U19233 : INV_X1 port map( I => Plaintext(33), ZN => n8666);
   U19234 : XOR2_X1 port map( A1 => n8666, A2 => Key(33), Z => n10058);
   U19237 : NOR2_X1 port map( A1 => n25787, A2 => n8678, ZN => n16670);
   U19239 : OAI21_X1 port map( A1 => n25798, A2 => n26753, B => n12611, ZN => 
                           n25799);
   U19240 : NAND2_X1 port map( A1 => n25782, A2 => n26753, ZN => n17222);
   U19243 : INV_X2 port map( I => n8681, ZN => n21253);
   U19245 : XOR2_X1 port map( A1 => n31491, A2 => n25619, Z => n23307);
   U19247 : XOR2_X1 port map( A1 => n19589, A2 => n13826, Z => n8685);
   U19249 : XOR2_X1 port map( A1 => n19644, A2 => n19368, Z => n19446);
   U19252 : INV_X1 port map( I => n29130, ZN => n19337);
   U19253 : XOR2_X1 port map( A1 => n29130, A2 => n25167, Z => n13843);
   U19255 : XOR2_X1 port map( A1 => n31279, A2 => n1432, Z => n13854);
   U19259 : INV_X2 port map( I => n8694, ZN => n23695);
   U19261 : XOR2_X1 port map( A1 => Plaintext(166), A2 => Key(166), Z => n18860
                           );
   U19262 : NAND2_X1 port map( A1 => n4683, A2 => n8010, ZN => n16543);
   U19263 : XOR2_X1 port map( A1 => n24539, A2 => n24454, Z => n24398);
   U19268 : XOR2_X1 port map( A1 => n8707, A2 => n24869, Z => Ciphertext(115));
   U19269 : OAI21_X1 port map( A1 => n8766, A2 => n25515, B => n25509, ZN => 
                           n8708);
   U19270 : NOR2_X1 port map( A1 => n8766, A2 => n25516, ZN => n8709);
   U19272 : XOR2_X1 port map( A1 => n8718, A2 => n9263, Z => n8715);
   U19274 : AOI21_X1 port map( A1 => n28736, A2 => n7555, B => n25129, ZN => 
                           n8722);
   U19277 : INV_X1 port map( I => n19164, ZN => n9652);
   U19278 : INV_X1 port map( I => n8237, ZN => n15029);
   U19279 : XOR2_X1 port map( A1 => n28889, A2 => n11490, Z => n19785);
   U19281 : XOR2_X1 port map( A1 => n29838, A2 => n16696, Z => n16949);
   U19282 : XOR2_X1 port map( A1 => n29838, A2 => n25091, Z => n20709);
   U19283 : AOI21_X1 port map( A1 => n17814, A2 => n33480, B => n25902, ZN => 
                           n17621);
   U19284 : NOR2_X1 port map( A1 => n11754, A2 => n1090, ZN => n8731);
   U19285 : NAND2_X2 port map( A1 => n21597, A2 => n21596, ZN => n22210);
   U19287 : NAND2_X1 port map( A1 => n13663, A2 => n11918, ZN => n8737);
   U19290 : AOI21_X1 port map( A1 => n8212, A2 => n8742, B => n33672, ZN => 
                           n14500);
   U19295 : XOR2_X1 port map( A1 => n8747, A2 => n8745, Z => n10171);
   U19296 : XOR2_X1 port map( A1 => n10729, A2 => n8746, Z => n8745);
   U19297 : XOR2_X1 port map( A1 => n11332, A2 => n1193, Z => n8746);
   U19300 : XOR2_X1 port map( A1 => n11166, A2 => n22210, Z => n8750);
   U19307 : XOR2_X1 port map( A1 => n19677, A2 => n8755, Z => n8754);
   U19313 : XOR2_X1 port map( A1 => n8765, A2 => n8763, Z => n10463);
   U19314 : XOR2_X1 port map( A1 => n23190, A2 => n8764, Z => n8763);
   U19315 : XOR2_X1 port map( A1 => n29235, A2 => n1064, Z => n8764);
   U19316 : XOR2_X1 port map( A1 => n29217, A2 => n29299, Z => n23190);
   U19317 : NAND2_X1 port map( A1 => n8770, A2 => n31522, ZN => n8769);
   U19318 : XOR2_X1 port map( A1 => n19739, A2 => n19211, Z => n8771);
   U19320 : XOR2_X1 port map( A1 => n31755, A2 => n12620, Z => n8772);
   U19322 : NAND2_X1 port map( A1 => n17655, A2 => n30316, ZN => n8773);
   U19323 : XOR2_X1 port map( A1 => n32894, A2 => n1427, Z => n8774);
   U19326 : NAND2_X1 port map( A1 => n31161, A2 => n1172, ZN => n8782);
   U19327 : XOR2_X1 port map( A1 => n8791, A2 => n12355, Z => n10350);
   U19335 : XOR2_X1 port map( A1 => n12958, A2 => n8806, Z => n8808);
   U19338 : XOR2_X1 port map( A1 => n23163, A2 => n8812, Z => n8811);
   U19339 : XOR2_X1 port map( A1 => n23260, A2 => n16533, Z => n8812);
   U19342 : XOR2_X1 port map( A1 => Plaintext(79), A2 => Key(79), Z => n16881);
   U19346 : XOR2_X1 port map( A1 => n14858, A2 => n1065, Z => n8826);
   U19348 : XNOR2_X1 port map( A1 => Plaintext(119), A2 => Key(119), ZN => 
                           n8832);
   U19350 : XOR2_X1 port map( A1 => n8845, A2 => n8843, Z => n17641);
   U19352 : XOR2_X1 port map( A1 => n32870, A2 => n24618, Z => n8844);
   U19363 : NAND2_X1 port map( A1 => n8860, A2 => n18738, ZN => n18124);
   U19364 : NAND2_X1 port map( A1 => n25744, A2 => n1597, ZN => n25740);
   U19365 : NAND2_X1 port map( A1 => n25737, A2 => n25748, ZN => n25742);
   U19366 : XOR2_X1 port map( A1 => n30314, A2 => n22274, Z => n8861);
   U19369 : NOR3_X1 port map( A1 => n18261, A2 => n30365, A3 => n25979, ZN => 
                           n8876);
   U19375 : XOR2_X1 port map( A1 => n23247, A2 => n8883, Z => n8882);
   U19379 : INV_X2 port map( I => n34169, ZN => n25590);
   U19380 : OR2_X1 port map( A1 => n34169, A2 => n8892, Z => n25529);
   U19383 : XOR2_X1 port map( A1 => n24624, A2 => n8895, Z => n8894);
   U19384 : XOR2_X1 port map( A1 => n24625, A2 => n13556, Z => n8896);
   U19385 : XOR2_X1 port map( A1 => n9217, A2 => n609, Z => n8899);
   U19386 : INV_X2 port map( I => n8899, ZN => n21056);
   U19387 : NOR2_X1 port map( A1 => n8901, A2 => n25587, ZN => n10395);
   U19388 : MUX2_X1 port map( I0 => n24075, I1 => n24127, S => n1235, Z => 
                           n24078);
   U19391 : XOR2_X1 port map( A1 => n24689, A2 => n25065, Z => n17325);
   U19392 : XOR2_X1 port map( A1 => n24689, A2 => n24964, Z => n10195);
   U19393 : XOR2_X1 port map( A1 => n23209, A2 => n1196, Z => n8916);
   U19394 : XOR2_X1 port map( A1 => n23257, A2 => n15497, Z => n8917);
   U19395 : XOR2_X1 port map( A1 => n24764, A2 => n25036, Z => n8920);
   U19396 : XOR2_X1 port map( A1 => n4028, A2 => n480, Z => n8922);
   U19397 : NAND2_X1 port map( A1 => n8207, A2 => n28196, ZN => n16279);
   U19398 : NAND2_X1 port map( A1 => n25154, A2 => n8926, ZN => n25140);
   U19400 : OAI21_X1 port map( A1 => n16273, A2 => n8207, B => n8925, ZN => 
                           n25160);
   U19402 : INV_X2 port map( I => n8933, ZN => n12168);
   U19403 : NAND2_X1 port map( A1 => n5966, A2 => n12168, ZN => n8934);
   U19406 : NOR2_X1 port map( A1 => n8944, A2 => n32193, ZN => n22529);
   U19408 : INV_X2 port map( I => n9626, ZN => n21452);
   U19414 : NAND2_X2 port map( A1 => n14773, A2 => n14772, ZN => n22871);
   U19416 : XOR2_X1 port map( A1 => n15114, A2 => n1197, Z => n8974);
   U19417 : XOR2_X1 port map( A1 => n8976, A2 => n13190, Z => n8975);
   U19418 : XOR2_X1 port map( A1 => n23503, A2 => n28927, Z => n8976);
   U19421 : XOR2_X1 port map( A1 => n21964, A2 => n1065, Z => n8992);
   U19424 : XOR2_X1 port map( A1 => n22036, A2 => n17723, Z => n9000);
   U19425 : INV_X1 port map( I => n20515, ZN => n20174);
   U19426 : XOR2_X1 port map( A1 => n9005, A2 => n9004, Z => n11051);
   U19429 : INV_X2 port map( I => n11051, ZN => n15110);
   U19432 : XOR2_X1 port map( A1 => n23419, A2 => n24861, Z => n9011);
   U19433 : XOR2_X1 port map( A1 => n23359, A2 => n15897, Z => n9013);
   U19435 : XOR2_X1 port map( A1 => n11836, A2 => n9021, Z => n9020);
   U19436 : XOR2_X1 port map( A1 => n11897, A2 => n16301, Z => n9021);
   U19443 : XOR2_X1 port map( A1 => n8347, A2 => n14557, Z => n9038);
   U19445 : NAND2_X1 port map( A1 => n936, A2 => n26566, ZN => n20313);
   U19446 : MUX2_X1 port map( I0 => n20578, I1 => n20579, S => n8528, Z => 
                           n20585);
   U19447 : XOR2_X1 port map( A1 => n19719, A2 => n9045, Z => n9044);
   U19448 : XOR2_X1 port map( A1 => n19763, A2 => n25104, Z => n9045);
   U19452 : INV_X2 port map( I => n9064, ZN => n12952);
   U19454 : NAND2_X1 port map( A1 => n24308, A2 => n11041, ZN => n12575);
   U19458 : XOR2_X1 port map( A1 => n9907, A2 => n24953, Z => n9087);
   U19459 : XOR2_X1 port map( A1 => n16237, A2 => n25319, Z => n12084);
   U19460 : XOR2_X1 port map( A1 => n22114, A2 => n1307, Z => n22115);
   U19463 : XOR2_X1 port map( A1 => n19616, A2 => n18902, Z => n18903);
   U19465 : XOR2_X1 port map( A1 => n13586, A2 => n16672, Z => n9092);
   U19467 : NAND2_X1 port map( A1 => n19997, A2 => n19986, ZN => n9098);
   U19469 : XOR2_X1 port map( A1 => n19641, A2 => n25224, Z => n9101);
   U19470 : XOR2_X1 port map( A1 => n19686, A2 => n15117, Z => n9102);
   U19476 : XOR2_X1 port map( A1 => n16351, A2 => n19787, Z => n9116);
   U19479 : XNOR2_X1 port map( A1 => Plaintext(114), A2 => Key(114), ZN => 
                           n9118);
   U19487 : XOR2_X1 port map( A1 => n343, A2 => n22173, Z => n21961);
   U19492 : AOI22_X1 port map( A1 => n19336, A2 => n12815, B1 => n12316, B2 => 
                           n16699, ZN => n9134);
   U19495 : XOR2_X1 port map( A1 => n21926, A2 => n13303, Z => n9136);
   U19496 : XOR2_X1 port map( A1 => n19530, A2 => n32981, Z => n9138);
   U19497 : XOR2_X1 port map( A1 => n9141, A2 => n16402, Z => n13856);
   U19499 : NOR2_X1 port map( A1 => n31969, A2 => n27600, ZN => n20359);
   U19500 : NAND2_X1 port map( A1 => n10312, A2 => n31969, ZN => n20239);
   U19501 : NAND2_X1 port map( A1 => n19865, A2 => n31969, ZN => n13246);
   U19502 : XOR2_X1 port map( A1 => n23206, A2 => n23207, Z => n9154);
   U19509 : AOI21_X2 port map( A1 => n11470, A2 => n9174, B => n18651, ZN => 
                           n11085);
   U19513 : NAND2_X1 port map( A1 => n11754, A2 => n31155, ZN => n16090);
   U19514 : NAND2_X1 port map( A1 => n1238, A2 => n24118, ZN => n9178);
   U19515 : INV_X1 port map( I => n25818, ZN => n25822);
   U19517 : NOR2_X1 port map( A1 => n9182, A2 => n9181, ZN => n9180);
   U19518 : NAND2_X2 port map( A1 => n18491, A2 => n9183, ZN => n18990);
   U19520 : XOR2_X1 port map( A1 => n9185, A2 => n16390, Z => n12580);
   U19521 : INV_X2 port map( I => n19255, ZN => n19256);
   U19531 : NAND2_X1 port map( A1 => n12143, A2 => n9219, ZN => n12430);
   U19533 : XOR2_X1 port map( A1 => n26562, A2 => n32881, Z => n14902);
   U19536 : XOR2_X1 port map( A1 => n9231, A2 => n9988, Z => n9230);
   U19538 : OAI21_X1 port map( A1 => n14503, A2 => n21662, B => n32898, ZN => 
                           n13803);
   U19543 : INV_X2 port map( I => n9239, ZN => n11944);
   U19545 : XOR2_X1 port map( A1 => n16693, A2 => n15147, Z => n9241);
   U19547 : NAND2_X1 port map( A1 => n830, A2 => n4770, ZN => n9249);
   U19549 : NOR2_X2 port map( A1 => n9014, A2 => n14005, ZN => n9255);
   U19553 : XOR2_X1 port map( A1 => n16586, A2 => n4975, Z => n19522);
   U19555 : XOR2_X1 port map( A1 => n24787, A2 => n25131, Z => n9281);
   U19557 : NAND2_X2 port map( A1 => n14161, A2 => n14005, ZN => n20219);
   U19560 : XOR2_X1 port map( A1 => n9290, A2 => n22099, Z => n22165);
   U19561 : INV_X1 port map( I => n8386, ZN => n9305);
   U19566 : INV_X1 port map( I => n10325, ZN => n9296);
   U19568 : XOR2_X1 port map( A1 => n26931, A2 => n22273, Z => n9298);
   U19574 : NAND2_X1 port map( A1 => n11264, A2 => n9302, ZN => n19882);
   U19576 : XOR2_X1 port map( A1 => n9303, A2 => n16662, Z => n10557);
   U19577 : XOR2_X1 port map( A1 => n9303, A2 => n1343, Z => n20702);
   U19578 : XOR2_X1 port map( A1 => n9308, A2 => n7603, Z => n9307);
   U19579 : XOR2_X1 port map( A1 => n9309, A2 => n9310, Z => n11238);
   U19580 : XOR2_X1 port map( A1 => n9311, A2 => n22310, Z => n9309);
   U19581 : XOR2_X1 port map( A1 => n16971, A2 => n21887, Z => n9310);
   U19584 : XOR2_X1 port map( A1 => n19464, A2 => n11361, Z => n9325);
   U19588 : AND3_X1 port map( A1 => n23950, A2 => n10187, A3 => n33659, Z => 
                           n9345);
   U19589 : XOR2_X1 port map( A1 => n23234, A2 => n9349, Z => n9347);
   U19591 : XOR2_X1 port map( A1 => n23438, A2 => n30557, Z => n9349);
   U19595 : XOR2_X1 port map( A1 => n14211, A2 => n9362, Z => n9361);
   U19596 : XOR2_X1 port map( A1 => n19682, A2 => n16680, Z => n9362);
   U19607 : AOI21_X2 port map( A1 => n13112, A2 => n13111, B => n13110, ZN => 
                           n19283);
   U19609 : XOR2_X1 port map( A1 => n24441, A2 => n24505, Z => n9385);
   U19610 : NAND3_X2 port map( A1 => n24278, A2 => n14288, A3 => n24279, ZN => 
                           n24475);
   U19611 : XOR2_X1 port map( A1 => n21949, A2 => n9388, Z => n9387);
   U19612 : XOR2_X1 port map( A1 => n22033, A2 => n25669, Z => n9388);
   U19616 : XOR2_X1 port map( A1 => n16838, A2 => n544, Z => n11995);
   U19619 : XOR2_X1 port map( A1 => n9412, A2 => n17679, Z => n21949);
   U19620 : XOR2_X1 port map( A1 => n9412, A2 => n25751, Z => n22142);
   U19625 : XOR2_X1 port map( A1 => Plaintext(132), A2 => Key(132), Z => n9437)
                           ;
   U19628 : INV_X2 port map( I => n9920, ZN => n23862);
   U19633 : INV_X2 port map( I => n9437, ZN => n18537);
   U19639 : NAND2_X1 port map( A1 => n9446, A2 => n22946, ZN => n16921);
   U19640 : XOR2_X1 port map( A1 => n22182, A2 => n9447, Z => n16617);
   U19641 : XOR2_X1 port map( A1 => n9960, A2 => n27281, Z => n9447);
   U19657 : XOR2_X1 port map( A1 => n11751, A2 => n1403, Z => n9475);
   U19662 : INV_X2 port map( I => n9486, ZN => n25763);
   U19663 : XOR2_X1 port map( A1 => n16838, A2 => n9488, Z => n9487);
   U19664 : XOR2_X1 port map( A1 => n24533, A2 => n27157, Z => n9488);
   U19668 : NAND2_X2 port map( A1 => n21089, A2 => n21090, ZN => n21687);
   U19670 : XOR2_X1 port map( A1 => n9504, A2 => n27137, Z => n9503);
   U19671 : XOR2_X1 port map( A1 => n18453, A2 => n25881, Z => n9504);
   U19672 : XOR2_X1 port map( A1 => n1305, A2 => n27180, Z => n9505);
   U19673 : XOR2_X1 port map( A1 => n20736, A2 => n20996, Z => n20738);
   U19674 : XOR2_X1 port map( A1 => n9507, A2 => n20542, Z => n10788);
   U19675 : NOR2_X1 port map( A1 => n13548, A2 => n13514, ZN => n9513);
   U19678 : XOR2_X1 port map( A1 => n29312, A2 => n9527, Z => n9526);
   U19680 : XOR2_X1 port map( A1 => n9533, A2 => n9529, Z => n9535);
   U19681 : XOR2_X1 port map( A1 => n9532, A2 => n9530, Z => n9529);
   U19682 : XOR2_X1 port map( A1 => n22210, A2 => n9531, Z => n9530);
   U19685 : NAND2_X2 port map( A1 => n9540, A2 => n9539, ZN => n19335);
   U19687 : AOI21_X1 port map( A1 => n33594, A2 => n22641, B => n22645, ZN => 
                           n9544);
   U19690 : XOR2_X1 port map( A1 => n23397, A2 => n9551, Z => n9550);
   U19691 : XOR2_X1 port map( A1 => n15183, A2 => n25693, Z => n9551);
   U19692 : INV_X2 port map( I => n9564, ZN => n11957);
   U19694 : XOR2_X1 port map( A1 => n27015, A2 => n9568, Z => n9567);
   U19696 : XOR2_X1 port map( A1 => n9209, A2 => n24809, Z => n9573);
   U19697 : XOR2_X1 port map( A1 => n24808, A2 => n10583, Z => n9574);
   U19705 : XOR2_X1 port map( A1 => n29718, A2 => n1192, Z => n9599);
   U19709 : XOR2_X1 port map( A1 => n9606, A2 => n9604, Z => n17218);
   U19710 : XOR2_X1 port map( A1 => n27375, A2 => n9605, Z => n9604);
   U19711 : NOR2_X1 port map( A1 => n9612, A2 => n25235, ZN => n9609);
   U19715 : NAND2_X1 port map( A1 => n22414, A2 => n9617, ZN => n15581);
   U19716 : XOR2_X1 port map( A1 => n9623, A2 => n9621, Z => n22394);
   U19717 : XOR2_X1 port map( A1 => n9622, A2 => n21967, Z => n9621);
   U19718 : XOR2_X1 port map( A1 => n31457, A2 => n13651, Z => n9622);
   U19719 : XOR2_X1 port map( A1 => n22183, A2 => n14994, Z => n9623);
   U19721 : XOR2_X1 port map( A1 => n10169, A2 => n453, Z => n9634);
   U19726 : INV_X2 port map( I => n9640, ZN => n19998);
   U19727 : XOR2_X1 port map( A1 => n19168, A2 => n18915, Z => n9641);
   U19729 : NAND2_X1 port map( A1 => n25193, A2 => n27149, ZN => n13266);
   U19730 : AOI21_X1 port map( A1 => n830, A2 => n25194, B => n27149, ZN => 
                           n9675);
   U19733 : XOR2_X1 port map( A1 => n6484, A2 => n25156, Z => n9650);
   U19736 : AND2_X1 port map( A1 => n3148, A2 => n23995, Z => n9658);
   U19737 : NAND3_X1 port map( A1 => n31960, A2 => n7182, A3 => n27954, ZN => 
                           n9896);
   U19740 : XOR2_X1 port map( A1 => n9665, A2 => n16472, Z => n10986);
   U19743 : XOR2_X1 port map( A1 => n13777, A2 => n23232, Z => n9672);
   U19745 : NOR2_X1 port map( A1 => n25985, A2 => n9677, ZN => n10853);
   U19747 : XOR2_X1 port map( A1 => n11860, A2 => n21582, Z => n9679);
   U19749 : NOR2_X1 port map( A1 => n1358, A2 => n13327, ZN => n11013);
   U19750 : NOR2_X1 port map( A1 => n29338, A2 => n1358, ZN => n14693);
   U19753 : AOI22_X1 port map( A1 => n9696, A2 => n29085, B1 => n27123, B2 => 
                           n9247, ZN => n9695);
   U19754 : NAND3_X1 port map( A1 => n13266, A2 => n4781, A3 => n9698, ZN => 
                           n9697);
   U19755 : NAND2_X1 port map( A1 => n10858, A2 => n4953, ZN => n9698);
   U19759 : NAND2_X1 port map( A1 => n13245, A2 => n9703, ZN => n9705);
   U19760 : NAND3_X1 port map( A1 => n29085, A2 => n786, A3 => n9247, ZN => 
                           n9704);
   U19761 : XOR2_X1 port map( A1 => n646, A2 => n27171, Z => n14818);
   U19762 : XOR2_X1 port map( A1 => n12821, A2 => n646, Z => n23075);
   U19763 : XOR2_X1 port map( A1 => n1262, A2 => n646, Z => n23469);
   U19765 : INV_X1 port map( I => n14179, ZN => n15661);
   U19767 : NOR2_X1 port map( A1 => n9729, A2 => n18711, ZN => n13566);
   U19768 : NOR2_X1 port map( A1 => n1835, A2 => n9729, ZN => n18317);
   U19773 : OAI21_X1 port map( A1 => n22807, A2 => n3614, B => n851, ZN => 
                           n22809);
   U19774 : NAND2_X1 port map( A1 => n15457, A2 => n3614, ZN => n12782);
   U19775 : NAND2_X1 port map( A1 => n22403, A2 => n22678, ZN => n9739);
   U19779 : XOR2_X1 port map( A1 => n22158, A2 => n22205, Z => n10626);
   U19783 : XOR2_X1 port map( A1 => n22137, A2 => n11863, Z => n9758);
   U19789 : XOR2_X1 port map( A1 => n11897, A2 => n16698, Z => n9764);
   U19791 : XOR2_X1 port map( A1 => n32660, A2 => n24923, Z => n24578);
   U19792 : XOR2_X1 port map( A1 => n32660, A2 => n15653, Z => n24453);
   U19793 : XOR2_X1 port map( A1 => Plaintext(23), A2 => Key(23), Z => n9930);
   U19795 : NOR2_X1 port map( A1 => n11943, A2 => n16320, ZN => n9768);
   U19799 : XOR2_X1 port map( A1 => n9782, A2 => n9780, Z => n9798);
   U19800 : XOR2_X1 port map( A1 => n9781, A2 => n15963, Z => n9780);
   U19801 : XOR2_X1 port map( A1 => n23450, A2 => n16160, Z => n9781);
   U19803 : NOR2_X2 port map( A1 => n13384, A2 => n14552, ZN => n23196);
   U19808 : NOR2_X1 port map( A1 => n28581, A2 => n9793, ZN => n11658);
   U19810 : OAI22_X1 port map( A1 => n9811, A2 => n8886, B1 => n21585, B2 => 
                           n9793, ZN => n10825);
   U19811 : NAND2_X1 port map( A1 => n12095, A2 => n9793, ZN => n11656);
   U19813 : NOR2_X1 port map( A1 => n953, A2 => n4868, ZN => n18573);
   U19817 : XOR2_X1 port map( A1 => n9819, A2 => n9820, Z => n9818);
   U19818 : XOR2_X1 port map( A1 => n32286, A2 => n19703, Z => n9820);
   U19819 : XOR2_X1 port map( A1 => n19426, A2 => n16381, Z => n9822);
   U19826 : XOR2_X1 port map( A1 => n9843, A2 => n17986, Z => n23248);
   U19827 : NAND2_X1 port map( A1 => n9847, A2 => n9846, ZN => n9933);
   U19830 : NAND2_X1 port map( A1 => n31155, A2 => n24117, ZN => n10118);
   U19831 : NAND2_X1 port map( A1 => n1238, A2 => n24225, ZN => n12068);
   U19834 : XOR2_X1 port map( A1 => n20727, A2 => n1428, Z => n13339);
   U19838 : XOR2_X1 port map( A1 => n9863, A2 => n23242, Z => n23447);
   U19841 : XOR2_X1 port map( A1 => n23255, A2 => n9867, Z => n9866);
   U19853 : INV_X2 port map( I => n14676, ZN => n15089);
   U19856 : NOR2_X1 port map( A1 => n16908, A2 => n12144, ZN => n16907);
   U19859 : OR2_X1 port map( A1 => n20556, A2 => n20236, Z => n20170);
   U19865 : XOR2_X1 port map( A1 => n11304, A2 => n9878, Z => n9877);
   U19866 : XOR2_X1 port map( A1 => n16708, A2 => n25038, Z => n9878);
   U19869 : XOR2_X1 port map( A1 => n24846, A2 => n25772, Z => n17296);
   U19872 : INV_X2 port map( I => n11413, ZN => n11676);
   U19874 : XOR2_X1 port map( A1 => n9904, A2 => n19513, Z => n19514);
   U19878 : XOR2_X1 port map( A1 => n9907, A2 => n11370, Z => n24546);
   U19887 : XOR2_X1 port map( A1 => n16081, A2 => n24374, Z => n9928);
   U19888 : INV_X2 port map( I => n9929, ZN => n19857);
   U19890 : NAND3_X1 port map( A1 => n25867, A2 => n700, A3 => n10062, ZN => 
                           n11253);
   U19902 : NOR2_X2 port map( A1 => n13071, A2 => n13070, ZN => n9951);
   U19903 : XOR2_X1 port map( A1 => n30943, A2 => n19479, Z => n9955);
   U19906 : XOR2_X1 port map( A1 => n356, A2 => n25054, Z => n12918);
   U19907 : XOR2_X1 port map( A1 => n24750, A2 => n356, Z => n13824);
   U19909 : INV_X2 port map( I => n9968, ZN => n11898);
   U19910 : XOR2_X1 port map( A1 => n9969, A2 => n13438, Z => Ciphertext(2));
   U19913 : INV_X1 port map( I => n19322, ZN => n19324);
   U19916 : OAI21_X2 port map( A1 => n29282, A2 => n14004, B => n9978, ZN => 
                           n20630);
   U19918 : OAI21_X1 port map( A1 => n25613, A2 => n9982, B => n9981, ZN => 
                           n10265);
   U19920 : XOR2_X1 port map( A1 => n15275, A2 => n20996, Z => n9984);
   U19921 : INV_X1 port map( I => n20479, ZN => n9985);
   U19923 : XOR2_X1 port map( A1 => n17040, A2 => n13388, Z => n9993);
   U19924 : NOR2_X1 port map( A1 => n21825, A2 => n9994, ZN => n21829);
   U19926 : NAND2_X1 port map( A1 => n30878, A2 => n28288, ZN => n10764);
   U19930 : NAND3_X1 port map( A1 => n10011, A2 => n10385, A3 => n16520, ZN => 
                           n10010);
   U19936 : XOR2_X1 port map( A1 => Plaintext(148), A2 => Key(148), Z => n15519
                           );
   U19939 : INV_X1 port map( I => Plaintext(83), ZN => n10044);
   U19940 : XOR2_X1 port map( A1 => n10044, A2 => Key(83), Z => n18575);
   U19943 : AOI21_X2 port map( A1 => n12837, A2 => n14537, B => n10055, ZN => 
                           n19108);
   U19946 : INV_X2 port map( I => n10058, ZN => n13514);
   U19947 : XOR2_X1 port map( A1 => Plaintext(35), A2 => Key(35), Z => n13531);
   U19951 : AOI21_X1 port map( A1 => n17489, A2 => n14108, B => n10062, ZN => 
                           n17488);
   U19952 : XOR2_X1 port map( A1 => n770, A2 => n16263, Z => n10064);
   U19957 : INV_X2 port map( I => n21228, ZN => n21443);
   U19959 : XOR2_X1 port map( A1 => n19517, A2 => n26005, Z => n10077);
   U19961 : NAND2_X1 port map( A1 => n23868, A2 => n844, ZN => n12603);
   U19963 : XOR2_X1 port map( A1 => n10082, A2 => n1405, Z => Ciphertext(160));
   U19965 : XOR2_X1 port map( A1 => n10084, A2 => n32814, Z => n24698);
   U19967 : XOR2_X1 port map( A1 => n10088, A2 => n10090, Z => n25710);
   U19968 : XOR2_X1 port map( A1 => n24597, A2 => n10089, Z => n10088);
   U19969 : XOR2_X1 port map( A1 => n24556, A2 => n24382, Z => n10090);
   U19972 : NAND2_X1 port map( A1 => n11046, A2 => n10097, ZN => n24864);
   U19973 : INV_X1 port map( I => n10099, ZN => n10098);
   U19975 : NAND2_X2 port map( A1 => n20316, A2 => n20315, ZN => n20872);
   U19977 : XOR2_X1 port map( A1 => n15710, A2 => n23453, Z => n23180);
   U19978 : NOR2_X1 port map( A1 => n28344, A2 => n18349, ZN => n12013);
   U19979 : XNOR2_X1 port map( A1 => Plaintext(40), A2 => Key(40), ZN => n10114
                           );
   U19980 : NOR2_X1 port map( A1 => n24225, A2 => n24118, ZN => n10119);
   U19983 : XOR2_X1 port map( A1 => n32791, A2 => n24917, Z => n10122);
   U19985 : XOR2_X1 port map( A1 => n19634, A2 => n24623, Z => n10123);
   U19986 : INV_X2 port map( I => n17820, ZN => n19290);
   U19987 : XOR2_X1 port map( A1 => n10130, A2 => n13517, Z => n10129);
   U19992 : INV_X2 port map( I => n657, ZN => n23868);
   U19993 : NOR2_X1 port map( A1 => n29246, A2 => n10145, ZN => n10542);
   U19995 : XOR2_X1 port map( A1 => n23521, A2 => n12122, Z => n10150);
   U19999 : XOR2_X1 port map( A1 => n22198, A2 => n25054, Z => n10155);
   U20000 : OAI21_X2 port map( A1 => n21607, A2 => n21776, B => n18163, ZN => 
                           n22198);
   U20002 : XOR2_X1 port map( A1 => n10157, A2 => n25735, Z => Ciphertext(158))
                           ;
   U20004 : XOR2_X1 port map( A1 => n20819, A2 => n10159, Z => n15338);
   U20008 : XOR2_X1 port map( A1 => n27180, A2 => n25570, Z => n10165);
   U20009 : INV_X2 port map( I => n10171, ZN => n25628);
   U20012 : XOR2_X1 port map( A1 => n22157, A2 => n16237, Z => n10370);
   U20013 : NAND3_X1 port map( A1 => n11931, A2 => n27262, A3 => n10174, ZN => 
                           n10268);
   U20017 : XOR2_X1 port map( A1 => n19341, A2 => n25009, Z => n10180);
   U20018 : NOR2_X1 port map( A1 => n10182, A2 => n10181, ZN => n18590);
   U20021 : XOR2_X1 port map( A1 => n21924, A2 => n21577, Z => n10184);
   U20027 : XOR2_X1 port map( A1 => n24428, A2 => n10195, Z => n10194);
   U20029 : NAND2_X2 port map( A1 => n17118, A2 => n24610, ZN => n10199);
   U20031 : XOR2_X1 port map( A1 => n9706, A2 => n24895, Z => n20712);
   U20032 : XOR2_X1 port map( A1 => n10201, A2 => n16657, Z => n14656);
   U20033 : AND2_X1 port map( A1 => n629, A2 => n10206, Z => n10908);
   U20034 : AOI21_X2 port map( A1 => n10208, A2 => n18403, B => n10207, ZN => 
                           n16354);
   U20035 : INV_X2 port map( I => n10209, ZN => n18219);
   U20036 : OAI21_X1 port map( A1 => n4289, A2 => n816, B => n20570, ZN => 
                           n20573);
   U20041 : XOR2_X1 port map( A1 => n29320, A2 => n11603, Z => n10237);
   U20042 : XOR2_X1 port map( A1 => n29320, A2 => n25728, Z => n24443);
   U20043 : XOR2_X1 port map( A1 => n29320, A2 => n24507, Z => n24508);
   U20044 : AOI21_X1 port map( A1 => n824, A2 => n10227, B => n13568, ZN => 
                           n17981);
   U20052 : XOR2_X1 port map( A1 => n10087, A2 => n13075, Z => n10249);
   U20053 : NOR2_X1 port map( A1 => n974, A2 => n10281, ZN => n24131);
   U20054 : NAND2_X1 port map( A1 => n2575, A2 => n10254, ZN => n14870);
   U20058 : XOR2_X1 port map( A1 => n19710, A2 => n25086, Z => n10262);
   U20059 : NAND3_X1 port map( A1 => n29659, A2 => n28010, A3 => n15519, ZN => 
                           n18438);
   U20060 : OAI22_X1 port map( A1 => n10843, A2 => n29659, B1 => n17321, B2 => 
                           n959, ZN => n10842);
   U20062 : XOR2_X1 port map( A1 => n22079, A2 => n10270, Z => n22082);
   U20063 : XOR2_X1 port map( A1 => n32881, A2 => n2353, Z => n10270);
   U20068 : XOR2_X1 port map( A1 => n24624, A2 => n11699, Z => n10276);
   U20069 : XOR2_X1 port map( A1 => n22014, A2 => n1392, Z => n10278);
   U20071 : XNOR2_X1 port map( A1 => Plaintext(180), A2 => Key(180), ZN => 
                           n10284);
   U20072 : INV_X2 port map( I => n10287, ZN => n10533);
   U20077 : NAND2_X1 port map( A1 => n12487, A2 => n10301, ZN => n12486);
   U20078 : OAI22_X1 port map( A1 => n16836, A2 => n14954, B1 => n28658, B2 => 
                           n10301, ZN => n12302);
   U20079 : NOR2_X1 port map( A1 => n1322, A2 => n21832, ZN => n21835);
   U20080 : XOR2_X1 port map( A1 => n12828, A2 => n10304, Z => n16332);
   U20081 : XOR2_X1 port map( A1 => n22300, A2 => n12084, Z => n10304);
   U20082 : XOR2_X1 port map( A1 => n23368, A2 => n10308, Z => n23127);
   U20083 : MUX2_X1 port map( I0 => n20360, I1 => n27600, S => n29553, Z => 
                           n20240);
   U20088 : XOR2_X1 port map( A1 => n572, A2 => n14916, Z => n10320);
   U20092 : NOR2_X1 port map( A1 => n30558, A2 => n10325, ZN => n18885);
   U20094 : XOR2_X1 port map( A1 => n8356, A2 => n24964, Z => n10328);
   U20096 : XOR2_X1 port map( A1 => n27801, A2 => n27950, Z => n24445);
   U20101 : XOR2_X1 port map( A1 => n9145, A2 => n14727, Z => n15588);
   U20103 : XOR2_X1 port map( A1 => n15293, A2 => n15408, Z => n10347);
   U20104 : INV_X2 port map( I => n10350, ZN => n15318);
   U20105 : OR2_X1 port map( A1 => n12691, A2 => n11608, Z => n10358);
   U20118 : XOR2_X1 port map( A1 => n30571, A2 => n16634, Z => n21457);
   U20119 : XOR2_X1 port map( A1 => n156, A2 => n1194, Z => n10399);
   U20121 : XOR2_X1 port map( A1 => n33219, A2 => n25213, Z => n10412);
   U20123 : AND2_X1 port map( A1 => n11346, A2 => n1775, Z => n10416);
   U20127 : XOR2_X1 port map( A1 => n22284, A2 => n22283, Z => n10421);
   U20129 : INV_X2 port map( I => n10426, ZN => n19724);
   U20130 : INV_X2 port map( I => n10430, ZN => n11900);
   U20132 : XOR2_X1 port map( A1 => n25993, A2 => n1431, Z => n10434);
   U20134 : NAND2_X1 port map( A1 => n17368, A2 => n14213, ZN => n10485);
   U20135 : NAND2_X1 port map( A1 => n12877, A2 => n14213, ZN => n12533);
   U20136 : OAI21_X1 port map( A1 => n16443, A2 => n26158, B => n10449, ZN => 
                           n10448);
   U20139 : XOR2_X1 port map( A1 => n848, A2 => n29155, Z => n10459);
   U20141 : XOR2_X1 port map( A1 => n11762, A2 => n22083, Z => n10461);
   U20147 : XOR2_X1 port map( A1 => n19731, A2 => n10467, Z => n10466);
   U20148 : XOR2_X1 port map( A1 => n19375, A2 => n1369, Z => n10467);
   U20150 : NOR2_X1 port map( A1 => n5455, A2 => n7492, ZN => n12144);
   U20153 : XOR2_X1 port map( A1 => n12414, A2 => n1198, Z => n10474);
   U20157 : NOR2_X2 port map( A1 => n10491, A2 => n10490, ZN => n22130);
   U20161 : INV_X2 port map( I => n10505, ZN => n21398);
   U20163 : XOR2_X1 port map( A1 => n20893, A2 => n10508, Z => n10507);
   U20164 : XOR2_X1 port map( A1 => n20970, A2 => n1338, Z => n10508);
   U20165 : INV_X2 port map( I => n10514, ZN => n19991);
   U20167 : XOR2_X1 port map( A1 => n24429, A2 => n15473, Z => n10515);
   U20168 : XOR2_X1 port map( A1 => n30795, A2 => n7879, Z => n24429);
   U20169 : XOR2_X1 port map( A1 => n10585, A2 => n15815, Z => n10516);
   U20173 : XOR2_X1 port map( A1 => n10525, A2 => n22712, Z => n15116);
   U20177 : NOR2_X1 port map( A1 => n71, A2 => n20103, ZN => n16980);
   U20178 : NAND2_X1 port map( A1 => n15551, A2 => n71, ZN => n20105);
   U20179 : XOR2_X1 port map( A1 => n10539, A2 => n13419, Z => n24529);
   U20180 : XOR2_X1 port map( A1 => n24635, A2 => n10539, Z => n16394);
   U20182 : OAI21_X2 port map( A1 => n10548, A2 => n10756, B => n10547, ZN => 
                           n10755);
   U20185 : XOR2_X1 port map( A1 => n29312, A2 => n10553, Z => n10552);
   U20189 : INV_X2 port map( I => n16881, ZN => n16948);
   U20190 : NAND2_X2 port map( A1 => n11247, A2 => n10566, ZN => n24970);
   U20191 : NAND2_X1 port map( A1 => n18035, A2 => n12323, ZN => n10571);
   U20193 : NAND2_X1 port map( A1 => n20580, A2 => n26566, ZN => n20584);
   U20195 : XOR2_X1 port map( A1 => n32399, A2 => n16685, Z => n10581);
   U20197 : XOR2_X1 port map( A1 => n2864, A2 => n10584, Z => n10583);
   U20198 : XOR2_X1 port map( A1 => n10587, A2 => n16533, Z => Ciphertext(69));
   U20200 : AND2_X1 port map( A1 => n30234, A2 => n8365, Z => n10589);
   U20205 : NOR2_X1 port map( A1 => n24590, A2 => n30018, ZN => n10600);
   U20206 : INV_X1 port map( I => n24590, ZN => n10603);
   U20207 : NOR2_X1 port map( A1 => n10606, A2 => n10605, ZN => n10604);
   U20213 : XOR2_X1 port map( A1 => n22056, A2 => n17679, Z => n22268);
   U20215 : XOR2_X1 port map( A1 => n11694, A2 => n1309, Z => n11884);
   U20216 : XOR2_X1 port map( A1 => n31105, A2 => n9960, Z => n21879);
   U20217 : XOR2_X1 port map( A1 => n7828, A2 => n15775, Z => n10616);
   U20220 : XOR2_X1 port map( A1 => n10626, A2 => n13956, Z => n11600);
   U20225 : XOR2_X1 port map( A1 => n16076, A2 => n10773, Z => n17915);
   U20227 : XOR2_X1 port map( A1 => n9536, A2 => n10650, Z => n10649);
   U20229 : NOR2_X1 port map( A1 => n13509, A2 => n7007, ZN => n10658);
   U20231 : NAND2_X1 port map( A1 => n21424, A2 => n6855, ZN => n15564);
   U20232 : NOR2_X1 port map( A1 => n30854, A2 => n21424, ZN => n21337);
   U20233 : OAI21_X1 port map( A1 => n21243, A2 => n30854, B => n11912, ZN => 
                           n17803);
   U20234 : MUX2_X1 port map( I0 => n20071, I1 => n31080, S => n729, Z => 
                           n20072);
   U20235 : XOR2_X1 port map( A1 => n19666, A2 => n10662, Z => n10661);
   U20236 : XOR2_X1 port map( A1 => n29312, A2 => n1193, Z => n10662);
   U20239 : NAND2_X1 port map( A1 => n18747, A2 => n10665, ZN => n17874);
   U20240 : NAND2_X1 port map( A1 => n16487, A2 => n10665, ZN => n14706);
   U20241 : NOR2_X1 port map( A1 => n12575, A2 => n12574, ZN => n10666);
   U20244 : XOR2_X1 port map( A1 => n22211, A2 => n22226, Z => n22242);
   U20245 : XNOR2_X1 port map( A1 => n10675, A2 => n10674, ZN => n10673);
   U20263 : XOR2_X1 port map( A1 => n10704, A2 => n10701, Z => n10725);
   U20264 : XOR2_X1 port map( A1 => n10703, A2 => n10702, Z => n10701);
   U20265 : XOR2_X1 port map( A1 => n17362, A2 => n25038, Z => n10702);
   U20272 : OAI21_X2 port map( A1 => n6303, A2 => n14955, B => n10721, ZN => 
                           n12561);
   U20273 : XOR2_X1 port map( A1 => n17213, A2 => n15708, Z => n10722);
   U20274 : XOR2_X1 port map( A1 => n19586, A2 => n461, Z => n10723);
   U20275 : XOR2_X1 port map( A1 => n10727, A2 => n17205, Z => n17203);
   U20276 : XOR2_X1 port map( A1 => n10728, A2 => n34160, Z => n10727);
   U20277 : XOR2_X1 port map( A1 => n17697, A2 => n1429, Z => n10728);
   U20284 : XOR2_X1 port map( A1 => n20857, A2 => n20905, Z => n10737);
   U20285 : XOR2_X1 port map( A1 => n19626, A2 => n19708, Z => n10738);
   U20288 : NOR2_X1 port map( A1 => n17110, A2 => n25292, ZN => n10744);
   U20289 : NOR2_X1 port map( A1 => n10748, A2 => n17110, ZN => n10747);
   U20291 : AOI22_X2 port map( A1 => n10763, A2 => n23850, B1 => n14664, B2 => 
                           n10762, ZN => n24299);
   U20302 : XOR2_X1 port map( A1 => n2353, A2 => n22248, Z => n17219);
   U20303 : NOR2_X2 port map( A1 => n11493, A2 => n19953, ZN => n11984);
   U20307 : XOR2_X1 port map( A1 => n10800, A2 => n10797, Z => n17144);
   U20308 : XOR2_X1 port map( A1 => n10799, A2 => n10798, Z => n10797);
   U20309 : XOR2_X1 port map( A1 => n20848, A2 => n16679, Z => n10798);
   U20313 : XOR2_X1 port map( A1 => n10810, A2 => n19591, Z => n10809);
   U20315 : XOR2_X1 port map( A1 => n28848, A2 => n25191, Z => n10814);
   U20316 : AND2_X1 port map( A1 => n25066, A2 => n10822, Z => n10821);
   U20322 : NOR2_X1 port map( A1 => n13304, A2 => n18048, ZN => n21387);
   U20335 : XOR2_X1 port map( A1 => n19763, A2 => n17091, Z => n10866);
   U20337 : XOR2_X1 port map( A1 => n10873, A2 => n14979, Z => n10872);
   U20341 : XOR2_X1 port map( A1 => n20916, A2 => n10878, Z => n10877);
   U20344 : XOR2_X1 port map( A1 => n2353, A2 => n24953, Z => n10887);
   U20345 : XOR2_X1 port map( A1 => n10889, A2 => n18190, Z => n10888);
   U20346 : XOR2_X1 port map( A1 => n30212, A2 => n25801, Z => n19340);
   U20347 : NAND3_X1 port map( A1 => n20569, A2 => n29069, A3 => n4289, ZN => 
                           n11761);
   U20351 : INV_X2 port map( I => n10900, ZN => n16442);
   U20353 : NAND2_X2 port map( A1 => n10910, A2 => n10909, ZN => n19199);
   U20354 : XOR2_X1 port map( A1 => n10915, A2 => n15029, Z => n10914);
   U20356 : XOR2_X1 port map( A1 => n15031, A2 => n4400, Z => n10917);
   U20357 : INV_X1 port map( I => n24004, ZN => n13984);
   U20358 : NAND2_X1 port map( A1 => n31096, A2 => n24004, ZN => n14889);
   U20361 : INV_X2 port map( I => n10932, ZN => n16633);
   U20362 : INV_X2 port map( I => n10936, ZN => n16534);
   U20364 : XOR2_X1 port map( A1 => n10945, A2 => n10944, Z => n25308);
   U20366 : XOR2_X1 port map( A1 => n10946, A2 => n24895, Z => n12779);
   U20367 : XOR2_X1 port map( A1 => n10946, A2 => n22056, Z => n21948);
   U20369 : OAI22_X2 port map( A1 => n17581, A2 => n3219, B1 => n15086, B2 => 
                           n15085, ZN => n24636);
   U20373 : MUX2_X1 port map( I0 => n802, I1 => n22766, S => n9293, Z => n22767
                           );
   U20379 : XOR2_X1 port map( A1 => n12614, A2 => n10961, Z => n10960);
   U20380 : XOR2_X1 port map( A1 => n14952, A2 => n960, Z => n10961);
   U20385 : XOR2_X1 port map( A1 => n10979, A2 => n24943, Z => n21661);
   U20386 : XOR2_X1 port map( A1 => n22303, A2 => n10979, Z => n22155);
   U20391 : XOR2_X1 port map( A1 => n19517, A2 => n10986, Z => n10985);
   U20392 : NAND2_X1 port map( A1 => n26830, A2 => n19229, ZN => n15845);
   U20395 : XOR2_X1 port map( A1 => n22244, A2 => n10990, Z => n10989);
   U20396 : XOR2_X1 port map( A1 => n22291, A2 => n10991, Z => n10990);
   U20397 : INV_X1 port map( I => n24968, ZN => n10991);
   U20398 : NAND2_X2 port map( A1 => n16364, A2 => n19810, ZN => n20429);
   U20400 : XOR2_X1 port map( A1 => n23526, A2 => n23525, Z => n23931);
   U20409 : INV_X2 port map( I => n11006, ZN => n12657);
   U20410 : XOR2_X1 port map( A1 => n27138, A2 => n32918, Z => n19700);
   U20411 : XOR2_X1 port map( A1 => n32889, A2 => n21016, Z => n11012);
   U20417 : XOR2_X1 port map( A1 => n22085, A2 => n11028, Z => n11027);
   U20418 : INV_X1 port map( I => n16636, ZN => n11028);
   U20422 : XOR2_X1 port map( A1 => n400, A2 => n25036, Z => n19638);
   U20425 : NAND2_X1 port map( A1 => n16291, A2 => n25276, ZN => n25280);
   U20427 : XOR2_X1 port map( A1 => n10870, A2 => n16438, Z => n15775);
   U20431 : NAND3_X1 port map( A1 => n32941, A2 => n13499, A3 => n33721, ZN => 
                           n20051);
   U20433 : XOR2_X1 port map( A1 => n20985, A2 => n12957, Z => n20896);
   U20434 : XOR2_X1 port map( A1 => n7256, A2 => n16685, Z => n24628);
   U20441 : NOR2_X1 port map( A1 => n23578, A2 => n12287, ZN => n11095);
   U20442 : NAND3_X1 port map( A1 => n14232, A2 => n23958, A3 => n11096, ZN => 
                           n23959);
   U20443 : MUX2_X1 port map( I0 => n21252, I1 => n17437, S => n1337, Z => 
                           n21254);
   U20444 : AOI22_X1 port map( A1 => n16017, A2 => n30283, B1 => n14677, B2 => 
                           n11107, ZN => n24036);
   U20449 : XOR2_X1 port map( A1 => n20982, A2 => n25648, Z => n11118);
   U20451 : XOR2_X1 port map( A1 => n11128, A2 => n15460, Z => n11124);
   U20453 : XOR2_X1 port map( A1 => n22128, A2 => n2353, Z => n11126);
   U20455 : XOR2_X1 port map( A1 => n11130, A2 => n11129, Z => n13080);
   U20456 : XOR2_X1 port map( A1 => n19441, A2 => n19442, Z => n11129);
   U20457 : XOR2_X1 port map( A1 => n13829, A2 => n12453, Z => n11130);
   U20460 : INV_X1 port map( I => n17110, ZN => n14509);
   U20461 : NOR2_X1 port map( A1 => n34109, A2 => n25247, ZN => n11136);
   U20466 : NOR2_X1 port map( A1 => n14376, A2 => n11147, ZN => n11146);
   U20467 : XOR2_X1 port map( A1 => n23190, A2 => n12123, Z => n11148);
   U20468 : XOR2_X1 port map( A1 => n23363, A2 => n23189, Z => n23276);
   U20470 : NAND2_X1 port map( A1 => n17661, A2 => n23806, ZN => n11159);
   U20472 : XOR2_X1 port map( A1 => n25969, A2 => n25908, Z => n20482);
   U20474 : INV_X1 port map( I => n21811, ZN => n14917);
   U20475 : AOI21_X2 port map( A1 => n21809, A2 => n2801, B => n11167, ZN => 
                           n11166);
   U20476 : XOR2_X1 port map( A1 => n24638, A2 => n25252, Z => n11170);
   U20477 : XOR2_X1 port map( A1 => n24455, A2 => n24600, Z => n11171);
   U20480 : INV_X2 port map( I => n11175, ZN => n22640);
   U20484 : XOR2_X1 port map( A1 => n23393, A2 => n26701, Z => n11194);
   U20491 : XOR2_X1 port map( A1 => n11206, A2 => n21886, Z => n21997);
   U20497 : AND3_X1 port map( A1 => n26026, A2 => n17828, A3 => n23104, Z => 
                           n17585);
   U20498 : XOR2_X1 port map( A1 => n11225, A2 => n11223, Z => n12906);
   U20503 : XOR2_X1 port map( A1 => n23453, A2 => n1402, Z => n11227);
   U20511 : INV_X1 port map( I => n25285, ZN => n25279);
   U20512 : NAND2_X1 port map( A1 => n18483, A2 => n9549, ZN => n15165);
   U20513 : INV_X2 port map( I => n24565, ZN => n25295);
   U20520 : INV_X2 port map( I => n11281, ZN => n11916);
   U20523 : XOR2_X1 port map( A1 => n23532, A2 => n25735, Z => n16263);
   U20526 : NOR2_X1 port map( A1 => n11734, A2 => n11966, ZN => n11285);
   U20527 : XOR2_X1 port map( A1 => n11290, A2 => n14481, Z => n11289);
   U20532 : XOR2_X1 port map( A1 => n11297, A2 => n29707, Z => n14079);
   U20534 : XOR2_X1 port map( A1 => n11297, A2 => n31687, Z => n24423);
   U20535 : XOR2_X1 port map( A1 => n11297, A2 => n16671, Z => n24048);
   U20536 : NAND2_X1 port map( A1 => n11302, A2 => n743, ZN => n19219);
   U20542 : XOR2_X1 port map( A1 => Plaintext(156), A2 => Key(156), Z => n14159
                           );
   U20543 : OR2_X1 port map( A1 => n18543, A2 => n18858, Z => n11318);
   U20548 : XOR2_X1 port map( A1 => n24642, A2 => n24861, Z => n24517);
   U20549 : INV_X2 port map( I => n15401, ZN => n23755);
   U20550 : XOR2_X1 port map( A1 => n22616, A2 => n11326, Z => n13132);
   U20551 : NAND3_X2 port map( A1 => n21757, A2 => n11719, A3 => n15410, ZN => 
                           n22096);
   U20552 : XOR2_X1 port map( A1 => n20989, A2 => n11339, Z => n11338);
   U20553 : XOR2_X1 port map( A1 => n20904, A2 => n16672, Z => n11339);
   U20555 : INV_X2 port map( I => n11348, ZN => n14290);
   U20556 : XOR2_X1 port map( A1 => n11353, A2 => n11351, Z => n11910);
   U20558 : XOR2_X1 port map( A1 => n11354, A2 => n19707, Z => n11353);
   U20560 : XOR2_X1 port map( A1 => n11357, A2 => n11356, Z => n11355);
   U20561 : XOR2_X1 port map( A1 => n22189, A2 => n30954, Z => n11356);
   U20562 : XOR2_X1 port map( A1 => n2896, A2 => n4342, Z => n11357);
   U20566 : NOR2_X1 port map( A1 => n25082, A2 => n11360, ZN => n25094);
   U20568 : XOR2_X1 port map( A1 => n19494, A2 => n25288, Z => n11361);
   U20569 : NAND3_X1 port map( A1 => n15434, A2 => n15005, A3 => n14545, ZN => 
                           n13933);
   U20570 : INV_X2 port map( I => n11364, ZN => n16317);
   U20574 : XOR2_X1 port map( A1 => n11722, A2 => n25720, Z => n24639);
   U20580 : XOR2_X1 port map( A1 => Plaintext(26), A2 => Key(26), Z => n11599);
   U20581 : XNOR2_X1 port map( A1 => Plaintext(103), A2 => Key(103), ZN => 
                           n11379);
   U20583 : NOR2_X1 port map( A1 => n27188, A2 => n18151, ZN => n12235);
   U20585 : NAND2_X1 port map( A1 => n962, A2 => n11390, ZN => n14543);
   U20588 : XOR2_X1 port map( A1 => n11568, A2 => n22728, Z => n23745);
   U20589 : NOR2_X2 port map( A1 => n6783, A2 => n12290, ZN => n12238);
   U20595 : OAI21_X2 port map( A1 => n24485, A2 => n29629, B => n11429, ZN => 
                           n24960);
   U20596 : XOR2_X1 port map( A1 => n19564, A2 => n11433, Z => n11432);
   U20597 : XOR2_X1 port map( A1 => n15117, A2 => n25324, Z => n11433);
   U20601 : NOR2_X1 port map( A1 => n16627, A2 => n22435, ZN => n11443);
   U20602 : XOR2_X1 port map( A1 => n14214, A2 => n17551, Z => n11450);
   U20603 : XNOR2_X1 port map( A1 => n19408, A2 => n19398, ZN => n18072);
   U20604 : INV_X2 port map( I => n11451, ZN => n16627);
   U20608 : XOR2_X1 port map( A1 => n26562, A2 => n20389, Z => n18113);
   U20609 : NAND2_X1 port map( A1 => n10181, A2 => n11459, ZN => n14695);
   U20611 : XOR2_X1 port map( A1 => Plaintext(177), A2 => Key(177), Z => n18873
                           );
   U20613 : NOR2_X1 port map( A1 => n10673, A2 => n499, ZN => n23633);
   U20614 : OAI21_X1 port map( A1 => n17947, A2 => n4254, B => n20486, ZN => 
                           n11465);
   U20615 : INV_X1 port map( I => n11468, ZN => n25153);
   U20616 : OAI22_X1 port map( A1 => n25166, A2 => n25174, B1 => n25179, B2 => 
                           n11468, ZN => n12457);
   U20617 : OAI21_X2 port map( A1 => n14971, A2 => n33904, B => n24463, ZN => 
                           n24956);
   U20618 : XOR2_X1 port map( A1 => n30628, A2 => n1196, Z => n11476);
   U20620 : XOR2_X1 port map( A1 => n11485, A2 => n11484, Z => n11483);
   U20622 : XOR2_X1 port map( A1 => n16693, A2 => n705, Z => n11485);
   U20624 : INV_X1 port map( I => n21258, ZN => n21255);
   U20626 : XOR2_X1 port map( A1 => n19541, A2 => n17072, Z => n11488);
   U20630 : XOR2_X1 port map( A1 => n1045, A2 => n13826, Z => n17213);
   U20632 : XOR2_X1 port map( A1 => n11504, A2 => n25506, Z => n23167);
   U20635 : NAND2_X2 port map( A1 => n19040, A2 => n19042, ZN => n13925);
   U20638 : XOR2_X1 port map( A1 => n19495, A2 => n11523, Z => n11522);
   U20639 : XOR2_X1 port map( A1 => n30193, A2 => n1419, Z => n11523);
   U20640 : XOR2_X1 port map( A1 => n17552, A2 => n15983, Z => n11524);
   U20641 : XOR2_X1 port map( A1 => n13810, A2 => n11526, Z => n11525);
   U20642 : XOR2_X1 port map( A1 => n24675, A2 => n7603, Z => n11526);
   U20643 : XOR2_X1 port map( A1 => n11529, A2 => n11528, Z => n22486);
   U20645 : XOR2_X1 port map( A1 => n16457, A2 => n17174, Z => n11529);
   U20646 : XOR2_X1 port map( A1 => n11532, A2 => n11531, Z => n11530);
   U20647 : XOR2_X1 port map( A1 => n13970, A2 => n13331, Z => n11531);
   U20651 : XOR2_X1 port map( A1 => n16513, A2 => n11544, Z => n11543);
   U20652 : XOR2_X1 port map( A1 => n16349, A2 => n19649, Z => n11544);
   U20655 : NOR2_X1 port map( A1 => n25391, A2 => n32884, ZN => n25392);
   U20657 : XOR2_X1 port map( A1 => n11558, A2 => n16649, Z => Ciphertext(91));
   U20659 : XOR2_X1 port map( A1 => n22032, A2 => n16703, Z => n11819);
   U20662 : NOR2_X1 port map( A1 => n11567, A2 => n30089, ZN => n23597);
   U20664 : XOR2_X1 port map( A1 => n9434, A2 => n30943, Z => n11574);
   U20665 : XOR2_X1 port map( A1 => n11578, A2 => n516, Z => n11577);
   U20668 : XOR2_X1 port map( A1 => n18401, A2 => Key(172), Z => n18847);
   U20673 : AND2_X1 port map( A1 => n11601, A2 => n21070, Z => n12933);
   U20676 : INV_X1 port map( I => n16674, ZN => n11603);
   U20677 : XOR2_X1 port map( A1 => n19772, A2 => n11604, Z => n19775);
   U20678 : XOR2_X1 port map( A1 => n22790, A2 => n11611, Z => n11610);
   U20679 : XOR2_X1 port map( A1 => n10773, A2 => n1393, Z => n11611);
   U20680 : XOR2_X1 port map( A1 => n23318, A2 => n23273, Z => n22790);
   U20681 : XOR2_X1 port map( A1 => n23173, A2 => n23460, Z => n11612);
   U20682 : NOR2_X1 port map( A1 => n13175, A2 => n24110, ZN => n11613);
   U20684 : INV_X2 port map( I => n11620, ZN => n22476);
   U20686 : XNOR2_X1 port map( A1 => n471, A2 => n11631, ZN => n11630);
   U20687 : XOR2_X1 port map( A1 => n17840, A2 => n19536, Z => n11631);
   U20689 : XOR2_X1 port map( A1 => Plaintext(74), A2 => Key(74), Z => n11773);
   U20692 : XOR2_X1 port map( A1 => n33453, A2 => n15816, Z => n17095);
   U20693 : XOR2_X1 port map( A1 => n33453, A2 => n23191, Z => n14967);
   U20698 : NAND2_X1 port map( A1 => n24250, A2 => n28553, ZN => n17409);
   U20702 : XOR2_X1 port map( A1 => n19780, A2 => n24964, Z => n11661);
   U20705 : XOR2_X1 port map( A1 => n1369, A2 => n876, Z => n11663);
   U20709 : NAND2_X2 port map( A1 => n11675, A2 => n12187, ZN => n24393);
   U20710 : XOR2_X1 port map( A1 => n18356, A2 => Key(18), Z => n18654);
   U20712 : NOR2_X1 port map( A1 => n1334, A2 => n11814, ZN => n11680);
   U20713 : XOR2_X1 port map( A1 => n24676, A2 => n16533, Z => n11681);
   U20714 : NAND2_X2 port map( A1 => n11686, A2 => n11682, ZN => n15296);
   U20715 : XOR2_X1 port map( A1 => n11689, A2 => n11690, Z => n16784);
   U20716 : XOR2_X1 port map( A1 => n20894, A2 => n15652, Z => n11690);
   U20719 : XOR2_X1 port map( A1 => n24652, A2 => n15779, Z => n11699);
   U20726 : XOR2_X1 port map( A1 => n5932, A2 => n25990, Z => n14363);
   U20727 : XOR2_X1 port map( A1 => n31508, A2 => n25991, Z => n24651);
   U20733 : XOR2_X1 port map( A1 => n22063, A2 => n16479, Z => n11750);
   U20736 : INV_X1 port map( I => n23263, ZN => n11766);
   U20739 : XOR2_X1 port map( A1 => n17091, A2 => n33918, Z => n19481);
   U20740 : XNOR2_X1 port map( A1 => n17091, A2 => n19337, ZN => n15157);
   U20741 : INV_X2 port map( I => n11773, ZN => n18559);
   U20743 : XOR2_X1 port map( A1 => n14656, A2 => n11776, Z => n11775);
   U20744 : XOR2_X1 port map( A1 => n24836, A2 => n14533, Z => n11782);
   U20745 : XOR2_X1 port map( A1 => n32310, A2 => n27920, Z => n11783);
   U20747 : XOR2_X1 port map( A1 => n17301, A2 => n16507, Z => n11803);
   U20749 : XOR2_X1 port map( A1 => n27252, A2 => n15415, Z => n13739);
   U20751 : XOR2_X1 port map( A1 => n20954, A2 => n20955, Z => n14854);
   U20752 : XOR2_X1 port map( A1 => n19445, A2 => n33587, Z => n11817);
   U20756 : XOR2_X1 port map( A1 => n11841, A2 => n11843, Z => n11844);
   U20757 : XOR2_X1 port map( A1 => n11842, A2 => n24637, Z => n11841);
   U20759 : INV_X2 port map( I => n11844, ZN => n12042);
   U20761 : XNOR2_X1 port map( A1 => n15047, A2 => n15048, ZN => n11847);
   U20763 : NAND3_X2 port map( A1 => n11854, A2 => n22458, A3 => n11853, ZN => 
                           n23086);
   U20764 : NAND2_X1 port map( A1 => n17670, A2 => n11855, ZN => n19547);
   U20767 : NAND2_X1 port map( A1 => n15797, A2 => n15796, ZN => n11860);
   U20768 : NAND3_X2 port map( A1 => n17101, A2 => n16048, A3 => n20373, ZN => 
                           n12424);
   U20772 : XOR2_X1 port map( A1 => n11869, A2 => n14401, Z => n14400);
   U20773 : XOR2_X1 port map( A1 => n24805, A2 => n5268, Z => n24668);
   U20777 : OAI21_X1 port map( A1 => n694, A2 => n25322, B => n16041, ZN => 
                           n15854);
   U20778 : NAND3_X1 port map( A1 => n32867, A2 => n16041, A3 => n694, ZN => 
                           n25309);
   U20779 : INV_X2 port map( I => n11877, ZN => n18035);
   U20781 : XOR2_X1 port map( A1 => n18348, A2 => Key(37), Z => n18548);
   U20787 : INV_X1 port map( I => n33848, ZN => n20034);
   U20788 : NAND4_X1 port map( A1 => n11214, A2 => n12642, A3 => n12640, A4 => 
                           n12641, ZN => n21546);
   U20789 : NOR2_X1 port map( A1 => n20944, A2 => n21181, ZN => n15321);
   U20790 : AOI22_X1 port map( A1 => n24780, A2 => n24874, B1 => n10770, B2 => 
                           n15719, ZN => n15234);
   U20792 : NOR2_X1 port map( A1 => n1205, A2 => n24998, ZN => n14837);
   U20793 : NAND3_X1 port map( A1 => n1291, A2 => n29336, A3 => n855, ZN => 
                           n14772);
   U20794 : NAND2_X1 port map( A1 => n13962, A2 => n31161, ZN => n15135);
   U20797 : INV_X1 port map( I => n12257, ZN => n15062);
   U20798 : NAND2_X1 port map( A1 => n18437, A2 => n958, ZN => n16207);
   U20799 : NOR2_X1 port map( A1 => n18007, A2 => n18427, ZN => n18428);
   U20802 : INV_X1 port map( I => n19412, ZN => n19592);
   U20804 : NOR2_X1 port map( A1 => n12244, A2 => n20338, ZN => n12843);
   U20805 : INV_X1 port map( I => n20574, ZN => n12812);
   U20818 : INV_X1 port map( I => n18623, ZN => n18771);
   U20821 : INV_X1 port map( I => n18423, ZN => n17102);
   U20824 : NAND2_X1 port map( A1 => n14828, A2 => n13738, ZN => n17231);
   U20834 : INV_X1 port map( I => n20842, ZN => n17759);
   U20839 : NAND4_X1 port map( A1 => n13285, A2 => n13284, A3 => n19892, A4 => 
                           n13283, ZN => n13282);
   U20844 : INV_X1 port map( I => n17672, ZN => n20266);
   U20847 : INV_X1 port map( I => n20351, ZN => n12367);
   U20850 : NAND2_X1 port map( A1 => n14156, A2 => n9437, ZN => n13788);
   U20852 : NOR2_X1 port map( A1 => n962, A2 => n14926, ZN => n12291);
   U20854 : NAND2_X1 port map( A1 => n16226, A2 => n29256, ZN => n14174);
   U20855 : NAND2_X1 port map( A1 => n21365, A2 => n20945, ZN => n20705);
   U20858 : NAND2_X1 port map( A1 => n19258, A2 => n19257, ZN => n19259);
   U20865 : NAND2_X1 port map( A1 => n957, A2 => n12956, ZN => n18519);
   U20874 : NAND2_X1 port map( A1 => n18439, A2 => n19355, ZN => n17996);
   U20875 : NOR2_X1 port map( A1 => n13390, A2 => n28386, ZN => n18439);
   U20878 : NAND2_X1 port map( A1 => n18825, A2 => n17553, ZN => n14859);
   U20880 : NAND3_X1 port map( A1 => n15417, A2 => n1048, A3 => n15780, ZN => 
                           n18452);
   U20881 : NAND2_X1 port map( A1 => n19271, A2 => n19265, ZN => n15780);
   U20882 : INV_X1 port map( I => n21379, ZN => n21178);
   U20883 : OAI21_X1 port map( A1 => n16905, A2 => n13319, B => n13581, ZN => 
                           n13580);
   U20885 : NAND3_X1 port map( A1 => n14384, A2 => n8029, A3 => n31042, ZN => 
                           n21519);
   U20886 : OAI21_X1 port map( A1 => n17078, A2 => n14640, B => n15171, ZN => 
                           n21521);
   U20889 : NOR2_X1 port map( A1 => n14008, A2 => n15752, ZN => n15635);
   U20892 : NAND2_X1 port map( A1 => n22478, A2 => n22377, ZN => n13186);
   U20898 : NAND2_X1 port map( A1 => n16493, A2 => n16105, ZN => n16262);
   U20899 : INV_X1 port map( I => n19368, ZN => n17104);
   U20902 : NOR2_X1 port map( A1 => n13561, A2 => n14253, ZN => n13587);
   U20907 : AOI21_X1 port map( A1 => n23778, A2 => n8547, B => n23776, ZN => 
                           n13140);
   U20908 : NAND2_X1 port map( A1 => n28367, A2 => n23871, ZN => n23876);
   U20917 : INV_X1 port map( I => n12720, ZN => n13825);
   U20918 : INV_X1 port map( I => n24356, ZN => n24493);
   U20919 : NAND2_X1 port map( A1 => n17047, A2 => n17037, ZN => n17046);
   U20922 : INV_X1 port map( I => n20454, ZN => n14086);
   U20925 : NAND2_X1 port map( A1 => n868, A2 => n20525, ZN => n20276);
   U20927 : INV_X1 port map( I => n20350, ZN => n12366);
   U20931 : INV_X1 port map( I => n25856, ZN => n14557);
   U20934 : INV_X1 port map( I => n18882, ZN => n17478);
   U20936 : INV_X1 port map( I => n18695, ZN => n18697);
   U20937 : NOR2_X1 port map( A1 => n30271, A2 => n12006, ZN => n15141);
   U20938 : AOI22_X1 port map( A1 => n14271, A2 => n15589, B1 => n7690, B2 => 
                           n3931, ZN => n14270);
   U20939 : NOR2_X1 port map( A1 => n15261, A2 => n14721, ZN => n14271);
   U20943 : NAND2_X1 port map( A1 => n15874, A2 => n21398, ZN => n16258);
   U20946 : INV_X1 port map( I => n17822, ZN => n14305);
   U20947 : NAND2_X1 port map( A1 => n14290, A2 => n1335, ZN => n15160);
   U20950 : NOR2_X1 port map( A1 => n21073, A2 => n29255, ZN => n16844);
   U20951 : INV_X1 port map( I => n16545, ZN => n16544);
   U20958 : INV_X1 port map( I => n21362, ZN => n14903);
   U20963 : AOI21_X1 port map( A1 => n16403, A2 => n18801, B => n18785, ZN => 
                           n18629);
   U20964 : NAND2_X1 port map( A1 => n828, A2 => n18775, ZN => n18624);
   U20966 : NOR2_X1 port map( A1 => n13254, A2 => n12317, ZN => n13408);
   U20970 : NOR2_X1 port map( A1 => n1048, A2 => n31726, ZN => n18975);
   U20972 : NOR2_X1 port map( A1 => n19097, A2 => n19098, ZN => n14030);
   U20973 : NAND2_X1 port map( A1 => n21095, A2 => n8190, ZN => n21295);
   U20975 : AOI21_X1 port map( A1 => n26782, A2 => n15838, B => n21793, ZN => 
                           n21791);
   U20977 : NOR2_X1 port map( A1 => n14488, A2 => n29497, ZN => n14487);
   U20978 : NOR2_X1 port map( A1 => n14489, A2 => n21412, ZN => n14488);
   U20981 : NAND3_X1 port map( A1 => n21084, A2 => n28406, A3 => n17985, ZN => 
                           n13315);
   U20987 : NAND3_X1 port map( A1 => n9, A2 => n15956, A3 => n18829, ZN => 
                           n17135);
   U20993 : NAND2_X1 port map( A1 => n16624, A2 => n16417, ZN => n12799);
   U20995 : AOI21_X1 port map( A1 => n10828, A2 => n19165, B => n19308, ZN => 
                           n15930);
   U20997 : NAND2_X1 port map( A1 => n17737, A2 => n17736, ZN => n17735);
   U21009 : NAND2_X1 port map( A1 => n19037, A2 => n2901, ZN => n14455);
   U21010 : NAND2_X1 port map( A1 => n16916, A2 => n27587, ZN => n12645);
   U21013 : INV_X1 port map( I => n33698, ZN => n19767);
   U21014 : NAND3_X1 port map( A1 => n19255, A2 => n19143, A3 => n1180, ZN => 
                           n18528);
   U21018 : NOR2_X1 port map( A1 => n30205, A2 => n137, ZN => n13485);
   U21022 : INV_X1 port map( I => n22536, ZN => n12844);
   U21031 : NAND2_X1 port map( A1 => n20255, A2 => n16951, ZN => n13380);
   U21040 : INV_X1 port map( I => n22619, ZN => n15349);
   U21042 : NAND2_X1 port map( A1 => n7957, A2 => n708, ZN => n22253);
   U21044 : INV_X1 port map( I => n23218, ZN => n23250);
   U21046 : NAND2_X1 port map( A1 => n19947, A2 => n15110, ZN => n15109);
   U21047 : OAI21_X1 port map( A1 => n11958, A2 => n20056, B => n14099, ZN => 
                           n17945);
   U21051 : NAND2_X1 port map( A1 => n23637, A2 => n13137, ZN => n13136);
   U21054 : NOR2_X1 port map( A1 => n23797, A2 => n14193, ZN => n15187);
   U21057 : INV_X1 port map( I => n23490, ZN => n17194);
   U21058 : INV_X1 port map( I => n23583, ZN => n14523);
   U21061 : OAI21_X1 port map( A1 => n23653, A2 => n8547, B => n13140, ZN => 
                           n13139);
   U21066 : NAND2_X1 port map( A1 => n13905, A2 => n23759, ZN => n13904);
   U21068 : INV_X1 port map( I => n23958, ZN => n23957);
   U21073 : INV_X1 port map( I => n16634, ZN => n15000);
   U21074 : INV_X1 port map( I => n13698, ZN => n16826);
   U21075 : INV_X1 port map( I => n13060, ZN => n12513);
   U21077 : INV_X1 port map( I => n11974, ZN => n14020);
   U21081 : NOR2_X1 port map( A1 => n24975, A2 => n25012, ZN => n14992);
   U21084 : NAND2_X1 port map( A1 => n13349, A2 => n4993, ZN => n24733);
   U21089 : NOR2_X1 port map( A1 => n15756, A2 => n16451, ZN => n15755);
   U21091 : NOR2_X1 port map( A1 => n15770, A2 => n28136, ZN => n15757);
   U21092 : INV_X2 port map( I => n17044, ZN => n25536);
   U21093 : NOR2_X1 port map( A1 => n11900, A2 => n11090, ZN => n13323);
   U21097 : NAND2_X1 port map( A1 => n965, A2 => n24960, ZN => n14933);
   U21099 : OAI21_X1 port map( A1 => n12783, A2 => n33434, B => n12204, ZN => 
                           n12203);
   U21100 : NAND2_X1 port map( A1 => n24972, A2 => n8622, ZN => n12204);
   U21101 : NAND2_X1 port map( A1 => n24969, A2 => n24970, ZN => n13737);
   U21103 : INV_X1 port map( I => n14638, ZN => n14637);
   U21104 : NAND2_X1 port map( A1 => n1074, A2 => n72, ZN => n15858);
   U21109 : INV_X1 port map( I => n20953, ZN => n20997);
   U21110 : NAND3_X1 port map( A1 => n20498, A2 => n20497, A3 => n30869, ZN => 
                           n16759);
   U21115 : NAND2_X1 port map( A1 => n20461, A2 => n20462, ZN => n13546);
   U21116 : INV_X1 port map( I => n20773, ZN => n12732);
   U21117 : NAND2_X1 port map( A1 => n13700, A2 => n21182, ZN => n12913);
   U21119 : NAND3_X1 port map( A1 => n14486, A2 => n14485, A3 => n16584, ZN => 
                           n14294);
   U21120 : NAND2_X1 port map( A1 => n10182, A2 => n11459, ZN => n15575);
   U21125 : NOR2_X1 port map( A1 => n18797, A2 => n16420, ZN => n17926);
   U21128 : NOR2_X1 port map( A1 => n1017, A2 => n21267, ZN => n21064);
   U21134 : INV_X1 port map( I => n12654, ZN => n14860);
   U21136 : OAI21_X1 port map( A1 => n14802, A2 => n21379, B => n7007, ZN => 
                           n21179);
   U21139 : NAND2_X1 port map( A1 => n13506, A2 => n21424, ZN => n17666);
   U21141 : NOR2_X1 port map( A1 => n13149, A2 => n21634, ZN => n13148);
   U21143 : NOR2_X1 port map( A1 => n21366, A2 => n21365, ZN => n12348);
   U21146 : AOI21_X1 port map( A1 => n6783, A2 => n962, B => n12290, ZN => 
                           n12197);
   U21148 : NOR2_X1 port map( A1 => n9423, A2 => n19355, ZN => n16750);
   U21152 : AOI21_X1 port map( A1 => n13787, A2 => n9437, B => n18638, ZN => 
                           n13201);
   U21155 : NAND2_X1 port map( A1 => n19268, A2 => n18974, ZN => n18449);
   U21158 : NAND2_X1 port map( A1 => n16487, A2 => n18706, ZN => n18708);
   U21159 : NOR2_X1 port map( A1 => n33078, A2 => n19178, ZN => n14426);
   U21160 : NOR2_X1 port map( A1 => n4016, A2 => n19348, ZN => n19218);
   U21164 : AOI21_X1 port map( A1 => n15874, A2 => n27955, B => n21143, ZN => 
                           n15024);
   U21165 : NAND3_X1 port map( A1 => n29552, A2 => n6176, A3 => n21772, ZN => 
                           n14868);
   U21169 : NAND2_X1 port map( A1 => n31826, A2 => n26021, ZN => n12507);
   U21171 : NOR2_X1 port map( A1 => n21052, A2 => n21257, ZN => n14643);
   U21172 : NAND2_X1 port map( A1 => n8631, A2 => n2738, ZN => n14853);
   U21175 : INV_X1 port map( I => n22021, ZN => n22162);
   U21178 : NAND2_X1 port map( A1 => n15774, A2 => n21812, ZN => n13167);
   U21182 : AOI21_X1 port map( A1 => n19323, A2 => n19317, B => n19324, ZN => 
                           n12384);
   U21183 : AND2_X1 port map( A1 => n6416, A2 => n16538, Z => n14696);
   U21184 : INV_X1 port map( I => n17165, ZN => n18865);
   U21188 : AOI21_X1 port map( A1 => n18432, A2 => n18433, B => n18743, ZN => 
                           n13501);
   U21191 : INV_X1 port map( I => n18135, ZN => n12928);
   U21193 : NAND2_X1 port map( A1 => n19114, A2 => n19115, ZN => n13227);
   U21196 : NOR2_X1 port map( A1 => n17455, A2 => n9721, ZN => n14999);
   U21204 : NAND2_X1 port map( A1 => n16447, A2 => n22403, ZN => n15204);
   U21205 : NAND2_X1 port map( A1 => n22678, A2 => n22562, ZN => n13710);
   U21206 : INV_X1 port map( I => n19878, ZN => n13987);
   U21209 : NAND2_X1 port map( A1 => n33561, A2 => n29013, ZN => n15737);
   U21211 : NOR2_X1 port map( A1 => n18803, A2 => n16403, ZN => n12175);
   U21214 : NOR2_X1 port map( A1 => n3626, A2 => n3790, ZN => n12590);
   U21218 : NOR2_X1 port map( A1 => n6275, A2 => n33264, ZN => n15267);
   U21220 : INV_X1 port map( I => n28638, ZN => n17293);
   U21221 : INV_X1 port map( I => n32057, ZN => n17291);
   U21222 : NOR2_X1 port map( A1 => n20059, A2 => n17608, ZN => n19420);
   U21227 : NOR2_X1 port map( A1 => n12112, A2 => n22610, ZN => n14157);
   U21229 : NOR2_X1 port map( A1 => n15008, A2 => n22570, ZN => n14081);
   U21233 : NAND2_X1 port map( A1 => n22503, A2 => n34125, ZN => n12254);
   U21234 : AOI21_X1 port map( A1 => n15322, A2 => n701, B => n22434, ZN => 
                           n14591);
   U21237 : NAND2_X1 port map( A1 => n873, A2 => n19819, ZN => n13451);
   U21239 : INV_X1 port map( I => n20133, ZN => n20025);
   U21240 : OAI21_X1 port map( A1 => n19987, A2 => n16623, B => n14440, ZN => 
                           n19339);
   U21241 : NOR2_X1 port map( A1 => n19986, A2 => n19998, ZN => n14622);
   U21242 : NOR2_X1 port map( A1 => n19308, A2 => n19165, ZN => n17526);
   U21248 : INV_X1 port map( I => n20079, ZN => n19803);
   U21261 : NOR2_X1 port map( A1 => n137, A2 => n31964, ZN => n14160);
   U21271 : NAND2_X1 port map( A1 => n15230, A2 => n6996, ZN => n20400);
   U21274 : NAND2_X1 port map( A1 => n13499, A2 => n16144, ZN => n14265);
   U21276 : NAND2_X1 port map( A1 => n22490, A2 => n22489, ZN => n12930);
   U21279 : AND2_X1 port map( A1 => n16078, A2 => n23003, Z => n11929);
   U21280 : NAND2_X1 port map( A1 => n23848, A2 => n23847, ZN => n13576);
   U21282 : NOR2_X1 port map( A1 => n20239, A2 => n20238, ZN => n17317);
   U21283 : NAND2_X1 port map( A1 => n1255, A2 => n14164, ZN => n13982);
   U21287 : OAI22_X1 port map( A1 => n17665, A2 => n13125, B1 => n16431, B2 => 
                           n23951, ZN => n17664);
   U21298 : NAND3_X1 port map( A1 => n23528, A2 => n23933, A3 => n23681, ZN => 
                           n12546);
   U21299 : NAND2_X1 port map( A1 => n23698, A2 => n23867, ZN => n13138);
   U21301 : NOR2_X1 port map( A1 => n13048, A2 => n24276, ZN => n13047);
   U21304 : NAND3_X1 port map( A1 => n16343, A2 => n16496, A3 => n29965, ZN => 
                           n23131);
   U21308 : NOR2_X1 port map( A1 => n24150, A2 => n797, ZN => n12189);
   U21312 : NAND2_X1 port map( A1 => n23718, A2 => n13031, ZN => n14924);
   U21317 : NAND3_X1 port map( A1 => n23770, A2 => n11567, A3 => n23769, ZN => 
                           n15402);
   U21318 : INV_X1 port map( I => n12775, ZN => n12774);
   U21329 : NOR2_X1 port map( A1 => n24153, A2 => n1245, ZN => n16983);
   U21331 : NOR2_X1 port map( A1 => n25013, A2 => n31274, ZN => n14021);
   U21333 : NAND2_X1 port map( A1 => n17110, A2 => n7081, ZN => n25197);
   U21336 : AOI21_X1 port map( A1 => n17038, A2 => n25539, B => n24667, ZN => 
                           n16828);
   U21337 : INV_X1 port map( I => n25876, ZN => n17762);
   U21340 : OAI21_X1 port map( A1 => n25398, A2 => n25403, B => n25397, ZN => 
                           n15882);
   U21342 : NOR2_X1 port map( A1 => n31783, A2 => n25198, ZN => n15705);
   U21350 : NOR2_X1 port map( A1 => n11090, A2 => n25582, ZN => n15598);
   U21351 : OAI21_X1 port map( A1 => n11945, A2 => n17118, B => n15046, ZN => 
                           n24462);
   U21354 : NAND2_X1 port map( A1 => n24955, A2 => n24956, ZN => n14932);
   U21357 : NAND2_X1 port map( A1 => n30302, A2 => n25375, ZN => n15478);
   U21361 : OAI21_X1 port map( A1 => n14454, A2 => n15084, B => n15223, ZN => 
                           n17771);
   U21365 : NOR2_X1 port map( A1 => n27118, A2 => n1223, ZN => n15673);
   U21371 : INV_X1 port map( I => n17594, ZN => n15332);
   U21372 : NAND3_X1 port map( A1 => n14627, A2 => n15641, A3 => n25145, ZN => 
                           n14631);
   U21373 : NOR2_X1 port map( A1 => n25199, A2 => n12476, ZN => n25147);
   U21374 : NAND2_X1 port map( A1 => n966, A2 => n25214, ZN => n25215);
   U21375 : NAND2_X1 port map( A1 => n25231, A2 => n25398, ZN => n17924);
   U21376 : NOR2_X1 port map( A1 => n15770, A2 => n17717, ZN => n15896);
   U21379 : NAND2_X1 port map( A1 => n25369, A2 => n25376, ZN => n16246);
   U21380 : NAND2_X1 port map( A1 => n24863, A2 => n9858, ZN => n16187);
   U21381 : AOI21_X1 port map( A1 => n25564, A2 => n17655, B => n25582, ZN => 
                           n13322);
   U21382 : NAND3_X1 port map( A1 => n25752, A2 => n25707, A3 => n25620, ZN => 
                           n25580);
   U21385 : NAND2_X1 port map( A1 => n13768, A2 => n20236, ZN => n12224);
   U21391 : NAND2_X1 port map( A1 => n15006, A2 => n20417, ZN => n20274);
   U21398 : NOR2_X1 port map( A1 => n33515, A2 => n13759, ZN => n13786);
   U21399 : NAND2_X1 port map( A1 => n13880, A2 => n20524, ZN => n12345);
   U21402 : INV_X1 port map( I => n20498, ZN => n16762);
   U21404 : NOR2_X1 port map( A1 => n2618, A2 => n30987, ZN => n17758);
   U21405 : NOR2_X1 port map( A1 => n31835, A2 => n865, ZN => n16505);
   U21406 : NAND3_X1 port map( A1 => n17971, A2 => n28502, A3 => n21251, ZN => 
                           n20935);
   U21407 : NAND3_X1 port map( A1 => n779, A2 => n16933, A3 => n21249, ZN => 
                           n20936);
   U21413 : INV_X1 port map( I => n17984, ZN => n16780);
   U21415 : NOR2_X1 port map( A1 => n21473, A2 => n27532, ZN => n12275);
   U21418 : INV_X1 port map( I => n13872, ZN => n21458);
   U21424 : NAND2_X1 port map( A1 => n17687, A2 => n18738, ZN => n18531);
   U21425 : NAND2_X1 port map( A1 => n28171, A2 => n878, ZN => n12807);
   U21426 : NAND2_X1 port map( A1 => n882, A2 => n28707, ZN => n15927);
   U21429 : OAI21_X1 port map( A1 => n18843, A2 => n746, B => n25981, ZN => 
                           n16713);
   U21430 : NAND2_X1 port map( A1 => n19321, A2 => n19322, ZN => n19232);
   U21436 : AOI22_X1 port map( A1 => n12130, A2 => n30271, B1 => n13846, B2 => 
                           n18699, ZN => n15196);
   U21438 : NOR2_X1 port map( A1 => n13200, A2 => n19180, ZN => n19182);
   U21440 : INV_X1 port map( I => n19507, ZN => n12683);
   U21443 : NAND2_X1 port map( A1 => n21668, A2 => n918, ZN => n14673);
   U21445 : NAND2_X1 port map( A1 => n17547, A2 => n7553, ZN => n12786);
   U21446 : INV_X1 port map( I => n14950, ZN => n14949);
   U21449 : NAND2_X1 port map( A1 => n16519, A2 => n16165, ZN => n12712);
   U21450 : NAND2_X1 port map( A1 => n27336, A2 => n432, ZN => n16863);
   U21455 : INV_X1 port map( I => n34040, ZN => n19263);
   U21456 : NAND2_X1 port map( A1 => n19269, A2 => n19265, ZN => n15505);
   U21459 : NOR2_X1 port map( A1 => n18581, A2 => n17419, ZN => n13036);
   U21460 : NOR2_X1 port map( A1 => n16403, A2 => n18785, ZN => n18786);
   U21461 : NAND2_X1 port map( A1 => n4677, A2 => n18801, ZN => n18787);
   U21462 : NAND2_X1 port map( A1 => n746, A2 => n15873, ZN => n16867);
   U21463 : NAND2_X1 port map( A1 => n16370, A2 => n6783, ZN => n12196);
   U21471 : NAND2_X1 port map( A1 => n19181, A2 => n19118, ZN => n13012);
   U21475 : OAI21_X1 port map( A1 => n18467, A2 => n18468, B => n945, ZN => 
                           n13708);
   U21477 : NAND2_X1 port map( A1 => n18532, A2 => n17166, ZN => n15583);
   U21479 : AOI21_X1 port map( A1 => n15685, A2 => n18254, B => n18434, ZN => 
                           n18709);
   U21480 : INV_X1 port map( I => n18704, ZN => n15685);
   U21481 : NOR2_X1 port map( A1 => n33205, A2 => n16287, ZN => n17359);
   U21495 : NOR2_X1 port map( A1 => n919, A2 => n21687, ZN => n12332);
   U21497 : NOR2_X1 port map( A1 => n13500, A2 => n21641, ZN => n13613);
   U21500 : NOR2_X1 port map( A1 => n16519, A2 => n16165, ZN => n14503);
   U21501 : OAI21_X1 port map( A1 => n21840, A2 => n16987, B => n26163, ZN => 
                           n13815);
   U21504 : NOR2_X1 port map( A1 => n29854, A2 => n9076, ZN => n15680);
   U21509 : INV_X1 port map( I => n22160, ZN => n17968);
   U21512 : NAND2_X1 port map( A1 => n21731, A2 => n15655, ZN => n12939);
   U21516 : NOR2_X1 port map( A1 => n14976, A2 => n14172, ZN => n20093);
   U21523 : INV_X1 port map( I => n22220, ZN => n12681);
   U21528 : NOR2_X1 port map( A1 => n31017, A2 => n34103, ZN => n13655);
   U21529 : AOI21_X1 port map( A1 => n19862, A2 => n16579, B => n19863, ZN => 
                           n18002);
   U21530 : NOR3_X1 port map( A1 => n34103, A2 => n14458, A3 => n31017, ZN => 
                           n14282);
   U21534 : NAND3_X1 port map( A1 => n14747, A2 => n11959, A3 => n3486, ZN => 
                           n13570);
   U21535 : NOR3_X1 port map( A1 => n20142, A2 => n11911, A3 => n11248, ZN => 
                           n12851);
   U21540 : INV_X1 port map( I => n19984, ZN => n12397);
   U21541 : AOI21_X1 port map( A1 => n22803, A2 => n22983, B => n16140, ZN => 
                           n12596);
   U21546 : NOR2_X1 port map( A1 => n22805, A2 => n14420, ZN => n14419);
   U21549 : NAND2_X1 port map( A1 => n22798, A2 => n23053, ZN => n22868);
   U21551 : INV_X1 port map( I => n23336, ZN => n14583);
   U21552 : NAND3_X1 port map( A1 => n11980, A2 => n13892, A3 => n16486, ZN => 
                           n15577);
   U21554 : NAND2_X1 port map( A1 => n13575, A2 => n22780, ZN => n13574);
   U21558 : OAI21_X1 port map( A1 => n3184, A2 => n3183, B => n22781, ZN => 
                           n16716);
   U21559 : NOR2_X1 port map( A1 => n28948, A2 => n17084, ZN => n14603);
   U21562 : AOI21_X1 port map( A1 => n31684, A2 => n13061, B => n29013, ZN => 
                           n14989);
   U21564 : NAND2_X1 port map( A1 => n26232, A2 => n20577, ZN => n20579);
   U21565 : OAI21_X1 port map( A1 => n20153, A2 => n11199, B => n20150, ZN => 
                           n15350);
   U21568 : NAND2_X1 port map( A1 => n19812, A2 => n20018, ZN => n19814);
   U21575 : NAND2_X1 port map( A1 => n22952, A2 => n2479, ZN => n13004);
   U21578 : NAND2_X1 port map( A1 => n28277, A2 => n25994, ZN => n13251);
   U21582 : AOI21_X1 port map( A1 => n13995, A2 => n23106, B => n14131, ZN => 
                           n14552);
   U21588 : INV_X1 port map( I => n23375, ZN => n23260);
   U21596 : INV_X1 port map( I => n23507, ZN => n13287);
   U21605 : NAND2_X1 port map( A1 => n16167, A2 => n20510, ZN => n14366);
   U21607 : NOR2_X1 port map( A1 => n20228, A2 => n7242, ZN => n20516);
   U21609 : NOR2_X1 port map( A1 => n20337, A2 => n20531, ZN => n14261);
   U21611 : OAI21_X1 port map( A1 => n15806, A2 => n22865, B => n989, ZN => 
                           n22707);
   U21614 : INV_X1 port map( I => n16076, ZN => n23321);
   U21616 : NAND2_X1 port map( A1 => n20240, A2 => n27386, ZN => n16857);
   U21619 : INV_X1 port map( I => n24226, ZN => n24042);
   U21621 : NAND3_X1 port map( A1 => n24325, A2 => n7361, A3 => n24245, ZN => 
                           n24079);
   U21622 : INV_X1 port map( I => n24276, ZN => n24195);
   U21625 : OR3_X1 port map( A1 => n27430, A2 => n24304, A3 => n12904, Z => 
                           n11937);
   U21628 : NAND2_X1 port map( A1 => n13082, A2 => n32737, ZN => n12629);
   U21639 : AOI21_X1 port map( A1 => n12189, A2 => n2913, B => n12188, ZN => 
                           n12187);
   U21643 : OAI21_X1 port map( A1 => n791, A2 => n26916, B => n12357, ZN => 
                           n23626);
   U21645 : NOR2_X1 port map( A1 => n24270, A2 => n11768, ZN => n14502);
   U21646 : INV_X1 port map( I => n3935, ZN => n14938);
   U21650 : NAND3_X1 port map( A1 => n14889, A2 => n28694, A3 => n16621, ZN => 
                           n14888);
   U21651 : OAI21_X1 port map( A1 => n28694, A2 => n17261, B => n13260, ZN => 
                           n24229);
   U21652 : NAND2_X1 port map( A1 => n1786, A2 => n1850, ZN => n15254);
   U21654 : INV_X1 port map( I => n24816, ZN => n18217);
   U21656 : INV_X1 port map( I => n24403, ZN => n12240);
   U21657 : NAND2_X1 port map( A1 => n317, A2 => n15880, ZN => n14139);
   U21659 : INV_X1 port map( I => n25584, ZN => n18196);
   U21661 : NOR2_X1 port map( A1 => n10755, A2 => n14752, ZN => n24912);
   U21662 : NAND2_X1 port map( A1 => n25258, A2 => n17273, ZN => n14511);
   U21663 : NOR2_X1 port map( A1 => n14960, A2 => n8622, ZN => n16383);
   U21665 : NAND2_X1 port map( A1 => n18151, A2 => n28096, ZN => n15185);
   U21666 : NOR2_X1 port map( A1 => n1209, A2 => n32897, ZN => n25496);
   U21667 : INV_X1 port map( I => n25058, ZN => n25050);
   U21673 : NAND2_X1 port map( A1 => n25705, A2 => n11944, ZN => n13359);
   U21675 : AOI21_X1 port map( A1 => n32856, A2 => n25615, B => n9982, ZN => 
                           n25618);
   U21677 : INV_X1 port map( I => n25224, ZN => n25225);
   U21679 : NAND2_X1 port map( A1 => n14780, A2 => n26447, ZN => n12215);
   U21681 : NAND2_X1 port map( A1 => n25605, A2 => n831, ZN => n13996);
   U21685 : OAI21_X1 port map( A1 => n24911, A2 => n10755, B => n14752, ZN => 
                           n24906);
   U21688 : NAND2_X1 port map( A1 => n25861, A2 => n18022, ZN => n18020);
   U21689 : OAI21_X1 port map( A1 => n25052, A2 => n28070, B => n17744, ZN => 
                           n17743);
   U21690 : NAND2_X1 port map( A1 => n15479, A2 => n15478, ZN => n25356);
   U21693 : AOI21_X1 port map( A1 => n3843, A2 => n24965, B => n13627, ZN => 
                           n12202);
   U21694 : AOI21_X1 port map( A1 => n28736, A2 => n14810, B => n28200, ZN => 
                           n12250);
   U21695 : OAI21_X1 port map( A1 => n14634, A2 => n14638, B => n1420, ZN => 
                           n14633);
   U21696 : NAND2_X1 port map( A1 => n27183, A2 => n1074, ZN => n17708);
   U21699 : NAND2_X1 port map( A1 => n25516, A2 => n32897, ZN => n16468);
   U21702 : INV_X1 port map( I => n24447, ZN => n25705);
   U21704 : XOR2_X1 port map( A1 => Plaintext(145), A2 => Key(145), Z => n11905
                           );
   U21706 : INV_X1 port map( I => n21305, ZN => n21131);
   U21708 : AND2_X1 port map( A1 => n22664, A2 => n14307, Z => n11928);
   U21711 : AND2_X1 port map( A1 => n3843, A2 => n24965, Z => n11939);
   U21714 : AND2_X1 port map( A1 => n25705, A2 => n25707, Z => n11951);
   U21715 : OR2_X1 port map( A1 => n20039, A2 => n20040, Z => n11952);
   U21719 : OR2_X1 port map( A1 => n20411, A2 => n28261, Z => n11964);
   U21721 : NOR2_X1 port map( A1 => n13894, A2 => n13893, ZN => n11980);
   U21723 : XNOR2_X1 port map( A1 => n20822, A2 => n13093, ZN => n11982);
   U21724 : INV_X1 port map( I => n19355, ZN => n15842);
   U21727 : OR2_X1 port map( A1 => n24610, A2 => n680, Z => n11994);
   U21728 : XNOR2_X1 port map( A1 => n33293, A2 => n25827, ZN => n11996);
   U21729 : AND2_X1 port map( A1 => n25884, A2 => n25872, Z => n11999);
   U21733 : NOR2_X1 port map( A1 => n24112, A2 => n24289, ZN => n12002);
   U21737 : XNOR2_X1 port map( A1 => n23430, A2 => n25224, ZN => n12014);
   U21738 : AND2_X1 port map( A1 => n27166, A2 => n13622, Z => n12016);
   U21739 : AND2_X1 port map( A1 => n781, A2 => n1351, Z => n12021);
   U21740 : AND2_X1 port map( A1 => n969, A2 => n24194, Z => n12022);
   U21741 : AND2_X1 port map( A1 => n16933, A2 => n21249, Z => n12029);
   U21742 : AND2_X1 port map( A1 => n16413, A2 => n11944, Z => n12030);
   U21743 : NAND3_X1 port map( A1 => n16688, A2 => n1096, A3 => n24218, ZN => 
                           n24043);
   U21747 : OR2_X2 port map( A1 => n12384, A2 => n12382, Z => n12048);
   U21750 : OR2_X1 port map( A1 => n14458, A2 => n31017, Z => n12053);
   U21756 : XNOR2_X1 port map( A1 => n31499, A2 => n24417, ZN => n12059);
   U21757 : XNOR2_X1 port map( A1 => n17145, A2 => n22041, ZN => n12062);
   U21758 : AND2_X1 port map( A1 => n15909, A2 => n18757, Z => n12065);
   U21759 : INV_X1 port map( I => n25916, ZN => n25926);
   U21761 : INV_X1 port map( I => n16778, ZN => n25400);
   U21765 : INV_X1 port map( I => n22412, ZN => n22639);
   U21766 : XNOR2_X1 port map( A1 => n22029, A2 => n25722, ZN => n12082);
   U21770 : INV_X1 port map( I => n11944, ZN => n25706);
   U21775 : INV_X1 port map( I => n24168, ZN => n24194);
   U21777 : XNOR2_X1 port map( A1 => n22034, A2 => n22035, ZN => n12101);
   U21778 : INV_X1 port map( I => n23639, ZN => n23873);
   U21779 : XNOR2_X1 port map( A1 => n8298, A2 => n23436, ZN => n12104);
   U21784 : INV_X1 port map( I => n23132, ZN => n14464);
   U21789 : AND2_X1 port map( A1 => n23487, A2 => n23486, Z => n12122);
   U21790 : INV_X1 port map( I => n18973, ZN => n19271);
   U21791 : XNOR2_X1 port map( A1 => n15130, A2 => n25086, ZN => n12123);
   U21792 : XNOR2_X1 port map( A1 => n34078, A2 => n16551, ZN => n12124);
   U21795 : XNOR2_X1 port map( A1 => n22130, A2 => n24869, ZN => n12127);
   U21798 : XNOR2_X1 port map( A1 => n19736, A2 => n24968, ZN => n12136);
   U21799 : XNOR2_X1 port map( A1 => n19566, A2 => n16523, ZN => n12137);
   U21802 : AND2_X1 port map( A1 => n20456, A2 => n14086, Z => n12139);
   U21804 : INV_X1 port map( I => n13401, ZN => n21059);
   U21805 : XNOR2_X1 port map( A1 => n19630, A2 => n25476, ZN => n12141);
   U21806 : INV_X1 port map( I => n27698, ZN => n19808);
   U21809 : INV_X2 port map( I => n16682, ZN => n22634);
   U21810 : INV_X1 port map( I => n16587, ZN => n15566);
   U21811 : INV_X1 port map( I => n8548, ZN => n17723);
   U21813 : INV_X1 port map( I => n25545, ZN => n15816);
   U21815 : INV_X1 port map( I => n16687, ZN => n17986);
   U21816 : INV_X1 port map( I => n25864, ZN => n18019);
   U21817 : INV_X1 port map( I => n16550, ZN => n13394);
   U21818 : INV_X1 port map( I => n8487, ZN => n16438);
   U21821 : INV_X1 port map( I => n16698, ZN => n14648);
   U21822 : INV_X1 port map( I => n16507, ZN => n13091);
   U21824 : INV_X1 port map( I => n16597, ZN => n16038);
   U21826 : INV_X1 port map( I => n25086, ZN => n13331);
   U21827 : INV_X1 port map( I => n24962, ZN => n15415);
   U21828 : INV_X1 port map( I => n16533, ZN => n18102);
   U21829 : INV_X2 port map( I => n13567, ZN => n15255);
   U21834 : INV_X2 port map( I => n16310, ZN => n17813);
   U21835 : NAND2_X1 port map( A1 => n27651, A2 => n25119, ZN => n12163);
   U21836 : XNOR2_X1 port map( A1 => Plaintext(164), A2 => Key(164), ZN => 
                           n12166);
   U21837 : XOR2_X1 port map( A1 => n20983, A2 => n12171, Z => n12170);
   U21838 : XOR2_X1 port map( A1 => n20758, A2 => n20621, Z => n12172);
   U21839 : XNOR2_X1 port map( A1 => n18083, A2 => n19374, ZN => n12182);
   U21840 : XOR2_X1 port map( A1 => n4975, A2 => n32367, Z => n19751);
   U21841 : NAND2_X1 port map( A1 => n17525, A2 => n1850, ZN => n18132);
   U21843 : XOR2_X1 port map( A1 => n14841, A2 => n14136, Z => n12185);
   U21846 : XOR2_X1 port map( A1 => n23391, A2 => n25911, Z => n12200);
   U21850 : NAND2_X1 port map( A1 => n28263, A2 => n28669, ZN => n12209);
   U21852 : XOR2_X1 port map( A1 => n12223, A2 => n12410, Z => n12409);
   U21854 : NOR2_X1 port map( A1 => n22590, A2 => n12236, ZN => n17584);
   U21855 : XOR2_X1 port map( A1 => n22028, A2 => n16548, Z => n16816);
   U21857 : XOR2_X1 port map( A1 => n24741, A2 => n12240, Z => n12239);
   U21858 : NAND2_X2 port map( A1 => n14674, A2 => n14673, ZN => n21726);
   U21860 : XOR2_X1 port map( A1 => n12252, A2 => n25252, Z => n18108);
   U21861 : XOR2_X1 port map( A1 => n12252, A2 => n14583, Z => n14582);
   U21872 : XOR2_X1 port map( A1 => n19764, A2 => n17600, Z => n12283);
   U21873 : XOR2_X1 port map( A1 => n12286, A2 => n12285, Z => n12284);
   U21874 : XOR2_X1 port map( A1 => n5348, A2 => n24953, Z => n12285);
   U21875 : XOR2_X1 port map( A1 => n28813, A2 => n12494, Z => n12286);
   U21877 : XOR2_X1 port map( A1 => n23279, A2 => n23278, Z => n12288);
   U21879 : NAND2_X1 port map( A1 => n28450, A2 => n15864, ZN => n14524);
   U21880 : NAND2_X1 port map( A1 => n534, A2 => n28450, ZN => n21873);
   U21882 : AND2_X1 port map( A1 => n12085, A2 => n15057, Z => n12300);
   U21884 : NAND3_X2 port map( A1 => n19955, A2 => n19956, A3 => n19954, ZN => 
                           n14858);
   U21885 : NAND2_X2 port map( A1 => n12616, A2 => n12553, ZN => n16173);
   U21887 : XOR2_X1 port map( A1 => n12313, A2 => n27125, Z => n16972);
   U21888 : NOR2_X1 port map( A1 => n25676, A2 => n12314, ZN => n25677);
   U21891 : NOR2_X1 port map( A1 => n12315, A2 => n15456, ZN => n15729);
   U21892 : NAND3_X1 port map( A1 => n12727, A2 => n22715, A3 => n12315, ZN => 
                           n22717);
   U21893 : OAI21_X1 port map( A1 => n18727, A2 => n11123, B => n18726, ZN => 
                           n18729);
   U21897 : NAND2_X1 port map( A1 => n12325, A2 => n21400, ZN => n21096);
   U21901 : MUX2_X1 port map( I0 => n32900, I1 => n12329, S => n10822, Z => 
                           n25081);
   U21904 : XOR2_X1 port map( A1 => n11324, A2 => n12387, Z => n12331);
   U21905 : INV_X2 port map( I => n12960, ZN => n16375);
   U21913 : XOR2_X1 port map( A1 => n21007, A2 => n27169, Z => n13395);
   U21916 : NAND2_X2 port map( A1 => n14990, A2 => n22833, ZN => n16799);
   U21917 : XOR2_X1 port map( A1 => n24422, A2 => n24215, Z => n12355);
   U21918 : XNOR2_X1 port map( A1 => n24522, A2 => n24618, ZN => n24422);
   U21920 : NAND2_X1 port map( A1 => n26516, A2 => n30146, ZN => n23659);
   U21921 : INV_X2 port map( I => n15518, ZN => n25891);
   U21924 : XOR2_X1 port map( A1 => n12376, A2 => n25131, Z => n21050);
   U21927 : XOR2_X1 port map( A1 => n19723, A2 => n19667, Z => n12380);
   U21928 : XOR2_X1 port map( A1 => n19584, A2 => n13682, Z => n12381);
   U21929 : AOI21_X1 port map( A1 => n27131, A2 => n12383, B => n19274, ZN => 
                           n12382);
   U21930 : NAND2_X1 port map( A1 => n19318, A2 => n19275, ZN => n12383);
   U21932 : INV_X1 port map( I => n12390, ZN => n12392);
   U21934 : NOR2_X1 port map( A1 => n20105, A2 => n12398, ZN => n20454);
   U21936 : NOR2_X1 port map( A1 => n14913, A2 => n33295, ZN => n12402);
   U21937 : MUX2_X1 port map( I0 => n24086, I1 => n24085, S => n14913, Z => 
                           n12403);
   U21940 : XOR2_X1 port map( A1 => n19577, A2 => n19380, Z => n12411);
   U21949 : XOR2_X1 port map( A1 => n12456, A2 => n1413, Z => Ciphertext(63));
   U21951 : XOR2_X1 port map( A1 => n12462, A2 => n612, Z => n12461);
   U21952 : XOR2_X1 port map( A1 => n4057, A2 => n32695, Z => n12462);
   U21953 : XOR2_X1 port map( A1 => n30489, A2 => n4295, Z => n21898);
   U21961 : XOR2_X1 port map( A1 => n13814, A2 => n1198, Z => n12475);
   U21962 : XOR2_X1 port map( A1 => n12944, A2 => n12942, Z => n25188);
   U21963 : INV_X2 port map( I => n22638, ZN => n22636);
   U21965 : XOR2_X1 port map( A1 => n5381, A2 => n12491, Z => n22948);
   U21967 : XOR2_X1 port map( A1 => n12493, A2 => n24966, Z => n24389);
   U21968 : XOR2_X1 port map( A1 => n12494, A2 => n25098, Z => n20684);
   U21969 : XOR2_X1 port map( A1 => n12494, A2 => n25549, Z => n20971);
   U21972 : AOI21_X1 port map( A1 => n827, A2 => n32485, B => n12502, ZN => 
                           n19346);
   U21976 : INV_X2 port map( I => n17074, ZN => n24466);
   U21977 : XOR2_X1 port map( A1 => n13849, A2 => n12513, Z => n12512);
   U21985 : NAND2_X1 port map( A1 => n12169, A2 => n12541, ZN => n12540);
   U21987 : NOR2_X2 port map( A1 => n24114, A2 => n16356, ZN => n23608);
   U21990 : XOR2_X1 port map( A1 => n348, A2 => n24386, Z => n12552);
   U21996 : MUX2_X1 port map( I0 => n32397, I1 => n12561, S => n21646, Z => 
                           n15748);
   U22002 : XOR2_X1 port map( A1 => n12573, A2 => n13932, Z => n13931);
   U22006 : INV_X2 port map( I => n12584, ZN => n21305);
   U22008 : NAND2_X1 port map( A1 => n1175, A2 => n12585, ZN => n16591);
   U22009 : NOR2_X1 port map( A1 => n25961, A2 => n12585, ZN => n16361);
   U22017 : XOR2_X1 port map( A1 => n12610, A2 => n25191, Z => n19380);
   U22021 : NAND2_X1 port map( A1 => n16603, A2 => n23886, ZN => n12615);
   U22025 : OAI21_X1 port map( A1 => n4016, A2 => n14194, B => n19348, ZN => 
                           n19000);
   U22026 : XOR2_X1 port map( A1 => n702, A2 => n17430, Z => n12620);
   U22029 : XOR2_X1 port map( A1 => n24836, A2 => n24764, Z => n12628);
   U22033 : XOR2_X1 port map( A1 => n24750, A2 => n16602, Z => n12636);
   U22036 : OAI21_X2 port map( A1 => n13891, A2 => n13890, B => n13889, ZN => 
                           n19408);
   U22040 : NOR2_X1 port map( A1 => n13210, A2 => n949, ZN => n12649);
   U22048 : XOR2_X1 port map( A1 => n17912, A2 => n12665, Z => n24625);
   U22050 : XOR2_X1 port map( A1 => n20959, A2 => n12673, Z => n12672);
   U22051 : XOR2_X1 port map( A1 => n12675, A2 => n27423, Z => n13519);
   U22054 : INV_X1 port map( I => n23905, ZN => n16238);
   U22055 : OR2_X1 port map( A1 => n14974, A2 => n12680, Z => n15943);
   U22058 : NAND2_X2 port map( A1 => n25871, A2 => n25885, ZN => n12699);
   U22059 : NAND3_X1 port map( A1 => n941, A2 => n821, A3 => n17608, ZN => 
                           n12704);
   U22061 : NOR2_X2 port map( A1 => n18920, A2 => n18921, ZN => n12707);
   U22063 : XOR2_X1 port map( A1 => n13844, A2 => n26002, Z => n12717);
   U22064 : XOR2_X1 port map( A1 => n12721, A2 => n16482, Z => n20797);
   U22065 : XOR2_X1 port map( A1 => n12721, A2 => n16507, Z => n20915);
   U22066 : NAND3_X1 port map( A1 => n22715, A2 => n851, A3 => n12729, ZN => 
                           n22716);
   U22067 : OAI21_X1 port map( A1 => n22807, A2 => n12729, B => n16458, ZN => 
                           n15101);
   U22068 : XOR2_X1 port map( A1 => n12731, A2 => n20774, Z => n21375);
   U22069 : XOR2_X1 port map( A1 => n20772, A2 => n12732, Z => n12731);
   U22073 : NOR2_X2 port map( A1 => n21386, A2 => n21385, ZN => n21630);
   U22075 : XOR2_X1 port map( A1 => n9145, A2 => n31687, Z => n24792);
   U22076 : INV_X2 port map( I => n12735, ZN => n18110);
   U22078 : XOR2_X1 port map( A1 => n23155, A2 => n23414, Z => n23537);
   U22079 : NAND2_X1 port map( A1 => n6842, A2 => n12747, ZN => n21069);
   U22081 : XOR2_X1 port map( A1 => n20995, A2 => n17793, Z => n12749);
   U22082 : XOR2_X1 port map( A1 => n4728, A2 => n16527, Z => n15573);
   U22083 : NAND3_X1 port map( A1 => n16699, A2 => n19335, A3 => n14597, ZN => 
                           n12755);
   U22085 : XOR2_X1 port map( A1 => n22189, A2 => n22056, Z => n12760);
   U22087 : XOR2_X1 port map( A1 => n34120, A2 => n23425, Z => n12765);
   U22094 : NOR2_X2 port map( A1 => n17378, A2 => n17379, ZN => n13627);
   U22095 : NAND2_X1 port map( A1 => n21642, A2 => n29234, ZN => n21473);
   U22096 : XOR2_X1 port map( A1 => n12800, A2 => n16548, Z => n24354);
   U22097 : XOR2_X1 port map( A1 => n12795, A2 => n12057, Z => n15237);
   U22100 : XOR2_X1 port map( A1 => Plaintext(169), A2 => Key(169), Z => n15966
                           );
   U22101 : XOR2_X1 port map( A1 => n15913, A2 => n19514, Z => n12803);
   U22103 : NAND2_X1 port map( A1 => n12812, A2 => n29069, ZN => n18270);
   U22106 : OAI21_X2 port map( A1 => n12432, A2 => n12816, B => n14942, ZN => 
                           n24164);
   U22107 : NAND2_X2 port map( A1 => n6072, A2 => n1125, ZN => n22439);
   U22108 : XOR2_X1 port map( A1 => n12821, A2 => n25131, Z => n17500);
   U22115 : NOR2_X1 port map( A1 => n12587, A2 => n30291, ZN => n21606);
   U22116 : NOR2_X1 port map( A1 => n2575, A2 => n30291, ZN => n21759);
   U22119 : XOR2_X1 port map( A1 => n30171, A2 => n24943, Z => n15993);
   U22120 : OR2_X1 port map( A1 => n15022, A2 => n21761, Z => n12853);
   U22121 : AOI21_X2 port map( A1 => n12855, A2 => n26386, B => n21606, ZN => 
                           n21952);
   U22122 : INV_X2 port map( I => n23579, ZN => n23833);
   U22123 : OR2_X1 port map( A1 => n24219, A2 => n16554, Z => n12861);
   U22124 : XOR2_X1 port map( A1 => Plaintext(45), A2 => Key(45), Z => n18777);
   U22125 : XOR2_X1 port map( A1 => n28977, A2 => n27125, Z => n13741);
   U22126 : XOR2_X1 port map( A1 => n20730, A2 => n20842, Z => n20732);
   U22131 : XOR2_X1 port map( A1 => n14215, A2 => n19559, Z => n12896);
   U22136 : XOR2_X1 port map( A1 => n24761, A2 => n16584, Z => n12905);
   U22137 : XOR2_X1 port map( A1 => n23517, A2 => n12955, Z => n12954);
   U22138 : INV_X1 port map( I => n12907, ZN => n12908);
   U22141 : XOR2_X1 port map( A1 => n12915, A2 => n13529, Z => n21965);
   U22142 : XOR2_X1 port map( A1 => n20704, A2 => n12916, Z => n20931);
   U22143 : XOR2_X1 port map( A1 => n20768, A2 => n20703, Z => n12916);
   U22145 : XOR2_X1 port map( A1 => Plaintext(121), A2 => Key(121), Z => n14409
                           );
   U22146 : XOR2_X1 port map( A1 => n24793, A2 => n12918, Z => n14065);
   U22147 : OAI21_X1 port map( A1 => n16600, A2 => n2217, B => n6660, ZN => 
                           n12919);
   U22150 : XOR2_X1 port map( A1 => n23529, A2 => n12922, Z => n12921);
   U22154 : XOR2_X1 port map( A1 => n24473, A2 => n18042, Z => n12936);
   U22157 : XOR2_X1 port map( A1 => n24838, A2 => n12943, Z => n12942);
   U22159 : XOR2_X1 port map( A1 => n24835, A2 => n24834, Z => n12944);
   U22160 : XOR2_X1 port map( A1 => n11751, A2 => n12945, Z => n24835);
   U22163 : NAND3_X1 port map( A1 => n30375, A2 => n20028, A3 => n28423, ZN => 
                           n19905);
   U22164 : MUX2_X1 port map( I0 => n19805, I1 => n19806, S => n19724, Z => 
                           n19807);
   U22165 : AOI21_X1 port map( A1 => n30271, A2 => n13846, B => n27687, ZN => 
                           n18390);
   U22167 : XOR2_X1 port map( A1 => n23262, A2 => n23444, Z => n12955);
   U22168 : NOR2_X1 port map( A1 => n12956, A2 => n18848, ZN => n18593);
   U22169 : NOR2_X1 port map( A1 => n12956, A2 => n17184, ZN => n18594);
   U22170 : OAI21_X1 port map( A1 => n15967, A2 => n12956, B => n18846, ZN => 
                           n18734);
   U22171 : NAND2_X1 port map( A1 => n31972, A2 => n10283, ZN => n18870);
   U22173 : XOR2_X1 port map( A1 => n12957, A2 => n24426, Z => n13404);
   U22174 : XOR2_X1 port map( A1 => n20720, A2 => n12957, Z => n20721);
   U22175 : XOR2_X1 port map( A1 => n23438, A2 => n12934, Z => n23283);
   U22177 : XOR2_X1 port map( A1 => n12959, A2 => n18072, Z => n12958);
   U22178 : XOR2_X1 port map( A1 => n28908, A2 => n25541, Z => n12959);
   U22179 : XOR2_X1 port map( A1 => n22000, A2 => n22002, Z => n12962);
   U22182 : XOR2_X1 port map( A1 => n32648, A2 => n20905, Z => n13179);
   U22184 : XOR2_X1 port map( A1 => n27211, A2 => n12969, Z => n12971);
   U22186 : NOR2_X1 port map( A1 => n12973, A2 => n28869, ZN => n21121);
   U22188 : AOI21_X1 port map( A1 => n7203, A2 => n33295, B => n24139, ZN => 
                           n12985);
   U22191 : INV_X2 port map( I => n13177, ZN => n21095);
   U22192 : NAND3_X1 port map( A1 => n19255, A2 => n19143, A3 => n19252, ZN => 
                           n12993);
   U22193 : NOR2_X2 port map( A1 => n19791, A2 => n19790, ZN => n20582);
   U22196 : NOR2_X1 port map( A1 => n9484, A2 => n868, ZN => n13880);
   U22198 : XOR2_X1 port map( A1 => n19676, A2 => n29515, Z => n19677);
   U22199 : XOR2_X1 port map( A1 => n33749, A2 => n29515, Z => n19377);
   U22201 : INV_X2 port map( I => n13022, ZN => n17731);
   U22203 : NAND2_X1 port map( A1 => n18738, A2 => n18737, ZN => n13024);
   U22204 : NOR2_X1 port map( A1 => n2378, A2 => n13032, ZN => n24446);
   U22205 : NAND2_X1 port map( A1 => n15155, A2 => n13032, ZN => n25714);
   U22208 : XOR2_X1 port map( A1 => n20820, A2 => n13041, Z => n17576);
   U22209 : XOR2_X1 port map( A1 => n13041, A2 => n25079, Z => n20988);
   U22214 : XOR2_X1 port map( A1 => n13065, A2 => n16662, Z => Ciphertext(66));
   U22215 : INV_X1 port map( I => n13067, ZN => n15795);
   U22216 : NOR2_X1 port map( A1 => n3880, A2 => n24084, ZN => n16100);
   U22217 : AND2_X1 port map( A1 => n3880, A2 => n16286, Z => n15010);
   U22220 : INV_X1 port map( I => n22303, ZN => n13075);
   U22221 : NOR2_X1 port map( A1 => n18781, A2 => n10080, ZN => n13076);
   U22223 : INV_X2 port map( I => n13080, ZN => n17711);
   U22226 : XOR2_X1 port map( A1 => n24524, A2 => n13086, Z => n13085);
   U22228 : NOR2_X1 port map( A1 => n20439, A2 => n14863, ZN => n13090);
   U22229 : XOR2_X1 port map( A1 => n13106, A2 => n13095, Z => n19554);
   U22232 : XOR2_X1 port map( A1 => n19379, A2 => n24065, Z => n13099);
   U22233 : NAND2_X1 port map( A1 => n8412, A2 => n24271, ZN => n15899);
   U22234 : NOR2_X1 port map( A1 => n23555, A2 => n23806, ZN => n17701);
   U22237 : NAND2_X1 port map( A1 => n32874, A2 => n25795, ZN => n15304);
   U22238 : NAND2_X1 port map( A1 => n15242, A2 => n1009, ZN => n15676);
   U22239 : NAND2_X1 port map( A1 => n17467, A2 => n27382, ZN => n20932);
   U22244 : OAI21_X1 port map( A1 => n14312, A2 => n10700, B => n15143, ZN => 
                           n17617);
   U22250 : NOR2_X1 port map( A1 => n19874, A2 => n20092, ZN => n15383);
   U22251 : NAND2_X1 port map( A1 => n16957, A2 => n28763, ZN => n17038);
   U22252 : OAI21_X1 port map( A1 => n20065, A2 => n16630, B => n10413, ZN => 
                           n15311);
   U22255 : NOR3_X1 port map( A1 => n834, A2 => n25865, A3 => n29063, ZN => 
                           n14872);
   U22258 : NAND2_X1 port map( A1 => n23889, A2 => n23888, ZN => n17257);
   U22267 : BUF_X2 port map( I => n19618, Z => n20154);
   U22271 : OAI21_X1 port map( A1 => n16694, A2 => n13852, B => n19863, ZN => 
                           n17061);
   U22272 : NAND2_X1 port map( A1 => n14960, A2 => n13627, ZN => n13935);
   U22273 : NAND2_X1 port map( A1 => n8919, A2 => n14845, ZN => n15699);
   U22275 : NAND2_X1 port map( A1 => n953, A2 => n17649, ZN => n17736);
   U22276 : NAND2_X1 port map( A1 => n21713, A2 => n727, ZN => n21478);
   U22283 : NOR2_X1 port map( A1 => n22468, A2 => n15089, ZN => n15939);
   U22286 : NAND2_X1 port map( A1 => n23822, A2 => n23942, ZN => n13668);
   U22289 : INV_X1 port map( I => n23933, ZN => n13102);
   U22290 : OAI21_X1 port map( A1 => n28010, A2 => n4194, B => n16181, ZN => 
                           n13111);
   U22291 : NAND2_X1 port map( A1 => n338, A2 => n16987, ZN => n21844);
   U22292 : NOR2_X2 port map( A1 => n13265, A2 => n20934, ZN => n13114);
   U22293 : OAI21_X1 port map( A1 => n17644, A2 => n29523, B => n13115, ZN => 
                           n21591);
   U22298 : XOR2_X1 port map( A1 => n600, A2 => n20700, Z => n13122);
   U22299 : XNOR2_X1 port map( A1 => n17871, A2 => n30322, ZN => n13123);
   U22300 : NAND2_X1 port map( A1 => n29270, A2 => n13125, ZN => n23642);
   U22301 : AOI21_X1 port map( A1 => n16431, A2 => n13125, B => n354, ZN => 
                           n16281);
   U22306 : NAND2_X1 port map( A1 => n12871, A2 => n17074, ZN => n24606);
   U22309 : NOR2_X2 port map( A1 => n17935, A2 => n16818, ZN => n23003);
   U22317 : XOR2_X1 port map( A1 => n20753, A2 => n13179, Z => n13178);
   U22320 : XOR2_X1 port map( A1 => n20786, A2 => n16655, Z => n13181);
   U22324 : MUX2_X1 port map( I0 => n13186, I1 => n13185, S => n900, Z => 
                           n17249);
   U22330 : XOR2_X1 port map( A1 => n30273, A2 => n13209, Z => n13208);
   U22331 : XOR2_X1 port map( A1 => n23464, A2 => n23414, Z => n13214);
   U22334 : XOR2_X1 port map( A1 => n2073, A2 => n16555, Z => n13222);
   U22338 : XOR2_X1 port map( A1 => n23497, A2 => n23180, Z => n13234);
   U22340 : XOR2_X1 port map( A1 => n23181, A2 => n17934, Z => n13235);
   U22346 : MUX2_X1 port map( I0 => n14756, I1 => n842, S => n299, Z => n13261)
                           ;
   U22358 : XOR2_X1 port map( A1 => n16175, A2 => n17998, Z => n13293);
   U22359 : XOR2_X1 port map( A1 => n20972, A2 => n20971, Z => n13294);
   U22361 : NAND2_X2 port map( A1 => n14521, A2 => n23959, ZN => n16868);
   U22362 : XOR2_X1 port map( A1 => n27151, A2 => n2864, Z => n13299);
   U22363 : NAND2_X2 port map( A1 => n13302, A2 => n13301, ZN => n14980);
   U22364 : XOR2_X1 port map( A1 => n33150, A2 => n16612, Z => n13303);
   U22369 : NOR2_X1 port map( A1 => n9191, A2 => n30313, ZN => n13312);
   U22370 : NAND3_X1 port map( A1 => n17985, A2 => n30313, A3 => n18035, ZN => 
                           n13313);
   U22372 : INV_X2 port map( I => n18110, ZN => n13319);
   U22374 : NAND2_X1 port map( A1 => n10700, A2 => n25968, ZN => n17510);
   U22376 : NAND2_X1 port map( A1 => n13329, A2 => n8787, ZN => n13328);
   U22377 : NAND3_X1 port map( A1 => n16066, A2 => n27500, A3 => n794, ZN => 
                           n23609);
   U22380 : XOR2_X1 port map( A1 => n13336, A2 => n21028, Z => n17440);
   U22384 : AOI21_X2 port map( A1 => n23222, A2 => n23223, B => n23221, ZN => 
                           n24276);
   U22391 : XOR2_X1 port map( A1 => n19445, A2 => n15117, Z => n19373);
   U22393 : XOR2_X1 port map( A1 => n20960, A2 => n13357, Z => n14930);
   U22403 : XOR2_X1 port map( A1 => n6462, A2 => n15779, Z => n15778);
   U22404 : XOR2_X1 port map( A1 => n13375, A2 => n13372, Z => n17768);
   U22405 : XOR2_X1 port map( A1 => n13373, A2 => n13374, Z => n13372);
   U22406 : XOR2_X1 port map( A1 => n15183, A2 => n16674, Z => n13373);
   U22407 : XOR2_X1 port map( A1 => n13638, A2 => n27613, Z => n13374);
   U22409 : XOR2_X1 port map( A1 => n16053, A2 => n25195, Z => n13388);
   U22410 : XOR2_X1 port map( A1 => n28262, A2 => n13394, Z => n13393);
   U22412 : XOR2_X1 port map( A1 => n13405, A2 => n13404, Z => n13403);
   U22413 : XOR2_X1 port map( A1 => n20996, A2 => n14858, Z => n13405);
   U22414 : INV_X1 port map( I => n13407, ZN => n21416);
   U22415 : INV_X2 port map( I => n12317, ZN => n18785);
   U22419 : XOR2_X1 port map( A1 => n24403, A2 => n13419, Z => n23551);
   U22420 : NOR2_X1 port map( A1 => n17339, A2 => n27033, ZN => n19126);
   U22421 : NOR2_X1 port map( A1 => n17339, A2 => n32414, ZN => n18985);
   U22423 : NOR2_X1 port map( A1 => n17382, A2 => n15719, ZN => n17770);
   U22424 : NOR2_X1 port map( A1 => n17382, A2 => n14454, ZN => n13429);
   U22426 : XOR2_X1 port map( A1 => n13439, A2 => n13441, Z => n16777);
   U22427 : XOR2_X1 port map( A1 => n19546, A2 => n13440, Z => n13439);
   U22428 : XOR2_X1 port map( A1 => n13826, A2 => n25064, Z => n13440);
   U22430 : XOR2_X1 port map( A1 => n19463, A2 => n19772, Z => n19545);
   U22439 : XOR2_X1 port map( A1 => n13454, A2 => n13453, Z => n13452);
   U22440 : XOR2_X1 port map( A1 => n33468, A2 => n4295, Z => n13454);
   U22442 : OR2_X1 port map( A1 => n23975, A2 => n23976, Z => n13459);
   U22444 : NOR2_X1 port map( A1 => n8320, A2 => n13483, ZN => n25544);
   U22446 : NAND3_X1 port map( A1 => n24059, A2 => n14501, A3 => n13394, ZN => 
                           n13467);
   U22447 : INV_X1 port map( I => n13469, ZN => n13468);
   U22448 : AOI21_X1 port map( A1 => n14501, A2 => n24059, B => n13394, ZN => 
                           n13469);
   U22452 : XOR2_X1 port map( A1 => n16060, A2 => n25648, Z => n21938);
   U22457 : NAND2_X1 port map( A1 => n950, A2 => n19116, ZN => n13494);
   U22458 : XOR2_X1 port map( A1 => n13498, A2 => n23450, Z => n13497);
   U22462 : XOR2_X1 port map( A1 => n22264, A2 => n25218, Z => n22265);
   U22463 : XOR2_X1 port map( A1 => n22264, A2 => n25693, Z => n14979);
   U22470 : XOR2_X1 port map( A1 => n23300, A2 => n23299, Z => n13517);
   U22471 : NAND2_X2 port map( A1 => n22054, A2 => n22053, ZN => n23300);
   U22474 : XOR2_X1 port map( A1 => n13527, A2 => n13394, Z => Ciphertext(124))
                           ;
   U22475 : AOI21_X1 port map( A1 => n25556, A2 => n33414, B => n16853, ZN => 
                           n13528);
   U22476 : INV_X1 port map( I => n25542, ZN => n25556);
   U22477 : XOR2_X1 port map( A1 => n30331, A2 => n14526, Z => n13529);
   U22479 : XOR2_X1 port map( A1 => n32871, A2 => n13545, Z => n24637);
   U22480 : XOR2_X1 port map( A1 => n24421, A2 => n13545, Z => n24415);
   U22483 : NOR2_X1 port map( A1 => n17328, A2 => n20563, ZN => n20564);
   U22487 : NAND2_X1 port map( A1 => n13558, A2 => n22971, ZN => n22972);
   U22489 : OAI21_X1 port map( A1 => n2635, A2 => n13558, B => n13191, ZN => 
                           n15753);
   U22490 : NAND2_X1 port map( A1 => n23106, A2 => n13558, ZN => n22804);
   U22493 : XOR2_X1 port map( A1 => n32084, A2 => n13564, Z => n22178);
   U22495 : XOR2_X1 port map( A1 => n13586, A2 => n24532, Z => n17309);
   U22496 : XOR2_X1 port map( A1 => n30795, A2 => n13586, Z => n24828);
   U22497 : XOR2_X1 port map( A1 => n25969, A2 => n24869, Z => n13590);
   U22498 : NOR2_X1 port map( A1 => n11198, A2 => n13591, ZN => n17155);
   U22500 : XOR2_X1 port map( A1 => n24830, A2 => n25506, Z => n13595);
   U22501 : XOR2_X1 port map( A1 => n15588, A2 => n24815, Z => n13596);
   U22502 : XOR2_X1 port map( A1 => n24513, A2 => n24512, Z => n24815);
   U22506 : XOR2_X1 port map( A1 => n13606, A2 => n16613, Z => n20864);
   U22507 : XOR2_X1 port map( A1 => n13606, A2 => n1431, Z => n15652);
   U22508 : NAND2_X2 port map( A1 => n13609, A2 => n13608, ZN => n20158);
   U22511 : NOR2_X1 port map( A1 => n24965, A2 => n13627, ZN => n17331);
   U22512 : INV_X2 port map( I => n15514, ZN => n14133);
   U22514 : NAND2_X1 port map( A1 => n19824, A2 => n1165, ZN => n19825);
   U22519 : XOR2_X1 port map( A1 => Plaintext(117), A2 => Key(117), Z => n13719
                           );
   U22522 : NOR2_X1 port map( A1 => n13319, A2 => n21167, ZN => n13680);
   U22523 : XOR2_X1 port map( A1 => n13681, A2 => n1434, Z => n15793);
   U22524 : XOR2_X1 port map( A1 => n32367, A2 => n25864, Z => n13682);
   U22529 : XOR2_X1 port map( A1 => n19384, A2 => n17091, Z => n13689);
   U22542 : NAND2_X1 port map( A1 => n30682, A2 => n19048, ZN => n19016);
   U22544 : AOI21_X1 port map( A1 => n13736, A2 => n24970, B => n13934, ZN => 
                           n13735);
   U22545 : NAND2_X1 port map( A1 => n32493, A2 => n992, ZN => n22436);
   U22546 : XOR2_X1 port map( A1 => n11862, A2 => n25619, Z => n13740);
   U22547 : XOR2_X1 port map( A1 => n968, A2 => n15161, Z => n13742);
   U22550 : XOR2_X1 port map( A1 => n24770, A2 => n24993, Z => n13745);
   U22556 : OAI21_X1 port map( A1 => n31921, A2 => n29539, B => n13763, ZN => 
                           n16188);
   U22557 : NAND3_X1 port map( A1 => n17177, A2 => n19866, A3 => n1395, ZN => 
                           n13765);
   U22558 : INV_X1 port map( I => n13767, ZN => n13766);
   U22559 : AOI21_X1 port map( A1 => n17177, A2 => n19866, B => n1395, ZN => 
                           n13767);
   U22562 : AND2_X1 port map( A1 => n13785, A2 => n13537, Z => n13784);
   U22566 : XOR2_X1 port map( A1 => n24783, A2 => n24668, Z => n13794);
   U22568 : INV_X2 port map( I => n17047, ZN => n25334);
   U22569 : MUX2_X1 port map( I0 => n33110, I1 => n33583, S => n31807, Z => 
                           n23222);
   U22571 : NOR2_X1 port map( A1 => n31716, A2 => n17189, ZN => n13809);
   U22572 : XOR2_X1 port map( A1 => n32753, A2 => n26931, Z => n22131);
   U22573 : MUX2_X1 port map( I0 => n23624, I1 => n23625, S => n791, Z => 
                           n23627);
   U22574 : XOR2_X1 port map( A1 => n17188, A2 => n24964, Z => n13812);
   U22575 : XOR2_X1 port map( A1 => n8347, A2 => n19718, Z => n15557);
   U22576 : XOR2_X1 port map( A1 => n13817, A2 => n19411, Z => n15679);
   U22577 : XOR2_X1 port map( A1 => n32271, A2 => n13826, Z => n19430);
   U22586 : INV_X1 port map( I => n15139, ZN => n13845);
   U22589 : XOR2_X1 port map( A1 => n19405, A2 => n13854, Z => n13853);
   U22590 : XNOR2_X1 port map( A1 => n19658, A2 => n19461, ZN => n19405);
   U22591 : XOR2_X1 port map( A1 => n19574, A2 => n19480, Z => n13855);
   U22592 : XOR2_X1 port map( A1 => n16727, A2 => n19353, Z => n19480);
   U22596 : OR2_X1 port map( A1 => n22721, A2 => n28849, Z => n13861);
   U22599 : OAI22_X1 port map( A1 => n15655, A2 => n920, B1 => n27024, B2 => 
                           n13872, ZN => n21275);
   U22601 : XOR2_X1 port map( A1 => n16891, A2 => n13877, Z => n13876);
   U22602 : XOR2_X1 port map( A1 => n27423, A2 => n25929, Z => n13877);
   U22604 : AND2_X1 port map( A1 => n25542, A2 => n31236, Z => n13883);
   U22607 : XOR2_X1 port map( A1 => n5348, A2 => n20825, Z => n20799);
   U22608 : XOR2_X1 port map( A1 => n20764, A2 => n13887, Z => n13886);
   U22609 : XOR2_X1 port map( A1 => n20843, A2 => n25074, Z => n13887);
   U22610 : XOR2_X1 port map( A1 => Plaintext(63), A2 => Key(63), Z => n16596);
   U22611 : INV_X1 port map( I => n13895, ZN => n13893);
   U22613 : XOR2_X1 port map( A1 => n28687, A2 => n25190, Z => n13898);
   U22615 : XOR2_X1 port map( A1 => n21009, A2 => n20924, Z => n13901);
   U22616 : XOR2_X1 port map( A1 => n13902, A2 => n12797, Z => Ciphertext(185))
                           ;
   U22618 : XOR2_X1 port map( A1 => n27252, A2 => n25182, Z => n13907);
   U22619 : XOR2_X1 port map( A1 => n14908, A2 => n4157, Z => n13909);
   U22623 : XOR2_X1 port map( A1 => n27481, A2 => n16322, Z => n13927);
   U22624 : XOR2_X1 port map( A1 => n23271, A2 => n23291, Z => n13928);
   U22627 : INV_X2 port map( I => n13931, ZN => n23855);
   U22631 : INV_X1 port map( I => n13944, ZN => n15946);
   U22633 : XOR2_X1 port map( A1 => n22108, A2 => n25224, Z => n13956);
   U22634 : NAND2_X1 port map( A1 => n8371, A2 => n14334, ZN => n19811);
   U22639 : NOR2_X1 port map( A1 => n14392, A2 => n22791, ZN => n22759);
   U22644 : NOR3_X1 port map( A1 => n17066, A2 => n17065, A3 => n17068, ZN => 
                           n17067);
   U22646 : NAND3_X1 port map( A1 => n25613, A2 => n11931, A3 => n9982, ZN => 
                           n25609);
   U22650 : NAND3_X1 port map( A1 => n16783, A2 => n25561, A3 => n16704, ZN => 
                           n13979);
   U22655 : XOR2_X1 port map( A1 => n22202, A2 => n22146, Z => n15686);
   U22656 : XOR2_X1 port map( A1 => n22284, A2 => n18113, Z => n15548);
   U22659 : NOR2_X1 port map( A1 => n25254, A2 => n17273, ZN => n15094);
   U22664 : NAND2_X1 port map( A1 => n21866, A2 => n21736, ZN => n16235);
   U22665 : OAI21_X1 port map( A1 => n21189, A2 => n21321, B => n14023, ZN => 
                           n14022);
   U22666 : OAI21_X1 port map( A1 => n25808, A2 => n25811, B => n14009, ZN => 
                           n25810);
   U22674 : OR2_X1 port map( A1 => n20099, A2 => n19990, Z => n14019);
   U22675 : XOR2_X1 port map( A1 => n19596, A2 => n19595, Z => n19601);
   U22678 : NAND2_X2 port map( A1 => n21191, A2 => n14022, ZN => n21872);
   U22680 : XOR2_X1 port map( A1 => n14908, A2 => n16110, Z => n14916);
   U22688 : XOR2_X1 port map( A1 => n22169, A2 => n21924, Z => n17919);
   U22691 : NAND3_X1 port map( A1 => n25773, A2 => n25788, A3 => n25796, ZN => 
                           n25768);
   U22693 : NOR2_X1 port map( A1 => n10364, A2 => n18662, ZN => n17910);
   U22696 : XOR2_X1 port map( A1 => n14043, A2 => n14494, Z => n17518);
   U22697 : XOR2_X1 port map( A1 => n618, A2 => n21661, Z => n14043);
   U22699 : OR2_X1 port map( A1 => n30949, A2 => n23938, Z => n15238);
   U22700 : XOR2_X1 port map( A1 => n15612, A2 => n23374, Z => n23936);
   U22701 : INV_X2 port map( I => n15613, ZN => n23533);
   U22703 : NAND2_X1 port map( A1 => n20609, A2 => n20608, ZN => n14050);
   U22704 : NAND2_X1 port map( A1 => n20610, A2 => n33397, ZN => n14051);
   U22705 : XOR2_X1 port map( A1 => n28262, A2 => n2616, Z => n20639);
   U22706 : XOR2_X1 port map( A1 => n14053, A2 => n4047, Z => n15099);
   U22708 : NAND2_X1 port map( A1 => n828, A2 => n18774, ZN => n14056);
   U22713 : XOR2_X1 port map( A1 => n14070, A2 => n25274, Z => Ciphertext(86));
   U22721 : AND2_X1 port map( A1 => n19243, A2 => n877, Z => n14699);
   U22723 : NAND2_X1 port map( A1 => n16156, A2 => n11774, ZN => n14100);
   U22725 : XOR2_X1 port map( A1 => n16128, A2 => n24696, Z => n24697);
   U22729 : INV_X2 port map( I => n18090, ZN => n20113);
   U22733 : XNOR2_X1 port map( A1 => n15787, A2 => n19654, ZN => n18051);
   U22738 : OAI21_X1 port map( A1 => n29815, A2 => n16872, B => n16871, ZN => 
                           n16870);
   U22739 : OR3_X1 port map( A1 => n20335, A2 => n30130, A3 => n20158, Z => 
                           n20159);
   U22741 : XOR2_X1 port map( A1 => n14391, A2 => n19617, Z => n19618);
   U22742 : XOR2_X1 port map( A1 => n22137, A2 => n22138, Z => n22140);
   U22744 : AOI21_X1 port map( A1 => n22338, A2 => n906, B => n22645, ZN => 
                           n14145);
   U22746 : XOR2_X1 port map( A1 => n29876, A2 => n3727, Z => n14146);
   U22748 : NAND2_X1 port map( A1 => n1385, A2 => n18990, ZN => n14148);
   U22749 : NAND2_X1 port map( A1 => n25471, A2 => n25472, ZN => n14149);
   U22750 : INV_X1 port map( I => n25057, ZN => n25045);
   U22751 : OR2_X1 port map( A1 => n25058, A2 => n25057, Z => n25043);
   U22753 : AND2_X1 port map( A1 => n2061, A2 => n6533, Z => n14150);
   U22754 : XOR2_X1 port map( A1 => n17309, A2 => n24355, Z => n17308);
   U22756 : XOR2_X1 port map( A1 => n14370, A2 => n14154, Z => n23352);
   U22760 : NAND2_X2 port map( A1 => n14657, A2 => n14660, ZN => n19255);
   U22762 : NAND2_X1 port map( A1 => n28070, A2 => n25062, ZN => n17741);
   U22764 : XOR2_X1 port map( A1 => n20912, A2 => n20914, Z => n15035);
   U22766 : OR2_X1 port map( A1 => n5394, A2 => n20940, Z => n15925);
   U22769 : NAND3_X1 port map( A1 => n17403, A2 => n15134, A3 => n17402, ZN => 
                           n17401);
   U22771 : NOR2_X2 port map( A1 => n19912, A2 => n19913, ZN => n14187);
   U22774 : INV_X2 port map( I => n14190, ZN => n23871);
   U22776 : NAND2_X1 port map( A1 => n23876, A2 => n801, ZN => n16325);
   U22777 : NOR2_X1 port map( A1 => n24137, A2 => n15011, ZN => n14196);
   U22782 : XOR2_X1 port map( A1 => n24806, A2 => n14203, Z => n14202);
   U22783 : XOR2_X1 port map( A1 => n24764, A2 => n26000, Z => n14203);
   U22786 : XOR2_X1 port map( A1 => n19561, A2 => n25993, Z => n14211);
   U22795 : INV_X2 port map( I => n18763, ZN => n18768);
   U22797 : XOR2_X1 port map( A1 => n24648, A2 => n14578, Z => n14239);
   U22798 : XOR2_X1 port map( A1 => n29190, A2 => n19718, Z => n14242);
   U22799 : XOR2_X1 port map( A1 => n23376, A2 => n16373, Z => n23289);
   U22804 : NOR2_X1 port map( A1 => n14438, A2 => n32253, ZN => n14437);
   U22807 : XOR2_X1 port map( A1 => n28864, A2 => n20892, Z => n15525);
   U22808 : NAND3_X1 port map( A1 => n15073, A2 => n15074, A3 => n17986, ZN => 
                           n14257);
   U22809 : INV_X1 port map( I => n14259, ZN => n14258);
   U22813 : AND2_X1 port map( A1 => n1218, A2 => n25183, Z => n14276);
   U22814 : XOR2_X1 port map( A1 => n24762, A2 => n14279, Z => n14277);
   U22816 : XOR2_X1 port map( A1 => n33447, A2 => n24759, Z => n14279);
   U22818 : XOR2_X1 port map( A1 => n22180, A2 => n14299, Z => n14298);
   U22820 : XOR2_X1 port map( A1 => n14316, A2 => n14315, Z => n19532);
   U22824 : NAND2_X1 port map( A1 => n19078, A2 => n31254, ZN => n19079);
   U22825 : XOR2_X1 port map( A1 => n5772, A2 => n24962, Z => n21022);
   U22826 : XOR2_X1 port map( A1 => n5772, A2 => n25519, Z => n20914);
   U22827 : XOR2_X1 port map( A1 => n5772, A2 => n25827, Z => n20166);
   U22833 : XOR2_X1 port map( A1 => n14349, A2 => n23185, Z => n14348);
   U22834 : XOR2_X1 port map( A1 => n29462, A2 => n33293, Z => n14349);
   U22839 : XOR2_X1 port map( A1 => n14364, A2 => n14361, Z => n15294);
   U22840 : XOR2_X1 port map( A1 => n14362, A2 => n14363, Z => n14361);
   U22842 : XOR2_X1 port map( A1 => n24685, A2 => n24443, Z => n14364);
   U22843 : OR2_X1 port map( A1 => n20434, A2 => n20432, Z => n14368);
   U22844 : XOR2_X1 port map( A1 => n19624, A2 => n25549, Z => n17009);
   U22848 : XOR2_X1 port map( A1 => n33574, A2 => n17301, Z => n14385);
   U22849 : NAND2_X1 port map( A1 => n16554, A2 => n24219, ZN => n14444);
   U22850 : NAND2_X1 port map( A1 => n16554, A2 => n24218, ZN => n23602);
   U22854 : INV_X2 port map( I => n14409, ZN => n16249);
   U22856 : INV_X2 port map( I => n18429, ZN => n18822);
   U22857 : NOR2_X1 port map( A1 => n1245, A2 => n29634, ZN => n16800);
   U22858 : XOR2_X1 port map( A1 => n21726, A2 => n25079, Z => n14416);
   U22859 : XOR2_X1 port map( A1 => n22294, A2 => n22064, Z => n14422);
   U22860 : XOR2_X1 port map( A1 => n20225, A2 => n20226, Z => n14429);
   U22864 : XOR2_X1 port map( A1 => n27126, A2 => n13091, Z => n14435);
   U22867 : XOR2_X1 port map( A1 => n23488, A2 => n29299, Z => n14442);
   U22869 : NAND3_X1 port map( A1 => n30279, A2 => n714, A3 => n3232, ZN => 
                           n14607);
   U22875 : NAND2_X1 port map( A1 => n14451, A2 => n14450, ZN => n14449);
   U22877 : NAND2_X2 port map( A1 => n23571, A2 => n23572, ZN => n15663);
   U22882 : NAND3_X2 port map( A1 => n14472, A2 => n14471, A3 => n14470, ZN => 
                           n14682);
   U22884 : OR2_X1 port map( A1 => n14683, A2 => n1355, Z => n14472);
   U22885 : NAND2_X1 port map( A1 => n23643, A2 => n3760, ZN => n23644);
   U22886 : NAND2_X1 port map( A1 => n14478, A2 => n17163, ZN => n21979);
   U22890 : XOR2_X1 port map( A1 => n1261, A2 => n23203, Z => n14481);
   U22891 : XOR2_X1 port map( A1 => n23503, A2 => n16523, Z => n14492);
   U22893 : XOR2_X1 port map( A1 => n22197, A2 => n22239, Z => n21813);
   U22895 : XOR2_X1 port map( A1 => n14506, A2 => n14504, Z => n21869);
   U22896 : XOR2_X1 port map( A1 => n21838, A2 => n14505, Z => n14504);
   U22897 : XOR2_X1 port map( A1 => n22243, A2 => n27180, Z => n14505);
   U22898 : XOR2_X1 port map( A1 => n33969, A2 => n31513, Z => n14507);
   U22900 : NAND2_X1 port map( A1 => n25338, A2 => n14509, ZN => n25341);
   U22903 : XOR2_X1 port map( A1 => n14517, A2 => n14519, Z => n16845);
   U22904 : XOR2_X1 port map( A1 => n20827, A2 => n14930, Z => n14519);
   U22910 : INV_X2 port map( I => n14534, ZN => n14556);
   U22912 : XOR2_X1 port map( A1 => n29235, A2 => n24943, Z => n23316);
   U22918 : XOR2_X1 port map( A1 => n24809, A2 => n24417, Z => n14578);
   U22920 : XOR2_X1 port map( A1 => n23219, A2 => n14586, Z => n14580);
   U22921 : XOR2_X1 port map( A1 => n14584, A2 => n14582, Z => n14581);
   U22922 : XOR2_X1 port map( A1 => n23266, A2 => n25880, Z => n14586);
   U22923 : XOR2_X1 port map( A1 => n15374, A2 => n15372, Z => n15399);
   U22926 : XOR2_X1 port map( A1 => n28730, A2 => n1407, Z => n15900);
   U22927 : INV_X1 port map( I => n14717, ZN => n17225);
   U22929 : NAND2_X1 port map( A1 => n24154, A2 => n31883, ZN => n23117);
   U22931 : XOR2_X1 port map( A1 => n20917, A2 => n16642, Z => n14646);
   U22933 : AND2_X1 port map( A1 => n18638, A2 => n18539, Z => n14653);
   U22934 : INV_X2 port map( I => n14661, ZN => n16489);
   U22937 : NAND2_X1 port map( A1 => n31907, A2 => n14365, ZN => n20508);
   U22944 : XOR2_X1 port map( A1 => n14682, A2 => n16454, Z => n20810);
   U22945 : XOR2_X1 port map( A1 => n22123, A2 => n21952, Z => n14684);
   U22947 : XOR2_X1 port map( A1 => n21998, A2 => n21953, Z => n14685);
   U22954 : XOR2_X1 port map( A1 => n20794, A2 => n20793, Z => n14701);
   U22955 : NAND2_X2 port map( A1 => n18225, A2 => n18224, ZN => n16093);
   U22961 : NOR2_X1 port map( A1 => n16627, A2 => n11895, ZN => n14713);
   U22962 : XOR2_X1 port map( A1 => n12459, A2 => n7717, Z => n14716);
   U22965 : XOR2_X1 port map( A1 => n8491, A2 => n1396, Z => n15368);
   U22966 : OAI21_X1 port map( A1 => n20112, A2 => n20045, B => n16812, ZN => 
                           n17609);
   U22967 : XOR2_X1 port map( A1 => n23179, A2 => n24763, Z => n24634);
   U22968 : XOR2_X1 port map( A1 => n19537, A2 => n32046, Z => n14744);
   U22970 : XOR2_X1 port map( A1 => n23355, A2 => n7045, Z => n14748);
   U22973 : XOR2_X1 port map( A1 => n22196, A2 => n16631, Z => n14754);
   U22979 : XOR2_X1 port map( A1 => n23330, A2 => n14782, Z => n14781);
   U22980 : XOR2_X1 port map( A1 => n29299, A2 => n1410, Z => n14782);
   U22981 : XOR2_X1 port map( A1 => n23507, A2 => n23209, Z => n23330);
   U22982 : XOR2_X1 port map( A1 => n20776, A2 => n25319, Z => n14784);
   U22984 : XOR2_X1 port map( A1 => n22201, A2 => n16578, Z => n14787);
   U22985 : XOR2_X1 port map( A1 => n23437, A2 => n23329, Z => n14791);
   U22989 : NOR2_X1 port map( A1 => n32590, A2 => n14805, ZN => n16532);
   U22991 : XOR2_X1 port map( A1 => n21017, A2 => n20915, Z => n14809);
   U22992 : INV_X2 port map( I => n14814, ZN => n14815);
   U22995 : XOR2_X1 port map( A1 => n22139, A2 => n4342, Z => n16036);
   U22996 : XOR2_X1 port map( A1 => n14820, A2 => n15702, Z => n15701);
   U22998 : NAND2_X1 port map( A1 => n7486, A2 => n20555, ZN => n20297);
   U23002 : XOR2_X1 port map( A1 => Plaintext(95), A2 => Key(95), Z => n15955);
   U23005 : XOR2_X1 port map( A1 => n21913, A2 => n910, Z => n14833);
   U23007 : AND2_X1 port map( A1 => n19936, A2 => n14834, Z => n15382);
   U23010 : NAND3_X1 port map( A1 => n2551, A2 => n28395, A3 => n1647, ZN => 
                           n21724);
   U23012 : XOR2_X1 port map( A1 => n24504, A2 => n477, Z => n14842);
   U23014 : XOR2_X1 port map( A1 => n22238, A2 => n1404, Z => n21930);
   U23015 : XOR2_X1 port map( A1 => n22238, A2 => n16438, Z => n22041);
   U23016 : NOR2_X1 port map( A1 => n14863, A2 => n20494, ZN => n19804);
   U23018 : NOR2_X1 port map( A1 => n26585, A2 => n14863, ZN => n20437);
   U23020 : NOR2_X2 port map( A1 => n14866, A2 => n16469, ZN => n14865);
   U23022 : XOR2_X1 port map( A1 => n27179, A2 => n16550, Z => n15049);
   U23027 : XOR2_X1 port map( A1 => n24425, A2 => n14884, Z => n14883);
   U23028 : XOR2_X1 port map( A1 => n24813, A2 => n14885, Z => n14884);
   U23029 : XOR2_X1 port map( A1 => n14887, A2 => n17643, Z => n16938);
   U23030 : XOR2_X1 port map( A1 => n11668, A2 => n25126, Z => n23495);
   U23032 : OAI21_X1 port map( A1 => n14893, A2 => n14892, B => n100, ZN => 
                           n17810);
   U23033 : OR2_X1 port map( A1 => n21440, A2 => n8115, Z => n14896);
   U23034 : XOR2_X1 port map( A1 => Key(105), A2 => Plaintext(105), Z => n14898
                           );
   U23035 : INV_X2 port map( I => n14898, ZN => n16732);
   U23036 : XOR2_X1 port map( A1 => n14902, A2 => n21112, Z => n14901);
   U23038 : NOR2_X1 port map( A1 => n25863, A2 => n14915, ZN => n25861);
   U23044 : XOR2_X1 port map( A1 => n24790, A2 => n25161, Z => n14920);
   U23046 : XOR2_X1 port map( A1 => n24816, A2 => n28898, Z => n24818);
   U23049 : XOR2_X1 port map( A1 => n24473, A2 => n15674, Z => n14935);
   U23050 : XOR2_X1 port map( A1 => n17301, A2 => n14938, Z => n14937);
   U23051 : XOR2_X1 port map( A1 => n2896, A2 => n25324, Z => n17187);
   U23060 : NOR2_X1 port map( A1 => n19874, A2 => n14976, ZN => n16065);
   U23065 : NAND2_X1 port map( A1 => n13300, A2 => n1154, ZN => n20178);
   U23069 : XOR2_X1 port map( A1 => n19733, A2 => n19467, Z => n14985);
   U23071 : XOR2_X1 port map( A1 => n12594, A2 => n17063, Z => n16344);
   U23072 : XOR2_X1 port map( A1 => n12594, A2 => n25161, Z => n22233);
   U23073 : XOR2_X1 port map( A1 => n22251, A2 => n12594, Z => n22018);
   U23074 : XOR2_X1 port map( A1 => n23506, A2 => n23407, Z => n22387);
   U23075 : XOR2_X1 port map( A1 => n11370, A2 => n25126, Z => n24476);
   U23076 : XOR2_X1 port map( A1 => n156, A2 => n28411, Z => n14994);
   U23078 : NAND2_X1 port map( A1 => n1350, A2 => n15005, ZN => n20420);
   U23079 : NAND2_X1 port map( A1 => n20419, A2 => n1352, ZN => n15006);
   U23083 : NOR2_X1 port map( A1 => n15027, A2 => n20463, ZN => n20352);
   U23086 : XOR2_X1 port map( A1 => n19423, A2 => n24953, Z => n15031);
   U23088 : XOR2_X1 port map( A1 => n20911, A2 => n15037, Z => n15036);
   U23089 : XOR2_X1 port map( A1 => n3799, A2 => n348, Z => n15037);
   U23090 : XOR2_X1 port map( A1 => n20925, A2 => n591, Z => n15048);
   U23094 : XOR2_X1 port map( A1 => n29644, A2 => n16674, Z => n19669);
   U23099 : XOR2_X1 port map( A1 => n31584, A2 => n20872, Z => n15083);
   U23102 : XOR2_X1 port map( A1 => n19634, A2 => n19633, Z => n19635);
   U23104 : XOR2_X1 port map( A1 => n23138, A2 => n15099, Z => n16283);
   U23105 : OR2_X1 port map( A1 => n21963, A2 => n15103, Z => n22418);
   U23107 : XOR2_X1 port map( A1 => n15106, A2 => n16730, Z => n16711);
   U23109 : OR2_X1 port map( A1 => n19947, A2 => n19857, Z => n15111);
   U23110 : INV_X2 port map( I => n15115, ZN => n17598);
   U23111 : XOR2_X1 port map( A1 => Key(71), A2 => Plaintext(71), Z => n15115);
   U23113 : XOR2_X1 port map( A1 => n438, A2 => n16373, Z => n15121);
   U23115 : INV_X1 port map( I => n16676, ZN => n23612);
   U23117 : NAND2_X1 port map( A1 => n15124, A2 => n25251, ZN => n16582);
   U23119 : NAND2_X1 port map( A1 => n21719, A2 => n17227, ZN => n15127);
   U23124 : INV_X1 port map( I => Plaintext(101), ZN => n17548);
   U23128 : NAND2_X2 port map( A1 => n15140, A2 => n15196, ZN => n19115);
   U23136 : XOR2_X1 port map( A1 => n15153, A2 => n16753, Z => n16756);
   U23138 : NAND2_X1 port map( A1 => n25527, A2 => n28096, ZN => n15156);
   U23142 : NAND2_X1 port map( A1 => n20626, A2 => n14005, ZN => n15173);
   U23147 : NAND2_X1 port map( A1 => n21707, A2 => n21512, ZN => n21482);
   U23150 : INV_X1 port map( I => n21071, ZN => n21427);
   U23151 : INV_X1 port map( I => n16558, ZN => n22635);
   U23154 : XOR2_X1 port map( A1 => n1130, A2 => n21938, Z => n21940);
   U23156 : NAND2_X2 port map( A1 => n18143, A2 => n22499, ZN => n22955);
   U23158 : XOR2_X1 port map( A1 => Plaintext(87), A2 => Key(87), Z => n15194);
   U23163 : BUF_X4 port map( I => n24459, Z => n25582);
   U23164 : XOR2_X1 port map( A1 => n15205, A2 => n15701, Z => n20015);
   U23166 : XOR2_X1 port map( A1 => Plaintext(13), A2 => Key(13), Z => n16914);
   U23167 : AND2_X1 port map( A1 => n22984, A2 => n22985, Z => n15208);
   U23169 : XOR2_X1 port map( A1 => n16586, A2 => n11889, Z => n19502);
   U23173 : INV_X1 port map( I => Key(118), ZN => n16378);
   U23175 : NAND2_X1 port map( A1 => n20205, A2 => n8206, ZN => n18171);
   U23177 : INV_X2 port map( I => n15229, ZN => n18098);
   U23178 : NOR3_X1 port map( A1 => n26350, A2 => n10700, A3 => n14312, ZN => 
                           n18716);
   U23179 : NAND2_X1 port map( A1 => n21791, A2 => n21790, ZN => n21796);
   U23181 : NOR2_X1 port map( A1 => n24610, A2 => n680, ZN => n15231);
   U23182 : XOR2_X1 port map( A1 => Plaintext(161), A2 => Key(161), Z => n15347
                           );
   U23183 : NAND2_X2 port map( A1 => n17196, A2 => n17195, ZN => n25916);
   U23189 : INV_X2 port map( I => n15235, ZN => n16704);
   U23190 : NOR2_X1 port map( A1 => n15722, A2 => n15238, ZN => n17180);
   U23191 : MUX2_X1 port map( I0 => n23549, I1 => n23548, S => n16066, Z => 
                           n23550);
   U23192 : XOR2_X1 port map( A1 => n23512, A2 => n6901, Z => n15307);
   U23193 : XOR2_X1 port map( A1 => Key(107), A2 => Plaintext(107), Z => n15240
                           );
   U23199 : AND3_X1 port map( A1 => n21181, A2 => n21182, A3 => n4076, Z => 
                           n16282);
   U23201 : XOR2_X1 port map( A1 => n17141, A2 => n12101, Z => n17140);
   U23203 : INV_X1 port map( I => Plaintext(124), ZN => n17622);
   U23204 : XOR2_X1 port map( A1 => n19580, A2 => n27137, Z => n19582);
   U23207 : OAI21_X2 port map( A1 => n19623, A2 => n19622, B => n19621, ZN => 
                           n20310);
   U23208 : NAND3_X1 port map( A1 => n24878, A2 => n24877, A3 => n24876, ZN => 
                           n24880);
   U23210 : INV_X1 port map( I => n17525, ZN => n15274);
   U23211 : AND3_X1 port map( A1 => n24316, A2 => n16305, A3 => n26938, Z => 
                           n16304);
   U23214 : NAND2_X1 port map( A1 => n15413, A2 => n15412, ZN => n21483);
   U23219 : XNOR2_X1 port map( A1 => n31374, A2 => n25364, ZN => n17106);
   U23221 : XOR2_X1 port map( A1 => n15292, A2 => n25560, Z => Ciphertext(125))
                           ;
   U23222 : INV_X2 port map( I => n15294, ZN => n15295);
   U23224 : INV_X1 port map( I => n23282, ZN => n15305);
   U23228 : NOR2_X1 port map( A1 => n832, A2 => n27189, ZN => n25733);
   U23232 : XOR2_X1 port map( A1 => n24691, A2 => n12969, Z => n15334);
   U23236 : INV_X1 port map( I => n20851, ZN => n15337);
   U23238 : XOR2_X1 port map( A1 => n29190, A2 => n25364, Z => n23207);
   U23240 : XOR2_X1 port map( A1 => n23168, A2 => n15370, Z => n15346);
   U23241 : INV_X2 port map( I => n15347, ZN => n18720);
   U23242 : OR2_X1 port map( A1 => n18720, A2 => n16614, Z => n15348);
   U23244 : XOR2_X1 port map( A1 => n8491, A2 => n32813, Z => n15744);
   U23245 : XOR2_X1 port map( A1 => n11481, A2 => n30309, Z => n18190);
   U23246 : XOR2_X1 port map( A1 => n20183, A2 => n24991, Z => n15352);
   U23249 : INV_X1 port map( I => n15364, ZN => n22803);
   U23251 : XOR2_X1 port map( A1 => n23297, A2 => n16581, Z => n15370);
   U23252 : XOR2_X1 port map( A1 => n23150, A2 => n25669, Z => n15373);
   U23254 : XOR2_X1 port map( A1 => n17407, A2 => n24855, Z => n25201);
   U23257 : INV_X2 port map( I => n15384, ZN => n21923);
   U23259 : XOR2_X1 port map( A1 => n17918, A2 => n15386, Z => n17917);
   U23260 : XOR2_X1 port map( A1 => n22130, A2 => n25772, Z => n15386);
   U23266 : XOR2_X1 port map( A1 => n207, A2 => n15415, Z => n18105);
   U23268 : INV_X2 port map( I => n25710, ZN => n25760);
   U23269 : XOR2_X1 port map( A1 => n14428, A2 => n25500, Z => n21010);
   U23270 : XOR2_X1 port map( A1 => n5149, A2 => n15420, Z => n15419);
   U23271 : XOR2_X1 port map( A1 => n702, A2 => n16597, Z => n15420);
   U23272 : XOR2_X1 port map( A1 => n5482, A2 => n24527, Z => n21905);
   U23273 : INV_X1 port map( I => n15421, ZN => n22754);
   U23274 : MUX2_X1 port map( I0 => n23000, I1 => n13159, S => n15421, Z => 
                           n23006);
   U23279 : XOR2_X1 port map( A1 => n15432, A2 => n15431, Z => n15430);
   U23280 : XOR2_X1 port map( A1 => n16076, A2 => n16584, Z => n15431);
   U23284 : NAND2_X1 port map( A1 => n15442, A2 => n21239, ZN => n15441);
   U23286 : XOR2_X1 port map( A1 => n27151, A2 => n24809, Z => n15452);
   U23287 : XOR2_X1 port map( A1 => n21945, A2 => n25880, Z => n15460);
   U23292 : XOR2_X1 port map( A1 => n15329, A2 => n22970, Z => n23153);
   U23293 : XOR2_X1 port map( A1 => n23152, A2 => n23154, Z => n15470);
   U23294 : XOR2_X1 port map( A1 => n460, A2 => n15471, Z => n15472);
   U23296 : NAND2_X1 port map( A1 => n23855, A2 => n4177, ZN => n15475);
   U23298 : NAND2_X2 port map( A1 => n25336, A2 => n15480, ZN => n25368);
   U23301 : XOR2_X1 port map( A1 => n23399, A2 => n23217, Z => n15489);
   U23303 : INV_X2 port map( I => n15496, ZN => n15528);
   U23310 : XOR2_X1 port map( A1 => n23284, A2 => n23283, Z => n15515);
   U23311 : XOR2_X1 port map( A1 => n15517, A2 => n11370, Z => n15987);
   U23313 : XOR2_X1 port map( A1 => n15526, A2 => n15523, Z => n21233);
   U23314 : XOR2_X1 port map( A1 => n15525, A2 => n15524, Z => n15523);
   U23315 : XOR2_X1 port map( A1 => n20733, A2 => n25208, Z => n15524);
   U23318 : XOR2_X1 port map( A1 => n20975, A2 => n1070, Z => n15538);
   U23319 : XOR2_X1 port map( A1 => n15875, A2 => n15540, Z => n15539);
   U23320 : XOR2_X1 port map( A1 => n20821, A2 => n30303, Z => n15540);
   U23324 : XOR2_X1 port map( A1 => n24515, A2 => n24815, Z => n15543);
   U23328 : INV_X2 port map( I => n23352, ZN => n23764);
   U23331 : XOR2_X1 port map( A1 => n22062, A2 => n22060, Z => n15561);
   U23332 : XOR2_X1 port map( A1 => n21048, A2 => n31584, Z => n15562);
   U23333 : XOR2_X1 port map( A1 => n19513, A2 => n15566, Z => n15565);
   U23338 : NAND3_X2 port map( A1 => n15579, A2 => n21983, A3 => n15578, ZN => 
                           n23209);
   U23339 : XOR2_X1 port map( A1 => Plaintext(165), A2 => Key(165), Z => n17167
                           );
   U23340 : NOR2_X1 port map( A1 => n31533, A2 => n2928, ZN => n15590);
   U23341 : NAND2_X2 port map( A1 => n15594, A2 => n15592, ZN => n20395);
   U23342 : NOR2_X1 port map( A1 => n6842, A2 => n5480, ZN => n21244);
   U23343 : NAND2_X1 port map( A1 => n13506, A2 => n6842, ZN => n21633);
   U23348 : NAND2_X1 port map( A1 => n10183, A2 => n9234, ZN => n15644);
   U23351 : XOR2_X1 port map( A1 => n15668, A2 => n15667, Z => n15666);
   U23352 : XOR2_X1 port map( A1 => n20869, A2 => n21018, Z => n15667);
   U23354 : XOR2_X1 port map( A1 => n24816, A2 => n15671, Z => n24452);
   U23356 : INV_X2 port map( I => n16939, ZN => n16451);
   U23360 : INV_X2 port map( I => n18071, ZN => n18743);
   U23361 : XOR2_X1 port map( A1 => n15788, A2 => n19447, Z => n19449);
   U23363 : XOR2_X1 port map( A1 => n23210, A2 => n23212, Z => n15691);
   U23365 : XOR2_X1 port map( A1 => n15978, A2 => n25054, Z => n15702);
   U23367 : XOR2_X1 port map( A1 => n30183, A2 => n24839, Z => n15707);
   U23370 : XOR2_X1 port map( A1 => Plaintext(171), A2 => Key(171), Z => n17029
                           );
   U23374 : XOR2_X1 port map( A1 => n21994, A2 => n1398, Z => n15725);
   U23382 : INV_X2 port map( I => n15754, ZN => n25238);
   U23385 : XOR2_X1 port map( A1 => n32893, A2 => n1394, Z => n15761);
   U23386 : INV_X1 port map( I => n24823, ZN => n15765);
   U23387 : OAI21_X2 port map( A1 => n15896, A2 => n15771, B => n15769, ZN => 
                           n25258);
   U23392 : XOR2_X1 port map( A1 => n15792, A2 => n7511, Z => n15791);
   U23395 : XOR2_X1 port map( A1 => n10522, A2 => n15802, Z => n15801);
   U23398 : XOR2_X1 port map( A1 => n19703, A2 => n15816, Z => n15815);
   U23399 : XOR2_X1 port map( A1 => n15817, A2 => n20357, Z => n21225);
   U23402 : XOR2_X1 port map( A1 => n19483, A2 => n25879, Z => n15819);
   U23405 : XOR2_X1 port map( A1 => n22164, A2 => n15822, Z => n15821);
   U23407 : OR2_X1 port map( A1 => n21603, A2 => n31960, Z => n15828);
   U23408 : NOR2_X1 port map( A1 => n21629, A2 => n21630, ZN => n15840);
   U23409 : XOR2_X1 port map( A1 => n15861, A2 => n24644, Z => n15860);
   U23410 : XOR2_X1 port map( A1 => n25182, A2 => n12969, Z => n15861);
   U23419 : MUX2_X1 port map( I0 => n24256, I1 => n24255, S => n15876, Z => 
                           n24259);
   U23424 : XOR2_X1 port map( A1 => n15183, A2 => n16636, Z => n15886);
   U23425 : XNOR2_X1 port map( A1 => n5932, A2 => n6547, ZN => n15887);
   U23426 : XOR2_X1 port map( A1 => n21027, A2 => n15890, Z => n15889);
   U23427 : XOR2_X1 port map( A1 => n20641, A2 => n20921, Z => n15890);
   U23428 : XOR2_X1 port map( A1 => n20919, A2 => n20922, Z => n15891);
   U23429 : XOR2_X1 port map( A1 => n646, A2 => n23430, Z => n15897);
   U23431 : NAND3_X1 port map( A1 => n22754, A2 => n806, A3 => n13159, ZN => 
                           n22755);
   U23433 : XOR2_X1 port map( A1 => n19378, A2 => n27672, Z => n15904);
   U23434 : INV_X1 port map( I => n15909, ZN => n18762);
   U23435 : AOI21_X1 port map( A1 => n15909, A2 => n18499, B => n33472, ZN => 
                           n18503);
   U23436 : XOR2_X1 port map( A1 => Plaintext(69), A2 => Key(69), Z => n18498);
   U23437 : XOR2_X1 port map( A1 => n15913, A2 => n19602, Z => n19613);
   U23440 : INV_X1 port map( I => n15929, ZN => n17318);
   U23443 : XOR2_X1 port map( A1 => n24546, A2 => n545, Z => n15934);
   U23445 : NOR2_X1 port map( A1 => n19124, A2 => n8233, ZN => n19125);
   U23450 : NAND3_X1 port map( A1 => n25845, A2 => n25844, A3 => n25846, ZN => 
                           n15947);
   U23451 : XOR2_X1 port map( A1 => n24777, A2 => n15949, Z => n15948);
   U23452 : XOR2_X1 port map( A1 => n12969, A2 => n7511, Z => n15949);
   U23454 : XOR2_X1 port map( A1 => n15959, A2 => n16657, Z => Ciphertext(168))
                           ;
   U23455 : XOR2_X1 port map( A1 => n400, A2 => n25716, Z => n19376);
   U23456 : XOR2_X1 port map( A1 => n11891, A2 => n25208, Z => n15963);
   U23457 : XOR2_X1 port map( A1 => Plaintext(125), A2 => Key(125), Z => n17143
                           );
   U23458 : NOR2_X1 port map( A1 => n17184, A2 => n18845, ZN => n15967);
   U23459 : INV_X2 port map( I => n17029, ZN => n17184);
   U23461 : XOR2_X1 port map( A1 => n9327, A2 => n19507, Z => n19415);
   U23462 : XOR2_X1 port map( A1 => n22072, A2 => n34150, Z => n15969);
   U23463 : NAND2_X1 port map( A1 => n15976, A2 => n3183, ZN => n22051);
   U23466 : XOR2_X1 port map( A1 => n19408, A2 => n17551, Z => n15983);
   U23468 : XOR2_X1 port map( A1 => n15992, A2 => n15994, Z => n16129);
   U23469 : XOR2_X1 port map( A1 => n15993, A2 => n20902, Z => n15992);
   U23470 : XOR2_X1 port map( A1 => n21997, A2 => n15998, Z => n16000);
   U23471 : XOR2_X1 port map( A1 => n22030, A2 => n22305, Z => n15998);
   U23472 : XOR2_X1 port map( A1 => n21998, A2 => n21999, Z => n15999);
   U23473 : XOR2_X1 port map( A1 => n19378, A2 => n30411, Z => n16005);
   U23474 : XOR2_X1 port map( A1 => n23367, A2 => n23368, Z => n16010);
   U23477 : AOI22_X1 port map( A1 => n24615, A2 => n33434, B1 => n16383, B2 => 
                           n1208, ZN => n16021);
   U23478 : XOR2_X1 port map( A1 => n16302, A2 => n16997, Z => n16996);
   U23481 : XOR2_X1 port map( A1 => n16036, A2 => n17529, Z => n16035);
   U23482 : OAI21_X1 port map( A1 => n20608, A2 => n20606, B => n16481, ZN => 
                           n20368);
   U23487 : NAND2_X1 port map( A1 => n24912, A2 => n24911, ZN => n17883);
   U23489 : INV_X1 port map( I => n24144, ZN => n16039);
   U23491 : NAND2_X1 port map( A1 => n23815, A2 => n354, ZN => n23818);
   U23494 : XOR2_X1 port map( A1 => n322, A2 => n25669, Z => n17991);
   U23497 : AND2_X1 port map( A1 => n19614, A2 => n4587, Z => n19622);
   U23498 : INV_X2 port map( I => n16062, ZN => n25701);
   U23501 : XOR2_X1 port map( A1 => n19533, A2 => n19532, Z => n19833);
   U23512 : XOR2_X1 port map( A1 => n16104, A2 => n16697, Z => Ciphertext(46));
   U23518 : AOI21_X2 port map( A1 => n21156, A2 => n27543, B => n21155, ZN => 
                           n22072);
   U23519 : XNOR2_X1 port map( A1 => n19708, A2 => n24514, ZN => n18082);
   U23523 : NAND2_X1 port map( A1 => n11892, A2 => n11804, ZN => n17076);
   U23524 : XOR2_X1 port map( A1 => n28813, A2 => n25161, Z => n16773);
   U23526 : XOR2_X1 port map( A1 => n24695, A2 => n24357, Z => n16416);
   U23530 : OR2_X1 port map( A1 => n25912, A2 => n25922, Z => n25920);
   U23535 : OAI22_X1 port map( A1 => n18624, A2 => n16522, B1 => n828, B2 => 
                           n18623, ZN => n16156);
   U23539 : XOR2_X1 port map( A1 => n23363, A2 => n23535, Z => n16162);
   U23541 : AOI21_X1 port map( A1 => n25281, A2 => n733, B => n17876, ZN => 
                           n17875);
   U23544 : XOR2_X1 port map( A1 => n20907, A2 => n21036, Z => n16191);
   U23545 : INV_X1 port map( I => n15116, ZN => n23595);
   U23546 : XOR2_X1 port map( A1 => n21900, A2 => n21899, Z => n21901);
   U23553 : NAND2_X1 port map( A1 => n18785, A2 => n32108, ZN => n18367);
   U23555 : XOR2_X1 port map( A1 => n21923, A2 => n22012, Z => n21281);
   U23556 : INV_X2 port map( I => n16220, ZN => n16766);
   U23557 : XOR2_X1 port map( A1 => Plaintext(56), A2 => Key(56), Z => n16220);
   U23559 : XOR2_X1 port map( A1 => Plaintext(143), A2 => Key(143), Z => n18071
                           );
   U23561 : NAND2_X2 port map( A1 => n24709, A2 => n24708, ZN => n25820);
   U23563 : XOR2_X1 port map( A1 => n20930, A2 => n17106, Z => n17957);
   U23564 : XOR2_X1 port map( A1 => n16237, A2 => n30275, Z => n18149);
   U23565 : NAND2_X1 port map( A1 => n19089, A2 => n5760, ZN => n19090);
   U23572 : INV_X1 port map( I => n1053, ZN => n19361);
   U23574 : XOR2_X1 port map( A1 => n19689, A2 => n19690, Z => n19695);
   U23578 : INV_X2 port map( I => n16277, ZN => n22433);
   U23581 : XOR2_X1 port map( A1 => n16284, A2 => n16581, Z => Ciphertext(92));
   U23586 : INV_X1 port map( I => n22873, ZN => n22916);
   U23590 : XOR2_X1 port map( A1 => Plaintext(89), A2 => Key(89), Z => n16310);
   U23591 : OAI21_X1 port map( A1 => n25745, A2 => n25746, B => n25744, ZN => 
                           n25747);
   U23597 : XOR2_X1 port map( A1 => Key(81), A2 => Plaintext(81), Z => n18613);
   U23603 : NAND2_X1 port map( A1 => n21760, A2 => n21759, ZN => n21765);
   U23604 : INV_X1 port map( I => n19108, ZN => n18930);
   U23613 : INV_X1 port map( I => n29269, ZN => n23932);
   U23615 : XOR2_X1 port map( A1 => n16378, A2 => n18382, Z => n18818);
   U23616 : INV_X1 port map( I => n32874, ZN => n25773);
   U23617 : XOR2_X1 port map( A1 => n4400, A2 => n16081, Z => n19787);
   U23618 : XOR2_X1 port map( A1 => n17042, A2 => n17041, Z => n17119);
   U23625 : NAND2_X1 port map( A1 => n16412, A2 => n16411, ZN => n18169);
   U23630 : XOR2_X1 port map( A1 => n19628, A2 => n16437, Z => n19631);
   U23631 : XOR2_X1 port map( A1 => n29030, A2 => n16438, Z => n16437);
   U23632 : XOR2_X1 port map( A1 => n22154, A2 => n21884, Z => n16439);
   U23633 : XOR2_X1 port map( A1 => n7879, A2 => n25282, Z => n24769);
   U23634 : XOR2_X1 port map( A1 => n20984, A2 => n20593, Z => n20600);
   U23638 : XOR2_X1 port map( A1 => n16242, A2 => n21889, Z => n16457);
   U23642 : XOR2_X1 port map( A1 => n17434, A2 => n17435, Z => n20064);
   U23644 : OR2_X1 port map( A1 => n23753, A2 => n11922, Z => n23727);
   U23650 : BUF_X2 port map( I => n20015, Z => n16491);
   U23655 : NOR2_X1 port map( A1 => n18196, A2 => n18195, ZN => n18194);
   U23657 : XOR2_X1 port map( A1 => n26794, A2 => n16672, Z => n16513);
   U23661 : OR3_X1 port map( A1 => n1141, A2 => n29497, A3 => n929, Z => n17171
                           );
   U23665 : XOR2_X1 port map( A1 => n16541, A2 => n30993, Z => Ciphertext(147))
                           ;
   U23669 : AOI22_X1 port map( A1 => n21065, A2 => n29460, B1 => n21064, B2 => 
                           n28642, ZN => n16553);
   U23671 : XOR2_X1 port map( A1 => Plaintext(17), A2 => Key(17), Z => n18198);
   U23681 : NAND3_X1 port map( A1 => n25365, A2 => n750, A3 => n25366, ZN => 
                           n25372);
   U23692 : NAND2_X1 port map( A1 => n16937, A2 => n25322, ZN => n16660);
   U23699 : XOR2_X1 port map( A1 => n21997, A2 => n21920, Z => n17452);
   U23701 : XOR2_X1 port map( A1 => n16689, A2 => n22179, Z => n22589);
   U23703 : XOR2_X1 port map( A1 => n21951, A2 => n21949, Z => n16692);
   U23704 : INV_X2 port map( I => n16695, ZN => n18064);
   U23707 : XOR2_X1 port map( A1 => Plaintext(55), A2 => Key(55), Z => n16819);
   U23708 : BUF_X2 port map( I => Key(191), Z => n16703);
   U23709 : XOR2_X1 port map( A1 => n24768, A2 => n29274, Z => n16730);
   U23710 : INV_X2 port map( I => n16711, ZN => n25145);
   U23713 : XOR2_X1 port map( A1 => n12, A2 => n30301, Z => n16718);
   U23714 : NOR2_X1 port map( A1 => n11930, A2 => n16432, ZN => n16724);
   U23715 : XOR2_X1 port map( A1 => n19502, A2 => n19501, Z => n16734);
   U23717 : XOR2_X1 port map( A1 => n8109, A2 => n16738, Z => n16737);
   U23718 : XOR2_X1 port map( A1 => n18216, A2 => n24671, Z => n16739);
   U23724 : XOR2_X1 port map( A1 => n16754, A2 => n17576, Z => n16753);
   U23725 : INV_X2 port map( I => n16756, ZN => n21203);
   U23727 : XOR2_X1 port map( A1 => n17555, A2 => n16604, Z => n16767);
   U23733 : INV_X2 port map( I => n16776, ZN => n23575);
   U23734 : NAND2_X1 port map( A1 => n17079, A2 => n16780, ZN => n17982);
   U23735 : NAND2_X1 port map( A1 => n17079, A2 => n13401, ZN => n17983);
   U23739 : OAI21_X1 port map( A1 => n21259, A2 => n16652, B => n21257, ZN => 
                           n21260);
   U23741 : AND2_X1 port map( A1 => n16819, A2 => n16766, Z => n18486);
   U23742 : XOR2_X1 port map( A1 => n13602, A2 => n10766, Z => n16823);
   U23744 : XOR2_X1 port map( A1 => n28163, A2 => n16649, Z => n20827);
   U23745 : NAND2_X1 port map( A1 => n20325, A2 => n28011, ZN => n17514);
   U23748 : XOR2_X1 port map( A1 => n19550, A2 => n27137, Z => n16841);
   U23750 : XOR2_X1 port map( A1 => n19474, A2 => n16690, Z => n19475);
   U23751 : INV_X1 port map( I => n16448, ZN => n20821);
   U23753 : MUX2_X1 port map( I0 => n18943, I1 => n18944, S => n18995, Z => 
                           n18947);
   U23756 : XOR2_X1 port map( A1 => n11166, A2 => n22198, Z => n17258);
   U23757 : XOR2_X1 port map( A1 => n16869, A2 => n25545, Z => Ciphertext(121))
                           ;
   U23758 : NAND3_X1 port map( A1 => n1049, A2 => n29815, A3 => n19326, ZN => 
                           n16871);
   U23759 : AOI21_X1 port map( A1 => n20627, A2 => n7280, B => n14005, ZN => 
                           n16883);
   U23760 : INV_X2 port map( I => n16885, ZN => n22435);
   U23762 : XOR2_X1 port map( A1 => n17913, A2 => n17915, Z => n16887);
   U23765 : XOR2_X1 port map( A1 => Plaintext(75), A2 => Key(75), Z => n16899);
   U23766 : INV_X2 port map( I => n16899, ZN => n18774);
   U23768 : XOR2_X1 port map( A1 => n22015, A2 => n16911, Z => n16910);
   U23769 : INV_X2 port map( I => n16913, ZN => n18151);
   U23770 : NAND2_X2 port map( A1 => n16926, A2 => n16928, ZN => n23453);
   U23773 : XOR2_X1 port map( A1 => n26701, A2 => n24748, Z => n23279);
   U23776 : XOR2_X1 port map( A1 => n22013, A2 => n26000, Z => n16945);
   U23777 : XOR2_X1 port map( A1 => n22303, A2 => n21994, Z => n16946);
   U23783 : XOR2_X1 port map( A1 => n22141, A2 => n24231, Z => n16974);
   U23784 : INV_X2 port map( I => n16996, ZN => n20103);
   U23785 : XOR2_X1 port map( A1 => n19567, A2 => n12137, Z => n16997);
   U23787 : XOR2_X1 port map( A1 => n23440, A2 => n17013, Z => n17012);
   U23788 : XOR2_X1 port map( A1 => n10773, A2 => n16613, Z => n17013);
   U23791 : XOR2_X1 port map( A1 => n20722, A2 => n20724, Z => n17026);
   U23796 : XOR2_X1 port map( A1 => n24666, A2 => n17049, Z => n17048);
   U23797 : XOR2_X1 port map( A1 => n16128, A2 => n705, Z => n17049);
   U23798 : INV_X2 port map( I => n17050, ZN => n23735);
   U23802 : MUX2_X1 port map( I0 => n27143, I1 => n13896, S => n16072, Z => 
                           n21199);
   U23803 : XOR2_X1 port map( A1 => n29312, A2 => n16636, Z => n17072);
   U23804 : XOR2_X1 port map( A1 => Plaintext(88), A2 => Key(88), Z => n18569);
   U23806 : AOI21_X1 port map( A1 => n16337, A2 => n23763, B => n17087, ZN => 
                           n17086);
   U23807 : XOR2_X1 port map( A1 => n19698, A2 => n17091, Z => n17090);
   U23812 : OR2_X1 port map( A1 => n751, A2 => n25627, Z => n17108);
   U23814 : XOR2_X1 port map( A1 => n17115, A2 => n8139, Z => Ciphertext(16));
   U23818 : XOR2_X1 port map( A1 => n19766, A2 => n12103, Z => n17125);
   U23819 : INV_X2 port map( I => n17127, ZN => n19867);
   U23821 : XOR2_X1 port map( A1 => n5380, A2 => n1433, Z => n23340);
   U23822 : NAND2_X1 port map( A1 => n17134, A2 => n31959, ZN => n23542);
   U23823 : INV_X2 port map( I => n24726, ZN => n25885);
   U23828 : XOR2_X1 port map( A1 => n22067, A2 => n22198, Z => n17145);
   U23830 : NOR2_X1 port map( A1 => n27597, A2 => n10831, ZN => n17363);
   U23831 : MUX2_X1 port map( I0 => n19856, I1 => n17365, S => n10831, Z => 
                           n17364);
   U23832 : NAND2_X2 port map( A1 => n20189, A2 => n20191, ZN => n20531);
   U23833 : XOR2_X1 port map( A1 => n24518, A2 => n24444, Z => n17159);
   U23835 : NAND2_X1 port map( A1 => n6638, A2 => n12548, ZN => n17162);
   U23836 : OR2_X1 port map( A1 => n22636, A2 => n22637, Z => n17163);
   U23838 : XNOR2_X1 port map( A1 => Plaintext(90), A2 => Key(90), ZN => n17168
                           );
   U23839 : NAND3_X1 port map( A1 => n33972, A2 => n29497, A3 => n21414, ZN => 
                           n17172);
   U23841 : XOR2_X1 port map( A1 => n33572, A2 => n29951, Z => n17174);
   U23843 : XOR2_X1 port map( A1 => n22108, A2 => n22055, Z => n22152);
   U23844 : XOR2_X1 port map( A1 => n17188, A2 => n23413, Z => n23415);
   U23845 : XOR2_X1 port map( A1 => n17193, A2 => n17192, Z => n20133);
   U23847 : XOR2_X1 port map( A1 => n30305, A2 => n28806, Z => n19729);
   U23848 : NAND2_X1 port map( A1 => n25899, A2 => n18219, ZN => n17196);
   U23851 : XOR2_X1 port map( A1 => n30284, A2 => n17206, Z => n17205);
   U23852 : INV_X1 port map( I => n22029, ZN => n17206);
   U23853 : XOR2_X1 port map( A1 => n17207, A2 => n17258, Z => n22090);
   U23857 : OAI21_X2 port map( A1 => n21390, A2 => n17217, B => n17215, ZN => 
                           n21849);
   U23859 : XOR2_X1 port map( A1 => n4554, A2 => n23478, Z => n17235);
   U23860 : NAND2_X1 port map( A1 => n17237, A2 => n20401, ZN => n20574);
   U23861 : XOR2_X1 port map( A1 => n1004, A2 => n1306, Z => n17244);
   U23865 : INV_X2 port map( I => n17255, ZN => n17582);
   U23866 : XOR2_X1 port map( A1 => n21961, A2 => n21962, Z => n17259);
   U23872 : XOR2_X1 port map( A1 => n20668, A2 => n17282, Z => n17281);
   U23873 : XOR2_X1 port map( A1 => n21044, A2 => n20586, Z => n17282);
   U23875 : INV_X1 port map( I => n17289, ZN => n17290);
   U23876 : NAND2_X1 port map( A1 => n32063, A2 => n24955, ZN => n24957);
   U23881 : XOR2_X1 port map( A1 => n24674, A2 => n24429, Z => n17307);
   U23882 : NAND2_X1 port map( A1 => n24103, A2 => n17310, ZN => n23664);
   U23885 : XOR2_X1 port map( A1 => n24526, A2 => n16038, Z => n24542);
   U23886 : XOR2_X1 port map( A1 => n24526, A2 => n14648, Z => n24752);
   U23887 : AND2_X1 port map( A1 => n18965, A2 => n18955, Z => n17320);
   U23888 : NOR2_X2 port map( A1 => n19273, A2 => n19272, ZN => n19772);
   U23890 : XOR2_X1 port map( A1 => n30443, A2 => n17324, Z => n17323);
   U23891 : INV_X1 port map( I => n25827, ZN => n17324);
   U23894 : NOR2_X1 port map( A1 => n14312, A2 => n947, ZN => n18982);
   U23895 : XOR2_X1 port map( A1 => n29312, A2 => n16402, Z => n19750);
   U23896 : XNOR2_X1 port map( A1 => n23336, A2 => n23335, ZN => n23446);
   U23897 : XOR2_X1 port map( A1 => n17353, A2 => n23445, Z => n17351);
   U23899 : XOR2_X1 port map( A1 => n31908, A2 => n19342, Z => n17355);
   U23900 : XOR2_X1 port map( A1 => n19588, A2 => n19340, Z => n17356);
   U23902 : NOR2_X1 port map( A1 => n25590, A2 => n26912, ZN => n17367);
   U23904 : XOR2_X1 port map( A1 => n17380, A2 => n17381, Z => n20117);
   U23905 : XOR2_X1 port map( A1 => n19739, A2 => n12136, Z => n17381);
   U23906 : OR2_X1 port map( A1 => n25316, A2 => n1074, Z => n17383);
   U23907 : XOR2_X1 port map( A1 => n26582, A2 => n16642, Z => n18015);
   U23909 : NAND2_X1 port map( A1 => n25546, A2 => n25542, ZN => n17402);
   U23915 : AND2_X1 port map( A1 => n21349, A2 => n21348, Z => n17418);
   U23916 : NOR2_X1 port map( A1 => n17419, A2 => n18722, ZN => n18301);
   U23920 : XOR2_X1 port map( A1 => n17436, A2 => n19706, Z => n17435);
   U23921 : XOR2_X1 port map( A1 => n31450, A2 => n1191, Z => n17436);
   U23923 : INV_X4 port map( I => n18923, ZN => n17445);
   U23924 : MUX2_X1 port map( I0 => n18719, I1 => n18718, S => n18855, Z => 
                           n17446);
   U23925 : NAND2_X2 port map( A1 => n18734, A2 => n18735, ZN => n18980);
   U23926 : INV_X2 port map( I => n17450, ZN => n22332);
   U23928 : XOR2_X1 port map( A1 => n23168, A2 => n23167, Z => n17457);
   U23933 : XOR2_X1 port map( A1 => Key(0), A2 => Plaintext(0), Z => n18882);
   U23938 : XOR2_X1 port map( A1 => n6547, A2 => n16697, Z => n24375);
   U23939 : XOR2_X1 port map( A1 => n6547, A2 => n24839, Z => n24840);
   U23944 : XOR2_X1 port map( A1 => n22033, A2 => n22205, Z => n17529);
   U23953 : NAND2_X1 port map( A1 => n17630, A2 => n22472, ZN => n17567);
   U23954 : NAND3_X1 port map( A1 => n13746, A2 => n17569, A3 => n22472, ZN => 
                           n17568);
   U23955 : XOR2_X1 port map( A1 => n24597, A2 => n17571, Z => n17570);
   U23956 : XOR2_X1 port map( A1 => n24596, A2 => n24595, Z => n17572);
   U23960 : XOR2_X1 port map( A1 => Plaintext(44), A2 => Key(44), Z => n18076);
   U23961 : INV_X1 port map( I => n25911, ZN => n17600);
   U23962 : XOR2_X1 port map( A1 => n16319, A2 => n25519, Z => n18144);
   U23963 : XOR2_X1 port map( A1 => n16319, A2 => n30954, Z => n24451);
   U23964 : XOR2_X1 port map( A1 => n16319, A2 => n25324, Z => n24671);
   U23966 : XOR2_X1 port map( A1 => n12, A2 => n16423, Z => n24481);
   U23968 : XOR2_X1 port map( A1 => n19463, A2 => n19412, Z => n17613);
   U23972 : NOR2_X2 port map( A1 => n18741, A2 => n18740, ZN => n19262);
   U23976 : XOR2_X1 port map( A1 => n34120, A2 => n16671, Z => n17628);
   U23978 : NOR2_X1 port map( A1 => n25495, A2 => n30935, ZN => n25498);
   U23979 : OAI21_X1 port map( A1 => n25496, A2 => n30935, B => n17636, ZN => 
                           n25497);
   U23982 : XOR2_X1 port map( A1 => n20868, A2 => n20867, Z => n17643);
   U23984 : XNOR2_X1 port map( A1 => Plaintext(100), A2 => Key(100), ZN => 
                           n17649);
   U23985 : XOR2_X1 port map( A1 => n19730, A2 => n17651, Z => n17650);
   U23986 : XOR2_X1 port map( A1 => n19779, A2 => n25832, Z => n17651);
   U23988 : OR2_X1 port map( A1 => n20651, A2 => n23191, Z => n17658);
   U23989 : NOR2_X1 port map( A1 => n25057, A2 => n25058, ZN => n17744);
   U23992 : NOR2_X1 port map( A1 => n17675, A2 => n19794, ZN => n20209);
   U23993 : XOR2_X1 port map( A1 => n25249, A2 => n16548, Z => Ciphertext(78));
   U23994 : XOR2_X1 port map( A1 => n17679, A2 => n22032, Z => n22035);
   U23996 : INV_X2 port map( I => n17683, ZN => n25012);
   U23999 : XOR2_X1 port map( A1 => n27148, A2 => n27995, Z => n17704);
   U24001 : XOR2_X1 port map( A1 => n24646, A2 => n25457, Z => n17705);
   U24004 : NAND3_X1 port map( A1 => n6072, A2 => n32483, A3 => n22584, ZN => 
                           n17718);
   U24007 : XNOR2_X1 port map( A1 => n33373, A2 => n20699, ZN => n20868);
   U24009 : XOR2_X1 port map( A1 => n17738, A2 => n20675, Z => n21136);
   U24012 : OR2_X1 port map( A1 => n25059, A2 => n28070, Z => n17742);
   U24013 : XOR2_X1 port map( A1 => n17752, A2 => n17754, Z => n24368);
   U24014 : XOR2_X1 port map( A1 => n24673, A2 => n17755, Z => n17754);
   U24015 : XOR2_X1 port map( A1 => n24531, A2 => n24801, Z => n17755);
   U24016 : XOR2_X1 port map( A1 => n22165, A2 => n22163, Z => n17765);
   U24017 : INV_X2 port map( I => n17768, ZN => n23942);
   U24018 : NAND2_X1 port map( A1 => n17781, A2 => n15046, ZN => n17778);
   U24020 : NAND2_X1 port map( A1 => n17810, A2 => n945, ZN => n18897);
   U24026 : NAND2_X1 port map( A1 => n31533, A2 => n2928, ZN => n17809);
   U24027 : XOR2_X1 port map( A1 => n19637, A2 => n1366, Z => n19639);
   U24029 : NAND2_X1 port map( A1 => n28528, A2 => n17817, ZN => n18359);
   U24032 : XOR2_X1 port map( A1 => n15844, A2 => n29728, Z => n17834);
   U24033 : XOR2_X1 port map( A1 => n17837, A2 => n21035, Z => n20660);
   U24035 : XOR2_X1 port map( A1 => n17844, A2 => n25619, Z => Ciphertext(137))
                           ;
   U24037 : OR2_X1 port map( A1 => n25488, A2 => n25478, Z => n17850);
   U24043 : XOR2_X1 port map( A1 => n24687, A2 => n24688, Z => n17869);
   U24044 : XOR2_X1 port map( A1 => n17875, A2 => n27672, Z => Ciphertext(87));
   U24045 : NAND2_X1 port map( A1 => n23899, A2 => n4069, ZN => n17881);
   U24046 : OR2_X1 port map( A1 => n24908, A2 => n6154, Z => n17884);
   U24047 : INV_X2 port map( I => n17886, ZN => n24610);
   U24049 : INV_X2 port map( I => n17903, ZN => n25755);
   U24050 : XOR2_X1 port map( A1 => n24825, A2 => n24401, Z => n17904);
   U24052 : XNOR2_X1 port map( A1 => n17919, A2 => n17917, ZN => n17916);
   U24054 : XOR2_X1 port map( A1 => n17933, A2 => n293, Z => Ciphertext(74));
   U24055 : XOR2_X1 port map( A1 => n23259, A2 => n25856, Z => n17934);
   U24057 : XOR2_X1 port map( A1 => n24491, A2 => n18138, Z => n17938);
   U24061 : NOR2_X1 port map( A1 => n17948, A2 => n25446, ZN => n25424);
   U24065 : NAND2_X1 port map( A1 => n739, A2 => n23889, ZN => n17949);
   U24069 : XOR2_X1 port map( A1 => n14337, A2 => n26751, Z => n17958);
   U24072 : XOR2_X1 port map( A1 => Plaintext(134), A2 => Key(134), Z => n17970
                           );
   U24074 : AOI21_X1 port map( A1 => n31435, A2 => n3241, B => n28365, ZN => 
                           n17977);
   U24075 : NAND2_X1 port map( A1 => n23807, A2 => n23848, ZN => n17978);
   U24076 : XOR2_X1 port map( A1 => n25181, A2 => n25182, Z => Ciphertext(65));
   U24082 : XOR2_X1 port map( A1 => n20970, A2 => n32052, Z => n17998);
   U24083 : XOR2_X1 port map( A1 => n21040, A2 => n25009, Z => n18010);
   U24084 : XOR2_X1 port map( A1 => n28806, A2 => n24966, Z => n18011);
   U24086 : AND2_X1 port map( A1 => n22610, A2 => n22634, Z => n18013);
   U24089 : XOR2_X1 port map( A1 => n20957, A2 => n20682, Z => n18024);
   U24092 : XOR2_X1 port map( A1 => n19445, A2 => n24917, Z => n18031);
   U24093 : NAND2_X1 port map( A1 => n16345, A2 => n21463, ZN => n18034);
   U24095 : NOR2_X1 port map( A1 => n21812, A2 => n21811, ZN => n18043);
   U24103 : INV_X2 port map( I => n18075, ZN => n25198);
   U24105 : XNOR2_X1 port map( A1 => Plaintext(46), A2 => Key(46), ZN => n18085
                           );
   U24111 : XOR2_X1 port map( A1 => n18096, A2 => n20959, Z => n18095);
   U24112 : XOR2_X1 port map( A1 => n30163, A2 => n31233, Z => n18096);
   U24113 : XOR2_X1 port map( A1 => n23166, A2 => n18108, Z => n18107);
   U24115 : NAND2_X1 port map( A1 => n842, A2 => n667, ZN => n23629);
   U24117 : INV_X1 port map( I => n23079, ZN => n18129);
   U24118 : NAND2_X1 port map( A1 => n18827, A2 => n18489, ZN => n18130);
   U24119 : NOR2_X1 port map( A1 => n18146, A2 => n24197, ZN => n18145);
   U24120 : XOR2_X1 port map( A1 => n18149, A2 => n18148, Z => n21815);
   U24121 : XOR2_X1 port map( A1 => n22240, A2 => n16602, Z => n18148);
   U24122 : INV_X2 port map( I => n18155, ZN => n25119);
   U24124 : XOR2_X1 port map( A1 => n19619, A2 => n112, Z => n18165);
   U24125 : XOR2_X1 port map( A1 => n24513, A2 => n15742, Z => n18173);
   U24128 : OAI21_X1 port map( A1 => n4146, A2 => n25697, B => n25699, ZN => 
                           n18195);
   U24132 : XOR2_X1 port map( A1 => n322, A2 => n18217, Z => n18216);
   U24133 : INV_X2 port map( I => n18220, ZN => n24436);
   U24135 : XOR2_X1 port map( A1 => n29890, A2 => n19769, Z => n19770);
   U24137 : XOR2_X1 port map( A1 => n19741, A2 => n25161, Z => n18231);
   U24140 : NAND2_X1 port map( A1 => n19971, A2 => n18237, ZN => n18236);
   U24141 : NAND2_X1 port map( A1 => n19900, A2 => n19899, ZN => n18237);
   U24142 : XOR2_X1 port map( A1 => n18238, A2 => n19685, Z => n20108);
   U24143 : XOR2_X1 port map( A1 => n19681, A2 => n19680, Z => n18238);
   U24149 : XOR2_X1 port map( A1 => Plaintext(141), A2 => Key(141), Z => n18314
                           );
   U24152 : OAI22_X1 port map( A1 => n25248, A2 => n27429, B1 => n25247, B2 => 
                           n25246, ZN => n25249);
   U24156 : BUF_X2 port map( I => n18569, Z => n18493);
   U24158 : INV_X1 port map( I => n20616, ZN => n20363);
   U24161 : BUF_X2 port map( I => n21100, Z => n21307);
   U24163 : NAND4_X1 port map( A1 => n23998, A2 => n23997, A3 => n23922, A4 => 
                           n23921, ZN => n23934);
   U24166 : XOR2_X1 port map( A1 => Key(72), A2 => Plaintext(72), Z => n18773);
   U24167 : INV_X1 port map( I => n18773, ZN => n18770);
   U24168 : INV_X1 port map( I => Plaintext(59), ZN => n18275);
   U24169 : XOR2_X1 port map( A1 => n18275, A2 => Key(59), Z => n18763);
   U24171 : INV_X1 port map( I => Plaintext(64), ZN => n18280);
   U24172 : INV_X1 port map( I => Plaintext(62), ZN => n18281);
   U24173 : XOR2_X1 port map( A1 => n18281, A2 => Key(62), Z => n18780);
   U24174 : INV_X1 port map( I => Plaintext(80), ZN => n18282);
   U24175 : XOR2_X1 port map( A1 => n18282, A2 => Key(80), Z => n18283);
   U24176 : INV_X1 port map( I => Plaintext(66), ZN => n18286);
   U24177 : XOR2_X1 port map( A1 => n18286, A2 => Key(66), Z => n18756);
   U24178 : XOR2_X1 port map( A1 => Key(67), A2 => Plaintext(67), Z => n18335);
   U24180 : INV_X1 port map( I => Plaintext(68), ZN => n18287);
   U24181 : XOR2_X1 port map( A1 => n18287, A2 => Key(68), Z => n18293);
   U24182 : NAND2_X1 port map( A1 => n18338, A2 => n18605, ZN => n18294);
   U24183 : NAND2_X1 port map( A1 => n32437, A2 => n19108, ZN => n18297);
   U24186 : XOR2_X1 port map( A1 => Key(85), A2 => Plaintext(85), Z => n18323);
   U24189 : XOR2_X1 port map( A1 => Key(150), A2 => Plaintext(150), Z => n18540
                           );
   U24190 : XOR2_X1 port map( A1 => Key(155), A2 => Plaintext(155), Z => n18300
                           );
   U24191 : XOR2_X1 port map( A1 => Key(154), A2 => Plaintext(154), Z => n18580
                           );
   U24192 : XOR2_X1 port map( A1 => Key(152), A2 => Plaintext(152), Z => n18541
                           );
   U24193 : INV_X1 port map( I => n18302, ZN => n18304);
   U24195 : XOR2_X1 port map( A1 => Key(137), A2 => Plaintext(137), Z => n18310
                           );
   U24196 : INV_X1 port map( I => n18314, ZN => n18747);
   U24197 : INV_X1 port map( I => Plaintext(142), ZN => n18313);
   U24198 : XOR2_X1 port map( A1 => n18313, A2 => Key(142), Z => n18434);
   U24199 : XOR2_X1 port map( A1 => Key(139), A2 => Plaintext(139), Z => n18707
                           );
   U24200 : INV_X1 port map( I => Plaintext(130), ZN => n18315);
   U24201 : OAI21_X1 port map( A1 => n1439, A2 => n18317, B => n18316, ZN => 
                           n18320);
   U24202 : XOR2_X1 port map( A1 => Key(131), A2 => Plaintext(131), Z => n18392
                           );
   U24203 : MUX2_X1 port map( I0 => n18492, I1 => n18566, S => n18324, Z => 
                           n18327);
   U24205 : NOR2_X1 port map( A1 => n18328, A2 => n16564, ZN => n18331);
   U24208 : AOI21_X1 port map( A1 => n18840, A2 => n1181, B => n30937, ZN => 
                           n18347);
   U24209 : NAND2_X1 port map( A1 => n26181, A2 => n19052, ZN => n18346);
   U24211 : NAND3_X1 port map( A1 => n18339, A2 => n18779, A3 => n10080, ZN => 
                           n18341);
   U24214 : XOR2_X1 port map( A1 => Key(39), A2 => Plaintext(39), Z => n18649);
   U24215 : INV_X1 port map( I => Plaintext(37), ZN => n18348);
   U24216 : INV_X1 port map( I => Plaintext(30), ZN => n18350);
   U24220 : INV_X1 port map( I => Plaintext(8), ZN => n18354);
   U24222 : XOR2_X1 port map( A1 => Key(11), A2 => Plaintext(11), Z => n18674);
   U24223 : INV_X1 port map( I => Plaintext(18), ZN => n18356);
   U24224 : XOR2_X1 port map( A1 => Key(21), A2 => Plaintext(21), Z => n18357);
   U24226 : NAND2_X1 port map( A1 => n18793, A2 => n26810, ZN => n18361);
   U24227 : INV_X1 port map( I => Plaintext(48), ZN => n18364);
   U24228 : INV_X1 port map( I => Plaintext(49), ZN => n18365);
   U24230 : XOR2_X1 port map( A1 => Key(42), A2 => Plaintext(42), Z => n18811);
   U24231 : OAI21_X1 port map( A1 => n8422, A2 => n18779, B => n6215, ZN => 
                           n18368);
   U24232 : NAND2_X1 port map( A1 => n18368, A2 => n18618, ZN => n18372);
   U24235 : NOR2_X1 port map( A1 => n12074, A2 => n18642, ZN => n18375);
   U24236 : NAND2_X1 port map( A1 => n18378, A2 => n18377, ZN => n18379);
   U24237 : INV_X1 port map( I => Plaintext(118), ZN => n18382);
   U24238 : NOR2_X1 port map( A1 => n956, A2 => n18459, ZN => n18387);
   U24241 : XOR2_X1 port map( A1 => Key(113), A2 => Plaintext(113), Z => n18696
                           );
   U24242 : XOR2_X1 port map( A1 => Key(108), A2 => Plaintext(108), Z => n18831
                           );
   U24243 : XOR2_X1 port map( A1 => Key(109), A2 => Plaintext(109), Z => n18700
                           );
   U24245 : XOR2_X1 port map( A1 => Key(123), A2 => Plaintext(123), Z => n18429
                           );
   U24246 : INV_X1 port map( I => Plaintext(120), ZN => n18393);
   U24249 : INV_X1 port map( I => Plaintext(3), ZN => n18395);
   U24250 : XOR2_X1 port map( A1 => n18395, A2 => Key(3), Z => n18888);
   U24251 : XOR2_X1 port map( A1 => Key(1), A2 => Plaintext(1), Z => n18660);
   U24252 : INV_X1 port map( I => Plaintext(183), ZN => n18396);
   U24254 : XOR2_X1 port map( A1 => Key(181), A2 => Plaintext(181), Z => n18688
                           );
   U24255 : INV_X1 port map( I => Plaintext(184), ZN => n18398);
   U24256 : XOR2_X1 port map( A1 => Key(187), A2 => Plaintext(187), Z => n18844
                           );
   U24257 : INV_X2 port map( I => n18844, ZN => n18681);
   U24258 : XOR2_X1 port map( A1 => Key(173), A2 => Plaintext(173), Z => n18402
                           );
   U24259 : INV_X1 port map( I => Plaintext(172), ZN => n18401);
   U24261 : XOR2_X1 port map( A1 => Key(167), A2 => Plaintext(167), Z => n18861
                           );
   U24262 : XOR2_X1 port map( A1 => Key(162), A2 => Plaintext(162), Z => n18862
                           );
   U24263 : INV_X1 port map( I => Plaintext(163), ZN => n18404);
   U24265 : NAND2_X1 port map( A1 => n10182, A2 => n18101, ZN => n18406);
   U24267 : NAND2_X1 port map( A1 => n31821, A2 => n18726, ZN => n18408);
   U24274 : NAND3_X1 port map( A1 => n18720, A2 => n16614, A3 => n8411, ZN => 
                           n18416);
   U24275 : NAND2_X2 port map( A1 => n18417, A2 => n18416, ZN => n19318);
   U24276 : NAND2_X1 port map( A1 => n33432, A2 => n19318, ZN => n18418);
   U24277 : NAND3_X1 port map( A1 => n19321, A2 => n18419, A3 => n18418, ZN => 
                           n18420);
   U24278 : NOR2_X1 port map( A1 => n19158, A2 => n14811, ZN => n18425);
   U24280 : INV_X1 port map( I => n18831, ZN => n18427);
   U24281 : INV_X1 port map( I => n18434, ZN => n18746);
   U24282 : NAND2_X1 port map( A1 => n8208, A2 => n6359, ZN => n18437);
   U24284 : NOR2_X1 port map( A1 => n18446, A2 => n18797, ZN => n18444);
   U24287 : NAND2_X1 port map( A1 => n18454, A2 => n17725, ZN => n18456);
   U24288 : NOR2_X1 port map( A1 => n18456, A2 => n18455, ZN => n18458);
   U24289 : NOR2_X1 port map( A1 => n18995, A2 => n18976, ZN => n18468);
   U24292 : NOR2_X1 port map( A1 => n18994, A2 => n100, ZN => n18467);
   U24294 : NOR2_X1 port map( A1 => n18006, A2 => n18699, ZN => n18471);
   U24298 : NAND2_X1 port map( A1 => n16585, A2 => n18811, ZN => n18479);
   U24300 : NOR3_X1 port map( A1 => n18481, A2 => n17597, A3 => n14093, ZN => 
                           n18482);
   U24301 : NOR2_X1 port map( A1 => n16417, A2 => n10080, ZN => n18483);
   U24302 : NAND2_X1 port map( A1 => n18601, A2 => n18755, ZN => n18501);
   U24303 : NAND2_X1 port map( A1 => n18761, A2 => n18605, ZN => n18500);
   U24304 : AOI21_X1 port map( A1 => n18501, A2 => n18500, B => n27940, ZN => 
                           n18502);
   U24305 : OR2_X1 port map( A1 => n18899, A2 => n19088, Z => n18504);
   U24306 : NOR2_X1 port map( A1 => n17516, A2 => n15888, ZN => n18507);
   U24308 : NAND2_X1 port map( A1 => n16732, A2 => n33941, ZN => n18512);
   U24310 : NOR2_X1 port map( A1 => n18845, A2 => n18731, ZN => n18520);
   U24311 : OAI21_X1 port map( A1 => n957, A2 => n18520, B => n18519, ZN => 
                           n18524);
   U24312 : NOR2_X1 port map( A1 => n17184, A2 => n18847, ZN => n18521);
   U24316 : NAND2_X1 port map( A1 => n18704, A2 => n18743, ZN => n18536);
   U24320 : NAND2_X1 port map( A1 => n18349, A2 => n18548, ZN => n18550);
   U24321 : MUX2_X1 port map( I0 => n18550, I1 => n18549, S => n17114, Z => 
                           n18551);
   U24323 : AOI21_X1 port map( A1 => n18559, A2 => n18623, B => n27129, ZN => 
                           n18561);
   U24324 : NAND2_X1 port map( A1 => n18774, A2 => n18771, ZN => n18560);
   U24329 : NOR2_X1 port map( A1 => n18848, A2 => n17030, ZN => n18596);
   U24330 : NOR2_X1 port map( A1 => n18402, A2 => n18846, ZN => n18595);
   U24332 : INV_X1 port map( I => n19158, ZN => n18599);
   U24333 : OAI21_X1 port map( A1 => n18599, A2 => n14812, B => n12548, ZN => 
                           n18600);
   U24335 : NOR2_X1 port map( A1 => n18618, A2 => n1430, ZN => n18619);
   U24336 : NOR2_X1 port map( A1 => n13254, A2 => n17937, ZN => n18627);
   U24337 : INV_X1 port map( I => n18821, ZN => n18632);
   U24341 : NOR2_X1 port map( A1 => n18683, A2 => n5700, ZN => n18651);
   U24343 : AOI22_X1 port map( A1 => n18798, A2 => n31724, B1 => n18797, B2 => 
                           n18655, ZN => n18656);
   U24344 : NOR2_X1 port map( A1 => n18656, A2 => n16420, ZN => n18657);
   U24345 : AOI21_X1 port map( A1 => n31971, A2 => n28675, B => n18687, ZN => 
                           n18664);
   U24346 : NOR2_X1 port map( A1 => n18866, A2 => n18871, ZN => n18663);
   U24347 : NOR2_X1 port map( A1 => n18664, A2 => n18663, ZN => n18666);
   U24351 : NAND2_X1 port map( A1 => n18692, A2 => n711, ZN => n18693);
   U24354 : NAND2_X1 port map( A1 => n18853, A2 => n15211, ZN => n18719);
   U24355 : AOI21_X1 port map( A1 => n18720, A2 => n16614, B => n18307, ZN => 
                           n18721);
   U24358 : NOR2_X1 port map( A1 => n18736, A2 => n17687, ZN => n18741);
   U24359 : NOR2_X1 port map( A1 => n18747, A2 => n18742, ZN => n18744);
   U24360 : NAND2_X1 port map( A1 => n18747, A2 => n18746, ZN => n18748);
   U24362 : NAND2_X1 port map( A1 => n14093, A2 => n18755, ZN => n18757);
   U24364 : NAND2_X1 port map( A1 => n18762, A2 => n18761, ZN => n19095);
   U24365 : NOR2_X1 port map( A1 => n18775, A2 => n18770, ZN => n18772);
   U24367 : NAND2_X1 port map( A1 => n31095, A2 => n1430, ZN => n18781);
   U24369 : NAND2_X1 port map( A1 => n18798, A2 => n18797, ZN => n18799);
   U24371 : XOR2_X1 port map( A1 => n9665, A2 => n24869, Z => n18814);
   U24373 : NOR2_X1 port map( A1 => n785, A2 => n18515, ZN => n18819);
   U24374 : NAND2_X1 port map( A1 => n18819, A2 => n16393, ZN => n19041);
   U24375 : NOR2_X1 port map( A1 => n171, A2 => n4868, ZN => n18825);
   U24376 : NAND2_X1 port map( A1 => n18829, A2 => n18827, ZN => n18828);
   U24378 : INV_X1 port map( I => n18921, ZN => n18836);
   U24379 : NAND3_X1 port map( A1 => n32784, A2 => n18836, A3 => n31324, ZN => 
                           n18838);
   U24380 : NOR2_X1 port map( A1 => n18848, A2 => n18847, ZN => n18851);
   U24385 : XOR2_X1 port map( A1 => n29030, A2 => n16454, Z => n18898);
   U24387 : NAND2_X1 port map( A1 => n19315, A2 => n825, ZN => n18904);
   U24388 : XOR2_X1 port map( A1 => n32262, A2 => n25038, Z => n18915);
   U24390 : NOR2_X1 port map( A1 => n28935, A2 => n18923, ZN => n18925);
   U24392 : XOR2_X1 port map( A1 => n28806, A2 => n25910, Z => n18932);
   U24394 : NAND3_X1 port map( A1 => n30959, A2 => n18939, A3 => n31949, ZN => 
                           n18940);
   U24396 : XOR2_X1 port map( A1 => n30443, A2 => n25519, Z => n18948);
   U24402 : NOR2_X1 port map( A1 => n31850, A2 => n16288, ZN => n18984);
   U24403 : NOR2_X1 port map( A1 => n14498, A2 => n18990, ZN => n18989);
   U24407 : INV_X1 port map( I => n13925, ZN => n19017);
   U24411 : NAND3_X1 port map( A1 => n10124, A2 => n745, A3 => n19196, ZN => 
                           n19024);
   U24413 : NAND2_X1 port map( A1 => n14130, A2 => n19202, ZN => n19028);
   U24414 : NAND2_X1 port map( A1 => n19301, A2 => n26600, ZN => n19027);
   U24415 : NAND3_X1 port map( A1 => n19028, A2 => n730, A3 => n19027, ZN => 
                           n19031);
   U24416 : NOR2_X1 port map( A1 => n16354, A2 => n16093, ZN => n19029);
   U24417 : INV_X1 port map( I => n19040, ZN => n19045);
   U24418 : INV_X1 port map( I => n19041, ZN => n19044);
   U24419 : INV_X1 port map( I => n19042, ZN => n19043);
   U24420 : NOR3_X1 port map( A1 => n19045, A2 => n19044, A3 => n19043, ZN => 
                           n19047);
   U24422 : NOR3_X1 port map( A1 => n1053, A2 => n19109, A3 => n19063, ZN => 
                           n19064);
   U24424 : NOR2_X1 port map( A1 => n19318, A2 => n19275, ZN => n19068);
   U24425 : NOR2_X1 port map( A1 => n19317, A2 => n30894, ZN => n19067);
   U24426 : INV_X1 port map( I => n19356, ZN => n19069);
   U24427 : NAND2_X1 port map( A1 => n19069, A2 => n6516, ZN => n19071);
   U24428 : NAND2_X1 port map( A1 => n15842, A2 => n6516, ZN => n19070);
   U24429 : AOI22_X1 port map( A1 => n19071, A2 => n19281, B1 => n19070, B2 => 
                           n19354, ZN => n19072);
   U24432 : INV_X1 port map( I => n19094, ZN => n19098);
   U24433 : AOI22_X1 port map( A1 => n19126, A2 => n31850, B1 => n19125, B2 => 
                           n7968, ZN => n19131);
   U24434 : XOR2_X1 port map( A1 => n19651, A2 => n16727, Z => n19447);
   U24435 : NOR2_X1 port map( A1 => n7810, A2 => n1379, ZN => n19134);
   U24437 : OAI21_X1 port map( A1 => n19137, A2 => n744, B => n25971, ZN => 
                           n19141);
   U24438 : NOR2_X1 port map( A1 => n19257, A2 => n19258, ZN => n19139);
   U24439 : NOR2_X1 port map( A1 => n19255, A2 => n19143, ZN => n19144);
   U24440 : NAND2_X1 port map( A1 => n4747, A2 => n25961, ZN => n19150);
   U24442 : NAND2_X1 port map( A1 => n16007, A2 => n19160, ZN => n19161);
   U24445 : XOR2_X1 port map( A1 => n19474, A2 => n16561, Z => n19193);
   U24446 : XOR2_X1 port map( A1 => n19384, A2 => n25815, Z => n19211);
   U24448 : MUX2_X1 port map( I0 => n19275, I1 => n30894, S => n19318, Z => 
                           n19233);
   U24449 : NAND2_X1 port map( A1 => n11940, A2 => n26603, ZN => n19240);
   U24450 : NAND3_X1 port map( A1 => n19243, A2 => n19242, A3 => n877, ZN => 
                           n19246);
   U24455 : MUX2_X1 port map( I0 => n19318, I1 => n27132, S => n19275, Z => 
                           n19277);
   U24456 : NAND2_X1 port map( A1 => n19322, A2 => n19320, ZN => n19276);
   U24457 : OAI21_X2 port map( A1 => n19278, A2 => n19277, B => n19276, ZN => 
                           n19641);
   U24459 : INV_X1 port map( I => n19292, ZN => n19293);
   U24460 : OAI21_X1 port map( A1 => n746, A2 => n19295, B => n19294, ZN => 
                           n19296);
   U24462 : NOR2_X1 port map( A1 => n19302, A2 => n19301, ZN => n19303);
   U24466 : XOR2_X1 port map( A1 => n19412, A2 => n15117, Z => n19342);
   U24467 : XOR2_X1 port map( A1 => n19625, A2 => n25074, Z => n19344);
   U24468 : XOR2_X1 port map( A1 => n11218, A2 => n19344, Z => n19345);
   U24470 : INV_X1 port map( I => n19349, ZN => n19347);
   U24471 : NAND2_X1 port map( A1 => n19347, A2 => n19346, ZN => n19351);
   U24472 : NAND2_X1 port map( A1 => n19349, A2 => n27941, ZN => n19350);
   U24474 : NAND2_X1 port map( A1 => n19361, A2 => n16444, ZN => n19362);
   U24475 : NAND2_X1 port map( A1 => n19363, A2 => n19362, ZN => n19366);
   U24477 : XOR2_X1 port map( A1 => n30212, A2 => n25929, Z => n19372);
   U24478 : XOR2_X1 port map( A1 => n19373, A2 => n19372, Z => n19374);
   U24483 : XOR2_X1 port map( A1 => n19630, A2 => n16550, Z => n19390);
   U24484 : XOR2_X1 port map( A1 => n19755, A2 => n16619, Z => n19394);
   U24486 : XOR2_X1 port map( A1 => n15028, A2 => n25720, Z => n19397);
   U24487 : XOR2_X1 port map( A1 => n19644, A2 => n24231, Z => n19401);
   U24488 : XOR2_X1 port map( A1 => n19405, A2 => n19549, Z => n19407);
   U24489 : XOR2_X1 port map( A1 => n19409, A2 => n19754, Z => n19411);
   U24491 : XOR2_X1 port map( A1 => n19412, A2 => n19589, Z => n19507);
   U24492 : XOR2_X1 port map( A1 => n29890, A2 => n16423, Z => n19413);
   U24493 : XOR2_X1 port map( A1 => n19414, A2 => n19415, Z => n19419);
   U24494 : NAND3_X1 port map( A1 => n29156, A2 => n19799, A3 => n19886, ZN => 
                           n19422);
   U24495 : XOR2_X1 port map( A1 => n19416, A2 => n25358, Z => n19417);
   U24497 : XOR2_X1 port map( A1 => n19684, A2 => n19427, Z => n19428);
   U24498 : XOR2_X1 port map( A1 => n19429, A2 => n19428, Z => n19796);
   U24500 : XOR2_X1 port map( A1 => n19711, A2 => n19434, Z => n19435);
   U24504 : NAND3_X1 port map( A1 => n25997, A2 => n12038, A3 => n11913, ZN => 
                           n19460);
   U24505 : XOR2_X1 port map( A1 => n19649, A2 => n25722, Z => n19465);
   U24506 : XOR2_X1 port map( A1 => n16138, A2 => n16604, Z => n19471);
   U24508 : XOR2_X1 port map( A1 => n15787, A2 => n25079, Z => n19487);
   U24509 : XOR2_X1 port map( A1 => n19509, A2 => n16390, Z => n19496);
   U24510 : XOR2_X1 port map( A1 => n19498, A2 => n19524, Z => n19500);
   U24511 : XOR2_X1 port map( A1 => n28399, A2 => n16653, Z => n19501);
   U24512 : INV_X1 port map( I => Key(2), ZN => n24831);
   U24514 : XOR2_X1 port map( A1 => n19508, A2 => n34077, Z => n19511);
   U24515 : XOR2_X1 port map( A1 => n19509, A2 => n24895, Z => n19510);
   U24516 : XOR2_X1 port map( A1 => n19511, A2 => n19510, Z => n19512);
   U24517 : XOR2_X1 port map( A1 => n19755, A2 => n24833, Z => n19516);
   U24519 : XOR2_X1 port map( A1 => n19764, A2 => n19524, Z => n19525);
   U24520 : XOR2_X1 port map( A1 => n19699, A2 => n19525, Z => n19526);
   U24521 : INV_X1 port map( I => n19530, ZN => n19531);
   U24522 : INV_X1 port map( I => n19833, ZN => n20040);
   U24523 : OAI21_X1 port map( A1 => n20040, A2 => n1169, B => n19834, ZN => 
                           n19534);
   U24524 : XOR2_X1 port map( A1 => n19736, A2 => n19539, Z => n19540);
   U24527 : XOR2_X1 port map( A1 => n19754, A2 => n16634, Z => n19559);
   U24528 : XOR2_X1 port map( A1 => n30766, A2 => n25554, Z => n19573);
   U24529 : XOR2_X1 port map( A1 => n19589, A2 => n24738, Z => n19590);
   U24530 : XOR2_X1 port map( A1 => n19591, A2 => n19590, Z => n19596);
   U24531 : XOR2_X1 port map( A1 => n15844, A2 => n19592, Z => n19593);
   U24532 : XOR2_X1 port map( A1 => n19594, A2 => n19593, Z => n19595);
   U24534 : XOR2_X1 port map( A1 => n19676, A2 => n25641, Z => n19602);
   U24535 : INV_X1 port map( I => n19603, ZN => n19607);
   U24536 : AOI22_X1 port map( A1 => n19607, A2 => n19606, B1 => n19605, B2 => 
                           n19604, ZN => n19609);
   U24537 : XOR2_X1 port map( A1 => n29718, A2 => n19609, Z => n19610);
   U24538 : XOR2_X1 port map( A1 => n19611, A2 => n19610, Z => n19612);
   U24539 : XOR2_X1 port map( A1 => n19612, A2 => n19613, Z => n19829);
   U24540 : XOR2_X1 port map( A1 => n12048, A2 => n16530, Z => n19615);
   U24543 : XOR2_X1 port map( A1 => n30411, A2 => n19649, Z => n19653);
   U24545 : XOR2_X1 port map( A1 => n32697, A2 => n25436, Z => n19655);
   U24549 : XOR2_X1 port map( A1 => n19661, A2 => n24417, Z => n19663);
   U24554 : NAND2_X1 port map( A1 => n18199, A2 => n19899, ZN => n20107);
   U24556 : XOR2_X1 port map( A1 => n19682, A2 => n25091, Z => n19683);
   U24557 : XOR2_X1 port map( A1 => n19684, A2 => n19683, Z => n19685);
   U24558 : XOR2_X1 port map( A1 => n32271, A2 => n19691, Z => n19694);
   U24560 : XOR2_X1 port map( A1 => n19696, A2 => n25610, Z => n19697);
   U24562 : XOR2_X1 port map( A1 => n19712, A2 => n16662, Z => n19713);
   U24563 : INV_X1 port map( I => Key(27), ZN => n19718);
   U24569 : XOR2_X1 port map( A1 => n19751, A2 => n19750, Z => n19752);
   U24570 : OAI21_X1 port map( A1 => n31683, A2 => n26368, B => n20112, ZN => 
                           n19761);
   U24573 : XOR2_X1 port map( A1 => n19771, A2 => n19770, Z => n19777);
   U24574 : XOR2_X1 port map( A1 => n19773, A2 => n25751, Z => n19774);
   U24575 : XOR2_X1 port map( A1 => n19775, A2 => n19774, Z => n19776);
   U24576 : XOR2_X1 port map( A1 => n19777, A2 => n19776, Z => n20083);
   U24577 : XOR2_X1 port map( A1 => n8571, A2 => n25040, Z => n19786);
   U24578 : AOI21_X1 port map( A1 => n19789, A2 => n20085, B => n16664, ZN => 
                           n19790);
   U24580 : NAND3_X1 port map( A1 => n20034, A2 => n20032, A3 => n19971, ZN => 
                           n19810);
   U24582 : INV_X1 port map( I => n20083, ZN => n20007);
   U24585 : NOR2_X1 port map( A1 => n15394, A2 => n17299, ZN => n19831);
   U24594 : NAND2_X1 port map( A1 => n27600, A2 => n11453, ZN => n19865);
   U24597 : AOI21_X2 port map( A1 => n19872, A2 => n821, B => n19871, ZN => 
                           n20521);
   U24598 : NAND2_X1 port map( A1 => n29339, A2 => n16491, ZN => n19875);
   U24599 : INV_X1 port map( I => n19933, ZN => n19876);
   U24601 : NAND3_X1 port map( A1 => n2606, A2 => n20096, A3 => n3915, ZN => 
                           n20293);
   U24605 : MUX2_X1 port map( I0 => n19896, I1 => n12682, S => n20136, Z => 
                           n20229);
   U24606 : NAND2_X1 port map( A1 => n16595, A2 => n20021, ZN => n19897);
   U24609 : NOR3_X1 port map( A1 => n19912, A2 => n19913, A3 => n12142, ZN => 
                           n19911);
   U24611 : INV_X1 port map( I => n8259, ZN => n19917);
   U24617 : NOR2_X1 port map( A1 => n4254, A2 => n20486, ZN => n19957);
   U24619 : INV_X1 port map( I => n20631, ZN => n19972);
   U24620 : NAND2_X1 port map( A1 => n19965, A2 => n20018, ZN => n19968);
   U24621 : AOI21_X1 port map( A1 => n20033, A2 => n2795, B => n16243, ZN => 
                           n19970);
   U24623 : NAND2_X1 port map( A1 => n19819, A2 => n32745, ZN => n19975);
   U24629 : XOR2_X1 port map( A1 => n20693, A2 => n16602, Z => n20005);
   U24630 : XOR2_X1 port map( A1 => n20722, A2 => n20005, Z => n20050);
   U24631 : OAI21_X1 port map( A1 => n20020, A2 => n20019, B => n20119, ZN => 
                           n20024);
   U24638 : INV_X1 port map( I => n20060, ZN => n20063);
   U24640 : INV_X1 port map( I => n20070, ZN => n20073);
   U24644 : MUX2_X1 port map( I0 => n20122, I1 => n20121, S => n14334, Z => 
                           n20127);
   U24645 : NOR2_X2 port map( A1 => n20127, A2 => n20126, ZN => n20460);
   U24650 : NAND2_X1 port map( A1 => n20266, A2 => n28376, ZN => n20163);
   U24651 : XOR2_X1 port map( A1 => n20868, A2 => n20166, Z => n20167);
   U24652 : XOR2_X1 port map( A1 => n20168, A2 => n20167, Z => n21258);
   U24653 : MUX2_X1 port map( I0 => n13768, I1 => n16374, S => n20556, Z => 
                           n20169);
   U24656 : NAND2_X1 port map( A1 => n28414, A2 => n20499, ZN => n20175);
   U24659 : INV_X1 port map( I => n20188, ZN => n20193);
   U24660 : INV_X1 port map( I => n20190, ZN => n20192);
   U24663 : INV_X1 port map( I => n20209, ZN => n20210);
   U24666 : NAND2_X1 port map( A1 => n4254, A2 => n20221, ZN => n20222);
   U24667 : XOR2_X1 port map( A1 => n20729, A2 => n20784, Z => n20226);
   U24668 : XOR2_X1 port map( A1 => n20715, A2 => n16548, Z => n20225);
   U24669 : NAND3_X1 port map( A1 => n20520, A2 => n16218, A3 => n20556, ZN => 
                           n20237);
   U24670 : XOR2_X1 port map( A1 => n20733, A2 => n25252, Z => n20241);
   U24672 : INV_X1 port map( I => n16050, ZN => n20255);
   U24673 : NAND2_X1 port map( A1 => n16951, A2 => n11182, ZN => n20256);
   U24675 : AOI22_X1 port map( A1 => n20651, A2 => n20271, B1 => n28575, B2 => 
                           n20270, ZN => n20272);
   U24676 : MUX2_X1 port map( I0 => n20273, I1 => n1157, S => n15434, Z => 
                           n20275);
   U24679 : INV_X1 port map( I => n20280, ZN => n20281);
   U24681 : INV_X1 port map( I => n16515, ZN => n20284);
   U24682 : NAND4_X1 port map( A1 => n20294, A2 => n20291, A3 => n20292, A4 => 
                           n20293, ZN => n20296);
   U24685 : NAND2_X1 port map( A1 => n12872, A2 => n6230, ZN => n20314);
   U24686 : XOR2_X1 port map( A1 => n3009, A2 => n16619, Z => n20318);
   U24687 : NAND3_X1 port map( A1 => n818, A2 => n710, A3 => n20335, ZN => 
                           n20336);
   U24690 : XOR2_X1 port map( A1 => n33969, A2 => n25358, Z => n20356);
   U24691 : XOR2_X1 port map( A1 => n21038, A2 => n20356, Z => n20357);
   U24695 : INV_X1 port map( I => n25428, ZN => n20389);
   U24703 : AOI21_X1 port map( A1 => n20562, A2 => n30931, B => n20523, ZN => 
                           n20415);
   U24706 : OAI21_X2 port map( A1 => n20422, A2 => n20421, B => n20420, ZN => 
                           n21043);
   U24707 : NAND2_X1 port map( A1 => n17329, A2 => n4647, ZN => n20424);
   U24708 : INV_X1 port map( I => n20431, ZN => n20432);
   U24709 : INV_X1 port map( I => n20433, ZN => n20434);
   U24710 : INV_X1 port map( I => n20495, ZN => n20440);
   U24712 : NAND2_X1 port map( A1 => n4468, A2 => n31768, ZN => n20446);
   U24714 : INV_X1 port map( I => n20453, ZN => n20456);
   U24716 : NAND3_X1 port map( A1 => n29695, A2 => n20489, A3 => n28812, ZN => 
                           n20490);
   U24717 : NOR2_X1 port map( A1 => n20495, A2 => n20494, ZN => n20496);
   U24719 : XOR2_X1 port map( A1 => n20920, A2 => n7705, Z => n20513);
   U24720 : XOR2_X1 port map( A1 => n20824, A2 => n16581, Z => n20512);
   U24721 : XOR2_X1 port map( A1 => n20512, A2 => n20513, Z => n20514);
   U24724 : XOR2_X1 port map( A1 => n21046, A2 => n16497, Z => n20542);
   U24725 : XOR2_X1 port map( A1 => n20586, A2 => n2616, Z => n20588);
   U24732 : NAND4_X1 port map( A1 => n20625, A2 => n20624, A3 => n20623, A4 => 
                           n20622, ZN => n20626);
   U24735 : XOR2_X1 port map( A1 => n32162, A2 => n25126, Z => n20640);
   U24736 : XOR2_X1 port map( A1 => n20690, A2 => n16504, Z => n20642);
   U24737 : XOR2_X1 port map( A1 => n32791, A2 => n24861, Z => n20645);
   U24738 : XOR2_X1 port map( A1 => n20984, A2 => n20647, Z => n20649);
   U24741 : XOR2_X1 port map( A1 => n20658, A2 => n24417, Z => n20659);
   U24742 : XOR2_X1 port map( A1 => n20660, A2 => n20659, Z => n20661);
   U24743 : XOR2_X1 port map( A1 => n20857, A2 => n25783, Z => n20663);
   U24746 : XOR2_X1 port map( A1 => n20747, A2 => n8487, Z => n20667);
   U24748 : XOR2_X1 port map( A1 => n5348, A2 => n25191, Z => n20672);
   U24749 : XOR2_X1 port map( A1 => n20673, A2 => n20672, Z => n20675);
   U24751 : XOR2_X1 port map( A1 => n21016, A2 => n16697, Z => n20682);
   U24753 : XOR2_X1 port map( A1 => n20775, A2 => n25054, Z => n20694);
   U24754 : XOR2_X1 port map( A1 => n20695, A2 => n20694, Z => n20696);
   U24755 : XOR2_X1 port map( A1 => n25619, A2 => n20720, Z => n20697);
   U24757 : XOR2_X1 port map( A1 => n20743, A2 => n20702, Z => n20704);
   U24758 : XOR2_X1 port map( A1 => n20848, A2 => n24623, Z => n20703);
   U24759 : XOR2_X1 port map( A1 => n20837, A2 => n16604, Z => n20706);
   U24761 : XOR2_X1 port map( A1 => n10522, A2 => n20756, Z => n20707);
   U24762 : XOR2_X1 port map( A1 => n20851, A2 => n16578, Z => n20719);
   U24763 : XOR2_X1 port map( A1 => n20917, A2 => n20836, Z => n20724);
   U24764 : XOR2_X1 port map( A1 => n21029, A2 => n16671, Z => n20731);
   U24766 : XOR2_X1 port map( A1 => n21019, A2 => n25182, Z => n20737);
   U24768 : INV_X1 port map( I => n23239, ZN => n25213);
   U24769 : XOR2_X1 port map( A1 => n32749, A2 => n16680, Z => n20744);
   U24770 : XOR2_X1 port map( A1 => n14132, A2 => n25728, Z => n20749);
   U24772 : XOR2_X1 port map( A1 => n21001, A2 => n24514, Z => n20759);
   U24775 : XOR2_X1 port map( A1 => n1342, A2 => n16555, Z => n20770);
   U24776 : XOR2_X1 port map( A1 => n20771, A2 => n20770, Z => n20774);
   U24778 : INV_X1 port map( I => n21402, ZN => n20795);
   U24779 : XOR2_X1 port map( A1 => n29241, A2 => n18019, Z => n20793);
   U24784 : XOR2_X1 port map( A1 => n30219, A2 => n25288, Z => n20815);
   U24789 : XOR2_X1 port map( A1 => n28864, A2 => n20839, Z => n20840);
   U24790 : XOR2_X1 port map( A1 => n20841, A2 => n20840, Z => n20846);
   U24791 : XOR2_X1 port map( A1 => n20843, A2 => n24907, Z => n20844);
   U24792 : XOR2_X1 port map( A1 => n20919, A2 => n20844, Z => n20845);
   U24793 : XOR2_X1 port map( A1 => n20845, A2 => n20846, Z => n21389);
   U24795 : XOR2_X1 port map( A1 => n21024, A2 => n20183, Z => n20865);
   U24796 : XOR2_X1 port map( A1 => n20865, A2 => n20864, Z => n20866);
   U24797 : NAND2_X1 port map( A1 => n20880, A2 => n6408, ZN => n20875);
   U24800 : XOR2_X1 port map( A1 => n1023, A2 => n25040, Z => n20908);
   U24802 : NOR2_X1 port map( A1 => n20909, A2 => n31760, ZN => n20910);
   U24803 : XOR2_X1 port map( A1 => n32478, A2 => n24992, Z => n20922);
   U24804 : XOR2_X1 port map( A1 => n20926, A2 => n16575, Z => n20927);
   U24805 : AOI21_X1 port map( A1 => n21363, A2 => n20932, B => n21182, ZN => 
                           n20934);
   U24806 : NAND2_X1 port map( A1 => n21363, A2 => n27382, ZN => n20933);
   U24808 : NOR2_X1 port map( A1 => n27773, A2 => n20945, ZN => n20944);
   U24812 : XOR2_X1 port map( A1 => n20975, A2 => n25641, Z => n20976);
   U24813 : XOR2_X1 port map( A1 => n20985, A2 => n25064, Z => n20986);
   U24814 : XOR2_X1 port map( A1 => n28687, A2 => n24999, Z => n20995);
   U24815 : XOR2_X1 port map( A1 => n20996, A2 => n20997, Z => n20998);
   U24817 : XOR2_X1 port map( A1 => n21001, A2 => n24374, Z => n21002);
   U24818 : XOR2_X1 port map( A1 => n21003, A2 => n21002, Z => n21004);
   U24819 : XOR2_X1 port map( A1 => n21005, A2 => n21004, Z => n21068);
   U24820 : INV_X1 port map( I => n21068, ZN => n21424);
   U24821 : XOR2_X1 port map( A1 => n21029, A2 => n25506, Z => n21030);
   U24822 : XOR2_X1 port map( A1 => n21031, A2 => n21030, Z => n21032);
   U24825 : NOR2_X1 port map( A1 => n16034, A2 => n8490, ZN => n21066);
   U24827 : NOR2_X1 port map( A1 => n5480, A2 => n21075, ZN => n21076);
   U24828 : NAND2_X1 port map( A1 => n21160, A2 => n4145, ZN => n21088);
   U24829 : MUX2_X1 port map( I0 => n21088, I1 => n32452, S => n26777, Z => 
                           n21090);
   U24831 : NAND2_X1 port map( A1 => n21206, A2 => n15874, ZN => n21098);
   U24832 : NAND3_X1 port map( A1 => n21289, A2 => n21143, A3 => n21396, ZN => 
                           n21097);
   U24833 : INV_X1 port map( I => n21100, ZN => n21303);
   U24837 : NAND2_X1 port map( A1 => n925, A2 => n6451, ZN => n21110);
   U24838 : INV_X1 port map( I => n24514, ZN => n25849);
   U24839 : XOR2_X1 port map( A1 => n8291, A2 => n25849, Z => n21112);
   U24841 : NAND2_X1 port map( A1 => n11187, A2 => n4381, ZN => n21118);
   U24842 : NAND2_X1 port map( A1 => n21306, A2 => n21307, ZN => n21129);
   U24845 : NAND3_X1 port map( A1 => n16034, A2 => n28642, A3 => n31965, ZN => 
                           n21137);
   U24846 : NAND2_X1 port map( A1 => n16222, A2 => n21592, ZN => n21594);
   U24849 : NOR2_X1 port map( A1 => n28190, A2 => n21379, ZN => n21159);
   U24854 : NAND2_X1 port map( A1 => n21439, A2 => n17832, ZN => n21226);
   U24857 : NOR2_X1 port map( A1 => n9186, A2 => n21237, ZN => n21634);
   U24861 : XOR2_X1 port map( A1 => n22147, A2 => n16680, Z => n21280);
   U24862 : NAND2_X1 port map( A1 => n1312, A2 => n1136, ZN => n21282);
   U24866 : MUX2_X1 port map( I0 => n21305, I1 => n21304, S => n21306, Z => 
                           n21310);
   U24875 : NAND2_X1 port map( A1 => n1328, A2 => n17416, ZN => n21346);
   U24877 : NAND3_X1 port map( A1 => n21340, A2 => n26542, A3 => n21339, ZN => 
                           n21345);
   U24880 : NOR2_X1 port map( A1 => n21369, A2 => n11966, ZN => n21370);
   U24883 : NOR3_X1 port map( A1 => n27711, A2 => n922, A3 => n6408, ZN => 
                           n21385);
   U24884 : NAND2_X1 port map( A1 => n21392, A2 => n21391, ZN => n21393);
   U24885 : NAND2_X1 port map( A1 => n8587, A2 => n812, ZN => n21394);
   U24890 : MUX2_X1 port map( I0 => n21469, I1 => n21467, S => n21793, Z => 
                           n21472);
   U24892 : NAND3_X1 port map( A1 => n21470, A2 => n21469, A3 => n8079, ZN => 
                           n21471);
   U24893 : NAND2_X1 port map( A1 => n21933, A2 => n21932, ZN => n21477);
   U24895 : NOR2_X1 port map( A1 => n21934, A2 => n28895, ZN => n21475);
   U24899 : MUX2_X1 port map( I0 => n21613, I1 => n21482, S => n21755, Z => 
                           n21485);
   U24900 : INV_X1 port map( I => n31765, ZN => n21487);
   U24902 : INV_X1 port map( I => n21497, ZN => n21502);
   U24903 : INV_X1 port map( I => n21498, ZN => n21501);
   U24904 : INV_X1 port map( I => n21499, ZN => n21500);
   U24905 : NOR3_X1 port map( A1 => n21502, A2 => n21501, A3 => n21500, ZN => 
                           n21503);
   U24912 : NOR2_X1 port map( A1 => n30677, A2 => n21532, ZN => n21534);
   U24914 : NAND2_X1 port map( A1 => n21539, A2 => n21857, ZN => n21540);
   U24917 : XOR2_X1 port map( A1 => n30495, A2 => n16705, Z => n21582);
   U24918 : OAI21_X1 port map( A1 => n31978, A2 => n21628, B => n2217, ZN => 
                           n21608);
   U24919 : INV_X1 port map( I => n21614, ZN => n21615);
   U24920 : NOR2_X1 port map( A1 => n21616, A2 => n21615, ZN => n21621);
   U24921 : INV_X1 port map( I => n21617, ZN => n21618);
   U24922 : NOR2_X1 port map( A1 => n21619, A2 => n21618, ZN => n21620);
   U24924 : INV_X1 port map( I => n21633, ZN => n21635);
   U24925 : NOR2_X1 port map( A1 => n21635, A2 => n21634, ZN => n21639);
   U24926 : NAND4_X1 port map( A1 => n31511, A2 => n21639, A3 => n21637, A4 => 
                           n21638, ZN => n21640);
   U24927 : NAND2_X1 port map( A1 => n30506, A2 => n15864, ZN => n21648);
   U24928 : XOR2_X1 port map( A1 => n3550, A2 => n25282, Z => n21650);
   U24929 : XOR2_X1 port map( A1 => n8291, A2 => n24992, Z => n21658);
   U24930 : NAND3_X1 port map( A1 => n21850, A2 => n21763, A3 => n15022, ZN => 
                           n21684);
   U24932 : OAI21_X1 port map( A1 => n26474, A2 => n21730, B => n920, ZN => 
                           n21731);
   U24936 : NAND2_X1 port map( A1 => n27649, A2 => n21755, ZN => n21753);
   U24938 : NAND2_X1 port map( A1 => n12587, A2 => n21763, ZN => n21760);
   U24939 : XOR2_X1 port map( A1 => n22086, A2 => n16550, Z => n21768);
   U24942 : NAND2_X1 port map( A1 => n21811, A2 => n21808, ZN => n21809);
   U24943 : XOR2_X1 port map( A1 => n21916, A2 => n21813, Z => n21814);
   U24944 : XOR2_X1 port map( A1 => n21815, A2 => n21814, Z => n22677);
   U24945 : INV_X1 port map( I => n21824, ZN => n21825);
   U24946 : INV_X1 port map( I => n21826, ZN => n21828);
   U24947 : INV_X1 port map( I => n21831, ZN => n21836);
   U24948 : NOR2_X1 port map( A1 => n11890, A2 => n25815, ZN => n21833);
   U24949 : OAI21_X1 port map( A1 => n1009, A2 => n15242, B => n21833, ZN => 
                           n21834);
   U24950 : OAI22_X1 port map( A1 => n21836, A2 => n25815, B1 => n21835, B2 => 
                           n21834, ZN => n21837);
   U24951 : AOI21_X1 port map( A1 => n25815, A2 => n34016, B => n21837, ZN => 
                           n21838);
   U24952 : INV_X1 port map( I => n21857, ZN => n21861);
   U24955 : XOR2_X1 port map( A1 => n21875, A2 => n21874, Z => n21881);
   U24956 : XOR2_X1 port map( A1 => n21878, A2 => n21879, Z => n21880);
   U24959 : XOR2_X1 port map( A1 => n22188, A2 => n25827, Z => n21884);
   U24960 : INV_X1 port map( I => n24417, ZN => n24435);
   U24961 : XOR2_X1 port map( A1 => n30306, A2 => n24435, Z => n21887);
   U24962 : XOR2_X1 port map( A1 => n16355, A2 => n22197, Z => n21888);
   U24963 : XOR2_X1 port map( A1 => n21923, A2 => n16687, Z => n21893);
   U24964 : INV_X1 port map( I => n12785, ZN => n21894);
   U24969 : XOR2_X1 port map( A1 => n21906, A2 => n21905, Z => n21907);
   U24970 : XOR2_X1 port map( A1 => n22044, A2 => n24748, Z => n21915);
   U24975 : XOR2_X1 port map( A1 => n22111, A2 => n22018, Z => n21939);
   U24976 : XOR2_X1 port map( A1 => n21940, A2 => n21939, Z => n21941);
   U24978 : XOR2_X1 port map( A1 => n21948, A2 => n21947, Z => n21950);
   U24979 : XOR2_X1 port map( A1 => n27180, A2 => n25104, Z => n21953);
   U24980 : NAND2_X1 port map( A1 => n22641, A2 => n33594, ZN => n21957);
   U24981 : XOR2_X1 port map( A1 => n21959, A2 => n22123, Z => n21960);
   U24982 : XOR2_X1 port map( A1 => n22226, A2 => n18019, Z => n21962);
   U24983 : XOR2_X1 port map( A1 => n22295, A2 => n16555, Z => n21967);
   U24985 : NAND2_X1 port map( A1 => n28124, A2 => n22489, ZN => n21972);
   U24990 : NAND2_X1 port map( A1 => n21979, A2 => n16240, ZN => n21980);
   U24991 : NAND3_X1 port map( A1 => n33007, A2 => n33115, A3 => n17930, ZN => 
                           n21983);
   U24993 : XOR2_X1 port map( A1 => n30495, A2 => n25735, Z => n21988);
   U24994 : XOR2_X1 port map( A1 => n22291, A2 => n25465, Z => n21999);
   U24997 : XOR2_X1 port map( A1 => n22239, A2 => n16507, Z => n22006);
   U25002 : XOR2_X1 port map( A1 => n22145, A2 => n25856, Z => n22022);
   U25005 : XOR2_X1 port map( A1 => n22251, A2 => n16581, Z => n22038);
   U25006 : XOR2_X1 port map( A1 => n22039, A2 => n22038, Z => n22040);
   U25007 : XOR2_X1 port map( A1 => n26957, A2 => n16402, Z => n22045);
   U25009 : NAND2_X1 port map( A1 => n22741, A2 => n22780, ZN => n22053);
   U25010 : XOR2_X1 port map( A1 => n7477, A2 => n25519, Z => n22057);
   U25011 : INV_X1 port map( I => n22185, ZN => n22058);
   U25012 : XOR2_X1 port map( A1 => n32885, A2 => n22058, Z => n22060);
   U25013 : XOR2_X1 port map( A1 => n28848, A2 => n25074, Z => n22062);
   U25019 : XOR2_X1 port map( A1 => n29011, A2 => n25500, Z => n22083);
   U25020 : XOR2_X1 port map( A1 => n32404, A2 => n22086, Z => n22088);
   U25021 : XOR2_X1 port map( A1 => n17555, A2 => n25373, Z => n22087);
   U25022 : XOR2_X1 port map( A1 => n22088, A2 => n22087, Z => n22089);
   U25023 : XOR2_X1 port map( A1 => n22090, A2 => n22089, Z => n22662);
   U25024 : XOR2_X1 port map( A1 => n22201, A2 => n25911, Z => n22093);
   U25025 : XOR2_X1 port map( A1 => n22093, A2 => n22259, Z => n22094);
   U25026 : XOR2_X1 port map( A1 => n16649, A2 => n27850, Z => n22103);
   U25027 : XOR2_X1 port map( A1 => n22104, A2 => n22103, Z => n22107);
   U25031 : XOR2_X1 port map( A1 => n22295, A2 => n16654, Z => n22133);
   U25034 : XOR2_X1 port map( A1 => n3550, A2 => n16666, Z => n22146);
   U25035 : INV_X1 port map( I => n22579, ZN => n22452);
   U25036 : XOR2_X1 port map( A1 => n28848, A2 => n24966, Z => n22151);
   U25037 : XOR2_X1 port map( A1 => n22162, A2 => n25049, Z => n22163);
   U25038 : XOR2_X1 port map( A1 => n17555, A2 => n16674, Z => n22174);
   U25039 : XOR2_X1 port map( A1 => n22175, A2 => n22174, Z => n22176);
   U25042 : XOR2_X1 port map( A1 => n22318, A2 => n25071, Z => n22181);
   U25049 : XOR2_X1 port map( A1 => n22238, A2 => n16502, Z => n22241);
   U25051 : MUX2_X1 port map( I0 => n22254, I1 => n22253, S => n28424, Z => 
                           n22258);
   U25052 : XOR2_X1 port map( A1 => n22260, A2 => n25783, Z => n22261);
   U25054 : NOR2_X1 port map( A1 => n28924, A2 => n32078, ZN => n22297);
   U25055 : XOR2_X1 port map( A1 => n22308, A2 => n25881, Z => n22309);
   U25056 : XOR2_X1 port map( A1 => n32154, A2 => n16655, Z => n22319);
   U25060 : NOR2_X1 port map( A1 => n22745, A2 => n27166, ZN => n22328);
   U25068 : NAND2_X1 port map( A1 => n11930, A2 => n22599, ZN => n22356);
   U25074 : XOR2_X1 port map( A1 => n23367, A2 => n25091, Z => n22384);
   U25075 : XOR2_X1 port map( A1 => n22385, A2 => n22384, Z => n22386);
   U25076 : XOR2_X1 port map( A1 => n22387, A2 => n22386, Z => n22617);
   U25079 : AOI21_X1 port map( A1 => n22408, A2 => n22534, B => n909, ZN => 
                           n22409);
   U25081 : NAND2_X1 port map( A1 => n22644, A2 => n33594, ZN => n22422);
   U25084 : NAND3_X1 port map( A1 => n22604, A2 => n17960, A3 => n14728, ZN => 
                           n22426);
   U25085 : NAND2_X1 port map( A1 => n16503, A2 => n22923, ZN => n22458);
   U25086 : NAND2_X1 port map( A1 => n22460, A2 => n5379, ZN => n22461);
   U25090 : NOR2_X1 port map( A1 => n22681, A2 => n11926, ZN => n22471);
   U25092 : NAND2_X1 port map( A1 => n22546, A2 => n1282, ZN => n22480);
   U25094 : OAI21_X1 port map( A1 => n14493, A2 => n22689, B => n15746, ZN => 
                           n22498);
   U25100 : XOR2_X1 port map( A1 => n9153, A2 => n25079, Z => n22515);
   U25101 : XOR2_X1 port map( A1 => n22516, A2 => n22515, Z => n22517);
   U25105 : NAND2_X1 port map( A1 => n22562, A2 => n16447, ZN => n22561);
   U25109 : NAND2_X1 port map( A1 => n22659, A2 => n22658, ZN => n22575);
   U25110 : INV_X1 port map( I => n22806, ZN => n22581);
   U25111 : NOR3_X1 port map( A1 => n22724, A2 => n22581, A3 => n22723, ZN => 
                           n22582);
   U25114 : XOR2_X1 port map( A1 => n23393, A2 => n16551, Z => n22616);
   U25119 : OAI21_X1 port map( A1 => n14183, A2 => n23072, B => n28970, ZN => 
                           n22692);
   U25121 : INV_X1 port map( I => n22697, ZN => n22698);
   U25122 : OAI21_X1 port map( A1 => n7181, A2 => n7881, B => n22827, ZN => 
                           n22706);
   U25123 : XOR2_X1 port map( A1 => n23328, A2 => n23363, Z => n22711);
   U25124 : MUX2_X1 port map( I0 => n30365, I1 => n26667, S => n23100, Z => 
                           n22710);
   U25125 : XOR2_X1 port map( A1 => n22711, A2 => n8298, Z => n22712);
   U25126 : XOR2_X1 port map( A1 => n23230, A2 => n25428, Z => n22719);
   U25127 : XOR2_X1 port map( A1 => n23373, A2 => n22719, Z => n22728);
   U25128 : NAND2_X1 port map( A1 => n6012, A2 => n23109, ZN => n22726);
   U25134 : MUX2_X1 port map( I0 => n22740, I1 => n22739, S => n3184, Z => 
                           n22743);
   U25136 : MUX2_X1 port map( I0 => n23583, I1 => n23745, S => n23770, Z => 
                           n22765);
   U25138 : NAND3_X1 port map( A1 => n22757, A2 => n23042, A3 => n13474, ZN => 
                           n22758);
   U25143 : XOR2_X1 port map( A1 => n23274, A2 => n25038, Z => n22799);
   U25149 : XOR2_X1 port map( A1 => n23467, A2 => n25064, Z => n22841);
   U25152 : INV_X1 port map( I => n3183, ZN => n22888);
   U25153 : OAI21_X1 port map( A1 => n29175, A2 => n3183, B => n22849, ZN => 
                           n22851);
   U25157 : XOR2_X1 port map( A1 => n23258, A2 => n25610, Z => n22867);
   U25158 : XOR2_X1 port map( A1 => n23439, A2 => n23189, Z => n22875);
   U25159 : XOR2_X1 port map( A1 => n23331, A2 => n22875, Z => n22877);
   U25161 : XOR2_X1 port map( A1 => n23274, A2 => n16472, Z => n22896);
   U25165 : NAND2_X1 port map( A1 => n22921, A2 => n22920, ZN => n22929);
   U25166 : INV_X1 port map( I => n22922, ZN => n22928);
   U25167 : INV_X1 port map( I => n22923, ZN => n22925);
   U25168 : OAI21_X1 port map( A1 => n31267, A2 => n22925, B => n22924, ZN => 
                           n22927);
   U25169 : NOR3_X1 port map( A1 => n22929, A2 => n22928, A3 => n22927, ZN => 
                           n22931);
   U25171 : XOR2_X1 port map( A1 => n23511, A2 => n23125, Z => n22934);
   U25172 : XOR2_X1 port map( A1 => n22935, A2 => n22934, Z => n22936);
   U25173 : NAND2_X1 port map( A1 => n22940, A2 => n27694, ZN => n22942);
   U25174 : INV_X2 port map( I => n32860, ZN => n23203);
   U25175 : XOR2_X1 port map( A1 => n23203, A2 => n1067, Z => n22954);
   U25177 : NOR2_X1 port map( A1 => n14129, A2 => n22965, ZN => n22966);
   U25178 : NAND2_X1 port map( A1 => n31935, A2 => n28680, ZN => n22996);
   U25179 : INV_X1 port map( I => n23007, ZN => n23008);
   U25180 : INV_X1 port map( I => n23011, ZN => n23012);
   U25181 : NOR2_X1 port map( A1 => n23013, A2 => n23012, ZN => n23014);
   U25182 : XOR2_X1 port map( A1 => n7070, A2 => n721, Z => n23023);
   U25184 : XOR2_X1 port map( A1 => n29217, A2 => n24833, Z => n23022);
   U25185 : XOR2_X1 port map( A1 => n23023, A2 => n23022, Z => n23024);
   U25187 : XOR2_X1 port map( A1 => n8659, A2 => n23376, Z => n23039);
   U25188 : XOR2_X1 port map( A1 => n27875, A2 => n25554, Z => n23038);
   U25189 : XOR2_X1 port map( A1 => n23038, A2 => n23039, Z => n23040);
   U25190 : NAND3_X1 port map( A1 => n27612, A2 => n1108, A3 => n28277, ZN => 
                           n23054);
   U25191 : NAND2_X1 port map( A1 => n1269, A2 => n26231, ZN => n23060);
   U25194 : XOR2_X1 port map( A1 => n23420, A2 => n16423, Z => n23076);
   U25195 : XOR2_X1 port map( A1 => n23075, A2 => n23076, Z => n23077);
   U25197 : NAND2_X1 port map( A1 => n14602, A2 => n17639, ZN => n23089);
   U25200 : XOR2_X1 port map( A1 => n24992, A2 => n11891, Z => n23118);
   U25201 : XOR2_X1 port map( A1 => n23122, A2 => n32893, Z => n23123);
   U25204 : XOR2_X1 port map( A1 => n13321, A2 => n16697, Z => n23139);
   U25205 : XOR2_X1 port map( A1 => n23344, A2 => n23139, Z => n23140);
   U25207 : XOR2_X1 port map( A1 => n24953, A2 => n3519, Z => n23146);
   U25210 : XOR2_X1 port map( A1 => n27763, A2 => n16666, Z => n23154);
   U25211 : INV_X1 port map( I => n23530, ZN => n23162);
   U25212 : XOR2_X1 port map( A1 => n32050, A2 => n23474, Z => n23163);
   U25216 : NAND2_X1 port map( A1 => n12658, A2 => n31796, ZN => n23177);
   U25217 : OAI21_X1 port map( A1 => n24385, A2 => n24383, B => n24384, ZN => 
                           n23179);
   U25218 : XOR2_X1 port map( A1 => n23420, A2 => n24231, Z => n23185);
   U25222 : XOR2_X1 port map( A1 => n3868, A2 => n25324, Z => n23198);
   U25223 : XOR2_X1 port map( A1 => n23454, A2 => n23346, Z => n23205);
   U25225 : XOR2_X1 port map( A1 => n24759, A2 => n23211, Z => n23212);
   U25226 : OAI21_X1 port map( A1 => n757, A2 => n32998, B => n23823, ZN => 
                           n23223);
   U25227 : XOR2_X1 port map( A1 => n23216, A2 => n24966, Z => n23217);
   U25228 : XOR2_X1 port map( A1 => n7045, A2 => n30315, Z => n23226);
   U25229 : XOR2_X1 port map( A1 => n23385, A2 => n23227, Z => n23228);
   U25230 : XOR2_X1 port map( A1 => n27875, A2 => n25282, Z => n23231);
   U25231 : XOR2_X1 port map( A1 => n32899, A2 => n16479, Z => n23232);
   U25233 : XOR2_X1 port map( A1 => n848, A2 => n25549, Z => n23243);
   U25234 : XOR2_X1 port map( A1 => n23250, A2 => n25910, Z => n23251);
   U25236 : XOR2_X1 port map( A1 => n24707, A2 => n11891, Z => n23268);
   U25237 : XOR2_X1 port map( A1 => n23298, A2 => n23268, Z => n23269);
   U25238 : XOR2_X1 port map( A1 => n5512, A2 => n5211, Z => n23278);
   U25239 : XOR2_X1 port map( A1 => n26656, A2 => n23287, Z => n23288);
   U25240 : XOR2_X1 port map( A1 => n27708, A2 => n23413, Z => n23303);
   U25241 : XOR2_X1 port map( A1 => n7363, A2 => n25311, Z => n23302);
   U25242 : XOR2_X1 port map( A1 => n23303, A2 => n23302, Z => n23304);
   U25243 : XOR2_X1 port map( A1 => n26656, A2 => n31513, Z => n23310);
   U25248 : XOR2_X1 port map( A1 => n23328, A2 => n25878, Z => n23329);
   U25249 : XOR2_X1 port map( A1 => n16160, A2 => n24514, Z => n23338);
   U25250 : NAND2_X1 port map( A1 => n23871, A2 => n27163, ZN => n24186);
   U25252 : NOR2_X1 port map( A1 => n23726, A2 => n23348, ZN => n23971);
   U25253 : NOR2_X1 port map( A1 => n23510, A2 => n23721, ZN => n23350);
   U25254 : NAND2_X1 port map( A1 => n23351, A2 => n16337, ZN => n23353);
   U25256 : XOR2_X1 port map( A1 => n16530, A2 => n23405, Z => n23356);
   U25258 : XOR2_X1 port map( A1 => n15130, A2 => n25206, Z => n23364);
   U25259 : XOR2_X1 port map( A1 => n23371, A2 => n25191, Z => n23372);
   U25260 : XOR2_X1 port map( A1 => n23373, A2 => n23372, Z => n23374);
   U25265 : INV_X1 port map( I => n23395, ZN => n23396);
   U25266 : XOR2_X1 port map( A1 => n33971, A2 => n23396, Z => n23397);
   U25267 : XOR2_X1 port map( A1 => n16631, A2 => n23405, Z => n23406);
   U25269 : XOR2_X1 port map( A1 => n23420, A2 => n25493, Z => n23421);
   U25272 : XOR2_X1 port map( A1 => n23429, A2 => n23430, Z => n23432);
   U25273 : XOR2_X1 port map( A1 => n33293, A2 => n24937, Z => n23431);
   U25274 : XOR2_X1 port map( A1 => n23431, A2 => n23432, Z => n23433);
   U25275 : XOR2_X1 port map( A1 => n27708, A2 => n16612, Z => n23436);
   U25276 : XOR2_X1 port map( A1 => n23467, A2 => n25560, Z => n23468);
   U25277 : INV_X1 port map( I => n23485, ZN => n23481);
   U25278 : INV_X1 port map( I => n23479, ZN => n23483);
   U25279 : NOR2_X1 port map( A1 => n23483, A2 => n25545, ZN => n23480);
   U25280 : OAI21_X1 port map( A1 => n23481, A2 => n23482, B => n23480, ZN => 
                           n23487);
   U25281 : NOR2_X1 port map( A1 => n23482, A2 => n15816, ZN => n23484);
   U25282 : AOI22_X1 port map( A1 => n23485, A2 => n23484, B1 => n23483, B2 => 
                           n25545, ZN => n23486);
   U25283 : XOR2_X1 port map( A1 => n982, A2 => n23511, Z => n23512);
   U25284 : XOR2_X1 port map( A1 => n31554, A2 => n8487, Z => n23513);
   U25287 : XOR2_X1 port map( A1 => n10773, A2 => n24869, Z => n23523);
   U25288 : XOR2_X1 port map( A1 => n23524, A2 => n23523, Z => n23525);
   U25289 : NAND2_X1 port map( A1 => n26290, A2 => n23527, ZN => n23528);
   U25293 : NAND2_X1 port map( A1 => n23540, A2 => n13343, ZN => n23548);
   U25294 : XOR2_X1 port map( A1 => n23552, A2 => n23551, Z => n23553);
   U25295 : XOR2_X1 port map( A1 => n23554, A2 => n23553, Z => n24359);
   U25301 : NAND2_X1 port map( A1 => n16186, A2 => n23917, ZN => n23573);
   U25307 : NOR2_X1 port map( A1 => n23770, A2 => n23768, ZN => n23598);
   U25308 : AOI21_X1 port map( A1 => n23778, A2 => n11392, B => n23775, ZN => 
                           n23604);
   U25309 : NAND3_X1 port map( A1 => n24220, A2 => n1096, A3 => n24218, ZN => 
                           n23606);
   U25310 : NAND2_X1 port map( A1 => n791, A2 => n24219, ZN => n23605);
   U25312 : NOR2_X1 port map( A1 => n24289, A2 => n24110, ZN => n23618);
   U25317 : NAND3_X1 port map( A1 => n16388, A2 => n29272, A3 => n28510, ZN => 
                           n23636);
   U25322 : INV_X1 port map( I => n23655, ZN => n23656);
   U25324 : NAND2_X1 port map( A1 => n13308, A2 => n11621, ZN => n23670);
   U25325 : MUX2_X1 port map( I0 => n24142, I1 => n24144, S => n319, Z => 
                           n23680);
   U25329 : NAND2_X1 port map( A1 => n13549, A2 => n1253, ZN => n23676);
   U25338 : OAI21_X1 port map( A1 => n29269, A2 => n23527, B => n23717, ZN => 
                           n23718);
   U25339 : NAND3_X1 port map( A1 => n23765, A2 => n1101, A3 => n23352, ZN => 
                           n23724);
   U25340 : INV_X1 port map( I => n23728, ZN => n23731);
   U25343 : MUX2_X1 port map( I0 => n23735, I1 => n29865, S => n23736, Z => 
                           n23740);
   U25344 : AOI21_X2 port map( A1 => n23740, A2 => n28676, B => n23739, ZN => 
                           n24072);
   U25347 : NAND3_X1 port map( A1 => n23776, A2 => n8547, A3 => n23775, ZN => 
                           n23780);
   U25348 : XOR2_X1 port map( A1 => n24638, A2 => n16705, Z => n23790);
   U25350 : NOR2_X1 port map( A1 => n14975, A2 => n16238, ZN => n23784);
   U25353 : NAND2_X1 port map( A1 => n23797, A2 => n23857, ZN => n23799);
   U25357 : INV_X1 port map( I => n23868, ZN => n23869);
   U25358 : NAND2_X1 port map( A1 => n23870, A2 => n31179, ZN => n23978);
   U25360 : INV_X1 port map( I => n23929, ZN => n23922);
   U25361 : INV_X1 port map( I => n23928, ZN => n23921);
   U25364 : INV_X1 port map( I => n23966, ZN => n23969);
   U25365 : INV_X1 port map( I => n23967, ZN => n23968);
   U25366 : INV_X1 port map( I => n23971, ZN => n23972);
   U25367 : NAND3_X1 port map( A1 => n23974, A2 => n23973, A3 => n23972, ZN => 
                           n23975);
   U25370 : INV_X1 port map( I => n24183, ZN => n23994);
   U25374 : XOR2_X1 port map( A1 => n24992, A2 => n24520, Z => n24021);
   U25379 : NOR2_X1 port map( A1 => n24305, A2 => n14252, ZN => n24032);
   U25380 : NAND2_X1 port map( A1 => n24114, A2 => n24040, ZN => n24041);
   U25381 : XOR2_X1 port map( A1 => n24513, A2 => n31687, Z => n24049);
   U25382 : XOR2_X1 port map( A1 => n24049, A2 => n24048, Z => n24050);
   U25384 : INV_X1 port map( I => n24065, ZN => n24993);
   U25388 : MUX2_X1 port map( I0 => n33540, I1 => n33680, S => n24243, Z => 
                           n24076);
   U25389 : NAND3_X1 port map( A1 => n890, A2 => n10987, A3 => n24326, ZN => 
                           n24081);
   U25390 : NOR2_X1 port map( A1 => n890, A2 => n24128, ZN => n24082);
   U25392 : XOR2_X1 port map( A1 => n24786, A2 => n12969, Z => n24089);
   U25395 : XOR2_X1 port map( A1 => n16679, A2 => n24622, Z => n24098);
   U25396 : NOR2_X1 port map( A1 => n24878, A2 => n24974, ZN => n24099);
   U25399 : INV_X1 port map( I => n24174, ZN => n24607);
   U25402 : NAND4_X1 port map( A1 => n24189, A2 => n24188, A3 => n24187, A4 => 
                           n24186, ZN => n24190);
   U25403 : NAND2_X1 port map( A1 => n9368, A2 => n32349, ZN => n24208);
   U25405 : XOR2_X1 port map( A1 => n24474, A2 => n24707, Z => n24215);
   U25406 : NAND2_X1 port map( A1 => n32737, A2 => n24225, ZN => n24227);
   U25407 : INV_X1 port map( I => n24231, ZN => n25259);
   U25408 : XOR2_X1 port map( A1 => n4728, A2 => n16636, Z => n24241);
   U25411 : NAND3_X1 port map( A1 => n24265, A2 => n31096, A3 => n16621, ZN => 
                           n24266);
   U25412 : XOR2_X1 port map( A1 => n25450, A2 => n11332, Z => n24267);
   U25413 : XOR2_X1 port map( A1 => n24394, A2 => n31687, Z => n24281);
   U25414 : XOR2_X1 port map( A1 => n24475, A2 => n25910, Z => n24280);
   U25417 : NAND2_X1 port map( A1 => n28240, A2 => n319, ZN => n24300);
   U25418 : NAND2_X1 port map( A1 => n24300, A2 => n1241, ZN => n24301);
   U25420 : INV_X1 port map( I => n24330, ZN => n24333);
   U25421 : INV_X1 port map( I => n24331, ZN => n24332);
   U25425 : XOR2_X1 port map( A1 => n25436, A2 => n24592, Z => n24355);
   U25431 : XOR2_X1 port map( A1 => n24761, A2 => n30540, Z => n24371);
   U25432 : INV_X1 port map( I => n24374, ZN => n25567);
   U25433 : NOR2_X1 port map( A1 => n25620, A2 => n25752, ZN => n24378);
   U25436 : XOR2_X1 port map( A1 => n24686, A2 => n25086, Z => n24387);
   U25437 : XOR2_X1 port map( A1 => n24814, A2 => n24391, Z => n24392);
   U25441 : XOR2_X1 port map( A1 => n25218, A2 => n11868, Z => n24402);
   U25443 : XOR2_X1 port map( A1 => n24786, A2 => n25578, Z => n24410);
   U25444 : XOR2_X1 port map( A1 => n24411, A2 => n24410, Z => n24412);
   U25446 : XOR2_X1 port map( A1 => n887, A2 => n24620, Z => n24428);
   U25449 : XOR2_X1 port map( A1 => n24962, A2 => n24753, Z => n24444);
   U25451 : XOR2_X1 port map( A1 => n24453, A2 => n24547, Z => n24457);
   U25453 : INV_X1 port map( I => n16757, ZN => n25564);
   U25456 : OAI21_X1 port map( A1 => n18264, A2 => n8758, B => n32012, ZN => 
                           n24485);
   U25458 : XOR2_X1 port map( A1 => n24781, A2 => n24622, Z => n24491);
   U25459 : NAND2_X1 port map( A1 => n24498, A2 => n15409, ZN => n24501);
   U25460 : NAND2_X1 port map( A1 => n24499, A2 => n15409, ZN => n24500);
   U25462 : NAND2_X1 port map( A1 => n32798, A2 => n28136, ZN => n24506);
   U25464 : XOR2_X1 port map( A1 => n24660, A2 => n24514, Z => n24515);
   U25465 : XOR2_X1 port map( A1 => n24518, A2 => n24517, Z => n24519);
   U25467 : XOR2_X1 port map( A1 => n24522, A2 => n27385, Z => n24523);
   U25469 : OAI21_X1 port map( A1 => n16650, A2 => n25397, B => n25343, ZN => 
                           n24557);
   U25470 : XOR2_X1 port map( A1 => n24937, A2 => n24559, Z => n24560);
   U25475 : NOR2_X1 port map( A1 => n11409, A2 => n24570, ZN => n24584);
   U25476 : INV_X1 port map( I => n24572, ZN => n24583);
   U25477 : NAND2_X1 port map( A1 => n33761, A2 => n25229, ZN => n24580);
   U25478 : MUX2_X1 port map( I0 => n24581, I1 => n24580, S => n32864, Z => 
                           n24582);
   U25482 : NOR2_X1 port map( A1 => n24969, A2 => n24970, ZN => n24615);
   U25485 : INV_X1 port map( I => n24623, ZN => n25065);
   U25488 : INV_X1 port map( I => n24655, ZN => n24657);
   U25489 : XOR2_X1 port map( A1 => n24658, A2 => n24659, Z => n24662);
   U25491 : INV_X1 port map( I => n24664, ZN => n24665);
   U25492 : XOR2_X1 port map( A1 => n31713, A2 => n24665, Z => n24666);
   U25499 : INV_X1 port map( I => Key(10), ZN => n25864);
   U25500 : XOR2_X1 port map( A1 => n24836, A2 => n24686, Z => n24688);
   U25502 : INV_X1 port map( I => n16523, ZN => n24696);
   U25503 : XOR2_X1 port map( A1 => n24698, A2 => n24697, Z => n24699);
   U25505 : NAND3_X2 port map( A1 => n24704, A2 => n24703, A3 => n24702, ZN => 
                           n25478);
   U25506 : NOR2_X1 port map( A1 => n25403, A2 => n25400, ZN => n24705);
   U25507 : INV_X1 port map( I => n25701, ZN => n24713);
   U25509 : NOR2_X1 port map( A1 => n25816, A2 => n11003, ZN => n24721);
   U25510 : INV_X1 port map( I => n25804, ZN => n25805);
   U25511 : NAND2_X1 port map( A1 => n25805, A2 => n4450, ZN => n24720);
   U25514 : XOR2_X1 port map( A1 => n24741, A2 => n24999, Z => n24742);
   U25515 : XOR2_X1 port map( A1 => n24743, A2 => n24742, Z => n24744);
   U25516 : XOR2_X1 port map( A1 => n24745, A2 => n24744, Z => n25022);
   U25518 : XOR2_X1 port map( A1 => n30307, A2 => n25500, Z => n24757);
   U25521 : XOR2_X1 port map( A1 => n24801, A2 => n16622, Z => n24802);
   U25522 : XOR2_X1 port map( A1 => n24817, A2 => n24818, Z => n24822);
   U25523 : XOR2_X1 port map( A1 => n24819, A2 => n25288, Z => n24820);
   U25524 : XOR2_X1 port map( A1 => n12800, A2 => n24833, Z => n24834);
   U25526 : XOR2_X1 port map( A1 => n31713, A2 => n24869, Z => n24848);
   U25527 : NAND2_X1 port map( A1 => n25148, A2 => n17005, ZN => n24856);
   U25529 : XOR2_X1 port map( A1 => n24862, A2 => n24861, Z => Ciphertext(149))
                           ;
   U25531 : INV_X1 port map( I => n25529, ZN => n24865);
   U25533 : NAND2_X1 port map( A1 => n15046, A2 => n11898, ZN => n24876);
   U25534 : NAND2_X1 port map( A1 => n15046, A2 => n24973, ZN => n24879);
   U25536 : OR2_X1 port map( A1 => n27651, A2 => n25019, Z => n24882);
   U25537 : NAND3_X1 port map( A1 => n25019, A2 => n5202, A3 => n560, ZN => 
                           n24886);
   U25539 : NAND3_X1 port map( A1 => n24884, A2 => n25114, A3 => n16025, ZN => 
                           n24885);
   U25542 : NAND3_X1 port map( A1 => n1201, A2 => n24938, A3 => n965, ZN => 
                           n24897);
   U25544 : NOR3_X1 port map( A1 => n24905, A2 => n10755, A3 => n24902, ZN => 
                           n24899);
   U25545 : AOI21_X1 port map( A1 => n24916, A2 => n24908, B => n24899, ZN => 
                           n24901);
   U25546 : XOR2_X1 port map( A1 => n24901, A2 => n28575, Z => Ciphertext(1));
   U25547 : OAI22_X1 port map( A1 => n24928, A2 => n24927, B1 => n24936, B2 => 
                           n24926, ZN => n24929);
   U25548 : AOI21_X1 port map( A1 => n24931, A2 => n24930, B => n24929, ZN => 
                           n24932);
   U25549 : XOR2_X1 port map( A1 => n24932, A2 => n15409, Z => Ciphertext(10));
   U25550 : NAND2_X1 port map( A1 => n24939, A2 => n24938, ZN => n24942);
   U25551 : INV_X1 port map( I => n28662, ZN => n24940);
   U25552 : AOI22_X1 port map( A1 => n24942, A2 => n24955, B1 => n24941, B2 => 
                           n24940, ZN => n24945);
   U25553 : XOR2_X1 port map( A1 => n24945, A2 => n24944, Z => Ciphertext(12));
   U25554 : OAI21_X1 port map( A1 => n24948, A2 => n24947, B => n24946, ZN => 
                           n24949);
   U25557 : OAI21_X1 port map( A1 => n24958, A2 => n965, B => n24954, ZN => 
                           n24961);
   U25558 : NAND2_X1 port map( A1 => n24957, A2 => n24956, ZN => n24959);
   U25562 : XOR2_X1 port map( A1 => n25000, A2 => n1415, Z => Ciphertext(31));
   U25564 : NOR2_X1 port map( A1 => n25050, A2 => n25057, ZN => n25029);
   U25565 : NOR2_X1 port map( A1 => n25121, A2 => n8210, ZN => n25024);
   U25566 : NAND3_X1 port map( A1 => n25025, A2 => n25120, A3 => n25152, ZN => 
                           n25028);
   U25567 : NAND2_X1 port map( A1 => n25026, A2 => n16293, ZN => n25027);
   U25569 : NOR2_X1 port map( A1 => n32760, A2 => n32106, ZN => n25031);
   U25571 : OAI21_X1 port map( A1 => n25063, A2 => n25044, B => n25057, ZN => 
                           n25034);
   U25572 : NAND2_X1 port map( A1 => n25035, A2 => n25034, ZN => n25037);
   U25573 : XOR2_X1 port map( A1 => n25037, A2 => n25036, Z => Ciphertext(36));
   U25576 : NAND2_X1 port map( A1 => n25058, A2 => n25051, ZN => n25042);
   U25579 : MUX2_X1 port map( I0 => n25062, I1 => n31640, S => n25057, Z => 
                           n25053);
   U25580 : XOR2_X1 port map( A1 => n25055, A2 => n25054, Z => Ciphertext(40));
   U25582 : NAND2_X1 port map( A1 => n25078, A2 => n16809, ZN => n25070);
   U25585 : AOI21_X1 port map( A1 => n25105, A2 => n25100, B => n32857, ZN => 
                           n25084);
   U25587 : XOR2_X1 port map( A1 => n25087, A2 => n13331, Z => Ciphertext(48));
   U25588 : INV_X1 port map( I => n25088, ZN => n25090);
   U25590 : INV_X1 port map( I => n25094, ZN => n25095);
   U25591 : INV_X1 port map( I => n25185, ZN => n25183);
   U25593 : NAND2_X1 port map( A1 => n25187, A2 => n8219, ZN => n25132);
   U25596 : NOR2_X1 port map( A1 => n14627, A2 => n15641, ZN => n25143);
   U25597 : NAND2_X1 port map( A1 => n7765, A2 => n25175, ZN => n25155);
   U25598 : OAI22_X1 port map( A1 => n25180, A2 => n25153, B1 => n25158, B2 => 
                           n25155, ZN => n25157);
   U25599 : XOR2_X1 port map( A1 => n25157, A2 => n25156, Z => Ciphertext(61));
   U25600 : INV_X1 port map( I => n25161, ZN => n25162);
   U25601 : XOR2_X1 port map( A1 => n25163, A2 => n25162, Z => Ciphertext(62));
   U25602 : NAND2_X1 port map( A1 => n25165, A2 => n25175, ZN => n25166);
   U25603 : NAND3_X1 port map( A1 => n25170, A2 => n25169, A3 => n25168, ZN => 
                           n25171);
   U25607 : NOR2_X1 port map( A1 => n25339, A2 => n25232, ZN => n25196);
   U25608 : XOR2_X1 port map( A1 => n25219, A2 => n1414, Z => Ciphertext(76));
   U25609 : OAI21_X1 port map( A1 => n16650, A2 => n25400, B => n14246, ZN => 
                           n25231);
   U25610 : NOR2_X1 port map( A1 => n25253, A2 => n25237, ZN => n25248);
   U25611 : OAI21_X1 port map( A1 => n25977, A2 => n32601, B => n9162, ZN => 
                           n25243);
   U25612 : NAND3_X1 port map( A1 => n31268, A2 => n1224, A3 => n33493, ZN => 
                           n25245);
   U25613 : XOR2_X1 port map( A1 => n25255, A2 => n16602, Z => Ciphertext(82));
   U25614 : AOI21_X1 port map( A1 => n733, A2 => n25279, B => n25278, ZN => 
                           n25265);
   U25615 : NAND2_X1 port map( A1 => n25284, A2 => n28532, ZN => n25264);
   U25616 : NAND3_X1 port map( A1 => n13985, A2 => n25302, A3 => n25261, ZN => 
                           n25262);
   U25617 : XOR2_X1 port map( A1 => n25267, A2 => n26000, Z => Ciphertext(84));
   U25619 : NAND2_X1 port map( A1 => n25279, A2 => n25278, ZN => n25268);
   U25622 : NAND2_X1 port map( A1 => n16291, A2 => n25278, ZN => n25272);
   U25626 : OAI21_X1 port map( A1 => n7081, A2 => n11132, B => n25290, ZN => 
                           n25294);
   U25627 : NAND2_X1 port map( A1 => n11132, A2 => n25339, ZN => n25291);
   U25628 : NAND3_X1 port map( A1 => n17110, A2 => n25292, A3 => n25291, ZN => 
                           n25293);
   U25634 : NAND3_X1 port map( A1 => n17110, A2 => n32659, A3 => n25339, ZN => 
                           n25340);
   U25636 : NOR2_X1 port map( A1 => n25352, A2 => n25375, ZN => n25349);
   U25637 : INV_X1 port map( I => n25368, ZN => n25379);
   U25639 : NOR2_X1 port map( A1 => n25367, A2 => n25368, ZN => n25354);
   U25640 : NAND2_X1 port map( A1 => n25352, A2 => n25361, ZN => n25353);
   U25644 : NAND2_X1 port map( A1 => n30276, A2 => n25376, ZN => n25365);
   U25645 : NAND3_X1 port map( A1 => n30400, A2 => n30302, A3 => n25368, ZN => 
                           n25370);
   U25647 : AOI21_X1 port map( A1 => n25376, A2 => n25375, B => n30276, ZN => 
                           n25377);
   U25651 : NAND2_X1 port map( A1 => n25331, A2 => n25562, ZN => n25383);
   U25656 : OAI21_X1 port map( A1 => n25430, A2 => n25425, B => n25445, ZN => 
                           n25416);
   U25658 : NAND2_X1 port map( A1 => n16650, A2 => n25400, ZN => n25401);
   U25664 : XOR2_X1 port map( A1 => n25417, A2 => n1394, Z => Ciphertext(102));
   U25667 : NAND2_X1 port map( A1 => n25425, A2 => n25429, ZN => n25419);
   U25671 : AOI22_X1 port map( A1 => n29280, A2 => n25453, B1 => n25424, B2 => 
                           n25437, ZN => n25427);
   U25674 : NAND2_X1 port map( A1 => n29280, A2 => n25437, ZN => n25449);
   U25677 : NAND3_X1 port map( A1 => n25452, A2 => n25446, A3 => n25455, ZN => 
                           n25447);
   U25681 : NOR2_X1 port map( A1 => n25462, A2 => n6310, ZN => n25459);
   U25684 : XOR2_X1 port map( A1 => n25467, A2 => n1404, Z => n25468);
   U25685 : NAND3_X1 port map( A1 => n25468, A2 => n25470, A3 => n25475, ZN => 
                           n25485);
   U25686 : INV_X1 port map( I => n25482, ZN => n25472);
   U25692 : NAND3_X1 port map( A1 => n25477, A2 => n4183, A3 => n25476, ZN => 
                           n25481);
   U25693 : NAND3_X1 port map( A1 => n25479, A2 => n1404, A3 => n6310, ZN => 
                           n25480);
   U25695 : XOR2_X1 port map( A1 => n25494, A2 => n1065, Z => Ciphertext(113));
   U25696 : OAI21_X1 port map( A1 => n2480, A2 => n32897, B => n8766, ZN => 
                           n25499);
   U25697 : INV_X1 port map( I => n32897, ZN => n25495);
   U25698 : OAI21_X1 port map( A1 => n25499, A2 => n25498, B => n25497, ZN => 
                           n25501);
   U25699 : XOR2_X1 port map( A1 => n25501, A2 => n25500, Z => Ciphertext(114))
                           ;
   U25701 : NAND2_X1 port map( A1 => n749, A2 => n32897, ZN => n25514);
   U25702 : NAND2_X1 port map( A1 => n25561, A2 => n16783, ZN => n25522);
   U25706 : NAND2_X1 port map( A1 => n25550, A2 => n15134, ZN => n25543);
   U25707 : NAND3_X1 port map( A1 => n25550, A2 => n31647, A3 => n8320, ZN => 
                           n25547);
   U25709 : NAND2_X1 port map( A1 => n25707, A2 => n11944, ZN => n25579);
   U25711 : NAND3_X1 port map( A1 => n25593, A2 => n12042, A3 => n837, ZN => 
                           n25594);
   U25719 : NAND2_X1 port map( A1 => n11931, A2 => n25615, ZN => n25608);
   U25723 : XOR2_X1 port map( A1 => n25642, A2 => n16472, Z => Ciphertext(139))
                           ;
   U25731 : AOI21_X1 port map( A1 => n34094, A2 => n3883, B => n26322, ZN => 
                           n25667);
   U25732 : NAND3_X1 port map( A1 => n25691, A2 => n25687, A3 => n32879, ZN => 
                           n25672);
   U25735 : AOI21_X1 port map( A1 => n17120, A2 => n33976, B => n25760, ZN => 
                           n25676);
   U25736 : NAND3_X1 port map( A1 => n25680, A2 => n26447, A3 => n25679, ZN => 
                           n25683);
   U25738 : NAND3_X1 port map( A1 => n33386, A2 => n10376, A3 => n25731, ZN => 
                           n25718);
   U25739 : NAND2_X1 port map( A1 => n25719, A2 => n25718, ZN => n25721);
   U25740 : XOR2_X1 port map( A1 => n25721, A2 => n25720, Z => Ciphertext(152))
                           ;
   U25742 : NAND3_X1 port map( A1 => n25731, A2 => n16494, A3 => n25729, ZN => 
                           n25726);
   U25744 : OAI21_X1 port map( A1 => n13640, A2 => n16494, B => n25729, ZN => 
                           n25730);
   U25745 : NAND2_X1 port map( A1 => n25746, A2 => n32863, ZN => n25737);
   U25746 : OAI21_X1 port map( A1 => n25743, A2 => n27164, B => n25738, ZN => 
                           n25741);
   U25747 : INV_X1 port map( I => n25743, ZN => n25749);
   U25749 : NAND3_X1 port map( A1 => n25788, A2 => n25781, A3 => n12611, ZN => 
                           n25770);
   U25750 : NAND2_X1 port map( A1 => n25763, A2 => n146, ZN => n25764);
   U25751 : NOR2_X1 port map( A1 => n32874, A2 => n25795, ZN => n25798);
   U25752 : AOI21_X1 port map( A1 => n25775, A2 => n12611, B => n25774, ZN => 
                           n25776);
   U25753 : OAI21_X1 port map( A1 => n25798, A2 => n25777, B => n25776, ZN => 
                           n25778);
   U25754 : XOR2_X1 port map( A1 => n25778, A2 => n17063, Z => Ciphertext(164))
                           ;
   U25755 : INV_X1 port map( I => n25780, ZN => n25782);
   U25756 : INV_X1 port map( I => n25784, ZN => n25785);
   U25757 : OAI21_X1 port map( A1 => n11899, A2 => n25786, B => n25785, ZN => 
                           n25787);
   U25758 : NAND2_X1 port map( A1 => n25789, A2 => n25788, ZN => n25792);
   U25763 : XOR2_X1 port map( A1 => n25802, A2 => n25801, Z => Ciphertext(167))
                           ;
   U25764 : NOR2_X1 port map( A1 => n4450, A2 => n25804, ZN => n25803);
   U25765 : OAI21_X1 port map( A1 => n25823, A2 => n25805, B => n11003, ZN => 
                           n25808);
   U25766 : XOR2_X1 port map( A1 => n25810, A2 => n32981, Z => Ciphertext(170))
                           ;
   U25767 : NAND2_X1 port map( A1 => n25817, A2 => n25816, ZN => n25821);
   U25768 : AOI21_X1 port map( A1 => n25823, A2 => n25804, B => n25822, ZN => 
                           n25824);
   U25769 : OAI22_X1 port map( A1 => n25826, A2 => n25825, B1 => n9181, B2 => 
                           n25824, ZN => n25828);
   U25770 : XOR2_X1 port map( A1 => n25828, A2 => n25827, Z => Ciphertext(173))
                           ;
   U25771 : OAI21_X1 port map( A1 => n25834, A2 => n25851, B => n14199, ZN => 
                           n25830);
   U25772 : NOR3_X1 port map( A1 => n16673, A2 => n10897, A3 => n25851, ZN => 
                           n25829);
   U25774 : XOR2_X1 port map( A1 => n25833, A2 => n1064, Z => Ciphertext(174));
   U25775 : NOR2_X1 port map( A1 => n25851, A2 => n13049, ZN => n25835);
   U25776 : OAI22_X1 port map( A1 => n25836, A2 => n25852, B1 => n25835, B2 => 
                           n25853, ZN => n25837);
   U25777 : XOR2_X1 port map( A1 => n25837, A2 => n16654, Z => Ciphertext(175))
                           ;
   U25779 : NOR2_X1 port map( A1 => n25838, A2 => n25901, ZN => n25841);
   U25780 : NOR4_X1 port map( A1 => n25843, A2 => n31979, A3 => n25841, A4 => 
                           n25840, ZN => n25847);
   U25784 : INV_X1 port map( I => n25923, ZN => n25906);
   U25785 : MUX2_X1 port map( I0 => n25922, I1 => n25925, S => n25915, Z => 
                           n25909);
   U25787 : AOI21_X1 port map( A1 => n25923, A2 => n14359, B => n25922, ZN => 
                           n25924);
   U6220 : INV_X2 port map( I => n23944, ZN => n1256);
   U322 : INV_X2 port map( I => n23275, ZN => n721);
   U5017 : INV_X4 port map( I => n10302, ZN => n6003);
   U20459 : INV_X4 port map( I => n25232, ZN => n11132);
   U923 : INV_X2 port map( I => n19300, ZN => n730);
   U1607 : BUF_X2 port map( I => n22390, Z => n15260);
   U6339 : INV_X4 port map( I => n17394, ZN => n992);
   U7806 : INV_X4 port map( I => n28202, ZN => n24335);
   U944 : NAND2_X2 port map( A1 => n5119, A2 => n5118, ZN => n19103);
   U5101 : NAND2_X2 port map( A1 => n27619, A2 => n26445, ZN => n21550);
   U668 : NAND2_X2 port map( A1 => n21095, A2 => n9322, ZN => n12811);
   U1745 : NAND2_X2 port map( A1 => n725, A2 => n14540, ZN => n7746);
   U2920 : NAND2_X2 port map( A1 => n24120, A2 => n1775, ZN => n23791);
   U799 : INV_X2 port map( I => n20228, ZN => n20325);
   U6586 : NOR2_X2 port map( A1 => n19269, A2 => n19265, ZN => n19226);
   U203 : INV_X4 port map( I => n23540, ZN => n24114);
   U5929 : AOI21_X2 port map( A1 => n17239, A2 => n18922, B => n17238, ZN => 
                           n15991);
   U10570 : INV_X2 port map( I => n24198, ZN => n16712);
   U287 : INV_X4 port map( I => n13297, ZN => n23828);
   U4738 : BUF_X2 port map( I => n24360, Z => n25884);
   U4497 : OAI21_X2 port map( A1 => n2633, A2 => n2634, B => n23137, ZN => 
                           n2631);
   U8397 : AOI22_X2 port map( A1 => n20506, A2 => n14367, B1 => n10057, B2 => 
                           n20435, ZN => n6775);
   U107 : INV_X2 port map( I => n18156, ZN => n18154);
   U4429 : INV_X2 port map( I => n17535, ZN => n25711);
   U4446 : INV_X2 port map( I => n25962, ZN => n15770);
   U4784 : AOI22_X2 port map( A1 => n9813, A2 => n801, B1 => n9812, B2 => 
                           n27163, ZN => n5258);
   U990 : NAND2_X2 port map( A1 => n12327, A2 => n7164, ZN => n18577);
   U751 : AOI21_X2 port map( A1 => n11809, A2 => n125, B => n11808, ZN => 
                           n12147);
   U1673 : NAND2_X2 port map( A1 => n24925, A2 => n24927, ZN => n24922);
   U5851 : INV_X2 port map( I => n15733, ZN => n21379);
   U553 : OAI22_X2 port map( A1 => n11981, A2 => n21876, B1 => n13345, B2 => 
                           n8602, ZN => n21702);
   U208 : INV_X2 port map( I => n24234, ZN => n24130);
   U5996 : INV_X2 port map( I => n33094, ZN => n18006);
   U7575 : NOR2_X2 port map( A1 => n18005, A2 => n18470, ZN => n17253);
   U793 : NAND2_X2 port map( A1 => n15310, A2 => n15311, ZN => n20463);
   U23623 : INV_X2 port map( I => n16401, ZN => n17405);
   U803 : OAI21_X2 port map( A1 => n937, A2 => n28876, B => n27343, ZN => 
                           n19931);
   U4485 : NAND2_X2 port map( A1 => n8614, A2 => n23852, ZN => n12722);
   U859 : INV_X2 port map( I => n12517, ZN => n16298);
   U983 : INV_X2 port map( I => n18588, ZN => n17687);
   U304 : INV_X2 port map( I => n9199, ZN => n13773);
   U1001 : INV_X2 port map( I => n17030, ZN => n12956);
   U9851 : AOI22_X2 port map( A1 => n29423, A2 => n17495, B1 => n20052, B2 => 
                           n1358, ZN => n3827);
   U8103 : BUF_X2 port map( I => n9170, Z => n1842);
   U5052 : NAND2_X2 port map( A1 => n22997, A2 => n22996, ZN => n23489);
   U12247 : INV_X2 port map( I => n6215, ZN => n9549);
   U922 : BUF_X4 port map( I => n14233, Z => n29);
   U8115 : AOI21_X2 port map( A1 => n15315, A2 => n32076, B => n14822, ZN => 
                           n15314);
   U6685 : NOR2_X2 port map( A1 => n18798, A2 => n18797, ZN => n18896);
   U363 : NAND2_X2 port map( A1 => n31937, A2 => n4084, ZN => n23067);
   U118 : INV_X2 port map( I => n3339, ZN => n16589);
   U7276 : NAND2_X2 port map( A1 => n1355, A2 => n15282, ZN => n20506);
   U206 : NOR2_X2 port map( A1 => n15179, A2 => n24254, ZN => n17801);
   U9205 : INV_X2 port map( I => n14726, ZN => n23843);
   U8727 : NOR2_X2 port map( A1 => n9631, A2 => n8309, ZN => n10784);
   U9747 : OAI21_X2 port map( A1 => n5589, A2 => n5592, B => n27785, ZN => 
                           n5588);
   U1566 : NAND2_X2 port map( A1 => n2141, A2 => n24243, ZN => n24127);
   U4948 : NAND2_X2 port map( A1 => n15051, A2 => n1573, ZN => n2270);
   U5772 : OAI21_X2 port map( A1 => n15464, A2 => n3567, B => n10282, ZN => 
                           n10386);
   U529 : NOR2_X2 port map( A1 => n7641, A2 => n14541, ZN => n22047);
   U4575 : NOR2_X2 port map( A1 => n16512, A2 => n31874, ZN => n20880);
   U1907 : AOI21_X2 port map( A1 => n32064, A2 => n17162, B => n12549, ZN => 
                           n1871);
   U399 : OAI21_X2 port map( A1 => n11614, A2 => n17630, B => n22472, ZN => 
                           n23079);
   U9838 : NAND2_X2 port map( A1 => n13986, A2 => n8549, ZN => n20294);
   U6679 : INV_X4 port map( I => n5327, ZN => n951);
   U8704 : BUF_X2 port map( I => n10423, Z => n4017);
   U3581 : INV_X2 port map( I => n10414, ZN => n16789);
   U4253 : NAND2_X2 port map( A1 => n4645, A2 => n4644, ZN => n5625);
   U959 : INV_X2 port map( I => n10228, ZN => n10229);
   U569 : INV_X2 port map( I => n21767, ZN => n914);
   U403 : INV_X2 port map( I => n7881, ZN => n1275);
   U17706 : NOR2_X2 port map( A1 => n828, A2 => n28987, ZN => n11815);
   U4535 : INV_X2 port map( I => n10258, ZN => n16529);
   U1007 : NAND2_X2 port map( A1 => n829, A2 => n1188, ZN => n8788);
   U209 : INV_X4 port map( I => n9964, ZN => n16688);
   U839 : INV_X2 port map( I => n9724, ZN => n9748);
   U103 : INV_X2 port map( I => n17523, ZN => n25699);
   U6466 : BUF_X2 port map( I => n21375, Z => n16421);
   U747 : NAND2_X2 port map( A1 => n1351, A2 => n9025, ZN => n20406);
   U9357 : AOI21_X2 port map( A1 => n22431, A2 => n22626, B => n17123, ZN => 
                           n17122);
   U666 : INV_X2 port map( I => n11847, ZN => n12654);
   U11620 : OAI21_X2 port map( A1 => n12582, A2 => n12407, B => n10000, ZN => 
                           n14966);
   U8844 : BUF_X2 port map( I => Key(147), Z => n25815);
   U13130 : NOR2_X2 port map( A1 => n8212, A2 => n17370, ZN => n12892);
   U5370 : NAND2_X2 port map( A1 => n12338, A2 => n901, ZN => n22523);
   U1003 : INV_X2 port map( I => n16849, ZN => n4259);
   U4576 : INV_X2 port map( I => n21389, ZN => n21147);
   U2783 : INV_X1 port map( I => n21224, ZN => n8115);
   U5523 : INV_X2 port map( I => n18643, ZN => n4626);
   U5390 : OAI21_X2 port map( A1 => n9312, A2 => n9313, B => n17385, ZN => 
                           n2490);
   U565 : INV_X2 port map( I => n21122, ZN => n913);
   U117 : INV_X1 port map( I => n12358, ZN => n716);
   U241 : OAI21_X2 port map( A1 => n144, A2 => n10068, B => n23940, ZN => n2448
                           );
   U3422 : NAND2_X2 port map( A1 => n14280, A2 => n13379, ZN => n7228);
   U4804 : INV_X4 port map( I => n23806, ZN => n1100);
   U493 : INV_X2 port map( I => n31932, ZN => n11917);
   U232 : INV_X2 port map( I => n5317, ZN => n5318);
   U22011 : NAND2_X2 port map( A1 => n3891, A2 => n12586, ZN => n22834);
   U6492 : OAI21_X2 port map( A1 => n16174, A2 => n20515, B => n20517, ZN => 
                           n10731);
   U1170 : INV_X2 port map( I => n7746, ZN => n17149);
   U865 : INV_X4 port map( I => n16317, ZN => n15665);
   U9771 : AOI21_X2 port map( A1 => n12089, A2 => n20333, B => n12880, ZN => 
                           n12879);
   U730 : OAI21_X2 port map( A1 => n29444, A2 => n16070, B => n1157, ZN => 
                           n4772);
   U8662 : AOI22_X2 port map( A1 => n13806, A2 => n26350, B1 => n10700, B2 => 
                           n14312, ZN => n3920);
   U5401 : INV_X2 port map( I => n29523, ZN => n21859);
   U7302 : NAND2_X2 port map( A1 => n33091, A2 => n20158, ZN => n20333);
   U704 : INV_X2 port map( I => n6684, ZN => n21085);
   U13709 : NAND2_X2 port map( A1 => n11947, A2 => n9436, ZN => n25205);
   U7053 : OAI21_X2 port map( A1 => n8274, A2 => n21607, B => n21775, ZN => 
                           n21609);
   U353 : AOI21_X2 port map( A1 => n1274, A2 => n2580, B => n2579, ZN => n4543)
                           ;
   U5609 : OR2_X2 port map( A1 => n17499, A2 => n24447, Z => n17092);
   U8434 : NAND2_X2 port map( A1 => n1153, A2 => n28028, ZN => n14177);
   U236 : NOR2_X2 port map( A1 => n23170, A2 => n23169, ZN => n24060);
   U6618 : INV_X4 port map( I => n2080, ZN => n19315);
   U5657 : INV_X2 port map( I => n11041, ZN => n23714);
   U211 : INV_X2 port map( I => n18077, ZN => n17310);
   U4543 : INV_X2 port map( I => n22363, ZN => n22588);
   U1658 : OAI21_X2 port map( A1 => n23758, A2 => n23757, B => n28671, ZN => 
                           n11418);
   U4352 : INV_X2 port map( I => n27134, ZN => n1208);
   U491 : INV_X2 port map( I => n17140, ZN => n22428);
   U9729 : OAI21_X2 port map( A1 => n12010, A2 => n20321, B => n18078, ZN => 
                           n13851);
   U5805 : INV_X4 port map( I => n32082, ZN => n22576);
   U3614 : INV_X2 port map( I => n24002, ZN => n767);
   U10547 : NAND2_X2 port map( A1 => n6632, A2 => n6633, ZN => n3380);
   U6149 : NOR2_X2 port map( A1 => n3222, A2 => n24248, ZN => n14972);
   U698 : INV_X2 port map( I => n13921, ZN => n12747);
   U4989 : INV_X2 port map( I => n9163, ZN => n12039);
   U46 : NAND2_X2 port map( A1 => n9754, A2 => n1462, ZN => n25513);
   U7949 : AOI21_X2 port map( A1 => n23085, A2 => n22884, B => n17668, ZN => 
                           n8455);
   U8469 : INV_X4 port map( I => n32240, ZN => n1153);
   U342 : NAND2_X2 port map( A1 => n8226, A2 => n11467, ZN => n12181);
   U5184 : INV_X2 port map( I => n18139, ZN => n8376);
   U6593 : OAI21_X2 port map( A1 => n15050, A2 => n19248, B => n4591, ZN => 
                           n14757);
   U6564 : INV_X4 port map( I => n4577, ZN => n17670);
   U1623 : INV_X1 port map( I => n8558, ZN => n1617);
   U7660 : BUF_X2 port map( I => Key(113), Z => n25064);
   U11202 : INV_X1 port map( I => n22656, ZN => n1286);
   U4508 : INV_X4 port map( I => n1485, ZN => n22977);
   U5083 : INV_X2 port map( I => n632, ZN => n15752);
   U4627 : BUF_X4 port map( I => n5545, Z => n1053);
   U8705 : BUF_X4 port map( I => n19222, Z => n16185);
   U4849 : NAND2_X2 port map( A1 => n18210, A2 => n18209, ZN => n21646);
   U11253 : NAND2_X2 port map( A1 => n21276, A2 => n21277, ZN => n15385);
   U6485 : NAND2_X2 port map( A1 => n14731, A2 => n11086, ZN => n19826);
   U545 : INV_X2 port map( I => n21821, ZN => n1317);
   U10111 : OAI21_X2 port map( A1 => n18772, A2 => n5805, B => n18771, ZN => 
                           n5311);
   U5426 : OAI22_X2 port map( A1 => n20475, A2 => n33288, B1 => n7394, B2 => 
                           n12758, ZN => n12757);
   U9992 : NAND2_X2 port map( A1 => n19085, A2 => n1046, ZN => n18405);
   U8181 : INV_X1 port map( I => n8602, ZN => n8569);
   U571 : NAND2_X2 port map( A1 => n27532, A2 => n11401, ZN => n21643);
   U5264 : OAI22_X2 port map( A1 => n12054, A2 => n29866, B1 => n24153, B2 => 
                           n26314, ZN => n3918);
   U6665 : NOR2_X2 port map( A1 => n6295, A2 => n328, ZN => n9090);
   U3434 : INV_X4 port map( I => n17306, ZN => n834);
   U1283 : INV_X1 port map( I => n13020, ZN => n9346);
   U5923 : AOI21_X2 port map( A1 => n3391, A2 => n19603, B => n19195, ZN => 
                           n19780);
   U6584 : NAND2_X2 port map( A1 => n3390, A2 => n3389, ZN => n19603);
   U9483 : AOI21_X2 port map( A1 => n13188, A2 => n33322, B => n13187, ZN => 
                           n21725);
   U7493 : INV_X2 port map( I => n14624, ZN => n9423);
   U5153 : INV_X2 port map( I => n4632, ZN => n10831);
   U2517 : INV_X2 port map( I => n11966, ZN => n812);
   U8755 : NOR2_X2 port map( A1 => n18445, A2 => n18444, ZN => n2099);
   U7567 : OAI21_X2 port map( A1 => n18798, A2 => n7899, B => n17843, ZN => 
                           n18445);
   U7179 : INV_X2 port map( I => n11601, ZN => n12363);
   U15105 : OAI21_X2 port map( A1 => n12367, A2 => n12366, B => n1023, ZN => 
                           n12365);
   U5931 : NAND2_X2 port map( A1 => n13011, A2 => n13012, ZN => n13481);
   U1714 : NOR2_X2 port map( A1 => n6219, A2 => n21359, ZN => n10313);
   U7265 : INV_X4 port map( I => n31522, ZN => n1026);
   U769 : INV_X2 port map( I => n20445, ZN => n20381);
   U4236 : NAND2_X2 port map( A1 => n4361, A2 => n4360, ZN => n4362);
   U10216 : BUF_X2 port map( I => Key(182), Z => n25735);
   U961 : OAI21_X2 port map( A1 => n18766, A2 => n14284, B => n18765, ZN => 
                           n18769);
   U4639 : NAND2_X2 port map( A1 => n1183, A2 => n7216, ZN => n12327);
   U9749 : NAND2_X2 port map( A1 => n1026, A2 => n20257, ZN => n3556);
   U6621 : BUF_X4 port map( I => n16960, Z => n8862);
   U7609 : OR2_X2 port map( A1 => n17558, A2 => n16450, Z => n12989);
   U947 : INV_X2 port map( I => n16960, ZN => n19116);
   U5128 : INV_X2 port map( I => n20526, ZN => n868);
   U6414 : INV_X2 port map( I => n21581, ZN => n16127);
   U22830 : INV_X4 port map( I => n14339, ZN => n18073);
   U12115 : AOI21_X2 port map( A1 => n17422, A2 => n28707, B => n3018, ZN => 
                           n10909);
   U5062 : BUF_X4 port map( I => n13679, Z => n803);
   U6622 : OAI21_X2 port map( A1 => n12065, A2 => n18759, B => n15281, ZN => 
                           n19094);
   U5733 : INV_X2 port map( I => n23267, ZN => n14077);
   U5461 : INV_X2 port map( I => n19418, ZN => n20059);
   U9266 : INV_X2 port map( I => n985, ZN => n7047);
   U5079 : INV_X2 port map( I => n1299, ZN => n22388);
   U4614 : OAI21_X2 port map( A1 => n26081, A2 => n26518, B => n8211, ZN => 
                           n18668);
   U9046 : AOI21_X2 port map( A1 => n12353, A2 => n24152, B => n3903, ZN => 
                           n3902);
   U5820 : NAND3_X2 port map( A1 => n17983, A2 => n17982, A3 => n1652, ZN => 
                           n14642);
   U4744 : INV_X2 port map( I => n9164, ZN => n17824);
   U11568 : INV_X4 port map( I => n17971, ZN => n4518);
   U1700 : NAND2_X2 port map( A1 => n14244, A2 => n14247, ZN => n14243);
   U388 : INV_X2 port map( I => n6874, ZN => n9954);
   U465 : INV_X2 port map( I => n17518, ZN => n22690);
   U4898 : AOI22_X2 port map( A1 => n18877, A2 => n961, B1 => n14658, B2 => 
                           n18101, ZN => n18939);
   U225 : INV_X2 port map( I => n31155, ZN => n24225);
   U3574 : INV_X2 port map( I => n10284, ZN => n18871);
   U4076 : NAND2_X2 port map( A1 => n16982, A2 => n23117, ZN => n24763);
   U9945 : INV_X2 port map( I => n17662, ZN => n20142);
   U5173 : NOR2_X2 port map( A1 => n13202, A2 => n13201, ZN => n13673);
   U6083 : INV_X2 port map( I => n25118, ZN => n25116);
   U1823 : NAND2_X1 port map( A1 => n14344, A2 => n15406, ZN => n10);
   U4442 : INV_X2 port map( I => n11622, ZN => n11947);
   U4243 : INV_X2 port map( I => n9553, ZN => n15050);
   U6231 : AOI21_X2 port map( A1 => n4155, A2 => n27612, B => n6099, ZN => 
                           n5593);
   U4058 : OR2_X2 port map( A1 => n9120, A2 => n23668, Z => n15550);
   U7234 : INV_X2 port map( I => n32648, ZN => n2789);
   U6979 : NAND2_X2 port map( A1 => n5453, A2 => n5744, ZN => n5448);
   U896 : NAND2_X2 port map( A1 => n379, A2 => n9787, ZN => n7438);
   U953 : NAND2_X2 port map( A1 => n2684, A2 => n2683, ZN => n19020);
   U4651 : BUF_X2 port map( I => Key(0), Z => n25206);
   U511 : INV_X2 port map( I => n22047, ZN => n21996);
   U5943 : INV_X4 port map( I => n10700, ZN => n947);
   U10213 : INV_X2 port map( I => n10664, ZN => n10665);
   U6681 : AOI22_X2 port map( A1 => n12238, A2 => n6891, B1 => n18553, B2 => 
                           n18891, ZN => n14844);
   U1491 : NAND4_X1 port map( A1 => n24497, A2 => n16502, A3 => n24495, A4 => 
                           n24496, ZN => n24502);
   U3620 : INV_X4 port map( I => n676, ZN => n11306);
   U5791 : NOR2_X2 port map( A1 => n22537, A2 => n22428, ZN => n22407);
   U8401 : AOI21_X2 port map( A1 => n12139, A2 => n33154, B => n20455, ZN => 
                           n20458);
   U9303 : NOR2_X2 port map( A1 => n772, A2 => n25994, ZN => n22760);
   U4905 : CLKBUF_X4 port map( I => n12282, Z => n6783);
   U3905 : INV_X2 port map( I => n24117, ZN => n24223);
   U24874 : NAND2_X2 port map( A1 => n13921, A2 => n27193, ZN => n21336);
   U4382 : INV_X2 port map( I => n2536, ZN => n7273);
   U6540 : OAI21_X2 port map( A1 => n822, A2 => n3626, B => n13346, ZN => 
                           n20006);
   U5792 : BUF_X2 port map( I => n22589, Z => n16562);
   U7365 : NAND3_X2 port map( A1 => n6644, A2 => n14172, A3 => n20066, ZN => 
                           n6643);
   U14244 : NAND2_X1 port map( A1 => n22572, A2 => n1298, ZN => n14775);
   U7270 : OAI21_X2 port map( A1 => n8353, A2 => n16182, B => n7056, ZN => 
                           n7055);
   U5858 : NAND2_X2 port map( A1 => n4648, A2 => n4266, ZN => n20423);
   U18858 : AOI21_X2 port map( A1 => n16221, A2 => n28404, B => n8303, ZN => 
                           n16106);
   U4478 : INV_X2 port map( I => n5306, ZN => n9625);
   U5035 : INV_X2 port map( I => n23576, ZN => n14207);
   U843 : INV_X2 port map( I => n12182, ZN => n822);
   U897 : NAND2_X2 port map( A1 => n28386, A2 => n13390, ZN => n19281);
   U607 : NAND2_X2 port map( A1 => n14397, A2 => n7182, ZN => n21846);
   U3598 : NOR2_X2 port map( A1 => n7310, A2 => n3909, ZN => n8084);
   U6724 : BUF_X2 port map( I => Key(70), Z => n16697);
   U4023 : OR2_X1 port map( A1 => n893, A2 => n23834, Z => n12020);
   U4189 : INV_X2 port map( I => n7119, ZN => n21322);
   U2340 : INV_X1 port map( I => n22307, ZN => n16700);
   U6419 : AOI21_X2 port map( A1 => n1142, A2 => n5049, B => n5047, ZN => n9396
                           );
   U6573 : AOI21_X2 port map( A1 => n16336, A2 => n16335, B => n15239, ZN => 
                           n18937);
   U795 : BUF_X4 port map( I => n20305, Z => n15434);
   U1733 : INV_X2 port map( I => n19788, ZN => n20009);
   U6581 : NOR2_X2 port map( A1 => n19004, A2 => n7176, ZN => n7283);
   U18831 : INV_X1 port map( I => n8277, ZN => n23717);
   U855 : INV_X4 port map( I => n20009, ZN => n9876);
   U4185 : NAND3_X2 port map( A1 => n7667, A2 => n21429, A3 => n7430, ZN => 
                           n21614);
   U1629 : NAND2_X2 port map( A1 => n13872, A2 => n16327, ZN => n12626);
   U6139 : NAND2_X2 port map( A1 => n24154, A2 => n16799, ZN => n17112);
   U5261 : NOR2_X2 port map( A1 => n5632, A2 => n7778, ZN => n10104);
   U5428 : BUF_X4 port map( I => n14980, Z => n13300);
   U25416 : AOI21_X2 port map( A1 => n33444, A2 => n15520, B => n24010, ZN => 
                           n24296);
   U6650 : INV_X4 port map( I => n19330, ZN => n880);
   U4126 : INV_X2 port map( I => n3773, ZN => n17161);
   U659 : INV_X2 port map( I => n9663, ZN => n21441);
   U7952 : AOI21_X2 port map( A1 => n15915, A2 => n899, B => n22769, ZN => 
                           n15914);
   U24701 : NOR2_X2 port map( A1 => n420, A2 => n29069, ZN => n20403);
   U111 : INV_X2 port map( I => n6143, ZN => n25409);
   U4696 : AOI22_X2 port map( A1 => n25328, A2 => n25406, B1 => n25329, B2 => 
                           n25410, ZN => n6411);
   U18918 : NAND2_X1 port map( A1 => n13917, A2 => n10293, ZN => n13916);
   U5190 : INV_X2 port map( I => n18498, ZN => n18601);
   U4988 : INV_X1 port map( I => n25628, ZN => n755);
   U6706 : INV_X2 port map( I => n18293, ZN => n18605);
   U4193 : BUF_X2 port map( I => n26448, Z => n8757);
   U10790 : NOR2_X1 port map( A1 => n13068, A2 => n10993, ZN => n23539);
   U14983 : NAND2_X1 port map( A1 => n21261, A2 => n21054, ZN => n10656);
   U9585 : INV_X4 port map( I => n9076, ZN => n21730);
   U6568 : INV_X2 port map( I => n19375, ZN => n12998);
   U24604 : NAND2_X1 port map( A1 => n8558, A2 => n15593, ZN => n19896);
   U3797 : INV_X1 port map( I => n3933, ZN => n21143);
   U7139 : INV_X4 port map( I => n17416, ZN => n21812);
   U17871 : OAI21_X2 port map( A1 => n8735, A2 => n829, B => n8737, ZN => n8734
                           );
   U6412 : INV_X2 port map( I => n16327, ZN => n920);
   U6313 : NAND2_X2 port map( A1 => n12613, A2 => n7964, ZN => n11161);
   U4844 : INV_X2 port map( I => n16222, ZN => n15838);
   U466 : INV_X2 port map( I => n5975, ZN => n8409);
   U18231 : OAI21_X2 port map( A1 => n16185, A2 => n28147, B => n4, ZN => n7436
                           );
   U5217 : AOI22_X2 port map( A1 => n31974, A2 => n25633, B1 => n25582, B2 => 
                           n25632, ZN => n15599);
   U946 : INV_X2 port map( I => n19360, ZN => n19109);
   U20868 : INV_X1 port map( I => n21353, ZN => n21172);
   U13467 : AND2_X2 port map( A1 => n13272, A2 => n11720, Z => n12337);
   U5054 : NAND3_X2 port map( A1 => n22937, A2 => n27694, A3 => n30925, ZN => 
                           n22852);
   U1155 : BUF_X4 port map( I => n9159, Z => n7144);
   U9785 : AOI22_X2 port map( A1 => n5029, A2 => n16182, B1 => n32035, B2 => 
                           n20603, ZN => n5027);
   U14381 : INV_X4 port map( I => n3483, ZN => n5741);
   U3036 : INV_X1 port map( I => n24561, ZN => n304);
   U4847 : INV_X4 port map( I => n16278, ZN => n5546);
   U9323 : INV_X4 port map( I => n22785, ZN => n7310);
   U11601 : NAND2_X1 port map( A1 => n14266, A2 => n20531, ZN => n14262);
   U828 : NAND2_X2 port map( A1 => n10831, A2 => n563, ZN => n19855);
   U9690 : INV_X4 port map( I => n11915, ZN => n7830);
   U24170 : NAND3_X2 port map( A1 => n34140, A2 => n28757, A3 => n18642, ZN => 
                           n18278);
   U6251 : OAI21_X2 port map( A1 => n5972, A2 => n5252, B => n17161, ZN => 
                           n5971);
   U4178 : NAND2_X2 port map( A1 => n2569, A2 => n2568, ZN => n9999);
   U5125 : INV_X2 port map( I => n14720, ZN => n14719);
   U4388 : NOR2_X2 port map( A1 => n25639, A2 => n25638, ZN => n25640);
   U6219 : INV_X2 port map( I => n3874, ZN => n846);
   U6386 : NAND2_X2 port map( A1 => n1137, A2 => n21816, ZN => n21820);
   U4850 : INV_X2 port map( I => n21225, ZN => n15261);
   U6431 : NOR2_X2 port map( A1 => n164, A2 => n7430, ZN => n21120);
   U5358 : AOI21_X2 port map( A1 => n22605, A2 => n22604, B => n22603, ZN => 
                           n14045);
   U8626 : AOI22_X2 port map( A1 => n13377, A2 => n28386, B1 => n19359, B2 => 
                           n19229, ZN => n13940);
   U22241 : AOI21_X2 port map( A1 => n6511, A2 => n28935, B => n18912, ZN => 
                           n18914);
   U5464 : INV_X4 port map( I => n10059, ZN => n11959);
   U6187 : NAND2_X2 port map( A1 => n23756, A2 => n26115, ZN => n7885);
   U4197 : BUF_X2 port map( I => n21136, Z => n16034);
   U9907 : NAND2_X2 port map( A1 => n7804, A2 => n19450, ZN => n3309);
   U5675 : INV_X4 port map( I => n12841, ZN => n24052);
   U775 : NAND2_X2 port map( A1 => n20213, A2 => n14564, ZN => n20631);
   U5480 : BUF_X2 port map( I => n9319, Z => n4714);
   U16652 : NAND2_X2 port map( A1 => n26600, A2 => n16093, ZN => n19302);
   U7470 : AOI22_X2 port map( A1 => n12052, A2 => n26181, B1 => n19007, B2 => 
                           n19052, ZN => n19008);
   U7230 : INV_X2 port map( I => n26448, ZN => n1022);
   U7889 : INV_X4 port map( I => n667, ZN => n23901);
   U3525 : INV_X1 port map( I => n3994, ZN => n24924);
   U13316 : OAI21_X2 port map( A1 => n2479, A2 => n28853, B => n805, ZN => 
                           n2404);
   U1354 : NOR2_X2 port map( A1 => n2734, A2 => n2732, ZN => n2731);
   U5981 : NAND2_X2 port map( A1 => n13548, A2 => n13514, ZN => n15018);
   U4254 : OR2_X2 port map( A1 => n18585, A2 => n12191, Z => n11970);
   U3626 : INV_X2 port map( I => n27154, ZN => n6263);
   U47 : NAND2_X2 port map( A1 => n25151, A2 => n34057, ZN => n25172);
   U21608 : NOR2_X2 port map( A1 => n28836, A2 => n34052, ZN => n17228);
   U10187 : BUF_X2 port map( I => n16462, Z => n6295);
   U8464 : INV_X4 port map( I => n1636, ZN => n20523);
   U7605 : INV_X2 port map( I => n11918, ZN => n18714);
   U11939 : INV_X2 port map( I => n16777, ZN => n3486);
   U2928 : BUF_X4 port map( I => n18300, Z => n18722);
   U929 : INV_X2 port map( I => n18980, ZN => n19257);
   U8598 : NAND3_X2 port map( A1 => n761, A2 => n11959, A3 => n9724, ZN => 
                           n4050);
   U4265 : BUF_X2 port map( I => n11605, Z => n2990);
   U12972 : INV_X2 port map( I => n8741, ZN => n9665);
   U11537 : OR2_X2 port map( A1 => n16938, A2 => n16743, Z => n21087);
   U6008 : BUF_X2 port map( I => Key(126), Z => n16561);
   U7859 : INV_X4 port map( I => n23843, ZN => n5373);
   U17098 : NAND2_X2 port map( A1 => n7830, A2 => n6082, ZN => n8256);
   U9215 : INV_X4 port map( I => n5191, ZN => n6661);
   U8653 : NOR2_X2 port map( A1 => n8051, A2 => n16485, ZN => n8831);
   U6997 : NAND2_X2 port map( A1 => n8131, A2 => n3063, ZN => n22531);
   U10910 : AOI21_X2 port map( A1 => n17149, A2 => n17148, B => n4652, ZN => 
                           n4651);
   U3538 : INV_X4 port map( I => n22641, ZN => n906);
   U15433 : AOI21_X2 port map( A1 => n14478, A2 => n29360, B => n29626, ZN => 
                           n15328);
   U13792 : NAND2_X2 port map( A1 => n1350, A2 => n2843, ZN => n11838);
   U7154 : INV_X2 port map( I => n17956, ZN => n7238);
   U10041 : INV_X2 port map( I => n19280, ZN => n13377);
   U3275 : NAND2_X2 port map( A1 => n6071, A2 => n27947, ZN => n365);
   U8218 : OAI22_X2 port map( A1 => n5048, A2 => n16779, B1 => n1142, B2 => 
                           n5049, ZN => n13292);
   U63 : INV_X2 port map( I => n25397, ZN => n14247);
   U9143 : OAI21_X2 port map( A1 => n16540, A2 => n33103, B => n16539, ZN => 
                           n1819);
   U6644 : INV_X4 port map( I => n8802, ZN => n879);
   U9296 : INV_X2 port map( I => n11626, ZN => n8479);
   U4407 : OR3_X2 port map( A1 => n1224, A2 => n33493, A3 => n31268, Z => 
                           n25109);
   U10762 : AOI21_X2 port map( A1 => n13342, A2 => n23510, B => n23918, ZN => 
                           n8983);
   U7737 : OR2_X2 port map( A1 => n24870, A2 => n8492, Z => n25149);
   U24482 : OAI21_X2 port map( A1 => n20078, A2 => n1163, B => n19381, ZN => 
                           n19382);
   U4893 : NOR3_X2 port map( A1 => n9511, A2 => n29683, A3 => n9514, ZN => 
                           n9509);
   U18961 : NAND2_X1 port map( A1 => n15129, A2 => n16228, ZN => n21545);
   U151 : NAND3_X1 port map( A1 => n11963, A2 => n24212, A3 => n24211, ZN => 
                           n17420);
   U22628 : INV_X2 port map( I => n23855, ZN => n23797);
   U3609 : INV_X2 port map( I => n23860, ZN => n2752);
   U6352 : INV_X1 port map( I => n11629, ZN => n10931);
   U9066 : INV_X2 port map( I => n24244, ZN => n1233);
   U5096 : NAND3_X1 port map( A1 => n8584, A2 => n8360, A3 => n17472, ZN => 
                           n1772);
   U10086 : NAND2_X2 port map( A1 => n24, A2 => n8335, ZN => n19328);
   U7765 : AOI21_X2 port map( A1 => n9257, A2 => n7203, B => n15010, ZN => 
                           n9256);
   U564 : INV_X2 port map( I => n14691, ZN => n17139);
   U8646 : OAI21_X2 port map( A1 => n4218, A2 => n4217, B => n27818, ZN => 
                           n4361);
   U11986 : NAND2_X2 port map( A1 => n13938, A2 => n29437, ZN => n13937);
   U894 : NAND2_X2 port map( A1 => n8862, A2 => n24, ZN => n15397);
   U14002 : INV_X2 port map( I => n5035, ZN => n8967);
   U6698 : INV_X2 port map( I => n16420, ZN => n7899);
   U15307 : OR2_X2 port map( A1 => n21330, A2 => n7453, Z => n21429);
   U20976 : OAI21_X2 port map( A1 => n16016, A2 => n21781, B => n17021, ZN => 
                           n16014);
   U7573 : INV_X2 port map( I => n13514, ZN => n18793);
   U9409 : NOR2_X2 port map( A1 => n239, A2 => n904, ZN => n2794);
   U5245 : INV_X2 port map( I => n25385, ZN => n25331);
   U2658 : INV_X2 port map( I => n3629, ZN => n11691);
   U7013 : NAND2_X2 port map( A1 => n16884, A2 => n1296, ZN => n7817);
   U5272 : INV_X1 port map( I => n7778, ZN => n24012);
   U10253 : BUF_X2 port map( I => Key(134), Z => n24707);
   U5434 : INV_X2 port map( I => n4693, ZN => n1156);
   U9614 : NAND3_X2 port map( A1 => n8256, A2 => n27230, A3 => n1335, ZN => 
                           n1882);
   U4432 : NAND2_X2 port map( A1 => n24723, A2 => n25905, ZN => n25838);
   U5137 : AOI21_X2 port map( A1 => n19918, A2 => n19917, B => n19916, ZN => 
                           n20526);
   U20250 : INV_X2 port map( I => n10681, ZN => n17201);
   U14432 : INV_X2 port map( I => n276, ZN => n21522);
   U14547 : NAND2_X1 port map( A1 => n17056, A2 => n25996, ZN => n5634);
   U4258 : INV_X2 port map( I => n18631, ZN => n16352);
   U5515 : INV_X2 port map( I => n5473, ZN => n953);
   U5740 : AOI21_X2 port map( A1 => n12107, A2 => n27865, B => n6591, ZN => 
                           n14466);
   U7632 : INV_X2 port map( I => n16585, ZN => n18228);
   U11698 : NAND2_X2 port map( A1 => n11838, A2 => n15434, ZN => n10321);
   U5492 : INV_X2 port map( I => n5455, ZN => n825);
   U5134 : NAND2_X2 port map( A1 => n1815, A2 => n13772, ZN => n4693);
   U6509 : INV_X2 port map( I => n14564, ZN => n9062);
   U7280 : AOI22_X2 port map( A1 => n20323, A2 => n5471, B1 => n8268, B2 => 
                           n15661, ZN => n13850);
   U5206 : NAND2_X2 port map( A1 => n11019, A2 => n25915, ZN => n14170);
   U7898 : INV_X4 port map( I => n11821, ZN => n1257);
   U4238 : INV_X2 port map( I => n11302, ZN => n946);
   U7143 : NAND2_X2 port map( A1 => n21120, A2 => n21429, ZN => n21499);
   U11293 : NAND2_X2 port map( A1 => n8006, A2 => n34087, ZN => n1543);
   U21194 : NOR2_X2 port map( A1 => n19883, A2 => n8616, ZN => n17574);
   U7781 : OAI21_X2 port map( A1 => n15179, A2 => n27436, B => n24253, ZN => 
                           n3604);
   U16330 : INV_X2 port map( I => n9690, ZN => n5073);
   U9999 : AOI21_X2 port map( A1 => n19034, A2 => n19088, B => n10867, ZN => 
                           n7316);
   U4218 : INV_X2 port map( I => n20110, ZN => n19971);
   U3197 : INV_X2 port map( I => n25473, ZN => n25470);
   U7174 : INV_X2 port map( I => n13304, ZN => n17956);
   U995 : NAND2_X1 port map( A1 => n6890, A2 => n10669, ZN => n5560);
   U5742 : NOR2_X2 port map( A1 => n30960, A2 => n15851, ZN => n3689);
   U850 : INV_X2 port map( I => n20142, ZN => n20036);
   U10963 : OAI21_X2 port map( A1 => n11925, A2 => n16919, B => n32766, ZN => 
                           n16918);
   U8853 : BUF_X2 port map( I => Key(129), Z => n16578);
   U9577 : INV_X2 port map( I => n12452, ZN => n21673);
   U4756 : OAI22_X2 port map( A1 => n11064, A2 => n8731, B1 => n10687, B2 => 
                           n24223, ZN => n9966);
   U7147 : AOI22_X2 port map( A1 => n11487, A2 => n21255, B1 => n8757, B2 => 
                           n4633, ZN => n7754);
   U36 : INV_X2 port map( I => n7702, ZN => n25915);
   U19164 : AND2_X2 port map( A1 => n10058, A2 => n18139, Z => n9514);
   U830 : INV_X2 port map( I => n33264, ZN => n6961);
   U9694 : INV_X2 port map( I => n18049, ZN => n21428);
   U4399 : NOR2_X2 port map( A1 => n13052, A2 => n6425, ZN => n13051);
   U4979 : BUF_X4 port map( I => n25885, Z => n4318);
   U19124 : OR2_X1 port map( A1 => n20029, A2 => n19961, Z => n16923);
   U8092 : INV_X1 port map( I => n22662, ZN => n22660);
   U4907 : INV_X2 port map( I => n16782, ZN => n13738);
   U8972 : OAI21_X2 port map( A1 => n14922, A2 => n1213, B => n16169, ZN => 
                           n11786);
   U25538 : INV_X2 port map( I => n24883, ZN => n25114);
   U16068 : INV_X2 port map( I => n4718, ZN => n15038);
   U7166 : AOI21_X2 port map( A1 => n21369, A2 => n1148, B => n17522, ZN => 
                           n4786);
   U12107 : AOI21_X2 port map( A1 => n4043, A2 => n17874, B => n16358, ZN => 
                           n13502);
   U8345 : BUF_X2 port map( I => n6556, Z => n3236);
   U6932 : NAND2_X2 port map( A1 => n22814, A2 => n4678, ZN => n9844);
   U16468 : NOR3_X1 port map( A1 => n7224, A2 => n7225, A3 => n5239, ZN => 
                           n18137);
   U5983 : NOR2_X2 port map( A1 => n18676, A2 => n12290, ZN => n18553);
   U13028 : INV_X2 port map( I => n15502, ZN => n19269);
   U323 : AND2_X2 port map( A1 => n5971, A2 => n11669, Z => n11668);
   U18570 : INV_X4 port map( I => n7965, ZN => n17764);
   U4295 : BUF_X2 port map( I => Key(170), Z => n16598);
   U4502 : BUF_X4 port map( I => n13415, Z => n5381);
   U22012 : AOI21_X2 port map( A1 => n29435, A2 => n21763, B => n21762, ZN => 
                           n21764);
   U716 : INV_X2 port map( I => n28813, ZN => n1023);
   U1854 : INV_X4 port map( I => n6416, ZN => n15902);
   U7407 : AND2_X2 port map( A1 => n10863, A2 => n571, Z => n12075);
   U3589 : OAI21_X2 port map( A1 => n29435, A2 => n21762, B => n6751, ZN => 
                           n12845);
   U16150 : INV_X1 port map( I => n22110, ZN => n13802);
   U10970 : NAND2_X1 port map( A1 => n3826, A2 => n27984, ZN => n10970);
   U23233 : AOI22_X2 port map( A1 => n15335, A2 => n16072, B1 => n4989, B2 => 
                           n21406, ZN => n21299);
   U7423 : INV_X4 port map( I => n20156, ZN => n940);
   U11267 : INV_X2 port map( I => n8291, ZN => n1310);
   U4688 : INV_X2 port map( I => n5412, ZN => n25922);
   U9003 : INV_X4 port map( I => n9127, ZN => n5387);
   U7582 : NAND2_X2 port map( A1 => n15108, A2 => n18018, ZN => n18574);
   U16901 : INV_X4 port map( I => n25981, ZN => n5834);
   U18746 : INV_X2 port map( I => n15009, ZN => n14457);
   U16955 : AOI21_X2 port map( A1 => n5896, A2 => n22606, B => n2858, ZN => 
                           n5958);
   U23056 : INV_X4 port map( I => n22427, ZN => n22534);
   U696 : INV_X2 port map( I => n17731, ZN => n1332);
   U3424 : INV_X4 port map( I => n19942, ZN => n1164);
   U19059 : OAI21_X1 port map( A1 => n8710, A2 => n8709, B => n8708, ZN => 
                           n8707);
   U22888 : NAND2_X1 port map( A1 => n29216, A2 => n28876, ZN => n14479);
   U8083 : INV_X1 port map( I => n645, ZN => n22368);
   U6893 : BUF_X2 port map( I => n14398, Z => n8525);
   U15560 : OR2_X2 port map( A1 => n10390, A2 => n8469, Z => n21061);
   U9891 : NOR2_X2 port map( A1 => n10072, A2 => n20149, ZN => n5550);
   U4687 : INV_X4 port map( I => n15483, ZN => n16041);
   U4715 : INV_X2 port map( I => n9941, ZN => n2886);
   U8634 : NAND2_X1 port map( A1 => n2599, A2 => n2935, ZN => n2598);
   U4173 : BUF_X2 port map( I => n21630, Z => n16601);
   U8852 : BUF_X2 port map( I => Key(108), Z => n25878);
   U4652 : CLKBUF_X2 port map( I => Key(39), Z => n25167);
   U12251 : BUF_X2 port map( I => Key(22), Z => n16551);
   U12265 : BUF_X2 port map( I => Key(112), Z => n16454);
   U4654 : CLKBUF_X2 port map( I => Key(84), Z => n16612);
   U7662 : BUF_X2 port map( I => Key(154), Z => n16605);
   U8869 : BUF_X2 port map( I => Key(109), Z => n25038);
   U6000 : BUF_X2 port map( I => Key(130), Z => n25450);
   U4290 : CLKBUF_X2 port map( I => Key(123), Z => n24487);
   U4276 : CLKBUF_X2 port map( I => Key(88), Z => n16631);
   U8866 : BUF_X2 port map( I => Key(114), Z => n25311);
   U8864 : BUF_X2 port map( I => Key(142), Z => n16674);
   U8845 : BUF_X2 port map( I => Key(48), Z => n25541);
   U6001 : BUF_X2 port map( I => Key(169), Z => n25355);
   U10252 : BUF_X2 port map( I => Key(76), Z => n25693);
   U4306 : CLKBUF_X2 port map( I => Key(34), Z => n16502);
   U4294 : CLKBUF_X2 port map( I => Key(184), Z => n8487);
   U5532 : BUF_X2 port map( I => Key(85), Z => n16523);
   U10223 : BUF_X2 port map( I => Key(31), Z => n16584);
   U4323 : CLKBUF_X2 port map( I => Key(52), Z => n16550);
   U7673 : BUF_X2 port map( I => Key(24), Z => n16619);
   U4301 : CLKBUF_X2 port map( I => Key(94), Z => n16355);
   U7674 : BUF_X2 port map( I => Key(90), Z => n16662);
   U5531 : BUF_X2 port map( I => Key(166), Z => n16604);
   U8862 : BUF_X2 port map( I => Key(138), Z => n25500);
   U12258 : BUF_X2 port map( I => Key(148), Z => n16636);
   U10232 : BUF_X2 port map( I => Key(61), Z => n25879);
   U2766 : CLKBUF_X2 port map( I => Key(173), Z => n16390);
   U8863 : BUF_X2 port map( I => Key(64), Z => n16322);
   U6012 : BUF_X2 port map( I => Key(49), Z => n24759);
   U10235 : BUF_X2 port map( I => Key(30), Z => n24833);
   U4319 : CLKBUF_X2 port map( I => Key(162), Z => n25641);
   U7669 : BUF_X2 port map( I => Key(172), Z => n16527);
   U4302 : CLKBUF_X2 port map( I => Key(3), Z => n24065);
   U4902 : BUF_X2 port map( I => n18882, Z => n17477);
   U2900 : INV_X1 port map( I => n270, ZN => n17597);
   U6717 : CLKBUF_X4 port map( I => n17189, Z => n1439);
   U4267 : CLKBUF_X2 port map( I => n11905, Z => n4194);
   U12253 : INV_X1 port map( I => n16504, ZN => n1392);
   U12252 : INV_X1 port map( I => n25274, ZN => n1391);
   U979 : INV_X2 port map( I => n18485, ZN => n18767);
   U12179 : CLKBUF_X1 port map( I => n12120, Z => n16426);
   U12118 : INV_X1 port map( I => n13466, ZN => n18749);
   U10080 : INV_X2 port map( I => n4392, ZN => n5813);
   U1929 : CLKBUF_X4 port map( I => n8802, Z => n24);
   U5176 : INV_X2 port map( I => n33986, ZN => n764);
   U21483 : NAND2_X1 port map( A1 => n19354, A2 => n19355, ZN => n14708);
   U23965 : NAND2_X1 port map( A1 => n18904, A2 => n32932, ZN => n17606);
   U10005 : NAND2_X1 port map( A1 => n824, A2 => n10229, ZN => n10855);
   U21154 : NAND2_X1 port map( A1 => n15869, A2 => n18449, ZN => n15418);
   U1531 : AOI21_X1 port map( A1 => n19366, A2 => n19365, B => n19364, ZN => 
                           n19367);
   U11931 : CLKBUF_X2 port map( I => n10696, Z => n4233);
   U11885 : INV_X1 port map( I => n5267, ZN => n5405);
   U8558 : NAND2_X1 port map( A1 => n20111, A2 => n32408, ZN => n7580);
   U11742 : INV_X1 port map( I => n20576, ZN => n7706);
   U788 : INV_X2 port map( I => n15043, ZN => n20338);
   U1243 : CLKBUF_X4 port map( I => n20339, Z => n384);
   U8386 : NAND2_X1 port map( A1 => n20554, A2 => n20553, ZN => n20557);
   U24702 : NAND2_X1 port map( A1 => n20540, A2 => n782, ZN => n20408);
   U4579 : NOR2_X1 port map( A1 => n1961, A2 => n6134, ZN => n1960);
   U2571 : AOI21_X1 port map( A1 => n5835, A2 => n15898, B => n184, ZN => n183)
                           ;
   U4581 : BUF_X4 port map( I => n20968, Z => n5024);
   U7228 : BUF_X2 port map( I => n20931, Z => n21365);
   U23648 : INV_X2 port map( I => n21189, ZN => n21419);
   U23736 : NOR2_X1 port map( A1 => n28642, A2 => n1017, ZN => n21065);
   U8200 : NAND2_X1 port map( A1 => n8457, A2 => n21736, ZN => n21737);
   U11317 : NAND2_X1 port map( A1 => n9350, A2 => n27532, ZN => n9448);
   U9489 : NAND3_X1 port map( A1 => n21753, A2 => n1316, A3 => n21752, ZN => 
                           n21757);
   U11270 : NAND2_X1 port map( A1 => n6937, A2 => n6935, ZN => n6600);
   U5091 : INV_X1 port map( I => n22100, ZN => n9290);
   U16077 : INV_X1 port map( I => n15825, ZN => n22214);
   U4160 : CLKBUF_X2 port map( I => n15606, Z => n3977);
   U4545 : BUF_X2 port map( I => n22662, Z => n16483);
   U8095 : BUF_X2 port map( I => n22412, Z => n16240);
   U4152 : CLKBUF_X2 port map( I => n21869, Z => n16447);
   U4137 : BUF_X2 port map( I => n22565, Z => n16490);
   U11173 : BUF_X2 port map( I => n11986, Z => n4100);
   U9442 : INV_X1 port map( I => n15805, ZN => n22663);
   U11197 : NOR2_X1 port map( A1 => n12530, A2 => n22403, ZN => n22333);
   U4539 : INV_X2 port map( I => n16166, ZN => n22484);
   U8043 : NOR2_X1 port map( A1 => n8098, A2 => n1842, ZN => n7662);
   U4121 : CLKBUF_X4 port map( I => n14600, Z => n897);
   U1887 : INV_X2 port map( I => n23103, ZN => n11399);
   U25186 : INV_X1 port map( I => n23027, ZN => n23029);
   U9246 : NAND2_X1 port map( A1 => n10790, A2 => n30573, ZN => n4780);
   U1109 : CLKBUF_X2 port map( I => n14612, Z => n6461);
   U7910 : BUF_X2 port map( I => n11205, Z => n8659);
   U1307 : INV_X1 port map( I => n23246, ZN => n5316);
   U5048 : INV_X1 port map( I => n13216, ZN => n11776);
   U4106 : CLKBUF_X2 port map( I => n23925, Z => n16121);
   U25290 : NAND2_X1 port map( A1 => n23691, A2 => n23857, ZN => n23543);
   U10827 : BUF_X2 port map( I => n17245, Z => n13549);
   U10719 : INV_X1 port map( I => n7524, ZN => n9137);
   U196 : INV_X2 port map( I => n4821, ZN => n14399);
   U17285 : INV_X2 port map( I => n24177, ZN => n8062);
   U5678 : INV_X2 port map( I => n24060, ZN => n792);
   U25391 : NAND2_X1 port map( A1 => n24139, A2 => n24141, ZN => n24086);
   U194 : NAND2_X1 port map( A1 => n17277, A2 => n24288, ZN => n3767);
   U10609 : NOR2_X1 port map( A1 => n794, A2 => n16356, ZN => n17066);
   U13127 : INV_X1 port map( I => n13306, ZN => n24277);
   U10508 : INV_X1 port map( I => n24842, ZN => n3544);
   U5594 : BUF_X2 port map( I => n11973, Z => n8307);
   U3559 : CLKBUF_X4 port map( I => n12871, Z => n12358);
   U18573 : INV_X2 port map( I => n13763, ZN => n9858);
   U6766 : NAND2_X1 port map( A1 => n4407, A2 => n33976, ZN => n8194);
   U8934 : NAND2_X1 port map( A1 => n7678, A2 => n8608, ZN => n7647);
   U1508 : OAI21_X1 port map( A1 => n3922, A2 => n15598, B => n25630, ZN => 
                           n15597);
   U8950 : NAND2_X1 port map( A1 => n25027, A2 => n25028, ZN => n1549);
   U10394 : OR2_X1 port map( A1 => n17782, A2 => n17778, Z => n14309);
   U8927 : CLKBUF_X4 port map( I => n25478, Z => n6310);
   U4689 : CLKBUF_X4 port map( I => n5412, Z => n5411);
   U25691 : NAND2_X1 port map( A1 => n25479, A2 => n6310, ZN => n25477);
   U10263 : INV_X1 port map( I => n10385, ZN => n10009);
   U10248 : CLKBUF_X2 port map( I => Key(55), Z => n16479);
   U4322 : BUF_X2 port map( I => Key(136), Z => n16482);
   U4318 : BUF_X2 port map( I => Key(139), Z => n25772);
   U4303 : BUF_X2 port map( I => Key(181), Z => n16613);
   U7672 : BUF_X2 port map( I => Key(73), Z => n23191);
   U4284 : BUF_X2 port map( I => Key(4), Z => n25218);
   U4307 : BUF_X2 port map( I => Key(16), Z => n16653);
   U8857 : BUF_X2 port map( I => Key(67), Z => n16649);
   U12269 : BUF_X2 port map( I => Key(186), Z => n16634);
   U4297 : BUF_X2 port map( I => Key(163), Z => n25908);
   U4908 : CLKBUF_X2 port map( I => Key(12), Z => n25266);
   U4277 : CLKBUF_X2 port map( I => Key(26), Z => n24907);
   U4282 : CLKBUF_X2 port map( I => Key(11), Z => n25009);
   U24366 : OAI21_X1 port map( A1 => n18775, A2 => n18774, B => n18773, ZN => 
                           n18776);
   U1367 : INV_X1 port map( I => n21662, ZN => n10345);
   U8056 : AOI21_X1 port map( A1 => n22503, A2 => n628, B => n3063, ZN => 
                           n11737);
   U1496 : INV_X1 port map( I => n22897, ZN => n10885);
   U10750 : INV_X1 port map( I => n23930, ZN => n9262);
   U9208 : NOR2_X1 port map( A1 => n7073, A2 => n17373, ZN => n3873);
   U134 : NAND2_X2 port map( A1 => n3547, A2 => n2361, ZN => n24370);
   U935 : BUF_X4 port map( I => n16047, Z => n5760);
   U11576 : INV_X2 port map( I => n8028, ZN => n5394);
   U11426 : OAI21_X2 port map( A1 => n21382, A2 => n21383, B => n15985, ZN => 
                           n21386);
   U7592 : OAI21_X2 port map( A1 => n18755, A2 => n18605, B => n18761, ZN => 
                           n18607);
   U22408 : INV_X2 port map( I => n17970, ZN => n18638);
   U11312 : OAI21_X2 port map( A1 => n8706, A2 => n8705, B => n34087, ZN => 
                           n2355);
   U21769 : INV_X4 port map( I => n26891, ZN => n16485);
   U9724 : OAI21_X2 port map( A1 => n12809, A2 => n28085, B => n12808, ZN => 
                           n20287);
   U17395 : AOI22_X2 port map( A1 => n14573, A2 => n14334, B1 => n16092, B2 => 
                           n14575, ZN => n14084);
   U21015 : OAI21_X2 port map( A1 => n20019, A2 => n16595, B => n14083, ZN => 
                           n14573);
   U5514 : NAND2_X1 port map( A1 => n16450, A2 => n17649, ZN => n5328);
   U22855 : INV_X2 port map( I => n31012, ZN => n18702);
   U8821 : NAND2_X1 port map( A1 => n18706, A2 => n18535, ZN => n18432);
   U22396 : INV_X2 port map( I => n13360, ZN => n16181);
   U2642 : INV_X1 port map( I => n18811, ZN => n7496);
   U1052 : INV_X2 port map( I => n18638, ZN => n955);
   U5192 : INV_X1 port map( I => n17649, ZN => n18572);
   U24268 : AOI21_X1 port map( A1 => n18848, A2 => n18845, B => n18730, ZN => 
                           n18409);
   U21441 : OAI21_X1 port map( A1 => n16995, A2 => n955, B => n14651, ZN => 
                           n14328);
   U12170 : AOI21_X1 port map( A1 => n28731, A2 => n4194, B => n27958, ZN => 
                           n10843);
   U6684 : NAND2_X1 port map( A1 => n18891, A2 => n6783, ZN => n14874);
   U10145 : NOR2_X1 port map( A1 => n18679, A2 => n10669, ZN => n5586);
   U20800 : INV_X1 port map( I => n12006, ZN => n18698);
   U5512 : NOR2_X1 port map( A1 => n10283, A2 => n10284, ZN => n18692);
   U5187 : NOR2_X1 port map( A1 => n32901, A2 => n12951, ZN => n18832);
   U7589 : AOI21_X1 port map( A1 => n16352, A2 => n31012, B => n18701, ZN => 
                           n13949);
   U13035 : NOR2_X1 port map( A1 => n2107, A2 => n962, ZN => n15694);
   U5972 : NOR2_X1 port map( A1 => n13466, A2 => n29659, ZN => n13110);
   U976 : AOI21_X1 port map( A1 => n18804, A2 => n17114, B => n11880, ZN => 
                           n18810);
   U14843 : NAND2_X1 port map( A1 => n18409, A2 => n18410, ZN => n3844);
   U7536 : OAI21_X1 port map( A1 => n14666, A2 => n15902, B => n10133, ZN => 
                           n10208);
   U5988 : OAI21_X1 port map( A1 => n14651, A2 => n18637, B => n18638, ZN => 
                           n5459);
   U20823 : OAI21_X1 port map( A1 => n18616, A2 => n12837, B => n10043, ZN => 
                           n18422);
   U5969 : NAND2_X1 port map( A1 => n7682, A2 => n7681, ZN => n18074);
   U7563 : INV_X1 port map( I => n12989, ZN => n18824);
   U12084 : INV_X1 port map( I => n19224, ZN => n1380);
   U8701 : INV_X2 port map( I => n4016, ZN => n12502);
   U924 : INV_X2 port map( I => n34107, ZN => n19228);
   U6625 : INV_X1 port map( I => n2150, ZN => n19096);
   U13321 : INV_X1 port map( I => n12468, ZN => n2412);
   U3309 : NAND3_X1 port map( A1 => n2150, A2 => n18769, A3 => n17905, ZN => 
                           n19200);
   U6608 : INV_X1 port map( I => n14597, ZN => n18993);
   U5493 : INV_X1 port map( I => n19348, ZN => n19217);
   U24430 : OAI22_X1 port map( A1 => n19076, A2 => n19196, B1 => n19075, B2 => 
                           n27726, ZN => n19077);
   U16522 : OAI21_X1 port map( A1 => n5813, A2 => n10203, B => n19200, ZN => 
                           n13890);
   U7520 : OAI21_X1 port map( A1 => n880, A2 => n19116, B => n879, ZN => n8864)
                           ;
   U22024 : NAND2_X1 port map( A1 => n4016, A2 => n19348, ZN => n16335);
   U1467 : NOR2_X1 port map( A1 => n19364, A2 => n19064, ZN => n19065);
   U18070 : NAND2_X1 port map( A1 => n1386, A2 => n11302, ZN => n7133);
   U9993 : INV_X1 port map( I => n18123, ZN => n3059);
   U9995 : NAND3_X1 port map( A1 => n9318, A2 => n19210, A3 => n4202, ZN => 
                           n9317);
   U4274 : BUF_X2 port map( I => Key(15), Z => n25049);
   U24295 : AOI21_X1 port map( A1 => n18474, A2 => n28147, B => n1378, ZN => 
                           n18478);
   U875 : INV_X1 port map( I => n4704, ZN => n8571);
   U11961 : CLKBUF_X2 port map( I => n19520, Z => n16586);
   U9959 : INV_X1 port map( I => n5127, ZN => n9988);
   U22449 : NAND2_X1 port map( A1 => n13477, A2 => n13480, ZN => n13479);
   U6003 : BUF_X2 port map( I => Key(190), Z => n16530);
   U1304 : INV_X1 port map( I => n19763, ZN => n1364);
   U13705 : NOR2_X1 port map( A1 => n2780, A2 => n20155, ZN => n13912);
   U7333 : NOR2_X1 port map( A1 => n5188, A2 => n19921, ZN => n1957);
   U2738 : BUF_X2 port map( I => n16646, Z => n12682);
   U2452 : INV_X1 port map( I => n6200, ZN => n10750);
   U22451 : NOR3_X1 port map( A1 => n19799, A2 => n19867, A3 => n19886, ZN => 
                           n13489);
   U5899 : INV_X1 port map( I => n18142, ZN => n20143);
   U7383 : NAND3_X1 port map( A1 => n1167, A2 => n20080, A3 => n1359, ZN => 
                           n2052);
   U5903 : INV_X1 port map( I => n565, ZN => n19794);
   U2873 : NOR2_X1 port map( A1 => n27655, A2 => n19900, ZN => n20111);
   U4220 : INV_X1 port map( I => n16105, ZN => n20013);
   U821 : INV_X1 port map( I => n8816, ZN => n1166);
   U14421 : NOR2_X1 port map( A1 => n11959, A2 => n5073, ZN => n3526);
   U1030 : AOI21_X1 port map( A1 => n20095, A2 => n579, B => n10439, ZN => 
                           n10394);
   U21027 : NAND3_X1 port map( A1 => n761, A2 => n3530, A3 => n15189, ZN => 
                           n13569);
   U11791 : NAND2_X1 port map( A1 => n20124, A2 => n20018, ZN => n17542);
   U9943 : OAI21_X1 port map( A1 => n14644, A2 => n19987, B => n5707, ZN => 
                           n20622);
   U21106 : INV_X1 port map( I => n20507, ZN => n17975);
   U9804 : NOR2_X1 port map( A1 => n1350, A2 => n2843, ZN => n20418);
   U24729 : NAND2_X1 port map( A1 => n7291, A2 => n20607, ZN => n20609);
   U21397 : NAND2_X1 port map( A1 => n20554, A2 => n7486, ZN => n13433);
   U4863 : INV_X1 port map( I => n20345, ZN => n760);
   U7272 : NOR2_X1 port map( A1 => n20517, A2 => n28011, ZN => n17297);
   U11707 : NOR2_X1 port map( A1 => n26424, A2 => n9025, ZN => n8869);
   U21403 : NOR2_X1 port map( A1 => n20334, A2 => n710, ZN => n12880);
   U11657 : OAI21_X1 port map( A1 => n782, A2 => n1863, B => n20342, ZN => 
                           n20349);
   U8417 : AOI22_X1 port map( A1 => n20531, A2 => n33721, B1 => n11055, B2 => 
                           n930, ZN => n11412);
   U24665 : NAND3_X1 port map( A1 => n111, A2 => n8998, A3 => n4468, ZN => 
                           n20217);
   U24718 : NAND3_X1 port map( A1 => n14731, A2 => n14719, A3 => n32747, ZN => 
                           n20504);
   U7282 : NAND2_X1 port map( A1 => n8868, A2 => n29628, ZN => n20350);
   U3031 : INV_X1 port map( I => n7330, ZN => n7960);
   U9682 : NAND2_X1 port map( A1 => n11733, A2 => n21391, ZN => n11732);
   U13593 : NOR2_X1 port map( A1 => n925, A2 => n1329, ZN => n2676);
   U5117 : NAND2_X1 port map( A1 => n601, A2 => n21221, ZN => n21060);
   U24848 : NAND3_X1 port map( A1 => n21147, A2 => n29901, A3 => n21218, ZN => 
                           n21148);
   U6426 : NOR3_X1 port map( A1 => n10837, A2 => n31614, A3 => n21387, ZN => 
                           n8560);
   U1500 : NOR2_X1 port map( A1 => n4274, A2 => n28668, ZN => n9816);
   U24801 : NAND2_X1 port map( A1 => n8028, A2 => n5395, ZN => n20909);
   U7195 : INV_X1 port map( I => n15874, ZN => n21289);
   U8253 : NAND3_X1 port map( A1 => n26971, A2 => n31614, A3 => n17956, ZN => 
                           n8170);
   U8249 : NAND2_X1 port map( A1 => n14853, A2 => n21151, ZN => n9378);
   U7199 : NOR2_X1 port map( A1 => n15002, A2 => n510, ZN => n9454);
   U630 : NAND2_X1 port map( A1 => n8170, A2 => n21148, ZN => n4863);
   U9572 : INV_X2 port map( I => n21789, ZN => n21653);
   U8228 : NAND2_X1 port map( A1 => n8457, A2 => n13652, ZN => n10357);
   U21419 : NAND2_X1 port map( A1 => n15838, A2 => n21653, ZN => n21467);
   U6407 : INV_X1 port map( I => n12827, ZN => n11394);
   U6404 : NAND2_X1 port map( A1 => n196, A2 => n27954, ZN => n21603);
   U4549 : OAI21_X1 port map( A1 => n11362, A2 => n10254, B => n26443, ZN => 
                           n14878);
   U9540 : AOI21_X1 port map( A1 => n16222, A2 => n21653, B => n21592, ZN => 
                           n3807);
   U9563 : INV_X1 port map( I => n21462, ZN => n21520);
   U9544 : OAI21_X1 port map( A1 => n3703, A2 => n17347, B => n1013, ZN => 
                           n3702);
   U8212 : NOR2_X1 port map( A1 => n14577, A2 => n14640, ZN => n21766);
   U7107 : NOR2_X1 port map( A1 => n1009, A2 => n2296, ZN => n15241);
   U1632 : OAI21_X1 port map( A1 => n17734, A2 => n29864, B => n28181, ZN => 
                           n21728);
   U11285 : NAND2_X1 port map( A1 => n27686, A2 => n13162, ZN => n13161);
   U9498 : AOI21_X1 port map( A1 => n21154, A2 => n21468, B => n21705, ZN => 
                           n21155);
   U11236 : INV_X1 port map( I => n9960, ZN => n11694);
   U8097 : INV_X2 port map( I => n4581, ZN => n16567);
   U21725 : INV_X1 port map( I => n22457, ZN => n22659);
   U6326 : INV_X1 port map( I => n8919, ZN => n4500);
   U21228 : NOR2_X1 port map( A1 => n9910, A2 => n26292, ZN => n18181);
   U463 : INV_X1 port map( I => n9592, ZN => n16745);
   U21801 : INV_X1 port map( I => n22428, ZN => n17626);
   U5782 : INV_X1 port map( I => n1125, ZN => n12236);
   U4834 : INV_X1 port map( I => n22610, ZN => n855);
   U17763 : INV_X1 port map( I => n16334, ZN => n17473);
   U5784 : AOI21_X1 port map( A1 => n22454, A2 => n22578, B => n15020, ZN => 
                           n15019);
   U9433 : NOR2_X1 port map( A1 => n468, A2 => n12733, ZN => n4560);
   U25095 : NAND2_X1 port map( A1 => n27638, A2 => n30014, ZN => n22502);
   U22129 : NAND3_X1 port map( A1 => n2471, A2 => n22574, A3 => n22657, ZN => 
                           n12887);
   U25059 : NOR2_X1 port map( A1 => n1842, A2 => n25947, ZN => n22325);
   U11195 : NOR2_X1 port map( A1 => n1001, A2 => n2132, ZN => n1523);
   U18985 : NAND2_X1 port map( A1 => n22650, A2 => n22651, ZN => n10928);
   U10938 : NOR2_X1 port map( A1 => n32766, A2 => n28313, ZN => n5096);
   U17711 : INV_X1 port map( I => n6605, ZN => n17327);
   U25137 : NAND2_X1 port map( A1 => n23043, A2 => n896, ZN => n22757);
   U7988 : INV_X1 port map( I => n3898, ZN => n17148);
   U391 : INV_X1 port map( I => n22655, ZN => n22895);
   U4816 : OAI21_X1 port map( A1 => n17161, A2 => n22977, B => n28227, ZN => 
                           n2078);
   U4505 : INV_X1 port map( I => n23262, ZN => n23443);
   U25120 : AOI21_X1 port map( A1 => n23158, A2 => n22693, B => n22692, ZN => 
                           n23425);
   U3610 : INV_X1 port map( I => n666, ZN => n23847);
   U22212 : NOR2_X1 port map( A1 => n14297, A2 => n23813, ZN => n13056);
   U6213 : INV_X1 port map( I => n4408, ZN => n16099);
   U3193 : INV_X2 port map( I => n23940, ZN => n23823);
   U22042 : INV_X1 port map( I => n28765, ZN => n23822);
   U7856 : NAND2_X1 port map( A1 => n895, A2 => n31890, ZN => n16211);
   U21286 : NAND2_X1 port map( A1 => n14164, A2 => n23578, ZN => n15642);
   U21285 : NAND2_X1 port map( A1 => n23824, A2 => n23825, ZN => n15615);
   U6898 : INV_X1 port map( I => n11922, ZN => n7895);
   U21320 : NOR2_X1 port map( A1 => n16496, A2 => n16343, ZN => n13364);
   U21291 : NAND3_X1 port map( A1 => n3241, A2 => n23848, A3 => n28365, ZN => 
                           n13173);
   U9186 : NOR2_X1 port map( A1 => n26641, A2 => n976, ZN => n14939);
   U12453 : OAI21_X1 port map( A1 => n1920, A2 => n15912, B => n26416, ZN => 
                           n5679);
   U21315 : INV_X1 port map( I => n24094, ZN => n24103);
   U181 : INV_X2 port map( I => n29977, ZN => n1237);
   U4473 : INV_X1 port map( I => n12904, ZN => n12903);
   U6830 : NAND2_X1 port map( A1 => n24315, A2 => n13232, ZN => n14336);
   U10579 : INV_X1 port map( I => n17801, ZN => n6632);
   U9096 : NAND3_X1 port map( A1 => n15179, A2 => n14399, A3 => n16868, ZN => 
                           n6633);
   U13663 : NAND2_X1 port map( A1 => n14663, A2 => n24316, ZN => n2745);
   U6121 : NAND2_X1 port map( A1 => n9581, A2 => n34137, ZN => n24059);
   U14790 : NAND3_X1 port map( A1 => n28120, A2 => n7068, A3 => n28784, ZN => 
                           n23989);
   U4750 : INV_X1 port map( I => n6484, ZN => n1230);
   U21085 : NAND2_X1 port map( A1 => n25897, A2 => n24607, ZN => n14108);
   U18574 : NAND2_X1 port map( A1 => n12042, A2 => n16397, ZN => n7973);
   U25737 : NAND2_X1 port map( A1 => n25701, A2 => n146, ZN => n25702);
   U21785 : INV_X1 port map( I => n17117, ZN => n24611);
   U6051 : NAND2_X1 port map( A1 => n25708, A2 => n16413, ZN => n13643);
   U1261 : OAI21_X1 port map( A1 => n25147, A2 => n25148, B => n25203, ZN => 
                           n9028);
   U21355 : INV_X1 port map( I => n25329, ZN => n24703);
   U5224 : NAND2_X1 port map( A1 => n25630, A2 => n8773, ZN => n11497);
   U8920 : NOR2_X1 port map( A1 => n27113, A2 => n5926, ZN => n10038);
   U21943 : NAND2_X1 port map( A1 => n25278, A2 => n12431, ZN => n17877);
   U2759 : INV_X1 port map( I => n7941, ZN => n5901);
   U8 : NAND3_X1 port map( A1 => n27113, A2 => n25577, A3 => n25575, ZN => 
                           n10039);
   U62 : NAND2_X1 port map( A1 => n13273, A2 => n14922, ZN => n3792);
   U100 : AND2_X1 port map( A1 => n1083, A2 => n25235, Z => n25134);
   U101 : AND2_X1 port map( A1 => n25695, A2 => n25628, Z => n6468);
   U119 : BUF_X2 port map( I => n25325, Z => n11366);
   U132 : NOR2_X1 port map( A1 => n3565, A2 => n9195, ZN => n26466);
   U136 : NAND2_X1 port map( A1 => n14495, A2 => n25119, ZN => n27625);
   U168 : INV_X1 port map( I => n24533, ZN => n7796);
   U182 : NAND3_X1 port map( A1 => n15876, A2 => n7150, A3 => n28296, ZN => 
                           n3545);
   U195 : NAND2_X1 port map( A1 => n23964, A2 => n10046, ZN => n27961);
   U245 : INV_X1 port map( I => n24072, ZN => n7891);
   U250 : BUF_X2 port map( I => n24014, Z => n16535);
   U259 : NOR2_X1 port map( A1 => n12904, A2 => n27430, ZN => n10778);
   U267 : OR2_X1 port map( A1 => n11041, A2 => n3421, Z => n11997);
   U297 : INV_X2 port map( I => n3880, ZN => n15011);
   U328 : OR2_X1 port map( A1 => n23918, A2 => n6869, Z => n26073);
   U339 : NAND2_X1 port map( A1 => n26716, A2 => n23675, ZN => n26211);
   U376 : OR2_X1 port map( A1 => n32998, A2 => n3004, Z => n26070);
   U382 : AOI22_X1 port map( A1 => n23902, A2 => n23843, B1 => n28034, B2 => 
                           n11067, ZN => n29081);
   U394 : OAI21_X1 port map( A1 => n23892, A2 => n32657, B => n26801, ZN => 
                           n23581);
   U398 : OR2_X1 port map( A1 => n16620, A2 => n4892, Z => n26074);
   U414 : NAND2_X1 port map( A1 => n28266, A2 => n29498, ZN => n26801);
   U441 : AOI21_X1 port map( A1 => n16343, A2 => n23832, B => n7005, ZN => 
                           n3448);
   U479 : CLKBUF_X2 port map( I => n29323, Z => n28297);
   U517 : NAND2_X1 port map( A1 => n4542, A2 => n4543, ZN => n29160);
   U540 : NAND2_X1 port map( A1 => n806, A2 => n4110, ZN => n26422);
   U547 : NOR2_X1 port map( A1 => n5982, A2 => n4399, ZN => n26994);
   U559 : NOR2_X1 port map( A1 => n22848, A2 => n31854, ZN => n22940);
   U572 : NAND2_X1 port map( A1 => n28680, A2 => n27752, ZN => n28327);
   U583 : OAI21_X1 port map( A1 => n29242, A2 => n27752, B => n22992, ZN => 
                           n9582);
   U618 : INV_X2 port map( I => n15704, ZN => n802);
   U683 : NAND2_X1 port map( A1 => n21972, A2 => n22277, ZN => n21975);
   U693 : AOI22_X1 port map( A1 => n22688, A2 => n2417, B1 => n6232, B2 => 
                           n2418, ZN => n28205);
   U703 : OR2_X1 port map( A1 => n22449, A2 => n16137, Z => n22973);
   U736 : OAI21_X1 port map( A1 => n10206, A2 => n28669, B => n32493, ZN => 
                           n1702);
   U754 : OR2_X1 port map( A1 => n6976, A2 => n1284, Z => n22449);
   U761 : NOR2_X1 port map( A1 => n27122, A2 => n22476, ZN => n27207);
   U789 : OAI21_X1 port map( A1 => n22670, A2 => n1127, B => n22558, ZN => 
                           n27357);
   U797 : NOR2_X1 port map( A1 => n22665, A2 => n22576, ZN => n15020);
   U824 : NAND2_X1 port map( A1 => n28924, A2 => n32078, ZN => n22420);
   U914 : OAI21_X1 port map( A1 => n3742, A2 => n26572, B => n13490, ZN => 
                           n5004);
   U915 : NAND3_X1 port map( A1 => n27707, A2 => n4331, A3 => n27706, ZN => 
                           n5075);
   U921 : NOR2_X1 port map( A1 => n26438, A2 => n21673, ZN => n26282);
   U962 : INV_X1 port map( I => n16194, ZN => n1325);
   U964 : NOR2_X1 port map( A1 => n21872, A2 => n7813, ZN => n13162);
   U982 : NOR2_X1 port map( A1 => n21865, A2 => n21738, ZN => n28068);
   U991 : NAND2_X1 port map( A1 => n27454, A2 => n17098, ZN => n11856);
   U1029 : AND2_X1 port map( A1 => n4234, A2 => n26163, Z => n12036);
   U1043 : NOR2_X1 port map( A1 => n1533, A2 => n21842, ZN => n27816);
   U1046 : NAND2_X1 port map( A1 => n14640, A2 => n29258, ZN => n15171);
   U1056 : INV_X1 port map( I => n15414, ZN => n1319);
   U1065 : NOR2_X1 port map( A1 => n21370, A2 => n26506, ZN => n26505);
   U1077 : NOR2_X1 port map( A1 => n13593, A2 => n21368, ZN => n26506);
   U1093 : AND2_X1 port map( A1 => n28668, A2 => n17341, Z => n11138);
   U1105 : NAND2_X1 port map( A1 => n17466, A2 => n27382, ZN => n27658);
   U1111 : NAND2_X1 port map( A1 => n9191, A2 => n15522, ZN => n26993);
   U1113 : NOR2_X1 port map( A1 => n4755, A2 => n17271, ZN => n2173);
   U1123 : NOR2_X1 port map( A1 => n5239, A2 => n8028, ZN => n26142);
   U1125 : NOR2_X1 port map( A1 => n6082, A2 => n21202, ZN => n14292);
   U1136 : NOR2_X1 port map( A1 => n29256, A2 => n4518, ZN => n26736);
   U1143 : NOR2_X1 port map( A1 => n21402, A2 => n12654, ZN => n28425);
   U1148 : AOI21_X1 port map( A1 => n17305, A2 => n4145, B => n17590, ZN => 
                           n12232);
   U1154 : NAND2_X1 port map( A1 => n21325, A2 => n21326, ZN => n27684);
   U1164 : NOR2_X1 port map( A1 => n2468, A2 => n5883, ZN => n26412);
   U1169 : INV_X1 port map( I => n21168, ZN => n27711);
   U1173 : NOR2_X1 port map( A1 => n21136, A2 => n31965, ZN => n28375);
   U1198 : NOR3_X1 port map( A1 => n6255, A2 => n6230, A3 => n26232, ZN => 
                           n19792);
   U1204 : NAND2_X1 port map( A1 => n20352, A2 => n1153, ZN => n26722);
   U1210 : NOR2_X1 port map( A1 => n17329, A2 => n17328, ZN => n12809);
   U1236 : AOI21_X1 port map( A1 => n20410, A2 => n20332, B => n6475, ZN => 
                           n7953);
   U1240 : AND2_X1 port map( A1 => n20345, A2 => n10717, Z => n20540);
   U1244 : AND2_X1 port map( A1 => n15230, A2 => n25966, Z => n5029);
   U1247 : NAND2_X1 port map( A1 => n2843, A2 => n14054, ZN => n20273);
   U1279 : OR2_X1 port map( A1 => n5781, A2 => n6610, Z => n27876);
   U1292 : OR2_X1 port map( A1 => n14179, A2 => n20450, Z => n5498);
   U1305 : BUF_X2 port map( I => n17236, Z => n29069);
   U1320 : NOR2_X1 port map( A1 => n28199, A2 => n27374, ZN => n27373);
   U1331 : NAND2_X1 port map( A1 => n28001, A2 => n875, ZN => n27569);
   U1332 : NAND3_X1 port map( A1 => n20043, A2 => n20157, A3 => n20156, ZN => 
                           n29225);
   U1339 : OR2_X1 port map( A1 => n28645, A2 => n26547, Z => n26007);
   U1346 : NAND2_X1 port map( A1 => n20068, A2 => n15110, ZN => n27716);
   U1349 : NAND3_X1 port map( A1 => n761, A2 => n20155, A3 => n3486, ZN => 
                           n19925);
   U1352 : NAND2_X1 port map( A1 => n729, A2 => n18126, ZN => n29034);
   U1356 : NAND2_X1 port map( A1 => n14589, A2 => n11959, ZN => n6067);
   U1363 : NAND2_X1 port map( A1 => n20147, A2 => n783, ZN => n27374);
   U1376 : NAND2_X1 port map( A1 => n15189, A2 => n20155, ZN => n9026);
   U1379 : AND2_X1 port map( A1 => n12179, A2 => n2391, Z => n26006);
   U1380 : NOR2_X1 port map( A1 => n8576, A2 => n27491, ZN => n9149);
   U1391 : NAND2_X1 port map( A1 => n12077, A2 => n14306, ZN => n9173);
   U1404 : NAND3_X1 port map( A1 => n19990, A2 => n12895, A3 => n28876, ZN => 
                           n3087);
   U1409 : NAND2_X1 port map( A1 => n579, A2 => n570, ZN => n28154);
   U1430 : NAND2_X1 port map( A1 => n11333, A2 => n575, ZN => n6859);
   U1434 : NOR2_X1 port map( A1 => n16193, A2 => n1161, ZN => n19939);
   U1437 : INV_X1 port map( I => n25997, ZN => n10805);
   U1449 : INV_X1 port map( I => n19399, ZN => n3195);
   U1453 : INV_X1 port map( I => n16349, ZN => n27825);
   U1463 : OAI21_X1 port map( A1 => n19260, A2 => n25971, B => n19257, ZN => 
                           n7419);
   U1480 : NOR2_X1 port map( A1 => n19261, A2 => n33206, ZN => n6343);
   U1483 : OAI22_X1 port map( A1 => n32932, A2 => n11000, B1 => n7492, B2 => 
                           n825, ZN => n26918);
   U1514 : OAI21_X1 port map( A1 => n28528, A2 => n10124, B => n3388, ZN => 
                           n19604);
   U1567 : BUF_X4 port map( I => n2150, Z => n26417);
   U1574 : OAI21_X1 port map( A1 => n26717, A2 => n18893, B => n13087, ZN => 
                           n18555);
   U1578 : OAI21_X1 port map( A1 => n13408, A2 => n4474, B => n4677, ZN => 
                           n28172);
   U1580 : NAND2_X1 port map( A1 => n18893, A2 => n10579, ZN => n28573);
   U1583 : NAND2_X1 port map( A1 => n7345, A2 => n14892, ZN => n1603);
   U1584 : OAI21_X1 port map( A1 => n18778, A2 => n18619, B => n16624, ZN => 
                           n15004);
   U1585 : AOI21_X1 port map( A1 => n12863, A2 => n10903, B => n7496, ZN => 
                           n18554);
   U1586 : AND2_X1 port map( A1 => n18805, A2 => n18806, Z => n26035);
   U1590 : OAI21_X1 port map( A1 => n18805, A2 => n18650, B => n27908, ZN => 
                           n9786);
   U1592 : NAND2_X1 port map( A1 => n3601, A2 => n27690, ZN => n9539);
   U1598 : OAI21_X1 port map( A1 => n18805, A2 => n17114, B => n17465, ZN => 
                           n27238);
   U1599 : NAND2_X1 port map( A1 => n27384, A2 => n6118, ZN => n6117);
   U1609 : NAND2_X1 port map( A1 => n25981, A2 => n18683, ZN => n19292);
   U1612 : NAND2_X1 port map( A1 => n18895, A2 => n16420, ZN => n27384);
   U1613 : NAND2_X1 port map( A1 => n26444, A2 => n6887, ZN => n4765);
   U1634 : NOR2_X1 port map( A1 => n18808, A2 => n16474, ZN => n27908);
   U1637 : NAND2_X1 port map( A1 => n18742, A2 => n18706, ZN => n18635);
   U1640 : NOR2_X1 port map( A1 => n12951, A2 => n12006, ZN => n13016);
   U1652 : BUF_X2 port map( I => n18780, Z => n16417);
   U1661 : OAI22_X2 port map( A1 => n30375, A2 => n20028, B1 => n16461, B2 => 
                           n16637, ZN => n19940);
   U1668 : INV_X2 port map( I => n4066, ZN => n6638);
   U1674 : NAND2_X2 port map( A1 => n18623, A2 => n27129, ZN => n11864);
   U1676 : NOR2_X1 port map( A1 => n18900, A2 => n28171, ZN => n28993);
   U1679 : INV_X2 port map( I => n19618, ZN => n20150);
   U1702 : INV_X2 port map( I => n22667, ZN => n13664);
   U1703 : INV_X2 port map( I => n22330, ZN => n22672);
   U1783 : OAI22_X2 port map( A1 => n20940, A2 => n3236, B1 => n5395, B2 => 
                           n7990, ZN => n5396);
   U1799 : AOI22_X2 port map( A1 => n1026, A2 => n7707, B1 => n7706, B2 => 
                           n26587, ZN => n7709);
   U1801 : NAND2_X1 port map( A1 => n3883, A2 => n734, ZN => n11213);
   U1835 : NAND2_X1 port map( A1 => n24585, A2 => n24588, ZN => n26217);
   U1839 : INV_X2 port map( I => n21992, ZN => n1714);
   U1856 : INV_X2 port map( I => n16267, ZN => n722);
   U1862 : BUF_X2 port map( I => n22679, Z => n16570);
   U1864 : AOI21_X2 port map( A1 => n5832, A2 => n31402, B => n722, ZN => 
                           n27451);
   U1865 : INV_X2 port map( I => n23866, ZN => n9741);
   U1871 : NAND3_X1 port map( A1 => n17333, A2 => n21712, A3 => n32904, ZN => 
                           n28995);
   U1917 : OAI21_X2 port map( A1 => n13170, A2 => n32298, B => n32299, ZN => 
                           n11675);
   U1935 : NAND2_X1 port map( A1 => n16955, A2 => n29180, ZN => n26370);
   U1939 : CLKBUF_X2 port map( I => n4908, Z => n27622);
   U1995 : NAND2_X1 port map( A1 => n9365, A2 => n25653, ZN => n7085);
   U2003 : OAI21_X1 port map( A1 => n10745, A2 => n10744, B => n25232, ZN => 
                           n10743);
   U2025 : BUF_X2 port map( I => n25723, Z => n9495);
   U2026 : INV_X1 port map( I => n27117, ZN => n17453);
   U2029 : CLKBUF_X2 port map( I => n27117, Z => n28784);
   U2033 : CLKBUF_X2 port map( I => n5544, Z => n5466);
   U2043 : NOR2_X1 port map( A1 => n4381, A2 => n28017, ZN => n21420);
   U2056 : OAI21_X1 port map( A1 => n5926, A2 => n6092, B => n25569, ZN => 
                           n6673);
   U2075 : NAND2_X1 port map( A1 => n14443, A2 => n6003, ZN => n17492);
   U2081 : CLKBUF_X2 port map( I => n2236, Z => n28734);
   U2090 : INV_X1 port map( I => n26848, ZN => n12643);
   U2123 : NOR2_X1 port map( A1 => n22619, A2 => n29314, ZN => n28320);
   U2140 : NOR2_X1 port map( A1 => n15011, A2 => n24141, ZN => n15052);
   U2143 : NOR2_X1 port map( A1 => n13627, A2 => n14960, ZN => n24967);
   U2149 : AND2_X1 port map( A1 => n12329, A2 => n32900, Z => n5867);
   U2174 : BUF_X2 port map( I => n24275, Z => n28120);
   U2176 : NAND2_X1 port map( A1 => n24277, A2 => n26247, ZN => n24278);
   U2178 : INV_X2 port map( I => n691, ZN => n13624);
   U2183 : AOI21_X1 port map( A1 => n24587, A2 => n753, B => n26217, ZN => 
                           n10609);
   U2184 : NAND2_X1 port map( A1 => n123, A2 => n17764, ZN => n13417);
   U2186 : AND2_X1 port map( A1 => n25062, A2 => n25057, Z => n3123);
   U2187 : AND2_X1 port map( A1 => n25063, A2 => n25062, Z => n16377);
   U2193 : OR2_X1 port map( A1 => n7915, A2 => n28343, Z => n23655);
   U2205 : OR3_X1 port map( A1 => n767, A2 => n24340, A3 => n24163, Z => n7091)
                           ;
   U2299 : NAND2_X1 port map( A1 => n25250, A2 => n7929, ZN => n15124);
   U2300 : NOR2_X1 port map( A1 => n25250, A2 => n7929, ZN => n5543);
   U2301 : NAND2_X1 port map( A1 => n7929, A2 => n25258, ZN => n25254);
   U2305 : OAI22_X1 port map( A1 => n25569, A2 => n13624, B1 => n25568, B2 => 
                           n6092, ZN => n6114);
   U2307 : NAND2_X1 port map( A1 => n9616, A2 => n5226, ZN => n24288);
   U2315 : NOR2_X1 port map( A1 => n8307, A2 => n25756, ZN => n26270);
   U2317 : OR2_X1 port map( A1 => n25709, A2 => n25756, Z => n26056);
   U2327 : NAND2_X1 port map( A1 => n25082, A2 => n11360, ZN => n25100);
   U2329 : NAND2_X1 port map( A1 => n25057, A2 => n25058, ZN => n27609);
   U2339 : NAND2_X1 port map( A1 => n3569, A2 => n547, ZN => n17023);
   U2363 : NOR2_X1 port map( A1 => n10097, A2 => n31921, ZN => n11181);
   U2364 : INV_X2 port map( I => n31921, ZN => n9862);
   U2370 : AOI21_X1 port map( A1 => n22626, A2 => n16170, B => n17955, ZN => 
                           n22627);
   U2374 : NOR2_X1 port map( A1 => n22982, A2 => n12586, ZN => n28318);
   U2385 : OR2_X1 port map( A1 => n29317, A2 => n13694, Z => n10293);
   U2396 : OR2_X1 port map( A1 => n10724, A2 => n17638, Z => n250);
   U2428 : NOR2_X1 port map( A1 => n13343, A2 => n4151, ZN => n17065);
   U2440 : NOR2_X1 port map( A1 => n23566, A2 => n769, ZN => n26464);
   U2443 : NOR2_X1 port map( A1 => n17373, A2 => n3874, ZN => n23675);
   U2447 : NOR2_X1 port map( A1 => n25900, A2 => n25867, ZN => n6981);
   U2453 : OAI21_X1 port map( A1 => n7935, A2 => n24157, B => n796, ZN => 
                           n17602);
   U2467 : NOR2_X1 port map( A1 => n1567, A2 => n2092, ZN => n27514);
   U2485 : INV_X1 port map( I => n25060, ZN => n25052);
   U2512 : AND2_X1 port map( A1 => n25699, A2 => n25696, Z => n12086);
   U2546 : OR2_X1 port map( A1 => n22816, A2 => n16315, Z => n15167);
   U2547 : INV_X1 port map( I => n24682, ZN => n9386);
   U2567 : NAND2_X1 port map( A1 => n5226, A2 => n11503, ZN => n17232);
   U2587 : NAND3_X1 port map( A1 => n9917, A2 => n25390, A3 => n24667, ZN => 
                           n14062);
   U2597 : OAI21_X1 port map( A1 => n17110, A2 => n25232, B => n5468, ZN => 
                           n6259);
   U2608 : BUF_X2 port map( I => n19624, Z => n27395);
   U2609 : OR2_X1 port map( A1 => n1511, A2 => n25973, Z => n1508);
   U2618 : NOR2_X1 port map( A1 => n21766, A2 => n6599, ZN => n3796);
   U2624 : NAND2_X1 port map( A1 => n12058, A2 => n1218, ZN => n24894);
   U2637 : NAND2_X1 port map( A1 => n15255, A2 => n17641, ZN => n8901);
   U2650 : INV_X2 port map( I => n31894, ZN => n23482);
   U2655 : NAND2_X1 port map( A1 => n7093, A2 => n24163, ZN => n2852);
   U2671 : INV_X1 port map( I => n25375, ZN => n25361);
   U2678 : NOR2_X1 port map( A1 => n20507, A2 => n16452, ZN => n17760);
   U2681 : BUF_X2 port map( I => n16831, Z => n28163);
   U2690 : INV_X1 port map( I => n12593, ZN => n24010);
   U2694 : CLKBUF_X4 port map( I => n22125, Z => n8356);
   U2700 : NAND3_X1 port map( A1 => n12005, A2 => n16152, A3 => n32298, ZN => 
                           n16409);
   U2715 : INV_X2 port map( I => n20819, ZN => n20658);
   U2716 : AND2_X1 port map( A1 => n19911, A2 => n12770, Z => n25941);
   U2732 : INV_X1 port map( I => n9159, ZN => n13345);
   U2733 : XOR2_X1 port map( A1 => n22121, A2 => n16622, Z => n25945);
   U2737 : INV_X2 port map( I => n10824, ZN => n22030);
   U2754 : INV_X2 port map( I => n14002, ZN => n23017);
   U2755 : INV_X1 port map( I => n22580, ZN => n9913);
   U2767 : NOR3_X2 port map( A1 => n12445, A2 => n17740, A3 => n12444, ZN => 
                           n27176);
   U2772 : INV_X2 port map( I => n23945, ZN => n1253);
   U2793 : NAND2_X2 port map( A1 => n27660, A2 => n27439, ZN => n27125);
   U2794 : INV_X2 port map( I => n24299, ZN => n24304);
   U2796 : INV_X1 port map( I => n25325, ZN => n25410);
   U2801 : INV_X2 port map( I => n25051, ZN => n28070);
   U2803 : INV_X2 port map( I => n31939, ZN => n27127);
   U2805 : NAND2_X2 port map( A1 => n11786, A2 => n13267, ZN => n27149);
   U2815 : NAND2_X1 port map( A1 => n802, A2 => n22876, ZN => n2028);
   U2825 : AND2_X1 port map( A1 => n14864, A2 => n13345, Z => n5078);
   U2846 : NAND2_X1 port map( A1 => n10717, A2 => n10106, ZN => n20342);
   U2853 : NOR2_X1 port map( A1 => n1718, A2 => n25628, ZN => n26563);
   U2864 : AND2_X1 port map( A1 => n25795, A2 => n8678, Z => n8676);
   U2880 : NAND2_X1 port map( A1 => n6544, A2 => n5546, ZN => n4358);
   U2898 : INV_X1 port map( I => n8533, ZN => n26493);
   U2906 : NOR2_X1 port map( A1 => n7811, A2 => n21872, ZN => n10492);
   U2909 : NAND2_X1 port map( A1 => n18727, A2 => n13279, ZN => n26398);
   U2910 : AND2_X2 port map( A1 => n18548, A2 => n18649, Z => n18804);
   U2939 : NAND2_X1 port map( A1 => n16194, A2 => n5016, ZN => n8360);
   U2951 : NAND2_X1 port map( A1 => n26244, A2 => n26242, ZN => n17083);
   U2955 : NAND2_X1 port map( A1 => n24251, A2 => n28553, ZN => n12551);
   U2977 : INV_X2 port map( I => n13614, ZN => n24421);
   U2987 : NAND3_X1 port map( A1 => n125, A2 => n12563, A3 => n20329, ZN => 
                           n12564);
   U2988 : NAND2_X1 port map( A1 => n15571, A2 => n24031, ZN => n15570);
   U3013 : NOR2_X1 port map( A1 => n15278, A2 => n20095, ZN => n15907);
   U3020 : CLKBUF_X1 port map( I => n19149, Z => n25959);
   U3022 : CLKBUF_X12 port map( I => n23944, Z => n16677);
   U3028 : INV_X1 port map( I => n15275, ZN => n26715);
   U3045 : NOR3_X1 port map( A1 => n32642, A2 => n21559, A3 => n6489, ZN => 
                           n8007);
   U3083 : NOR2_X1 port map( A1 => n12982, A2 => n3421, ZN => n27863);
   U3115 : NAND2_X1 port map( A1 => n17084, A2 => n23087, ZN => n26244);
   U3120 : NAND3_X1 port map( A1 => n26070, A2 => n31807, A3 => n33583, ZN => 
                           n2992);
   U3126 : NOR2_X1 port map( A1 => n19178, A2 => n29769, ZN => n27273);
   U3139 : AOI21_X1 port map( A1 => n12038, A2 => n25997, B => n19998, ZN => 
                           n26823);
   U3149 : AOI21_X2 port map( A1 => n17268, A2 => n11202, B => n34074, ZN => 
                           n10167);
   U3172 : NAND2_X1 port map( A1 => n12535, A2 => n28580, ZN => n12140);
   U3184 : NAND2_X1 port map( A1 => n3203, A2 => n21532, ZN => n12347);
   U3195 : AOI21_X1 port map( A1 => n14619, A2 => n16799, B => n839, ZN => 
                           n10112);
   U3253 : AND2_X2 port map( A1 => n15216, A2 => n15347, Z => n18543);
   U3259 : INV_X1 port map( I => n22970, ZN => n23259);
   U3279 : INV_X1 port map( I => n26750, ZN => n14373);
   U3290 : AND2_X2 port map( A1 => n21224, A2 => n14934, Z => n21317);
   U3307 : INV_X1 port map( I => n7810, ZN => n1050);
   U3308 : NAND3_X1 port map( A1 => n16274, A2 => n7810, A3 => n7680, ZN => 
                           n2585);
   U3312 : NAND2_X1 port map( A1 => n26806, A2 => n24244, ZN => n2324);
   U3319 : NAND2_X1 port map( A1 => n27685, A2 => n30832, ZN => n26283);
   U3322 : OR2_X2 port map( A1 => n10932, A2 => n14439, Z => n21451);
   U3328 : BUF_X4 port map( I => n22856, Z => n25979);
   U3342 : NAND2_X1 port map( A1 => n15829, A2 => n22990, ZN => n22619);
   U3343 : INV_X1 port map( I => n22990, ZN => n14977);
   U3373 : INV_X1 port map( I => n21232, ZN => n21132);
   U3376 : OR2_X2 port map( A1 => n21232, A2 => n21228, Z => n21302);
   U3377 : NAND2_X1 port map( A1 => n1289, A2 => n9617, ZN => n22336);
   U3380 : OAI21_X1 port map( A1 => n18146, A2 => n27430, B => n12903, ZN => 
                           n15571);
   U3396 : OAI21_X1 port map( A1 => n28157, A2 => n3340, B => n3515, ZN => 
                           n19003);
   U3428 : NAND2_X1 port map( A1 => n9630, A2 => n29288, ZN => n12613);
   U3451 : AND2_X2 port map( A1 => n10891, A2 => n495, Z => n18843);
   U3454 : INV_X1 port map( I => n495, ZN => n1389);
   U3457 : NAND2_X1 port map( A1 => n1318, A2 => n26439, ZN => n26438);
   U3475 : OAI22_X1 port map( A1 => n7219, A2 => n985, B1 => n7221, B2 => n9280
                           , ZN => n28402);
   U3487 : NAND3_X1 port map( A1 => n21284, A2 => n33889, A3 => n33147, ZN => 
                           n8866);
   U3490 : NOR2_X1 port map( A1 => n7068, A2 => n31461, ZN => n8665);
   U3493 : INV_X1 port map( I => n18076, ZN => n16372);
   U3494 : AOI22_X2 port map( A1 => n3522, A2 => n32021, B1 => n31551, B2 => 
                           n3521, ZN => n3520);
   U3512 : NAND3_X1 port map( A1 => n4071, A2 => n34013, A3 => n5275, ZN => 
                           n10290);
   U3517 : NAND3_X1 port map( A1 => n10106, A2 => n20344, A3 => n20345, ZN => 
                           n27225);
   U3519 : BUF_X2 port map( I => n7811, Z => n5383);
   U3529 : NAND2_X1 port map( A1 => n24276, A2 => n24168, ZN => n24167);
   U3532 : NAND2_X1 port map( A1 => n25066, A2 => n12329, ZN => n12487);
   U3533 : OAI21_X1 port map( A1 => n24139, A2 => n24138, B => n3880, ZN => 
                           n6978);
   U3539 : INV_X1 port map( I => n2643, ZN => n21468);
   U3566 : INV_X1 port map( I => n11217, ZN => n26540);
   U3567 : BUF_X4 port map( I => n10260, Z => n25985);
   U3602 : OAI21_X1 port map( A1 => n28659, A2 => n30904, B => n28318, ZN => 
                           n17175);
   U3605 : NAND2_X1 port map( A1 => n10360, A2 => n28697, ZN => n22985);
   U3634 : NAND2_X1 port map( A1 => n21070, A2 => n3192, ZN => n21328);
   U3641 : AND3_X2 port map( A1 => n21630, A2 => n21573, A3 => n21628, Z => 
                           n3798);
   U3647 : NOR2_X1 port map( A1 => n1327, A2 => n21707, ZN => n27648);
   U3768 : BUF_X2 port map( I => n10772, Z => n17906);
   U3772 : AND2_X2 port map( A1 => n33531, A2 => n15393, Z => n20148);
   U3814 : NAND2_X1 port map( A1 => n4755, A2 => n26345, ZN => n21081);
   U3832 : AOI21_X1 port map( A1 => n25410, A2 => n16528, B => n25411, ZN => 
                           n26892);
   U3843 : CLKBUF_X1 port map( I => n24276, Z => n26247);
   U3847 : AOI21_X1 port map( A1 => n27734, A2 => n23943, B => n13549, ZN => 
                           n23326);
   U3849 : NAND2_X1 port map( A1 => n23562, A2 => n33260, ZN => n7141);
   U3855 : NOR2_X1 port map( A1 => n23634, A2 => n28510, ZN => n28509);
   U3857 : CLKBUF_X1 port map( I => n9490, Z => n26290);
   U3872 : BUF_X2 port map( I => n31566, Z => n26231);
   U3875 : CLKBUF_X2 port map( I => n6593, Z => n27865);
   U3876 : BUF_X4 port map( I => n23051, Z => n25994);
   U3887 : CLKBUF_X2 port map( I => n10402, Z => n26292);
   U3897 : CLKBUF_X2 port map( I => n22036, Z => n28411);
   U3909 : CLKBUF_X1 port map( I => n14730, Z => n26899);
   U3911 : NAND2_X1 port map( A1 => n21850, A2 => n13490, ZN => n27005);
   U3918 : OAI21_X1 port map( A1 => n16147, A2 => n31958, B => n33766, ZN => 
                           n2720);
   U3922 : BUF_X2 port map( I => n16147, Z => n26904);
   U3937 : OAI21_X1 port map( A1 => n5026, A2 => n5030, B => n1160, ZN => n5025
                           );
   U3946 : NAND2_X1 port map( A1 => n17882, A2 => n1170, ZN => n4045);
   U3956 : CLKBUF_X2 port map( I => n6974, Z => n28889);
   U3981 : INV_X1 port map( I => n16649, ZN => n26002);
   U3990 : OAI22_X1 port map( A1 => n11134, A2 => n11136, B1 => n14510, B2 => 
                           n11133, ZN => n27047);
   U3992 : NAND3_X1 port map( A1 => n24946, A2 => n26199, A3 => n26197, ZN => 
                           n15249);
   U4001 : INV_X2 port map( I => n25723, ZN => n16494);
   U4014 : NAND2_X1 port map( A1 => n28738, A2 => n26892, ZN => n695);
   U4015 : BUF_X4 port map( I => n7198, Z => n25995);
   U4020 : NAND2_X1 port map( A1 => n30269, A2 => n26390, ZN => n28888);
   U4024 : NAND2_X1 port map( A1 => n11254, A2 => n11253, ZN => n17295);
   U4025 : NAND2_X1 port map( A1 => n26281, A2 => n31822, ZN => n14267);
   U4035 : NAND2_X1 port map( A1 => n25760, A2 => n24729, ZN => n12265);
   U4036 : INV_X1 port map( I => n28223, ZN => n24734);
   U4044 : CLKBUF_X1 port map( I => n15528, Z => n28634);
   U4066 : NOR2_X1 port map( A1 => n32017, A2 => n27982, ZN => n9398);
   U4070 : INV_X1 port map( I => n7511, ZN => n27791);
   U4072 : NAND2_X1 port map( A1 => n17069, A2 => n794, ZN => n27267);
   U4078 : NOR2_X1 port map( A1 => n7019, A2 => n1086, ZN => n7018);
   U4093 : NAND2_X1 port map( A1 => n31772, A2 => n27591, ZN => n6767);
   U4104 : NOR2_X1 port map( A1 => n6286, A2 => n1931, ZN => n27854);
   U4105 : CLKBUF_X2 port map( I => n24308, Z => n28590);
   U4119 : CLKBUF_X2 port map( I => n4821, Z => n27436);
   U4123 : CLKBUF_X2 port map( I => n24110, Z => n29010);
   U4128 : NAND2_X1 port map( A1 => n28509, A2 => n28507, ZN => n10383);
   U4129 : NAND2_X1 port map( A1 => n17086, A2 => n23766, ZN => n14587);
   U4134 : NAND2_X1 port map( A1 => n27078, A2 => n1253, ZN => n57);
   U4163 : NAND2_X1 port map( A1 => n23116, A2 => n23115, ZN => n26150);
   U4168 : CLKBUF_X2 port map( I => n23157, Z => n29068);
   U4174 : INV_X1 port map( I => n8674, ZN => n27321);
   U4187 : NAND2_X1 port map( A1 => n23917, A2 => n6869, ZN => n26533);
   U4331 : INV_X1 port map( I => n23458, ZN => n29220);
   U4335 : INV_X1 port map( I => n23494, ZN => n26924);
   U4342 : INV_X1 port map( I => n33265, ZN => n28492);
   U4348 : INV_X1 port map( I => n28402, ZN => n28401);
   U4349 : NOR2_X1 port map( A1 => n26026, A2 => n28227, ZN => n28862);
   U4353 : NAND2_X1 port map( A1 => n2028, A2 => n2029, ZN => n26336);
   U4362 : NAND2_X1 port map( A1 => n27191, A2 => n29176, ZN => n22054);
   U4365 : INV_X1 port map( I => n11084, ZN => n2031);
   U4379 : OAI21_X1 port map( A1 => n28778, A2 => n28777, B => n23055, ZN => 
                           n17458);
   U4381 : OAI21_X1 port map( A1 => n26106, A2 => n29174, B => n29173, ZN => 
                           n27191);
   U4383 : NAND2_X1 port map( A1 => n22051, A2 => n31824, ZN => n29176);
   U4391 : NAND2_X1 port map( A1 => n23029, A2 => n23028, ZN => n27079);
   U4392 : INV_X1 port map( I => n17707, ZN => n27969);
   U4397 : CLKBUF_X2 port map( I => n15633, Z => n28891);
   U4418 : OR2_X1 port map( A1 => n1271, A2 => n10528, Z => n26104);
   U4423 : AND2_X1 port map( A1 => n22780, A2 => n30925, Z => n26106);
   U4455 : CLKBUF_X2 port map( I => n3670, Z => n26169);
   U4466 : CLKBUF_X2 port map( I => n12700, Z => n27389);
   U4475 : CLKBUF_X8 port map( I => n15829, Z => n27752);
   U4481 : CLKBUF_X2 port map( I => n8040, Z => n26868);
   U4531 : CLKBUF_X2 port map( I => n14307, Z => n28635);
   U4570 : INV_X1 port map( I => n22217, ZN => n26845);
   U4590 : CLKBUF_X2 port map( I => n22172, Z => n28490);
   U4597 : INV_X1 port map( I => n22149, ZN => n28465);
   U4604 : AND2_X1 port map( A1 => n21597, A2 => n21596, Z => n27120);
   U4608 : NAND2_X1 port map( A1 => n26265, A2 => n26625, ZN => n13539);
   U4631 : NAND2_X1 port map( A1 => n26522, A2 => n27005, ZN => n7240);
   U4634 : NAND2_X1 port map( A1 => n3807, A2 => n15837, ZN => n15836);
   U4635 : NOR2_X1 port map( A1 => n26386, A2 => n13490, ZN => n14871);
   U4662 : OAI21_X1 port map( A1 => n21682, A2 => n2575, B => n26341, ZN => 
                           n21517);
   U4673 : NOR2_X1 port map( A1 => n21682, A2 => n2575, ZN => n3742);
   U4680 : NAND2_X1 port map( A1 => n21509, A2 => n21510, ZN => n26451);
   U4682 : NOR2_X1 port map( A1 => n16327, A2 => n12866, ZN => n17429);
   U4691 : CLKBUF_X2 port map( I => n21462, Z => n28838);
   U4707 : NAND2_X1 port map( A1 => n27720, A2 => n13313, ZN => n13310);
   U4708 : NAND2_X1 port map( A1 => n21255, A2 => n21259, ZN => n28255);
   U4710 : NAND2_X1 port map( A1 => n21255, A2 => n21257, ZN => n21256);
   U4711 : INV_X1 port map( I => n27198, ZN => n21292);
   U4718 : NAND2_X1 port map( A1 => n20935, A2 => n20938, ZN => n28298);
   U4724 : NAND2_X1 port map( A1 => n28501, A2 => n32357, ZN => n16934);
   U4725 : NOR2_X1 port map( A1 => n21325, A2 => n1146, ZN => n8012);
   U4739 : OR2_X1 port map( A1 => n10546, A2 => n16034, Z => n11700);
   U4742 : NAND2_X1 port map( A1 => n17455, A2 => n21295, ZN => n27305);
   U4763 : CLKBUF_X2 port map( I => n15226, Z => n26407);
   U4771 : NOR2_X1 port map( A1 => n7822, A2 => n510, ZN => n9879);
   U4778 : CLKBUF_X2 port map( I => n14029, Z => n26798);
   U4788 : CLKBUF_X2 port map( I => n6854, Z => n27193);
   U4796 : CLKBUF_X4 port map( I => n20946, Z => n29062);
   U4799 : INV_X1 port map( I => n8972, ZN => n27200);
   U4800 : INV_X1 port map( I => n10508, ZN => n20823);
   U4806 : NAND2_X1 port map( A1 => n20272, A2 => n17658, ZN => n27923);
   U4807 : CLKBUF_X2 port map( I => n20953, Z => n28823);
   U4831 : NAND2_X1 port map( A1 => n442, A2 => n1863, ZN => n26296);
   U4845 : INV_X1 port map( I => n20601, ZN => n27621);
   U4848 : NAND2_X1 port map( A1 => n1160, A2 => n10431, ZN => n27620);
   U4857 : NAND2_X1 port map( A1 => n20383, A2 => n15162, ZN => n26986);
   U4861 : NAND2_X1 port map( A1 => n20419, A2 => n14054, ZN => n19893);
   U4869 : NOR2_X1 port map( A1 => n27105, A2 => n5748, ZN => n443);
   U4871 : OR2_X1 port map( A1 => n710, A2 => n28261, Z => n12149);
   U4911 : NOR2_X1 port map( A1 => n27301, A2 => n19842, ZN => n27300);
   U4915 : NAND2_X1 port map( A1 => n26825, A2 => n26823, ZN => n28454);
   U4916 : OAI21_X1 port map( A1 => n12682, A2 => n20136, B => n28012, ZN => 
                           n19837);
   U4918 : NAND2_X1 port map( A1 => n3486, A2 => n27398, ZN => n7473);
   U4934 : NOR2_X1 port map( A1 => n31046, A2 => n16108, ZN => n27019);
   U4935 : NOR2_X1 port map( A1 => n29339, A2 => n1166, ZN => n20017);
   U4936 : NOR2_X1 port map( A1 => n6859, A2 => n17882, ZN => n27301);
   U4943 : AND2_X1 port map( A1 => n13488, A2 => n821, Z => n26093);
   U4965 : INV_X2 port map( I => n11969, ZN => n25997);
   U4973 : NAND2_X1 port map( A1 => n29135, A2 => n29134, ZN => n29133);
   U4987 : AOI21_X1 port map( A1 => n12649, A2 => n16669, B => n26043, ZN => 
                           n50);
   U4990 : INV_X1 port map( I => n10398, ZN => n29135);
   U4991 : NAND2_X1 port map( A1 => n28498, A2 => n18297, ZN => n18298);
   U4994 : NAND2_X1 port map( A1 => n14611, A2 => n12549, ZN => n28371);
   U4997 : NOR2_X1 port map( A1 => n19214, A2 => n29963, ZN => n28133);
   U5000 : NAND2_X1 port map( A1 => n19092, A2 => n19093, ZN => n27929);
   U5006 : INV_X2 port map( I => n2207, ZN => n5491);
   U5011 : OAI21_X1 port map( A1 => n13444, A2 => n958, B => n16207, ZN => 
                           n27857);
   U5016 : NAND2_X1 port map( A1 => n18851, A2 => n18730, ZN => n27762);
   U5030 : NAND2_X1 port map( A1 => n18850, A2 => n18849, ZN => n27761);
   U5033 : NAND2_X1 port map( A1 => n18662, A2 => n17477, ZN => n29239);
   U5034 : INV_X1 port map( I => n18858, ZN => n28102);
   U5041 : CLKBUF_X2 port map( I => n954, Z => n28707);
   U5047 : INV_X1 port map( I => n16691, ZN => n28422);
   U5050 : CLKBUF_X2 port map( I => n488, Z => n26810);
   U5053 : CLKBUF_X2 port map( I => n270, Z => n27940);
   U5056 : CLKBUF_X2 port map( I => n18811, Z => n28686);
   U5059 : INV_X1 port map( I => n25728, ZN => n28711);
   U5060 : CLKBUF_X2 port map( I => n10114, Z => n28344);
   U5061 : INV_X1 port map( I => n16527, ZN => n28462);
   U5063 : INV_X1 port map( I => n25282, ZN => n27672);
   U5068 : INV_X1 port map( I => n25079, ZN => n26001);
   U5069 : NAND2_X1 port map( A1 => n18662, A2 => n17478, ZN => n11406);
   U5092 : CLKBUF_X1 port map( I => n8386, Z => n28578);
   U5104 : AOI21_X1 port map( A1 => n15956, A2 => n18487, B => n9, ZN => n18488
                           );
   U5105 : NOR2_X1 port map( A1 => n18635, A2 => n18743, ZN => n16359);
   U5123 : AOI21_X1 port map( A1 => n10669, A2 => n18679, B => n10537, ZN => 
                           n10829);
   U5130 : NOR2_X1 port map( A1 => n4868, A2 => n5327, ZN => n5644);
   U5135 : NOR2_X1 port map( A1 => n18648, A2 => n18650, ZN => n2430);
   U5157 : NAND2_X1 port map( A1 => n2614, A2 => n16474, ZN => n26594);
   U5172 : NAND2_X1 port map( A1 => n31821, A2 => n18722, ZN => n18724);
   U5178 : AOI22_X1 port map( A1 => n16181, A2 => n28010, B1 => n29659, B2 => 
                           n13360, ZN => n13444);
   U5202 : INV_X1 port map( I => n5032, ZN => n3341);
   U5203 : NAND3_X1 port map( A1 => n7714, A2 => n9766, A3 => n7713, ZN => 
                           n12826);
   U5222 : NOR2_X1 port map( A1 => n745, A2 => n19021, ZN => n6059);
   U5223 : NOR2_X1 port map( A1 => n6846, A2 => n7995, ZN => n28929);
   U5235 : AND3_X1 port map( A1 => n27743, A2 => n13925, A3 => n949, Z => 
                           n26043);
   U5256 : NAND2_X1 port map( A1 => n14354, A2 => n13475, ZN => n274);
   U5283 : CLKBUF_X1 port map( I => n4632, Z => n294);
   U5316 : NOR2_X1 port map( A1 => n3790, A2 => n27805, ZN => n28419);
   U5327 : CLKBUF_X2 port map( I => n567, Z => n28423);
   U5339 : AND3_X1 port map( A1 => n16108, A2 => n1161, A3 => n13605, Z => 
                           n6073);
   U5340 : NAND2_X1 port map( A1 => n19456, A2 => n16681, ZN => n19846);
   U5374 : NOR2_X1 port map( A1 => n10613, A2 => n28904, ZN => n28269);
   U5405 : NAND2_X1 port map( A1 => n19906, A2 => n17790, ZN => n15256);
   U5412 : NOR2_X1 port map( A1 => n8031, A2 => n7577, ZN => n3750);
   U5423 : NAND2_X1 port map( A1 => n20564, A2 => n12263, ZN => n20568);
   U5435 : NOR2_X1 port map( A1 => n20418, A2 => n20417, ZN => n20422);
   U5444 : INV_X1 port map( I => n20917, ZN => n20809);
   U5447 : INV_X1 port map( I => n5724, ZN => n10109);
   U5486 : NOR2_X1 port map( A1 => n8190, A2 => n21095, ZN => n17841);
   U5504 : NOR2_X1 port map( A1 => n26677, A2 => n26635, ZN => n7225);
   U5513 : NAND2_X1 port map( A1 => n17832, A2 => n21317, ZN => n20373);
   U5521 : NAND2_X1 port map( A1 => n4683, A2 => n27684, ZN => n28549);
   U5537 : NAND2_X1 port map( A1 => n21752, A2 => n15414, ZN => n15412);
   U5538 : AOI21_X1 port map( A1 => n9699, A2 => n28037, B => n8197, ZN => 
                           n15905);
   U5546 : NAND3_X1 port map( A1 => n28737, A2 => n18218, A3 => n1019, ZN => 
                           n10555);
   U5563 : NAND2_X1 port map( A1 => n26993, A2 => n12643, ZN => n12641);
   U5569 : NAND2_X1 port map( A1 => n16544, A2 => n16543, ZN => n14950);
   U5587 : AND2_X1 port map( A1 => n32506, A2 => n21568, Z => n3315);
   U5588 : INV_X1 port map( I => n22291, ZN => n1903);
   U5595 : NOR2_X1 port map( A1 => n21736, A2 => n21867, ZN => n26298);
   U5600 : OAI22_X1 port map( A1 => n11848, A2 => n14917, B1 => n21346, B2 => 
                           n8140, ZN => n21347);
   U5605 : NAND3_X1 port map( A1 => n15127, A2 => n31954, A3 => n21741, ZN => 
                           n14041);
   U5607 : INV_X1 port map( I => n22005, ZN => n22086);
   U5614 : INV_X1 port map( I => n21937, ZN => n28941);
   U5623 : NAND2_X1 port map( A1 => n22484, A2 => n6297, ZN => n8594);
   U5637 : NOR2_X1 port map( A1 => n6297, A2 => n22641, ZN => n4300);
   U5674 : NAND3_X1 port map( A1 => n11250, A2 => n16334, A3 => n27959, ZN => 
                           n14069);
   U5681 : NOR2_X1 port map( A1 => n22664, A2 => n27415, ZN => n22437);
   U5684 : NOR2_X1 port map( A1 => n898, A2 => n32595, ZN => n10645);
   U5690 : NAND2_X1 port map( A1 => n7819, A2 => n28131, ZN => n135);
   U5706 : INV_X1 port map( I => n23051, ZN => n28555);
   U5710 : INV_X1 port map( I => n30234, ZN => n1267);
   U5719 : NAND2_X1 port map( A1 => n2937, A2 => n8308, ZN => n26590);
   U5725 : AOI21_X1 port map( A1 => n17707, A2 => n23026, B => n6190, ZN => 
                           n6189);
   U5743 : INV_X2 port map( I => n13694, ZN => n23158);
   U5748 : INV_X1 port map( I => n23196, ZN => n23216);
   U5757 : INV_X1 port map( I => n11897, ZN => n10218);
   U5761 : INV_X1 port map( I => n528, ZN => n26888);
   U5763 : INV_X1 port map( I => n23447, ZN => n27080);
   U5773 : INV_X1 port map( I => n29178, ZN => n15971);
   U5797 : NAND2_X1 port map( A1 => n23855, A2 => n29178, ZN => n9167);
   U5808 : INV_X1 port map( I => n9490, ZN => n10967);
   U5810 : INV_X1 port map( I => n23851, ZN => n8615);
   U5816 : NOR2_X1 port map( A1 => n27455, A2 => n1099, ZN => n14119);
   U5825 : INV_X1 port map( I => n14350, ZN => n300);
   U5837 : NOR2_X1 port map( A1 => n23940, A2 => n31807, ZN => n2563);
   U5845 : AND2_X1 port map( A1 => n6394, A2 => n30282, Z => n15017);
   U5846 : INV_X1 port map( I => n14193, ZN => n23544);
   U5866 : NAND2_X1 port map( A1 => n13260, A2 => n24004, ZN => n2865);
   U5885 : NOR3_X1 port map( A1 => n15011, A2 => n24084, A3 => n14913, ZN => 
                           n24035);
   U5896 : NOR2_X1 port map( A1 => n24288, A2 => n9625, ZN => n24108);
   U5898 : OAI21_X1 port map( A1 => n12402, A2 => n24140, B => n24087, ZN => 
                           n29184);
   U5920 : INV_X1 port map( I => n25115, ZN => n27650);
   U5946 : OR2_X1 port map( A1 => n10170, A2 => n27181, Z => n15459);
   U5958 : NOR2_X1 port map( A1 => n9198, A2 => n28096, ZN => n7806);
   U5963 : NOR2_X1 port map( A1 => n25900, A2 => n18219, ZN => n6325);
   U5975 : NAND2_X1 port map( A1 => n33919, A2 => n33915, ZN => n28562);
   U6014 : NOR2_X1 port map( A1 => n9611, A2 => n25234, ZN => n9610);
   U6038 : NOR2_X1 port map( A1 => n25390, A2 => n24867, ZN => n24672);
   U6052 : NAND2_X1 port map( A1 => n25316, A2 => n2236, ZN => n17028);
   U6054 : CLKBUF_X1 port map( I => n24909, Z => n14075);
   U6087 : INV_X1 port map( I => n25206, ZN => n27920);
   U6088 : NAND2_X1 port map( A1 => n25362, A2 => n25361, ZN => n28517);
   U6091 : AOI21_X1 port map( A1 => n7701, A2 => n25916, B => n5411, ZN => 
                           n11155);
   U6096 : INV_X1 port map( I => n25064, ZN => n16911);
   U6103 : XNOR2_X1 port map( A1 => n19518, A2 => n2980, ZN => n26004);
   U6105 : XNOR2_X1 port map( A1 => n19599, A2 => n25355, ZN => n26005);
   U6107 : OR2_X1 port map( A1 => n31721, A2 => n9831, Z => n26008);
   U6120 : AND2_X1 port map( A1 => n9329, A2 => n6129, Z => n26012);
   U6123 : AND2_X1 port map( A1 => n21400, A2 => n21398, Z => n26013);
   U6125 : AND2_X1 port map( A1 => n924, A2 => n1337, Z => n26014);
   U6127 : XNOR2_X1 port map( A1 => n16349, A2 => n702, ZN => n26016);
   U6135 : OR3_X1 port map( A1 => n11306, A2 => n11090, A3 => n25633, Z => 
                           n26022);
   U6138 : AND2_X1 port map( A1 => n11366, A2 => n25412, Z => n26023);
   U6143 : XNOR2_X1 port map( A1 => n6906, A2 => n25751, ZN => n26028);
   U6144 : XOR2_X1 port map( A1 => n33835, A2 => n23191, Z => n26029);
   U6145 : XNOR2_X1 port map( A1 => n20692, A2 => n16523, ZN => n26030);
   U6148 : XNOR2_X1 port map( A1 => n34016, A2 => n16506, ZN => n26031);
   U6154 : XNOR2_X1 port map( A1 => n19773, A2 => n24937, ZN => n26032);
   U6155 : AND2_X1 port map( A1 => n1672, A2 => n1671, Z => n26033);
   U6158 : INV_X1 port map( I => n8376, ZN => n18791);
   U6162 : AND2_X1 port map( A1 => n23754, A2 => n22617, Z => n26036);
   U6169 : AND2_X1 port map( A1 => n28958, A2 => n15528, Z => n26038);
   U6173 : CLKBUF_X2 port map( I => n5748, Z => n26730);
   U6182 : OR2_X1 port map( A1 => n20413, A2 => n20414, Z => n26041);
   U6186 : XNOR2_X1 port map( A1 => n356, A2 => n24573, ZN => n26045);
   U6192 : INV_X1 port map( I => n18557, ZN => n18775);
   U6211 : XOR2_X1 port map( A1 => n33835, A2 => n25908, Z => n26053);
   U6212 : XOR2_X1 port map( A1 => n12376, A2 => n24738, Z => n26054);
   U6214 : XNOR2_X1 port map( A1 => n19712, A2 => n24943, ZN => n26055);
   U6215 : XNOR2_X1 port map( A1 => n22226, A2 => n16691, ZN => n26057);
   U6221 : XNOR2_X1 port map( A1 => n20861, A2 => n16479, ZN => n26058);
   U6222 : XNOR2_X1 port map( A1 => n23476, A2 => n25167, ZN => n26059);
   U6225 : NAND2_X1 port map( A1 => n23842, A2 => n23887, ZN => n26060);
   U6226 : AND2_X1 port map( A1 => n25278, A2 => n16291, Z => n26061);
   U6232 : AND2_X1 port map( A1 => n16170, A2 => n16306, Z => n26065);
   U6234 : AND2_X1 port map( A1 => n12500, A2 => n13925, Z => n26067);
   U6235 : NAND2_X1 port map( A1 => n31915, A2 => n976, ZN => n26069);
   U6239 : OR2_X1 port map( A1 => n10724, A2 => n16166, Z => n26072);
   U6245 : XNOR2_X1 port map( A1 => n7653, A2 => n20820, ZN => n26075);
   U6250 : XNOR2_X1 port map( A1 => n27156, A2 => n25735, ZN => n26076);
   U6259 : AND3_X1 port map( A1 => n791, A2 => n9964, A3 => n24220, Z => n26079
                           );
   U6262 : CLKBUF_X4 port map( I => n1484, Z => n28227);
   U6267 : INV_X1 port map( I => n1484, ZN => n26160);
   U6279 : NOR2_X1 port map( A1 => n11051, A2 => n13080, ZN => n26083);
   U6284 : XNOR2_X1 port map( A1 => n12957, A2 => n9874, ZN => n26085);
   U6293 : XNOR2_X1 port map( A1 => n20732, A2 => n20731, ZN => n26087);
   U6294 : AND2_X2 port map( A1 => n19938, A2 => n16105, Z => n26088);
   U6311 : XNOR2_X1 port map( A1 => n17385, A2 => n25436, ZN => n26094);
   U6316 : XNOR2_X1 port map( A1 => n21994, A2 => n24623, ZN => n26096);
   U6323 : XNOR2_X1 port map( A1 => n22031, A2 => n25610, ZN => n26097);
   U6333 : XNOR2_X1 port map( A1 => n22130, A2 => n16472, ZN => n26100);
   U6337 : XNOR2_X1 port map( A1 => n4732, A2 => n25929, ZN => n26101);
   U6341 : XNOR2_X1 port map( A1 => n7477, A2 => n16423, ZN => n26103);
   U6347 : XNOR2_X1 port map( A1 => n7229, A2 => n12754, ZN => n26108);
   U6355 : INV_X1 port map( I => n11983, ZN => n29175);
   U6359 : XNOR2_X1 port map( A1 => n24629, A2 => n24628, ZN => n26111);
   U6369 : AND2_X2 port map( A1 => n31957, A2 => n4646, Z => n26113);
   U6372 : XNOR2_X1 port map( A1 => n227, A2 => n6924, ZN => n26115);
   U6374 : XNOR2_X1 port map( A1 => n16162, A2 => n23364, ZN => n26116);
   U6382 : XNOR2_X1 port map( A1 => n23467, A2 => n14526, ZN => n26118);
   U6385 : INV_X1 port map( I => n13308, ZN => n23559);
   U6389 : INV_X1 port map( I => n24327, ZN => n1093);
   U6390 : XOR2_X1 port map( A1 => n14645, A2 => n25693, Z => n26121);
   U6394 : XNOR2_X1 port map( A1 => n33971, A2 => n25450, ZN => n26123);
   U6397 : XNOR2_X1 port map( A1 => n32623, A2 => n13858, ZN => n26124);
   U6403 : OR2_X1 port map( A1 => n25659, A2 => n25657, Z => n26127);
   U6418 : XNOR2_X1 port map( A1 => n8269, A2 => n7808, ZN => n3393);
   U6421 : INV_X2 port map( I => n31451, ZN => n19107);
   U6422 : NAND2_X1 port map( A1 => n19063, A2 => n31451, ZN => n19062);
   U6448 : AND2_X1 port map( A1 => n32855, A2 => n10948, Z => n25611);
   U6463 : XOR2_X1 port map( A1 => n4397, A2 => n9505, Z => n4395);
   U6467 : XOR2_X1 port map( A1 => n22147, A2 => n28465, Z => n6396);
   U6475 : NAND2_X2 port map( A1 => n18032, A2 => n21279, ZN => n22147);
   U6488 : NAND2_X1 port map( A1 => n31654, A2 => n21777, ZN => n4211);
   U6489 : XOR2_X1 port map( A1 => n12422, A2 => n12032, Z => n13084);
   U6508 : NOR2_X2 port map( A1 => n29027, A2 => n29026, ZN => n987);
   U6542 : XOR2_X1 port map( A1 => n20779, A2 => n11374, Z => n26140);
   U6559 : AOI21_X1 port map( A1 => n24283, A2 => n16356, B => n4151, ZN => 
                           n3862);
   U6575 : XOR2_X1 port map( A1 => n10289, A2 => n23498, Z => n26145);
   U6576 : NOR2_X2 port map( A1 => n12358, A2 => n24466, ZN => n26334);
   U6607 : NAND2_X2 port map( A1 => n26150, A2 => n26073, ZN => n839);
   U6624 : INV_X2 port map( I => n26153, ZN => n19942);
   U6626 : XOR2_X1 port map( A1 => n9821, A2 => n9818, Z => n26153);
   U6630 : XOR2_X1 port map( A1 => n16035, A2 => n26154, Z => n16682);
   U6632 : XOR2_X1 port map( A1 => n21918, A2 => n21919, Z => n26154);
   U6645 : XOR2_X1 port map( A1 => n24394, A2 => n9907, Z => n24395);
   U6662 : NOR2_X2 port map( A1 => n11608, A2 => n12691, ZN => n12313);
   U6666 : INV_X2 port map( I => n15393, ZN => n27748);
   U6669 : XOR2_X1 port map( A1 => n11092, A2 => n11093, Z => n15393);
   U6676 : AOI21_X2 port map( A1 => n4926, A2 => n5700, B => n26156, ZN => 
                           n4508);
   U6759 : INV_X2 port map( I => n26162, ZN => n13989);
   U6773 : NAND2_X2 port map( A1 => n17960, A2 => n16375, ZN => n22505);
   U6774 : INV_X2 port map( I => n15053, ZN => n26633);
   U6802 : NAND2_X2 port map( A1 => n2902, A2 => n2692, ZN => n19212);
   U6803 : NAND2_X2 port map( A1 => n18309, A2 => n18308, ZN => n2692);
   U6809 : NAND3_X1 port map( A1 => n17373, A2 => n26775, A3 => n23945, ZN => 
                           n23677);
   U6821 : NAND2_X2 port map( A1 => n2771, A2 => n26165, ZN => n20926);
   U6824 : XOR2_X1 port map( A1 => n9790, A2 => n26168, Z => n11100);
   U6827 : XOR2_X1 port map( A1 => n22241, A2 => n12898, Z => n26168);
   U6829 : XOR2_X1 port map( A1 => n24512, A2 => n31866, Z => n26502);
   U6836 : INV_X2 port map( I => n26170, ZN => n5736);
   U6842 : NAND2_X2 port map( A1 => n9806, A2 => n9804, ZN => n25654);
   U6868 : XOR2_X1 port map( A1 => n9761, A2 => n26172, Z => n7657);
   U6870 : XOR2_X1 port map( A1 => n21034, A2 => n11424, Z => n26172);
   U6873 : XOR2_X1 port map( A1 => n23343, A2 => n27041, Z => n5314);
   U6917 : OAI21_X2 port map( A1 => n27802, A2 => n822, B => n16059, ZN => 
                           n3962);
   U6926 : XNOR2_X1 port map( A1 => n33699, A2 => n13519, ZN => n29108);
   U6957 : OR2_X1 port map( A1 => n20158, A2 => n26182, Z => n10615);
   U6958 : XOR2_X1 port map( A1 => n20893, A2 => n20890, Z => n1686);
   U6959 : XOR2_X1 port map( A1 => n20982, A2 => n20822, Z => n20893);
   U6960 : XOR2_X1 port map( A1 => n1944, A2 => n9880, Z => n11062);
   U7021 : NAND2_X1 port map( A1 => n6102, A2 => n23052, ZN => n6101);
   U7050 : INV_X2 port map( I => n24158, ZN => n9934);
   U7054 : OAI21_X2 port map( A1 => n7377, A2 => n7378, B => n16629, ZN => 
                           n7376);
   U7066 : XOR2_X1 port map( A1 => n5241, A2 => n5240, Z => n26194);
   U7076 : NAND2_X1 port map( A1 => n26198, A2 => n24955, ZN => n26197);
   U7077 : OR2_X1 port map( A1 => n24955, A2 => n24956, Z => n26199);
   U7080 : OAI22_X1 port map( A1 => n8073, A2 => n1075, B1 => n7554, B2 => 
                           n28736, ZN => n14764);
   U7090 : NAND2_X1 port map( A1 => n24244, A2 => n28374, ZN => n24075);
   U7095 : NOR2_X2 port map( A1 => n24330, A2 => n24331, ZN => n24244);
   U7102 : NAND2_X2 port map( A1 => n7447, A2 => n26202, ZN => n14864);
   U7105 : XOR2_X1 port map( A1 => n22203, A2 => n14787, Z => n14786);
   U7109 : XOR2_X1 port map( A1 => n32084, A2 => n22031, Z => n22203);
   U7123 : NAND3_X2 port map( A1 => n26204, A2 => n9147, A3 => n23981, ZN => 
                           n9145);
   U7141 : NOR2_X1 port map( A1 => n15070, A2 => n180, ZN => n28773);
   U7159 : OR2_X2 port map( A1 => n7918, A2 => n10390, Z => n1783);
   U7170 : XOR2_X1 port map( A1 => n7574, A2 => n26208, Z => n681);
   U7171 : INV_X1 port map( I => n25880, ZN => n26208);
   U7182 : XOR2_X1 port map( A1 => n12473, A2 => n17194, Z => n663);
   U7197 : XOR2_X1 port map( A1 => n3619, A2 => n3618, Z => n16961);
   U7217 : XOR2_X1 port map( A1 => n26215, A2 => n19388, Z => n15476);
   U7219 : XOR2_X1 port map( A1 => n19387, A2 => n19567, Z => n26215);
   U7220 : XOR2_X1 port map( A1 => n24654, A2 => n24683, Z => n16930);
   U7274 : NAND2_X1 port map( A1 => n16954, A2 => n15296, ZN => n28);
   U7303 : XOR2_X1 port map( A1 => n23457, A2 => n23404, Z => n23314);
   U7309 : NAND2_X2 port map( A1 => n14610, A2 => n22738, ZN => n23457);
   U7320 : AOI22_X2 port map( A1 => n26228, A2 => n20877, B1 => n21691, B2 => 
                           n5628, ZN => n22056);
   U7323 : NAND3_X2 port map( A1 => n31927, A2 => n21, A3 => n13115, ZN => 
                           n26228);
   U7349 : XOR2_X1 port map( A1 => n5856, A2 => n26233, Z => n11068);
   U7350 : XOR2_X1 port map( A1 => n4975, A2 => n3870, Z => n26233);
   U7395 : XOR2_X1 port map( A1 => n5563, A2 => n5562, Z => n26237);
   U7399 : NOR2_X2 port map( A1 => n26239, A2 => n26238, ZN => n2285);
   U7400 : NOR2_X2 port map( A1 => n5825, A2 => n17882, ZN => n26239);
   U7405 : NAND2_X1 port map( A1 => n27934, A2 => n8125, ZN => n5079);
   U7409 : OAI21_X2 port map( A1 => n26241, A2 => n23946, B => n23950, ZN => 
                           n3554);
   U7422 : NOR2_X2 port map( A1 => n154, A2 => n1337, ZN => n21099);
   U7457 : OAI22_X2 port map( A1 => n1857, A2 => n28784, B1 => n13324, B2 => 
                           n17453, ZN => n13586);
   U7480 : XOR2_X1 port map( A1 => Plaintext(82), A2 => Key(82), Z => n26249);
   U7490 : AOI21_X2 port map( A1 => n18970, A2 => n12645, B => n26250, ZN => 
                           n19710);
   U7533 : NAND2_X1 port map( A1 => n20481, A2 => n26566, ZN => n8171);
   U7542 : XOR2_X1 port map( A1 => n21946, A2 => n6245, Z => n26256);
   U7559 : NAND2_X2 port map( A1 => n27741, A2 => n32594, ZN => n13867);
   U7610 : NAND2_X1 port map( A1 => n18150, A2 => n18151, ZN => n12230);
   U7625 : XOR2_X1 port map( A1 => n26262, A2 => n15987, Z => n8522);
   U7633 : XOR2_X1 port map( A1 => n15986, A2 => n24373, Z => n26262);
   U7714 : XOR2_X1 port map( A1 => n11527, A2 => n11525, Z => n18150);
   U7727 : NAND2_X2 port map( A1 => n6432, A2 => n3894, ZN => n28942);
   U7728 : NAND3_X2 port map( A1 => n7961, A2 => n27627, A3 => n17992, ZN => 
                           n7330);
   U7733 : AOI21_X2 port map( A1 => n26268, A2 => n21430, B => n7666, ZN => 
                           n21617);
   U7761 : XOR2_X1 port map( A1 => n15787, A2 => n6488, Z => n6033);
   U7770 : XOR2_X1 port map( A1 => n16792, A2 => n6028, Z => n26272);
   U7778 : NAND2_X1 port map( A1 => n29048, A2 => n29050, ZN => n26275);
   U7783 : XOR2_X1 port map( A1 => n26276, A2 => n7328, Z => n20939);
   U7784 : XOR2_X1 port map( A1 => n14522, A2 => n20687, Z => n26276);
   U7795 : XOR2_X1 port map( A1 => n16080, A2 => n14404, Z => n5699);
   U7800 : XOR2_X1 port map( A1 => n19626, A2 => n14293, Z => n14404);
   U7808 : AOI21_X2 port map( A1 => n17272, A2 => n21171, B => n27424, ZN => 
                           n27379);
   U7813 : NAND2_X2 port map( A1 => n10232, A2 => n10233, ZN => n22014);
   U7825 : INV_X4 port map( I => n26640, ZN => n11940);
   U7829 : XOR2_X1 port map( A1 => n28411, A2 => n27850, Z => n4529);
   U7839 : INV_X2 port map( I => n26284, ZN => n22429);
   U7854 : OR2_X1 port map( A1 => n8044, A2 => n15518, Z => n24605);
   U7865 : INV_X1 port map( I => n26439, ZN => n21669);
   U7878 : AOI21_X2 port map( A1 => n3128, A2 => n12178, B => n26006, ZN => 
                           n26291);
   U7884 : XOR2_X1 port map( A1 => n26294, A2 => n24089, Z => n24090);
   U7885 : XOR2_X1 port map( A1 => n28258, A2 => n25619, Z => n26294);
   U7886 : XOR2_X1 port map( A1 => n26295, A2 => n16038, Z => Ciphertext(93));
   U7902 : NAND3_X2 port map( A1 => n17420, A2 => n24214, A3 => n17676, ZN => 
                           n24474);
   U7906 : OR2_X1 port map( A1 => n28199, A2 => n16568, Z => n9233);
   U7908 : XOR2_X1 port map( A1 => n30319, A2 => n3589, Z => n4003);
   U7913 : NAND2_X1 port map( A1 => n31636, A2 => n29335, ZN => n22573);
   U7923 : XOR2_X1 port map( A1 => n26300, A2 => n2363, Z => n3511);
   U7939 : AND2_X1 port map( A1 => n27378, A2 => n7965, Z => n26301);
   U7942 : OAI22_X1 port map( A1 => n25667, A2 => n25666, B1 => n734, B2 => 
                           n25668, ZN => n28052);
   U7945 : NOR2_X1 port map( A1 => n11981, A2 => n7144, ZN => n15215);
   U7965 : NAND3_X2 port map( A1 => n26304, A2 => n27761, A3 => n27762, ZN => 
                           n19206);
   U7966 : NAND3_X1 port map( A1 => n6312, A2 => n6313, A3 => n957, ZN => 
                           n26304);
   U7976 : NOR2_X2 port map( A1 => n4856, A2 => n4857, ZN => n18266);
   U7983 : XOR2_X1 port map( A1 => n29030, A2 => n4157, Z => n19491);
   U7995 : BUF_X2 port map( I => n7024, Z => n26305);
   U8004 : AOI21_X2 port map( A1 => n11436, A2 => n11437, B => n26307, ZN => 
                           n11439);
   U8018 : XOR2_X1 port map( A1 => n23266, A2 => n30272, Z => n6608);
   U8061 : XOR2_X1 port map( A1 => n27290, A2 => n3476, Z => n14142);
   U8065 : XOR2_X1 port map( A1 => n21033, A2 => n9762, Z => n9761);
   U8075 : OAI21_X2 port map( A1 => n26318, A2 => n18573, B => n29087, ZN => 
                           n5478);
   U8079 : NAND2_X2 port map( A1 => n951, A2 => n4868, ZN => n12490);
   U8084 : NAND2_X2 port map( A1 => n3181, A2 => n6555, ZN => n24347);
   U8106 : NAND2_X2 port map( A1 => n9917, A2 => n8105, ZN => n24867);
   U8107 : NAND3_X2 port map( A1 => n26362, A2 => n12215, A3 => n24860, ZN => 
                           n24862);
   U8112 : NAND2_X2 port map( A1 => n24436, A2 => n25696, ZN => n25627);
   U8123 : NAND2_X2 port map( A1 => n4075, A2 => n10056, ZN => n11988);
   U8126 : OAI21_X2 port map( A1 => n25539, A2 => n25536, B => n17046, ZN => 
                           n25297);
   U8134 : XOR2_X1 port map( A1 => n6548, A2 => n16958, Z => n20767);
   U8160 : AND2_X1 port map( A1 => n15968, A2 => n20676, Z => n26328);
   U8185 : XOR2_X1 port map( A1 => n30628, A2 => n22014, Z => n22027);
   U8189 : INV_X2 port map( I => n26330, ZN => n522);
   U8191 : XOR2_X1 port map( A1 => n5796, A2 => n13452, Z => n26330);
   U8216 : INV_X2 port map( I => n26334, ZN => n13326);
   U8225 : AND2_X1 port map( A1 => n30978, A2 => n13114, Z => n4433);
   U8237 : XOR2_X1 port map( A1 => n26338, A2 => n10052, Z => n10051);
   U8242 : OR2_X1 port map( A1 => n20344, A2 => n10717, Z => n20538);
   U8243 : NOR2_X1 port map( A1 => n26445, A2 => n432, ZN => n3168);
   U8271 : INV_X2 port map( I => n26340, ZN => n11762);
   U8279 : NAND2_X2 port map( A1 => n30995, A2 => n19224, ZN => n19060);
   U8337 : OAI22_X2 port map( A1 => n26355, A2 => n33635, B1 => n32951, B2 => 
                           n19185, ZN => n11385);
   U8347 : NAND2_X2 port map( A1 => n2612, A2 => n7687, ZN => n13219);
   U8350 : AOI21_X2 port map( A1 => n26357, A2 => n19868, B => n941, ZN => 
                           n19871);
   U8360 : NOR2_X2 port map( A1 => n4633, A2 => n8757, ZN => n5111);
   U8362 : NOR2_X2 port map( A1 => n14556, A2 => n21053, ZN => n4633);
   U8380 : XOR2_X1 port map( A1 => n5436, A2 => n5434, Z => n4060);
   U8391 : INV_X2 port map( I => n20555, ZN => n28166);
   U8392 : OAI22_X2 port map( A1 => n19881, A2 => n19880, B1 => n31046, B2 => 
                           n11119, ZN => n20555);
   U8410 : XOR2_X1 port map( A1 => n24440, A2 => n24664, Z => n24596);
   U8411 : OAI21_X2 port map( A1 => n2921, A2 => n7101, B => n13046, ZN => 
                           n24440);
   U8421 : NAND2_X1 port map( A1 => n12217, A2 => n25689, ZN => n26362);
   U8428 : NAND2_X2 port map( A1 => n11795, A2 => n7457, ZN => n22013);
   U8436 : XOR2_X1 port map( A1 => n23282, A2 => n2520, Z => n23408);
   U8453 : XOR2_X1 port map( A1 => n26365, A2 => n8537, Z => n9163);
   U8458 : BUF_X2 port map( I => n20117, Z => n26368);
   U8460 : OAI22_X2 port map( A1 => n26909, A2 => n2430, B1 => n2432, B2 => 
                           n16120, ZN => n11203);
   U8516 : INV_X2 port map( I => n15839, ZN => n28714);
   U8519 : XOR2_X1 port map( A1 => n7032, A2 => n7029, Z => n15839);
   U8525 : NOR2_X2 port map( A1 => n23754, A2 => n1099, ZN => n12432);
   U8530 : XOR2_X1 port map( A1 => n32581, A2 => n31374, Z => n20779);
   U8543 : INV_X1 port map( I => n19188, ZN => n26376);
   U8554 : NOR2_X1 port map( A1 => n18802, A2 => n33621, ZN => n26378);
   U8574 : AOI21_X2 port map( A1 => n20349, A2 => n760, B => n27227, ZN => 
                           n28813);
   U8583 : NAND2_X1 port map( A1 => n28366, A2 => n5288, ZN => n1864);
   U8589 : XOR2_X1 port map( A1 => n8071, A2 => n26423, Z => n23130);
   U8616 : XOR2_X1 port map( A1 => n3411, A2 => n3410, Z => n26385);
   U8618 : XOR2_X1 port map( A1 => n24479, A2 => n12969, Z => n24778);
   U8619 : NAND2_X2 port map( A1 => n12403, A2 => n29184, ZN => n12969);
   U8625 : NOR2_X2 port map( A1 => n8984, A2 => n8983, ZN => n26387);
   U8638 : NAND2_X1 port map( A1 => n25144, A2 => n17595, ZN => n16729);
   U8647 : NOR2_X2 port map( A1 => n3698, A2 => n3695, ZN => n14396);
   U8654 : AOI21_X2 port map( A1 => n2176, A2 => n21172, B => n2174, ZN => 
                           n15172);
   U8676 : XOR2_X1 port map( A1 => n10482, A2 => n9673, Z => n26388);
   U8710 : NAND2_X2 port map( A1 => n727, A2 => n7592, ZN => n21712);
   U8711 : NOR2_X2 port map( A1 => n1456, A2 => n1457, ZN => n7592);
   U8722 : NAND2_X2 port map( A1 => n26393, A2 => n22629, ZN => n4734);
   U8801 : NOR2_X1 port map( A1 => n6433, A2 => n31531, ZN => n13835);
   U8875 : AOI22_X2 port map( A1 => n26400, A2 => n28815, B1 => n24462, B2 => 
                           n8648, ZN => n14931);
   U8894 : XOR2_X1 port map( A1 => n32537, A2 => n22148, Z => n5105);
   U8904 : NAND3_X2 port map( A1 => n21505, A2 => n21510, A3 => n21506, ZN => 
                           n21706);
   U8910 : NOR2_X2 port map( A1 => n26772, A2 => n26408, ZN => n17720);
   U8921 : INV_X1 port map( I => n15786, ZN => n27098);
   U8931 : INV_X1 port map( I => n26585, ZN => n20439);
   U8941 : INV_X2 port map( I => n12948, ZN => n3874);
   U8946 : NAND2_X1 port map( A1 => n26775, A2 => n12948, ZN => n23943);
   U8952 : XOR2_X1 port map( A1 => n6539, A2 => n12950, Z => n12948);
   U8956 : AND2_X1 port map( A1 => n16811, A2 => n20117, Z => n19959);
   U8964 : INV_X2 port map( I => n11774, ZN => n5805);
   U8978 : INV_X2 port map( I => n2022, ZN => n26415);
   U8992 : AOI21_X2 port map( A1 => n1563, A2 => n26373, B => n27451, ZN => 
                           n23387);
   U8997 : INV_X2 port map( I => n26418, ZN => n18373);
   U8999 : XNOR2_X1 port map( A1 => Key(41), A2 => Plaintext(41), ZN => n26418)
                           ;
   U9009 : XOR2_X1 port map( A1 => n32537, A2 => n21923, Z => n21577);
   U9020 : NOR2_X1 port map( A1 => n8742, A2 => n9885, ZN => n3022);
   U9051 : XOR2_X1 port map( A1 => n23128, A2 => n23127, Z => n26423);
   U9104 : XOR2_X1 port map( A1 => n15161, A2 => n27125, Z => n26429);
   U9105 : XOR2_X1 port map( A1 => n12413, A2 => n19748, Z => n4701);
   U9128 : XOR2_X1 port map( A1 => n1259, A2 => n15130, Z => n6706);
   U9137 : INV_X1 port map( I => n32917, ZN => n840);
   U9142 : NAND2_X2 port map( A1 => n990, A2 => n30297, ZN => n11626);
   U9145 : INV_X4 port map( I => n10528, ZN => n990);
   U9150 : INV_X2 port map( I => n26433, ZN => n22427);
   U9163 : INV_X2 port map( I => n12701, ZN => n22982);
   U9164 : OAI21_X2 port map( A1 => n4503, A2 => n4504, B => n4502, ZN => 
                           n12701);
   U9169 : NAND3_X2 port map( A1 => n6251, A2 => n6250, A3 => n26916, ZN => 
                           n27439);
   U9174 : XOR2_X1 port map( A1 => n26435, A2 => n17991, Z => n17407);
   U9192 : NOR2_X1 port map( A1 => n7867, A2 => n25941, ZN => n8264);
   U9197 : XOR2_X1 port map( A1 => n19505, A2 => n9138, Z => n26436);
   U9198 : XOR2_X1 port map( A1 => n11884, A2 => n6396, Z => n6395);
   U9203 : NOR2_X2 port map( A1 => n18941, A2 => n18942, ZN => n19509);
   U9209 : NAND2_X1 port map( A1 => n11390, A2 => n14926, ZN => n11398);
   U9210 : NAND2_X1 port map( A1 => n7941, A2 => n26440, ZN => n434);
   U9222 : XOR2_X1 port map( A1 => n8762, A2 => n25598, Z => n10697);
   U9245 : NAND2_X1 port map( A1 => n2105, A2 => n6891, ZN => n26444);
   U9250 : NAND2_X1 port map( A1 => n8373, A2 => n26774, ZN => n20029);
   U9292 : XOR2_X1 port map( A1 => n23370, A2 => n26452, Z => n15612);
   U9293 : XOR2_X1 port map( A1 => n32975, A2 => n6169, Z => n26452);
   U9294 : NAND2_X1 port map( A1 => n22665, A2 => n22576, ZN => n26453);
   U9298 : XOR2_X1 port map( A1 => n28460, A2 => n8548, Z => n3621);
   U9308 : NAND2_X2 port map( A1 => n14272, A2 => n14270, ZN => n27954);
   U9310 : NOR2_X1 port map( A1 => n26455, A2 => n27648, ZN => n26690);
   U9311 : OAI21_X1 port map( A1 => n27649, A2 => n230, B => n32441, ZN => 
                           n26455);
   U9319 : XOR2_X1 port map( A1 => n3285, A2 => n3283, Z => n26774);
   U9327 : NAND2_X2 port map( A1 => n2593, A2 => n2595, ZN => n26600);
   U9330 : XOR2_X1 port map( A1 => n19490, A2 => n3415, Z => n26456);
   U9340 : NOR2_X1 port map( A1 => n1360, A2 => n1043, ZN => n10273);
   U9343 : NAND2_X2 port map( A1 => n18598, A2 => n26458, ZN => n19330);
   U9353 : XNOR2_X1 port map( A1 => n20801, A2 => n25881, ZN => n29054);
   U9400 : XOR2_X1 port map( A1 => n24390, A2 => n24472, Z => n17653);
   U9418 : NAND2_X2 port map( A1 => n13831, A2 => n26469, ZN => n19074);
   U9434 : OAI21_X2 port map( A1 => n15870, A2 => n9476, B => n1389, ZN => 
                           n26627);
   U9457 : AOI21_X2 port map( A1 => n18809, A2 => n18650, B => n26472, ZN => 
                           n28944);
   U9459 : AND2_X1 port map( A1 => n18648, A2 => n18349, Z => n26472);
   U9460 : NOR2_X2 port map( A1 => n2614, A2 => n18648, ZN => n18809);
   U9494 : OR2_X1 port map( A1 => n20393, A2 => n15468, Z => n26478);
   U9501 : NAND2_X2 port map( A1 => n24334, A2 => n3014, ZN => n28202);
   U9502 : NOR2_X2 port map( A1 => n1876, A2 => n1875, ZN => n24334);
   U9516 : XOR2_X1 port map( A1 => n20755, A2 => n26530, Z => n13857);
   U9521 : INV_X1 port map( I => n8121, ZN => n27768);
   U9522 : INV_X4 port map( I => n13412, ZN => n791);
   U9547 : XOR2_X1 port map( A1 => n8109, A2 => n24525, Z => n8113);
   U9562 : XOR2_X1 port map( A1 => n26484, A2 => n22247, Z => n8471);
   U9576 : XOR2_X1 port map( A1 => n13602, A2 => n27147, Z => n13727);
   U9578 : NAND2_X2 port map( A1 => n26485, A2 => n11037, ZN => n20849);
   U9592 : XOR2_X1 port map( A1 => n14682, A2 => n12671, Z => n20796);
   U9595 : AND2_X1 port map( A1 => n691, A2 => n8168, Z => n12508);
   U9604 : XOR2_X1 port map( A1 => n15726, A2 => n15725, Z => n26487);
   U9611 : XOR2_X1 port map( A1 => n5976, A2 => n29170, Z => n5975);
   U9630 : XOR2_X1 port map( A1 => n26490, A2 => n7652, Z => n446);
   U9634 : XOR2_X1 port map( A1 => n9665, A2 => n4314, Z => n26490);
   U9639 : XOR2_X1 port map( A1 => n26492, A2 => n21988, Z => n29259);
   U9641 : XOR2_X1 port map( A1 => n3723, A2 => n26493, Z => n26492);
   U9730 : AOI22_X2 port map( A1 => n16549, A2 => n22534, B1 => n12698, B2 => 
                           n17146, ZN => n12697);
   U9731 : OR2_X1 port map( A1 => n22655, A2 => n22951, Z => n22862);
   U9733 : XOR2_X1 port map( A1 => n26502, A2 => n7173, Z => n29275);
   U9748 : NAND2_X2 port map( A1 => n26505, A2 => n26504, ZN => n16194);
   U9810 : BUF_X2 port map( I => n20137, Z => n8558);
   U9828 : XOR2_X1 port map( A1 => n26511, A2 => n11542, Z => n8625);
   U9847 : INV_X2 port map( I => n26515, ZN => n16333);
   U9859 : BUF_X2 port map( I => n12356, Z => n26516);
   U9861 : AOI22_X2 port map( A1 => n27696, A2 => n14734, B1 => n29223, B2 => 
                           n19203, ZN => n8692);
   U9862 : XOR2_X1 port map( A1 => n22295, A2 => n18189, Z => n21944);
   U9886 : NAND2_X2 port map( A1 => n26520, A2 => n16915, ZN => n14831);
   U9896 : NAND2_X2 port map( A1 => n25033, A2 => n26521, ZN => n25044);
   U9902 : OAI21_X1 port map( A1 => n25031, A2 => n14055, B => n29334, ZN => 
                           n26521);
   U9922 : NAND2_X2 port map( A1 => n26524, A2 => n9453, ZN => n13652);
   U9936 : INV_X2 port map( I => n26525, ZN => n11513);
   U9940 : XNOR2_X1 port map( A1 => n11514, A2 => n26977, ZN => n26525);
   U9965 : NAND2_X2 port map( A1 => n12515, A2 => n31470, ZN => n20385);
   U9968 : AOI22_X2 port map( A1 => n3571, A2 => n3401, B1 => n32004, B2 => 
                           n23577, ZN => n24201);
   U10063 : NAND2_X2 port map( A1 => n6332, A2 => n18810, ZN => n2207);
   U10077 : XOR2_X1 port map( A1 => n25998, A2 => n28479, Z => n26534);
   U10095 : INV_X2 port map( I => n26537, ZN => n7965);
   U10153 : OR2_X1 port map( A1 => n14290, A2 => n21403, Z => n4920);
   U10154 : XOR2_X1 port map( A1 => n20848, A2 => n30304, Z => n20671);
   U10259 : XOR2_X1 port map( A1 => n12474, A2 => n23228, Z => n12473);
   U10261 : XOR2_X1 port map( A1 => n13864, A2 => n20715, Z => n5184);
   U10269 : NAND2_X2 port map( A1 => n9158, A2 => n9156, ZN => n849);
   U10290 : NAND2_X1 port map( A1 => n16111, A2 => n25790, ZN => n12308);
   U10323 : XOR2_X1 port map( A1 => n26552, A2 => n12552, Z => n5166);
   U10326 : XOR2_X1 port map( A1 => n20736, A2 => n31043, Z => n26552);
   U10327 : XOR2_X1 port map( A1 => n19449, A2 => n27824, Z => n8435);
   U10344 : AOI22_X2 port map( A1 => n3463, A2 => n3462, B1 => n26555, B2 => 
                           n28316, ZN => n3461);
   U10350 : XOR2_X1 port map( A1 => n3177, A2 => n3178, Z => n3176);
   U10360 : XOR2_X1 port map( A1 => n26556, A2 => n119, Z => n24174);
   U10362 : XOR2_X1 port map( A1 => n24405, A2 => n24649, Z => n26556);
   U10364 : OR2_X1 port map( A1 => n4632, A2 => n9469, Z => n18126);
   U10369 : XOR2_X1 port map( A1 => n4631, A2 => n29039, Z => n4632);
   U10379 : OAI21_X2 port map( A1 => n26557, A2 => n15849, B => n15850, ZN => 
                           n20329);
   U10385 : NOR2_X2 port map( A1 => n15614, A2 => n14014, ZN => n12904);
   U10407 : XOR2_X1 port map( A1 => n21006, A2 => n16636, Z => n27573);
   U10410 : OAI21_X2 port map( A1 => n4469, A2 => n4471, B => n20446, ZN => 
                           n21006);
   U10431 : XOR2_X1 port map( A1 => n23272, A2 => n25355, Z => n643);
   U10433 : AND2_X1 port map( A1 => n10599, A2 => n5822, Z => n4248);
   U10437 : OAI21_X2 port map( A1 => n26563, A2 => n6468, B => n33120, ZN => 
                           n6722);
   U10445 : AOI21_X2 port map( A1 => n14163, A2 => n33787, B => n14162, ZN => 
                           n8726);
   U10464 : XOR2_X1 port map( A1 => n23369, A2 => n27201, Z => n16776);
   U10478 : OAI22_X1 port map( A1 => n15167, A2 => n776, B1 => n22964, B2 => 
                           n15852, ZN => n22820);
   U10479 : OAI22_X2 port map( A1 => n26569, A2 => n17621, B1 => n7143, B2 => 
                           n25905, ZN => n5412);
   U10489 : XOR2_X1 port map( A1 => n5315, A2 => n5314, Z => n5527);
   U10494 : AOI22_X2 port map( A1 => n18807, A2 => n17465, B1 => n18809, B2 => 
                           n27909, ZN => n6332);
   U10496 : XOR2_X1 port map( A1 => n26571, A2 => n16634, Z => Ciphertext(162))
                           ;
   U10501 : AND2_X1 port map( A1 => n17370, A2 => n16699, Z => n6030);
   U10513 : NOR2_X1 port map( A1 => n16023, A2 => n30291, ZN => n26572);
   U10555 : NAND2_X2 port map( A1 => n26022, A2 => n26581, ZN => n25664);
   U10560 : XOR2_X1 port map( A1 => n2365, A2 => n7222, Z => n2364);
   U10567 : OAI21_X1 port map( A1 => n26290, A2 => n23862, B => n13068, ZN => 
                           n6235);
   U10584 : INV_X2 port map( I => n26583, ZN => n13829);
   U10591 : XOR2_X1 port map( A1 => n19520, A2 => n4157, Z => n26583);
   U10629 : AOI21_X2 port map( A1 => n15397, A2 => n13072, B => n15395, ZN => 
                           n19754);
   U10649 : AOI21_X2 port map( A1 => n26589, A2 => n26588, B => n10480, ZN => 
                           n24004);
   U10650 : NAND2_X1 port map( A1 => n17881, A2 => n32308, ZN => n26588);
   U10661 : NAND2_X2 port map( A1 => n3994, A2 => n14001, ZN => n24926);
   U10668 : AOI21_X2 port map( A1 => n28242, A2 => n13641, B => n718, ZN => 
                           n13636);
   U10682 : NAND2_X1 port map( A1 => n26829, A2 => n5141, ZN => n15422);
   U10685 : NOR2_X2 port map( A1 => n11861, A2 => n31317, ZN => n16016);
   U10692 : INV_X2 port map( I => n26593, ZN => n29279);
   U10693 : XOR2_X1 port map( A1 => n391, A2 => n13358, Z => n26593);
   U10694 : NAND2_X2 port map( A1 => n11199, A2 => n11198, ZN => n10072);
   U10713 : AOI22_X1 port map( A1 => n25812, A2 => n25816, B1 => n17642, B2 => 
                           n25811, ZN => n25813);
   U10731 : INV_X2 port map( I => n26597, ZN => n5961);
   U10755 : NOR2_X1 port map( A1 => n26611, A2 => n16115, ZN => n17115);
   U10757 : AOI21_X2 port map( A1 => n25951, A2 => n28347, B => n23796, ZN => 
                           n2234);
   U10795 : INV_X2 port map( I => n18373, ZN => n2614);
   U10832 : AND2_X1 port map( A1 => n32253, A2 => n26640, Z => n3643);
   U10888 : NAND2_X1 port map( A1 => n16187, A2 => n16188, ZN => n26614);
   U10896 : NAND2_X1 port map( A1 => n2728, A2 => n15038, ZN => n27064);
   U10905 : NOR2_X2 port map( A1 => n15376, A2 => n5160, ZN => n28525);
   U10917 : NOR2_X1 port map( A1 => n16954, A2 => n29980, ZN => n16953);
   U10924 : XOR2_X1 port map( A1 => n3599, A2 => n16504, Z => n26617);
   U10934 : NAND2_X2 port map( A1 => n14758, A2 => n9256, ZN => n24520);
   U10951 : NOR2_X2 port map( A1 => n29224, A2 => n25678, ZN => n25675);
   U10997 : XOR2_X1 port map( A1 => n23041, A2 => n23040, Z => n23720);
   U11006 : XOR2_X1 port map( A1 => n22237, A2 => n21931, Z => n10704);
   U11010 : OAI21_X1 port map( A1 => n22641, A2 => n22484, B => n9544, ZN => 
                           n27445);
   U11018 : OAI21_X1 port map( A1 => n9026, A2 => n9027, B => n19974, ZN => 
                           n26644);
   U11021 : INV_X1 port map( I => n26644, ZN => n7474);
   U11026 : AOI21_X1 port map( A1 => n3468, A2 => n17077, B => n1135, ZN => 
                           n26625);
   U11053 : INV_X4 port map( I => n25488, ZN => n25462);
   U11054 : NAND2_X1 port map( A1 => n4151, A2 => n13343, ZN => n28275);
   U11061 : INV_X2 port map( I => n26630, ZN => n3004);
   U11068 : NOR2_X2 port map( A1 => n27446, A2 => n26631, ZN => n24014);
   U11081 : XOR2_X1 port map( A1 => n20808, A2 => n20807, Z => n4849);
   U11086 : XOR2_X1 port map( A1 => n30219, A2 => n20869, Z => n20807);
   U11087 : NAND2_X2 port map( A1 => n3499, A2 => n28380, ZN => n3515);
   U11104 : AOI21_X1 port map( A1 => n17120, A2 => n754, B => n4407, ZN => 
                           n26637);
   U11130 : NAND2_X2 port map( A1 => n12650, A2 => n10100, ZN => n10099);
   U11133 : NOR2_X2 port map( A1 => n13502, A2 => n13501, ZN => n26640);
   U11152 : XOR2_X1 port map( A1 => n23471, A2 => n23472, Z => n26642);
   U11155 : XOR2_X1 port map( A1 => n26643, A2 => n17723, Z => Ciphertext(157))
                           ;
   U11163 : AOI22_X1 port map( A1 => n25750, A2 => n1979, B1 => n25734, B2 => 
                           n25733, ZN => n26643);
   U11181 : XOR2_X1 port map( A1 => n2875, A2 => n438, Z => n26646);
   U11198 : NAND3_X2 port map( A1 => n26648, A2 => n18536, A3 => n32530, ZN => 
                           n19284);
   U11203 : NAND2_X1 port map( A1 => n18256, A2 => n18745, ZN => n26648);
   U11218 : XOR2_X1 port map( A1 => n7452, A2 => n12805, Z => n7646);
   U11235 : AOI22_X2 port map( A1 => n28638, A2 => n29715, B1 => n3206, B2 => 
                           n13475, ZN => n19197);
   U11263 : XOR2_X1 port map( A1 => n26655, A2 => n22039, Z => n10816);
   U11272 : XOR2_X1 port map( A1 => n28730, A2 => n16060, Z => n26655);
   U11279 : NAND2_X2 port map( A1 => n4050, A2 => n4051, ZN => n13911);
   U11294 : NAND2_X2 port map( A1 => n9786, A2 => n9785, ZN => n19224);
   U11300 : NAND2_X2 port map( A1 => n5004, A2 => n10968, ZN => n4342);
   U11308 : XOR2_X1 port map( A1 => n24838, A2 => n24552, Z => n18188);
   U11360 : AOI21_X2 port map( A1 => n26007, A2 => n26741, B => n942, ZN => 
                           n26663);
   U11370 : XOR2_X1 port map( A1 => n12736, A2 => n26665, Z => n12735);
   U11372 : XOR2_X1 port map( A1 => n20858, A2 => n10737, Z => n26665);
   U11394 : NAND2_X1 port map( A1 => n17467, A2 => n34089, ZN => n12911);
   U11395 : INV_X1 port map( I => n26666, ZN => n27862);
   U11400 : NAND3_X1 port map( A1 => n25621, A2 => n11944, A3 => n25707, ZN => 
                           n26666);
   U11402 : XOR2_X1 port map( A1 => n27733, A2 => n23239, Z => n2048);
   U11406 : NAND2_X1 port map( A1 => n2107, A2 => n18676, ZN => n3586);
   U11424 : XOR2_X1 port map( A1 => n12495, A2 => n21921, Z => n6329);
   U11435 : XOR2_X1 port map( A1 => n29285, A2 => n7458, Z => n3237);
   U11458 : NAND2_X2 port map( A1 => n11560, A2 => n15836, ZN => n22032);
   U11462 : INV_X2 port map( I => n10791, ZN => n26677);
   U11464 : NAND2_X2 port map( A1 => n26635, A2 => n26677, ZN => n7990);
   U11465 : NOR2_X2 port map( A1 => n1156, A2 => n26278, ZN => n20321);
   U11466 : NOR2_X2 port map( A1 => n28381, A2 => n28382, ZN => n28380);
   U11467 : XOR2_X1 port map( A1 => n29072, A2 => n27823, Z => n7020);
   U11476 : OAI21_X2 port map( A1 => n31975, A2 => n20480, B => n26471, ZN => 
                           n20316);
   U11483 : AOI21_X2 port map( A1 => n1184, A2 => n13381, B => n26680, ZN => 
                           n6170);
   U11484 : NAND2_X2 port map( A1 => n14651, A2 => n18638, ZN => n6138);
   U11486 : NAND2_X2 port map( A1 => n1214, A2 => n25889, ZN => n7350);
   U11540 : XNOR2_X1 port map( A1 => n20680, A2 => n20693, ZN => n20859);
   U11575 : NAND2_X2 port map( A1 => n25995, A2 => n30288, ZN => n25882);
   U11589 : XOR2_X1 port map( A1 => n3143, A2 => n3144, Z => n15012);
   U11592 : NOR2_X1 port map( A1 => n2902, A2 => n2692, ZN => n14438);
   U11593 : NOR2_X1 port map( A1 => n22674, A2 => n22467, ZN => n8252);
   U11609 : XOR2_X1 port map( A1 => n26692, A2 => n8312, Z => n26691);
   U11616 : XOR2_X1 port map( A1 => n3175, A2 => n26693, Z => n22504);
   U11617 : XOR2_X1 port map( A1 => n21906, A2 => n25945, Z => n26693);
   U11632 : NAND2_X2 port map( A1 => n26696, A2 => n19882, ZN => n20515);
   U11664 : XOR2_X1 port map( A1 => n3399, A2 => n26702, Z => n577);
   U11695 : BUF_X2 port map( I => n709, Z => n26710);
   U11745 : XOR2_X1 port map( A1 => n26711, A2 => n16523, Z => Ciphertext(13));
   U11774 : OAI21_X2 port map( A1 => n10686, A2 => n15002, B => n151, ZN => 
                           n14996);
   U11801 : OR2_X1 port map( A1 => n13297, A2 => n5736, Z => n7386);
   U11821 : OR2_X1 port map( A1 => n26040, A2 => n26717, Z => n3179);
   U11840 : XOR2_X1 port map( A1 => n14215, A2 => n26055, Z => n4895);
   U11860 : XOR2_X1 port map( A1 => n10201, A2 => n16662, Z => n23412);
   U11888 : NAND2_X2 port map( A1 => n19298, A2 => n27831, ZN => n14606);
   U11895 : INV_X2 port map( I => n11570, ZN => n7929);
   U11902 : NAND2_X2 port map( A1 => n15768, A2 => n17924, ZN => n11570);
   U11906 : NOR2_X1 port map( A1 => n15094, A2 => n16348, ZN => n16347);
   U11907 : NAND2_X2 port map( A1 => n19006, A2 => n18939, ZN => n27077);
   U11922 : BUF_X2 port map( I => n24883, Z => n25019);
   U11930 : INV_X4 port map( I => n3004, ZN => n23940);
   U11947 : XOR2_X1 port map( A1 => n12595, A2 => n14901, Z => n15343);
   U11977 : NOR2_X1 port map( A1 => n21646, A2 => n28580, ZN => n21647);
   U11998 : XOR2_X1 port map( A1 => n29652, A2 => n15566, Z => n27643);
   U12015 : XOR2_X1 port map( A1 => n30306, A2 => n22243, Z => n28835);
   U12018 : INV_X2 port map( I => n26738, ZN => n17688);
   U12025 : XOR2_X1 port map( A1 => n26740, A2 => n17663, Z => n25115);
   U12026 : XOR2_X1 port map( A1 => n24788, A2 => n1226, Z => n26740);
   U12037 : NAND3_X2 port map( A1 => n12876, A2 => n12875, A3 => n1182, ZN => 
                           n26742);
   U12045 : NAND2_X1 port map( A1 => n10359, A2 => n25995, ZN => n26744);
   U12058 : NOR2_X1 port map( A1 => n20067, A2 => n13080, ZN => n27542);
   U12069 : OAI21_X1 port map( A1 => n12904, A2 => n24305, B => n26747, ZN => 
                           n24302);
   U12070 : AOI21_X1 port map( A1 => n27430, A2 => n12904, B => n1241, ZN => 
                           n26747);
   U12081 : NAND2_X1 port map( A1 => n867, A2 => n18078, ZN => n2512);
   U12094 : XOR2_X1 port map( A1 => n4955, A2 => n22790, Z => n14382);
   U12129 : INV_X2 port map( I => n19597, ZN => n26751);
   U12132 : AND2_X1 port map( A1 => n15149, A2 => n21147, Z => n11151);
   U12142 : NAND2_X1 port map( A1 => n3646, A2 => n7929, ZN => n7926);
   U12147 : XOR2_X1 port map( A1 => n26755, A2 => n15904, Z => n27824);
   U12149 : XOR2_X1 port map( A1 => n27825, A2 => n19448, Z => n26755);
   U12178 : NOR2_X2 port map( A1 => n2395, A2 => n7986, ZN => n2394);
   U12185 : INV_X1 port map( I => n2380, ZN => n26758);
   U12239 : NAND2_X2 port map( A1 => n4909, A2 => n4913, ZN => n5348);
   U12275 : XOR2_X1 port map( A1 => n13145, A2 => n24409, Z => n27951);
   U12295 : NOR2_X1 port map( A1 => n15456, A2 => n12315, ZN => n12118);
   U12301 : INV_X2 port map( I => n26761, ZN => n579);
   U12303 : XOR2_X1 port map( A1 => n5768, A2 => n503, Z => n26761);
   U12307 : NAND2_X2 port map( A1 => n26762, A2 => n3594, ZN => n16297);
   U12310 : NAND2_X2 port map( A1 => n3597, A2 => n3598, ZN => n22500);
   U12311 : XOR2_X1 port map( A1 => n10631, A2 => n13470, Z => n13309);
   U12315 : XOR2_X1 port map( A1 => n26765, A2 => n22102, Z => n4161);
   U12322 : OAI21_X1 port map( A1 => n2536, A2 => n14940, B => n25995, ZN => 
                           n5300);
   U12329 : NOR2_X2 port map( A1 => n7732, A2 => n11970, ZN => n13495);
   U12372 : NAND2_X2 port map( A1 => n25670, A2 => n25675, ZN => n25691);
   U12376 : OAI22_X2 port map( A1 => n9083, A2 => n17370, B1 => n18993, B2 => 
                           n13252, ZN => n26768);
   U12378 : XOR2_X1 port map( A1 => n110, A2 => n7025, Z => n7024);
   U12382 : AND2_X1 port map( A1 => n19857, A2 => n20067, Z => n27541);
   U12394 : INV_X1 port map( I => n28504, ZN => n15824);
   U12395 : OR2_X1 port map( A1 => n28504, A2 => n31967, Z => n16251);
   U12402 : OR2_X1 port map( A1 => n5410, A2 => n25995, Z => n7425);
   U12404 : AND3_X1 port map( A1 => n22505, A2 => n22524, A3 => n8314, Z => 
                           n29026);
   U12408 : INV_X2 port map( I => n23144, ZN => n23841);
   U12421 : NAND2_X2 port map( A1 => n15137, A2 => n30995, ZN => n18477);
   U12422 : INV_X1 port map( I => n21214, ZN => n21215);
   U12441 : XOR2_X1 port map( A1 => n23241, A2 => n23533, Z => n9863);
   U12450 : AND2_X1 port map( A1 => n8083, A2 => n12231, Z => n26780);
   U12456 : OR2_X1 port map( A1 => n23843, A2 => n31796, Z => n14350);
   U12475 : NOR2_X1 port map( A1 => n4006, A2 => n1109, ZN => n16927);
   U12492 : XOR2_X1 port map( A1 => n9843, A2 => n28927, Z => n23210);
   U12493 : NAND2_X2 port map( A1 => n4542, A2 => n4543, ZN => n9843);
   U12499 : NOR2_X2 port map( A1 => n10373, A2 => n1384, ZN => n12744);
   U12510 : XNOR2_X1 port map( A1 => Key(93), A2 => Plaintext(93), ZN => n26791
                           );
   U12521 : OAI21_X2 port map( A1 => n17320, A2 => n15378, B => n17319, ZN => 
                           n19436);
   U12526 : NAND2_X2 port map( A1 => n8286, A2 => n14551, ZN => n24218);
   U12548 : AND2_X1 port map( A1 => n20334, A2 => n28261, Z => n12089);
   U12557 : XNOR2_X1 port map( A1 => n10075, A2 => n22080, ZN => n26822);
   U12576 : NAND2_X2 port map( A1 => n26799, A2 => n16414, ZN => n22919);
   U12590 : INV_X1 port map( I => n5373, ZN => n28740);
   U12617 : NAND2_X1 port map( A1 => n7040, A2 => n25734, ZN => n7039);
   U12620 : INV_X2 port map( I => n27105, ZN => n20541);
   U12625 : XOR2_X1 port map( A1 => n15618, A2 => n26807, Z => n15617);
   U12626 : XOR2_X1 port map( A1 => n2477, A2 => n371, Z => n26807);
   U12630 : OAI21_X2 port map( A1 => n28347, A2 => n4177, B => n25996, ZN => 
                           n26808);
   U12632 : NOR2_X1 port map( A1 => n6816, A2 => n25128, ZN => n27518);
   U12661 : INV_X2 port map( I => n20305, ZN => n20419);
   U12664 : AOI21_X1 port map( A1 => n31821, A2 => n11123, B => n13279, ZN => 
                           n18303);
   U12668 : INV_X2 port map( I => n26812, ZN => n13496);
   U12676 : XOR2_X1 port map( A1 => n9636, A2 => n26815, Z => n20102);
   U12705 : XOR2_X1 port map( A1 => n5279, A2 => n5280, Z => n5287);
   U12712 : XOR2_X1 port map( A1 => n26821, A2 => n22082, Z => n10681);
   U12718 : XOR2_X1 port map( A1 => n22081, A2 => n26822, Z => n26821);
   U12730 : NOR2_X2 port map( A1 => n24498, A2 => n24499, ZN => n24750);
   U12732 : NAND2_X1 port map( A1 => n13747, A2 => n10805, ZN => n26825);
   U12745 : OAI22_X2 port map( A1 => n31079, A2 => n11637, B1 => n29077, B2 => 
                           n8454, ZN => n11634);
   U12750 : XOR2_X1 port map( A1 => n23426, A2 => n23427, Z => n10674);
   U12757 : NOR3_X1 port map( A1 => n28704, A2 => n1168, A3 => n17670, ZN => 
                           n26827);
   U12765 : XOR2_X1 port map( A1 => n21006, A2 => n6431, Z => n20748);
   U12770 : INV_X2 port map( I => n19284, ZN => n28721);
   U12776 : NAND2_X2 port map( A1 => n1680, A2 => n1679, ZN => n20467);
   U12782 : XOR2_X1 port map( A1 => n3195, A2 => n19691, Z => n3652);
   U12796 : NAND2_X1 port map( A1 => n16265, A2 => n16266, ZN => n21104);
   U12800 : AOI21_X2 port map( A1 => n14867, A2 => n25123, B => n16607, ZN => 
                           n14866);
   U12807 : NAND2_X2 port map( A1 => n7310, A2 => n13622, ZN => n22890);
   U12810 : OR2_X1 port map( A1 => n9406, A2 => n6908, Z => n6013);
   U12813 : OAI22_X2 port map( A1 => n26078, A2 => n9146, B1 => n24347, B2 => 
                           n29043, ZN => n29143);
   U12852 : XOR2_X1 port map( A1 => n21896, A2 => n26096, Z => n26842);
   U12858 : XOR2_X1 port map( A1 => n26844, A2 => n12461, Z => n27004);
   U12861 : XOR2_X1 port map( A1 => n22165, A2 => n26845, Z => n26844);
   U12872 : INV_X2 port map( I => n26846, ZN => n17971);
   U12877 : OAI21_X2 port map( A1 => n11106, A2 => n7656, B => n26432, ZN => 
                           n1862);
   U12881 : NAND2_X2 port map( A1 => n27765, A2 => n21140, ZN => n21592);
   U12884 : XOR2_X1 port map( A1 => n27613, A2 => n26582, Z => n23514);
   U12910 : NAND3_X1 port map( A1 => n33750, A2 => n630, A3 => n26305, ZN => 
                           n21909);
   U12911 : AOI22_X2 port map( A1 => n26855, A2 => n1773, B1 => n22375, B2 => 
                           n1282, ZN => n9575);
   U12915 : OAI21_X1 port map( A1 => n23026, A2 => n26169, B => n16280, ZN => 
                           n26856);
   U12924 : XOR2_X1 port map( A1 => n32861, A2 => n24738, Z => n23151);
   U12925 : INV_X1 port map( I => n5826, ZN => n27302);
   U12953 : NOR2_X1 port map( A1 => n14102, A2 => n750, ZN => n14101);
   U12956 : XOR2_X1 port map( A1 => n29220, A2 => n7382, Z => n26865);
   U12961 : AOI22_X2 port map( A1 => n19992, A2 => n16681, B1 => n19993, B2 => 
                           n19943, ZN => n28786);
   U12963 : AOI22_X1 port map( A1 => n25492, A2 => n30047, B1 => n138, B2 => 
                           n4183, ZN => n25494);
   U12964 : XOR2_X1 port map( A1 => n23417, A2 => n23444, Z => n23497);
   U12974 : OAI21_X2 port map( A1 => n26023, A2 => n28634, B => n6144, ZN => 
                           n25330);
   U12993 : XOR2_X1 port map( A1 => n9269, A2 => n30314, Z => n27055);
   U13007 : XOR2_X1 port map( A1 => n11324, A2 => n26869, Z => n6502);
   U13009 : XOR2_X1 port map( A1 => n23457, A2 => n16402, Z => n26869);
   U13017 : OAI21_X1 port map( A1 => n28166, A2 => n16374, B => n16218, ZN => 
                           n14876);
   U13036 : XOR2_X1 port map( A1 => n9006, A2 => n462, Z => n26872);
   U13047 : NAND3_X2 port map( A1 => n27437, A2 => n29404, A3 => n9055, ZN => 
                           n26875);
   U13050 : XOR2_X1 port map( A1 => n26877, A2 => n16479, Z => Ciphertext(79));
   U13064 : NOR2_X2 port map( A1 => n27683, A2 => n18435, ZN => n8606);
   U13069 : NAND2_X2 port map( A1 => n26885, A2 => n16028, ZN => n23189);
   U13072 : NOR2_X1 port map( A1 => n22808, A2 => n11308, ZN => n26886);
   U13074 : INV_X1 port map( I => n22809, ZN => n26887);
   U13137 : XOR2_X1 port map( A1 => n10087, A2 => n22046, Z => n7640);
   U13146 : NAND2_X1 port map( A1 => n8544, A2 => n9375, ZN => n5116);
   U13155 : AND2_X1 port map( A1 => n15704, A2 => n28077, Z => n28613);
   U13156 : INV_X2 port map( I => n26896, ZN => n29256);
   U13157 : XOR2_X1 port map( A1 => n16770, A2 => n11982, Z => n26896);
   U13169 : XOR2_X1 port map( A1 => n9038, A2 => n26897, Z => n9037);
   U13170 : XOR2_X1 port map( A1 => n15877, A2 => n15, Z => n26897);
   U13193 : AND2_X1 port map( A1 => n30506, A2 => n15863, Z => n27326);
   U13241 : NOR3_X2 port map( A1 => n13475, A2 => n17311, A3 => n948, ZN => 
                           n28175);
   U13250 : INV_X1 port map( I => n27561, ZN => n28913);
   U13251 : NAND3_X2 port map( A1 => n258, A2 => n4290, A3 => n8143, ZN => 
                           n9141);
   U13252 : NOR2_X1 port map( A1 => n21529, A2 => n21697, ZN => n26913);
   U13266 : NAND2_X1 port map( A1 => n26724, A2 => n758, ZN => n5481);
   U13274 : NAND2_X1 port map( A1 => n6910, A2 => n25394, ZN => n26917);
   U13286 : INV_X1 port map( I => n22401, ZN => n4983);
   U13291 : NAND2_X1 port map( A1 => n17477, A2 => n10325, ZN => n10366);
   U13323 : NAND2_X2 port map( A1 => n22965, A2 => n14129, ZN => n22814);
   U13336 : XOR2_X1 port map( A1 => n1971, A2 => n859, Z => n22292);
   U13338 : AOI22_X2 port map( A1 => n26921, A2 => n33460, B1 => n25297, B2 => 
                           n28763, ZN => n15483);
   U13347 : XOR2_X1 port map( A1 => n22193, A2 => n26922, Z => n17487);
   U13348 : XOR2_X1 port map( A1 => n16619, A2 => n30314, Z => n26922);
   U13350 : XOR2_X1 port map( A1 => n6396, A2 => n32154, Z => n11528);
   U13356 : NAND2_X2 port map( A1 => n22615, A2 => n11308, ZN => n4399);
   U13361 : XOR2_X1 port map( A1 => n4660, A2 => n26923, Z => n666);
   U13362 : XOR2_X1 port map( A1 => n26924, A2 => n23249, Z => n26923);
   U13385 : OAI21_X1 port map( A1 => n26051, A2 => n1318, B => n26927, ZN => 
                           n14674);
   U13399 : INV_X2 port map( I => n26930, ZN => n13308);
   U13414 : INV_X2 port map( I => n22048, ZN => n26931);
   U13422 : OAI22_X2 port map( A1 => n5694, A2 => n13605, B1 => n11120, B2 => 
                           n5693, ZN => n20634);
   U13426 : XOR2_X1 port map( A1 => n26934, A2 => n26933, Z => n27880);
   U13436 : XOR2_X1 port map( A1 => n5742, A2 => n26936, Z => n1708);
   U13437 : INV_X1 port map( I => n16604, ZN => n26936);
   U13442 : NAND2_X2 port map( A1 => n11873, A2 => n14623, ZN => n5742);
   U13448 : XOR2_X1 port map( A1 => n2981, A2 => n26004, Z => n2978);
   U13449 : NOR3_X2 port map( A1 => n34131, A2 => n3236, A3 => n31760, ZN => 
                           n6958);
   U13450 : OAI21_X2 port map( A1 => n6101, A2 => n4489, B => n26937, ZN => 
                           n22870);
   U13452 : INV_X2 port map( I => n9890, ZN => n26938);
   U13464 : AOI22_X2 port map( A1 => n6858, A2 => n6859, B1 => n16681, B2 => 
                           n19944, ZN => n8118);
   U13466 : XOR2_X1 port map( A1 => n12878, A2 => n17929, Z => n23245);
   U13469 : OAI22_X2 port map( A1 => n6964, A2 => n896, B1 => n13142, B2 => 
                           n6965, ZN => n17929);
   U13487 : OAI21_X2 port map( A1 => n14653, A2 => n14654, B => n13686, ZN => 
                           n27242);
   U13490 : AOI21_X2 port map( A1 => n21274, A2 => n21273, B => n21272, ZN => 
                           n16327);
   U13491 : AOI21_X2 port map( A1 => n22892, A2 => n23037, B => n899, ZN => 
                           n8149);
   U13512 : NAND2_X2 port map( A1 => n16663, A2 => n23542, ZN => n16066);
   U13513 : OR2_X1 port map( A1 => n4274, A2 => n27838, Z => n5684);
   U13517 : XOR2_X1 port map( A1 => n15560, A2 => n26941, Z => n12595);
   U13518 : XOR2_X1 port map( A1 => n26942, A2 => n22248, Z => n26941);
   U13527 : NAND2_X2 port map( A1 => n1602, A2 => n18977, ZN => n15074);
   U13529 : XOR2_X1 port map( A1 => n29162, A2 => n26945, Z => n28373);
   U13536 : XOR2_X1 port map( A1 => n17128, A2 => n32024, Z => n26945);
   U13539 : XOR2_X1 port map( A1 => n26947, A2 => n11289, Z => n29273);
   U13543 : XOR2_X1 port map( A1 => n5382, A2 => n26118, Z => n26947);
   U13546 : NAND3_X1 port map( A1 => n25788, A2 => n25796, A3 => n12611, ZN => 
                           n26948);
   U13547 : NAND2_X2 port map( A1 => n9323, A2 => n26950, ZN => n26949);
   U13563 : OAI21_X2 port map( A1 => n23722, A2 => n23349, B => n9443, ZN => 
                           n18077);
   U13565 : NOR2_X1 port map( A1 => n2512, A2 => n31873, ZN => n26953);
   U13575 : XOR2_X1 port map( A1 => n2388, A2 => n3727, Z => n2982);
   U13588 : NOR2_X2 port map( A1 => n772, A2 => n31129, ZN => n4489);
   U13592 : XOR2_X1 port map( A1 => n19709, A2 => n19397, Z => n17953);
   U13595 : XOR2_X1 port map( A1 => n22085, A2 => n26957, Z => n10873);
   U13611 : NAND2_X2 port map( A1 => n26958, A2 => n4854, ZN => n20374);
   U13617 : OAI21_X1 port map( A1 => n25556, A2 => n28760, B => n28759, ZN => 
                           n28758);
   U13619 : AOI21_X2 port map( A1 => n30502, A2 => n22706, B => n26960, ZN => 
                           n13814);
   U13631 : XOR2_X1 port map( A1 => n26426, A2 => n32893, Z => n27548);
   U13644 : NAND2_X2 port map( A1 => n25914, A2 => n25913, ZN => n25923);
   U13651 : XOR2_X1 port map( A1 => n23275, A2 => n24623, Z => n23174);
   U13652 : NOR2_X2 port map( A1 => n13289, A2 => n13288, ZN => n23275);
   U13665 : XOR2_X1 port map( A1 => n8893, A2 => n26111, Z => n8892);
   U13670 : NAND2_X2 port map( A1 => n13918, A2 => n11057, ZN => n27763);
   U13686 : XOR2_X1 port map( A1 => n24682, A2 => n13614, Z => n14897);
   U13689 : XOR2_X1 port map( A1 => n20736, A2 => n20953, Z => n20808);
   U13690 : OAI21_X2 port map( A1 => n5879, A2 => n5909, B => n12194, ZN => 
                           n17947);
   U13695 : NOR2_X2 port map( A1 => n27460, A2 => n19014, ZN => n19699);
   U13697 : NAND2_X1 port map( A1 => n12777, A2 => n23912, ZN => n26967);
   U13698 : XOR2_X1 port map( A1 => n9459, A2 => n21993, Z => n1713);
   U13731 : OR2_X1 port map( A1 => n3157, A2 => n30130, Z => n10613);
   U13740 : NOR2_X1 port map( A1 => n9690, A2 => n5074, ZN => n14589);
   U13741 : NAND2_X1 port map( A1 => n15228, A2 => n16098, ZN => n13971);
   U13746 : NAND2_X1 port map( A1 => n13766, A2 => n13765, ZN => n26974);
   U13752 : NAND2_X2 port map( A1 => n7474, A2 => n7473, ZN => n9025);
   U13756 : XOR2_X1 port map( A1 => n14296, A2 => n21023, Z => n26977);
   U13761 : INV_X2 port map( I => n26978, ZN => n700);
   U13763 : XOR2_X1 port map( A1 => n11171, A2 => n11169, Z => n26978);
   U13776 : NAND2_X1 port map( A1 => n21285, A2 => n29303, ZN => n27431);
   U13790 : INV_X2 port map( I => n26980, ZN => n1835);
   U13798 : XOR2_X1 port map( A1 => Plaintext(127), A2 => Key(127), Z => n26980
                           );
   U13814 : AND2_X1 port map( A1 => n5741, A2 => n24190, Z => n6770);
   U13828 : XOR2_X1 port map( A1 => n26983, A2 => n31912, Z => n616);
   U13829 : XOR2_X1 port map( A1 => n28490, A2 => n13612, Z => n26983);
   U13830 : XOR2_X1 port map( A1 => n28177, A2 => n2458, Z => n17826);
   U13853 : INV_X2 port map( I => n8040, ZN => n10360);
   U13872 : XOR2_X1 port map( A1 => n589, A2 => n3237, Z => n6556);
   U13887 : XOR2_X1 port map( A1 => n20449, A2 => n20748, Z => n1613);
   U13892 : NOR2_X2 port map( A1 => n11447, A2 => n11446, ZN => n6500);
   U13899 : NAND2_X1 port map( A1 => n24335, A2 => n24242, ZN => n11563);
   U13902 : OAI21_X2 port map( A1 => n26991, A2 => n27889, B => n904, ZN => 
                           n6836);
   U13903 : NAND3_X1 port map( A1 => n1896, A2 => n25717, A3 => n26992, ZN => 
                           n25719);
   U13905 : INV_X2 port map( I => n1102, ZN => n23393);
   U13909 : NOR2_X2 port map( A1 => n26995, A2 => n26994, ZN => n1102);
   U13914 : XOR2_X1 port map( A1 => n20049, A2 => n20050, Z => n21221);
   U13920 : AND2_X1 port map( A1 => n23944, A2 => n16961, Z => n16676);
   U13928 : NAND3_X2 port map( A1 => n7777, A2 => n5776, A3 => n664, ZN => 
                           n9220);
   U13929 : XOR2_X1 port map( A1 => n16303, A2 => n19682, Z => n19486);
   U13934 : XOR2_X1 port map( A1 => n19744, A2 => n3568, Z => n16303);
   U13936 : NAND3_X2 port map( A1 => n4212, A2 => n4211, A3 => n17021, ZN => 
                           n26998);
   U13942 : NAND2_X2 port map( A1 => n27752, A2 => n29314, ZN => n14978);
   U13951 : OAI21_X2 port map( A1 => n27865, A2 => n22904, B => n18177, ZN => 
                           n23247);
   U13957 : INV_X4 port map( I => n5073, ZN => n761);
   U13961 : NAND2_X2 port map( A1 => n14627, A2 => n15641, ZN => n2726);
   U13967 : NOR2_X2 port map( A1 => n777, A2 => n32898, ZN => n11756);
   U13973 : NOR2_X2 port map( A1 => n3312, A2 => n10572, ZN => n21350);
   U13975 : NAND2_X2 port map( A1 => n14719, A2 => n2821, ZN => n20428);
   U13977 : NOR2_X2 port map( A1 => n3527, A2 => n3525, ZN => n2821);
   U13997 : XOR2_X1 port map( A1 => n7535, A2 => n28144, Z => n10770);
   U13998 : OAI21_X2 port map( A1 => n27010, A2 => n11187, B => n21421, ZN => 
                           n14236);
   U14001 : XOR2_X1 port map( A1 => n27011, A2 => n721, Z => n23490);
   U14004 : INV_X2 port map( I => n27012, ZN => n599);
   U14006 : NOR2_X1 port map( A1 => n8270, A2 => n28847, ZN => n29080);
   U14011 : XOR2_X1 port map( A1 => n12924, A2 => n14077, Z => n12923);
   U14022 : XOR2_X1 port map( A1 => n27169, A2 => n27015, Z => n27014);
   U14025 : OR2_X1 port map( A1 => n579, A2 => n29250, Z => n10484);
   U14031 : INV_X4 port map( I => n9280, ZN => n5178);
   U14033 : XOR2_X1 port map( A1 => n3568, A2 => n14588, Z => n19726);
   U14035 : NAND2_X2 port map( A1 => n25440, A2 => n25441, ZN => n25429);
   U14040 : XOR2_X1 port map( A1 => n21992, A2 => n22013, Z => n13873);
   U14054 : XOR2_X1 port map( A1 => n20907, A2 => n21028, Z => n3617);
   U14075 : NOR2_X2 port map( A1 => n2705, A2 => n2706, ZN => n8506);
   U14082 : XOR2_X1 port map( A1 => n23507, A2 => n27708, Z => n4413);
   U14086 : AND2_X1 port map( A1 => n23968, A2 => n23969, Z => n27026);
   U14097 : NAND4_X1 port map( A1 => n25440, A2 => n25442, A3 => n25439, A4 => 
                           n25441, ZN => n25443);
   U14112 : NAND2_X2 port map( A1 => n13800, A2 => n14950, ZN => n6442);
   U14115 : NAND2_X2 port map( A1 => n5973, A2 => n22654, ZN => n23137);
   U14125 : OR2_X1 port map( A1 => n25675, A2 => n25686, Z => n25685);
   U14166 : NAND3_X1 port map( A1 => n17087, A2 => n23723, A3 => n23738, ZN => 
                           n28506);
   U14167 : XOR2_X1 port map( A1 => n6168, A2 => n24809, Z => n24405);
   U14169 : NAND2_X2 port map( A1 => n6167, A2 => n6166, ZN => n24809);
   U14170 : XOR2_X1 port map( A1 => n27613, A2 => n27126, Z => n27041);
   U14173 : XOR2_X1 port map( A1 => n27190, A2 => n22131, Z => n22136);
   U14174 : XOR2_X1 port map( A1 => n22192, A2 => n22130, Z => n27190);
   U14181 : XOR2_X1 port map( A1 => n3280, A2 => n27042, Z => n17799);
   U14183 : AOI22_X2 port map( A1 => n12886, A2 => n2990, B1 => n16318, B2 => 
                           n11323, ZN => n11322);
   U14195 : NAND2_X1 port map( A1 => n5327, A2 => n17649, ZN => n17553);
   U14204 : NAND2_X2 port map( A1 => n27044, A2 => n2992, ZN => n24315);
   U14212 : NAND2_X1 port map( A1 => n24168, A2 => n5454, ZN => n3984);
   U14219 : XOR2_X1 port map( A1 => n27047, A2 => n1424, Z => Ciphertext(80));
   U14224 : AOI22_X2 port map( A1 => n3297, A2 => n28649, B1 => n3296, B2 => 
                           n33132, ZN => n1565);
   U14228 : INV_X2 port map( I => n27050, ZN => n4577);
   U14229 : XOR2_X1 port map( A1 => n4578, A2 => n4579, Z => n27050);
   U14231 : XOR2_X1 port map( A1 => n16998, A2 => n23165, Z => n27052);
   U14232 : XOR2_X1 port map( A1 => n24621, A2 => n17325, Z => n13513);
   U14243 : XOR2_X1 port map( A1 => n20815, A2 => n21018, Z => n27054);
   U14252 : XOR2_X1 port map( A1 => n11836, A2 => n23295, Z => n11822);
   U14253 : XOR2_X1 port map( A1 => n23519, A2 => n23294, Z => n11836);
   U14283 : INV_X2 port map( I => n27058, ZN => n14083);
   U14307 : OR2_X1 port map( A1 => n7425, A2 => n25879, Z => n7265);
   U14315 : XOR2_X1 port map( A1 => n27063, A2 => n25319, Z => Ciphertext(94));
   U14318 : XOR2_X1 port map( A1 => n19483, A2 => n26002, Z => n19305);
   U14325 : AOI21_X2 port map( A1 => n27066, A2 => n11376, B => n22280, ZN => 
                           n22785);
   U14329 : OAI21_X2 port map( A1 => n8479, A2 => n29115, B => n27652, ZN => 
                           n27067);
   U14341 : XOR2_X1 port map( A1 => n22970, A2 => n30993, Z => n7011);
   U14344 : AOI21_X2 port map( A1 => n15730, A2 => n15729, B => n14680, ZN => 
                           n22970);
   U14350 : XOR2_X1 port map( A1 => n24456, A2 => n24457, Z => n27072);
   U14364 : INV_X2 port map( I => n7453, ZN => n21241);
   U14383 : NAND2_X2 port map( A1 => n27392, A2 => n29131, ZN => n24138);
   U14385 : XOR2_X1 port map( A1 => n27081, A2 => n27080, Z => n28151);
   U14387 : XOR2_X1 port map( A1 => n8432, A2 => n23243, Z => n27081);
   U14391 : XOR2_X1 port map( A1 => n3491, A2 => n27082, Z => n416);
   U14392 : XOR2_X1 port map( A1 => n33971, A2 => n26701, Z => n27082);
   U14393 : AND2_X1 port map( A1 => n28123, A2 => n15038, Z => n9734);
   U14414 : XOR2_X1 port map( A1 => n6151, A2 => n6152, Z => n14255);
   U14423 : XOR2_X1 port map( A1 => n30193, A2 => n9904, Z => n19575);
   U14431 : XOR2_X1 port map( A1 => n23313, A2 => n17500, Z => n12950);
   U14452 : INV_X1 port map( I => n22933, ZN => n27088);
   U14462 : XOR2_X1 port map( A1 => n1302, A2 => n22027, Z => n8680);
   U14475 : BUF_X2 port map( I => n11622, Z => n6034);
   U14492 : XOR2_X1 port map( A1 => n22043, A2 => n10155, Z => n10154);
   U14494 : XOR2_X1 port map( A1 => n22173, A2 => n22196, Z => n22043);
   U14502 : NAND2_X2 port map( A1 => n4167, A2 => n4168, ZN => n15043);
   U14507 : XOR2_X1 port map( A1 => n4448, A2 => n20908, Z => n27091);
   U14530 : OAI22_X1 port map( A1 => n10009, A2 => n10012, B1 => n10385, B2 => 
                           n30557, ZN => n27092);
   U14531 : NAND2_X2 port map( A1 => n17364, A2 => n14, ZN => n2843);
   U14534 : INV_X2 port map( I => n1696, ZN => n8100);
   U14537 : XOR2_X1 port map( A1 => n1698, A2 => n29079, Z => n1696);
   U14539 : NOR2_X1 port map( A1 => n14881, A2 => n22522, ZN => n27094);
   U14542 : XNOR2_X1 port map( A1 => n12789, A2 => n21994, ZN => n22193);
   U14563 : AOI21_X1 port map( A1 => n28973, A2 => n28972, B => n27532, ZN => 
                           n28494);
   U14580 : NOR2_X2 port map( A1 => n28455, A2 => n25902, ZN => n10085);
   U14582 : NAND3_X2 port map( A1 => n20290, A2 => n20289, A3 => n20292, ZN => 
                           n14821);
   U14586 : AOI21_X2 port map( A1 => n28167, A2 => n28166, B => n34132, ZN => 
                           n15749);
   U14590 : XOR2_X1 port map( A1 => n22311, A2 => n12621, Z => n8405);
   U14592 : XOR2_X1 port map( A1 => Key(47), A2 => Plaintext(47), Z => n28946);
   U14600 : XOR2_X1 port map( A1 => n15489, A2 => n15487, Z => n28765);
   U14607 : NOR2_X2 port map( A1 => n19135, A2 => n15126, ZN => n19654);
   U14619 : NAND2_X2 port map( A1 => n4801, A2 => n4804, ZN => n11193);
   U14629 : XOR2_X1 port map( A1 => n24792, A2 => n27100, Z => n17663);
   U14630 : XOR2_X1 port map( A1 => n24790, A2 => n27101, Z => n27100);
   U14631 : INV_X1 port map( I => n25648, ZN => n27101);
   U14645 : XOR2_X1 port map( A1 => n10172, A2 => n8562, Z => n10170);
   U14651 : XOR2_X1 port map( A1 => n12675, A2 => n24786, Z => n24817);
   U14653 : OAI21_X2 port map( A1 => n9658, A2 => n9659, B => n23996, ZN => 
                           n24786);
   U14658 : XOR2_X1 port map( A1 => n32880, A2 => n25436, Z => n15923);
   U14662 : XOR2_X1 port map( A1 => n24821, A2 => n24822, Z => n25242);
   U14670 : AOI21_X2 port map( A1 => n2726, A2 => n1218, B => n16276, ZN => 
                           n1547);
   U14678 : OAI21_X2 port map( A1 => n7147, A2 => n6427, B => n8603, ZN => 
                           n8602);
   U14687 : NAND2_X1 port map( A1 => n17273, A2 => n7925, ZN => n5568);
   U14689 : OAI22_X2 port map( A1 => n3529, A2 => n27111, B1 => n761, B2 => 
                           n2089, ZN => n3527);
   U14697 : NOR2_X2 port map( A1 => n4871, A2 => n28449, ZN => n23430);
   U14703 : OR2_X1 port map( A1 => n17239, A2 => n28705, Z => n12565);
   U14712 : INV_X4 port map( I => n27214, ZN => n7492);
   U14721 : INV_X2 port map( I => n11934, ZN => n16397);
   U14726 : OAI21_X1 port map( A1 => n25559, A2 => n14944, B => n28758, ZN => 
                           n15292);
   U14742 : NOR3_X1 port map( A1 => n24311, A2 => n7503, A3 => n9962, ZN => 
                           n27982);
   U14746 : NAND3_X2 port map( A1 => n24017, A2 => n24016, A3 => n24018, ZN => 
                           n27115);
   U14747 : NAND3_X1 port map( A1 => n24017, A2 => n24016, A3 => n24018, ZN => 
                           n24832);
   U14758 : INV_X1 port map( I => n28761, ZN => n28760);
   U14760 : NAND2_X1 port map( A1 => n16092, A2 => n16595, ZN => n29020);
   U14767 : NAND2_X1 port map( A1 => n28244, A2 => n28243, ZN => n25471);
   U14773 : NAND3_X1 port map( A1 => n4183, A2 => n25476, A3 => n25470, ZN => 
                           n28244);
   U14777 : NAND2_X1 port map( A1 => n25405, A2 => n25412, ZN => n28738);
   U14781 : NOR2_X1 port map( A1 => n15665, A2 => n8616, ZN => n29098);
   U14800 : NAND2_X1 port map( A1 => n16684, A2 => n20561, ZN => n19906);
   U14809 : AND2_X1 port map( A1 => n8238, A2 => n14195, Z => n5376);
   U14817 : NOR2_X1 port map( A1 => n25302, A2 => n25229, ZN => n1858);
   U14820 : OAI21_X1 port map( A1 => n14959, A2 => n4245, B => n26020, ZN => 
                           n25017);
   U14829 : INV_X1 port map( I => n23043, ZN => n28356);
   U14834 : OR2_X1 port map( A1 => n16425, A2 => n25570, Z => n11852);
   U14835 : INV_X2 port map( I => n30783, ZN => n2088);
   U14845 : AND2_X1 port map( A1 => n1218, A2 => n15641, Z => n25186);
   U14849 : NAND2_X1 port map( A1 => n25611, A2 => n25612, ZN => n10266);
   U14850 : INV_X1 port map( I => n9982, ZN => n25612);
   U14851 : NAND2_X1 port map( A1 => n750, A2 => n25368, ZN => n15479);
   U14852 : NAND3_X1 port map( A1 => n9731, A2 => n9733, A3 => n25323, ZN => 
                           n27330);
   U14855 : AOI22_X1 port map( A1 => n25539, A2 => n12088, B1 => n9917, B2 => 
                           n15481, ZN => n15480);
   U14856 : NAND2_X1 port map( A1 => n14454, A2 => n17382, ZN => n3033);
   U14865 : NOR2_X1 port map( A1 => n27926, A2 => n14454, ZN => n689);
   U14895 : AND2_X1 port map( A1 => n8555, A2 => n4415, Z => n4416);
   U14896 : NOR2_X1 port map( A1 => n17336, A2 => n32092, ZN => n17335);
   U14907 : NAND3_X1 port map( A1 => n25651, A2 => n25666, A3 => n7087, ZN => 
                           n7086);
   U14918 : INV_X1 port map( I => n24181, ZN => n14111);
   U14919 : NOR2_X1 port map( A1 => n25378, A2 => n25369, ZN => n25360);
   U14949 : NOR2_X1 port map( A1 => n27162, A2 => n25858, ZN => n405);
   U14951 : OR2_X1 port map( A1 => n15496, A2 => n25409, Z => n27119);
   U14952 : AND2_X1 port map( A1 => n5343, A2 => n17873, Z => n27121);
   U14957 : NAND2_X1 port map( A1 => n25394, A2 => n25238, ZN => n15756);
   U14958 : INV_X1 port map( I => n19122, ZN => n1055);
   U14962 : XOR2_X1 port map( A1 => n9623, A2 => n9621, Z => n27122);
   U14964 : NAND2_X1 port map( A1 => n31236, A2 => n25557, ZN => n28761);
   U14965 : OAI22_X1 port map( A1 => n25559, A2 => n25552, B1 => n25544, B2 => 
                           n25543, ZN => n16869);
   U14989 : INV_X1 port map( I => n11781, ZN => n5206);
   U14997 : NOR2_X1 port map( A1 => n4041, A2 => n3673, ZN => n14802);
   U15000 : NAND2_X2 port map( A1 => n3724, A2 => n3725, ZN => n27123);
   U15002 : AOI21_X1 port map( A1 => n24996, A2 => n7941, B => n5113, ZN => 
                           n12035);
   U15003 : CLKBUF_X4 port map( I => n25110, Z => n8219);
   U15011 : AOI21_X1 port map( A1 => n8248, A2 => n7809, B => n8178, ZN => 
                           n15973);
   U15037 : NAND2_X2 port map( A1 => n803, A2 => n29317, ZN => n22914);
   U15045 : NAND3_X1 port map( A1 => n25105, A2 => n787, A3 => n32857, ZN => 
                           n3824);
   U15046 : INV_X1 port map( I => n23403, ZN => n27552);
   U15048 : INV_X1 port map( I => n25617, ZN => n25602);
   U15062 : OR2_X1 port map( A1 => n8277, A2 => n9920, Z => n13068);
   U15063 : NAND2_X1 port map( A1 => n28904, A2 => n20545, ZN => n20548);
   U15080 : NAND2_X1 port map( A1 => n24780, A2 => n17382, ZN => n28520);
   U15081 : OAI21_X1 port map( A1 => n18648, A2 => n16474, B => n4200, ZN => 
                           n27561);
   U15107 : XNOR2_X1 port map( A1 => Plaintext(77), A2 => Key(77), ZN => n27129
                           );
   U15116 : NAND2_X1 port map( A1 => n13037, A2 => n13035, ZN => n27132);
   U15133 : AOI21_X1 port map( A1 => n21306, A2 => n21305, B => n21303, ZN => 
                           n21101);
   U15144 : NAND2_X2 port map( A1 => n9166, A2 => n9167, ZN => n28350);
   U15152 : OR2_X2 port map( A1 => n17378, A2 => n17379, Z => n27134);
   U15161 : NOR2_X1 port map( A1 => n29180, A2 => n33325, ZN => n13230);
   U15162 : NAND2_X2 port map( A1 => n723, A2 => n27719, ZN => n22897);
   U15168 : CLKBUF_X1 port map( I => n6552, Z => n5254);
   U15175 : AOI21_X1 port map( A1 => n17068, A2 => n24283, B => n16356, ZN => 
                           n24284);
   U15191 : NAND2_X1 port map( A1 => n24436, A2 => n25699, ZN => n17863);
   U15196 : OR2_X1 port map( A1 => n24919, A2 => n15569, Z => n17480);
   U15198 : INV_X1 port map( I => n24919, ZN => n1200);
   U15199 : XOR2_X1 port map( A1 => n10659, A2 => n11148, Z => n27136);
   U15201 : NAND2_X2 port map( A1 => n12597, A2 => n12596, ZN => n23332);
   U15204 : NAND3_X2 port map( A1 => n2870, A2 => n2868, A3 => n2867, ZN => 
                           n27137);
   U15207 : NAND3_X2 port map( A1 => n2870, A2 => n2868, A3 => n2867, ZN => 
                           n27138);
   U15228 : INV_X1 port map( I => n29121, ZN => n27277);
   U15230 : OR2_X2 port map( A1 => n495, A2 => n10891, Z => n9651);
   U15246 : NAND2_X1 port map( A1 => n6068, A2 => n6067, ZN => n27139);
   U15251 : OAI21_X1 port map( A1 => n29222, A2 => n10680, B => n14339, ZN => 
                           n3475);
   U15253 : NAND2_X1 port map( A1 => n10680, A2 => n809, ZN => n15812);
   U15267 : OR2_X2 port map( A1 => n11605, A2 => n4036, Z => n10578);
   U15276 : INV_X1 port map( I => n19335, ZN => n9538);
   U15278 : AOI21_X1 port map( A1 => n5491, A2 => n19335, B => n14597, ZN => 
                           n1452);
   U15289 : XOR2_X1 port map( A1 => n20740, A2 => n20739, Z => n27143);
   U15304 : NAND2_X1 port map( A1 => n25360, A2 => n25368, ZN => n28516);
   U15308 : XOR2_X1 port map( A1 => Key(92), A2 => Plaintext(92), Z => n27146);
   U15313 : NAND3_X2 port map( A1 => n8797, A2 => n10765, A3 => n10764, ZN => 
                           n27147);
   U15314 : OR2_X2 port map( A1 => n10000, A2 => n7116, Z => n10765);
   U15321 : INV_X2 port map( I => n16568, ZN => n20147);
   U15326 : INV_X1 port map( I => n22940, ZN => n22938);
   U15330 : OR2_X2 port map( A1 => n13862, A2 => n636, Z => n14231);
   U15335 : OAI21_X1 port map( A1 => n7361, A2 => n24327, B => n24245, ZN => 
                           n5286);
   U15341 : INV_X1 port map( I => n16053, ZN => n17051);
   U15355 : NOR2_X2 port map( A1 => n4665, A2 => n4664, ZN => n27151);
   U15371 : NAND2_X1 port map( A1 => n28801, A2 => n16280, ZN => n11494);
   U15374 : NAND2_X2 port map( A1 => n20364, A2 => n20363, ZN => n4225);
   U15378 : NAND2_X1 port map( A1 => n27188, A2 => n18151, ZN => n9197);
   U15389 : XOR2_X1 port map( A1 => n2366, A2 => n2364, Z => n27154);
   U15394 : NAND2_X1 port map( A1 => n16008, A2 => n19156, ZN => n28372);
   U15398 : XOR2_X1 port map( A1 => n15982, A2 => n27155, Z => n265);
   U15399 : XNOR2_X1 port map( A1 => n27115, A2 => n32981, ZN => n27155);
   U15402 : AOI21_X1 port map( A1 => n14813, A2 => n15437, B => n7188, ZN => 
                           n28403);
   U15403 : NAND2_X1 port map( A1 => n32898, A2 => n28099, ZN => n3043);
   U15404 : NAND2_X1 port map( A1 => n27127, A2 => n33681, ZN => n1890);
   U15411 : BUF_X4 port map( I => n20054, Z => n8616);
   U15424 : OAI21_X1 port map( A1 => n19051, A2 => n19000, B => n27877, ZN => 
                           n27156);
   U15435 : INV_X2 port map( I => n8721, ZN => n22599);
   U15437 : INV_X2 port map( I => n25145, ZN => n17595);
   U15442 : OAI21_X1 port map( A1 => n15376, A2 => n888, B => n33544, ZN => 
                           n15375);
   U15443 : NOR3_X1 port map( A1 => n12304, A2 => n25072, A3 => n25078, ZN => 
                           n27925);
   U15449 : AND2_X2 port map( A1 => n11063, A2 => n11272, Z => n15506);
   U15453 : INV_X2 port map( I => n33117, ZN => n741);
   U15460 : OR3_X2 port map( A1 => n1052, A2 => n26600, A3 => n7251, Z => 
                           n18123);
   U15466 : NOR2_X1 port map( A1 => n4405, A2 => n1379, ZN => n3243);
   U15467 : INV_X2 port map( I => n4405, ZN => n7415);
   U15484 : OAI21_X1 port map( A1 => n19058, A2 => n7345, B => n5625, ZN => 
                           n4914);
   U15501 : INV_X1 port map( I => n25789, ZN => n29168);
   U15507 : NOR2_X1 port map( A1 => n24969, A2 => n3843, ZN => n2129);
   U15523 : NOR2_X1 port map( A1 => n25221, A2 => n7515, ZN => n10941);
   U15526 : CLKBUF_X4 port map( I => n16045, Z => n28898);
   U15545 : NAND2_X1 port map( A1 => n20401, A2 => n20569, ZN => n27904);
   U15546 : NAND2_X1 port map( A1 => n6765, A2 => n21876, ZN => n27706);
   U15571 : OR2_X1 port map( A1 => n4019, A2 => n24148, Z => n8963);
   U15579 : NOR2_X1 port map( A1 => n11571, A2 => n7929, ZN => n25253);
   U15580 : INV_X2 port map( I => n6402, ZN => n1075);
   U15591 : OR2_X1 port map( A1 => n22781, A2 => n11383, Z => n11382);
   U15600 : AOI21_X1 port map( A1 => n28659, A2 => n28697, B => n8040, ZN => 
                           n8038);
   U15627 : XOR2_X1 port map( A1 => n11349, A2 => n7717, Z => n27165);
   U15628 : AND2_X2 port map( A1 => n28083, A2 => n4221, Z => n27166);
   U15676 : NAND3_X1 port map( A1 => n6997, A2 => n6995, A3 => n6994, ZN => 
                           n5415);
   U15683 : NAND2_X1 port map( A1 => n6431, A2 => n20755, ZN => n7951);
   U15692 : INV_X1 port map( I => n7093, ZN => n28715);
   U15701 : NAND2_X1 port map( A1 => n20045, A2 => n19907, ZN => n4143);
   U15706 : NAND2_X2 port map( A1 => n10486, A2 => n10489, ZN => n27169);
   U15709 : XOR2_X1 port map( A1 => n3819, A2 => n12672, Z => n27170);
   U15713 : OAI21_X1 port map( A1 => n5274, A2 => n22919, B => n32967, ZN => 
                           n11539);
   U15726 : NAND2_X1 port map( A1 => n6555, A2 => n29043, ZN => n15437);
   U15729 : AND2_X1 port map( A1 => n19724, A2 => n14082, Z => n19902);
   U15735 : NAND3_X2 port map( A1 => n60, A2 => n22943, A3 => n22942, ZN => 
                           n27171);
   U15737 : NOR2_X1 port map( A1 => n24164, A2 => n2826, ZN => n27525);
   U15739 : NOR2_X1 port map( A1 => n19249, A2 => n7810, ZN => n14332);
   U15751 : INV_X1 port map( I => n31394, ZN => n23442);
   U15755 : OAI22_X1 port map( A1 => n27719, A2 => n17211, B1 => n31325, B2 => 
                           n723, ZN => n3826);
   U15763 : NOR2_X1 port map( A1 => n23066, A2 => n23065, ZN => n10643);
   U15774 : INV_X1 port map( I => n23066, ZN => n1281);
   U15779 : INV_X2 port map( I => n12446, ZN => n12445);
   U15781 : INV_X2 port map( I => n14029, ZN => n4041);
   U15783 : NOR3_X1 port map( A1 => n7232, A2 => n7776, A3 => n7775, ZN => 
                           n27177);
   U15802 : AOI21_X2 port map( A1 => n5055, A2 => n5619, B => n5054, ZN => 
                           n27179);
   U15803 : NAND2_X2 port map( A1 => n21537, A2 => n8196, ZN => n27180);
   U15817 : NAND3_X1 port map( A1 => n25199, A2 => n32873, A3 => n9294, ZN => 
                           n7854);
   U15818 : INV_X2 port map( I => n32877, ZN => n15068);
   U15828 : NOR2_X1 port map( A1 => n12482, A2 => n17928, ZN => n152);
   U15829 : NAND2_X1 port map( A1 => n1161, A2 => n9759, ZN => n20014);
   U15833 : XOR2_X1 port map( A1 => n8747, A2 => n8745, Z => n27181);
   U15839 : NAND2_X2 port map( A1 => n27811, A2 => n4800, ZN => n27184);
   U15855 : INV_X1 port map( I => n25973, ZN => n12520);
   U15864 : OR2_X2 port map( A1 => n16778, A2 => n24565, Z => n25296);
   U15867 : OAI21_X1 port map( A1 => n1071, A2 => n27123, B => n9247, ZN => 
                           n11365);
   U15869 : NAND2_X1 port map( A1 => n27650, A2 => n24883, ZN => n27461);
   U15899 : NAND2_X1 port map( A1 => n10038, A2 => n32876, ZN => n37);
   U15902 : AOI21_X1 port map( A1 => n742, A2 => n741, B => n31961, ZN => 
                           n20161);
   U15905 : OR2_X1 port map( A1 => n31939, A2 => n25700, Z => n9805);
   U15906 : XNOR2_X1 port map( A1 => n7984, A2 => n28746, ZN => n27188);
   U15914 : NAND3_X2 port map( A1 => n8194, A2 => n8195, A3 => n12314, ZN => 
                           n1600);
   U15916 : AOI21_X1 port map( A1 => n7287, A2 => n23057, B => n3007, ZN => 
                           n2911);
   U15918 : NAND3_X2 port map( A1 => n26231, A2 => n31437, A3 => n28974, ZN => 
                           n8308);
   U15923 : AND2_X2 port map( A1 => n7043, A2 => n31939, Z => n7064);
   U15933 : INV_X1 port map( I => n18777, ZN => n954);
   U15937 : INV_X1 port map( I => n14899, ZN => n5980);
   U15951 : INV_X2 port map( I => n25023, ZN => n2092);
   U15952 : XOR2_X1 port map( A1 => n8939, A2 => n28663, Z => n25023);
   U15954 : MUX2_X1 port map( I0 => n33115, I1 => n22795, S => n13473, Z => 
                           n6964);
   U15975 : OAI21_X2 port map( A1 => n11091, A2 => n12743, B => n15015, ZN => 
                           n7146);
   U15988 : NOR2_X2 port map( A1 => n16165, A2 => n21662, ZN => n3379);
   U15991 : AOI21_X1 port map( A1 => n17595, A2 => n675, B => n25185, ZN => 
                           n17594);
   U15992 : INV_X2 port map( I => n27202, ZN => n2499);
   U15993 : XOR2_X1 port map( A1 => n2500, A2 => n2501, Z => n27202);
   U15995 : INV_X2 port map( I => n27203, ZN => n16792);
   U15996 : XOR2_X1 port map( A1 => n19651, A2 => n19384, Z => n27203);
   U16006 : OAI21_X2 port map( A1 => n27402, A2 => n22547, B => n22393, ZN => 
                           n22375);
   U16017 : AOI21_X1 port map( A1 => n25854, A2 => n14199, B => n10897, ZN => 
                           n25848);
   U16033 : NAND3_X1 port map( A1 => n25781, A2 => n16111, A3 => n32874, ZN => 
                           n25769);
   U16043 : NOR2_X1 port map( A1 => n10031, A2 => n15704, ZN => n27212);
   U16056 : NOR2_X2 port map( A1 => n7493, A2 => n27215, ZN => n27214);
   U16063 : NAND2_X2 port map( A1 => n27218, A2 => n11291, ZN => n196);
   U16064 : XOR2_X1 port map( A1 => n14250, A2 => n681, Z => n8562);
   U16069 : XOR2_X1 port map( A1 => n24617, A2 => n24421, Z => n14250);
   U16078 : XOR2_X1 port map( A1 => n27220, A2 => n17871, Z => n23319);
   U16102 : XOR2_X1 port map( A1 => n14796, A2 => n518, Z => n3812);
   U16118 : XOR2_X1 port map( A1 => n1902, A2 => n26031, Z => n27226);
   U16119 : BUF_X2 port map( I => n15455, Z => n27228);
   U16139 : NOR2_X2 port map( A1 => n24064, A2 => n16425, ZN => n24770);
   U16143 : XOR2_X1 port map( A1 => n27234, A2 => n23024, Z => n23746);
   U16147 : OR2_X2 port map( A1 => n9125, A2 => n27894, Z => n11752);
   U16148 : BUF_X2 port map( I => n16704, Z => n27236);
   U16161 : OAI21_X2 port map( A1 => n26035, A2 => n27238, B => n27237, ZN => 
                           n2080);
   U16169 : AND2_X1 port map( A1 => n6149, A2 => n31637, Z => n27590);
   U16172 : XOR2_X1 port map( A1 => n24372, A2 => n15982, Z => n28916);
   U16178 : AOI21_X1 port map( A1 => n1299, A2 => n16647, B => n857, ZN => 
                           n6064);
   U16190 : INV_X2 port map( I => n27244, ZN => n9234);
   U16196 : XOR2_X1 port map( A1 => n9235, A2 => n9679, Z => n27244);
   U16210 : AND2_X1 port map( A1 => n19315, A2 => n7197, Z => n28025);
   U16220 : NAND2_X1 port map( A1 => n11135, A2 => n15054, ZN => n11134);
   U16249 : NAND2_X2 port map( A1 => n18408, A2 => n27253, ZN => n13037);
   U16252 : NOR2_X1 port map( A1 => n17605, A2 => n27719, ZN => n17604);
   U16254 : AOI21_X1 port map( A1 => n21859, A2 => n21858, B => n21860, ZN => 
                           n18251);
   U16255 : INV_X2 port map( I => n27257, ZN => n11734);
   U16268 : NAND2_X1 port map( A1 => n5219, A2 => n27605, ZN => n5218);
   U16270 : NAND2_X1 port map( A1 => n17191, A2 => n26072, ZN => n13462);
   U16274 : NAND2_X2 port map( A1 => n15693, A2 => n15151, ZN => n7810);
   U16282 : NAND2_X2 port map( A1 => n27261, A2 => n18748, ZN => n19258);
   U16286 : XOR2_X1 port map( A1 => n10515, A2 => n15472, Z => n17523);
   U16300 : XOR2_X1 port map( A1 => n29415, A2 => n22042, Z => n27268);
   U16313 : NAND2_X1 port map( A1 => n17637, A2 => n1204, ZN => n17636);
   U16317 : XOR2_X1 port map( A1 => n9087, A2 => n8844, Z => n8843);
   U16321 : NAND2_X2 port map( A1 => n27271, A2 => n13422, ZN => n5942);
   U16328 : NAND2_X1 port map( A1 => n13421, A2 => n25588, ZN => n27271);
   U16335 : NAND2_X2 port map( A1 => n14425, A2 => n14423, ZN => n29130);
   U16339 : XOR2_X1 port map( A1 => n10815, A2 => n10814, Z => n10813);
   U16342 : XOR2_X1 port map( A1 => n19468, A2 => n27275, Z => n471);
   U16349 : XOR2_X1 port map( A1 => n28107, A2 => n27276, Z => n5640);
   U16352 : XOR2_X1 port map( A1 => n5847, A2 => n27277, Z => n27276);
   U16361 : NAND2_X1 port map( A1 => n27282, A2 => n27281, ZN => n7213);
   U16362 : INV_X1 port map( I => n24991, ZN => n27281);
   U16364 : XOR2_X1 port map( A1 => n28797, A2 => n1225, Z => n27283);
   U16369 : OAI22_X2 port map( A1 => n32095, A2 => n24304, B1 => n16039, B2 => 
                           n27284, ZN => n283);
   U16373 : OR2_X1 port map( A1 => n18145, A2 => n319, Z => n27284);
   U16387 : XOR2_X1 port map( A1 => n7131, A2 => n23516, Z => n27289);
   U16392 : NAND2_X2 port map( A1 => n15665, A2 => n8616, ZN => n17675);
   U16393 : NOR2_X2 port map( A1 => n19909, A2 => n870, ZN => n16132);
   U16397 : NOR2_X2 port map( A1 => n23560, A2 => n23561, ZN => n16305);
   U16407 : NAND2_X1 port map( A1 => n10435, A2 => n871, ZN => n10439);
   U16427 : NAND2_X2 port map( A1 => n27297, A2 => n21202, ZN => n5944);
   U16432 : NAND2_X2 port map( A1 => n7830, A2 => n21401, ZN => n27297);
   U16437 : OAI22_X2 port map( A1 => n1359, A2 => n20010, B1 => n16664, B2 => 
                           n12100, ZN => n3366);
   U16439 : AOI22_X2 port map( A1 => n12432, A2 => n28222, B1 => n23646, B2 => 
                           n23726, ZN => n27551);
   U16458 : NOR2_X1 port map( A1 => n18801, A2 => n32034, ZN => n4474);
   U16462 : INV_X2 port map( I => n17937, ZN => n18801);
   U16469 : XOR2_X1 port map( A1 => Plaintext(52), A2 => Key(52), Z => n17937);
   U16471 : NAND2_X2 port map( A1 => n28789, A2 => n14234, ZN => n28616);
   U16482 : NAND2_X2 port map( A1 => n27302, A2 => n27300, ZN => n20339);
   U16485 : NAND2_X2 port map( A1 => n5906, A2 => n21226, ZN => n2386);
   U16498 : XOR2_X1 port map( A1 => n29140, A2 => n8531, Z => n6689);
   U16508 : XOR2_X1 port map( A1 => n32809, A2 => n19716, Z => n8283);
   U16509 : XOR2_X1 port map( A1 => n19780, A2 => n8785, Z => n19716);
   U16513 : XOR2_X1 port map( A1 => n27308, A2 => n16696, Z => Ciphertext(133))
                           ;
   U16523 : OAI21_X1 port map( A1 => n27309, A2 => n24129, B => n24346, ZN => 
                           n3334);
   U16529 : INV_X2 port map( I => n27311, ZN => n6416);
   U16532 : XNOR2_X1 port map( A1 => Plaintext(176), A2 => Key(176), ZN => 
                           n27311);
   U16533 : XOR2_X1 port map( A1 => n27312, A2 => n22176, Z => n22363);
   U16553 : INV_X1 port map( I => n1533, ZN => n12041);
   U16554 : INV_X2 port map( I => n27315, ZN => n29116);
   U16558 : INV_X2 port map( I => n25473, ZN => n27315);
   U16568 : NAND2_X1 port map( A1 => n23853, A2 => n23852, ZN => n27320);
   U16582 : NOR2_X2 port map( A1 => n27334, A2 => n27662, ZN => n27660);
   U16587 : INV_X2 port map( I => n27324, ZN => n3601);
   U16591 : XOR2_X1 port map( A1 => Plaintext(27), A2 => Key(27), Z => n27324);
   U16592 : OAI22_X1 port map( A1 => n14564, A2 => n20630, B1 => n9062, B2 => 
                           n31471, ZN => n20216);
   U16607 : NOR2_X1 port map( A1 => n10217, A2 => n14080, ZN => n12528);
   U16615 : XOR2_X1 port map( A1 => n27330, A2 => n25324, Z => Ciphertext(95));
   U16627 : NAND2_X1 port map( A1 => n27332, A2 => n25977, ZN => n3225);
   U16630 : AND2_X2 port map( A1 => n24257, A2 => n4746, Z => n24232);
   U16639 : NOR3_X2 port map( A1 => n18805, A2 => n18349, A3 => n16122, ZN => 
                           n18374);
   U16688 : AOI21_X2 port map( A1 => n23669, A2 => n1250, B => n23953, ZN => 
                           n16842);
   U16689 : NAND2_X2 port map( A1 => n27731, A2 => n25021, ZN => n25057);
   U16702 : OAI21_X2 port map( A1 => n4422, A2 => n21367, B => n16311, ZN => 
                           n27337);
   U16725 : XOR2_X1 port map( A1 => n14613, A2 => n17914, Z => n17913);
   U16752 : XOR2_X1 port map( A1 => n4562, A2 => n4563, Z => n7022);
   U16758 : NAND3_X2 port map( A1 => n28672, A2 => n28670, A3 => n23651, ZN => 
                           n27341);
   U16769 : NAND2_X2 port map( A1 => n14890, A2 => n14888, ZN => n24790);
   U16773 : OR2_X1 port map( A1 => n33684, A2 => n21259, Z => n28256);
   U16777 : XOR2_X1 port map( A1 => n16002, A2 => n2452, Z => n27344);
   U16793 : XOR2_X1 port map( A1 => n6560, A2 => n6562, Z => n7738);
   U16794 : XNOR2_X1 port map( A1 => n28493, A2 => n28492, ZN => n27881);
   U16821 : NOR2_X2 port map( A1 => n24572, A2 => n24570, ZN => n12431);
   U16824 : NAND2_X2 port map( A1 => n16398, A2 => n16400, ZN => n24572);
   U16825 : INV_X1 port map( I => n4551, ZN => n27769);
   U16828 : OAI21_X1 port map( A1 => n11852, A2 => n24064, B => n27354, ZN => 
                           n9585);
   U16839 : XOR2_X1 port map( A1 => n20985, A2 => n15275, Z => n15668);
   U16877 : XOR2_X1 port map( A1 => n19734, A2 => n10810, Z => n7297);
   U16878 : XOR2_X1 port map( A1 => n19473, A2 => n13106, Z => n19734);
   U16887 : NAND2_X1 port map( A1 => n9663, A2 => n8243, ZN => n27358);
   U16890 : NAND2_X2 port map( A1 => n20441, A2 => n2650, ZN => n20917);
   U16898 : INV_X2 port map( I => n10835, ZN => n18059);
   U16900 : XOR2_X1 port map( A1 => n5529, A2 => n5530, Z => n10835);
   U16904 : XOR2_X1 port map( A1 => n10766, A2 => n31526, Z => n27361);
   U16919 : AND2_X1 port map( A1 => n23084, A2 => n23088, Z => n14192);
   U16920 : AND2_X1 port map( A1 => n667, A2 => n23843, Z => n13263);
   U16921 : NAND2_X2 port map( A1 => n27363, A2 => n20436, ZN => n3539);
   U16929 : XOR2_X1 port map( A1 => n16303, A2 => n19565, Z => n16302);
   U16935 : XOR2_X1 port map( A1 => n2750, A2 => n26016, Z => n27365);
   U16945 : AND2_X1 port map( A1 => n22955, A2 => n5035, Z => n22508);
   U16962 : NAND2_X1 port map( A1 => n25375, A2 => n25376, ZN => n4089);
   U16977 : XOR2_X1 port map( A1 => n28632, A2 => n21925, Z => n9267);
   U16993 : XOR2_X1 port map( A1 => n11143, A2 => n11144, Z => n11559);
   U17026 : XOR2_X1 port map( A1 => n3868, A2 => n2221, Z => n2367);
   U17041 : OAI21_X2 port map( A1 => n3604, A2 => n3603, B => n27381, ZN => 
                           n4665);
   U17042 : XNOR2_X1 port map( A1 => n1044, A2 => n8785, ZN => n28458);
   U17050 : NAND2_X1 port map( A1 => n22627, A2 => n22628, ZN => n22629);
   U17053 : NAND2_X2 port map( A1 => n2283, A2 => n11302, ZN => n19038);
   U17064 : OR2_X1 port map( A1 => n16868, A2 => n24257, Z => n9889);
   U17072 : INV_X4 port map( I => n29196, ZN => n10773);
   U17079 : XOR2_X1 port map( A1 => n23246, A2 => n27388, Z => n8069);
   U17083 : XOR2_X1 port map( A1 => n5904, A2 => n13638, Z => n27388);
   U17088 : AOI22_X2 port map( A1 => n15017, A2 => n976, B1 => n9734, B2 => 
                           n1249, ZN => n27392);
   U17108 : NOR2_X1 port map( A1 => n15189, A2 => n11959, ZN => n27398);
   U17130 : INV_X2 port map( I => n27401, ZN => n2019);
   U17131 : XOR2_X1 port map( A1 => Plaintext(149), A2 => Key(149), Z => n27401
                           );
   U17136 : NAND2_X2 port map( A1 => n27403, A2 => n18591, ZN => n8802);
   U17139 : AOI22_X2 port map( A1 => n1710, A2 => n11459, B1 => n1709, B2 => 
                           n14658, ZN => n27403);
   U17146 : NAND2_X1 port map( A1 => n27408, A2 => n32898, ZN => n9601);
   U17149 : NAND2_X1 port map( A1 => n21662, A2 => n4097, ZN => n27408);
   U17178 : AOI22_X2 port map( A1 => n18875, A2 => n10182, B1 => n1709, B2 => 
                           n18590, ZN => n18591);
   U17190 : NOR2_X2 port map( A1 => n28124, A2 => n17302, ZN => n12929);
   U17199 : XOR2_X1 port map( A1 => n8055, A2 => n29515, Z => n8054);
   U17234 : XOR2_X1 port map( A1 => Plaintext(112), A2 => Key(112), Z => n27428
                           );
   U17247 : OAI22_X2 port map( A1 => n2099, A2 => n18447, B1 => n18446, B2 => 
                           n18796, ZN => n19268);
   U17259 : XOR2_X1 port map( A1 => n23391, A2 => n16622, Z => n11835);
   U17262 : NAND2_X1 port map( A1 => n18844, A2 => n27747, ZN => n4925);
   U17273 : INV_X2 port map( I => n27435, ZN => n692);
   U17278 : NAND2_X2 port map( A1 => n8081, A2 => n6519, ZN => n23420);
   U17295 : NAND2_X2 port map( A1 => n6068, A2 => n6067, ZN => n20615);
   U17301 : INV_X2 port map( I => n27441, ZN => n13413);
   U17302 : OAI21_X1 port map( A1 => n16176, A2 => n27442, B => n782, ZN => 
                           n2771);
   U17312 : XOR2_X1 port map( A1 => n14337, A2 => n25428, Z => n27444);
   U17321 : INV_X2 port map( I => n27453, ZN => n3933);
   U17322 : AOI22_X1 port map( A1 => n15939, A2 => n12530, B1 => n14034, B2 => 
                           n22333, ZN => n14750);
   U17324 : XOR2_X1 port map( A1 => n4732, A2 => n18122, Z => n11427);
   U17326 : NOR2_X1 port map( A1 => n27456, A2 => n11201, ZN => n5002);
   U17328 : NAND2_X1 port map( A1 => n4999, A2 => n33425, ZN => n27456);
   U17344 : INV_X2 port map( I => n14577, ZN => n17078);
   U17348 : NAND2_X2 port map( A1 => n3924, A2 => n21067, ZN => n14577);
   U17351 : NOR2_X2 port map( A1 => n12341, A2 => n3380, ZN => n24682);
   U17374 : NAND2_X2 port map( A1 => n13390, A2 => n19355, ZN => n19280);
   U17380 : AND2_X1 port map( A1 => n28865, A2 => n22330, Z => n28456);
   U17390 : INV_X2 port map( I => n27471, ZN => n628);
   U17391 : XOR2_X1 port map( A1 => n3102, A2 => n3100, Z => n27471);
   U17419 : INV_X2 port map( I => n27475, ZN => n10059);
   U17420 : XOR2_X1 port map( A1 => n10060, A2 => n11488, Z => n27475);
   U17444 : INV_X4 port map( I => n29658, ZN => n28010);
   U17448 : XOR2_X1 port map( A1 => n10235, A2 => n10237, Z => n10236);
   U17473 : NAND2_X1 port map( A1 => n8336, A2 => n32862, ZN => n27480);
   U17482 : NOR2_X1 port map( A1 => n21170, A2 => n6957, ZN => n27482);
   U17484 : XOR2_X1 port map( A1 => n24616, A2 => n11722, Z => n15982);
   U17485 : NOR2_X2 port map( A1 => n11723, A2 => n11767, ZN => n24616);
   U17497 : INV_X2 port map( I => n27485, ZN => n9430);
   U17515 : XOR2_X1 port map( A1 => n27487, A2 => n16390, Z => Ciphertext(101))
                           ;
   U17520 : INV_X2 port map( I => n27490, ZN => n25339);
   U17525 : INV_X2 port map( I => n31468, ZN => n27491);
   U17529 : AOI21_X2 port map( A1 => n2878, A2 => n1610, B => n17396, ZN => 
                           n23967);
   U17537 : AND3_X1 port map( A1 => n15699, A2 => n29903, A3 => n32080, Z => 
                           n27993);
   U17541 : NAND2_X2 port map( A1 => n25999, A2 => n27033, ZN => n18753);
   U17543 : XOR2_X1 port map( A1 => n2331, A2 => n8456, Z => n10810);
   U17550 : XOR2_X1 port map( A1 => n9866, A2 => n9865, Z => n23696);
   U17583 : XOR2_X1 port map( A1 => n27505, A2 => n16636, Z => Ciphertext(28));
   U17587 : OAI22_X1 port map( A1 => n14318, A2 => n12035, B1 => n14320, B2 => 
                           n14322, ZN => n27505);
   U17603 : OR2_X1 port map( A1 => n23855, A2 => n9152, Z => n23690);
   U17616 : INV_X2 port map( I => n27147, ZN => n20857);
   U17618 : OAI21_X2 port map( A1 => n18472, A2 => n18471, B => n13846, ZN => 
                           n15148);
   U17621 : NAND2_X1 port map( A1 => n29376, A2 => n24069, ZN => n27735);
   U17625 : NAND2_X1 port map( A1 => n19053, A2 => n2581, ZN => n29102);
   U17634 : OAI22_X2 port map( A1 => n18622, A2 => n18331, B1 => n18330, B2 => 
                           n18329, ZN => n19053);
   U17635 : OAI21_X2 port map( A1 => n23798, A2 => n23570, B => n23797, ZN => 
                           n23571);
   U17636 : NOR2_X2 port map( A1 => n13963, A2 => n27509, ZN => n19222);
   U17657 : XNOR2_X1 port map( A1 => n19673, A2 => n11627, ZN => n29032);
   U17679 : XOR2_X1 port map( A1 => n24603, A2 => n24647, Z => n27516);
   U17680 : NAND2_X2 port map( A1 => n2929, A2 => n27517, ZN => n2928);
   U17689 : XNOR2_X1 port map( A1 => n32052, A2 => n20842, ZN => n20919);
   U17696 : INV_X2 port map( I => n7576, ZN => n27520);
   U17697 : NAND2_X2 port map( A1 => n10198, A2 => n16535, ZN => n7576);
   U17700 : NAND2_X1 port map( A1 => n21568, A2 => n3203, ZN => n21542);
   U17716 : NAND2_X1 port map( A1 => n27525, A2 => n7093, ZN => n7095);
   U17730 : INV_X2 port map( I => n14794, ZN => n27529);
   U17735 : XOR2_X1 port map( A1 => n24764, A2 => n13060, Z => n24687);
   U17742 : AND2_X1 port map( A1 => n25443, A2 => n25444, Z => n27531);
   U17751 : NOR2_X1 port map( A1 => n14912, A2 => n24141, ZN => n27534);
   U17756 : NAND2_X2 port map( A1 => n28944, A2 => n2680, ZN => n19289);
   U17760 : AND2_X1 port map( A1 => n7195, A2 => n30813, Z => n15632);
   U17771 : NOR2_X1 port map( A1 => n31894, A2 => n985, ZN => n5177);
   U17785 : XOR2_X1 port map( A1 => n27538, A2 => n2473, Z => n17829);
   U17788 : XOR2_X1 port map( A1 => n2476, A2 => n28513, Z => n27538);
   U17814 : XOR2_X1 port map( A1 => n9468, A2 => n24622, Z => n24768);
   U17826 : XOR2_X1 port map( A1 => n28940, A2 => n9387, Z => n622);
   U17853 : NAND2_X2 port map( A1 => n25739, A2 => n1597, ZN => n1979);
   U17855 : AOI21_X2 port map( A1 => n12989, A2 => n17557, B => n17649, ZN => 
                           n5052);
   U17892 : XOR2_X1 port map( A1 => n5149, A2 => n5148, Z => n5151);
   U17893 : XOR2_X1 port map( A1 => n19461, A2 => n17430, Z => n5149);
   U17894 : INV_X4 port map( I => n25116, ZN => n27651);
   U17897 : NOR2_X1 port map( A1 => n502, A2 => n5433, ZN => n6954);
   U17898 : AOI22_X2 port map( A1 => n28105, A2 => n28104, B1 => n9648, B2 => 
                           n7415, ZN => n27553);
   U17909 : OAI22_X1 port map( A1 => n10364, A2 => n18884, B1 => n18677, B2 => 
                           n17477, ZN => n4659);
   U17931 : XOR2_X1 port map( A1 => n5284, A2 => n10111, Z => n24803);
   U17948 : INV_X2 port map( I => n27563, ZN => n21505);
   U17950 : NOR2_X2 port map( A1 => n21265, A2 => n28375, ZN => n27563);
   U17976 : NAND2_X2 port map( A1 => n7942, A2 => n7943, ZN => n27566);
   U18012 : AOI21_X1 port map( A1 => n13200, A2 => n19178, B => n19181, ZN => 
                           n8906);
   U18026 : OR2_X1 port map( A1 => n24149, A2 => n32178, Z => n10446);
   U18027 : INV_X2 port map( I => n27570, ZN => n11821);
   U18035 : OAI21_X2 port map( A1 => n6511, A2 => n5119, B => n17445, ZN => 
                           n18912);
   U18036 : XOR2_X1 port map( A1 => n27571, A2 => n18269, Z => n15721);
   U18052 : XOR2_X1 port map( A1 => n27573, A2 => n29241, Z => n6079);
   U18088 : OAI21_X2 port map( A1 => n18749, A2 => n17073, B => n27582, ZN => 
                           n13160);
   U18114 : XNOR2_X1 port map( A1 => n22102, A2 => n25641, ZN => n27943);
   U18119 : XOR2_X1 port map( A1 => n28977, A2 => n26001, Z => n460);
   U18127 : XOR2_X1 port map( A1 => n19630, A2 => n4157, Z => n14817);
   U18130 : OAI21_X2 port map( A1 => n15629, A2 => n15842, B => n15627, ZN => 
                           n4157);
   U18131 : OAI21_X2 port map( A1 => n16318, A2 => n10579, B => n3179, ZN => 
                           n12886);
   U18172 : OR2_X2 port map( A1 => n29334, A2 => n15318, Z => n15051);
   U18175 : XOR2_X1 port map( A1 => n4287, A2 => n24810, Z => n29236);
   U18181 : OAI21_X2 port map( A1 => n27590, A2 => n27589, B => n27588, ZN => 
                           n13276);
   U18183 : INV_X4 port map( I => n33382, ZN => n27589);
   U18185 : NOR2_X2 port map( A1 => n31973, A2 => n8831, ZN => n8829);
   U18196 : NOR2_X1 port map( A1 => n5741, A2 => n24193, ZN => n27591);
   U18198 : XOR2_X1 port map( A1 => n27593, A2 => n9459, Z => n13833);
   U18199 : XOR2_X1 port map( A1 => n14237, A2 => n3030, Z => n27593);
   U18200 : NOR2_X2 port map( A1 => n10833, A2 => n16359, ZN => n16357);
   U18201 : NOR3_X2 port map( A1 => n32041, A2 => n24273, A3 => n13040, ZN => 
                           n24499);
   U18206 : AND2_X2 port map( A1 => n13960, A2 => n7702, Z => n690);
   U18210 : NAND2_X1 port map( A1 => n21663, A2 => n13828, ZN => n27594);
   U18218 : XOR2_X1 port map( A1 => n19784, A2 => n19783, Z => n16351);
   U18219 : INV_X2 port map( I => n29446, ZN => n27597);
   U18246 : AND2_X2 port map( A1 => n13391, A2 => n27745, Z => n14094);
   U18247 : OAI22_X2 port map( A1 => n16358, A2 => n18433, B1 => n18432, B2 => 
                           n5269, ZN => n27683);
   U18255 : INV_X2 port map( I => n25654, ZN => n25650);
   U18261 : NOR2_X2 port map( A1 => n13911, A2 => n27604, ZN => n9831);
   U18267 : XOR2_X1 port map( A1 => n12370, A2 => n21768, Z => n21769);
   U18277 : NAND2_X1 port map( A1 => n18184, A2 => n17416, ZN => n2802);
   U18295 : XOR2_X1 port map( A1 => n14094, A2 => n27607, Z => n15357);
   U18321 : NOR2_X1 port map( A1 => n8051, A2 => n947, ZN => n18715);
   U18358 : NAND2_X1 port map( A1 => n3181, A2 => n31862, ZN => n14813);
   U18389 : XOR2_X1 port map( A1 => n1714, A2 => n10979, Z => n9459);
   U18408 : NAND2_X2 port map( A1 => n28683, A2 => n14134, ZN => n20404);
   U18416 : INV_X1 port map( I => n17061, ZN => n28685);
   U18429 : NAND3_X1 port map( A1 => n19893, A2 => n14545, A3 => n19894, ZN => 
                           n27627);
   U18437 : OAI21_X2 port map( A1 => n31987, A2 => n18692, B => n952, ZN => 
                           n27628);
   U18438 : NOR2_X1 port map( A1 => n7418, A2 => n27629, ZN => n7420);
   U18441 : NOR2_X1 port map( A1 => n7417, A2 => n7415, ZN => n27629);
   U18488 : AOI22_X2 port map( A1 => n19902, A2 => n16637, B1 => n19903, B2 => 
                           n27938, ZN => n19904);
   U18491 : INV_X4 port map( I => n692, ZN => n25229);
   U18496 : BUF_X2 port map( I => n9592, Z => n27638);
   U18506 : AOI21_X2 port map( A1 => n2147, A2 => n19867, B => n2146, ZN => 
                           n14138);
   U18509 : NAND2_X1 port map( A1 => n18798, A2 => n7712, ZN => n7898);
   U18517 : NOR2_X1 port map( A1 => n18803, A2 => n12317, ZN => n27641);
   U18522 : XOR2_X1 port map( A1 => Plaintext(24), A2 => Key(24), Z => n15455);
   U18523 : INV_X2 port map( I => n27642, ZN => n632);
   U18526 : XOR2_X1 port map( A1 => n10461, A2 => n10462, Z => n27642);
   U18531 : XOR2_X1 port map( A1 => n27645, A2 => n32759, Z => n24855);
   U18535 : XOR2_X1 port map( A1 => n24645, A2 => n15671, Z => n27645);
   U18554 : BUF_X2 port map( I => n725, Z => n27652);
   U18564 : NAND2_X2 port map( A1 => n20619, A2 => n20620, ZN => n21029);
   U18569 : AOI21_X2 port map( A1 => n17542, A2 => n20024, B => n27654, ZN => 
                           n20345);
   U18575 : OAI22_X1 port map( A1 => n20123, A2 => n16595, B1 => n20022, B2 => 
                           n20021, ZN => n27654);
   U18576 : OR2_X2 port map( A1 => n22617, A2 => n15401, Z => n23753);
   U18611 : OR2_X1 port map( A1 => n25923, A2 => n14359, Z => n27659);
   U18613 : OAI22_X2 port map( A1 => n25348, A2 => n31941, B1 => n25347, B2 => 
                           n25346, ZN => n25376);
   U18616 : XOR2_X1 port map( A1 => n27664, A2 => n25131, Z => Ciphertext(59));
   U18618 : XOR2_X1 port map( A1 => n16200, A2 => n13907, Z => n4562);
   U18626 : AND2_X2 port map( A1 => n19053, A2 => n30663, Z => n12052);
   U18635 : OAI21_X2 port map( A1 => n7904, A2 => n7905, B => n22552, ZN => 
                           n27719);
   U18649 : NAND2_X2 port map( A1 => n15820, A2 => n21740, ZN => n22031);
   U18654 : OR2_X1 port map( A1 => n22641, A2 => n10725, Z => n5648);
   U18682 : XOR2_X1 port map( A1 => n17659, A2 => n27672, Z => n449);
   U18689 : AOI21_X2 port map( A1 => n13659, A2 => n15520, B => n29473, ZN => 
                           n13658);
   U18709 : NOR2_X1 port map( A1 => n298, A2 => n30281, ZN => n27680);
   U18733 : XOR2_X1 port map( A1 => n20958, A2 => n20959, Z => n8076);
   U18741 : BUF_X2 port map( I => n12951, Z => n27687);
   U18742 : NOR2_X2 port map( A1 => n10113, A2 => n865, ZN => n27688);
   U18752 : NAND2_X1 port map( A1 => n1279, A2 => n23017, ZN => n22963);
   U18753 : OR2_X1 port map( A1 => n22791, A2 => n14392, Z => n15391);
   U18755 : NAND3_X2 port map( A1 => n28442, A2 => n19024, A3 => n19026, ZN => 
                           n19658);
   U18767 : NAND2_X2 port map( A1 => n19302, A2 => n730, ZN => n27696);
   U18770 : NAND2_X2 port map( A1 => n23658, A2 => n23657, ZN => n12356);
   U18777 : NAND3_X1 port map( A1 => n867, A2 => n1156, A3 => n6679, ZN => 
                           n8996);
   U18784 : XOR2_X1 port map( A1 => n22195, A2 => n22193, Z => n11423);
   U18791 : XOR2_X1 port map( A1 => n27703, A2 => n1067, Z => Ciphertext(53));
   U18794 : AOI22_X1 port map( A1 => n3208, A2 => n25082, B1 => n1203, B2 => 
                           n5520, ZN => n27703);
   U18800 : NAND2_X2 port map( A1 => n16747, A2 => n19717, ZN => n6255);
   U18804 : XOR2_X1 port map( A1 => n702, A2 => n19539, Z => n17931);
   U18816 : NOR2_X2 port map( A1 => n18816, A2 => n18714, ZN => n27709);
   U18823 : XOR2_X1 port map( A1 => n28262, A2 => n20775, Z => n1848);
   U18828 : INV_X2 port map( I => n23157, ZN => n707);
   U18834 : INV_X2 port map( I => n20569, ZN => n816);
   U18843 : XOR2_X1 port map( A1 => n10685, A2 => n321, Z => n11172);
   U18850 : XOR2_X1 port map( A1 => n5402, A2 => n27717, Z => n5401);
   U18857 : OAI22_X2 port map( A1 => n19606, A2 => n3388, B1 => n9356, B2 => 
                           n826, ZN => n27718);
   U18862 : NAND2_X1 port map( A1 => n13312, A2 => n12323, ZN => n27720);
   U18873 : OR3_X1 port map( A1 => n4066, A2 => n19156, A3 => n18599, Z => 
                           n19160);
   U18878 : XOR2_X1 port map( A1 => n27721, A2 => n9475, Z => n3144);
   U18882 : XOR2_X1 port map( A1 => n3146, A2 => n24781, Z => n27721);
   U18892 : NAND2_X2 port map( A1 => n2903, A2 => n19934, ZN => n18078);
   U18906 : NAND2_X2 port map( A1 => n24179, A2 => n24178, ZN => n24512);
   U18913 : XOR2_X1 port map( A1 => n1612, A2 => n1613, Z => n21100);
   U18917 : NAND2_X2 port map( A1 => n7826, A2 => n27724, ZN => n13478);
   U18920 : OR2_X1 port map( A1 => n13481, A2 => n13482, Z => n27724);
   U18926 : XOR2_X1 port map( A1 => n26255, A2 => n11349, Z => n28541);
   U18936 : INV_X1 port map( I => n32052, ZN => n27729);
   U18944 : INV_X1 port map( I => n20674, ZN => n28803);
   U18952 : XOR2_X1 port map( A1 => n12801, A2 => n27728, Z => n5137);
   U18958 : NAND2_X2 port map( A1 => n6864, A2 => n19921, ZN => n19844);
   U18962 : NAND2_X2 port map( A1 => n12879, A2 => n20336, ZN => n20842);
   U18967 : INV_X2 port map( I => n27732, ZN => n10787);
   U18976 : XOR2_X1 port map( A1 => n15308, A2 => n24783, Z => n24173);
   U18980 : NAND3_X1 port map( A1 => n14795, A2 => n25222, A3 => n15340, ZN => 
                           n5174);
   U18983 : INV_X2 port map( I => n27736, ZN => n17305);
   U18992 : XOR2_X1 port map( A1 => n21992, A2 => n10205, Z => n7639);
   U19006 : XOR2_X1 port map( A1 => n16893, A2 => n30007, Z => n21986);
   U19011 : OAI21_X1 port map( A1 => n16749, A2 => n16750, B => n6516, ZN => 
                           n27745);
   U19017 : INV_X2 port map( I => n27747, ZN => n469);
   U19018 : XOR2_X1 port map( A1 => Plaintext(186), A2 => Key(186), Z => n27747
                           );
   U19025 : NAND2_X2 port map( A1 => n21956, A2 => n8853, ZN => n23301);
   U19033 : NAND2_X2 port map( A1 => n27756, A2 => n14924, ZN => n24087);
   U19034 : NOR2_X1 port map( A1 => n15330, A2 => n16276, ZN => n27758);
   U19035 : XOR2_X1 port map( A1 => n11337, A2 => n11338, Z => n13195);
   U19044 : NAND2_X2 port map( A1 => n1351, A2 => n20447, ZN => n20224);
   U19060 : XOR2_X1 port map( A1 => n23319, A2 => n3620, Z => n3619);
   U19068 : AOI22_X2 port map( A1 => n27769, A2 => n27768, B1 => n9506, B2 => 
                           n8120, ZN => n7925);
   U19085 : OAI22_X1 port map( A1 => n13568, A2 => n8450, B1 => n25985, B2 => 
                           n10227, ZN => n2517);
   U19086 : AOI21_X2 port map( A1 => n27775, A2 => n29329, B => n13835, ZN => 
                           n13834);
   U19094 : NAND2_X2 port map( A1 => n27776, A2 => n28084, ZN => n2902);
   U19097 : NAND2_X1 port map( A1 => n18303, A2 => n18304, ZN => n27776);
   U19100 : NAND2_X1 port map( A1 => n13953, A2 => n13952, ZN => n29095);
   U19102 : NOR2_X2 port map( A1 => n5704, A2 => n25975, ZN => n21716);
   U19126 : XOR2_X1 port map( A1 => n27375, A2 => n1592, Z => n27778);
   U19136 : AOI21_X1 port map( A1 => n7361, A2 => n24327, B => n28030, ZN => 
                           n28029);
   U19141 : AOI22_X2 port map( A1 => n23982, A2 => n28538, B1 => n5286, B2 => 
                           n24325, ZN => n24785);
   U19151 : AOI22_X2 port map( A1 => n12105, A2 => n28436, B1 => n14891, B2 => 
                           n5913, ZN => n14890);
   U19184 : NAND2_X2 port map( A1 => n10523, A2 => n20173, ZN => n17554);
   U19201 : INV_X2 port map( I => n27797, ZN => n18648);
   U19202 : XNOR2_X1 port map( A1 => Key(38), A2 => Plaintext(38), ZN => n27797
                           );
   U19209 : AND2_X1 port map( A1 => n18648, A2 => n18649, Z => n17113);
   U19214 : XOR2_X1 port map( A1 => n27243, A2 => n11897, Z => n22516);
   U19236 : XOR2_X1 port map( A1 => n5212, A2 => n27179, Z => n3491);
   U19242 : XOR2_X1 port map( A1 => n2362, A2 => n2363, Z => n2366);
   U19264 : XOR2_X1 port map( A1 => n412, A2 => n27804, Z => n2022);
   U19271 : XOR2_X1 port map( A1 => n1676, A2 => n26033, Z => n27804);
   U19273 : NAND2_X1 port map( A1 => n822, A2 => n13348, ZN => n27805);
   U19276 : XOR2_X1 port map( A1 => n11490, A2 => n19740, Z => n11222);
   U19302 : OAI22_X2 port map( A1 => n11050, A2 => n12680, B1 => n23786, B2 => 
                           n23785, ZN => n15692);
   U19328 : INV_X2 port map( I => n1266, ZN => n22953);
   U19333 : XOR2_X1 port map( A1 => n4291, A2 => n13298, Z => n14605);
   U19351 : INV_X2 port map( I => n27819, ZN => n16205);
   U19362 : OAI21_X1 port map( A1 => n3136, A2 => n24972, B => n3135, ZN => 
                           n3134);
   U19371 : XOR2_X1 port map( A1 => n15887, A2 => n24549, Z => n27823);
   U19376 : NOR2_X1 port map( A1 => n28954, A2 => n13735, ZN => n29004);
   U19399 : OR2_X1 port map( A1 => n8558, A2 => n20136, Z => n27829);
   U19413 : NAND2_X1 port map( A1 => n10501, A2 => n25608, ZN => n27833);
   U19427 : OAI22_X1 port map( A1 => n1376, A2 => n30501, B1 => n31254, B2 => 
                           n10943, ZN => n14354);
   U19438 : XOR2_X1 port map( A1 => n29262, A2 => n14684, Z => n335);
   U19449 : INV_X2 port map( I => n27838, ZN => n28668);
   U19450 : XNOR2_X1 port map( A1 => n7890, A2 => n28748, ZN => n27838);
   U19482 : OR2_X1 port map( A1 => n32747, A2 => n11086, Z => n28857);
   U19490 : XOR2_X1 port map( A1 => Plaintext(5), A2 => Key(5), Z => n27936);
   U19503 : XOR2_X1 port map( A1 => n28239, A2 => n21894, Z => n21896);
   U19522 : OAI22_X2 port map( A1 => n27845, A2 => n24285, B1 => n27500, B2 => 
                           n24284, ZN => n24478);
   U19523 : AND2_X1 port map( A1 => n28275, A2 => n4604, Z => n27845);
   U19526 : NAND2_X2 port map( A1 => n15965, A2 => n7736, ZN => n16144);
   U19530 : XOR2_X1 port map( A1 => n23366, A2 => n26116, Z => n28811);
   U19546 : XOR2_X1 port map( A1 => n227, A2 => n6924, Z => n2839);
   U19572 : XOR2_X1 port map( A1 => n22161, A2 => n22110, Z => n22019);
   U19575 : NAND2_X2 port map( A1 => n27857, A2 => n18438, ZN => n19355);
   U19597 : INV_X2 port map( I => n6168, ZN => n24526);
   U19598 : NAND2_X2 port map( A1 => n2939, A2 => n27998, ZN => n6168);
   U19599 : BUF_X2 port map( I => n23508, Z => n27860);
   U19600 : NOR2_X2 port map( A1 => n21, A2 => n21857, ZN => n21691);
   U19614 : NOR3_X1 port map( A1 => n6939, A2 => n25707, A3 => n25705, ZN => 
                           n27861);
   U19624 : XOR2_X1 port map( A1 => n17659, A2 => n20904, Z => n5282);
   U19626 : NAND2_X1 port map( A1 => n19287, A2 => n19021, ZN => n19026);
   U19660 : XNOR2_X1 port map( A1 => n8568, A2 => n16691, ZN => n29205);
   U19665 : NAND2_X2 port map( A1 => n27867, A2 => n13973, ZN => n13972);
   U19686 : NAND2_X2 port map( A1 => n580, A2 => n20614, ZN => n20455);
   U19720 : INV_X2 port map( I => n15734, ZN => n28190);
   U19724 : NOR2_X1 port map( A1 => n3495, A2 => n29158, ZN => n3494);
   U19735 : XOR2_X1 port map( A1 => n16590, A2 => n28457, Z => n578);
   U19738 : AND2_X1 port map( A1 => n21392, A2 => n27170, Z => n2602);
   U19752 : XOR2_X1 port map( A1 => n20982, A2 => n20891, Z => n20673);
   U19757 : NAND2_X1 port map( A1 => n27873, A2 => n27872, ZN => n25281);
   U19758 : NAND2_X1 port map( A1 => n30281, A2 => n25276, ZN => n27872);
   U19781 : OAI21_X2 port map( A1 => n12111, A2 => n16546, B => n14692, ZN => 
                           n28450);
   U19784 : XOR2_X1 port map( A1 => n22231, A2 => n29121, Z => n4763);
   U19790 : AND2_X1 port map( A1 => n14650, A2 => n14954, Z => n16810);
   U19807 : NOR2_X2 port map( A1 => n19301, A2 => n16354, ZN => n19085);
   U19809 : INV_X2 port map( I => n27883, ZN => n5191);
   U19815 : XOR2_X1 port map( A1 => n19558, A2 => n25998, Z => n27884);
   U19821 : NAND2_X1 port map( A1 => n28704, A2 => n4577, ZN => n18119);
   U19824 : NAND2_X2 port map( A1 => n1297, A2 => n22660, ZN => n22446);
   U19835 : XOR2_X1 port map( A1 => n16733, A2 => n32683, Z => n673);
   U19837 : AOI21_X2 port map( A1 => n24034, A2 => n24033, B => n24032, ZN => 
                           n16733);
   U19849 : AND2_X1 port map( A1 => n2180, A2 => n3994, Z => n24934);
   U19855 : NAND2_X2 port map( A1 => n14355, A2 => n274, ZN => n19698);
   U19875 : XOR2_X1 port map( A1 => n4944, A2 => n9434, Z => n27895);
   U19880 : MUX2_X1 port map( I0 => n27430, I1 => n12904, S => n24305, Z => 
                           n24034);
   U19883 : INV_X2 port map( I => n18146, ZN => n24305);
   U19884 : XOR2_X1 port map( A1 => n16989, A2 => n27896, Z => n11934);
   U19885 : XOR2_X1 port map( A1 => n673, A2 => n16394, Z => n27896);
   U19892 : NAND2_X2 port map( A1 => n8024, A2 => n30010, ZN => n19004);
   U19895 : NAND2_X2 port map( A1 => n10307, A2 => n10306, ZN => n8024);
   U19908 : NOR3_X2 port map( A1 => n10687, A2 => n13, A3 => n24042, ZN => 
                           n27899);
   U19929 : NAND2_X2 port map( A1 => n21617, A2 => n21614, ZN => n6489);
   U19933 : XOR2_X1 port map( A1 => n6373, A2 => n13844, Z => n23460);
   U19938 : INV_X2 port map( I => n27907, ZN => n29255);
   U19942 : XOR2_X1 port map( A1 => n6273, A2 => n8076, Z => n27907);
   U19948 : OAI21_X2 port map( A1 => n8222, A2 => n14081, B => n12472, ZN => 
                           n22968);
   U19962 : AOI21_X2 port map( A1 => n18478, A2 => n18477, B => n18476, ZN => 
                           n19461);
   U19964 : XOR2_X1 port map( A1 => n22037, A2 => n10887, Z => n8328);
   U19974 : NAND3_X2 port map( A1 => n15004, A2 => n437, A3 => n436, ZN => 
                           n19122);
   U19976 : NAND2_X2 port map( A1 => n27914, A2 => n26060, ZN => n14770);
   U19984 : NAND3_X1 port map( A1 => n53, A2 => n32481, A3 => n29774, ZN => 
                           n7834);
   U19994 : INV_X2 port map( I => n31324, ZN => n12500);
   U19997 : XOR2_X1 port map( A1 => n19433, A2 => n27919, Z => n3932);
   U19998 : XOR2_X1 port map( A1 => n33749, A2 => n27920, Z => n27919);
   U20003 : NAND2_X2 port map( A1 => n28309, A2 => n29667, ZN => n20283);
   U20015 : XOR2_X1 port map( A1 => n12048, A2 => n14908, Z => n19541);
   U20016 : NAND2_X2 port map( A1 => n13706, A2 => n13705, ZN => n19651);
   U20020 : XOR2_X1 port map( A1 => n14716, A2 => n27923, Z => n8249);
   U20048 : OR2_X1 port map( A1 => n20037, A2 => n27911, Z => n19835);
   U20049 : NAND2_X1 port map( A1 => n21204, A2 => n27955, ZN => n16197);
   U20051 : OAI21_X2 port map( A1 => n4539, A2 => n4538, B => n4536, ZN => 
                           n3421);
   U20057 : INV_X1 port map( I => n19460, ZN => n28453);
   U20070 : XOR2_X1 port map( A1 => n15028, A2 => n19424, Z => n19443);
   U20085 : NOR2_X1 port map( A1 => n18662, A2 => n18678, ZN => n18450);
   U20098 : NAND2_X2 port map( A1 => n27930, A2 => n27929, ZN => n4387);
   U20138 : INV_X2 port map( I => n27936, ZN => n18884);
   U20142 : BUF_X2 port map( I => n21842, Z => n27937);
   U20155 : INV_X2 port map( I => n21429, ZN => n27939);
   U20156 : XNOR2_X1 port map( A1 => n22211, A2 => n22210, ZN => n28873);
   U20186 : XOR2_X1 port map( A1 => n27946, A2 => n6328, Z => n6820);
   U20210 : NOR2_X1 port map( A1 => n6300, A2 => n22956, ZN => n16203);
   U20243 : XOR2_X1 port map( A1 => n14733, A2 => n15923, Z => n27952);
   U20246 : OAI21_X2 port map( A1 => n18407, A2 => n9401, B => n27953, ZN => 
                           n19322);
   U20266 : NOR3_X1 port map( A1 => n11845, A2 => n24315, A3 => n13232, ZN => 
                           n12188);
   U20270 : OAI21_X1 port map( A1 => n33721, A2 => n13499, B => n17878, ZN => 
                           n14266);
   U20279 : INV_X2 port map( I => n27957, ZN => n572);
   U20292 : INV_X2 port map( I => n27960, ZN => n29268);
   U20296 : NAND2_X1 port map( A1 => n27962, A2 => n27961, ZN => n2421);
   U20300 : INV_X1 port map( I => n24675, ZN => n27962);
   U20314 : XOR2_X1 port map( A1 => n7686, A2 => n7684, Z => n17450);
   U20320 : NOR2_X1 port map( A1 => n27963, A2 => n14490, ZN => n15818);
   U20332 : OAI21_X2 port map( A1 => n15841, A2 => n33783, B => n2778, ZN => 
                           n17515);
   U20343 : XOR2_X1 port map( A1 => n27968, A2 => n24993, Z => Ciphertext(27));
   U20360 : NAND3_X1 port map( A1 => n27969, A2 => n23027, A3 => n16976, ZN => 
                           n22749);
   U20375 : NAND2_X2 port map( A1 => n27972, A2 => n11448, ZN => n13553);
   U20390 : XOR2_X1 port map( A1 => n32286, A2 => n8548, Z => n12121);
   U20404 : OR2_X1 port map( A1 => n469, A2 => n26049, Z => n4927);
   U20415 : XOR2_X1 port map( A1 => n8053, A2 => n8054, Z => n27976);
   U20435 : NOR2_X1 port map( A1 => n676, A2 => n25564, ZN => n3922);
   U20446 : XOR2_X1 port map( A1 => n304, A2 => n24560, Z => n27977);
   U20447 : NAND2_X1 port map( A1 => n23825, A2 => n14164, ZN => n13721);
   U20452 : NOR2_X1 port map( A1 => n16849, A2 => n31579, ZN => n27980);
   U20473 : NAND2_X2 port map( A1 => n8962, A2 => n8963, ZN => n10510);
   U20489 : NOR2_X2 port map( A1 => n9500, A2 => n9502, ZN => n16458);
   U20493 : INV_X4 port map( I => n12700, ZN => n12586);
   U20494 : NAND2_X1 port map( A1 => n22983, A2 => n12700, ZN => n22800);
   U20495 : NOR2_X2 port map( A1 => n27994, A2 => n27993, ZN => n12700);
   U20501 : XOR2_X1 port map( A1 => n28163, A2 => n27995, Z => n453);
   U20505 : XOR2_X1 port map( A1 => n5472, A2 => n20836, Z => n20916);
   U20510 : NOR2_X1 port map( A1 => n23842, A2 => n23887, ZN => n28016);
   U20515 : XOR2_X1 port map( A1 => n12478, A2 => n16958, Z => n8526);
   U20524 : XOR2_X1 port map( A1 => n22023, A2 => n28000, Z => n110);
   U20533 : XOR2_X1 port map( A1 => n19515, A2 => n28004, Z => n16590);
   U20539 : XOR2_X1 port map( A1 => n28908, A2 => n26000, Z => n28004);
   U20544 : BUF_X2 port map( I => n22185, Z => n28005);
   U20557 : NAND2_X2 port map( A1 => n19839, A2 => n19838, ZN => n20507);
   U20565 : INV_X2 port map( I => n28014, ZN => n28865);
   U20572 : NOR2_X1 port map( A1 => n4182, A2 => n724, ZN => n6382);
   U20576 : OAI22_X1 port map( A1 => n9438, A2 => n14156, B1 => n955, B2 => 
                           n15406, ZN => n14652);
   U20623 : XOR2_X1 port map( A1 => n18050, A2 => n28027, Z => n18049);
   U20688 : XOR2_X1 port map( A1 => n3630, A2 => n3627, Z => n18197);
   U20695 : INV_X2 port map( I => n28034, ZN => n667);
   U20704 : NAND2_X2 port map( A1 => n13284, A2 => n13283, ZN => n20519);
   U20721 : OAI21_X2 port map( A1 => n7051, A2 => n21178, B => n28038, ZN => 
                           n21581);
   U20723 : XOR2_X1 port map( A1 => n2333, A2 => n2334, Z => n28039);
   U20775 : NAND2_X1 port map( A1 => n4425, A2 => n31914, ZN => n6244);
   U20796 : OR2_X1 port map( A1 => n11072, A2 => n19315, Z => n11070);
   U20816 : OAI21_X1 port map( A1 => n18587, A2 => n18532, B => n33205, ZN => 
                           n18530);
   U20826 : XOR2_X1 port map( A1 => n28052, A2 => n25669, Z => Ciphertext(143))
                           ;
   U20830 : INV_X2 port map( I => n21454, ZN => n6493);
   U20833 : NAND2_X1 port map( A1 => n780, A2 => n27912, ZN => n11292);
   U20840 : XOR2_X1 port map( A1 => n17804, A2 => n603, Z => n21454);
   U20863 : XNOR2_X1 port map( A1 => n12609, A2 => n6789, ZN => n28086);
   U20897 : XOR2_X1 port map( A1 => n28057, A2 => n18065, Z => n16695);
   U20903 : XOR2_X1 port map( A1 => n17958, A2 => n6376, Z => n28057);
   U20915 : NOR2_X2 port map( A1 => n11596, A2 => n14864, ZN => n28059);
   U20920 : XOR2_X1 port map( A1 => n22178, A2 => n22177, Z => n22179);
   U20960 : XOR2_X1 port map( A1 => n23496, A2 => n23118, Z => n28062);
   U20986 : NAND2_X2 port map( A1 => n14539, A2 => n12004, ZN => n12329);
   U21001 : XOR2_X1 port map( A1 => n6454, A2 => n22056, Z => n22312);
   U21029 : NAND2_X1 port map( A1 => n17673, A2 => n24565, ZN => n25344);
   U21039 : INV_X4 port map( I => n17855, ZN => n10031);
   U21052 : XOR2_X1 port map( A1 => n7411, A2 => n51, Z => n28072);
   U21090 : OAI21_X1 port map( A1 => n14331, A2 => n9553, B => n19249, ZN => 
                           n8672);
   U21095 : INV_X2 port map( I => n28078, ZN => n6860);
   U21096 : XOR2_X1 port map( A1 => Plaintext(160), A2 => Key(160), Z => n28078
                           );
   U21102 : XOR2_X1 port map( A1 => n17423, A2 => n14206, Z => n20773);
   U21130 : XNOR2_X1 port map( A1 => n9517, A2 => n19516, ZN => n28174);
   U21157 : AOI22_X1 port map( A1 => n18301, A2 => n13279, B1 => n18302, B2 => 
                           n18722, ZN => n28084);
   U21189 : INV_X2 port map( I => n12895, ZN => n20099);
   U21212 : XOR2_X1 port map( A1 => n24684, A2 => n6646, Z => n28093);
   U21230 : AND2_X1 port map( A1 => n15216, A2 => n6860, Z => n18858);
   U21231 : OAI21_X1 port map( A1 => n27719, A2 => n27007, B => n17408, ZN => 
                           n22825);
   U21235 : NOR2_X1 port map( A1 => n25760, A2 => n17120, ZN => n24437);
   U21243 : INV_X2 port map( I => n18150, ZN => n28096);
   U21253 : OR2_X1 port map( A1 => n18638, A2 => n9437, Z => n9438);
   U21255 : XOR2_X1 port map( A1 => n23233, A2 => n29231, Z => n28100);
   U21262 : NAND2_X2 port map( A1 => n11086, A2 => n12966, ZN => n20426);
   U21265 : NAND3_X1 port map( A1 => n28102, A2 => n18855, A3 => n26068, ZN => 
                           n5154);
   U21269 : XOR2_X1 port map( A1 => n23358, A2 => n23306, Z => n23236);
   U21277 : XOR2_X1 port map( A1 => n16128, A2 => n8548, Z => n24382);
   U21278 : NOR2_X2 port map( A1 => n7098, A2 => n7100, ZN => n16128);
   U21294 : INV_X2 port map( I => n3535, ZN => n28104);
   U21295 : INV_X2 port map( I => n19133, ZN => n28105);
   U21300 : INV_X2 port map( I => n30281, ZN => n1207);
   U21324 : AOI22_X1 port map( A1 => n20617, A2 => n32594, B1 => n7873, B2 => 
                           n20616, ZN => n20620);
   U21328 : XOR2_X1 port map( A1 => n28109, A2 => n8596, Z => n17638);
   U21335 : AOI21_X2 port map( A1 => n21672, A2 => n21673, B => n28111, ZN => 
                           n7641);
   U21343 : INV_X1 port map( I => n28114, ZN => n28113);
   U21344 : OAI21_X1 port map( A1 => n888, A2 => n23665, B => n23382, ZN => 
                           n28114);
   U21356 : XOR2_X1 port map( A1 => n28116, A2 => n16598, Z => Ciphertext(146))
                           ;
   U21363 : XOR2_X1 port map( A1 => n23244, A2 => n530, Z => n13131);
   U21368 : XOR2_X1 port map( A1 => n28118, A2 => n23276, Z => n10659);
   U21369 : INV_X1 port map( I => n23383, ZN => n28118);
   U21388 : NAND2_X2 port map( A1 => n7376, A2 => n3104, ZN => n10720);
   U21390 : XOR2_X1 port map( A1 => n9569, A2 => n9567, Z => n28121);
   U21408 : XOR2_X1 port map( A1 => n4414, A2 => n4411, Z => n28123);
   U21412 : OR2_X1 port map( A1 => n20527, A2 => n20566, Z => n28126);
   U21414 : XNOR2_X1 port map( A1 => n16946, A2 => n16945, ZN => n28751);
   U21439 : NAND2_X2 port map( A1 => n10234, A2 => n15640, ZN => n22255);
   U21464 : XOR2_X1 port map( A1 => n20983, A2 => n11118, Z => n28134);
   U21487 : NAND2_X2 port map( A1 => n14233, A2 => n14194, ZN => n19050);
   U21505 : INV_X2 port map( I => n28142, ZN => n2967);
   U21513 : NAND2_X2 port map( A1 => n3885, A2 => n6722, ZN => n25689);
   U21527 : NAND2_X1 port map( A1 => n24921, A2 => n24933, ZN => n24348);
   U21553 : XOR2_X1 port map( A1 => n10255, A2 => n28150, Z => n15496);
   U21555 : XOR2_X1 port map( A1 => n9307, A2 => n15452, Z => n28150);
   U21556 : INV_X2 port map( I => n28151, ZN => n11621);
   U21566 : INV_X2 port map( I => n16291, ZN => n733);
   U21580 : XOR2_X1 port map( A1 => n17775, A2 => n28152, Z => n8432);
   U21581 : XOR2_X1 port map( A1 => n23286, A2 => n23297, Z => n28152);
   U21589 : NAND3_X1 port map( A1 => n12952, A2 => n8527, A3 => n9580, ZN => 
                           n22513);
   U21592 : NAND2_X1 port map( A1 => n224, A2 => n19868, ZN => n19869);
   U21593 : OR2_X1 port map( A1 => n17971, A2 => n12670, Z => n4517);
   U21602 : NOR2_X1 port map( A1 => n24874, A2 => n28520, ZN => n28519);
   U21613 : AOI21_X1 port map( A1 => n28471, A2 => n20306, B => n28316, ZN => 
                           n20162);
   U21615 : XOR2_X1 port map( A1 => n28156, A2 => n25610, Z => Ciphertext(135))
                           ;
   U21632 : NAND2_X1 port map( A1 => n18251, A2 => n21740, ZN => n28158);
   U21633 : XOR2_X1 port map( A1 => n20686, A2 => n2976, Z => n2756);
   U21634 : XOR2_X1 port map( A1 => n20766, A2 => n20921, Z => n20686);
   U21638 : NAND2_X1 port map( A1 => n11406, A2 => n10670, ZN => n6380);
   U21669 : XOR2_X1 port map( A1 => n3739, A2 => n27171, Z => n13702);
   U21680 : NAND2_X2 port map( A1 => n7462, A2 => n882, ZN => n9555);
   U21682 : NAND2_X2 port map( A1 => n9805, A2 => n9363, ZN => n25765);
   U21683 : NAND2_X2 port map( A1 => n25701, A2 => n25703, ZN => n9363);
   U21684 : BUF_X2 port map( I => n22428, Z => n28170);
   U21691 : NAND2_X2 port map( A1 => n4472, A2 => n28172, ZN => n4016);
   U21698 : XOR2_X1 port map( A1 => n22023, A2 => n1992, Z => n1991);
   U21700 : NAND2_X1 port map( A1 => n17624, A2 => n21341, ZN => n10468);
   U21703 : OAI22_X2 port map( A1 => n5978, A2 => n21076, B1 => n9842, B2 => 
                           n21243, ZN => n5830);
   U21709 : XOR2_X1 port map( A1 => n28174, A2 => n12803, Z => n562);
   U21731 : XOR2_X1 port map( A1 => n20825, A2 => n25910, Z => n16775);
   U21732 : NAND2_X2 port map( A1 => n20233, A2 => n285, ZN => n20825);
   U21762 : XOR2_X1 port map( A1 => n28179, A2 => n10507, Z => n10505);
   U21776 : NOR2_X2 port map( A1 => n23749, A2 => n23757, ZN => n8330);
   U21780 : XOR2_X1 port map( A1 => n22229, A2 => n16971, Z => n5196);
   U21833 : XOR2_X1 port map( A1 => n24761, A2 => n1225, Z => n28188);
   U21853 : NAND2_X1 port map( A1 => n9858, A2 => n837, ZN => n11046);
   U21868 : NOR2_X2 port map( A1 => n18997, A2 => n18996, ZN => n28197);
   U21869 : NAND2_X2 port map( A1 => n3915, A2 => n20097, ZN => n19878);
   U21886 : XOR2_X1 port map( A1 => n5148, A2 => n16841, Z => n12750);
   U21889 : NAND2_X1 port map( A1 => n30937, A2 => n29102, ZN => n3091);
   U21945 : NAND2_X1 port map( A1 => n14795, A2 => n25215, ZN => n25217);
   U21950 : XOR2_X1 port map( A1 => n17126, A2 => n17125, Z => n17127);
   U21958 : OR2_X1 port map( A1 => n295, A2 => n16144, Z => n2622);
   U21964 : XOR2_X1 port map( A1 => n28216, A2 => n19492, Z => n6693);
   U21995 : NOR2_X2 port map( A1 => n10397, A2 => n8543, ZN => n10511);
   U21997 : OAI21_X2 port map( A1 => n9242, A2 => n32037, B => n32858, ZN => 
                           n9243);
   U22000 : INV_X1 port map( I => n5713, ZN => n28228);
   U22014 : XNOR2_X1 port map( A1 => n17400, A2 => n23519, ZN => n29194);
   U22015 : INV_X4 port map( I => n701, ZN => n28473);
   U22022 : AOI21_X2 port map( A1 => n11078, A2 => n977, B => n11077, ZN => 
                           n28235);
   U22030 : OAI21_X1 port map( A1 => n3915, A2 => n27832, B => n30692, ZN => 
                           n8549);
   U22034 : XOR2_X1 port map( A1 => n32052, A2 => n21028, Z => n2976);
   U22041 : INV_X2 port map( I => n28236, ZN => n9678);
   U22057 : NAND2_X2 port map( A1 => n17907, A2 => n12116, ZN => n19252);
   U22080 : BUF_X2 port map( I => n9342, Z => n28240);
   U22090 : OR2_X1 port map( A1 => n25470, A2 => n25476, Z => n28243);
   U22098 : XNOR2_X1 port map( A1 => Plaintext(146), A2 => Key(146), ZN => 
                           n28245);
   U22118 : NAND2_X2 port map( A1 => n10387, A2 => n10386, ZN => n28697);
   U22130 : XOR2_X1 port map( A1 => n19574, A2 => n16792, Z => n13780);
   U22134 : XOR2_X1 port map( A1 => n28251, A2 => n16698, Z => Ciphertext(141))
                           ;
   U22139 : NAND3_X1 port map( A1 => n28252, A2 => n15185, A3 => n15295, ZN => 
                           n15184);
   U22144 : INV_X1 port map( I => n12235, ZN => n28252);
   U22151 : OAI21_X2 port map( A1 => n23752, A2 => n7895, B => n31984, ZN => 
                           n6716);
   U22156 : BUF_X2 port map( I => n24755, Z => n28258);
   U22195 : INV_X2 port map( I => n15092, ZN => n28266);
   U22206 : NOR2_X1 port map( A1 => n25093, A2 => n32857, ZN => n28270);
   U22213 : XOR2_X1 port map( A1 => n21044, A2 => n16322, Z => n7138);
   U22227 : XOR2_X1 port map( A1 => n23337, A2 => n23338, Z => n14103);
   U22243 : NAND2_X2 port map( A1 => n10481, A2 => n10485, ZN => n14597);
   U22263 : NAND2_X2 port map( A1 => n16050, A2 => n34108, ZN => n2535);
   U22268 : NAND2_X1 port map( A1 => n27188, A2 => n28096, ZN => n28283);
   U22278 : AND2_X1 port map( A1 => n19451, A2 => n4180, Z => n3593);
   U22279 : NAND2_X2 port map( A1 => n7952, A2 => n7951, ZN => n20959);
   U22311 : BUF_X2 port map( I => n10001, Z => n28288);
   U22321 : XOR2_X1 port map( A1 => n28289, A2 => n12957, Z => n4021);
   U22322 : NAND2_X2 port map( A1 => n20275, A2 => n20274, ZN => n12957);
   U22342 : XOR2_X1 port map( A1 => n31043, A2 => n31966, Z => n8827);
   U22357 : NAND2_X1 port map( A1 => n19224, A2 => n5610, ZN => n4366);
   U22387 : AND2_X1 port map( A1 => n6474, A2 => n23872, Z => n9813);
   U22388 : AOI21_X1 port map( A1 => n6097, A2 => n25475, B => n28302, ZN => 
                           n6095);
   U22397 : OR2_X1 port map( A1 => n17151, A2 => n32082, Z => n29021);
   U22401 : NAND2_X2 port map( A1 => n17404, A2 => n32917, ZN => n24039);
   U22417 : OAI21_X2 port map( A1 => n8841, A2 => n8840, B => n28304, ZN => 
                           n5578);
   U22433 : OAI21_X2 port map( A1 => n5163, A2 => n1249, B => n9736, ZN => 
                           n28307);
   U22437 : OAI21_X2 port map( A1 => n933, A2 => n1636, B => n15213, ZN => 
                           n28309);
   U22450 : XOR2_X1 port map( A1 => n23290, A2 => n28311, Z => n29203);
   U22453 : XOR2_X1 port map( A1 => n14242, A2 => n23289, Z => n28311);
   U22460 : AOI21_X2 port map( A1 => n5851, A2 => n31102, B => n5849, ZN => 
                           n5848);
   U22467 : INV_X2 port map( I => n28312, ZN => n635);
   U22482 : OR2_X1 port map( A1 => n8457, A2 => n13652, Z => n12725);
   U22531 : NOR2_X1 port map( A1 => n11454, A2 => n2387, ZN => n28451);
   U22538 : XOR2_X1 port map( A1 => n29876, A2 => n16685, Z => n462);
   U22553 : XOR2_X1 port map( A1 => Plaintext(12), A2 => Key(12), Z => n28321);
   U22555 : AND2_X1 port map( A1 => n5191, A2 => n13413, Z => n23758);
   U22585 : NAND2_X1 port map( A1 => n25666, A2 => n25650, ZN => n25643);
   U22588 : NAND2_X2 port map( A1 => n25640, A2 => n15184, ZN => n25666);
   U22593 : XOR2_X1 port map( A1 => n28331, A2 => n16464, Z => Ciphertext(186))
                           ;
   U22600 : OR2_X1 port map( A1 => n9831, A2 => n14980, Z => n9833);
   U22603 : NAND2_X2 port map( A1 => n17405, A2 => n32745, ZN => n19820);
   U22614 : NAND2_X2 port map( A1 => n28332, A2 => n13865, ZN => n13864);
   U22637 : NAND2_X2 port map( A1 => n12586, A2 => n28697, ZN => n15364);
   U22640 : NAND2_X2 port map( A1 => n15696, A2 => n18074, ZN => n7680);
   U22641 : NOR2_X2 port map( A1 => n7726, A2 => n28796, ZN => n15696);
   U22654 : XOR2_X1 port map( A1 => n528, A2 => n23205, Z => n6294);
   U22660 : NAND2_X2 port map( A1 => n12863, A2 => n28686, ZN => n9667);
   U22662 : XOR2_X1 port map( A1 => n28903, A2 => n3635, Z => n2163);
   U22668 : NAND2_X2 port map( A1 => n4508, A2 => n4507, ZN => n28885);
   U22670 : NOR2_X1 port map( A1 => n19822, A2 => n9619, ZN => n28856);
   U22671 : NOR2_X1 port map( A1 => n18650, A2 => n18373, ZN => n16196);
   U22707 : NAND3_X1 port map( A1 => n1247, A2 => n27136, A3 => n23860, ZN => 
                           n5685);
   U22719 : XOR2_X1 port map( A1 => n9274, A2 => n5558, Z => n28354);
   U22720 : OR2_X1 port map( A1 => n7305, A2 => n15359, Z => n5621);
   U22727 : XOR2_X1 port map( A1 => n10865, A2 => n26003, Z => n10863);
   U22735 : XOR2_X1 port map( A1 => n20987, A2 => n20988, Z => n2820);
   U22759 : OR2_X1 port map( A1 => n22674, A2 => n10568, Z => n13105);
   U22773 : NOR2_X1 port map( A1 => n23847, A2 => n26114, ZN => n17980);
   U22775 : OAI21_X1 port map( A1 => n18775, A2 => n18556, B => n29074, ZN => 
                           n29073);
   U22779 : NAND3_X1 port map( A1 => n20014, A2 => n20013, A3 => n5267, ZN => 
                           n28366);
   U22792 : OR2_X1 port map( A1 => n627, A2 => n5379, Z => n2793);
   U22853 : INV_X2 port map( I => n28373, ZN => n1926);
   U22871 : NAND2_X2 port map( A1 => n11464, A2 => n20222, ZN => n20729);
   U22872 : NAND2_X2 port map( A1 => n16785, A2 => n21267, ZN => n21265);
   U22879 : OAI22_X2 port map( A1 => n1534, A2 => n21748, B1 => n1532, B2 => 
                           n1533, ZN => n22211);
   U22880 : XOR2_X1 port map( A1 => n28399, A2 => n16322, Z => n28859);
   U22902 : AND2_X1 port map( A1 => n2964, A2 => n2107, Z => n28381);
   U22905 : NOR2_X1 port map( A1 => n28383, A2 => n2107, ZN => n28382);
   U22950 : AOI21_X2 port map( A1 => n9686, A2 => n28838, B => n28393, ZN => 
                           n9691);
   U22975 : NAND2_X2 port map( A1 => n28397, A2 => n3794, ZN => n8515);
   U22976 : NAND2_X1 port map( A1 => n9957, A2 => n9402, ZN => n28397);
   U22978 : BUF_X2 port map( I => n19197, Z => n28399);
   U22986 : OAI21_X2 port map( A1 => n3797, A2 => n3796, B => n5997, ZN => 
                           n22005);
   U23013 : OAI22_X2 port map( A1 => n25767, A2 => n25766, B1 => n25764, B2 => 
                           n25765, ZN => n25795);
   U23019 : OR2_X1 port map( A1 => n14780, A2 => n29243, Z => n11518);
   U23043 : OAI22_X1 port map( A1 => n25207, A2 => n5173, B1 => n5043, B2 => 
                           n715, ZN => n5172);
   U23045 : INV_X2 port map( I => n28407, ZN => n29269);
   U23055 : INV_X2 port map( I => n9625, ZN => n28410);
   U23101 : XOR2_X1 port map( A1 => n22206, A2 => n28416, Z => n29162);
   U23103 : XOR2_X1 port map( A1 => n1308, A2 => n22205, Z => n28416);
   U23118 : NOR2_X1 port map( A1 => n3663, A2 => n12408, ZN => n28418);
   U23122 : AOI21_X2 port map( A1 => n12232, A2 => n12110, B => n28420, ZN => 
                           n206);
   U23125 : XOR2_X1 port map( A1 => n19522, A2 => n28421, Z => n12057);
   U23126 : XOR2_X1 port map( A1 => n28601, A2 => n28422, Z => n28421);
   U23129 : NOR2_X2 port map( A1 => n28426, A2 => n28425, ZN => n263);
   U23140 : XOR2_X1 port map( A1 => n22288, A2 => n22289, Z => n9911);
   U23143 : INV_X2 port map( I => n28430, ZN => n20080);
   U23155 : NAND3_X2 port map( A1 => n28437, A2 => n13867, A3 => n29676, ZN => 
                           n13865);
   U23160 : NAND3_X1 port map( A1 => n28438, A2 => n18855, A3 => n8411, ZN => 
                           n8554);
   U23170 : XNOR2_X1 port map( A1 => n22048, A2 => n22148, ZN => n21931);
   U23172 : XOR2_X1 port map( A1 => n9000, A2 => n1128, Z => n28441);
   U23187 : NAND2_X1 port map( A1 => n13426, A2 => n19021, ZN => n19022);
   U23188 : NAND2_X1 port map( A1 => n8227, A2 => n17817, ZN => n28442);
   U23195 : XOR2_X1 port map( A1 => n19579, A2 => n19480, Z => n17300);
   U23197 : XOR2_X1 port map( A1 => n28443, A2 => n5663, Z => n17214);
   U23216 : NAND2_X2 port map( A1 => n28444, A2 => n18452, ZN => n19764);
   U23239 : XOR2_X1 port map( A1 => n7160, A2 => n11476, Z => n28446);
   U23248 : NAND2_X1 port map( A1 => n28447, A2 => n18973, ZN => n16725);
   U23255 : XOR2_X1 port map( A1 => n9154, A2 => n6294, Z => n9152);
   U23261 : XOR2_X1 port map( A1 => n12422, A2 => n13496, Z => n28448);
   U23263 : NOR2_X1 port map( A1 => n18088, A2 => n15753, ZN => n28449);
   U23302 : XOR2_X1 port map( A1 => n15527, A2 => n28458, Z => n28457);
   U23312 : BUF_X2 port map( I => n23318, Z => n28460);
   U23317 : XOR2_X1 port map( A1 => n20639, A2 => n28461, Z => n16820);
   U23325 : XOR2_X1 port map( A1 => n29241, A2 => n28462, Z => n28461);
   U23334 : XOR2_X1 port map( A1 => n24455, A2 => n24454, Z => n24456);
   U23335 : XOR2_X1 port map( A1 => n8703, A2 => n14727, Z => n24454);
   U23337 : XOR2_X1 port map( A1 => n2483, A2 => n25993, Z => n15485);
   U23345 : NAND2_X2 port map( A1 => n14734, A2 => n28466, ZN => n19298);
   U23346 : OR2_X1 port map( A1 => n19296, A2 => n19297, Z => n28466);
   U23350 : XOR2_X1 port map( A1 => n27165, A2 => n12539, Z => n10582);
   U23353 : INV_X1 port map( I => n8519, ZN => n22553);
   U23357 : NAND2_X1 port map( A1 => n11451, A2 => n34161, ZN => n8519);
   U23373 : NAND2_X1 port map( A1 => n16627, A2 => n32532, ZN => n10244);
   U23381 : OR2_X1 port map( A1 => n701, A2 => n32532, Z => n22572);
   U23390 : NAND2_X1 port map( A1 => n25357, A2 => n25367, ZN => n28469);
   U23393 : NAND2_X1 port map( A1 => n25356, A2 => n30400, ZN => n28470);
   U23397 : XOR2_X1 port map( A1 => n19711, A2 => n7530, Z => n15527);
   U23400 : NAND2_X2 port map( A1 => n4914, A2 => n19059, ZN => n7530);
   U23401 : XOR2_X1 port map( A1 => n8715, A2 => n12212, Z => n8714);
   U23404 : NAND2_X2 port map( A1 => n5633, A2 => n5634, ZN => n16052);
   U23406 : NAND2_X2 port map( A1 => n28475, A2 => n28474, ZN => n22848);
   U23412 : OR2_X1 port map( A1 => n11737, A2 => n34125, Z => n28474);
   U23414 : NOR2_X2 port map( A1 => n22026, A2 => n3186, ZN => n28475);
   U23423 : NOR2_X2 port map( A1 => n23976, A2 => n23971, ZN => n888);
   U23430 : NAND2_X2 port map( A1 => n5371, A2 => n375, ZN => n6704);
   U23432 : XOR2_X1 port map( A1 => n7530, A2 => n16464, Z => n28479);
   U23438 : INV_X2 port map( I => n28480, ZN => n497);
   U23442 : XOR2_X1 port map( A1 => Plaintext(138), A2 => Key(138), Z => n28480
                           );
   U23444 : NOR2_X1 port map( A1 => n824, A2 => n9677, ZN => n12128);
   U23447 : NAND2_X2 port map( A1 => n16357, A2 => n18636, ZN => n19167);
   U23453 : XOR2_X1 port map( A1 => n24551, A2 => n6050, Z => n6054);
   U23467 : NAND2_X2 port map( A1 => n8203, A2 => n18534, ZN => n19285);
   U23476 : XOR2_X1 port map( A1 => n28482, A2 => n12185, Z => n14031);
   U23479 : XOR2_X1 port map( A1 => n23451, A2 => n13497, Z => n28482);
   U23480 : AOI21_X2 port map( A1 => n6482, A2 => n7090, B => n28483, ZN => 
                           n6835);
   U23483 : NOR2_X1 port map( A1 => n1284, A2 => n7090, ZN => n28483);
   U23493 : AOI21_X2 port map( A1 => n14696, A2 => n1709, B => n14694, ZN => 
                           n19006);
   U23496 : XOR2_X1 port map( A1 => n28486, A2 => n16911, Z => Ciphertext(41));
   U23510 : XOR2_X1 port map( A1 => n8691, A2 => n24412, Z => n11973);
   U23525 : NAND2_X1 port map( A1 => n5172, A2 => n5174, ZN => n17933);
   U23527 : AOI21_X2 port map( A1 => n11712, A2 => n10848, B => n8869, ZN => 
                           n9803);
   U23537 : NOR2_X2 port map( A1 => n25650, A2 => n25666, ZN => n9365);
   U23538 : OAI21_X1 port map( A1 => n22338, A2 => n16166, B => n22337, ZN => 
                           n22339);
   U23540 : INV_X2 port map( I => n28496, ZN => n561);
   U23547 : NAND2_X1 port map( A1 => n23833, A2 => n30252, ZN => n28497);
   U23558 : OAI22_X1 port map( A1 => n5043, A2 => n25216, B1 => n15359, B2 => 
                           n15462, ZN => n5577);
   U23582 : AOI22_X2 port map( A1 => n13238, A2 => n15376, B1 => n13237, B2 => 
                           n13459, ZN => n13236);
   U23583 : XNOR2_X1 port map( A1 => n23464, A2 => n23463, ZN => n287);
   U23592 : NAND2_X1 port map( A1 => n5438, A2 => n23655, ZN => n28503);
   U23593 : XOR2_X1 port map( A1 => n3781, A2 => n542, Z => n17703);
   U23610 : XOR2_X1 port map( A1 => n8795, A2 => n27174, Z => n28513);
   U23611 : INV_X2 port map( I => n28514, ZN => n11985);
   U23621 : NAND2_X2 port map( A1 => n13409, A2 => n13249, ZN => n22470);
   U23635 : XOR2_X1 port map( A1 => n19598, A2 => n2982, Z => n2981);
   U23654 : OAI21_X2 port map( A1 => n29123, A2 => n28525, B => n28524, ZN => 
                           n24789);
   U23656 : NAND2_X2 port map( A1 => n1869, A2 => n1870, ZN => n2483);
   U23662 : XOR2_X1 port map( A1 => n31499, A2 => n23180, Z => n23377);
   U23673 : AOI21_X2 port map( A1 => n3482, A2 => n3481, B => n28534, ZN => 
                           n3483);
   U23678 : NAND2_X2 port map( A1 => n1751, A2 => n28536, ZN => n6288);
   U23679 : NAND2_X1 port map( A1 => n25636, A2 => n24446, ZN => n28536);
   U23682 : NAND2_X2 port map( A1 => n22664, A2 => n22578, ZN => n5452);
   U23700 : NAND3_X1 port map( A1 => n28781, A2 => n4151, A3 => n28779, ZN => 
                           n3213);
   U23719 : INV_X2 port map( I => n562, ZN => n1169);
   U23720 : INV_X2 port map( I => n7677, ZN => n19474);
   U23722 : NAND2_X2 port map( A1 => n28540, A2 => n28539, ZN => n7677);
   U23730 : OAI21_X2 port map( A1 => n10259, A2 => n17981, B => n14113, ZN => 
                           n13826);
   U23732 : XOR2_X1 port map( A1 => n6624, A2 => n28542, Z => n17662);
   U23738 : XOR2_X1 port map( A1 => n19757, A2 => n18105, Z => n28542);
   U23755 : INV_X2 port map( I => n28545, ZN => n22606);
   U23774 : XOR2_X1 port map( A1 => n23335, A2 => n11891, Z => n23400);
   U23778 : OAI22_X2 port map( A1 => n5458, A2 => n5457, B1 => n18311, B2 => 
                           n5459, ZN => n10260);
   U23781 : XOR2_X1 port map( A1 => n21992, A2 => n30628, Z => n21891);
   U23799 : XOR2_X1 port map( A1 => n4601, A2 => Key(16), Z => n29061);
   U23801 : OAI22_X2 port map( A1 => n844, A2 => n23867, B1 => n33345, B2 => 
                           n11821, ZN => n1506);
   U23805 : XOR2_X1 port map( A1 => n23286, A2 => n24907, Z => n28552);
   U23810 : INV_X2 port map( I => n28554, ZN => n9953);
   U23834 : INV_X2 port map( I => n28560, ZN => n16528);
   U23840 : XOR2_X1 port map( A1 => n17097, A2 => n17094, Z => n28560);
   U23846 : NAND2_X1 port map( A1 => n32911, A2 => n5202, ZN => n7678);
   U23849 : XOR2_X1 port map( A1 => n17377, A2 => n14755, Z => n14753);
   U23854 : XOR2_X1 port map( A1 => n19662, A2 => n19663, Z => n19664);
   U23858 : NAND2_X1 port map( A1 => n16280, A2 => n3668, ZN => n3669);
   U23863 : NAND2_X1 port map( A1 => n24705, A2 => n16650, ZN => n28564);
   U23864 : OR2_X1 port map( A1 => n13194, A2 => n21313, Z => n28565);
   U23868 : XOR2_X1 port map( A1 => n28566, A2 => n17452, Z => n28979);
   U23880 : XOR2_X1 port map( A1 => n3041, A2 => n26097, Z => n28566);
   U23910 : NAND2_X2 port map( A1 => n3336, A2 => n3334, ZN => n24741);
   U23927 : OAI21_X2 port map( A1 => n1594, A2 => n857, B => n1001, ZN => 
                           n28567);
   U23936 : XOR2_X1 port map( A1 => n8921, A2 => n28571, Z => n2759);
   U23937 : XOR2_X1 port map( A1 => n3568, A2 => n2761, Z => n28571);
   U23958 : INV_X1 port map( I => n23191, ZN => n28575);
   U23990 : XOR2_X1 port map( A1 => n8680, A2 => n17119, Z => n22625);
   U23997 : XOR2_X1 port map( A1 => n32124, A2 => n18100, Z => n17141);
   U24030 : NOR2_X1 port map( A1 => n443, A2 => n30139, ZN => n442);
   U24034 : NAND2_X2 port map( A1 => n11957, A2 => n25710, ZN => n24712);
   U24040 : NOR2_X2 port map( A1 => n28586, A2 => n29221, ZN => n16309);
   U24051 : XNOR2_X1 port map( A1 => n9517, A2 => n7676, ZN => n29007);
   U24053 : XOR2_X1 port map( A1 => Plaintext(7), A2 => Key(7), Z => n8386);
   U24064 : NOR2_X1 port map( A1 => n4040, A2 => n14903, ZN => n4906);
   U24067 : INV_X2 port map( I => n28589, ZN => n639);
   U24071 : XOR2_X1 port map( A1 => n27145, A2 => n24836, Z => n12943);
   U24090 : XOR2_X1 port map( A1 => n19729, A2 => n28593, Z => n17192);
   U24091 : XOR2_X1 port map( A1 => n4400, A2 => n16581, Z => n28593);
   U24102 : XNOR2_X1 port map( A1 => n20707, A2 => n20708, ZN => n28594);
   U24106 : INV_X2 port map( I => n8088, ZN => n1333);
   U24107 : XOR2_X1 port map( A1 => n9815, A2 => n28595, Z => n8088);
   U24130 : OR2_X1 port map( A1 => n21490, A2 => n423, Z => n6146);
   U24139 : NAND2_X2 port map( A1 => n28602, A2 => n3378, ZN => n7940);
   U24146 : OAI21_X1 port map( A1 => n9252, A2 => n1158, B => n28603, ZN => 
                           n20617);
   U24148 : INV_X2 port map( I => n28605, ZN => n21403);
   U24160 : XOR2_X1 port map( A1 => n1306, A2 => n27185, Z => n28606);
   U24204 : OAI21_X2 port map( A1 => n5590, A2 => n12793, B => n5588, ZN => 
                           n20924);
   U24212 : INV_X2 port map( I => n28607, ZN => n21392);
   U24233 : INV_X2 port map( I => n28608, ZN => n651);
   U24285 : XOR2_X1 port map( A1 => n16242, A2 => n15795, Z => n28612);
   U24296 : OAI21_X2 port map( A1 => n4398, A2 => n14187, B => n8794, ZN => 
                           n8795);
   U24322 : XOR2_X1 port map( A1 => n24808, A2 => n553, Z => n2809);
   U24327 : AND2_X1 port map( A1 => n15021, A2 => n19088, Z => n28614);
   U24331 : OR2_X1 port map( A1 => n32883, A2 => n29215, Z => n21423);
   U24339 : INV_X2 port map( I => n28617, ZN => n12074);
   U24340 : XOR2_X1 port map( A1 => Plaintext(58), A2 => Key(58), Z => n28617);
   U24381 : NOR2_X1 port map( A1 => n7004, A2 => n13558, ZN => n7003);
   U24401 : NAND2_X1 port map( A1 => n14745, A2 => n16799, ZN => n28623);
   U24405 : INV_X2 port map( I => n28624, ZN => n14339);
   U24408 : XOR2_X1 port map( A1 => n6615, A2 => n28627, Z => n8228);
   U24409 : XOR2_X1 port map( A1 => n6614, A2 => n20744, Z => n28627);
   U24423 : XOR2_X1 port map( A1 => n4161, A2 => n618, Z => n28633);
   U24441 : XOR2_X1 port map( A1 => Plaintext(106), A2 => Key(106), Z => n13445
                           );
   U24461 : XOR2_X1 port map( A1 => n28636, A2 => n2045, Z => n10255);
   U24464 : XOR2_X1 port map( A1 => n10257, A2 => n24807, Z => n28636);
   U24546 : BUF_X2 port map( I => n8398, Z => n28641);
   U24566 : XOR2_X1 port map( A1 => n13419, A2 => n24553, Z => n24626);
   U24593 : INV_X2 port map( I => n15324, ZN => n28649);
   U24632 : NAND2_X1 port map( A1 => n28658, A2 => n25072, ZN => n28657);
   U24648 : XOR2_X1 port map( A1 => n23388, A2 => n27171, Z => n23255);
   U24649 : XOR2_X1 port map( A1 => n20788, A2 => n3705, Z => n6088);
   U24664 : NAND2_X2 port map( A1 => n10048, A2 => n18120, ZN => n24799);
   U24694 : XOR2_X1 port map( A1 => n2698, A2 => n2699, Z => n28663);
   U24698 : NAND2_X2 port map( A1 => n974, A2 => n10281, ZN => n6319);
   U24734 : NAND2_X2 port map( A1 => n33731, A2 => n1133, ZN => n7502);
   U24740 : INV_X1 port map( I => n17167, ZN => n28964);
   U24771 : XOR2_X1 port map( A1 => n28673, A2 => n3599, Z => n5324);
   U24773 : XOR2_X1 port map( A1 => n19408, A2 => n16520, Z => n28673);
   U24774 : AOI22_X1 port map( A1 => n5543, A2 => n17273, B1 => n7928, B2 => 
                           n25247, ZN => n4226);
   U24782 : NOR2_X1 port map( A1 => n19183, A2 => n19105, ZN => n15291);
   U24785 : NAND2_X2 port map( A1 => n28674, A2 => n18905, ZN => n16349);
   U24807 : XOR2_X1 port map( A1 => n7630, A2 => n26028, Z => n15669);
   U24852 : XOR2_X1 port map( A1 => n1085, A2 => n24689, Z => n5358);
   U24867 : NOR3_X2 port map( A1 => n29211, A2 => n26093, A3 => n13489, ZN => 
                           n20518);
   U24886 : NOR2_X2 port map( A1 => n28696, A2 => n11769, ZN => n14161);
   U24891 : OAI21_X2 port map( A1 => n8037, A2 => n8038, B => n12702, ZN => 
                           n13844);
   U24897 : NAND2_X2 port map( A1 => n28698, A2 => n1730, ZN => n6286);
   U24907 : XOR2_X1 port map( A1 => n5925, A2 => n26029, Z => n7374);
   U24915 : AND2_X1 port map( A1 => n9953, A2 => n639, Z => n15464);
   U24940 : XOR2_X1 port map( A1 => n15787, A2 => n15786, Z => n15788);
   U24992 : OR2_X1 port map( A1 => n11006, A2 => n19936, Z => n28852);
   U24999 : XOR2_X1 port map( A1 => n28708, A2 => n4158, Z => n14676);
   U25000 : XOR2_X1 port map( A1 => n22187, A2 => n15900, Z => n28708);
   U25001 : NAND2_X2 port map( A1 => n12599, A2 => n12598, ZN => n15230);
   U25015 : XOR2_X1 port map( A1 => n253, A2 => n28711, Z => n28710);
   U25028 : NAND3_X2 port map( A1 => n607, A2 => n28712, A3 => n10671, ZN => 
                           n11562);
   U25053 : XOR2_X1 port map( A1 => n10331, A2 => n24755, Z => n8109);
   U25067 : NAND2_X2 port map( A1 => n15058, A2 => n2270, ZN => n25006);
   U25078 : NAND2_X2 port map( A1 => n18910, A2 => n18909, ZN => n14120);
   U25083 : OAI21_X2 port map( A1 => n15486, A2 => n17311, B => n17819, ZN => 
                           n19599);
   U25117 : INV_X2 port map( I => n28723, ZN => n676);
   U25145 : XOR2_X1 port map( A1 => n2012, A2 => n2013, Z => n28723);
   U25147 : NAND2_X1 port map( A1 => n25664, A2 => n25650, ZN => n7087);
   U25148 : XOR2_X1 port map( A1 => n17219, A2 => n28724, Z => n11806);
   U25162 : XOR2_X1 port map( A1 => n1310, A2 => n6435, Z => n28724);
   U25203 : NAND3_X1 port map( A1 => n19597, A2 => n18668, A3 => n18669, ZN => 
                           n8716);
   U25209 : INV_X2 port map( I => n28731, ZN => n13360);
   U25213 : XOR2_X1 port map( A1 => Plaintext(147), A2 => Key(147), Z => n28731
                           );
   U25261 : AOI22_X2 port map( A1 => n2709, A2 => n4359, B1 => n2710, B2 => 
                           n21823, ZN => n22196);
   U25264 : XOR2_X1 port map( A1 => n28735, A2 => n25311, Z => Ciphertext(90));
   U25300 : XOR2_X1 port map( A1 => n14000, A2 => n24686, Z => n24783);
   U25305 : NOR2_X2 port map( A1 => n3256, A2 => n3257, ZN => n14000);
   U25356 : XOR2_X1 port map( A1 => n20787, A2 => n7113, Z => n28748);
   U25375 : INV_X2 port map( I => n28750, ZN => n25014);
   U25377 : AOI22_X2 port map( A1 => n18577, A2 => n3779, B1 => n14453, B2 => 
                           n18387, ZN => n7995);
   U25387 : XOR2_X1 port map( A1 => n9193, A2 => n28751, Z => n22414);
   U25423 : XOR2_X1 port map( A1 => n29190, A2 => n29206, Z => n28753);
   U25430 : OR2_X2 port map( A1 => n8251, A2 => n2450, Z => n23885);
   U25452 : OAI22_X2 port map( A1 => n28755, A2 => n8271, B1 => n414, B2 => 
                           n9651, ZN => n7233);
   U25454 : OAI21_X2 port map( A1 => n1059, A2 => n5834, B => n1659, ZN => 
                           n28755);
   U25494 : XNOR2_X1 port map( A1 => n19193, A2 => n11450, ZN => n29079);
   U25497 : INV_X2 port map( I => n10937, ZN => n14756);
   U25528 : INV_X2 port map( I => n28763, ZN => n8105);
   U25535 : XOR2_X1 port map( A1 => n16737, A2 => n16739, Z => n28763);
   U25570 : XOR2_X1 port map( A1 => n19495, A2 => n28769, Z => n11321);
   U25574 : XOR2_X1 port map( A1 => n19637, A2 => n28908, Z => n28769);
   U25586 : NAND2_X2 port map( A1 => n28770, A2 => n14100, ZN => n18626);
   U25595 : XOR2_X1 port map( A1 => n28771, A2 => n19551, Z => n3074);
   U25604 : XOR2_X1 port map( A1 => n1370, A2 => n3076, Z => n28771);
   U25643 : NAND2_X1 port map( A1 => n24283, A2 => n26387, ZN => n28779);
   U25654 : NOR2_X1 port map( A1 => n22577, A2 => n28635, ZN => n14220);
   U25659 : OAI21_X1 port map( A1 => n1200, A2 => n24934, B => n24933, ZN => 
                           n7787);
   U25660 : NAND2_X2 port map( A1 => n8778, A2 => n14001, ZN => n24919);
   U25662 : XOR2_X1 port map( A1 => n20733, A2 => n20891, Z => n20765);
   U25668 : XOR2_X1 port map( A1 => n12442, A2 => n15978, Z => n19666);
   U25670 : NAND2_X2 port map( A1 => n11777, A2 => n11778, ZN => n12442);
   U25675 : INV_X1 port map( I => n24283, ZN => n24040);
   U25687 : XNOR2_X1 port map( A1 => n22182, A2 => n22181, ZN => n29170);
   U25708 : XOR2_X1 port map( A1 => n28788, A2 => n4000, Z => n8190);
   U25710 : XOR2_X1 port map( A1 => n20758, A2 => n29832, Z => n28788);
   U25712 : OAI21_X2 port map( A1 => n18486, A2 => n14284, B => n18768, ZN => 
                           n28789);
   U25713 : NAND2_X2 port map( A1 => n7708, A2 => n7709, ZN => n7705);
   U25715 : OAI21_X1 port map( A1 => n32856, A2 => n9982, B => n28791, ZN => 
                           n25605);
   U25718 : AOI21_X1 port map( A1 => n1034, A2 => n27177, B => n9320, ZN => 
                           n5219);
   U25724 : OR2_X1 port map( A1 => n14331, A2 => n15050, Z => n259);
   U25727 : NAND2_X1 port map( A1 => n12195, A2 => n6213, ZN => n6212);
   U25729 : NAND2_X1 port map( A1 => n16785, A2 => n8490, ZN => n12195);
   U25730 : XOR2_X1 port map( A1 => n20806, A2 => n13590, Z => n13456);
   U25743 : NOR2_X1 port map( A1 => n7898, A2 => n9766, ZN => n28796);
   U25760 : NAND2_X1 port map( A1 => n7213, A2 => n7212, ZN => n28797);
   U25761 : INV_X2 port map( I => n9240, ZN => n25621);
   U25773 : XOR2_X1 port map( A1 => n8522, A2 => n17833, Z => n9240);
   U25786 : OR2_X1 port map( A1 => n20605, A2 => n7892, Z => n28799);
   U25790 : NAND2_X1 port map( A1 => n28800, A2 => n28580, ZN => n4123);
   U25791 : NOR2_X1 port map( A1 => n12535, A2 => n10720, ZN => n28800);
   U25798 : OAI21_X1 port map( A1 => n16193, A2 => n16493, B => n16105, ZN => 
                           n11502);
   U25799 : NAND2_X2 port map( A1 => n22773, A2 => n9075, ZN => n11891);
   U25803 : XOR2_X1 port map( A1 => n19629, A2 => n15978, Z => n19441);
   U25806 : XOR2_X1 port map( A1 => n8635, A2 => n16319, Z => n28807);
   U25813 : NAND2_X2 port map( A1 => n18514, A2 => n14393, ZN => n19178);
   U25816 : XOR2_X1 port map( A1 => n3190, A2 => n3191, Z => n3192);
   U25817 : XOR2_X1 port map( A1 => n20767, A2 => n21046, Z => n28814);
   U25821 : INV_X2 port map( I => n28816, ZN => n680);
   U25822 : XOR2_X1 port map( A1 => n28817, A2 => n23522, Z => n2972);
   U25823 : XOR2_X1 port map( A1 => n9843, A2 => n2974, Z => n28817);
   U25824 : AND2_X1 port map( A1 => n29207, A2 => n11966, Z => n4423);
   U25826 : NAND3_X1 port map( A1 => n24069, A2 => n1092, A3 => n25973, ZN => 
                           n3021);
   U25827 : XOR2_X1 port map( A1 => n28818, A2 => n2190, Z => n4338);
   U25828 : NAND2_X1 port map( A1 => n12291, A2 => n12290, ZN => n10127);
   U25835 : OAI21_X2 port map( A1 => n6051, A2 => n30307, B => n28830, ZN => 
                           n6050);
   U25842 : XOR2_X1 port map( A1 => n22202, A2 => n28835, Z => n4140);
   U25843 : XOR2_X1 port map( A1 => n28837, A2 => n24759, Z => Ciphertext(169))
                           ;
   U25844 : OAI22_X1 port map( A1 => n25825, A2 => n25812, B1 => n24721, B2 => 
                           n24720, ZN => n28837);
   U25850 : AND2_X1 port map( A1 => n20180, A2 => n20181, Z => n28844);
   U25861 : XOR2_X1 port map( A1 => n24562, A2 => n8112, Z => n8110);
   U25868 : NOR2_X1 port map( A1 => n25775, A2 => n15304, ZN => n28854);
   U25870 : NOR2_X2 port map( A1 => n3161, A2 => n3159, ZN => n23328);
   U25872 : NAND2_X2 port map( A1 => n415, A2 => n4595, ZN => n253);
   U25874 : NAND2_X2 port map( A1 => n13539, A2 => n13540, ZN => n22294);
   U25878 : INV_X2 port map( I => n16275, ZN => n21189);
   U25881 : XOR2_X1 port map( A1 => n24824, A2 => n28861, Z => n6328);
   U25882 : XOR2_X1 port map( A1 => n24839, A2 => n28422, Z => n28861);
   U25883 : NAND2_X2 port map( A1 => n15381, A2 => n11006, ZN => n6027);
   U25890 : NAND2_X2 port map( A1 => n15521, A2 => n23689, ZN => n4286);
   U25893 : XOR2_X1 port map( A1 => n28870, A2 => n8917, Z => n28975);
   U25898 : XOR2_X1 port map( A1 => n6058, A2 => n28873, Z => n28872);
   U25909 : XOR2_X1 port map( A1 => n28887, A2 => n24738, Z => Ciphertext(179))
                           ;
   U25911 : NAND2_X2 port map( A1 => n12686, A2 => n14590, ZN => n15704);
   U25912 : NAND2_X1 port map( A1 => n24920, A2 => n3994, ZN => n24930);
   U25917 : NAND2_X2 port map( A1 => n16807, A2 => n16806, ZN => n5889);
   U25918 : AOI22_X2 port map( A1 => n22784, A2 => n7746, B1 => n14212, B2 => 
                           n7747, ZN => n23444);
   U25922 : XOR2_X1 port map( A1 => n23456, A2 => n25373, Z => n22932);
   U25927 : XOR2_X1 port map( A1 => n23430, A2 => n3589, Z => n23254);
   U25935 : XOR2_X1 port map( A1 => n23263, A2 => n26059, Z => n28903);
   U25938 : XOR2_X1 port map( A1 => n20953, A2 => n16703, Z => n6507);
   U25939 : OAI22_X2 port map( A1 => n17002, A2 => n17003, B1 => n9255, B2 => 
                           n10978, ZN => n20953);
   U25940 : XOR2_X1 port map( A1 => n20956, A2 => n28909, Z => n8605);
   U25941 : XOR2_X1 port map( A1 => n8485, A2 => n14854, Z => n28909);
   U25942 : NOR2_X1 port map( A1 => n32877, A2 => n24060, ZN => n13600);
   U25946 : XOR2_X1 port map( A1 => n30443, A2 => n19508, Z => n19564);
   U25948 : NOR2_X2 port map( A1 => n13279, A2 => n18580, ZN => n29182);
   U25951 : XOR2_X1 port map( A1 => n28916, A2 => n11717, Z => n15777);
   U25956 : XOR2_X1 port map( A1 => n9141, A2 => n3929, Z => n6808);
   U25957 : NAND2_X1 port map( A1 => n25606, A2 => n27262, ZN => n28917);
   U25958 : XOR2_X1 port map( A1 => n27841, A2 => n6127, Z => n28918);
   U25961 : NAND2_X2 port map( A1 => n28921, A2 => n21265, ZN => n11214);
   U25972 : OAI21_X1 port map( A1 => n25685, A2 => n32879, B => n28931, ZN => 
                           n25692);
   U25973 : INV_X2 port map( I => n28932, ZN => n701);
   U25974 : XOR2_X1 port map( A1 => n14786, A2 => n4140, Z => n28932);
   U25975 : NOR2_X2 port map( A1 => n28933, A2 => n17910, ZN => n17907);
   U25976 : XOR2_X1 port map( A1 => n1761, A2 => n6726, Z => n6725);
   U25982 : INV_X2 port map( I => n4192, ZN => n9515);
   U25983 : OAI21_X2 port map( A1 => n28938, A2 => n28937, B => n16375, ZN => 
                           n17959);
   U25984 : NOR2_X1 port map( A1 => n22524, A2 => n16665, ZN => n28937);
   U25985 : NOR3_X1 port map( A1 => n16915, A2 => n18827, A3 => n18489, ZN => 
                           n18490);
   U25986 : XOR2_X1 port map( A1 => n13198, A2 => n28941, Z => n28940);
   U25991 : INV_X2 port map( I => n28946, ZN => n470);
   U25992 : NAND2_X2 port map( A1 => n14601, A2 => n28947, ZN => n23450);
   U25993 : OAI21_X1 port map( A1 => n22967, A2 => n22966, B => n28948, ZN => 
                           n28947);
   U25998 : NAND2_X1 port map( A1 => n23664, A2 => n14373, ZN => n15377);
   U25999 : XOR2_X1 port map( A1 => n28953, A2 => n20803, Z => n6683);
   U26001 : AOI21_X1 port map( A1 => n3006, A2 => n13737, B => n2103, ZN => 
                           n28954);
   U26002 : XOR2_X1 port map( A1 => n24632, A2 => n24853, Z => n24377);
   U26005 : NOR2_X1 port map( A1 => n5869, A2 => n8576, ZN => n14004);
   U26010 : OAI21_X2 port map( A1 => n8472, A2 => n8473, B => n1256, ZN => 
                           n28956);
   U26017 : XOR2_X1 port map( A1 => n18404, A2 => Key(163), Z => n18586);
   U26018 : XOR2_X1 port map( A1 => n24813, A2 => n8306, Z => n17096);
   U26021 : AND2_X1 port map( A1 => n22577, A2 => n22664, Z => n14221);
   U26024 : NAND2_X2 port map( A1 => n1897, A2 => n1900, ZN => n8903);
   U26025 : OAI21_X2 port map( A1 => n12021, A2 => n10848, B => n28967, ZN => 
                           n20351);
   U26027 : OAI22_X1 port map( A1 => n14933, A2 => n24958, B1 => n965, B2 => 
                           n14932, ZN => n16115);
   U26030 : NAND2_X1 port map( A1 => n11401, A2 => n21651, ZN => n28972);
   U26034 : XOR2_X1 port map( A1 => n28978, A2 => n30435, Z => n18269);
   U26036 : INV_X2 port map( I => n28979, ZN => n11932);
   U26037 : OAI22_X2 port map( A1 => n29147, A2 => n18381, B1 => n1179, B2 => 
                           n15137, ZN => n19399);
   U26048 : XOR2_X1 port map( A1 => n19371, A2 => n19426, Z => n4028);
   U26050 : NAND2_X1 port map( A1 => n5582, A2 => n20147, ZN => n28982);
   U26051 : NAND2_X1 port map( A1 => n981, A2 => n16431, ZN => n17665);
   U26052 : AOI21_X1 port map( A1 => n20606, A2 => n20130, B => n7292, ZN => 
                           n16481);
   U26056 : AOI21_X2 port map( A1 => n4477, A2 => n1275, B => n4476, ZN => 
                           n5904);
   U26059 : NAND2_X2 port map( A1 => n6025, A2 => n6026, ZN => n18988);
   U26060 : NOR2_X1 port map( A1 => n18978, A2 => n14812, ZN => n16008);
   U26066 : NAND2_X1 port map( A1 => n25666, A2 => n25653, ZN => n28992);
   U26070 : NAND2_X2 port map( A1 => n16274, A2 => n4436, ZN => n19133);
   U26071 : INV_X2 port map( I => n3815, ZN => n19594);
   U26072 : NAND2_X2 port map( A1 => n3055, A2 => n3056, ZN => n3815);
   U26074 : OR2_X1 port map( A1 => n22937, A2 => n31824, Z => n22943);
   U26078 : XOR2_X1 port map( A1 => n5378, A2 => n5539, Z => n28999);
   U26079 : XOR2_X1 port map( A1 => n23328, A2 => n10625, Z => n23464);
   U26080 : XOR2_X1 port map( A1 => n24841, A2 => n29000, Z => n6421);
   U26085 : OAI21_X2 port map( A1 => n29002, A2 => n29001, B => n21406, ZN => 
                           n5801);
   U26090 : XOR2_X1 port map( A1 => n5512, A2 => n27481, Z => n11325);
   U26091 : XOR2_X1 port map( A1 => n29004, A2 => n18122, Z => Ciphertext(23));
   U26092 : NAND3_X1 port map( A1 => n25314, A2 => n25315, A3 => n32867, ZN => 
                           n25318);
   U26098 : XOR2_X1 port map( A1 => n12764, A2 => n15346, Z => n12763);
   U26101 : XOR2_X1 port map( A1 => n8491, A2 => n12454, Z => n29009);
   U26103 : XOR2_X1 port map( A1 => n8129, A2 => n15305, Z => n29012);
   U26114 : XOR2_X1 port map( A1 => n12067, A2 => n12905, Z => n321);
   U26115 : XOR2_X1 port map( A1 => n26053, A2 => n19647, Z => n14060);
   U26116 : XOR2_X1 port map( A1 => n19371, A2 => n17342, Z => n19647);
   U26119 : XOR2_X1 port map( A1 => n29320, A2 => n30183, Z => n7471);
   U26120 : XOR2_X1 port map( A1 => n29028, A2 => n9822, Z => n9821);
   U26121 : XOR2_X1 port map( A1 => n12381, A2 => n12380, Z => n29029);
   U26122 : NAND3_X2 port map( A1 => n9728, A2 => n3269, A3 => n3272, ZN => 
                           n14049);
   U26125 : XOR2_X1 port map( A1 => n18200, A2 => n29032, Z => n18199);
   U26128 : NOR2_X1 port map( A1 => n14321, A2 => n7940, ZN => n8202);
   U26130 : XOR2_X1 port map( A1 => n24794, A2 => n24795, Z => n29033);
   U26131 : XOR2_X1 port map( A1 => n20687, A2 => n20834, Z => n7570);
   U26132 : XOR2_X1 port map( A1 => n8728, A2 => n12459, Z => n20834);
   U26134 : INV_X2 port map( I => n19951, ZN => n29035);
   U26137 : XOR2_X1 port map( A1 => n10738, A2 => n476, Z => n29039);
   U26146 : XOR2_X1 port map( A1 => n4236, A2 => n29046, Z => n7859);
   U26149 : AOI21_X1 port map( A1 => n3843, A2 => n13627, B => n29049, ZN => 
                           n29048);
   U26151 : NAND2_X1 port map( A1 => n29051, A2 => n7503, ZN => n7481);
   U26152 : NAND2_X1 port map( A1 => n17635, A2 => n13971, ZN => n8536);
   U26153 : NAND2_X2 port map( A1 => n10062, A2 => n25897, ZN => n7413);
   U26157 : XOR2_X1 port map( A1 => n20966, A2 => n29054, Z => n8496);
   U26159 : OAI21_X1 port map( A1 => n1207, A2 => n25284, B => n32882, ZN => 
                           n11294);
   U26162 : OR2_X1 port map( A1 => n29255, A2 => n10558, Z => n7148);
   U26166 : XOR2_X1 port map( A1 => n8630, A2 => n22066, Z => n29057);
   U26171 : INV_X2 port map( I => n29064, ZN => n9959);
   U26177 : NOR2_X1 port map( A1 => n28987, A2 => n18556, ZN => n10374);
   U26182 : NAND3_X2 port map( A1 => n6659, A2 => n14906, A3 => n16732, ZN => 
                           n29071);
   U26185 : OAI21_X2 port map( A1 => n29073, A2 => n18561, B => n18560, ZN => 
                           n19123);
   U26186 : NAND2_X1 port map( A1 => n18556, A2 => n16522, ZN => n29074);
   U26187 : INV_X2 port map( I => n29075, ZN => n23949);
   U26190 : OAI21_X1 port map( A1 => n25093, A2 => n25106, B => n18175, ZN => 
                           n29076);
   U26195 : NAND2_X1 port map( A1 => n828, A2 => n18776, ZN => n29149);
   U26200 : BUF_X2 port map( I => n498, Z => n29087);
   U26201 : XOR2_X1 port map( A1 => n29090, A2 => n5150, Z => n15621);
   U26207 : NOR2_X1 port map( A1 => n27637, A2 => n676, ZN => n29094);
   U26208 : AOI21_X1 port map( A1 => n29095, A2 => n25830, B => n25829, ZN => 
                           n25833);
   U26211 : INV_X1 port map( I => n3005, ZN => n29099);
   U26214 : OAI21_X1 port map( A1 => n11939, A2 => n17331, B => n13934, ZN => 
                           n17330);
   U26215 : NAND3_X1 port map( A1 => n24039, A2 => n23659, A3 => n14195, ZN => 
                           n23663);
   U26225 : XOR2_X1 port map( A1 => n19571, A2 => n31361, Z => n19492);
   U26226 : NOR2_X1 port map( A1 => n25005, A2 => n2876, ZN => n29110);
   U26228 : NAND2_X1 port map( A1 => n23715, A2 => n29498, ZN => n29111);
   U26235 : XOR2_X1 port map( A1 => n12212, A2 => n29119, Z => n8416);
   U26236 : XOR2_X1 port map( A1 => n14293, A2 => n11034, Z => n29119);
   U26238 : XOR2_X1 port map( A1 => n24024, A2 => n26126, Z => n15518);
   U26240 : XOR2_X1 port map( A1 => n2591, A2 => n2589, Z => n11348);
   U26241 : NAND2_X1 port map( A1 => n1951, A2 => n16809, ZN => n12485);
   U26243 : XOR2_X1 port map( A1 => n5380, A2 => n5381, Z => n5382);
   U26244 : NAND2_X2 port map( A1 => n29124, A2 => n14587, ZN => n8058);
   U26248 : AOI21_X1 port map( A1 => n5827, A2 => n5828, B => n575, ZN => n5826
                           );
   U26252 : NAND3_X1 port map( A1 => n30285, A2 => n25577, A3 => n6092, ZN => 
                           n4056);
   U26253 : INV_X1 port map( I => n13541, ZN => n29134);
   U26259 : XOR2_X1 port map( A1 => n3517, A2 => n3518, Z => n29139);
   U26262 : XOR2_X1 port map( A1 => n7759, A2 => n7761, Z => n8044);
   U26267 : XOR2_X1 port map( A1 => n29236, A2 => n6545, Z => n24470);
   U26268 : NAND2_X2 port map( A1 => n5311, A2 => n29149, ZN => n2150);
   U26269 : INV_X2 port map( I => n2971, ZN => n8787);
   U26272 : NAND2_X1 port map( A1 => n193, A2 => n13922, ZN => n29152);
   U26274 : BUF_X2 port map( I => n23530, Z => n29155);
   U26276 : INV_X2 port map( I => n32078, ZN => n29158);
   U26277 : XOR2_X1 port map( A1 => n29159, A2 => n8302, Z => n12517);
   U26278 : XOR2_X1 port map( A1 => n15527, A2 => n12519, Z => n29159);
   U26283 : NOR2_X2 port map( A1 => n3998, A2 => n13076, ZN => n10974);
   U26285 : XOR2_X1 port map( A1 => n7452, A2 => n29285, Z => n20740);
   U26287 : XOR2_X1 port map( A1 => n4419, A2 => n4418, Z => n4449);
   U26289 : XOR2_X1 port map( A1 => Plaintext(36), A2 => Key(36), Z => n4200);
   U26293 : OAI21_X2 port map( A1 => n1702, A2 => n10908, B => n1486, ZN => 
                           n1484);
   U26302 : XOR2_X1 port map( A1 => n28939, A2 => n24801, Z => n15471);
   U26303 : NAND2_X1 port map( A1 => n29172, A2 => n32441, ZN => n7789);
   U26304 : OAI21_X1 port map( A1 => n1319, A2 => n230, B => n6351, ZN => 
                           n29172);
   U26306 : XOR2_X1 port map( A1 => n12675, A2 => n24479, Z => n24644);
   U26312 : XOR2_X1 port map( A1 => n19634, A2 => n19675, Z => n19444);
   U26313 : NAND2_X2 port map( A1 => n19065, A2 => n7591, ZN => n19675);
   U26318 : XOR2_X1 port map( A1 => n29189, A2 => n25126, Z => Ciphertext(56));
   U26319 : AOI22_X1 port map( A1 => n25125, A2 => n25127, B1 => n12250, B2 => 
                           n12251, ZN => n29189);
   U26326 : AOI21_X2 port map( A1 => n13460, A2 => n30437, B => n10410, ZN => 
                           n29196);
   U26329 : NAND2_X2 port map( A1 => n252, A2 => n22397, ZN => n22396);
   U26334 : NAND2_X2 port map( A1 => n29634, A2 => n5317, ZN => n24005);
   U26340 : NAND2_X1 port map( A1 => n15115, A2 => n270, ZN => n18499);
   U26341 : NAND2_X1 port map( A1 => n24117, A2 => n30505, ZN => n9374);
   U26344 : INV_X2 port map( I => n29203, ZN => n16981);
   U26346 : XOR2_X1 port map( A1 => n23444, A2 => n25213, Z => n29206);
   U26349 : XOR2_X1 port map( A1 => n2484, A2 => n9361, Z => n4133);
   U26351 : AOI21_X1 port map( A1 => n1439, A2 => n18710, B => n328, ZN => 
                           n18509);
   U26352 : XOR2_X1 port map( A1 => Plaintext(128), A2 => Key(128), Z => n11707
                           );
   U26357 : XOR2_X1 port map( A1 => n30193, A2 => n19675, Z => n19432);
   U26359 : NAND2_X1 port map( A1 => n21538, A2 => n18235, ZN => n29212);
   U26362 : OAI21_X2 port map( A1 => n29214, A2 => n9095, B => n20875, ZN => 
                           n21857);
   U26366 : NAND3_X2 port map( A1 => n6564, A2 => n6567, A3 => n6563, ZN => 
                           n6974);
   U26374 : INV_X2 port map( I => n21193, ZN => n16440);
   U26375 : XOR2_X1 port map( A1 => n2524, A2 => n2526, Z => n21193);
   U26380 : XOR2_X1 port map( A1 => n9013, A2 => n9010, Z => n15917);
   U26381 : NOR2_X1 port map( A1 => n25130, A2 => n25124, ZN => n29227);
   U26382 : INV_X2 port map( I => n29228, ZN => n1850);
   U26385 : INV_X2 port map( I => n29230, ZN => n510);
   U26389 : NAND2_X2 port map( A1 => n25136, A2 => n25135, ZN => n25154);
   U26395 : BUF_X2 port map( I => n12792, Z => n29234);
   U26400 : OAI21_X2 port map( A1 => n15040, A2 => n8909, B => n8908, ZN => 
                           n19624);
   U26401 : NAND2_X2 port map( A1 => n20171, A2 => n20172, ZN => n20680);
   U26405 : XOR2_X1 port map( A1 => n6079, A2 => n6078, Z => n29244);
   U26406 : NOR2_X1 port map( A1 => n19257, A2 => n19137, ZN => n29245);
   U26413 : XOR2_X1 port map( A1 => n13645, A2 => n14293, Z => n12410);
   U26415 : INV_X2 port map( I => n12379, ZN => n13348);
   U26420 : INV_X2 port map( I => n2956, ZN => n3030);
   U26421 : XNOR2_X1 port map( A1 => n22206, A2 => n3583, ZN => n29260);
   U26423 : INV_X2 port map( I => n17109, ZN => n1289);
   U26425 : AOI21_X2 port map( A1 => n22020, A2 => n1117, B => n2257, ZN => 
                           n2256);
   U26428 : OR2_X1 port map( A1 => n22707, A2 => n32089, Z => n29266);
   U26431 : INV_X2 port map( I => n5880, ZN => n23860);
   U26438 : XNOR2_X1 port map( A1 => n1231, A2 => n16587, ZN => n29274);
   U26441 : INV_X1 port map( I => n25150, ZN => n25120);
   U26444 : INV_X2 port map( I => n5019, ZN => n16632);
   U1504 : AOI21_X2 port map( A1 => n18488, A2 => n14831, B => n18490, ZN => 
                           n9183);
   U1964 : INV_X2 port map( I => n19206, ZN => n7176);
   U6752 : AOI21_X2 port map( A1 => n6850, A2 => n31456, B => n6849, ZN => 
                           n2001);
   U8793 : NOR2_X2 port map( A1 => n17843, A2 => n18895, ZN => n14091);
   U12023 : INV_X2 port map( I => n26969, ZN => n1630);
   U3103 : OR2_X1 port map( A1 => n4378, A2 => n9064, Z => n12572);
   U8729 : OAI21_X2 port map( A1 => n15695, A2 => n18659, B => n2107, ZN => 
                           n15151);
   U15014 : INV_X2 port map( I => n14864, ZN => n17887);
   U7211 : INV_X2 port map( I => n3192, ZN => n11601);
   U22246 : INV_X2 port map( I => n21671, ZN => n21668);
   U11943 : INV_X2 port map( I => n15343, ZN => n8919);
   U2415 : NOR2_X2 port map( A1 => n4835, A2 => n30817, ZN => n11280);
   U4768 : BUF_X2 port map( I => n606, Z => n28869);
   U23141 : INV_X2 port map( I => n32532, ZN => n28472);
   U2323 : NAND2_X2 port map( A1 => n25756, A2 => n2967, ZN => n4708);
   U4471 : BUF_X2 port map( I => n9624, Z => n7546);
   U14451 : INV_X4 port map( I => n9678, ZN => n8197);
   U7067 : AOI22_X2 port map( A1 => n6447, A2 => n27178, B1 => n21720, B2 => 
                           n1007, ZN => n2393);
   U1274 : NAND2_X2 port map( A1 => n14049, A2 => n17544, ZN => n9808);
   U1357 : NOR2_X2 port map( A1 => n161, A2 => n29003, ZN => n12625);
   U18501 : NAND2_X2 port map( A1 => n14010, A2 => n13168, ZN => n18261);
   U1131 : NOR2_X2 port map( A1 => n26412, A2 => n26411, ZN => n2466);
   U9119 : AOI21_X2 port map( A1 => n2023, A2 => n1732, B => n1731, ZN => n1730
                           );
   U1053 : NAND2_X2 port map( A1 => n20302, A2 => n20075, ZN => n9588);
   U1036 : NOR2_X2 port map( A1 => n27529, A2 => n17716, ZN => n2395);
   U20028 : INV_X2 port map( I => n10197, ZN => n16136);
   U26110 : NAND3_X1 port map( A1 => n29020, A2 => n20022, A3 => n20021, ZN => 
                           n19657);
   U2707 : NOR2_X2 port map( A1 => n13969, A2 => n17299, ZN => n28199);
   U23943 : INV_X4 port map( I => n17522, ZN => n21367);
   U3486 : NOR2_X2 port map( A1 => n16569, A2 => n18007, ZN => n18835);
   U16423 : NAND3_X1 port map( A1 => n27296, A2 => n22913, A3 => n29317, ZN => 
                           n4711);
   U10180 : INV_X2 port map( I => n18101, ZN => n1572);
   U515 : AOI22_X2 port map( A1 => n22775, A2 => n15718, B1 => n18241, B2 => 
                           n31861, ZN => n22777);
   U20600 : OR2_X1 port map( A1 => n14329, A2 => n11443, Z => n11442);
   U1022 : INV_X2 port map( I => n21707, ZN => n27649);
   U15785 : INV_X2 port map( I => n19197, ZN => n9880);
   U6937 : BUF_X4 port map( I => n23003, Z => n13159);
   U11034 : NAND2_X2 port map( A1 => n18094, A2 => n14017, ZN => n16818);
   U8775 : NAND2_X2 port map( A1 => n18705, A2 => n18743, ZN => n18256);
   U718 : INV_X2 port map( I => n20652, ZN => n1340);
   U3578 : NOR2_X2 port map( A1 => n11460, A2 => n10182, ZN => n18407);
   U2337 : BUF_X4 port map( I => n21350, Z => n21566);
   U898 : NOR2_X2 port map( A1 => n19325, A2 => n9646, ZN => n19185);
   U5425 : OAI21_X2 port map( A1 => n20631, A2 => n20381, B => n8998, ZN => 
                           n8994);
   U1631 : NOR2_X1 port map( A1 => n14197, A2 => n14196, ZN => n14311);
   U1355 : OAI21_X2 port map( A1 => n3311, A2 => n9563, B => n7804, ZN => n1677
                           );
   U8307 : OR2_X1 port map( A1 => n22425, A2 => n22602, Z => n12334);
   U21451 : NOR2_X2 port map( A1 => n21781, A2 => n517, ZN => n12545);
   U12314 : OAI21_X2 port map( A1 => n1458, A2 => n17662, B => n14210, ZN => 
                           n11730);
   U1006 : INV_X2 port map( I => n17167, ZN => n18737);
   U15126 : INV_X2 port map( I => n20565, ZN => n20527);
   U1474 : OAI21_X2 port map( A1 => n13495, A2 => n5162, B => n24, ZN => n8863)
                           ;
   U7538 : NAND2_X2 port map( A1 => n12490, A2 => n18572, ZN => n18386);
   U10190 : INV_X2 port map( I => n18402, ZN => n18730);
   U6648 : NAND2_X2 port map( A1 => n9838, A2 => n18337, ZN => n9837);
   U1000 : NAND2_X2 port map( A1 => n18759, A2 => n18761, ZN => n9838);
   U1237 : INV_X1 port map( I => n16847, ZN => n10017);
   U1059 : NAND2_X2 port map( A1 => n5843, A2 => n13113, ZN => n1533);
   U827 : NOR2_X2 port map( A1 => n15381, A2 => n20066, ZN => n19935);
   U11996 : OAI21_X1 port map( A1 => n6779, A2 => n6780, B => n31139, ZN => 
                           n1654);
   U2615 : OAI21_X2 port map( A1 => n1647, A2 => n14641, B => n6599, ZN => 
                           n13188);
   U2673 : OAI21_X2 port map( A1 => n6133, A2 => n1125, B => n3970, ZN => n2407
                           );
   U4694 : NAND2_X2 port map( A1 => n883, A2 => n3800, ZN => n8542);
   U22865 : INV_X2 port map( I => n14439, ZN => n21239);
   U17993 : NAND2_X2 port map( A1 => n13657, A2 => n1039, ZN => n13656);
   U15431 : AOI21_X2 port map( A1 => n9654, A2 => n22353, B => n8918, ZN => 
                           n9224);
   U2720 : NAND2_X2 port map( A1 => n29173, A2 => n3184, ZN => n11383);
   U1135 : NOR2_X2 port map( A1 => n1889, A2 => n26997, ZN => n20751);
   U6350 : BUF_X2 port map( I => n8471, Z => n7957);
   U1494 : NAND2_X2 port map( A1 => n16740, A2 => n25971, ZN => n19261);
   U852 : INV_X4 port map( I => n14210, ZN => n1362);
   U1267 : INV_X2 port map( I => n30099, ZN => n2566);
   U23643 : INV_X2 port map( I => n16845, ZN => n21395);
   U393 : INV_X2 port map( I => n22983, ZN => n22836);
   U9338 : AOI21_X2 port map( A1 => n18013, A2 => n15853, B => n18012, ZN => 
                           n14856);
   U3359 : INV_X4 port map( I => n11985, ZN => n13985);
   U7224 : INV_X2 port map( I => n8700, ZN => n16639);
   U3964 : NOR2_X2 port map( A1 => n20377, A2 => n20450, ZN => n20202);
   U5992 : INV_X2 port map( I => n18459, ZN => n11380);
   U10892 : OR2_X2 port map( A1 => n15955, A2 => n28231, Z => n18563);
   U7398 : OAI22_X2 port map( A1 => n19960, A2 => n6748, B1 => n31906, B2 => 
                           n19961, ZN => n6733);
   U5500 : INV_X2 port map( I => n10423, ZN => n10015);
   U5809 : INV_X2 port map( I => n21726, ZN => n22201);
   U16885 : AOI21_X2 port map( A1 => n10374, A2 => n11864, B => n5805, ZN => 
                           n6025);
   U9919 : INV_X2 port map( I => n20150, ZN => n4587);
   U1303 : INV_X2 port map( I => n20374, ZN => n8268);
   U552 : INV_X2 port map( I => n21877, ZN => n1315);
   U7523 : INV_X4 port map( I => n7161, ZN => n18983);
   U10928 : INV_X1 port map( I => n30832, ZN => n27686);
   U5663 : NAND2_X2 port map( A1 => n10757, A2 => n10288, ZN => n28160);
   U8731 : OAI21_X2 port map( A1 => n31986, A2 => n2509, B => n711, ZN => n2508
                           );
   U6675 : INV_X2 port map( I => n17638, ZN => n22641);
   U810 : INV_X2 port map( I => n29101, ZN => n29261);
   U6741 : INV_X2 port map( I => n25107, ZN => n1203);
   U6046 : OAI21_X2 port map( A1 => n32038, A2 => n7771, B => n34057, ZN => 
                           n7770);
   U2522 : NAND2_X2 port map( A1 => n23017, A2 => n9377, ZN => n22882);
   U1990 : AOI21_X2 port map( A1 => n17112, A2 => n24005, B => n1245, ZN => 
                           n4521);
   U945 : INV_X2 port map( I => n11085, ZN => n19310);
   U2870 : NOR2_X2 port map( A1 => n8616, A2 => n20056, ZN => n17713);
   U1008 : INV_X4 port map( I => n29309, ZN => n711);
   U2493 : NAND2_X2 port map( A1 => n8657, A2 => n1141, ZN => n9906);
   U4210 : BUF_X4 port map( I => n20605, Z => n7577);
   U17914 : AOI21_X1 port map( A1 => n636, A2 => n1805, B => n28568, ZN => 
                           n13965);
   U21021 : OAI21_X2 port map( A1 => n17764, A2 => n996, B => n13664, ZN => 
                           n13414);
   U3889 : CLKBUF_X4 port map( I => n23130, Z => n23832);
   U9380 : NOR2_X2 port map( A1 => n15589, A2 => n5595, ZN => n21439);
   U3326 : BUF_X2 port map( I => n14834, Z => n375);
   U2202 : NOR2_X2 port map( A1 => n21763, A2 => n21761, ZN => n21762);
   U499 : INV_X2 port map( I => n27799, ZN => n23754);
   U5897 : INV_X2 port map( I => n11958, ZN => n20055);
   U3252 : INV_X2 port map( I => n20460, ZN => n20606);
   U6673 : NAND2_X2 port map( A1 => n12238, A2 => n18891, ZN => n6888);
   U4818 : NAND2_X2 port map( A1 => n18240, A2 => n1719, ZN => n22874);
   U21431 : NAND2_X2 port map( A1 => n31726, A2 => n18973, ZN => n15417);
   U2473 : NAND2_X2 port map( A1 => n1087, A2 => n24283, ZN => n4604);
   U3548 : INV_X2 port map( I => n16356, ZN => n1087);
   U10055 : INV_X2 port map( I => n27921, ZN => n17725);
   U9881 : NAND2_X1 port map( A1 => n16298, A2 => n20044, ZN => n14033);
   U8022 : INV_X1 port map( I => n1284, ZN => n16367);
   U5727 : INV_X4 port map( I => n13998, ZN => n23953);
   U951 : AOI21_X2 port map( A1 => n11719, A2 => n21754, B => n27649, ZN => 
                           n6728);
   U16351 : INV_X2 port map( I => n11515, ZN => n13367);
   U12674 : INV_X2 port map( I => n16297, ZN => n23101);
   U5284 : NAND2_X2 port map( A1 => n31982, A2 => n7190, ZN => n4375);
   U2961 : OR2_X1 port map( A1 => n4177, A2 => n28615, Z => n17055);
   U13296 : INV_X2 port map( I => n621, ZN => n22462);
   U506 : NAND2_X2 port map( A1 => n9243, A2 => n9244, ZN => n27126);
   U15176 : OAI22_X1 port map( A1 => n25320, A2 => n16041, B1 => n25312, B2 => 
                           n25322, ZN => n8629);
   U10703 : AOI22_X2 port map( A1 => n33104, A2 => n4069, B1 => n23705, B2 => 
                           n23897, ZN => n4536);
   U3839 : NAND2_X2 port map( A1 => n27377, A2 => n14118, ZN => n23976);
   U6672 : NAND2_X2 port map( A1 => n18759, A2 => n18601, ZN => n18289);
   U8623 : NAND2_X2 port map( A1 => n29378, A2 => n12502, ZN => n12798);
   U2959 : INV_X2 port map( I => n31095, ZN => n18618);
   U8077 : INV_X2 port map( I => n12490, ZN => n26318);
   U5191 : INV_X1 port map( I => n18540, ZN => n18723);
   U9075 : NOR2_X2 port map( A1 => n24139, A2 => n30969, ZN => n9257);
   U12491 : INV_X2 port map( I => n31671, ZN => n27097);
   U6075 : INV_X4 port map( I => n29063, ZN => n1214);
   U1201 : NOR2_X2 port map( A1 => n20406, A2 => n1349, ZN => n15714);
   U1017 : INV_X2 port map( I => n14640, ZN => n14641);
   U3148 : NOR2_X2 port map( A1 => n7317, A2 => n6473, ZN => n6494);
   U21488 : OAI21_X2 port map( A1 => n8683, A2 => n803, B => n8577, ZN => 
                           n28138);
   U5713 : NAND2_X2 port map( A1 => n8990, A2 => n22908, ZN => n16898);
   U1444 : INV_X2 port map( I => n28082, ZN => n1366);
   U12546 : NAND2_X2 port map( A1 => n1655, A2 => n1654, ZN => n11604);
   U10001 : NOR2_X2 port map( A1 => n18284, A2 => n18285, ZN => n18299);
   U5859 : INV_X4 port map( I => n5548, ZN => n12966);
   U2036 : NOR2_X2 port map( A1 => n11848, A2 => n21811, ZN => n9206);
   U4600 : OAI21_X2 port map( A1 => n12562, A2 => n861, B => n4123, ZN => 
                           n10491);
   U15643 : INV_X2 port map( I => n24645, ZN => n24559);
   U412 : INV_X2 port map( I => n29294, ZN => n23950);
   U907 : INV_X2 port map( I => n16354, ZN => n14734);
   U13465 : NAND2_X2 port map( A1 => n28831, A2 => n803, ZN => n8577);
   U4169 : AOI21_X2 port map( A1 => n23815, A2 => n6694, B => n8525, ZN => 
                           n26631);
   U10725 : NOR2_X2 port map( A1 => n9444, A2 => n23350, ZN => n9443);
   U6331 : BUF_X4 port map( I => n11208, Z => n10699);
   U2677 : INV_X2 port map( I => n17641, ZN => n25586);
   U285 : INV_X4 port map( I => n25987, ZN => n23938);
   U10835 : INV_X4 port map( I => n26606, ZN => n2858);
   U8942 : NAND2_X2 port map( A1 => n13643, A2 => n13359, ZN => n5810);
   U812 : AND2_X2 port map( A1 => n9630, A2 => n3392, Z => n26098);
   U3703 : NAND2_X2 port map( A1 => n15149, A2 => n31614, ZN => n2118);
   U2460 : NAND2_X1 port map( A1 => n14032, A2 => n17609, ZN => n27992);
   U1311 : BUF_X4 port map( I => n6997, Z => n25966);
   U5665 : OAI21_X2 port map( A1 => n14227, A2 => n18073, B => n16260, ZN => 
                           n15636);
   U3060 : AOI21_X2 port map( A1 => n23074, A2 => n23073, B => n8953, ZN => 
                           n13690);
   U4713 : NAND2_X2 port map( A1 => n13042, A2 => n14832, ZN => n3800);
   U4748 : INV_X2 port map( I => n5051, ZN => n12665);
   U13106 : BUF_X4 port map( I => n15144, Z => n26891);
   U5922 : OAI21_X2 port map( A1 => n32952, A2 => n4210, B => n4714, ZN => 
                           n5329);
   U715 : NOR2_X2 port map( A1 => n22343, A2 => n7090, ZN => n26991);
   U5422 : INV_X2 port map( I => n8795, ZN => n10766);
   U2699 : OAI21_X2 port map( A1 => n19144, A2 => n2871, B => n19254, ZN => 
                           n2870);
   U4599 : INV_X2 port map( I => n25966, ZN => n1160);
   U9206 : INV_X2 port map( I => n17373, ZN => n23826);
   U20627 : NAND3_X2 port map( A1 => n20038, A2 => n20039, A3 => n20135, ZN => 
                           n20042);
   U1373 : NOR2_X2 port map( A1 => n19451, A2 => n20056, ZN => n20053);
   U2519 : INV_X4 port map( I => n19724, ZN => n20028);
   U22284 : AOI21_X2 port map( A1 => n10273, A2 => n11350, B => n10271, ZN => 
                           n28285);
   U12832 : NAND2_X2 port map( A1 => n16842, A2 => n29372, ZN => n26834);
   U2840 : NOR3_X2 port map( A1 => n30692, A2 => n20097, A3 => n16630, ZN => 
                           n10241);
   U1193 : INV_X2 port map( I => n20837, ZN => n27015);
   U176 : INV_X2 port map( I => n30795, ZN => n968);
   U22939 : NOR2_X2 port map( A1 => n24062, A2 => n24156, ZN => n28391);
   U8047 : AOI21_X2 port map( A1 => n22689, A2 => n14493, B => n5769, ZN => 
                           n5770);
   U3124 : AND3_X1 port map( A1 => n22990, A2 => n29313, A3 => n15829, Z => 
                           n13430);
   U8867 : BUF_X2 port map( I => Key(116), Z => n25910);
   U12446 : NAND2_X2 port map( A1 => n27279, A2 => n16923, ZN => n6398);
   U3921 : INV_X2 port map( I => n920, ZN => n27024);
   U15897 : INV_X2 port map( I => n4236, ZN => n19784);
   U2883 : AND2_X1 port map( A1 => n6489, A2 => n6544, Z => n21855);
   U4033 : INV_X2 port map( I => n16442, ZN => n26390);
   U504 : INV_X2 port map( I => n23120, ZN => n1262);
   U5437 : INV_X2 port map( I => n7852, ZN => n20608);
   U7033 : INV_X4 port map( I => n22433, ZN => n22651);
   U10229 : BUF_X2 port map( I => Key(167), Z => n25929);
   U16428 : INV_X2 port map( I => n16392, ZN => n10862);
   U1402 : NOR2_X2 port map( A1 => n19820, A2 => n28600, ZN => n15246);
   U8774 : NAND2_X2 port map( A1 => n18764, A2 => n27981, ZN => n18766);
   U1179 : NAND2_X2 port map( A1 => n10280, A2 => n23030, ZN => n22738);
   U302 : INV_X2 port map( I => n5097, ZN => n11888);
   U3582 : INV_X2 port map( I => n13348, ZN => n1163);
   U13030 : INV_X4 port map( I => n11322, ZN => n19267);
   U24404 : AOI21_X2 port map( A1 => n18989, A2 => n18988, B => n19034, ZN => 
                           n18992);
   U8690 : NOR2_X2 port map( A1 => n1385, A2 => n19089, ZN => n19034);
   U1259 : INV_X2 port map( I => n9403, ZN => n1159);
   U5796 : INV_X2 port map( I => n14297, ZN => n3860);
   U17438 : INV_X1 port map( I => n13176, ZN => n24217);
   U931 : AOI21_X2 port map( A1 => n12545, A2 => n11861, B => n29434, ZN => 
                           n28155);
   U3101 : AOI21_X2 port map( A1 => n9192, A2 => n16751, B => n25186, ZN => 
                           n8481);
   U10536 : NAND2_X2 port map( A1 => n24296, A2 => n24297, ZN => n3780);
   U5668 : BUF_X4 port map( I => n9890, Z => n2913);
   U6223 : INV_X2 port map( I => n12821, ZN => n1980);
   U4245 : BUF_X4 port map( I => n19285, Z => n17311);
   U822 : BUF_X2 port map( I => n34162, Z => n28568);
   U8344 : CLKBUF_X4 port map( I => n8605, Z => n1146);
   U1503 : NAND2_X2 port map( A1 => n784, A2 => n13200, ZN => n27274);
   U14671 : OAI21_X2 port map( A1 => n27941, A2 => n15239, B => n10740, ZN => 
                           n10739);
   U13439 : NAND2_X1 port map( A1 => n14775, A2 => n2522, ZN => n14774);
   U4022 : INV_X2 port map( I => n16384, ZN => n16781);
   U2855 : OR2_X1 port map( A1 => n4146, A2 => n25628, Z => n277);
   U8093 : INV_X2 port map( I => n15617, ZN => n22658);
   U9615 : NAND3_X2 port map( A1 => n3852, A2 => n23021, A3 => n3851, ZN => 
                           n23202);
   U457 : INV_X2 port map( I => n28123, ZN => n4408);
   U1366 : INV_X2 port map( I => n567, ZN => n13994);
   U12825 : INV_X2 port map( I => n398, ZN => n16184);
   U2799 : INV_X2 port map( I => n23018, ZN => n1279);
   U7122 : INV_X4 port map( I => n21665, ZN => n1134);
   U3341 : NAND2_X2 port map( A1 => n28328, A2 => n31798, ZN => n15830);
   U10955 : INV_X2 port map( I => n2130, ZN => n22722);
   U2669 : AOI21_X2 port map( A1 => n21692, A2 => n21857, B => n2797, ZN => 
                           n15847);
   U9230 : NAND2_X2 port map( A1 => n3770, A2 => n896, ZN => n6965);
   U5598 : NOR2_X2 port map( A1 => n13030, A2 => n12036, ZN => n13029);
   U537 : NAND2_X2 port map( A1 => n9844, A2 => n6236, ZN => n26796);
   U6024 : INV_X2 port map( I => n25755, ZN => n1212);
   U1094 : AOI21_X2 port map( A1 => n7226, A2 => n21354, B => n2088, ZN => 
                           n3698);
   U7820 : AOI21_X2 port map( A1 => n8850, A2 => n27615, B => n8849, ZN => 
                           n8848);
   U1287 : NAND2_X2 port map( A1 => n16488, A2 => n12345, ZN => n12344);
   U7708 : NAND3_X1 port map( A1 => n4451, A2 => n24711, A3 => n4452, ZN => 
                           n3835);
   U5664 : NOR2_X2 port map( A1 => n14972, A2 => n24251, ZN => n17581);
   U10974 : NAND2_X2 port map( A1 => n12762, A2 => n23068, ZN => n14914);
   U6799 : NOR2_X2 port map( A1 => n16620, A2 => n23721, ZN => n11812);
   U123 : INV_X4 port map( I => n4490, ZN => n4407);
   U1994 : NAND3_X2 port map( A1 => n7086, A2 => n7085, A3 => n7084, ZN => 
                           n28251);
   U1005 : INV_X2 port map( I => n16819, ZN => n18485);
   U3277 : NAND2_X2 port map( A1 => n26750, A2 => n24106, ZN => n24093);
   U19409 : AOI21_X2 port map( A1 => n26600, A2 => n16354, B => n4656, ZN => 
                           n27831);
   U606 : INV_X4 port map( I => n34163, ZN => n22981);
   U4647 : INV_X2 port map( I => n18688, ZN => n10283);
   U7093 : BUF_X2 port map( I => n21626, Z => n6176);
   U26265 : OAI22_X2 port map( A1 => n1179, A2 => n9787, B1 => n1380, B2 => 
                           n15137, ZN => n29147);
   U1506 : AOI21_X2 port map( A1 => n15814, A2 => n15428, B => n21162, ZN => 
                           n7049);
   U6264 : INV_X2 port map( I => n6975, ZN => n1104);
   U4247 : BUF_X4 port map( I => n19283, Z => n13475);
   U4372 : OAI22_X2 port map( A1 => n26104, A2 => n29115, B1 => n23016, B2 => 
                           n28891, ZN => n13289);
   U7016 : NAND2_X2 port map( A1 => n2177, A2 => n16790, ZN => n26289);
   U17035 : INV_X2 port map( I => n29767, ZN => n14195);
   U6594 : INV_X4 port map( I => n4747, ZN => n1175);
   U6329 : INV_X2 port map( I => n11208, ZN => n21799);
   U41 : INV_X2 port map( I => n14960, ZN => n24972);
   U8717 : INV_X1 port map( I => n2902, ZN => n19035);
   U17631 : INV_X4 port map( I => n6899, ZN => n20489);
   U885 : INV_X2 port map( I => n5848, ZN => n22248);
   U6380 : NAND2_X2 port map( A1 => n3539, A2 => n21780, ZN => n21583);
   U12472 : NAND2_X2 port map( A1 => n10441, A2 => n10442, ZN => n22098);
   U15273 : INV_X1 port map( I => n31960, ZN => n15595);
   U9865 : OAI21_X2 port map( A1 => n20071, A2 => n729, B => n19888, ZN => 
                           n18036);
   U205 : OR2_X2 port map( A1 => n16552, A2 => n7171, Z => n24342);
   U3440 : AND2_X1 port map( A1 => n27921, A2 => n5889, Z => n6566);
   U26343 : NAND2_X1 port map( A1 => n20170, A2 => n20298, ZN => n29202);
   U10089 : NOR2_X2 port map( A1 => n10638, A2 => n10637, ZN => n7286);
   U5915 : INV_X2 port map( I => n13272, ZN => n18142);
   U5326 : BUF_X2 port map( I => n31906, Z => n28767);
   U24357 : OAI21_X2 port map( A1 => n18733, A2 => n18732, B => n18731, ZN => 
                           n18735);
   U5615 : INV_X2 port map( I => n17697, ZN => n22305);
   U1454 : NAND2_X2 port map( A1 => n1491, A2 => n26293, ZN => n19682);
   U6792 : NAND2_X2 port map( A1 => n23965, A2 => n13, ZN => n18120);
   U7186 : NAND2_X2 port map( A1 => n865, A2 => n2738, ZN => n21284);
   U8692 : INV_X2 port map( I => n27242, ZN => n13685);
   U5639 : OAI21_X2 port map( A1 => n22657, A2 => n22658, B => n16503, ZN => 
                           n5766);
   U2241 : NOR2_X2 port map( A1 => n28914, A2 => n654, ZN => n4538);
   U4287 : CLKBUF_X2 port map( I => Key(78), Z => n16504);
   U9064 : INV_X4 port map( I => n24335, ZN => n1235);
   U8433 : NOR2_X2 port map( A1 => n3317, A2 => n21572, ZN => n3316);
   U4030 : BUF_X4 port map( I => n18613, Z => n17223);
   U2201 : NAND2_X2 port map( A1 => n15022, A2 => n21761, ZN => n21850);
   U3820 : INV_X2 port map( I => n21095, ZN => n21408);
   U11605 : OAI21_X2 port map( A1 => n13915, A2 => n33902, B => n6083, ZN => 
                           n15142);
   U3989 : OR3_X1 port map( A1 => n18186, A2 => n1430, A3 => n6215, Z => n10975
                           );
   U1398 : OAI21_X2 port map( A1 => n11052, A2 => n26083, B => n11264, ZN => 
                           n29008);
   U6472 : OAI22_X2 port map( A1 => n10718, A2 => n9419, B1 => n5275, B2 => 
                           n20541, ZN => n9418);
   U8373 : NOR2_X2 port map( A1 => n26358, A2 => n17758, ZN => n7392);
   U5369 : OR2_X2 port map( A1 => n29395, A2 => n3567, Z => n9801);
   U7448 : INV_X1 port map( I => n4386, ZN => n4385);
   U8331 : INV_X2 port map( I => n13367, ZN => n1141);
   U5935 : NAND2_X2 port map( A1 => n12937, A2 => n4016, ZN => n13450);
   U24496 : INV_X2 port map( I => n19419, ZN => n19868);
   U9944 : BUF_X2 port map( I => n31671, Z => n11199);
   U21362 : OAI21_X2 port map( A1 => n27236, A2 => n16783, B => n25520, ZN => 
                           n25521);
   U1189 : NAND2_X2 port map( A1 => n10460, A2 => n7330, ZN => n7332);
   U12423 : INV_X2 port map( I => n16421, ZN => n26777);
   U26417 : INV_X1 port map( I => n21375, ZN => n21374);
   U895 : AOI22_X2 port map( A1 => n17428, A2 => n17773, B1 => n21459, B2 => 
                           n21458, ZN => n11795);
   U21138 : NAND2_X2 port map( A1 => n17699, A2 => n29062, ZN => n20947);
   U9928 : BUF_X4 port map( I => n15237, Z => n20135);
   U3554 : NOR2_X2 port map( A1 => n22705, A2 => n27007, ZN => n16236);
   U26192 : BUF_X4 port map( I => n16136, Z => n29078);
   U13001 : INV_X2 port map( I => n3084, ZN => n20589);
   U10117 : OAI21_X2 port map( A1 => n18517, A2 => n18878, B => n18112, ZN => 
                           n2704);
   U7354 : OAI21_X2 port map( A1 => n8421, A2 => n16243, B => n32408, ZN => 
                           n3825);
   U5097 : OAI21_X2 port map( A1 => n2443, A2 => n21716, B => n911, ZN => n2442
                           );
   U21201 : NOR2_X2 port map( A1 => n15872, A2 => n15506, ZN => n14692);
   U2848 : INV_X2 port map( I => n10717, ZN => n5275);
   U7226 : OR2_X2 port map( A1 => n21184, A2 => n13989, Z => n12756);
   U24283 : OAI21_X2 port map( A1 => n16466, A2 => n18672, B => n18441, ZN => 
                           n18443);
   U4842 : AOI21_X2 port map( A1 => n6121, A2 => n29938, B => n3972, ZN => 
                           n4965);
   U1431 : INV_X4 port map( I => n15110, ZN => n27715);
   U21005 : INV_X1 port map( I => n22490, ZN => n14671);
   U4632 : NOR2_X1 port map( A1 => n1014, A2 => n12028, ZN => n2743);
   U13097 : NOR2_X2 port map( A1 => n6446, A2 => n13685, ZN => n26890);
   U5611 : INV_X2 port map( I => n16896, ZN => n12370);
   U5572 : NOR2_X2 port map( A1 => n31927, A2 => n21, ZN => n2797);
   U2391 : AOI22_X2 port map( A1 => n11802, A2 => n1377, B1 => n26518, B2 => 
                           n10828, ZN => n11801);
   U5491 : INV_X2 port map( I => n19053, ZN => n1181);
   U5692 : OAI21_X2 port map( A1 => n983, A2 => n12259, B => n12910, ZN => 
                           n12909);
   U24023 : INV_X2 port map( I => n17799, ZN => n23813);
   U2824 : NOR2_X2 port map( A1 => n897, A2 => n22876, ZN => n12910);
   U11490 : INV_X2 port map( I => n5111, ZN => n3866);
   U1522 : INV_X2 port map( I => n18626, ZN => n19147);
   U15419 : INV_X1 port map( I => n18186, ZN => n16624);
   U18887 : AND2_X2 port map( A1 => n10303, A2 => n16332, Z => n22479);
   U21571 : NAND2_X2 port map( A1 => n4468, A2 => n15162, ZN => n12516);
   U5526 : INV_X4 port map( I => n18815, ZN => n785);
   U8735 : AOI21_X2 port map( A1 => n4843, A2 => n1188, B => n8043, ZN => n4644
                           );
   U19478 : INV_X2 port map( I => n9118, ZN => n11918);
   U15441 : NAND2_X1 port map( A1 => n10134, A2 => n33972, ZN => n7815);
   U5145 : OAI21_X2 port map( A1 => n18370, A2 => n18369, B => n12120, ZN => 
                           n18371);
   U4821 : NOR2_X1 port map( A1 => n26953, A2 => n12010, ZN => n8995);
   U1742 : OAI21_X2 port map( A1 => n10977, A2 => n18778, B => n10975, ZN => 
                           n3998);
   U19862 : INV_X1 port map( I => n16202, ZN => n28878);
   U23003 : INV_X1 port map( I => n24359, ZN => n14832);
   U5910 : NAND2_X2 port map( A1 => n23606, A2 => n23605, ZN => n16815);
   U12965 : AOI21_X1 port map( A1 => n864, A2 => n33139, B => n2061, ZN => 
                           n2060);
   U23628 : INV_X2 port map( I => n23696, ZN => n16431);
   U3439 : INV_X4 port map( I => n31967, ZN => n1347);
   U12943 : AOI21_X2 port map( A1 => n12865, A2 => n11215, B => n27608, ZN => 
                           n12642);
   U2424 : BUF_X4 port map( I => n31448, Z => n149);
   U1441 : INV_X2 port map( I => n29029, ZN => n12379);
   U1501 : AND2_X2 port map( A1 => n17201, A2 => n8452, Z => n22570);
   U2028 : INV_X4 port map( I => n20092, ZN => n15192);
   U10106 : AOI22_X2 port map( A1 => n18894, A2 => n31724, B1 => n18896, B2 => 
                           n6119, ZN => n6116);
   U10078 : INV_X2 port map( I => n17821, ZN => n20155);
   U5107 : NAND2_X2 port map( A1 => n497, A2 => n18747, ZN => n18433);
   U2464 : BUF_X2 port map( I => n519, Z => n154);
   U5638 : INV_X4 port map( I => n17960, ZN => n12338);
   U16864 : NOR2_X2 port map( A1 => n6699, A2 => n6698, ZN => n10946);
   U10833 : BUF_X2 port map( I => n23905, Z => n12680);
   U13667 : INV_X2 port map( I => n20080, ZN => n20084);
   U22425 : NAND2_X1 port map( A1 => n15191, A2 => n15190, ZN => n28776);
   U12317 : INV_X4 port map( I => n25980, ZN => n1458);
   U7044 : INV_X4 port map( I => n16124, ZN => n17960);
   U9101 : NAND2_X2 port map( A1 => n28296, A2 => n6476, ZN => n7151);
   U661 : INV_X4 port map( I => n27752, ZN => n28328);
   U4244 : BUF_X2 port map( I => n19360, Z => n16444);
   U1971 : OAI21_X2 port map( A1 => n26113, A2 => n16229, B => n21817, ZN => 
                           n5757);
   U1432 : BUF_X2 port map( I => n13510, Z => n29208);
   U12101 : AOI21_X2 port map( A1 => n18878, A2 => n18881, B => n6754, ZN => 
                           n6753);
   U17829 : NOR2_X2 port map( A1 => n18672, A2 => n18881, ZN => n6754);
   U1462 : OAI21_X2 port map( A1 => n19170, A2 => n19171, B => n948, ZN => 
                           n3245);
   U22400 : NOR2_X2 port map( A1 => n34005, A2 => n28721, ZN => n19170);
   U22728 : NOR2_X2 port map( A1 => n25974, A2 => n24251, ZN => n15086);
   U22647 : NAND2_X2 port map( A1 => n20139, A2 => n32141, ZN => n15594);
   U5166 : NOR3_X1 port map( A1 => n1053, A2 => n5889, A3 => n31451, ZN => 
                           n6565);
   U2908 : NAND2_X2 port map( A1 => n18722, A2 => n13279, ZN => n18582);
   U1326 : BUF_X4 port map( I => n1736, Z => n1632);
   U24810 : NAND2_X2 port map( A1 => n21451, A2 => n20950, ZN => n20951);
   U22817 : INV_X4 port map( I => n14458, ZN => n20000);
   U17258 : INV_X4 port map( I => n33740, ZN => n10757);
   U3811 : OR2_X1 port map( A1 => n31970, A2 => n3093, Z => n15284);
   U13638 : INV_X4 port map( I => n8924, ZN => n16473);
   U1981 : AOI22_X2 port map( A1 => n13210, A2 => n13925, B1 => n19046, B2 => 
                           n19047, ZN => n12601);
   U2676 : BUF_X2 port map( I => n23827, Z => n16467);
   U25782 : NAND3_X2 port map( A1 => n14925, A2 => n34149, A3 => n32590, ZN => 
                           n25913);
   U11206 : INV_X1 port map( I => n3911, ZN => n22552);
   U1233 : OAI21_X2 port map( A1 => n30602, A2 => n19256, B => n2703, ZN => 
                           n2124);
   U4695 : BUF_X2 port map( I => n14396, Z => n26337);
   U5814 : OAI21_X2 port map( A1 => n4668, A2 => n18043, B => n21808, ZN => 
                           n21727);
   U6142 : OR2_X1 port map( A1 => n3773, A2 => n22977, Z => n26026);
   U2148 : NAND2_X2 port map( A1 => n5481, A2 => n11399, ZN => n27975);
   U4858 : INV_X2 port map( I => n4740, ZN => n4755);
   U1680 : INV_X1 port map( I => n5511, ZN => n6901);
   U2996 : BUF_X4 port map( I => n11984, Z => n295);
   U7539 : NAND2_X2 port map( A1 => n9837, A2 => n9836, ZN => n4571);
   U725 : OAI22_X2 port map( A1 => n20416, A2 => n20415, B1 => n30931, B2 => 
                           n20414, ZN => n20860);
   U5057 : INV_X2 port map( I => n32595, ZN => n11059);
   U451 : NAND2_X2 port map( A1 => n22488, A2 => n31551, ZN => n75);
   U1302 : NOR3_X2 port map( A1 => n8619, A2 => n2625, A3 => n30152, ZN => 
                           n8618);
   U5392 : OR2_X1 port map( A1 => n15713, A2 => n16167, Z => n27299);
   U12749 : INV_X2 port map( I => n1850, ZN => n9294);
   U1412 : NAND2_X2 port map( A1 => n19884, A2 => n224, ZN => n26357);
   U15510 : OR2_X2 port map( A1 => n12654, A2 => n14290, Z => n7205);
   U4298 : BUF_X2 port map( I => Key(96), Z => n16657);
   U2518 : BUF_X2 port map( I => n19698, Z => n112);
   U2740 : BUF_X2 port map( I => n22625, Z => n16170);
   U5507 : BUF_X2 port map( I => n11272, Z => n6584);
   U11440 : NAND2_X2 port map( A1 => n18213, A2 => n29369, ZN => n18210);
   U2857 : OR2_X1 port map( A1 => n5736, A2 => n2163, Z => n3480);
   U21925 : INV_X1 port map( I => n16440, ZN => n28211);
   U129 : INV_X2 port map( I => n6545, ZN => n24771);
   U10689 : OAI21_X2 port map( A1 => n23682, A2 => n23681, B => n14124, ZN => 
                           n23685);
   U16763 : NOR2_X2 port map( A1 => n11730, A2 => n8775, ZN => n6631);
   U17263 : NAND2_X1 port map( A1 => n11213, A2 => n25658, ZN => n11212);
   U21252 : NOR2_X1 port map( A1 => n12377, A2 => n23034, ZN => n15191);
   U879 : INV_X2 port map( I => n18453, ZN => n1370);
   U389 : INV_X4 port map( I => n33115, ZN => n23045);
   U2808 : BUF_X2 port map( I => n14000, Z => n27841);
   U5 : NAND2_X1 port map( A1 => n11211, A2 => n34094, ZN => n28631);
   U17453 : NAND3_X1 port map( A1 => n18361, A2 => n17792, A3 => n18362, ZN => 
                           n18162);
   U6196 : INV_X2 port map( I => n893, ZN => n8835);
   U6982 : AOI22_X2 port map( A1 => n1669, A2 => n9580, B1 => n13079, B2 => 
                           n22599, ZN => n1668);
   U7162 : OAI21_X2 port map( A1 => n11405, A2 => n28869, B => n21431, ZN => 
                           n13150);
   U5067 : INV_X2 port map( I => n23000, ZN => n16078);
   U11161 : NOR2_X2 port map( A1 => n630, A2 => n28124, ZN => n3521);
   U6197 : INV_X1 port map( I => n14398, ZN => n13125);
   U14822 : NOR2_X2 port map( A1 => n18374, A2 => n18809, ZN => n9785);
   U3108 : INV_X4 port map( I => n635, ZN => n16137);
   U11717 : OAI22_X2 port map( A1 => n26008, A2 => n13537, B1 => n13759, B2 => 
                           n13538, ZN => n13783);
   U23824 : OR2_X2 port map( A1 => n5097, A2 => n29270, Z => n23819);
   U908 : OAI21_X2 port map( A1 => n27326, A2 => n864, B => n1, ZN => n3685);
   U9262 : OAI21_X2 port map( A1 => n32595, A2 => n1275, B => n30502, ZN => 
                           n13460);
   U10879 : NAND2_X1 port map( A1 => n8494, A2 => n17828, ZN => n4779);
   U5113 : INV_X2 port map( I => n606, ZN => n12925);
   U7345 : OAI21_X2 port map( A1 => n15737, A2 => n10340, B => n15735, ZN => 
                           n19912);
   U12921 : INV_X2 port map( I => n16510, ZN => n17717);
   U5535 : AOI22_X2 port map( A1 => n12992, A2 => n10686, B1 => n15002, B2 => 
                           n7512, ZN => n28664);
   U5452 : INV_X2 port map( I => n7014, ZN => n20071);
   U7659 : BUF_X2 port map( I => Key(13), Z => n16696);
   U18598 : AOI21_X2 port map( A1 => n18940, A2 => n19244, B => n27818, ZN => 
                           n18941);
   U7295 : NOR2_X2 port map( A1 => n13589, A2 => n17328, ZN => n20234);
   U18458 : INV_X2 port map( I => n10371, ZN => n15799);
   U2053 : OAI22_X2 port map( A1 => n25591, A2 => n10497, B1 => n9197, B2 => 
                           n13032, ZN => n28557);
   U8172 : NAND2_X2 port map( A1 => n21805, A2 => n3467, ZN => n7501);
   U899 : OAI21_X2 port map( A1 => n1766, A2 => n2283, B => n2280, ZN => n2279)
                           ;
   U5086 : INV_X2 port map( I => n15455, ZN => n26717);
   U1539 : CLKBUF_X4 port map( I => n19348, Z => n27941);
   U21250 : OR2_X1 port map( A1 => n22680, A2 => n32172, Z => n12531);
   U2052 : NAND2_X2 port map( A1 => n10497, A2 => n18151, ZN => n25636);
   U15707 : INV_X4 port map( I => n30885, ZN => n17348);
   U11812 : INV_X2 port map( I => n26278, ZN => n1357);
   U1906 : INV_X2 port map( I => n16781, ZN => n28671);
   U6658 : NAND2_X2 port map( A1 => n6888, A2 => n6889, ZN => n6266);
   U3406 : BUF_X4 port map( I => n8506, Z => n29118);
   U476 : INV_X2 port map( I => n6882, ZN => n5769);
   U7361 : NOR2_X2 port map( A1 => n19884, A2 => n19868, ZN => n20057);
   U11451 : NAND2_X2 port map( A1 => n1915, A2 => n1914, ZN => n1913);
   U5913 : NAND2_X2 port map( A1 => n7730, A2 => n1237, ZN => n6773);
   U13802 : INV_X1 port map( I => n18151, ZN => n28097);
   U3395 : INV_X2 port map( I => n24104, ZN => n15376);
   U3462 : OR2_X1 port map( A1 => n12452, A2 => n26439, Z => n28654);
   U22510 : NOR2_X2 port map( A1 => n31402, A2 => n7310, ZN => n14114);
   U5393 : OAI21_X2 port map( A1 => n31996, A2 => n13869, B => n26727, ZN => 
                           n10441);
   U3371 : INV_X2 port map( I => n31074, ZN => n19254);
   U11072 : OAI21_X1 port map( A1 => n6187, A2 => n28825, B => n5814, ZN => 
                           n2861);
   U11307 : NOR2_X1 port map( A1 => n11582, A2 => n3580, ZN => n3579);
   U18158 : INV_X2 port map( I => n20395, ZN => n7291);
   U13502 : INV_X4 port map( I => n11734, ZN => n21369);
   U11746 : NAND2_X1 port map( A1 => n24950, A2 => n24949, ZN => n26711);
   U14982 : INV_X4 port map( I => n12145, ZN => n16681);
   U2138 : NAND2_X1 port map( A1 => n25256, A2 => n7871, ZN => n26497);
   U3404 : AND2_X1 port map( A1 => n19252, A2 => n8506, Z => n18525);
   U2566 : NAND3_X1 port map( A1 => n25530, A2 => n25588, A3 => n25529, ZN => 
                           n25535);
   U904 : OAI22_X2 port map( A1 => n3468, A2 => n21660, B1 => n3467, B2 => 
                           n21659, ZN => n11053);
   U7670 : BUF_X2 port map( I => Key(17), Z => n25619);
   U5873 : INV_X2 port map( I => n20582, ZN => n12872);
   U8928 : NOR2_X2 port map( A1 => n9114, A2 => n23960, ZN => n9113);
   U6090 : INV_X2 port map( I => n16321, ZN => n7837);
   U20872 : NOR2_X1 port map( A1 => n15215, A2 => n8602, ZN => n12751);
   U15799 : NAND2_X1 port map( A1 => n17172, A2 => n17171, ZN => n4390);
   U9587 : INV_X2 port map( I => n21872, ZN => n21871);
   U3762 : INV_X4 port map( I => n10465, ZN => n3626);
   U17210 : NAND3_X1 port map( A1 => n20487, A2 => n20252, A3 => n5878, ZN => 
                           n11140);
   U21533 : OAI21_X2 port map( A1 => n9876, A2 => n12100, B => n20007, ZN => 
                           n17785);
   U22256 : NAND2_X1 port map( A1 => n15417, A2 => n19267, ZN => n15416);
   U2919 : INV_X4 port map( I => n11390, ZN => n2107);
   U2429 : NOR2_X1 port map( A1 => n27971, A2 => n5936, ZN => n5933);
   U2482 : INV_X1 port map( I => n32998, ZN => n10018);
   U4367 : NAND2_X2 port map( A1 => n27537, A2 => n26222, ZN => n6519);
   U15561 : AOI22_X2 port map( A1 => n21534, A2 => n21566, B1 => n29806, B2 => 
                           n21568, ZN => n8196);
   U16881 : NAND2_X1 port map( A1 => n27358, A2 => n6520, ZN => n2369);
   U10257 : BUF_X2 port map( I => Key(107), Z => n25578);
   U6093 : INV_X2 port map( I => n32317, ZN => n1232);
   U3659 : NOR2_X2 port map( A1 => n7176, A2 => n30010, ZN => n1494);
   U3179 : INV_X1 port map( I => n18874, ZN => n961);
   U3334 : NOR2_X2 port map( A1 => n30355, A2 => n2679, ZN => n2678);
   U21437 : OAI21_X2 port map( A1 => n15141, A2 => n18697, B => n33098, ZN => 
                           n15140);
   U20675 : INV_X2 port map( I => n20102, ZN => n12038);
   U15051 : NOR2_X2 port map( A1 => n5205, A2 => n30573, ZN => n28863);
   U3682 : OAI21_X2 port map( A1 => n10947, A2 => n11521, B => n25997, ZN => 
                           n18949);
   U10166 : BUF_X2 port map( I => n18434, Z => n18705);
   U12217 : INV_X2 port map( I => n10891, ZN => n18683);
   U8660 : NAND2_X1 port map( A1 => n28157, A2 => n19236, ZN => n2599);
   U5672 : AOI22_X2 port map( A1 => n7560, A2 => n16170, B1 => n17955, B2 => 
                           n7559, ZN => n27916);
   U25895 : AOI21_X2 port map( A1 => n17392, A2 => n17393, B => n3562, ZN => 
                           n8425);
   U5468 : INV_X1 port map( I => n14340, ZN => n27412);
   U11408 : NAND2_X1 port map( A1 => n11687, A2 => n16034, ZN => n11686);
   U4550 : NAND4_X2 port map( A1 => n21829, A2 => n21828, A3 => n21827, A4 => 
                           n21832, ZN => n17406);
   U1322 : NAND3_X2 port map( A1 => n13994, A2 => n20028, A3 => n16461, ZN => 
                           n12947);
   U18707 : INV_X4 port map( I => n8408, ZN => n27678);
   U8760 : OAI21_X2 port map( A1 => n18399, A2 => n2596, B => n29309, ZN => 
                           n2595);
   U23330 : INV_X4 port map( I => n15559, ZN => n17624);
   U6566 : INV_X1 port map( I => n16904, ZN => n873);
   U24080 : NAND2_X1 port map( A1 => n12572, A2 => n9065, ZN => n28592);
   U8091 : BUF_X4 port map( I => n29451, Z => n1297);
   U12104 : NAND2_X2 port map( A1 => n16338, A2 => n18576, ZN => n8461);
   U4912 : OAI21_X2 port map( A1 => n8931, A2 => n8930, B => n8929, ZN => n8928
                           );
   U11824 : NAND2_X2 port map( A1 => n3366, A2 => n32780, ZN => n17786);
   U14633 : NAND3_X1 port map( A1 => n9903, A2 => n24997, A3 => n9902, ZN => 
                           n4035);
   U17288 : OR2_X1 port map( A1 => n16777, A2 => n15189, Z => n4163);
   U8153 : BUF_X2 port map( I => n21860, Z => n3756);
   U4640 : INV_X2 port map( I => n497, ZN => n18742);
   U17538 : NAND2_X2 port map( A1 => n27981, A2 => n27980, ZN => n14234);
   U14489 : CLKBUF_X8 port map( I => n16051, Z => n27090);
   U637 : INV_X2 port map( I => n1104, ZN => n29115);
   U2640 : AOI21_X2 port map( A1 => n10199, A2 => n24361, B => n680, ZN => 
                           n15150);
   U23026 : NOR2_X1 port map( A1 => n8919, A2 => n16745, ZN => n14881);
   U1647 : INV_X4 port map( I => n18768, ZN => n27981);
   U276 : INV_X2 port map( I => n8125, ZN => n3165);
   U5042 : INV_X4 port map( I => n2450, ZN => n756);
   U6635 : AOI21_X2 port map( A1 => n6921, A2 => n32005, B => n6920, ZN => 
                           n6919);
   U1811 : INV_X1 port map( I => n14083, ZN => n20123);
   U11799 : NOR2_X2 port map( A1 => n15259, A2 => n15258, ZN => n14711);
   U12669 : INV_X2 port map( I => n9170, ZN => n1773);
   U20989 : NAND2_X2 port map( A1 => n19196, A2 => n3388, ZN => n19075);
   U3616 : AND2_X1 port map( A1 => n32595, A2 => n7881, Z => n10646);
   U12695 : NAND2_X1 port map( A1 => n32253, A2 => n19212, ZN => n26818);
   U2324 : NAND3_X1 port map( A1 => n28531, A2 => n25309, A3 => n25315, ZN => 
                           n28735);
   U21179 : INV_X2 port map( I => n15261, ZN => n17832);
   U1851 : BUF_X4 port map( I => n11513, Z => n8657);
   U11389 : INV_X4 port map( I => n1137, ZN => n2368);
   U23297 : NOR2_X2 port map( A1 => n28453, A2 => n7607, ZN => n28452);
   U21293 : NOR2_X1 port map( A1 => n13056, A2 => n23611, ZN => n13055);
   U15277 : INV_X2 port map( I => n25198, ZN => n25302);
   U7005 : INV_X2 port map( I => n8553, ZN => n10206);
   U5353 : NOR2_X2 port map( A1 => n10846, A2 => n14282, ZN => n7549);
   U2087 : AOI21_X2 port map( A1 => n11158, A2 => n11159, B => n11157, ZN => 
                           n4164);
   U167 : INV_X1 port map( I => n24499, ZN => n24497);
   U17441 : AOI22_X2 port map( A1 => n20285, A2 => n20284, B1 => n12263, B2 => 
                           n13589, ZN => n27478);
   U20507 : OAI22_X2 port map( A1 => n10317, A2 => n902, B1 => n10316, B2 => 
                           n1116, ZN => n10315);
   U2111 : NOR3_X2 port map( A1 => n15152, A2 => n883, A3 => n13050, ZN => 
                           n9114);
   U5802 : INV_X1 port map( I => n13704, ZN => n14253);
   U20056 : NOR2_X2 port map( A1 => n22658, A2 => n9515, ZN => n22923);
   U12622 : NOR2_X2 port map( A1 => n2023, A2 => n23859, ZN => n1731);
   U18652 : INV_X1 port map( I => n8074, ZN => n21300);
   U26358 : NAND2_X1 port map( A1 => n29212, A2 => n21540, ZN => n15820);
   U22432 : NOR2_X2 port map( A1 => n2678, A2 => n26083, ZN => n2677);
   U6011 : BUF_X2 port map( I => Key(81), Z => n16301);
   U21454 : NOR2_X1 port map( A1 => n28133, A2 => n28132, ZN => n6602);
   U5171 : BUF_X4 port map( I => n13673, Z => n13200);
   U18897 : OAI21_X2 port map( A1 => n22823, A2 => n10972, B => n22705, ZN => 
                           n10971);
   U19529 : NAND2_X2 port map( A1 => n9213, A2 => n9212, ZN => n14882);
   U9906 : NAND2_X2 port map( A1 => n12398, A2 => n19819, ZN => n12396);
   U18905 : NAND2_X1 port map( A1 => n8913, A2 => n8911, ZN => n10003);
   U15892 : AOI21_X1 port map( A1 => n27638, A2 => n29142, B => n4500, ZN => 
                           n8913);
   U8293 : OAI21_X2 port map( A1 => n21081, A2 => n21353, B => n3696, ZN => 
                           n3695);
   U3116 : INV_X2 port map( I => n15966, ZN => n18845);
   U1682 : INV_X2 port map( I => n219, ZN => n19993);
   U1947 : OAI21_X1 port map( A1 => n16954, A2 => n9793, B => n27338, ZN => 
                           n16955);
   U13354 : NAND3_X2 port map( A1 => n2621, A2 => n2622, A3 => n27755, ZN => 
                           n2620);
   U22210 : AOI22_X2 port map( A1 => n4318, A2 => n883, B1 => n25872, B2 => 
                           n13042, ZN => n14971);
   U4938 : BUF_X2 port map( I => n31161, Z => n29003);
   U12105 : NAND2_X2 port map( A1 => n9513, A2 => n7454, ZN => n9512);
   U5342 : AOI21_X2 port map( A1 => n22913, A2 => n5915, B => n803, ZN => n8943
                           );
   U21781 : BUF_X2 port map( I => n15144, Z => n14312);
   U230 : NAND2_X2 port map( A1 => n13974, A2 => n33557, ZN => n18127);
   U17790 : INV_X2 port map( I => n6693, ZN => n19456);
   U4403 : NAND2_X2 port map( A1 => n12856, A2 => n10392, ZN => n13555);
   U6906 : NAND2_X2 port map( A1 => n23047, A2 => n33007, ZN => n23048);
   U4102 : BUF_X2 port map( I => n16799, Z => n26314);
   U3787 : BUF_X2 port map( I => n5612, Z => n25990);
   U9632 : NOR2_X1 port map( A1 => n13692, A2 => n21357, ZN => n11678);
   U10122 : OAI21_X2 port map( A1 => n33098, A2 => n18698, B => n18833, ZN => 
                           n18514);
   U7178 : NAND2_X2 port map( A1 => n1145, A2 => n599, ZN => n13407);
   U9701 : NAND2_X2 port map( A1 => n30813, A2 => n926, ZN => n5469);
   U6627 : INV_X4 port map( I => n30010, ZN => n877);
   U15634 : NAND2_X2 port map( A1 => n12872, A2 => n6255, ZN => n7978);
   U4235 : CLKBUF_X4 port map( I => n7748, Z => n4236);
   U8384 : AOI21_X2 port map( A1 => n31975, A2 => n936, B => n12873, ZN => 
                           n18205);
   U5685 : OAI22_X2 port map( A1 => n9894, A2 => n33659, B1 => n29198, B2 => 
                           n9893, ZN => n23561);
   U7922 : NAND2_X2 port map( A1 => n27583, A2 => n10264, ZN => n27582);
   U18089 : NAND2_X2 port map( A1 => n10844, A2 => n17321, ZN => n27583);
   U8494 : INV_X2 port map( I => n26374, ZN => n24338);
   U7425 : INV_X2 port map( I => n27597, ZN => n19853);
   U631 : NAND3_X1 port map( A1 => n21449, A2 => n9518, A3 => n21451, ZN => 
                           n1965);
   U14814 : INV_X4 port map( I => n14931, ZN => n24955);
   U8591 : INV_X4 port map( I => n20103, ZN => n12398);
   U8180 : NOR2_X2 port map( A1 => n26955, A2 => n17701, ZN => n13603);
   U4283 : BUF_X2 port map( I => Key(156), Z => n25036);
   U10542 : NAND2_X1 port map( A1 => n13055, A2 => n8674, ZN => n26579);
   U4279 : BUF_X2 port map( I => Key(40), Z => n25476);
   U4321 : CLKBUF_X2 port map( I => Key(174), Z => n25716);
   U12281 : BUF_X2 port map( I => Key(46), Z => n16507);
   U12272 : BUF_X2 port map( I => Key(1), Z => n25545);
   U4316 : BUF_X2 port map( I => Key(141), Z => n16533);
   U4313 : CLKBUF_X2 port map( I => Key(120), Z => n16679);
   U4305 : BUF_X2 port map( I => Key(37), Z => n8548);
   U10256 : BUF_X2 port map( I => Key(100), Z => n16402);
   U8850 : BUF_X2 port map( I => Key(28), Z => n25373);
   U10218 : BUF_X2 port map( I => Key(42), Z => n24964);
   U7661 : BUF_X2 port map( I => Key(178), Z => n25728);
   U4310 : BUF_X2 port map( I => Key(180), Z => n16587);
   U6727 : BUF_X2 port map( I => Key(124), Z => n24748);
   U10205 : INV_X1 port map( I => n25720, ZN => n1428);
   U4268 : CLKBUF_X1 port map( I => n14159, Z => n8411);
   U3362 : CLKBUF_X4 port map( I => n5594, Z => n25981);
   U13955 : INV_X1 port map( I => n11605, ZN => n10095);
   U10215 : CLKBUF_X2 port map( I => n18314, Z => n18706);
   U6270 : BUF_X2 port map( I => n18674, Z => n16572);
   U21819 : INV_X1 port map( I => n25358, ZN => n15653);
   U6204 : INV_X2 port map( I => n27146, ZN => n16915);
   U3982 : CLKBUF_X2 port map( I => n18688, Z => n28675);
   U5724 : INV_X1 port map( I => n25071, ZN => n27995);
   U7606 : CLKBUF_X4 port map( I => n18293, Z => n18759);
   U18747 : NOR2_X1 port map( A1 => n732, A2 => n27691, ZN => n27690);
   U6686 : NOR2_X1 port map( A1 => n16417, A2 => n16624, ZN => n18340);
   U8740 : NOR2_X1 port map( A1 => n16328, A2 => n18482, ZN => n6252);
   U25592 : NAND2_X1 port map( A1 => n18625, A2 => n16522, ZN => n28770);
   U13211 : INV_X2 port map( I => n7134, ZN => n2283);
   U7532 : INV_X2 port map( I => n18257, ZN => n948);
   U12473 : INV_X2 port map( I => n8506, ZN => n7600);
   U10083 : OR2_X1 port map( A1 => n3388, A2 => n28528, Z => n3389);
   U1466 : NOR2_X1 port map( A1 => n16444, A2 => n19062, ZN => n19364);
   U7440 : OAI21_X1 port map( A1 => n3244, A2 => n3243, B => n19175, ZN => 
                           n3242);
   U11952 : INV_X1 port map( I => n19504, ZN => n8504);
   U3240 : CLKBUF_X2 port map( I => n19436, Z => n358);
   U14367 : INV_X1 port map( I => n33339, ZN => n16852);
   U3771 : CLKBUF_X1 port map( I => n20088, Z => n16108);
   U9948 : CLKBUF_X4 port map( I => n20102, Z => n10947);
   U11918 : INV_X1 port map( I => n4893, ZN => n8816);
   U14063 : NOR2_X1 port map( A1 => n20013, A2 => n13605, ZN => n27018);
   U11920 : BUF_X2 port map( I => n20083, Z => n16664);
   U5317 : INV_X1 port map( I => n4602, ZN => n11757);
   U19401 : NAND2_X1 port map( A1 => n28826, A2 => n8558, ZN => n27830);
   U11874 : NAND2_X1 port map( A1 => n12784, A2 => n11911, ZN => n6630);
   U24602 : NAND2_X1 port map( A1 => n30794, A2 => n28644, ZN => n19879);
   U14062 : OAI21_X1 port map( A1 => n27019, A2 => n27018, B => n20012, ZN => 
                           n19717);
   U5307 : AOI21_X1 port map( A1 => n10465, A2 => n822, B => n20076, ZN => 
                           n27846);
   U24406 : CLKBUF_X2 port map( I => n8057, Z => n28625);
   U2714 : INV_X2 port map( I => n9115, ZN => n20602);
   U1213 : NOR2_X1 port map( A1 => n32903, A2 => n14265, ZN => n14264);
   U22325 : INV_X1 port map( I => n10949, ZN => n28289);
   U19359 : NAND3_X1 port map( A1 => n26255, A2 => n13766, A3 => n13765, ZN => 
                           n1733);
   U3935 : CLKBUF_X2 port map( I => n7124, Z => n27285);
   U14827 : BUF_X2 port map( I => n21068, Z => n21243);
   U9712 : INV_X2 port map( I => n3879, ZN => n6520);
   U2448 : BUF_X2 port map( I => n21095, Z => n151);
   U1141 : INV_X1 port map( I => n26829, ZN => n21343);
   U19054 : OR2_X1 port map( A1 => n21141, A2 => n21373, Z => n27765);
   U2530 : INV_X2 port map( I => n21338, ZN => n14168);
   U5562 : INV_X2 port map( I => n12221, ZN => n17227);
   U1060 : CLKBUF_X4 port map( I => n16077, Z => n423);
   U5564 : INV_X2 port map( I => n15172, ZN => n6074);
   U3111 : INV_X2 port map( I => n29302, ZN => n15026);
   U12758 : CLKBUF_X4 port map( I => n21779, Z => n29084);
   U13059 : INV_X2 port map( I => n15863, ZN => n15864);
   U23949 : INV_X1 port map( I => n17547, ZN => n21785);
   U9530 : INV_X1 port map( I => n6231, ZN => n11924);
   U20683 : INV_X1 port map( I => n27560, ZN => n21732);
   U2903 : BUF_X2 port map( I => n8533, Z => n28848);
   U770 : BUF_X2 port map( I => n1289, Z => n28131);
   U4523 : BUF_X2 port map( I => n22597, Z => n8527);
   U796 : CLKBUF_X2 port map( I => n22362, Z => n28424);
   U4546 : NAND2_X1 port map( A1 => n9752, A2 => n9751, ZN => n10316);
   U18975 : CLKBUF_X4 port map( I => n7023, Z => n28124);
   U5082 : INV_X2 port map( I => n22645, ZN => n1292);
   U25071 : OAI21_X1 port map( A1 => n22368, A2 => n16225, B => n7023, ZN => 
                           n22369);
   U14138 : INV_X2 port map( I => n11916, ZN => n856);
   U25103 : NAND2_X1 port map( A1 => n22526, A2 => n16665, ZN => n22527);
   U15310 : NOR2_X1 port map( A1 => n27298, A2 => n5035, ZN => n9242);
   U1257 : OAI21_X1 port map( A1 => n11494, A2 => n22748, B => n3669, ZN => 
                           n4453);
   U10946 : INV_X1 port map( I => n22860, ZN => n14163);
   U6735 : NAND2_X1 port map( A1 => n26161, A2 => n26160, ZN => n2076);
   U10838 : INV_X1 port map( I => n23257, ZN => n6745);
   U4100 : INV_X2 port map( I => n9152, ZN => n14193);
   U4227 : CLKBUF_X2 port map( I => n29273, Z => n299);
   U22698 : CLKBUF_X2 port map( I => n28615, Z => n28347);
   U1760 : BUF_X4 port map( I => n8523, Z => n976);
   U4207 : BUF_X2 port map( I => n10954, Z => n29246);
   U4219 : BUF_X2 port map( I => n28765, Z => n26965);
   U10058 : AOI21_X1 port map( A1 => n26533, A2 => n23919, B => n29185, ZN => 
                           n8984);
   U7835 : NAND2_X1 port map( A1 => n23612, A2 => n16467, ZN => n23613);
   U10684 : NAND2_X1 port map( A1 => n15615, A2 => n15642, ZN => n15614);
   U21907 : NOR2_X1 port map( A1 => n23768, A2 => n27910, ZN => n12336);
   U26227 : NOR2_X1 port map( A1 => n32434, A2 => n29111, ZN => n4099);
   U17413 : NAND2_X1 port map( A1 => n10560, A2 => n8852, ZN => n8851);
   U2180 : NAND2_X1 port map( A1 => n23752, A2 => n23726, ZN => n26790);
   U1882 : CLKBUF_X4 port map( I => n13530, Z => n13268);
   U6693 : INV_X2 port map( I => n15663, ZN => n26158);
   U9029 : OAI22_X1 port map( A1 => n12022, A2 => n26247, B1 => n8665, B2 => 
                           n8663, ZN => n13144);
   U2000 : BUF_X2 port map( I => n10331, Z => n27950);
   U19559 : CLKBUF_X2 port map( I => n24753, Z => n27852);
   U1694 : CLKBUF_X4 port map( I => n91, Z => n28939);
   U4942 : INV_X1 port map( I => n25260, ZN => n11112);
   U4728 : NAND2_X1 port map( A1 => n24605, A2 => n24606, ZN => n3569);
   U4702 : INV_X1 port map( I => n12295, ZN => n25148);
   U10391 : NAND2_X1 port map( A1 => n24892, A2 => n31274, ZN => n24893);
   U15731 : NAND2_X1 port map( A1 => n14269, A2 => n14268, ZN => n12679);
   U14199 : NAND3_X1 port map( A1 => n28722, A2 => n26127, A3 => n25660, ZN => 
                           n16094);
   U10331 : INV_X2 port map( I => n2180, ZN => n15569);
   U8880 : INV_X1 port map( I => n24954, ZN => n11469);
   U5728 : BUF_X2 port map( I => n23476, Z => n29082);
   U16699 : NAND2_X2 port map( A1 => n26612, A2 => n31549, ZN => n4339);
   U1672 : INV_X2 port map( I => n26049, ZN => n5700);
   U10214 : BUF_X2 port map( I => n18873, Z => n11459);
   U13720 : BUF_X2 port map( I => n18397, Z => n18866);
   U6640 : OAI21_X1 port map( A1 => n18866, A2 => n29309, B => n18871, ZN => 
                           n18867);
   U24210 : NAND2_X1 port map( A1 => n18481, A2 => n18601, ZN => n18337);
   U24187 : INV_X1 port map( I => n18323, ZN => n18567);
   U6721 : INV_X1 port map( I => n18660, ZN => n18678);
   U5995 : BUF_X2 port map( I => n9930, Z => n9766);
   U22010 : INV_X2 port map( I => n28231, ZN => n18827);
   U4641 : INV_X1 port map( I => n469, ZN => n746);
   U5193 : INV_X2 port map( I => n4677, ZN => n8395);
   U23837 : INV_X1 port map( I => n17168, ZN => n18489);
   U4644 : INV_X1 port map( I => n10114, ZN => n18650);
   U2607 : INV_X1 port map( I => n18349, ZN => n18806);
   U10144 : NAND2_X1 port map( A1 => n34139, A2 => n18567, ZN => n4550);
   U4645 : INV_X1 port map( I => n8317, ZN => n18795);
   U6683 : NOR2_X1 port map( A1 => n1389, A2 => n4925, ZN => n26156);
   U18750 : INV_X1 port map( I => n10578, ZN => n27691);
   U6667 : NOR2_X1 port map( A1 => n16417, A2 => n12120, ZN => n18778);
   U8822 : INV_X1 port map( I => n4259, ZN => n17266);
   U13643 : NAND2_X1 port map( A1 => n16522, A2 => n18774, ZN => n26962);
   U10104 : NAND2_X1 port map( A1 => n10669, A2 => n9296, ZN => n10326);
   U3688 : INV_X1 port map( I => n17223, ZN => n17224);
   U985 : INV_X1 port map( I => n18860, ZN => n18532);
   U24372 : NAND2_X1 port map( A1 => n30371, A2 => n785, ZN => n18817);
   U6712 : INV_X1 port map( I => n18357, ZN => n18895);
   U8777 : NAND2_X1 port map( A1 => n10579, A2 => n2990, ZN => n6457);
   U24299 : OAI21_X1 port map( A1 => n18481, A2 => n18601, B => n18602, ZN => 
                           n18480);
   U13783 : AOI21_X1 port map( A1 => n955, A2 => n16995, B => n1184, ZN => 
                           n5458);
   U2233 : NAND3_X1 port map( A1 => n18332, A2 => n18489, A3 => n6256, ZN => 
                           n18334);
   U21122 : NAND2_X1 port map( A1 => n16249, A2 => n18822, ZN => n13946);
   U24356 : NOR2_X1 port map( A1 => n18730, A2 => n18846, ZN => n18732);
   U8787 : NOR2_X1 port map( A1 => n18759, A2 => n27940, ZN => n18606);
   U5189 : NAND2_X1 port map( A1 => n18532, A2 => n18588, ZN => n17599);
   U2237 : NAND3_X1 port map( A1 => n1659, A2 => n5700, A3 => n46, ZN => n7319)
                           ;
   U16162 : AOI22_X1 port map( A1 => n16196, A2 => n18648, B1 => n18373, B2 => 
                           n18804, ZN => n27237);
   U10098 : NOR2_X1 port map( A1 => n14843, A2 => n11397, ZN => n11396);
   U10140 : OAI21_X1 port map( A1 => n28010, A2 => n959, B => n27958, ZN => 
                           n16018);
   U5174 : NOR2_X1 port map( A1 => n18532, A2 => n18588, ZN => n18739);
   U10183 : INV_X1 port map( I => n12120, ZN => n18339);
   U2682 : INV_X1 port map( I => n10264, ZN => n18750);
   U9648 : NAND2_X1 port map( A1 => n18846, A2 => n18847, ZN => n18410);
   U8737 : OAI21_X1 port map( A1 => n6579, A2 => n18802, B => n8395, ZN => 
                           n4472);
   U6899 : AOI22_X1 port map( A1 => n18340, A2 => n18339, B1 => n1430, B2 => 
                           n6215, ZN => n26176);
   U24206 : OAI21_X1 port map( A1 => n27129, A2 => n28987, B => n18556, ZN => 
                           n18329);
   U7552 : NOR2_X1 port map( A1 => n11864, A2 => n18559, ZN => n18330);
   U2620 : OAI21_X1 port map( A1 => n17113, A2 => n12013, B => n18808, ZN => 
                           n2680);
   U7562 : NAND2_X1 port map( A1 => n18812, A2 => n2990, ZN => n2683);
   U15208 : NOR2_X1 port map( A1 => n15136, A2 => n4008, ZN => n18260);
   U1314 : BUF_X2 port map( I => n10579, Z => n3429);
   U8491 : BUF_X2 port map( I => n19049, Z => n28705);
   U6670 : AOI21_X1 port map( A1 => n17360, A2 => n18587, B => n18863, ZN => 
                           n13025);
   U3971 : INV_X2 port map( I => n9677, ZN => n13568);
   U18050 : NOR2_X1 port map( A1 => n19011, A2 => n5119, ZN => n7110);
   U21515 : INV_X1 port map( I => n14811, ZN => n18426);
   U19805 : NAND2_X1 port map( A1 => n9787, A2 => n19224, ZN => n12505);
   U5484 : NAND2_X1 port map( A1 => n1053, A2 => n31451, ZN => n18454);
   U22187 : INV_X2 port map( I => n19048, ZN => n16669);
   U7495 : INV_X1 port map( I => n16699, ZN => n19334);
   U15115 : NAND2_X1 port map( A1 => n13037, A2 => n13035, ZN => n27131);
   U21485 : NOR2_X1 port map( A1 => n13200, A2 => n19118, ZN => n14424);
   U22712 : INV_X1 port map( I => n19033, ZN => n4102);
   U7477 : NAND3_X1 port map( A1 => n7435, A2 => n7434, A3 => n1047, ZN => 
                           n7439);
   U7450 : AOI22_X1 port map( A1 => n9424, A2 => n9423, B1 => n18068, B2 => 
                           n26830, ZN => n9422);
   U5501 : BUF_X2 port map( I => n18980, Z => n16740);
   U16708 : NOR3_X1 port map( A1 => n18930, A2 => n16444, A3 => n1053, ZN => 
                           n18284);
   U3973 : BUF_X2 port map( I => n2581, Z => n26181);
   U13526 : AOI21_X1 port map( A1 => n15074, A2 => n15073, B => n17986, ZN => 
                           n14259);
   U5233 : NAND3_X1 port map( A1 => n19087, A2 => n19089, A3 => n1384, ZN => 
                           n10868);
   U21457 : NOR2_X1 port map( A1 => n19215, A2 => n2901, ZN => n28132);
   U900 : OAI21_X1 port map( A1 => n10013, A2 => n11080, B => n4017, ZN => 
                           n18910);
   U5481 : NOR2_X1 port map( A1 => n19332, A2 => n8335, ZN => n5162);
   U7999 : NOR2_X1 port map( A1 => n19359, A2 => n19356, ZN => n15629);
   U19389 : NAND2_X1 port map( A1 => n1180, A2 => n19255, ZN => n8910);
   U5490 : INV_X1 port map( I => n19080, ZN => n19171);
   U7509 : NOR2_X1 port map( A1 => n19116, A2 => n19330, ZN => n3784);
   U10330 : INV_X1 port map( I => n19148, ZN => n26554);
   U12769 : NAND3_X1 port map( A1 => n3365, A2 => n745, A3 => n3360, ZN => 
                           n1870);
   U7489 : AOI21_X1 port map( A1 => n32064, A2 => n15120, B => n16916, ZN => 
                           n19162);
   U9991 : INV_X1 port map( I => n12996, ZN => n5710);
   U21998 : INV_X1 port map( I => n12830, ZN => n12567);
   U5252 : INV_X1 port map( I => n19128, ZN => n15378);
   U12039 : INV_X1 port map( I => n11074, ZN => n17678);
   U5941 : NAND2_X1 port map( A1 => n12707, A2 => n16669, ZN => n3822);
   U21514 : NAND2_X1 port map( A1 => n16592, A2 => n16591, ZN => n18268);
   U5924 : NAND3_X1 port map( A1 => n18967, A2 => n11085, A3 => n19165, ZN => 
                           n11800);
   U20394 : AOI21_X1 port map( A1 => n19280, A2 => n32908, B => n26830, ZN => 
                           n19282);
   U2876 : NAND3_X1 port map( A1 => n34005, A2 => n29715, A3 => n17311, ZN => 
                           n19173);
   U12044 : OAI21_X1 port map( A1 => n18983, A2 => n19128, B => n18963, ZN => 
                           n18966);
   U15672 : OAI21_X1 port map( A1 => n764, A2 => n25985, B => n9677, ZN => 
                           n9709);
   U15974 : NOR2_X1 port map( A1 => n1378, A2 => n29146, ZN => n12532);
   U6188 : INV_X1 port map( I => n1180, ZN => n26288);
   U8621 : OAI21_X1 port map( A1 => n1382, A2 => n19004, B => n19210, ZN => 
                           n18942);
   U12330 : AOI22_X1 port map( A1 => n13495, A2 => n19116, B1 => n879, B2 => 
                           n5162, ZN => n28003);
   U19512 : INV_X1 port map( I => n19151, ZN => n9176);
   U18141 : NAND3_X1 port map( A1 => n16354, A2 => n19291, A3 => n7251, ZN => 
                           n19204);
   U7668 : BUF_X2 port map( I => Key(160), Z => n25054);
   U9966 : INV_X1 port map( I => n16727, ZN => n3076);
   U2889 : INV_X1 port map( I => n2073, ZN => n2761);
   U878 : INV_X1 port map( I => n2483, ZN => n6115);
   U4273 : BUF_X2 port map( I => Key(122), Z => n25358);
   U11959 : INV_X1 port map( I => n19644, ZN => n1916);
   U6100 : BUF_X2 port map( I => Key(45), Z => n25783);
   U4278 : BUF_X2 port map( I => Key(99), Z => n25554);
   U847 : INV_X1 port map( I => n20067, ZN => n823);
   U4925 : NAND2_X1 port map( A1 => n823, A2 => n19947, ZN => n28021);
   U19508 : INV_X2 port map( I => n10934, ZN => n14210);
   U8377 : INV_X2 port map( I => n4060, ZN => n5433);
   U3238 : INV_X1 port map( I => n577, ZN => n1041);
   U825 : INV_X2 port map( I => n17688, ZN => n20110);
   U24625 : INV_X1 port map( I => n29981, ZN => n19976);
   U5892 : INV_X2 port map( I => n1164, ZN => n7920);
   U2496 : INV_X2 port map( I => n16811, ZN => n16812);
   U837 : INV_X2 port map( I => n29253, ZN => n1036);
   U863 : INV_X1 port map( I => n26774, ZN => n875);
   U5347 : OAI22_X1 port map( A1 => n12038, A2 => n25997, B1 => n13747, B2 => 
                           n10947, ZN => n17371);
   U833 : INV_X1 port map( I => n20109, ZN => n20035);
   U9941 : INV_X1 port map( I => n16193, ZN => n20012);
   U16819 : NAND2_X1 port map( A1 => n5707, A2 => n19987, ZN => n14440);
   U7388 : NAND2_X1 port map( A1 => n3626, A2 => n20076, ZN => n3663);
   U5277 : NAND2_X1 port map( A1 => n12008, A2 => n10086, ZN => n8946);
   U11780 : AOI21_X1 port map( A1 => n19861, A2 => n7923, B => n1164, ZN => 
                           n7921);
   U21988 : INV_X2 port map( I => n19986, ZN => n28219);
   U20149 : INV_X1 port map( I => n20134, ZN => n20132);
   U7424 : INV_X1 port map( I => n3486, ZN => n3530);
   U11848 : NAND2_X1 port map( A1 => n16346, A2 => n17243, ZN => n3128);
   U8504 : NOR2_X1 port map( A1 => n9876, A2 => n8301, ZN => n2933);
   U13885 : NOR3_X1 port map( A1 => n20007, A2 => n20008, A3 => n20009, ZN => 
                           n2930);
   U5299 : NAND2_X1 port map( A1 => n1036, A2 => n31161, ZN => n8033);
   U8550 : OAI21_X1 port map( A1 => n5871, A2 => n5869, B => n31468, ZN => 
                           n3292);
   U9937 : INV_X1 port map( I => n4215, ZN => n17389);
   U20249 : NAND2_X1 port map( A1 => n584, A2 => n14559, ZN => n11475);
   U11804 : NAND2_X1 port map( A1 => n26088, A2 => n30794, ZN => n5288);
   U14929 : NAND2_X1 port map( A1 => n20132, A2 => n16461, ZN => n5931);
   U19858 : NOR2_X1 port map( A1 => n13987, A2 => n10241, ZN => n13986);
   U7385 : NAND2_X1 port map( A1 => n15278, A2 => n1166, ZN => n20292);
   U5338 : AND2_X1 port map( A1 => n10831, A2 => n33627, Z => n19952);
   U9898 : NOR2_X1 port map( A1 => n20154, A2 => n27097, ZN => n16307);
   U6528 : NOR2_X1 port map( A1 => n4215, A2 => n17243, ZN => n12078);
   U19422 : AOI21_X1 port map( A1 => n17243, A2 => n4233, B => n4215, ZN => 
                           n9139);
   U14805 : NAND3_X1 port map( A1 => n20100, A2 => n12895, A3 => n19990, ZN => 
                           n17035);
   U819 : OAI21_X1 port map( A1 => n29281, A2 => n25997, B => n12038, ZN => 
                           n13954);
   U5357 : NAND2_X1 port map( A1 => n19952, A2 => n19856, ZN => n12194);
   U11802 : OAI21_X1 port map( A1 => n32559, A2 => n13058, B => n19823, ZN => 
                           n10478);
   U8529 : NOR2_X1 port map( A1 => n19884, A2 => n19886, ZN => n19421);
   U1348 : NOR2_X1 port map( A1 => n12408, A2 => n3626, ZN => n27802);
   U21532 : NAND2_X1 port map( A1 => n17785, A2 => n20010, ZN => n17784);
   U2404 : INV_X1 port map( I => n20485, ZN => n1346);
   U806 : NAND2_X1 port map( A1 => n20006, A2 => n20078, ZN => n13107);
   U15780 : NAND2_X1 port map( A1 => n19998, A2 => n28219, ZN => n4367);
   U13038 : NAND3_X1 port map( A1 => n20100, A2 => n29216, A3 => n29944, ZN => 
                           n20623);
   U1310 : AOI21_X1 port map( A1 => n19986, A2 => n25997, B => n11521, ZN => 
                           n4368);
   U21264 : INV_X1 port map( I => n20312, ZN => n20578);
   U4594 : INV_X2 port map( I => n20492, ZN => n20494);
   U1298 : INV_X1 port map( I => n8374, ZN => n20525);
   U771 : INV_X2 port map( I => n31504, ZN => n12169);
   U22617 : NAND2_X1 port map( A1 => n17947, A2 => n20485, ZN => n17532);
   U23017 : NOR2_X1 port map( A1 => n20268, A2 => n14863, ZN => n20269);
   U3325 : INV_X1 port map( I => n9320, ZN => n1028);
   U1242 : INV_X2 port map( I => n15027, ZN => n27771);
   U8444 : NOR2_X1 port map( A1 => n935, A2 => n29628, ZN => n17414);
   U19867 : NAND2_X1 port map( A1 => n27105, A2 => n30643, ZN => n20347);
   U3199 : NAND2_X1 port map( A1 => n20268, A2 => n5781, ZN => n5670);
   U2892 : BUF_X2 port map( I => n20267, Z => n266);
   U6503 : NAND2_X1 port map( A1 => n9320, A2 => n14436, ZN => n20257);
   U22722 : BUF_X2 port map( I => n14049, Z => n28357);
   U14587 : INV_X2 port map( I => n5748, ZN => n782);
   U6504 : NAND2_X1 port map( A1 => n20268, A2 => n20210, ZN => n5782);
   U4830 : NAND2_X1 port map( A1 => n15169, A2 => n20590, ZN => n28893);
   U23091 : INV_X2 port map( I => n2928, ZN => n28414);
   U11727 : NOR2_X1 port map( A1 => n12771, A2 => n9484, ZN => n5061);
   U16049 : AOI21_X1 port map( A1 => n30971, A2 => n31873, B => n20379, ZN => 
                           n20380);
   U23485 : NAND3_X1 port map( A1 => n28893, A2 => n31967, A3 => n15824, ZN => 
                           n28485);
   U8414 : NOR2_X1 port map( A1 => n7978, A2 => n936, ZN => n12873);
   U16113 : OAI21_X1 port map( A1 => n20347, A2 => n26730, B => n27225, ZN => 
                           n27227);
   U26129 : INV_X1 port map( I => n17947, ZN => n17896);
   U24715 : NAND2_X1 port map( A1 => n1159, A2 => n30987, ZN => n20475);
   U13112 : NOR2_X1 port map( A1 => n31804, A2 => n31533, ZN => n5993);
   U9953 : INV_X1 port map( I => n31471, ZN => n1354);
   U14535 : INV_X1 port map( I => n3644, ZN => n12407);
   U22901 : AOI21_X1 port map( A1 => n15042, A2 => n15043, B => n28840, ZN => 
                           n15041);
   U8390 : OAI22_X1 port map( A1 => n29972, A2 => n20426, B1 => n16146, B2 => 
                           n20427, ZN => n1930);
   U15874 : NOR2_X1 port map( A1 => n1354, A2 => n4468, ZN => n4471);
   U23867 : NAND2_X1 port map( A1 => n817, A2 => n31804, ZN => n17270);
   U12457 : NAND3_X1 port map( A1 => n1351, A2 => n11312, A3 => n1349, ZN => 
                           n20407);
   U24661 : OAI21_X1 port map( A1 => n20202, A2 => n20201, B => n27887, ZN => 
                           n20203);
   U3535 : NOR2_X1 port map( A1 => n5003, A2 => n32504, ZN => n20164);
   U11737 : NOR2_X1 port map( A1 => n2965, A2 => n1159, ZN => n2764);
   U24658 : INV_X1 port map( I => n20462, ZN => n20187);
   U9719 : INV_X1 port map( I => n9303, ZN => n20871);
   U19160 : INV_X1 port map( I => n20755, ZN => n12674);
   U2704 : INV_X1 port map( I => n20939, ZN => n21270);
   U19708 : NOR2_X1 port map( A1 => n7007, A2 => n28190, ZN => n6303);
   U5115 : INV_X2 port map( I => n21170, ZN => n14803);
   U9718 : INV_X1 port map( I => n11733, ZN => n1148);
   U4754 : INV_X1 port map( I => n34157, ZN => n21167);
   U8306 : NOR2_X1 port map( A1 => n21398, A2 => n32625, ZN => n21206);
   U6435 : NOR2_X1 port map( A1 => n5049, A2 => n29255, ZN => n5047);
   U21135 : NOR2_X1 port map( A1 => n21165, A2 => n14803, ZN => n21086);
   U7165 : INV_X2 port map( I => n21428, ZN => n21341);
   U2645 : INV_X1 port map( I => n2118, ZN => n8267);
   U11538 : INV_X1 port map( I => n28190, ZN => n13509);
   U20930 : NOR2_X1 port map( A1 => n1334, A2 => n21270, ZN => n12243);
   U9698 : NAND2_X1 port map( A1 => n5141, A2 => n14168, ZN => n21340);
   U15904 : NAND3_X1 port map( A1 => n28502, A2 => n21079, A3 => n4518, ZN => 
                           n20938);
   U11542 : INV_X1 port map( I => n15751, ZN => n17093);
   U7185 : NOR2_X1 port map( A1 => n17640, A2 => n3106, ZN => n7378);
   U8254 : NOR2_X1 port map( A1 => n6451, A2 => n1736, ZN => n4569);
   U14558 : OAI21_X1 port map( A1 => n11151, A2 => n27842, B => n21217, ZN => 
                           n11150);
   U13282 : NAND2_X1 port map( A1 => n7196, A2 => n6520, ZN => n2568);
   U8383 : NOR2_X1 port map( A1 => n28502, A2 => n16933, ZN => n16484);
   U4751 : CLKBUF_X2 port map( I => n21170, Z => n26861);
   U8287 : NOR2_X1 port map( A1 => n21212, A2 => n6408, ZN => n18213);
   U24830 : INV_X1 port map( I => n31909, ZN => n21093);
   U5413 : NAND2_X1 port map( A1 => n21405, A2 => n4989, ZN => n4988);
   U8246 : OAI22_X1 port map( A1 => n20933, A2 => n21080, B1 => n21365, B2 => 
                           n21183, ZN => n13265);
   U632 : OAI21_X1 port map( A1 => n9454, A2 => n7822, B => n17455, ZN => n9453
                           );
   U16203 : NAND2_X1 port map( A1 => n8175, A2 => n21434, ZN => n27249);
   U9642 : NOR2_X1 port map( A1 => n20662, A2 => n4518, ZN => n4283);
   U7129 : OAI21_X1 port map( A1 => n8012, A2 => n16639, B => n7526, ZN => 
                           n21437);
   U15029 : NAND2_X1 port map( A1 => n7123, A2 => n7120, ZN => n5843);
   U3913 : NAND2_X1 port map( A1 => n2575, A2 => n21849, ZN => n26341);
   U23415 : NOR3_X1 port map( A1 => n21408, A2 => n4119, A3 => n30755, ZN => 
                           n15872);
   U9593 : AOI21_X1 port map( A1 => n7148, A2 => n8604, B => n8010, ZN => n6427
                           );
   U1032 : NOR2_X1 port map( A1 => n13133, A2 => n1136, ZN => n26175);
   U24342 : BUF_X2 port map( I => n21665, Z => n28618);
   U6368 : NAND3_X1 port map( A1 => n16577, A2 => n13133, A3 => n1312, ZN => 
                           n21667);
   U6399 : INV_X2 port map( I => n21463, ZN => n918);
   U14233 : AOI21_X1 port map( A1 => n15813, A2 => n10401, B => n11890, ZN => 
                           n27053);
   U597 : INV_X1 port map( I => n28232, ZN => n1328);
   U24913 : AOI21_X1 port map( A1 => n21690, A2 => n21859, B => n21857, ZN => 
                           n21538);
   U1016 : NAND3_X1 port map( A1 => n1328, A2 => n15772, A3 => n21811, ZN => 
                           n8174);
   U11968 : NOR2_X1 port map( A1 => n21709, A2 => n30441, ZN => n27383);
   U3649 : NAND2_X1 port map( A1 => n8276, A2 => n21707, ZN => n9055);
   U23200 : NOR2_X1 port map( A1 => n30885, A2 => n27635, ZN => n17347);
   U1015 : NOR2_X1 port map( A1 => n21629, A2 => n21628, ZN => n27991);
   U11957 : NOR2_X1 port map( A1 => n31954, A2 => n27178, ZN => n26731);
   U8183 : BUF_X2 port map( I => n8602, Z => n4331);
   U8196 : INV_X2 port map( I => n21779, ZN => n21781);
   U3251 : INV_X1 port map( I => n6489, ZN => n21853);
   U557 : NOR2_X1 port map( A1 => n21806, A2 => n6483, ZN => n279);
   U11404 : NAND2_X1 port map( A1 => n21690, A2 => n29523, ZN => n2708);
   U11337 : NAND2_X1 port map( A1 => n21164, A2 => n16577, ZN => n12994);
   U3590 : INV_X1 port map( I => n21715, ZN => n911);
   U4165 : INV_X1 port map( I => n14095, ZN => n21775);
   U4633 : INV_X1 port map( I => n7502, ZN => n28665);
   U22789 : NOR2_X1 port map( A1 => n30440, A2 => n31309, ZN => n21934);
   U940 : NAND3_X1 port map( A1 => n17644, A2 => n3756, A3 => n21857, ZN => 
                           n28159);
   U9505 : NAND3_X1 port map( A1 => n21800, A2 => n21801, A3 => n21799, ZN => 
                           n15640);
   U18456 : NAND2_X1 port map( A1 => n21678, A2 => n28203, ZN => n27630);
   U23082 : OAI21_X1 port map( A1 => n17472, A2 => n15026, B => n16194, ZN => 
                           n21495);
   U11322 : AOI21_X1 port map( A1 => n12102, A2 => n21686, B => n26513, ZN => 
                           n10490);
   U3432 : NAND2_X1 port map( A1 => n9119, A2 => n21655, ZN => n21936);
   U21170 : NAND2_X1 port map( A1 => n15091, A2 => n31085, ZN => n14012);
   U5396 : NOR2_X1 port map( A1 => n21622, A2 => n28387, ZN => n21561);
   U13782 : NAND2_X1 port map( A1 => n10028, A2 => n27619, ZN => n26979);
   U11282 : NOR2_X1 port map( A1 => n17164, A2 => n15319, ZN => n16164);
   U13910 : OAI21_X1 port map( A1 => n12626, A2 => n9076, B => n11619, ZN => 
                           n9088);
   U3902 : NAND2_X1 port map( A1 => n21819, A2 => n26904, ZN => n27103);
   U9515 : AOI21_X1 port map( A1 => n9666, A2 => n15091, B => n28618, ZN => 
                           n13804);
   U22785 : NAND2_X1 port map( A1 => n21934, A2 => n915, ZN => n21935);
   U524 : INV_X1 port map( I => n22172, ZN => n4723);
   U4839 : INV_X1 port map( I => n32055, ZN => n9065);
   U6356 : INV_X1 port map( I => n11100, ZN => n22543);
   U6318 : NAND2_X1 port map( A1 => n1122, A2 => n31931, ZN => n11575);
   U2572 : INV_X2 port map( I => n22543, ZN => n1124);
   U23842 : NAND2_X1 port map( A1 => n28472, A2 => n16627, ZN => n22571);
   U21002 : NAND2_X1 port map( A1 => n15752, A2 => n29451, ZN => n15008);
   U8027 : OAI21_X1 port map( A1 => n4055, A2 => n4054, B => n8527, ZN => n7610
                           );
   U9350 : NOR2_X1 port map( A1 => n18098, A2 => n12076, ZN => n17263);
   U20086 : NAND2_X1 port map( A1 => n22330, A2 => n14376, ZN => n10317);
   U782 : NOR2_X1 port map( A1 => n998, A2 => n22330, ZN => n17132);
   U3597 : INV_X2 port map( I => n22626, ZN => n1117);
   U4141 : INV_X1 port map( I => n8409, ZN => n22586);
   U4132 : INV_X1 port map( I => n30668, ZN => n1282);
   U492 : INV_X2 port map( I => n16205, ZN => n22689);
   U25106 : OAI21_X1 port map( A1 => n22565, A2 => n22561, B => n22560, ZN => 
                           n22566);
   U430 : NAND2_X1 port map( A1 => n15229, A2 => n22476, ZN => n13534);
   U724 : NAND3_X1 port map( A1 => n26878, A2 => n27378, A3 => n996, ZN => 
                           n26178);
   U17275 : OAI21_X1 port map( A1 => n22610, A2 => n29336, B => n22631, ZN => 
                           n22613);
   U8005 : NOR2_X1 port map( A1 => n22531, A2 => n9234, ZN => n9777);
   U18681 : NOR2_X1 port map( A1 => n7957, A2 => n1124, ZN => n8136);
   U21232 : OAI21_X1 port map( A1 => n17960, A2 => n16375, B => n1728, ZN => 
                           n22526);
   U9386 : INV_X1 port map( I => n9272, ZN => n8348);
   U2334 : NOR2_X1 port map( A1 => n16170, A2 => n25, ZN => n26862);
   U11069 : NAND2_X1 port map( A1 => n1113, A2 => n22923, ZN => n3854);
   U21922 : NAND2_X1 port map( A1 => n1294, A2 => n26884, ZN => n28206);
   U9438 : NAND2_X1 port map( A1 => n9271, A2 => n9234, ZN => n9270);
   U19882 : OAI22_X1 port map( A1 => n13417, A2 => n9913, B1 => n22667, B2 => 
                           n29078, ZN => n22723);
   U14894 : INV_X2 port map( I => n4908, ZN => n724);
   U6546 : OAI21_X1 port map( A1 => n26144, A2 => n26660, B => n14728, ZN => 
                           n26394);
   U9367 : AOI21_X1 port map( A1 => n8595, A2 => n30641, B => n4300, ZN => 
                           n4299);
   U4529 : NAND2_X1 port map( A1 => n22392, A2 => n22546, ZN => n14024);
   U1044 : NAND2_X1 port map( A1 => n22407, A2 => n22429, ZN => n17627);
   U15007 : INV_X1 port map( I => n23072, ZN => n8683);
   U6949 : NOR2_X1 port map( A1 => n22878, A2 => n31437, ZN => n2169);
   U9236 : NOR2_X1 port map( A1 => n14131, A2 => n2635, ZN => n6285);
   U9322 : INV_X1 port map( I => n6798, ZN => n1107);
   U590 : INV_X1 port map( I => n31637, ZN => n13778);
   U7972 : INV_X2 port map( I => n849, ZN => n7181);
   U6287 : INV_X1 port map( I => n5915, ZN => n23073);
   U615 : INV_X1 port map( I => n22968, ZN => n23083);
   U16802 : NOR2_X1 port map( A1 => n27622, A2 => n3163, ZN => n13917);
   U25193 : NAND3_X1 port map( A1 => n23070, A2 => n10641, A3 => n23069, ZN => 
                           n23071);
   U6261 : NOR2_X1 port map( A1 => n26724, A2 => n23104, ZN => n5972);
   U21545 : OAI21_X1 port map( A1 => n18241, A2 => n22916, B => n27090, ZN => 
                           n18047);
   U4409 : INV_X1 port map( I => n28214, ZN => n27409);
   U26084 : NOR2_X1 port map( A1 => n22798, A2 => n23053, ZN => n23050);
   U1427 : NAND2_X1 port map( A1 => n641, A2 => n11268, ZN => n6227);
   U16265 : NAND2_X1 port map( A1 => n32091, A2 => n10296, ZN => n22441);
   U19331 : NAND3_X1 port map( A1 => n15852, A2 => n15851, A3 => n30960, ZN => 
                           n13598);
   U22109 : NOR2_X1 port map( A1 => n22872, A2 => n31861, ZN => n12824);
   U14459 : OAI22_X1 port map( A1 => n10360, A2 => n3570, B1 => n3891, B2 => 
                           n12586, ZN => n22714);
   U10853 : INV_X1 port map( I => n15941, ZN => n2974);
   U10860 : INV_X1 port map( I => n12716, ZN => n3282);
   U312 : INV_X1 port map( I => n23475, ZN => n6262);
   U458 : INV_X1 port map( I => n28811, ZN => n662);
   U9134 : OAI21_X1 port map( A1 => n11887, A2 => n11933, B => n3004, ZN => 
                           n10069);
   U7887 : INV_X1 port map( I => n23719, ZN => n23919);
   U6218 : INV_X1 port map( I => n23567, ZN => n23849);
   U8286 : INV_X1 port map( I => n23683, ZN => n23681);
   U25891 : NAND2_X1 port map( A1 => n32998, A2 => n11933, ZN => n15490);
   U5789 : NAND2_X1 port map( A1 => n23491, A2 => n23712, ZN => n17520);
   U477 : INV_X1 port map( I => n10954, ZN => n11968);
   U2850 : OR2_X1 port map( A1 => n28611, A2 => n8166, Z => n8674);
   U5695 : NOR2_X1 port map( A1 => n23713, A2 => n23889, ZN => n23842);
   U413 : INV_X2 port map( I => n756, ZN => n28510);
   U10532 : NAND2_X1 port map( A1 => n23813, A2 => n663, ZN => n23692);
   U9216 : INV_X2 port map( I => n27455, ZN => n23752);
   U9199 : INV_X1 port map( I => n11567, ZN => n8095);
   U4113 : INV_X1 port map( I => n9430, ZN => n15912);
   U19075 : AND2_X1 port map( A1 => n7022, A2 => n2839, Z => n14092);
   U20458 : NOR2_X1 port map( A1 => n23864, A2 => n23527, ZN => n11131);
   U7815 : NAND2_X1 port map( A1 => n23894, A2 => n29068, ZN => n6249);
   U9180 : NAND2_X1 port map( A1 => n7915, A2 => n23778, ZN => n11393);
   U25320 : INV_X1 port map( I => n23646, ZN => n23647);
   U3881 : NOR2_X1 port map( A1 => n707, A2 => n8370, ZN => n655);
   U18362 : AOI21_X1 port map( A1 => n10193, A2 => n34008, B => n23897, ZN => 
                           n10560);
   U5831 : NAND2_X1 port map( A1 => n17520, A2 => n17234, ZN => n11491);
   U5711 : INV_X1 port map( I => n976, ZN => n1249);
   U10819 : NOR2_X1 port map( A1 => n13549, A2 => n27219, ZN => n8473);
   U6856 : NOR2_X1 port map( A1 => n8544, A2 => n14207, ZN => n11309);
   U404 : INV_X2 port map( I => n15423, ZN => n23850);
   U9139 : NAND2_X1 port map( A1 => n978, A2 => n8273, ZN => n15351);
   U4790 : INV_X1 port map( I => n14092, ZN => n23651);
   U2110 : OAI21_X1 port map( A1 => n13544, A2 => n13578, B => n17906, ZN => 
                           n7613);
   U25328 : NAND2_X1 port map( A1 => n11192, A2 => n16337, ZN => n28744);
   U6895 : NAND3_X1 port map( A1 => n16467, A2 => n846, A3 => n27219, ZN => 
                           n7075);
   U16858 : NAND3_X1 port map( A1 => n847, A2 => n23573, A3 => n5759, ZN => 
                           n23574);
   U21319 : NAND2_X1 port map( A1 => n23832, A2 => n23912, ZN => n17398);
   U21050 : NOR2_X1 port map( A1 => n8408, A2 => n17895, ZN => n17806);
   U2242 : NAND2_X1 port map( A1 => n32711, A2 => n654, ZN => n26384);
   U21292 : INV_X1 port map( I => n23923, ZN => n16118);
   U375 : INV_X1 port map( I => n32308, ZN => n26383);
   U8694 : INV_X1 port map( I => n26392, ZN => n26391);
   U348 : NOR2_X1 port map( A1 => n9797, A2 => n14207, ZN => n9769);
   U10741 : NAND2_X1 port map( A1 => n17618, A2 => n13503, ZN => n3484);
   U24025 : NOR2_X1 port map( A1 => n17807, A2 => n17806, ZN => n17805);
   U1627 : INV_X1 port map( I => n9919, ZN => n10530);
   U218 : INV_X1 port map( I => n6911, ZN => n24312);
   U3087 : CLKBUF_X2 port map( I => n24299, Z => n319);
   U26435 : BUF_X2 port map( I => n24314, Z => n7503);
   U6831 : INV_X2 port map( I => n3205, ZN => n9323);
   U204 : INV_X1 port map( I => n5199, ZN => n24245);
   U1655 : INV_X1 port map( I => n9342, ZN => n14252);
   U9113 : INV_X1 port map( I => n16799, ZN => n1089);
   U8289 : NAND2_X1 port map( A1 => n24243, A2 => n24242, ZN => n1480);
   U8049 : NAND2_X1 port map( A1 => n1089, A2 => n14619, ZN => n5615);
   U9049 : AOI21_X1 port map( A1 => n796, A2 => n10226, B => n970, ZN => n9282)
                           ;
   U20904 : NOR2_X1 port map( A1 => n24305, A2 => n24197, ZN => n16901);
   U2309 : NAND2_X1 port map( A1 => n27159, A2 => n24094, ZN => n13239);
   U9043 : NOR2_X1 port map( A1 => n16985, A2 => n1245, ZN => n5616);
   U4097 : INV_X1 port map( I => n14725, ZN => n27550);
   U15179 : INV_X1 port map( I => n3148, ZN => n3038);
   U9027 : NAND2_X1 port map( A1 => n24061, A2 => n10651, ZN => n11342);
   U4777 : NOR2_X1 port map( A1 => n3483, A2 => n24193, ZN => n24057);
   U3528 : NAND2_X1 port map( A1 => n27117, A2 => n24168, ZN => n13306);
   U4779 : NOR2_X1 port map( A1 => n10033, A2 => n24201, ZN => n7669);
   U14171 : OAI21_X1 port map( A1 => n7809, A2 => n30280, B => n16651, ZN => 
                           n5937);
   U5263 : NAND3_X1 port map( A1 => n24211, A2 => n24213, A3 => n24209, ZN => 
                           n6990);
   U8171 : NAND3_X1 port map( A1 => n24322, A2 => n29785, A3 => n24209, ZN => 
                           n6817);
   U10544 : NAND2_X1 port map( A1 => n28120, A2 => n13048, ZN => n13046);
   U10615 : INV_X1 port map( I => n11346, ZN => n10428);
   U15680 : NOR2_X1 port map( A1 => n24097, A2 => n24096, ZN => n5377);
   U7785 : NOR2_X1 port map( A1 => n14443, A2 => n17404, ZN => n7105);
   U2256 : OAI21_X1 port map( A1 => n32036, A2 => n7669, B => n24008, ZN => 
                           n7668);
   U7810 : NAND2_X1 port map( A1 => n8058, A2 => n24106, ZN => n23665);
   U3284 : NAND2_X1 port map( A1 => n11342, A2 => n11341, ZN => n11340);
   U14084 : NAND2_X1 port map( A1 => n6001, A2 => n27026, ZN => n12693);
   U18424 : NAND3_X1 port map( A1 => n1244, A2 => n29010, A3 => n24216, ZN => 
                           n10175);
   U23247 : NAND2_X1 port map( A1 => n23748, A2 => n27184, ZN => n24018);
   U9069 : NAND2_X1 port map( A1 => n10188, A2 => n31355, ZN => n8000);
   U3711 : NAND3_X1 port map( A1 => n24322, A2 => n13268, A3 => n29785, ZN => 
                           n24324);
   U25404 : NAND2_X1 port map( A1 => n24213, A2 => n13268, ZN => n24214);
   U1058 : NAND2_X1 port map( A1 => n2852, A2 => n29567, ZN => n2849);
   U11550 : AOI21_X1 port map( A1 => n14336, A2 => n24317, B => n32298, ZN => 
                           n2156);
   U22969 : NAND3_X1 port map( A1 => n1089, A2 => n12054, A3 => n14745, ZN => 
                           n15224);
   U10526 : INV_X1 port map( I => n24442, ZN => n10070);
   U173 : OR2_X1 port map( A1 => n6877, A2 => n4207, Z => n27153);
   U9015 : INV_X1 port map( I => n24839, ZN => n3233);
   U21655 : INV_X1 port map( I => n24522, ZN => n24658);
   U6784 : INV_X1 port map( I => n16319, ZN => n7466);
   U3744 : INV_X1 port map( I => n13695, ZN => n24642);
   U3027 : BUF_X2 port map( I => n25308, Z => n25962);
   U17370 : NOR2_X1 port map( A1 => n7413, A2 => n24607, ZN => n6326);
   U2117 : NOR2_X1 port map( A1 => n13532, A2 => n16397, ZN => n6691);
   U8419 : NAND2_X1 port map( A1 => n15719, A2 => n24874, ZN => n27926);
   U2261 : INV_X2 port map( I => n12676, ZN => n24725);
   U19329 : INV_X1 port map( I => n4885, ZN => n18264);
   U4424 : INV_X1 port map( I => n25012, ZN => n17684);
   U16251 : AOI21_X1 port map( A1 => n13050, A2 => n25872, B => n884, ZN => 
                           n4931);
   U4393 : NAND2_X1 port map( A1 => n16729, A2 => n16276, ZN => n16728);
   U26368 : NAND2_X1 port map( A1 => n4885, A2 => n32760, ZN => n11953);
   U25363 : NOR2_X1 port map( A1 => n4318, A2 => n25871, ZN => n23960);
   U4731 : NOR2_X1 port map( A1 => n13985, A2 => n18059, ZN => n5793);
   U2316 : NOR2_X1 port map( A1 => n717, A2 => n25756, ZN => n3275);
   U12928 : OAI21_X1 port map( A1 => n12086, A2 => n12926, B => n718, ZN => 
                           n3885);
   U15073 : INV_X1 port map( I => n1221, ZN => n27128);
   U7762 : NAND2_X1 port map( A1 => n2967, A2 => n26270, ZN => n24413);
   U19613 : NOR2_X1 port map( A1 => n27862, A2 => n27861, ZN => n28875);
   U52 : INV_X1 port map( I => n25712, ZN => n12314);
   U10317 : NAND2_X1 port map( A1 => n2536, A2 => n30288, ZN => n10359);
   U5554 : INV_X1 port map( I => n25664, ZN => n25659);
   U2146 : INV_X1 port map( I => n24970, ZN => n29049);
   U9260 : INV_X2 port map( I => n25689, ZN => n26447);
   U25541 : INV_X1 port map( I => n24956, ZN => n24938);
   U25495 : INV_X1 port map( I => n25490, ZN => n25475);
   U6035 : INV_X1 port map( I => n12611, ZN => n12309);
   U23695 : OAI21_X1 port map( A1 => n8676, A2 => n16670, B => n12611, ZN => 
                           n25793);
   U1 : OR2_X1 port map( A1 => n14208, A2 => n964, Z => n9902);
   U9 : NAND2_X1 port map( A1 => n25474, A2 => n25475, ZN => n30118);
   U11 : NAND3_X1 port map( A1 => n31647, A2 => n8320, A3 => n13483, ZN => 
                           n30134);
   U12 : NAND3_X1 port map( A1 => n14944, A2 => n15134, A3 => n31236, ZN => 
                           n8804);
   U13 : OR2_X1 port map( A1 => n27164, A2 => n1597, Z => n7040);
   U15 : OR2_X1 port map( A1 => n8515, A2 => n9956, Z => n30330);
   U34 : NOR2_X1 port map( A1 => n28070, A2 => n25060, ZN => n17728);
   U43 : INV_X1 port map( I => n25214, ZN => n25220);
   U58 : INV_X1 port map( I => n25665, ZN => n25658);
   U90 : OAI21_X1 port map( A1 => n31602, A2 => n31603, B => n33278, ZN => 
                           n29911);
   U124 : NOR2_X1 port map( A1 => n32571, A2 => n1212, ZN => n30876);
   U127 : NOR2_X1 port map( A1 => n17781, A2 => n11945, ZN => n31603);
   U131 : INV_X1 port map( I => n24471, ZN => n30461);
   U133 : NAND2_X1 port map( A1 => n14959, A2 => n25012, ZN => n30145);
   U135 : NOR2_X1 port map( A1 => n884, A2 => n13042, ZN => n31463);
   U137 : OR2_X1 port map( A1 => n25892, A2 => n25890, Z => n14042);
   U139 : NOR2_X1 port map( A1 => n883, A2 => n25885, ZN => n4930);
   U158 : NOR2_X1 port map( A1 => n24725, A2 => n13050, ZN => n31464);
   U163 : OAI21_X1 port map( A1 => n30998, A2 => n6691, B => n837, ZN => n30386
                           );
   U164 : INV_X2 port map( I => n547, ZN => n14268);
   U170 : OR2_X1 port map( A1 => n5897, A2 => n14454, Z => n29351);
   U171 : NOR2_X1 port map( A1 => n14055, A2 => n15318, ZN => n14484);
   U213 : NAND2_X1 port map( A1 => n25900, A2 => n25897, ZN => n24461);
   U231 : INV_X1 port map( I => n25700, ZN => n3565);
   U240 : CLKBUF_X2 port map( I => n25023, Z => n8210);
   U268 : INV_X1 port map( I => n24531, ZN => n29589);
   U295 : NAND3_X1 port map( A1 => n24124, A2 => n24182, A3 => n11463, ZN => 
                           n13204);
   U303 : NAND2_X1 port map( A1 => n12312, A2 => n6001, ZN => n29502);
   U316 : NAND2_X1 port map( A1 => n24162, A2 => n14592, ZN => n16859);
   U319 : CLKBUF_X1 port map( I => n4151, Z => n27500);
   U329 : NAND3_X1 port map( A1 => n17588, A2 => n1232, A3 => n17589, ZN => 
                           n17587);
   U335 : NOR2_X1 port map( A1 => n24039, A2 => n6001, ZN => n31016);
   U356 : OR2_X1 port map( A1 => n2444, A2 => n13175, Z => n10859);
   U357 : NAND2_X1 port map( A1 => n26314, A2 => n839, ZN => n5366);
   U369 : CLKBUF_X2 port map( I => n15536, Z => n29306);
   U373 : AND2_X1 port map( A1 => n1244, A2 => n24289, Z => n29293);
   U383 : NAND2_X1 port map( A1 => n14252, A2 => n319, ZN => n29512);
   U395 : INV_X1 port map( I => n24314, ZN => n10033);
   U406 : NAND2_X1 port map( A1 => n28350, A2 => n9214, ZN => n30280);
   U407 : CLKBUF_X2 port map( I => n14619, Z => n31883);
   U408 : CLKBUF_X1 port map( I => n14335, Z => n31271);
   U411 : NAND2_X1 port map( A1 => n28210, A2 => n23880, ZN => n23709);
   U424 : NAND2_X1 port map( A1 => n7993, A2 => n30251, ZN => n664);
   U426 : OAI21_X1 port map( A1 => n11131, A2 => n15446, B => n23932, ZN => 
                           n30898);
   U455 : OAI21_X1 port map( A1 => n27678, A2 => n23867, B => n10142, ZN => 
                           n17807);
   U461 : OAI21_X1 port map( A1 => n14513, A2 => n29590, B => n5417, ZN => 
                           n14990);
   U490 : AND2_X1 port map( A1 => n23904, A2 => n23905, Z => n17287);
   U496 : NAND3_X1 port map( A1 => n26074, A2 => n23721, A3 => n15095, ZN => 
                           n28194);
   U497 : NAND2_X1 port map( A1 => n31696, A2 => n739, ZN => n25954);
   U503 : INV_X1 port map( I => n23590, ZN => n14746);
   U514 : NOR2_X1 port map( A1 => n14975, A2 => n12680, ZN => n30620);
   U521 : INV_X1 port map( I => n17694, ZN => n31175);
   U523 : OAI21_X1 port map( A1 => n16786, A2 => n14297, B => n23852, ZN => 
                           n29682);
   U543 : OR2_X1 port map( A1 => n23720, A2 => n23719, Z => n23510);
   U568 : NOR2_X1 port map( A1 => n23887, A2 => n23840, ZN => n23632);
   U570 : NOR2_X1 port map( A1 => n29240, A2 => n23713, ZN => n31158);
   U588 : INV_X1 port map( I => n23720, ZN => n23917);
   U605 : AOI22_X1 port map( A1 => n3173, A2 => n23100, B1 => n3174, B2 => n986
                           , ZN => n3172);
   U622 : AND2_X1 port map( A1 => n30231, A2 => n16280, Z => n16975);
   U629 : NAND2_X1 port map( A1 => n5874, A2 => n23111, ZN => n30123);
   U638 : AND2_X1 port map( A1 => n22832, A2 => n31943, Z => n17064);
   U646 : NOR2_X1 port map( A1 => n17828, A2 => n31549, ZN => n31548);
   U647 : NOR3_X1 port map( A1 => n28957, A2 => n28801, A3 => n22748, ZN => 
                           n30247);
   U651 : NAND2_X1 port map( A1 => n23083, A2 => n7802, ZN => n23084);
   U664 : NAND2_X1 port map( A1 => n16254, A2 => n30476, ZN => n27834);
   U675 : OAI21_X1 port map( A1 => n15039, A2 => n32119, B => n33675, ZN => 
                           n5619);
   U700 : OAI22_X1 port map( A1 => n22761, A2 => n641, B1 => n15704, B2 => 
                           n15301, ZN => n10404);
   U719 : CLKBUF_X2 port map( I => n26898, Z => n30976);
   U733 : NOR2_X1 port map( A1 => n3163, A2 => n29317, ZN => n23074);
   U786 : NAND2_X2 port map( A1 => n30762, A2 => n30349, ZN => n31637);
   U790 : OR2_X1 port map( A1 => n22587, A2 => n1125, Z => n29406);
   U791 : OR2_X1 port map( A1 => n13710, A2 => n15089, Z => n12019);
   U808 : NAND3_X1 port map( A1 => n31559, A2 => n22646, A3 => n4459, ZN => 
                           n9156);
   U844 : NAND3_X1 port map( A1 => n858, A2 => n22670, A3 => n29495, ZN => 
                           n1516);
   U860 : NAND2_X1 port map( A1 => n22681, A2 => n10354, ZN => n17569);
   U873 : NAND2_X1 port map( A1 => n22647, A2 => n5961, ZN => n31559);
   U887 : NOR2_X1 port map( A1 => n18062, A2 => n22651, ZN => n29583);
   U892 : NOR2_X1 port map( A1 => n17960, A2 => n22524, ZN => n26144);
   U911 : OR2_X1 port map( A1 => n11895, A2 => n32532, Z => n22200);
   U916 : NOR3_X1 port map( A1 => n5769, A2 => n355, A3 => n31931, ZN => n28661
                           );
   U917 : AOI21_X1 port map( A1 => n1000, A2 => n22681, B => n10282, ZN => 
                           n17269);
   U925 : OAI21_X1 port map( A1 => n6257, A2 => n28424, B => n29342, ZN => 
                           n31363);
   U928 : OR2_X1 port map( A1 => n16277, A2 => n13704, Z => n22648);
   U932 : AND2_X1 port map( A1 => n22670, A2 => n1127, Z => n29371);
   U933 : AND2_X1 port map( A1 => n22636, A2 => n12043, Z => n29355);
   U937 : NAND2_X1 port map( A1 => n10725, A2 => n22645, ZN => n29562);
   U939 : NAND2_X1 port map( A1 => n31838, A2 => n11083, ZN => n118);
   U941 : AND2_X1 port map( A1 => n15089, A2 => n32172, Z => n12556);
   U949 : INV_X1 port map( I => n22670, ZN => n30106);
   U957 : NOR2_X1 port map( A1 => n17960, A2 => n1728, ZN => n15033);
   U989 : NAND2_X1 port map( A1 => n10622, A2 => n10568, ZN => n9752);
   U1020 : BUF_X2 port map( I => n11907, Z => n29304);
   U1037 : INV_X1 port map( I => n22232, ZN => n2863);
   U1041 : INV_X1 port map( I => n3704, ZN => n30087);
   U1045 : INV_X1 port map( I => n3634, ZN => n26863);
   U1047 : INV_X1 port map( I => n22227, ZN => n30747);
   U1068 : OAI21_X1 port map( A1 => n10215, A2 => n11081, B => n21673, ZN => 
                           n17681);
   U1071 : AND2_X1 port map( A1 => n21465, A2 => n1134, Z => n29455);
   U1073 : AOI21_X1 port map( A1 => n31511, A2 => n21786, B => n1323, ZN => 
                           n4687);
   U1078 : NAND2_X1 port map( A1 => n15091, A2 => n21581, ZN => n31089);
   U1084 : AND2_X1 port map( A1 => n2575, A2 => n16023, Z => n29435);
   U1095 : AND2_X1 port map( A1 => n32252, A2 => n27635, Z => n29407);
   U1096 : AND2_X1 port map( A1 => n17098, A2 => n21463, Z => n10215);
   U1098 : NOR2_X1 port map( A1 => n17472, A2 => n29302, ZN => n10028);
   U1114 : NAND3_X1 port map( A1 => n861, A2 => n21687, A3 => n21688, ZN => 
                           n31121);
   U1116 : AND2_X1 port map( A1 => n30506, A2 => n28429, Z => n12279);
   U1118 : NOR2_X1 port map( A1 => n21717, A2 => n26710, ZN => n7986);
   U1130 : NOR2_X1 port map( A1 => n21645, A2 => n21646, ZN => n21091);
   U1134 : NAND2_X1 port map( A1 => n11861, A2 => n21583, ZN => n3588);
   U1137 : OR2_X1 port map( A1 => n21687, A2 => n21688, Z => n12102);
   U1138 : NOR2_X1 port map( A1 => n28729, A2 => n12394, ZN => n29796);
   U1144 : AOI22_X1 port map( A1 => n1008, A2 => n8313, B1 => n21799, B2 => 
                           n21797, ZN => n31026);
   U1174 : NAND2_X1 port map( A1 => n30326, A2 => n21553, ZN => n21678);
   U1175 : NAND2_X1 port map( A1 => n21716, A2 => n21715, ZN => n7276);
   U1186 : OR2_X1 port map( A1 => n5170, A2 => n9999, Z => n2337);
   U1200 : OR2_X1 port map( A1 => n29258, A2 => n1652, Z => n11796);
   U1208 : NOR3_X1 port map( A1 => n27560, A2 => n29854, A3 => n21730, ZN => 
                           n29943);
   U1224 : INV_X1 port map( I => n9666, ZN => n11729);
   U1226 : NAND2_X1 port map( A1 => n21755, A2 => n26451, ZN => n30902);
   U1229 : OR2_X1 port map( A1 => n26445, A2 => n27336, Z => n16864);
   U1232 : NOR2_X1 port map( A1 => n31511, A2 => n21786, ZN => n11938);
   U1278 : NOR2_X1 port map( A1 => n27563, A2 => n29777, ZN => n21509);
   U1289 : NAND2_X1 port map( A1 => n12340, A2 => n21183, ZN => n30700);
   U1290 : NOR2_X1 port map( A1 => n10921, A2 => n21127, ZN => n31677);
   U1306 : OAI21_X1 port map( A1 => n21396, A2 => n27955, B => n3933, ZN => 
                           n31815);
   U1308 : NOR2_X1 port map( A1 => n21306, A2 => n21303, ZN => n30544);
   U1334 : NAND2_X1 port map( A1 => n3933, A2 => n29303, ZN => n21286);
   U1337 : INV_X1 port map( I => n21506, ZN => n29777);
   U1340 : INV_X1 port map( I => n4683, ZN => n728);
   U1341 : NAND2_X1 port map( A1 => n16639, A2 => n320, ZN => n7526);
   U1393 : NOR2_X1 port map( A1 => n28037, A2 => n21253, ZN => n15932);
   U1399 : OR2_X1 port map( A1 => n31614, A2 => n349, Z => n31613);
   U1400 : NOR2_X1 port map( A1 => n11734, A2 => n1148, ZN => n30863);
   U1406 : AOI21_X1 port map( A1 => n11187, A2 => n21189, B => n2822, ZN => 
                           n14023);
   U1407 : OR2_X1 port map( A1 => n21442, A2 => n21100, Z => n21304);
   U1414 : OAI21_X1 port map( A1 => n21307, A2 => n21443, B => n21306, ZN => 
                           n21308);
   U1428 : INV_X1 port map( I => n21270, ZN => n31476);
   U1485 : CLKBUF_X2 port map( I => n21356, Z => n28701);
   U1486 : BUF_X2 port map( I => n21165, Z => n27075);
   U1498 : OR2_X1 port map( A1 => n9405, A2 => n9626, Z => n31004);
   U1499 : BUF_X2 port map( I => n21432, Z => n320);
   U1515 : INV_X1 port map( I => n13092, ZN => n30543);
   U1533 : NAND3_X1 port map( A1 => n10765, A2 => n8797, A3 => n10764, ZN => 
                           n31608);
   U1534 : INV_X1 port map( I => n6500, ZN => n30430);
   U1535 : OR2_X1 port map( A1 => n14177, A2 => n32329, Z => n7956);
   U1560 : NAND3_X1 port map( A1 => n16004, A2 => n9688, A3 => n8087, ZN => 
                           n30197);
   U1561 : NAND2_X1 port map( A1 => n3644, A2 => n31047, ZN => n5413);
   U1563 : NAND2_X1 port map( A1 => n16132, A2 => n20523, ZN => n30414);
   U1600 : INV_X1 port map( I => n31211, ZN => n31210);
   U1626 : OR2_X1 port map( A1 => n20471, A2 => n29337, Z => n2766);
   U1635 : NAND2_X1 port map( A1 => n30425, A2 => n32504, ZN => n2767);
   U1642 : INV_X1 port map( I => n20537, ZN => n31250);
   U1645 : OAI22_X1 port map( A1 => n20528, A2 => n13499, B1 => n13599, B2 => 
                           n11984, ZN => n31022);
   U1646 : NOR2_X1 port map( A1 => n8206, A2 => n27771, ZN => n30471);
   U1650 : NOR2_X1 port map( A1 => n28626, A2 => n741, ZN => n29724);
   U1654 : OAI21_X1 port map( A1 => n2879, A2 => n14187, B => n33530, ZN => 
                           n7867);
   U1684 : NAND2_X1 port map( A1 => n7242, A2 => n6530, ZN => n15833);
   U1687 : CLKBUF_X2 port map( I => n2928, Z => n31804);
   U1691 : NAND2_X1 port map( A1 => n8770, A2 => n14436, ZN => n3787);
   U1693 : NAND3_X1 port map( A1 => n31721, A2 => n13759, A3 => n20310, ZN => 
                           n29983);
   U1708 : BUF_X2 port map( I => n20384, Z => n30594);
   U1711 : INV_X1 port map( I => n20345, ZN => n30138);
   U1715 : NOR2_X1 port map( A1 => n20463, A2 => n20371, ZN => n20464);
   U1729 : BUF_X2 port map( I => n20581, Z => n6230);
   U1731 : INV_X1 port map( I => n19909, ZN => n29668);
   U1744 : NAND2_X1 port map( A1 => n15286, A2 => n31766, ZN => n15285);
   U1759 : OAI21_X1 port map( A1 => n8421, A2 => n19971, B => n31164, ZN => 
                           n8759);
   U1767 : NOR3_X1 port map( A1 => n20010, A2 => n20008, A3 => n9876, ZN => 
                           n9341);
   U1772 : NAND3_X1 port map( A1 => n20028, A2 => n20025, A3 => n1042, ZN => 
                           n19735);
   U1774 : AOI22_X1 port map( A1 => n1361, A2 => n11893, B1 => n3591, B2 => 
                           n19794, ZN => n3590);
   U1777 : NOR2_X1 port map( A1 => n34153, A2 => n20100, ZN => n19562);
   U1780 : NOR2_X1 port map( A1 => n30064, A2 => n16966, ZN => n16979);
   U1792 : NOR2_X1 port map( A1 => n20136, A2 => n20037, ZN => n31766);
   U1795 : NAND2_X1 port map( A1 => n10072, A2 => n19979, ZN => n31443);
   U1808 : NAND3_X1 port map( A1 => n18089, A2 => n7804, A3 => n31445, ZN => 
                           n8015);
   U1812 : INV_X1 port map( I => n875, ZN => n29840);
   U1817 : INV_X2 port map( I => n19867, ZN => n17608);
   U1818 : AND2_X1 port map( A1 => n29153, A2 => n4224, Z => n29358);
   U1829 : INV_X1 port map( I => n10413, ZN => n8147);
   U1845 : AND2_X1 port map( A1 => n20113, A2 => n19907, Z => n29373);
   U1855 : NOR2_X1 port map( A1 => n27808, A2 => n16812, ZN => n31697);
   U1860 : INV_X1 port map( I => n13650, ZN => n30017);
   U1869 : NOR2_X1 port map( A1 => n19901, A2 => n19900, ZN => n5999);
   U1875 : CLKBUF_X2 port map( I => n12040, Z => n6532);
   U1878 : INV_X1 port map( I => n1368, ZN => n30819);
   U1879 : INV_X1 port map( I => n19764, ZN => n31646);
   U1886 : INV_X1 port map( I => n27138, ZN => n29689);
   U1895 : NAND2_X1 port map( A1 => n5709, A2 => n5710, ZN => n31573);
   U1926 : NAND2_X1 port map( A1 => n16874, A2 => n30789, ZN => n16873);
   U1930 : INV_X1 port map( I => n29781, ZN => n31217);
   U1932 : NAND2_X1 port map( A1 => n18977, A2 => n8092, ZN => n30660);
   U1933 : AOI21_X1 port map( A1 => n27743, A2 => n28705, B => n16669, ZN => 
                           n12498);
   U1945 : AND2_X1 port map( A1 => n30663, A2 => n339, Z => n10013);
   U1962 : CLKBUF_X2 port map( I => n19332, Z => n28404);
   U1968 : NAND2_X1 port map( A1 => n29815, A2 => n7687, ZN => n30789);
   U1972 : NOR2_X1 port map( A1 => n1384, A2 => n31352, ZN => n31351);
   U1975 : NAND2_X1 port map( A1 => n16960, A2 => n8335, ZN => n19333);
   U1978 : BUF_X2 port map( I => n8606, Z => n26830);
   U1999 : NAND3_X1 port map( A1 => n29684, A2 => n3364, A3 => n29683, ZN => 
                           n3361);
   U2001 : NAND3_X1 port map( A1 => n26398, A2 => n18581, A3 => n18724, ZN => 
                           n26591);
   U2005 : NOR2_X1 port map( A1 => n18578, A2 => n30866, ZN => n11319);
   U2008 : AOI22_X1 port map( A1 => n485, A2 => n18571, B1 => n5753, B2 => 
                           n4868, ZN => n5751);
   U2011 : NAND3_X1 port map( A1 => n26717, A2 => n3601, A3 => n10579, ZN => 
                           n2684);
   U2018 : NAND2_X1 port map( A1 => n15956, A2 => n31519, ZN => n18491);
   U2020 : NOR2_X1 port map( A1 => n469, A2 => n25981, ZN => n8271);
   U2030 : NOR2_X1 port map( A1 => n1188, A2 => n8739, ZN => n7977);
   U2031 : OAI22_X1 port map( A1 => n16247, A2 => n16352, B1 => n18822, B2 => 
                           n18820, ZN => n30001);
   U2035 : NAND3_X1 port map( A1 => n18635, A2 => n5269, A3 => n6037, ZN => 
                           n18636);
   U2038 : NAND2_X1 port map( A1 => n17582, A2 => n16948, ZN => n31339);
   U2044 : OR2_X1 port map( A1 => n18574, A2 => n18617, Z => n8821);
   U2045 : NOR2_X1 port map( A1 => n6256, A2 => n13738, ZN => n31519);
   U2048 : AND2_X1 port map( A1 => n18586, A2 => n28964, Z => n17165);
   U2051 : NOR2_X1 port map( A1 => n18822, A2 => n16249, ZN => n30698);
   U2058 : NOR2_X1 port map( A1 => n18867, A2 => n31986, ZN => n30908);
   U2059 : OAI21_X1 port map( A1 => n3601, A2 => n26040, B => n27228, ZN => 
                           n11323);
   U2060 : NAND3_X1 port map( A1 => n1188, A2 => n8739, A3 => n18639, ZN => 
                           n18640);
   U2061 : NOR2_X1 port map( A1 => n16569, A2 => n12006, ZN => n18469);
   U2064 : CLKBUF_X1 port map( I => n15966, Z => n26155);
   U2091 : BUF_X1 port map( I => n18186, Z => n30744);
   U2097 : AOI21_X2 port map( A1 => n18324, A2 => n34139, B => n180, ZN => 
                           n12214);
   U2099 : BUF_X4 port map( I => n24257, Z => n6476);
   U2106 : OAI22_X2 port map( A1 => n10731, A2 => n17228, B1 => n15832, B2 => 
                           n20516, ZN => n30304);
   U2107 : OAI21_X2 port map( A1 => n13300, A2 => n33301, B => n13830, ZN => 
                           n20311);
   U2113 : NOR2_X2 port map( A1 => n18487, A2 => n18827, ZN => n18462);
   U2114 : BUF_X2 port map( I => n15955, Z => n14828);
   U2121 : NAND2_X2 port map( A1 => n29398, A2 => n19225, ZN => n13938);
   U2124 : BUF_X2 port map( I => n17237, Z => n8454);
   U2125 : BUF_X4 port map( I => n2396, Z => n2141);
   U2127 : AOI21_X2 port map( A1 => n1373, A2 => n11940, B => n1764, ZN => 
                           n1763);
   U2129 : AND2_X1 port map( A1 => n18768, A2 => n16849, Z => n18376);
   U2142 : BUF_X4 port map( I => n18722, Z => n29602);
   U2154 : OR2_X1 port map( A1 => n10568, A2 => n28014, Z => n22466);
   U2161 : OAI21_X2 port map( A1 => n12590, A2 => n20079, B => n6444, ZN => 
                           n26961);
   U2170 : INV_X2 port map( I => n14789, ZN => n27545);
   U2171 : NAND2_X1 port map( A1 => n30976, A2 => n5374, ZN => n29621);
   U2177 : INV_X2 port map( I => n26445, ZN => n28435);
   U2198 : AOI21_X2 port map( A1 => n1287, A2 => n30405, B => n29232, ZN => 
                           n27565);
   U2200 : NAND3_X2 port map( A1 => n12053, A2 => n14283, A3 => n1039, ZN => 
                           n31319);
   U2210 : AND2_X1 port map( A1 => n21306, A2 => n21305, Z => n29382);
   U2218 : NAND2_X2 port map( A1 => n15830, A2 => n22992, ZN => n30388);
   U2230 : INV_X2 port map( I => n23156, ZN => n18133);
   U2231 : AOI21_X2 port map( A1 => n1170, A2 => n19456, B => n16681, ZN => 
                           n6858);
   U2232 : BUF_X2 port map( I => n18696, Z => n16569);
   U2234 : INV_X4 port map( I => n7287, ZN => n23055);
   U2245 : OR2_X1 port map( A1 => n18696, A2 => n18831, Z => n13015);
   U2246 : OR2_X1 port map( A1 => n23540, A2 => n24283, Z => n28781);
   U2254 : INV_X2 port map( I => n28091, ZN => n30737);
   U2266 : INV_X2 port map( I => n25201, ZN => n25200);
   U2268 : INV_X4 port map( I => n16651, ZN => n29056);
   U2270 : INV_X2 port map( I => n29153, ZN => n6962);
   U2274 : OAI22_X1 port map( A1 => n16254, A2 => n6360, B1 => n6012, B2 => 
                           n16022, ZN => n5874);
   U2275 : OAI21_X1 port map( A1 => n23708, A2 => n16238, B => n14974, ZN => 
                           n12509);
   U2283 : NAND2_X1 port map( A1 => n12837, A2 => n17223, ZN => n18029);
   U2284 : NAND2_X1 port map( A1 => n17582, A2 => n17223, ZN => n16338);
   U2285 : INV_X1 port map( I => n17223, ZN => n29751);
   U2286 : CLKBUF_X2 port map( I => n10469, Z => n7371);
   U2291 : NAND3_X1 port map( A1 => n1290, A2 => n6478, A3 => n8409, ZN => 
                           n22555);
   U2293 : INV_X1 port map( I => n25903, ZN => n29771);
   U2295 : NAND2_X1 port map( A1 => n31801, A2 => n7093, ZN => n29584);
   U2303 : NAND2_X1 port map( A1 => n5417, A2 => n15038, ZN => n30515);
   U2321 : OAI21_X1 port map( A1 => n29261, A2 => n900, B => n22476, ZN => 
                           n30383);
   U2331 : AOI21_X1 port map( A1 => n15757, A2 => n11556, B => n15755, ZN => 
                           n15769);
   U2336 : NOR2_X1 port map( A1 => n17120, A2 => n30221, ZN => n31245);
   U2338 : AND2_X1 port map( A1 => n33007, A2 => n22795, Z => n29438);
   U2345 : INV_X1 port map( I => n10111, ZN => n24781);
   U2352 : NAND2_X1 port map( A1 => n29107, A2 => n23058, ZN => n14418);
   U2357 : INV_X2 port map( I => n25736, ZN => n25744);
   U2358 : NAND2_X1 port map( A1 => n14721, A2 => n21223, ZN => n21316);
   U2360 : NOR3_X1 port map( A1 => n26868, A2 => n14188, A3 => n28697, ZN => 
                           n16140);
   U2395 : NOR2_X1 port map( A1 => n18764, A2 => n18767, ZN => n31521);
   U2397 : NAND2_X1 port map( A1 => n30369, A2 => n25211, ZN => n10942);
   U2406 : NAND2_X1 port map( A1 => n6483, A2 => n21721, ZN => n14076);
   U2416 : CLKBUF_X2 port map( I => n24914, Z => n27248);
   U2417 : OAI22_X1 port map( A1 => n12615, A2 => n23144, B1 => n17257, B2 => 
                           n6479, ZN => n26392);
   U2431 : INV_X1 port map( I => n12329, ZN => n25076);
   U2439 : INV_X1 port map( I => n661, ZN => n4892);
   U2444 : CLKBUF_X4 port map( I => n16141, Z => n12);
   U2454 : NOR2_X1 port map( A1 => n13985, A2 => n25198, ZN => n1861);
   U2463 : AOI21_X1 port map( A1 => n16117, A2 => n5056, B => n13073, ZN => 
                           n18221);
   U2480 : OAI21_X1 port map( A1 => n7655, A2 => n1215, B => n27342, ZN => 
                           n1859);
   U2495 : NAND2_X1 port map( A1 => n13268, A2 => n24210, ZN => n24321);
   U2521 : OAI21_X1 port map( A1 => n28473, A2 => n28472, B => n22435, ZN => 
                           n11441);
   U2537 : OAI21_X1 port map( A1 => n15359, A2 => n25214, B => n15339, ZN => 
                           n30369);
   U2544 : AND2_X1 port map( A1 => n29304, A2 => n8275, Z => n4812);
   U2545 : NAND3_X1 port map( A1 => n27123, A2 => n29085, A3 => n1071, ZN => 
                           n4768);
   U2548 : OAI21_X1 port map( A1 => n16097, A2 => n23848, B => n23847, ZN => 
                           n10762);
   U2554 : BUF_X2 port map( I => n23567, Z => n23848);
   U2574 : INV_X1 port map( I => n9664, ZN => n10483);
   U2584 : BUF_X2 port map( I => n4599, Z => n3898);
   U2593 : NOR2_X1 port map( A1 => n15054, A2 => n2191, ZN => n7928);
   U2599 : BUF_X2 port map( I => n24147, Z => n4019);
   U2623 : NAND2_X1 port map( A1 => n2746, A2 => n2745, ZN => n30110);
   U2626 : BUF_X2 port map( I => n5128, Z => n4781);
   U2628 : NAND2_X1 port map( A1 => n25132, A2 => n1083, ZN => n31780);
   U2630 : INV_X1 port map( I => n1083, ZN => n31779);
   U2644 : INV_X2 port map( I => n25867, ZN => n790);
   U2646 : NOR3_X1 port map( A1 => n29706, A2 => n13049, A3 => n25847, ZN => 
                           n15944);
   U2666 : OAI21_X1 port map( A1 => n24715, A2 => n16323, B => n9195, ZN => 
                           n24716);
   U2670 : NOR2_X1 port map( A1 => n16323, A2 => n25701, ZN => n24449);
   U2679 : OR2_X1 port map( A1 => n9163, A2 => n9164, Z => n27376);
   U2687 : NOR2_X1 port map( A1 => n11575, A2 => n6882, ZN => n642);
   U2702 : AND2_X1 port map( A1 => n17927, A2 => n10858, Z => n9655);
   U2758 : NOR2_X1 port map( A1 => n19857, A2 => n17711, ZN => n11903);
   U2768 : NAND2_X1 port map( A1 => n31920, A2 => n4490, ZN => n24711);
   U2770 : OAI21_X1 port map( A1 => n16467, A2 => n9391, B => n7073, ZN => 
                           n7505);
   U2771 : NAND2_X1 port map( A1 => n27479, A2 => n13709, ZN => n12293);
   U2780 : NAND2_X1 port map( A1 => n22422, A2 => n906, ZN => n30639);
   U2790 : NOR2_X1 port map( A1 => n11299, A2 => n12363, ZN => n12372);
   U2810 : AND2_X1 port map( A1 => n9199, A2 => n651, Z => n13666);
   U2817 : NOR2_X1 port map( A1 => n6910, A2 => n25394, ZN => n25347);
   U2822 : NOR2_X1 port map( A1 => n30139, A2 => n1863, ZN => n31286);
   U2823 : NAND2_X1 port map( A1 => n6668, A2 => n2042, ZN => n6667);
   U2826 : INV_X1 port map( I => n19509, ZN => n8456);
   U2838 : AND2_X1 port map( A1 => n14335, A2 => n3860, Z => n1978);
   U2841 : AND2_X1 port map( A1 => n14335, A2 => n31294, Z => n31293);
   U2842 : AND2_X1 port map( A1 => n6595, A2 => n8766, Z => n8710);
   U2845 : INV_X1 port map( I => n11334, ZN => n6133);
   U2849 : NOR2_X1 port map( A1 => n11334, A2 => n22584, ZN => n17007);
   U2879 : NAND2_X1 port map( A1 => n15550, A2 => n13050, ZN => n12677);
   U2894 : BUF_X2 port map( I => n25221, Z => n28651);
   U2915 : CLKBUF_X2 port map( I => n29157, Z => n31722);
   U2916 : NAND3_X1 port map( A1 => n30328, A2 => n24927, A3 => n2180, ZN => 
                           n24350);
   U2921 : CLKBUF_X1 port map( I => n11931, Z => n27057);
   U2922 : NOR2_X1 port map( A1 => n11931, A2 => n10504, ZN => n25617);
   U2923 : CLKBUF_X2 port map( I => n14865, Z => n254);
   U2925 : INV_X1 port map( I => n14865, ZN => n25003);
   U2950 : NAND2_X1 port map( A1 => n29253, A2 => n8100, ZN => n13962);
   U2953 : NAND2_X1 port map( A1 => n12677, A2 => n25884, ZN => n24463);
   U2954 : NAND2_X1 port map( A1 => n25884, A2 => n14832, ZN => n4932);
   U2965 : AND2_X1 port map( A1 => n25973, A2 => n24251, Z => n29376);
   U2971 : NOR2_X1 port map( A1 => n25060, A2 => n25051, ZN => n25063);
   U2976 : NAND3_X1 port map( A1 => n12974, A2 => n842, A3 => n14756, ZN => 
                           n16947);
   U2979 : NOR2_X1 port map( A1 => n25980, A2 => n14210, ZN => n12784);
   U2981 : AND2_X1 port map( A1 => n7748, A2 => n1984, Z => n1983);
   U2985 : AND3_X1 port map( A1 => n5760, A2 => n18990, A3 => n18017, Z => 
                           n10867);
   U2989 : BUF_X2 port map( I => n18017, Z => n28171);
   U3002 : AOI21_X1 port map( A1 => n21811, A2 => n28181, B => n1328, ZN => 
                           n21349);
   U3017 : AOI22_X1 port map( A1 => n891, A2 => n3506, B1 => n29576, B2 => 
                           n28410, ZN => n6106);
   U3019 : AOI22_X1 port map( A1 => n10567, A2 => n790, B1 => n18219, B2 => 
                           n790, ZN => n10566);
   U3026 : NOR2_X1 port map( A1 => n16041, A2 => n72, ZN => n16937);
   U3030 : INV_X2 port map( I => n16041, ZN => n25312);
   U3040 : NAND2_X1 port map( A1 => n31916, A2 => n29268, ZN => n23616);
   U3056 : INV_X1 port map( I => n13159, ZN => n16817);
   U3077 : OAI21_X1 port map( A1 => n16149, A2 => n22576, B => n16567, ZN => 
                           n6657);
   U3112 : NOR3_X1 port map( A1 => n1119, A2 => n1926, A3 => n1805, ZN => n1887
                           );
   U3125 : OAI21_X1 port map( A1 => n1165, A2 => n13061, B => n31684, ZN => 
                           n14988);
   U3131 : NAND3_X1 port map( A1 => n15736, A2 => n31684, A3 => n1165, ZN => 
                           n15735);
   U3132 : NOR2_X1 port map( A1 => n1165, A2 => n29152, ZN => n15306);
   U3152 : OAI21_X1 port map( A1 => n15189, A2 => n20155, B => n3486, ZN => 
                           n6069);
   U3156 : INV_X1 port map( I => n5988, ZN => n25575);
   U3157 : AOI22_X1 port map( A1 => n19117, A2 => n28404, B1 => n19154, B2 => 
                           n8862, ZN => n12368);
   U3162 : OAI21_X1 port map( A1 => n880, A2 => n879, B => n19154, ZN => n16221
                           );
   U3169 : NOR2_X1 port map( A1 => n11366, A2 => n16528, ZN => n30372);
   U3182 : NOR2_X1 port map( A1 => n17894, A2 => n25901, ZN => n4205);
   U3186 : AND2_X1 port map( A1 => n386, A2 => n30089, Z => n15404);
   U3191 : NOR2_X1 port map( A1 => n7195, A2 => n21441, ZN => n2689);
   U3196 : OAI21_X1 port map( A1 => n31195, A2 => n7195, B => n21441, ZN => 
                           n7196);
   U3198 : AOI21_X1 port map( A1 => n796, A2 => n10226, B => n7935, ZN => 
                           n11341);
   U3208 : NOR2_X1 port map( A1 => n21864, A2 => n21865, ZN => n8619);
   U3225 : NAND4_X1 port map( A1 => n3052, A2 => n3057, A3 => n3051, A4 => 
                           n18123, ZN => n3056);
   U3226 : NAND2_X1 port map( A1 => n15283, A2 => n30586, ZN => n12319);
   U3227 : INV_X1 port map( I => n19754, ZN => n26230);
   U3243 : OAI22_X1 port map( A1 => n24988, A2 => n713, B1 => n24994, B2 => 
                           n4525, ZN => n24989);
   U3248 : NAND2_X1 port map( A1 => n6500, A2 => n11617, ZN => n30551);
   U3250 : AOI21_X1 port map( A1 => n21587, A2 => n26766, B => n30806, ZN => 
                           n21589);
   U3267 : NOR3_X1 port map( A1 => n1211, A2 => n28338, A3 => n1212, ZN => 
                           n13296);
   U3271 : AOI21_X1 port map( A1 => n6763, A2 => n3340, B => n7134, ZN => n3343
                           );
   U3273 : INV_X2 port map( I => n6763, ZN => n31139);
   U3291 : BUF_X2 port map( I => n15255, Z => n26912);
   U3298 : INV_X1 port map( I => n15255, ZN => n25588);
   U3299 : NAND3_X1 port map( A1 => n15255, A2 => n11820, A3 => n34169, ZN => 
                           n25534);
   U3305 : OAI21_X1 port map( A1 => n4281, A2 => n28265, B => n30527, ZN => 
                           n7538);
   U3311 : BUF_X2 port map( I => n32309, Z => n4281);
   U3313 : NAND3_X1 port map( A1 => n15278, A2 => n10484, A3 => n19933, ZN => 
                           n1813);
   U3332 : NAND2_X1 port map( A1 => n26447, A2 => n27173, ZN => n28931);
   U3336 : NAND2_X1 port map( A1 => n791, A2 => n16688, ZN => n6250);
   U3337 : INV_X1 port map( I => n5932, ZN => n15264);
   U3344 : NOR2_X1 port map( A1 => n25637, A2 => n2378, ZN => n25638);
   U3346 : CLKBUF_X2 port map( I => n21455, Z => n29088);
   U3347 : CLKBUF_X2 port map( I => n3880, Z => n30969);
   U3348 : NAND2_X1 port map( A1 => n24084, A2 => n3880, ZN => n14677);
   U3354 : NAND2_X1 port map( A1 => n33722, A2 => n23813, ZN => n31294);
   U3363 : INV_X1 port map( I => n25816, ZN => n25826);
   U3374 : INV_X1 port map( I => n23924, ZN => n23736);
   U3386 : OAI21_X1 port map( A1 => n20437, A2 => n20438, B => n30099, ZN => 
                           n2650);
   U3391 : OAI22_X1 port map( A1 => n26520, A2 => n18827, B1 => n18489, B2 => 
                           n18487, ZN => n17251);
   U3392 : NAND2_X1 port map( A1 => n18487, A2 => n18827, ZN => n18332);
   U3393 : INV_X2 port map( I => n26791, ZN => n18487);
   U3394 : AOI21_X1 port map( A1 => n11888, A2 => n354, B => n8217, ZN => 
                           n13503);
   U3402 : NAND2_X1 port map( A1 => n32063, A2 => n24956, ZN => n24954);
   U3403 : NOR2_X1 port map( A1 => n1201, A2 => n32063, ZN => n8639);
   U3416 : INV_X1 port map( I => n23266, ZN => n23445);
   U3430 : INV_X1 port map( I => n14031, ZN => n1247);
   U3443 : AND2_X2 port map( A1 => n11913, A2 => n16, Z => n29281);
   U3445 : AND2_X1 port map( A1 => n29022, A2 => n20100, Z => n29283);
   U3447 : INV_X1 port map( I => n8713, ZN => n19921);
   U3449 : BUF_X2 port map( I => n8713, Z => n1826);
   U3461 : XNOR2_X1 port map( A1 => n10949, A2 => n6906, ZN => n29285);
   U3465 : NOR2_X2 port map( A1 => n7954, A2 => n7955, ZN => n6431);
   U3470 : INV_X1 port map( I => n20882, ZN => n21391);
   U3485 : INV_X2 port map( I => n14045, ZN => n853);
   U3497 : XNOR2_X1 port map( A1 => n23224, A2 => n16691, ZN => n29291);
   U3502 : INV_X2 port map( I => n6169, ZN => n14136);
   U3513 : INV_X2 port map( I => n4286, ZN => n15520);
   U3520 : INV_X2 port map( I => n23301, ZN => n30380);
   U3527 : INV_X4 port map( I => n25756, ZN => n1211);
   U3543 : BUF_X2 port map( I => n7242, Z => n28836);
   U3550 : AND2_X2 port map( A1 => n9490, A2 => n8277, Z => n15446);
   U3560 : INV_X1 port map( I => n4110, ZN => n22830);
   U3572 : NAND3_X1 port map( A1 => n16835, A2 => n700, A3 => n25867, ZN => 
                           n11254);
   U3573 : INV_X1 port map( I => n6255, ZN => n20481);
   U3584 : BUF_X2 port map( I => n29471, Z => n29294);
   U3585 : OAI21_X1 port map( A1 => n5272, A2 => n836, B => n25901, ZN => n5271
                           );
   U3617 : INV_X1 port map( I => n23808, ZN => n31483);
   U3627 : AOI21_X1 port map( A1 => n5670, A2 => n5779, B => n26585, ZN => 
                           n5669);
   U3629 : OR2_X2 port map( A1 => n28545, A2 => n26606, Z => n22646);
   U3632 : NAND2_X1 port map( A1 => n20527, A2 => n16515, ZN => n17392);
   U3648 : INV_X2 port map( I => n11372, ZN => n13273);
   U3650 : NAND2_X1 port map( A1 => n11372, A2 => n25977, ZN => n3791);
   U3651 : AND2_X2 port map( A1 => n9280, A2 => n9951, Z => n22843);
   U3654 : NAND3_X1 port map( A1 => n30902, A2 => n21512, A3 => n9057, ZN => 
                           n27437);
   U3657 : NOR2_X1 port map( A1 => n21755, A2 => n21512, ZN => n8276);
   U3674 : INV_X2 port map( I => n6669, ZN => n17077);
   U3676 : NAND2_X1 port map( A1 => n31911, A2 => n31309, ZN => n21801);
   U3687 : OAI22_X1 port map( A1 => n17255, A2 => n18617, B1 => n17062, B2 => 
                           n16948, ZN => n31333);
   U3696 : NAND2_X1 port map( A1 => n15108, A2 => n18617, ZN => n14536);
   U3701 : AND2_X1 port map( A1 => n1119, A2 => n13862, Z => n1594);
   U3733 : INV_X1 port map( I => n24621, ZN => n31088);
   U3741 : NOR2_X1 port map( A1 => n18546, A2 => n1185, ZN => n9510);
   U3743 : INV_X1 port map( I => n18546, ZN => n18647);
   U3746 : NOR2_X1 port map( A1 => n18546, A2 => n26810, ZN => n18363);
   U3753 : NOR2_X2 port map( A1 => n21321, A2 => n21322, ZN => n21190);
   U3761 : NOR2_X1 port map( A1 => n18110, A2 => n16129, ZN => n13582);
   U3778 : AOI21_X1 port map( A1 => n1041, A2 => n20097, B => n16789, ZN => 
                           n17442);
   U3794 : INV_X1 port map( I => n13720, ZN => n798);
   U3806 : BUF_X4 port map( I => n17278, Z => n29299);
   U3815 : NAND2_X1 port map( A1 => n12902, A2 => n20311, ZN => n31188);
   U3822 : AOI21_X2 port map( A1 => n17639, A2 => n14603, B => n14602, ZN => 
                           n14601);
   U3823 : NAND2_X2 port map( A1 => n12836, A2 => n9439, ZN => n27218);
   U3833 : NAND2_X1 port map( A1 => n11368, A2 => n20423, ZN => n26399);
   U3853 : INV_X1 port map( I => n19057, ZN => n1387);
   U3864 : INV_X2 port map( I => n14954, ZN => n10822);
   U3865 : NAND2_X1 port map( A1 => n12329, A2 => n14954, ZN => n25067);
   U3880 : NAND2_X1 port map( A1 => n10883, A2 => n27007, ZN => n39);
   U3883 : INV_X1 port map( I => n27007, ZN => n29635);
   U3885 : NAND2_X1 port map( A1 => n27007, A2 => n22824, ZN => n17605);
   U3886 : AND2_X2 port map( A1 => n27007, A2 => n22592, Z => n22823);
   U3899 : OAI21_X1 port map( A1 => n14168, A2 => n21072, B => n5141, ZN => 
                           n31025);
   U3914 : BUF_X2 port map( I => n10631, Z => n31508);
   U3933 : NOR2_X1 port map( A1 => n15864, A2 => n30506, ZN => n12280);
   U3948 : BUF_X2 port map( I => n16710, Z => n28378);
   U3962 : AND3_X1 port map( A1 => n21568, A2 => n21569, A3 => n30389, Z => 
                           n21570);
   U3976 : NOR4_X1 port map( A1 => n22729, A2 => n22730, A3 => n22731, A4 => 
                           n22732, ZN => n12055);
   U3980 : INV_X1 port map( I => n5454, ZN => n13048);
   U3983 : AOI21_X1 port map( A1 => n14620, A2 => n20261, B => n32747, ZN => 
                           n1929);
   U4005 : AOI21_X1 port map( A1 => n16688, A2 => n16554, B => n24219, ZN => 
                           n12357);
   U4006 : CLKBUF_X12 port map( I => n16554, Z => n26916);
   U4029 : NOR2_X1 port map( A1 => n1323, A2 => n7868, ZN => n17547);
   U4032 : OR2_X2 port map( A1 => n10438, A2 => n4735, Z => n7561);
   U4049 : OR3_X2 port map( A1 => n11208, A2 => n12211, A3 => n8313, Z => n5309
                           );
   U4077 : NAND2_X1 port map( A1 => n16018, A2 => n16181, ZN => n5428);
   U4079 : NOR3_X1 port map( A1 => n16181, A2 => n489, A3 => n29658, ZN => 
                           n9631);
   U4080 : OAI22_X1 port map( A1 => n19333, A2 => n28404, B1 => n19331, B2 => 
                           n8862, ZN => n26503);
   U4090 : NAND2_X1 port map( A1 => n1094, A2 => n13412, ZN => n1640);
   U4120 : BUF_X4 port map( I => n15536, Z => n29307);
   U4122 : INV_X1 port map( I => n23438, ZN => n29231);
   U4124 : INV_X1 port map( I => n12652, ZN => n5157);
   U4136 : INV_X1 port map( I => n18283, ZN => n12837);
   U4139 : BUF_X2 port map( I => n18283, Z => n18617);
   U4140 : AOI21_X2 port map( A1 => n28278, A2 => n34046, B => n11890, ZN => 
                           n12794);
   U4149 : NAND2_X1 port map( A1 => n16688, A2 => n24220, ZN => n23624);
   U4175 : INV_X1 port map( I => n21551, ZN => n30511);
   U4182 : OAI21_X2 port map( A1 => n20057, A2 => n20058, B => n19867, ZN => 
                           n27840);
   U4188 : OAI22_X1 port map( A1 => n11199, A2 => n20154, B1 => n11198, B2 => 
                           n19926, ZN => n19918);
   U4194 : NOR2_X1 port map( A1 => n20157, A2 => n20156, ZN => n16795);
   U4202 : NAND3_X1 port map( A1 => n30934, A2 => n33687, A3 => n34139, ZN => 
                           n11919);
   U4211 : OAI21_X1 port map( A1 => n18567, A2 => n34139, B => n12154, ZN => 
                           n12153);
   U4225 : NAND2_X1 port map( A1 => n23956, A2 => n23955, ZN => n14521);
   U4249 : OR3_X2 port map( A1 => n25121, A2 => n1567, A3 => n16293, Z => 
                           n24889);
   U4288 : OAI22_X1 port map( A1 => n11311, A2 => n781, B1 => n20447, B2 => 
                           n26424, ZN => n7955);
   U4338 : INV_X2 port map( I => n20756, ZN => n6218);
   U4345 : INV_X1 port map( I => n27077, ZN => n1382);
   U4356 : NAND3_X1 port map( A1 => n15646, A2 => n24780, A3 => n24983, ZN => 
                           n4216);
   U4357 : INV_X2 port map( I => n24780, ZN => n15084);
   U4371 : CLKBUF_X4 port map( I => n25146, Z => n1786);
   U4385 : NOR2_X1 port map( A1 => n21832, A2 => n5170, ZN => n12161);
   U4413 : NOR2_X1 port map( A1 => n14839, A2 => n24163, ZN => n29568);
   U4415 : INV_X1 port map( I => n23333, ZN => n28323);
   U4434 : NAND2_X2 port map( A1 => n583, A2 => n9288, ZN => n30530);
   U4450 : NOR2_X2 port map( A1 => n25985, A2 => n33335, ZN => n19146);
   U4462 : NOR2_X1 port map( A1 => n22361, A2 => n4135, ZN => n26609);
   U4468 : AND2_X1 port map( A1 => n31637, A2 => n22361, Z => n29430);
   U4472 : INV_X2 port map( I => n20450, ZN => n20378);
   U4479 : OR2_X2 port map( A1 => n32055, A2 => n9064, Z => n22600);
   U4483 : INV_X1 port map( I => n18184, ZN => n21808);
   U4487 : INV_X1 port map( I => n18411, ZN => n18848);
   U4488 : BUF_X2 port map( I => n18411, Z => n18846);
   U4491 : INV_X1 port map( I => n18078, ZN => n9783);
   U4504 : NAND2_X1 port map( A1 => n23079, A2 => n22885, ZN => n31712);
   U4514 : NOR2_X1 port map( A1 => n20160, A2 => n14138, ZN => n26555);
   U4517 : OAI22_X1 port map( A1 => n4683, A2 => n1146, B1 => n8010, B2 => 
                           n5049, ZN => n8175);
   U4522 : BUF_X4 port map( I => n31951, Z => n19926);
   U4525 : NAND2_X1 port map( A1 => n5889, A2 => n27921, ZN => n19363);
   U4528 : AND2_X2 port map( A1 => n15343, A2 => n22521, Z => n22522);
   U4540 : INV_X1 port map( I => n21198, ZN => n21405);
   U4563 : INV_X1 port map( I => n30637, ZN => n16190);
   U4565 : NAND2_X1 port map( A1 => n15692, A2 => n23877, ZN => n9975);
   U4573 : NOR2_X1 port map( A1 => n4820, A2 => n23742, ZN => n30172);
   U4582 : NAND2_X1 port map( A1 => n13759, A2 => n8087, ZN => n13785);
   U4583 : AOI21_X1 port map( A1 => n8087, A2 => n33515, B => n9688, ZN => 
                           n13830);
   U4589 : OAI21_X1 port map( A1 => n13509, A2 => n17313, B => n26133, ZN => 
                           n14955);
   U4601 : NAND2_X1 port map( A1 => n19057, A2 => n7345, ZN => n8092);
   U4613 : AND2_X2 port map( A1 => n25894, A2 => n9125, Z => n28910);
   U4624 : AND2_X2 port map( A1 => n8899, A2 => n595, Z => n7721);
   U4636 : NAND2_X1 port map( A1 => n20529, A2 => n30637, ZN => n20528);
   U4653 : NOR2_X1 port map( A1 => n20529, A2 => n30637, ZN => n20196);
   U4655 : NAND2_X1 port map( A1 => n19088, A2 => n18990, ZN => n31352);
   U4667 : CLKBUF_X12 port map( I => n18869, Z => n29308);
   U4668 : BUF_X4 port map( I => n18869, Z => n29309);
   U4685 : INV_X1 port map( I => n5414, ZN => n31059);
   U4697 : INV_X2 port map( I => n5440, ZN => n6072);
   U4699 : NAND2_X1 port map( A1 => n5440, A2 => n5441, ZN => n11334);
   U4705 : NAND2_X1 port map( A1 => n22586, A2 => n33320, ZN => n22587);
   U4709 : NAND2_X1 port map( A1 => n12421, A2 => n2821, ZN => n19830);
   U4735 : INV_X1 port map( I => n27503, ZN => n21080);
   U4740 : NAND2_X1 port map( A1 => n29655, A2 => n27931, ZN => n14460);
   U4743 : OR2_X2 port map( A1 => n8469, A2 => n4568, Z => n8467);
   U4746 : NAND2_X1 port map( A1 => n5433, A2 => n1168, ZN => n13058);
   U4758 : NAND2_X1 port map( A1 => n5433, A2 => n17670, ZN => n4744);
   U4767 : INV_X1 port map( I => n12040, ZN => n19987);
   U4776 : BUF_X4 port map( I => n2041, Z => n29312);
   U4782 : NAND2_X1 port map( A1 => n16621, A2 => n24180, ZN => n27786);
   U4783 : CLKBUF_X12 port map( I => n30410, Z => n29313);
   U4789 : BUF_X4 port map( I => n30410, Z => n29314);
   U4795 : CLKBUF_X4 port map( I => n4669, Z => n29315);
   U4798 : CLKBUF_X12 port map( I => n16354, Z => n14130);
   U4817 : AOI21_X1 port map( A1 => n21357, A2 => n12037, B => n21358, ZN => 
                           n30226);
   U4823 : NOR2_X1 port map( A1 => n12863, A2 => n10903, ZN => n12663);
   U4827 : OAI22_X1 port map( A1 => n7497, A2 => n10903, B1 => n7495, B2 => 
                           n12863, ZN => n27215);
   U4846 : AOI22_X1 port map( A1 => n18595, A2 => n18731, B1 => n18845, B2 => 
                           n18596, ZN => n26458);
   U4853 : CLKBUF_X4 port map( I => n20064, Z => n16630);
   U4873 : INV_X1 port map( I => n16022, ZN => n6360);
   U4914 : NOR2_X1 port map( A1 => n22865, A2 => n4084, ZN => n12578);
   U4919 : INV_X2 port map( I => n4084, ZN => n10641);
   U4920 : BUF_X4 port map( I => n29321, Z => n29322);
   U4921 : NAND3_X1 port map( A1 => n16490, A2 => n32172, A3 => n15089, ZN => 
                           n21882);
   U4923 : OAI21_X1 port map( A1 => n22678, A2 => n15089, B => n16570, ZN => 
                           n15911);
   U4926 : NOR2_X1 port map( A1 => n16563, A2 => n2839, ZN => n23757);
   U4931 : INV_X2 port map( I => n432, ZN => n17472);
   U4933 : NOR2_X1 port map( A1 => n432, A2 => n16194, ZN => n31557);
   U4955 : NAND2_X1 port map( A1 => n20630, A2 => n14564, ZN => n30496);
   U4958 : NOR2_X1 port map( A1 => n30326, A2 => n12827, ZN => n13332);
   U4974 : OAI22_X1 port map( A1 => n6671, A2 => n12517, B1 => n19908, B2 => 
                           n16298, ZN => n6377);
   U4975 : CLKBUF_X4 port map( I => n7552, Z => n53);
   U4986 : NOR2_X1 port map( A1 => n29253, A2 => n17967, ZN => n8108);
   U4998 : INV_X2 port map( I => n17967, ZN => n7804);
   U5020 : BUF_X2 port map( I => n20152, Z => n8259);
   U5037 : NAND2_X1 port map( A1 => n29118, A2 => n26969, ZN => n9441);
   U5064 : INV_X2 port map( I => n5696, ZN => n14183);
   U5070 : NAND2_X1 port map( A1 => n6453, A2 => n3103, ZN => n14555);
   U5078 : INV_X2 port map( I => n21870, ZN => n12394);
   U5098 : NOR2_X1 port map( A1 => n18078, A2 => n6679, ZN => n20223);
   U5110 : CLKBUF_X12 port map( I => n18586, Z => n18587);
   U5121 : OR3_X2 port map( A1 => n27619, A2 => n26445, A3 => n27336, Z => n615
                           );
   U5129 : INV_X2 port map( I => n27726, ZN => n826);
   U5131 : NAND2_X1 port map( A1 => n29302, A2 => n16194, ZN => n21494);
   U5147 : NOR2_X1 port map( A1 => n21211, A2 => n16906, ZN => n12066);
   U5149 : NAND2_X1 port map( A1 => n14402, A2 => n7287, ZN => n31790);
   U5158 : BUF_X4 port map( I => n22909, Z => n29329);
   U5165 : NOR2_X1 port map( A1 => n16249, A2 => n18820, ZN => n12976);
   U5169 : NOR2_X1 port map( A1 => n9484, A2 => n2958, ZN => n9483);
   U5188 : NAND2_X1 port map( A1 => n31837, A2 => n11789, ZN => n8279);
   U5196 : INV_X1 port map( I => n11789, ZN => n24222);
   U5198 : BUF_X2 port map( I => n2600, Z => n29331);
   U5204 : NAND3_X1 port map( A1 => n13751, A2 => n5915, A3 => n14183, ZN => 
                           n3160);
   U5228 : CLKBUF_X12 port map( I => n18763, Z => n16559);
   U5232 : NAND2_X1 port map( A1 => n28028, A2 => n20534, ZN => n6925);
   U5265 : NAND2_X1 port map( A1 => n1239, A2 => n24262, ZN => n16574);
   U5268 : INV_X2 port map( I => n24262, ZN => n26950);
   U5278 : INV_X1 port map( I => n17015, ZN => n23785);
   U5282 : INV_X1 port map( I => n17927, ZN => n830);
   U5291 : OAI22_X1 port map( A1 => n15944, A2 => n25848, B1 => n25857, B2 => 
                           n14915, ZN => n30808);
   U5293 : NAND2_X1 port map( A1 => n27057, A2 => n12049, ZN => n30831);
   U5308 : INV_X2 port map( I => n24965, ZN => n24969);
   U5325 : NAND2_X1 port map( A1 => n29593, A2 => n7688, ZN => n4900);
   U5334 : INV_X1 port map( I => n29594, ZN => n29593);
   U5348 : NAND2_X1 port map( A1 => n9857, A2 => n9859, ZN => n9856);
   U5384 : INV_X1 port map( I => n24878, ZN => n31602);
   U5387 : BUF_X2 port map( I => n25762, Z => n17120);
   U5411 : CLKBUF_X1 port map( I => n679, Z => n30308);
   U5415 : INV_X1 port map( I => n24390, ZN => n30883);
   U5419 : INV_X1 port map( I => n14727, ZN => n24660);
   U5431 : NAND2_X1 port map( A1 => n16901, A2 => n29512, ZN => n13660);
   U5446 : AND2_X1 port map( A1 => n24244, A2 => n1235, Z => n29387);
   U5451 : NOR2_X1 port map( A1 => n15996, A2 => n11200, ZN => n31033);
   U5455 : AND3_X1 port map( A1 => n6003, A2 => n33868, A3 => n24095, Z => 
                           n29397);
   U5466 : OR2_X1 port map( A1 => n30270, A2 => n31772, Z => n273);
   U5469 : NOR2_X1 port map( A1 => n27826, A2 => n9323, ZN => n27971);
   U5502 : CLKBUF_X2 port map( I => n14770, Z => n29985);
   U5503 : INV_X1 port map( I => n9368, ZN => n31544);
   U5506 : CLKBUF_X2 port map( I => n4655, Z => n31355);
   U5511 : CLKBUF_X2 port map( I => n15663, Z => n29655);
   U5525 : AND2_X1 port map( A1 => n27392, A2 => n29131, Z => n30283);
   U5540 : INV_X1 port map( I => n27184, ZN => n31615);
   U5547 : INV_X1 port map( I => n29590, ZN => n12399);
   U5550 : NAND2_X1 port map( A1 => n7475, A2 => n14133, ZN => n30886);
   U5553 : OAI21_X1 port map( A1 => n7088, A2 => n26965, B => n2447, ZN => 
                           n31247);
   U5556 : NAND2_X1 port map( A1 => n18152, A2 => n23940, ZN => n29708);
   U5565 : AND2_X1 port map( A1 => n27474, A2 => n30408, Z => n29368);
   U5570 : INV_X1 port map( I => n6309, ZN => n23954);
   U5583 : NAND2_X1 port map( A1 => n13291, A2 => n31916, ZN => n31601);
   U5586 : INV_X1 port map( I => n299, ZN => n30408);
   U5619 : CLKBUF_X4 port map( I => n27996, Z => n31491);
   U5621 : NAND2_X1 port map( A1 => n14417, A2 => n13977, ZN => n29614);
   U5629 : NOR2_X1 port map( A1 => n30868, A2 => n10296, ZN => n17464);
   U5632 : NOR2_X1 port map( A1 => n1277, A2 => n15577, ZN => n30968);
   U5633 : AOI22_X1 port map( A1 => n23104, A2 => n26724, B1 => n5448, B2 => 
                           n22582, ZN => n22591);
   U5634 : NAND3_X1 port map( A1 => n15391, A2 => n22873, A3 => n15390, ZN => 
                           n393);
   U5647 : BUF_X2 port map( I => n849, Z => n30437);
   U5659 : NAND2_X1 port map( A1 => n31363, A2 => n10288, ZN => n6540);
   U5666 : NAND2_X1 port map( A1 => n31315, A2 => n22680, ZN => n4156);
   U5699 : CLKBUF_X2 port map( I => n9953, Z => n31019);
   U5705 : BUF_X2 port map( I => n27160, Z => n22524);
   U5712 : CLKBUF_X4 port map( I => n11110, Z => n29335);
   U5720 : INV_X1 port map( I => n22213, ZN => n31331);
   U5723 : OAI21_X1 port map( A1 => n29408, A2 => n21475, B => n21936, ZN => 
                           n21481);
   U5726 : AND2_X1 port map( A1 => n21477, A2 => n28895, Z => n29408);
   U5729 : NAND2_X1 port map( A1 => n7813, A2 => n29796, ZN => n30622);
   U5732 : NOR2_X1 port map( A1 => n29433, A2 => n29943, ZN => n3908);
   U5734 : NOR2_X1 port map( A1 => n21785, A2 => n7553, ZN => n30374);
   U5741 : CLKBUF_X4 port map( I => n1917, Z => n31616);
   U5758 : NOR2_X1 port map( A1 => n21282, A2 => n28618, ZN => n31073);
   U5759 : NAND2_X1 port map( A1 => n31557, A2 => n31458, ZN => n31572);
   U5760 : NOR2_X1 port map( A1 => n9601, A2 => n13213, ZN => n13212);
   U5764 : NAND2_X1 port map( A1 => n21278, A2 => n29827, ZN => n21279);
   U5767 : INV_X2 port map( I => n5863, ZN => n7813);
   U5768 : NAND2_X1 port map( A1 => n21, A2 => n30033, ZN => n21539);
   U5774 : CLKBUF_X2 port map( I => n12535, Z => n30243);
   U5776 : NAND2_X1 port map( A1 => n12725, A2 => n31334, ZN => n12724);
   U5779 : CLKBUF_X4 port map( I => n6533, Z => n31765);
   U5819 : INV_X1 port map( I => n31484, ZN => n16925);
   U5821 : INV_X1 port map( I => n2802, ZN => n29931);
   U5822 : AND3_X1 port map( A1 => n21733, A2 => n26474, A3 => n13872, Z => 
                           n29433);
   U5824 : NAND2_X1 port map( A1 => n16257, A2 => n16258, ZN => n29711);
   U5836 : INV_X1 port map( I => n21316, ZN => n14230);
   U5844 : OAI21_X1 port map( A1 => n12325, A2 => n3933, B => n21400, ZN => 
                           n15113);
   U5852 : NOR2_X1 port map( A1 => n6277, A2 => n21302, ZN => n18207);
   U5853 : NAND2_X1 port map( A1 => n21167, A2 => n16905, ZN => n30005);
   U5854 : INV_X1 port map( I => n20880, ZN => n30006);
   U5857 : NAND2_X1 port map( A1 => n1334, A2 => n31476, ZN => n31475);
   U5871 : BUF_X2 port map( I => n3106, Z => n26635);
   U5874 : NAND2_X1 port map( A1 => n17439, A2 => n925, ZN => n1785);
   U5880 : INV_X1 port map( I => n20972, ZN => n29810);
   U5884 : BUF_X2 port map( I => n21220, Z => n15149);
   U5890 : INV_X1 port map( I => n2756, ZN => n29833);
   U5891 : INV_X1 port map( I => n20978, ZN => n31235);
   U5919 : CLKBUF_X2 port map( I => n8728, Z => n29838);
   U5926 : OR2_X1 port map( A1 => n20247, A2 => n7394, Z => n1684);
   U5932 : NOR2_X1 port map( A1 => n30915, A2 => n20317, ZN => n17732);
   U5934 : NOR2_X1 port map( A1 => n30414, A2 => n30413, ZN => n20282);
   U5937 : INV_X1 port map( I => n1354, ZN => n31470);
   U5938 : INV_X1 port map( I => n931, ZN => n30545);
   U5945 : CLKBUF_X2 port map( I => n6531, Z => n31863);
   U5947 : CLKBUF_X2 port map( I => n9115, Z => n30878);
   U5951 : CLKBUF_X2 port map( I => n4693, Z => n31873);
   U5952 : INV_X2 port map( I => n6996, ZN => n16182);
   U5998 : CLKBUF_X2 port map( I => n19849, Z => n31742);
   U6016 : CLKBUF_X4 port map( I => n17711, Z => n30355);
   U6019 : INV_X4 port map( I => n29882, ZN => n20010);
   U6041 : CLKBUF_X2 port map( I => n19389, Z => n31410);
   U6043 : NAND2_X1 port map( A1 => n30710, A2 => n3341, ZN => n19239);
   U6044 : NOR2_X1 port map( A1 => n19011, A2 => n7995, ZN => n30401);
   U6045 : INV_X1 port map( I => n19205, ZN => n9316);
   U6061 : BUF_X2 port map( I => n11477, Z => n4210);
   U6063 : BUF_X4 port map( I => n13320, Z => n25968);
   U6069 : AOI21_X1 port map( A1 => n12132, A2 => n18701, B => n29366, ZN => 
                           n8551);
   U6071 : INV_X1 port map( I => n18462, ZN => n31903);
   U6076 : OAI21_X1 port map( A1 => n17478, A2 => n31428, B => n31427, ZN => 
                           n12116);
   U6082 : OAI21_X1 port map( A1 => n8411, A2 => n16614, B => n18307, ZN => 
                           n30866);
   U6085 : INV_X1 port map( I => n9836, ZN => n18338);
   U6092 : NAND3_X1 port map( A1 => n3152, A2 => n2990, A3 => n18893, ZN => 
                           n30919);
   U6095 : CLKBUF_X2 port map( I => n18018, Z => n31115);
   U6102 : INV_X1 port map( I => n24966, ZN => n30881);
   U6110 : INV_X1 port map( I => n24923, ZN => n31513);
   U6117 : BUF_X2 port map( I => n18557, Z => n28987);
   U6124 : INV_X1 port map( I => n25450, ZN => n29851);
   U6130 : INV_X1 port map( I => n16520, ZN => n30557);
   U6132 : CLKBUF_X2 port map( I => n8317, Z => n31724);
   U6136 : INV_X1 port map( I => n25195, ZN => n30954);
   U6137 : INV_X1 port map( I => n16653, ZN => n30018);
   U6163 : NAND2_X1 port map( A1 => n18730, A2 => n18846, ZN => n6313);
   U6164 : OAI21_X1 port map( A1 => n16370, A2 => n962, B => n6783, ZN => 
                           n12199);
   U6165 : NAND2_X1 port map( A1 => n1186, A2 => n18822, ZN => n16247);
   U6183 : NOR2_X1 port map( A1 => n18835, A2 => n32901, ZN => n13013);
   U6195 : NOR2_X1 port map( A1 => n10578, A2 => n11941, ZN => n2734);
   U6201 : BUF_X2 port map( I => n16766, Z => n28238);
   U6205 : INV_X1 port map( I => n7320, ZN => n9174);
   U6224 : CLKBUF_X2 port map( I => n29061, Z => n28548);
   U6227 : INV_X1 port map( I => n9514, ZN => n17792);
   U6228 : NAND2_X1 port map( A1 => n18792, A2 => n13514, ZN => n29684);
   U6240 : NAND2_X1 port map( A1 => n19315, A2 => n11000, ZN => n10999);
   U6241 : NOR2_X1 port map( A1 => n10857, A2 => n13568, ZN => n10856);
   U6246 : INV_X2 port map( I => n19154, ZN => n2040);
   U6247 : NAND2_X1 port map( A1 => n7415, A2 => n14332, ZN => n19247);
   U6271 : CLKBUF_X2 port map( I => n7134, Z => n1386);
   U6273 : INV_X2 port map( I => n27807, ZN => n26518);
   U6274 : NAND2_X1 port map( A1 => n27077, A2 => n5789, ZN => n19210);
   U6277 : INV_X1 port map( I => n6488, ZN => n1367);
   U6280 : INV_X1 port map( I => n16429, ZN => n31750);
   U6281 : NAND2_X1 port map( A1 => n19190, A2 => n19261, ZN => n28540);
   U6289 : NAND2_X1 port map( A1 => n15239, A2 => n19218, ZN => n19352);
   U6297 : OAI21_X1 port map( A1 => n1630, A2 => n19176, B => n12993, ZN => 
                           n1629);
   U6300 : AOI21_X1 port map( A1 => n18908, A2 => n26181, B => n16353, ZN => 
                           n18909);
   U6304 : INV_X1 port map( I => n2499, ZN => n29727);
   U6306 : INV_X1 port map( I => n19343, ZN => n30258);
   U6307 : INV_X1 port map( I => n15913, ZN => n17220);
   U6317 : NAND2_X1 port map( A1 => n20000, A2 => n14457, ZN => n13654);
   U6325 : NAND2_X1 port map( A1 => n1043, A2 => n11350, ZN => n5642);
   U6327 : CLKBUF_X2 port map( I => n20011, Z => n30794);
   U6328 : INV_X1 port map( I => n30600, ZN => n8687);
   U6336 : OAI21_X1 port map( A1 => n15192, A2 => n19874, B => n149, ZN => 
                           n12669);
   U6357 : NAND2_X1 port map( A1 => n29373, A2 => n31694, ZN => n31693);
   U6358 : NAND2_X1 port map( A1 => n28021, A2 => n20068, ZN => n28020);
   U6371 : NAND2_X1 port map( A1 => n5999, A2 => n20033, ZN => n4201);
   U6379 : NAND2_X1 port map( A1 => n20017, A2 => n15278, ZN => n30072);
   U6388 : INV_X1 port map( I => n20107, ZN => n31164);
   U6395 : OAI21_X1 port map( A1 => n19808, A2 => n15278, B => n8816, ZN => 
                           n10742);
   U6396 : NAND2_X1 port map( A1 => n20090, A2 => n19879, ZN => n19881);
   U6398 : INV_X2 port map( I => n34151, ZN => n729);
   U6423 : NAND2_X1 port map( A1 => n15953, A2 => n9484, ZN => n30464);
   U6429 : CLKBUF_X2 port map( I => n10414, Z => n3915);
   U6432 : NAND3_X1 port map( A1 => n2879, A2 => n31504, A3 => n20524, ZN => 
                           n31563);
   U6433 : AND2_X1 port map( A1 => n17647, A2 => n6230, Z => n29409);
   U6437 : NAND2_X1 port map( A1 => n28288, A2 => n6997, ZN => n7056);
   U6440 : INV_X1 port map( I => n20536, ZN => n20535);
   U6442 : AOI21_X1 port map( A1 => n33288, A2 => n20472, B => n32504, ZN => 
                           n20165);
   U6446 : INV_X2 port map( I => n8903, ZN => n1349);
   U6450 : NAND2_X1 port map( A1 => n9115, A2 => n6996, ZN => n12583);
   U6452 : NAND2_X1 port map( A1 => n8702, A2 => n9854, ZN => n31496);
   U6453 : OAI21_X1 port map( A1 => n818, A2 => n710, B => n20334, ZN => n20048
                           );
   U6454 : NOR2_X1 port map( A1 => n10718, A2 => n10716, ZN => n10715);
   U6456 : NAND2_X1 port map( A1 => n32068, A2 => n20452, ZN => n15662);
   U6468 : OAI21_X1 port map( A1 => n1160, A2 => n27621, B => n27620, ZN => 
                           n2754);
   U6478 : INV_X1 port map( I => n20863, ZN => n29734);
   U6490 : NOR2_X1 port map( A1 => n21060, A2 => n4568, ZN => n10921);
   U6491 : NAND2_X1 port map( A1 => n29255, A2 => n26712, ZN => n6337);
   U6493 : NAND2_X1 port map( A1 => n21203, A2 => n3933, ZN => n21204);
   U6495 : INV_X1 port map( I => n29802, ZN => n13700);
   U6496 : AND2_X1 port map( A1 => n4145, A2 => n32452, Z => n29361);
   U6502 : NAND2_X1 port map( A1 => n8197, A2 => n924, ZN => n1555);
   U6505 : INV_X1 port map( I => n31197, ZN => n30816);
   U6510 : NOR2_X1 port map( A1 => n21113, A2 => n1332, ZN => n27539);
   U6516 : NOR2_X1 port map( A1 => n18218, A2 => n31030, ZN => n7845);
   U6523 : NAND2_X1 port map( A1 => n14721, A2 => n8115, ZN => n14087);
   U6524 : NAND3_X1 port map( A1 => n20883, A2 => n21369, A3 => n1148, ZN => 
                           n20884);
   U6531 : NOR2_X1 port map( A1 => n21358, A2 => n11814, ZN => n6307);
   U6541 : NAND2_X1 port map( A1 => n21211, A2 => n13319, ZN => n20874);
   U6547 : NAND2_X1 port map( A1 => n30227, A2 => n30226, ZN => n30225);
   U6552 : INV_X1 port map( I => n21147, ZN => n17217);
   U6561 : NOR2_X1 port map( A1 => n3140, A2 => n30885, ZN => n27836);
   U6562 : AOI21_X1 port map( A1 => n16755, A2 => n27955, B => n21400, ZN => 
                           n16257);
   U6563 : NAND2_X1 port map( A1 => n4293, A2 => n31613, ZN => n31612);
   U6565 : AOI21_X1 port map( A1 => n30006, A2 => n30005, B => n21209, ZN => 
                           n29214);
   U6572 : INV_X1 port map( I => n11861, ZN => n31653);
   U6578 : AOI21_X1 port map( A1 => n10345, A2 => n16519, B => n777, ZN => 
                           n10344);
   U6579 : INV_X1 port map( I => n16605, ZN => n30007);
   U6597 : INV_X1 port map( I => n2576, ZN => n21682);
   U6601 : NAND2_X1 port map( A1 => n31475, A2 => n31474, ZN => n21274);
   U6603 : INV_X2 port map( I => n5795, ZN => n1135);
   U6617 : NAND2_X1 port map( A1 => n18055, A2 => n21, ZN => n30608);
   U6634 : OAI21_X1 port map( A1 => n21696, A2 => n30769, B => n1013, ZN => 
                           n21699);
   U6651 : NAND2_X1 port map( A1 => n15748, A2 => n26513, ZN => n10232);
   U6663 : INV_X1 port map( I => n10519, ZN => n22244);
   U6664 : INV_X2 port map( I => n22092, ZN => n14289);
   U6671 : INV_X1 port map( I => n1716, ZN => n29896);
   U6674 : OAI21_X1 port map( A1 => n13371, A2 => n22220, B => n13370, ZN => 
                           n22246);
   U6695 : INV_X1 port map( I => n22565, ZN => n22468);
   U6696 : NOR3_X1 port map( A1 => n22543, A2 => n10757, A3 => n252, ZN => 
                           n7236);
   U6716 : CLKBUF_X4 port map( I => n632, Z => n14227);
   U6730 : NOR2_X1 port map( A1 => n22682, A2 => n9802, ZN => n3455);
   U6732 : NAND3_X1 port map( A1 => n900, A2 => n11920, A3 => n22476, ZN => 
                           n14017);
   U6744 : NAND2_X1 port map( A1 => n29335, A2 => n22435, ZN => n31634);
   U6748 : NOR2_X1 port map( A1 => n16986, A2 => n9370, ZN => n22026);
   U6750 : OAI21_X1 port map( A1 => n29461, A2 => n15635, B => n29222, ZN => 
                           n28894);
   U6753 : NOR2_X1 port map( A1 => n29508, A2 => n22574, ZN => n10121);
   U6769 : INV_X1 port map( I => n22560, ZN => n31315);
   U6781 : AOI22_X1 port map( A1 => n12281, A2 => n10288, B1 => n22542, B2 => 
                           n22397, ZN => n22299);
   U6791 : NAND3_X1 port map( A1 => n29222, A2 => n18073, A3 => n10680, ZN => 
                           n12472);
   U6793 : NAND2_X1 port map( A1 => n15033, A2 => n8314, ZN => n15032);
   U6797 : INV_X2 port map( I => n7004, ZN => n14131);
   U6808 : NAND2_X1 port map( A1 => n2635, A2 => n13191, ZN => n2638);
   U6818 : NAND2_X1 port map( A1 => n14131, A2 => n23106, ZN => n15280);
   U6835 : OAI22_X1 port map( A1 => n22502, A2 => n32449, B1 => n13874, B2 => 
                           n30014, ZN => n26772);
   U6847 : NAND3_X1 port map( A1 => n29610, A2 => n4113, A3 => n22791, ZN => 
                           n22776);
   U6848 : AOI21_X1 port map( A1 => n3783, A2 => n28801, B => n30247, ZN => 
                           n9075);
   U6852 : INV_X1 port map( I => n9185, ZN => n31056);
   U6857 : CLKBUF_X2 port map( I => n8762, Z => n29235);
   U6863 : INV_X1 port map( I => n14464, ZN => n29675);
   U6864 : INV_X1 port map( I => n23331, ZN => n23509);
   U6866 : NAND2_X1 port map( A1 => n23873, A2 => n23872, ZN => n23874);
   U6867 : AOI21_X1 port map( A1 => n27298, A2 => n8967, B => n22957, ZN => 
                           n22904);
   U6869 : INV_X1 port map( I => n23742, ZN => n23768);
   U6877 : INV_X1 port map( I => n23778, ZN => n975);
   U6883 : INV_X1 port map( I => n8045, ZN => n11960);
   U6884 : NAND2_X1 port map( A1 => n1252, A2 => n23603, ZN => n14039);
   U6886 : NOR2_X1 port map( A1 => n23611, A2 => n33144, ZN => n1892);
   U6887 : NAND2_X1 port map( A1 => n23647, A2 => n26790, ZN => n28303);
   U6891 : INV_X1 port map( I => n28615, ZN => n23691);
   U6896 : INV_X2 port map( I => n9828, ZN => n16686);
   U6900 : CLKBUF_X2 port map( I => n23924, Z => n1101);
   U6903 : OAI21_X1 port map( A1 => n15187, A2 => n15186, B => n23691, ZN => 
                           n23572);
   U6907 : NAND3_X1 port map( A1 => n23799, A2 => n23798, A3 => n23800, ZN => 
                           n23802);
   U6908 : NAND2_X1 port map( A1 => n23855, A2 => n652, ZN => n23856);
   U6912 : INV_X2 port map( I => n23603, ZN => n23776);
   U6923 : NAND2_X1 port map( A1 => n793, A2 => n6713, ZN => n5132);
   U6928 : AND2_X1 port map( A1 => n11438, A2 => n29748, Z => n29379);
   U6936 : NAND2_X1 port map( A1 => n23707, A2 => n23786, ZN => n23711);
   U6947 : NOR2_X1 port map( A1 => n30283, A2 => n24087, ZN => n11107);
   U6964 : OAI22_X1 port map( A1 => n7068, A2 => n24196, B1 => n13048, B2 => 
                           n969, ZN => n13324);
   U6972 : AND2_X1 port map( A1 => n24234, A2 => n7581, Z => n8004);
   U6978 : CLKBUF_X4 port map( I => n13508, Z => n7828);
   U6981 : INV_X1 port map( I => n14897, ZN => n1226);
   U6988 : INV_X1 port map( I => n24427, ZN => n29639);
   U6992 : NAND2_X1 port map( A1 => n16113, A2 => n25870, ZN => n24732);
   U7006 : CLKBUF_X4 port map( I => n16757, Z => n11090);
   U7011 : NAND2_X1 port map( A1 => n26917, A2 => n15770, ZN => n25396);
   U7015 : NAND2_X1 port map( A1 => n25870, A2 => n4993, ZN => n11718);
   U7023 : NAND2_X1 port map( A1 => n419, A2 => n11366, ZN => n16339);
   U7027 : AOI21_X1 port map( A1 => n24955, A2 => n24956, B => n24947, ZN => 
                           n29664);
   U7029 : OAI21_X1 port map( A1 => n25204, A2 => n32601, B => n25205, ZN => 
                           n18259);
   U7031 : CLKBUF_X1 port map( I => n11974, Z => n4245);
   U7034 : INV_X1 port map( I => n29664, ZN => n29663);
   U7056 : CLKBUF_X1 port map( I => n25258, Z => n27429);
   U7060 : INV_X2 port map( I => n5128, ZN => n786);
   U7062 : CLKBUF_X1 port map( I => Key(158), Z => n16705);
   U7071 : XNOR2_X1 port map( A1 => n5150, A2 => n14648, ZN => n29341);
   U7074 : XNOR2_X1 port map( A1 => n19580, A2 => n32796, ZN => n29343);
   U7075 : XNOR2_X1 port map( A1 => n23271, A2 => n16653, ZN => n29344);
   U7084 : XNOR2_X1 port map( A1 => n27423, A2 => n25108, ZN => n29345);
   U7086 : XNOR2_X1 port map( A1 => n24635, A2 => n16654, ZN => n29346);
   U7087 : XNOR2_X1 port map( A1 => n16237, A2 => n28711, ZN => n29347);
   U7088 : XNOR2_X1 port map( A1 => n24617, A2 => n25735, ZN => n29348);
   U7089 : OR2_X1 port map( A1 => n32021, A2 => n31551, Z => n29349);
   U7092 : AND2_X1 port map( A1 => n24293, A2 => n5632, Z => n29352);
   U7096 : AND2_X1 port map( A1 => n14980, A2 => n31721, Z => n29354);
   U7103 : OR2_X1 port map( A1 => n28293, A2 => n1170, Z => n29359);
   U7112 : AND2_X1 port map( A1 => n20263, A2 => n16146, Z => n29363);
   U7113 : AND2_X1 port map( A1 => n3791, A2 => n6034, Z => n29364);
   U7120 : OR2_X1 port map( A1 => n17694, A2 => n11968, Z => n29367);
   U7132 : OR2_X2 port map( A1 => n28197, A2 => n33232, Z => n29378);
   U7136 : OR2_X1 port map( A1 => n28669, A2 => n10206, Z => n29380);
   U7140 : AND2_X1 port map( A1 => n21779, A2 => n31654, Z => n29383);
   U7144 : OR2_X1 port map( A1 => n26547, A2 => n1596, Z => n29385);
   U7149 : XNOR2_X1 port map( A1 => n24598, A2 => n29416, ZN => n29386);
   U7153 : OR2_X1 port map( A1 => n28833, A2 => n5615, Z => n29389);
   U7155 : OR2_X1 port map( A1 => n22659, A2 => n22658, Z => n29390);
   U7160 : AND2_X1 port map( A1 => n28801, A2 => n11235, Z => n29391);
   U7161 : AND3_X1 port map( A1 => n6012, A2 => n16254, A3 => n23110, Z => 
                           n29392);
   U7163 : AND2_X1 port map( A1 => n17077, A2 => n21579, Z => n29393);
   U7176 : INV_X1 port map( I => n3106, ZN => n4971);
   U7183 : XNOR2_X1 port map( A1 => n17586, A2 => n12082, ZN => n29400);
   U7190 : INV_X1 port map( I => n10124, ZN => n29730);
   U7191 : AND2_X1 port map( A1 => n24436, A2 => n25695, Z => n29402);
   U7192 : OR3_X2 port map( A1 => n7753, A2 => n26622, A3 => n15414, Z => 
                           n29404);
   U7194 : AND2_X1 port map( A1 => n15465, A2 => n21866, Z => n29405);
   U7196 : INV_X1 port map( I => n19283, ZN => n30932);
   U7201 : XNOR2_X1 port map( A1 => n20885, A2 => n25716, ZN => n29412);
   U7202 : XNOR2_X1 port map( A1 => n21043, A2 => n30007, ZN => n29413);
   U7212 : XNOR2_X1 port map( A1 => n34150, A2 => n16533, ZN => n29415);
   U7221 : XNOR2_X1 port map( A1 => n24616, A2 => n24907, ZN => n29416);
   U7222 : XNOR2_X1 port map( A1 => n27167, A2 => n16653, ZN => n29417);
   U7223 : XNOR2_X1 port map( A1 => n34150, A2 => n24065, ZN => n29418);
   U7225 : XNOR2_X1 port map( A1 => n23153, A2 => n14464, ZN => n29420);
   U7229 : AND2_X1 port map( A1 => n17828, A2 => n26160, Z => n29421);
   U7241 : XNOR2_X1 port map( A1 => n19651, A2 => n19658, ZN => n29426);
   U7242 : XNOR2_X1 port map( A1 => n8497, A2 => n513, ZN => n29428);
   U7251 : INV_X2 port map( I => n16132, ZN => n15213);
   U7256 : XNOR2_X1 port map( A1 => n19727, A2 => n18814, ZN => n29441);
   U7257 : XNOR2_X1 port map( A1 => n34082, A2 => n25560, ZN => n29442);
   U7261 : INV_X1 port map( I => n18199, ZN => n19900);
   U7267 : XNOR2_X1 port map( A1 => n4107, A2 => n27361, ZN => n29443);
   U7281 : XNOR2_X1 port map( A1 => n9102, A2 => n9101, ZN => n29445);
   U7288 : XNOR2_X1 port map( A1 => n3665, A2 => n5920, ZN => n29446);
   U7289 : XNOR2_X1 port map( A1 => n10224, A2 => n1365, ZN => n29447);
   U7290 : OR2_X1 port map( A1 => n19226, A2 => n19227, Z => n29448);
   U7293 : XOR2_X1 port map( A1 => n21916, A2 => n21915, Z => n29450);
   U7294 : XOR2_X1 port map( A1 => n30070, A2 => n22094, Z => n29451);
   U7300 : AND2_X2 port map( A1 => n6357, A2 => n9999, Z => n29454);
   U7306 : XNOR2_X1 port map( A1 => n22076, A2 => n24937, ZN => n29457);
   U7310 : XNOR2_X1 port map( A1 => n22154, A2 => n22152, ZN => n29458);
   U7316 : INV_X1 port map( I => n27160, ZN => n28915);
   U7318 : NOR2_X1 port map( A1 => n632, A2 => n22662, ZN => n29461);
   U7324 : XNOR2_X1 port map( A1 => n2899, A2 => n2898, ZN => n29463);
   U7325 : OR2_X1 port map( A1 => n8381, A2 => n5211, Z => n29464);
   U7328 : XNOR2_X1 port map( A1 => n11427, A2 => n11426, ZN => n29467);
   U7334 : INV_X1 port map( I => n12375, ZN => n808);
   U7337 : CLKBUF_X2 port map( I => n16536, Z => n6479);
   U7340 : AND2_X1 port map( A1 => n17394, A2 => n13318, Z => n29469);
   U7351 : INV_X1 port map( I => n5736, ZN => n13281);
   U7352 : XOR2_X1 port map( A1 => n281, A2 => n15515, Z => n29472);
   U7363 : NOR2_X1 port map( A1 => n2855, A2 => n23767, ZN => n29474);
   U7364 : XNOR2_X1 port map( A1 => n24819, A2 => n24632, ZN => n29475);
   U7366 : CLKBUF_X2 port map( I => n24975, Z => n31274);
   U7373 : NAND2_X1 port map( A1 => n10430, A2 => n27072, ZN => n29476);
   U7376 : NAND2_X2 port map( A1 => n2550, A2 => n6409, ZN => n11557);
   U7377 : NOR2_X1 port map( A1 => n4135, A2 => n29325, ZN => n29477);
   U7379 : XOR2_X1 port map( A1 => n19726, A2 => n12718, Z => n29487);
   U7387 : INV_X2 port map( I => n28196, ZN => n7765);
   U7397 : NAND2_X2 port map( A1 => n25170, A2 => n25168, ZN => n28196);
   U7406 : XOR2_X1 port map( A1 => n11423, A2 => n11421, Z => n11451);
   U7408 : NOR3_X1 port map( A1 => n21865, A2 => n21738, A3 => n13652, ZN => 
                           n30806);
   U7414 : OAI21_X2 port map( A1 => n29358, A2 => n29480, B => n8927, ZN => 
                           n9097);
   U7416 : INV_X1 port map( I => n576, ZN => n29480);
   U7419 : INV_X2 port map( I => n33373, ZN => n29481);
   U7430 : NOR3_X1 port map( A1 => n11516, A2 => n9430, A3 => n7993, ZN => 
                           n5777);
   U7435 : XOR2_X1 port map( A1 => n5431, A2 => n30171, Z => n29482);
   U7436 : INV_X4 port map( I => n29483, ZN => n9677);
   U7437 : NOR2_X2 port map( A1 => n10842, A2 => n4267, ZN => n29483);
   U7443 : NAND2_X1 port map( A1 => n896, A2 => n23045, ZN => n22400);
   U7447 : NAND3_X1 port map( A1 => n9962, A2 => n10033, A3 => n24311, ZN => 
                           n12318);
   U7452 : OAI21_X2 port map( A1 => n29654, A2 => n30233, B => n31960, ZN => 
                           n6123);
   U7460 : NOR3_X2 port map( A1 => n11411, A2 => n2085, A3 => n2084, ZN => 
                           n23306);
   U7462 : XOR2_X1 port map( A1 => n29485, A2 => n24486, Z => n31005);
   U7464 : XOR2_X1 port map( A1 => n24488, A2 => n24771, Z => n29485);
   U7465 : XOR2_X1 port map( A1 => n7537, A2 => n24603, Z => n28144);
   U7482 : XOR2_X1 port map( A1 => n27977, A2 => n24564, Z => n17673);
   U7483 : OR2_X1 port map( A1 => n23086, A2 => n4834, Z => n4833);
   U7488 : XOR2_X1 port map( A1 => n29486, A2 => n29487, Z => n8327);
   U7496 : NAND2_X2 port map( A1 => n29488, A2 => n28875, ZN => n25653);
   U7499 : OAI21_X2 port map( A1 => n15355, A2 => n15354, B => n25706, ZN => 
                           n29488);
   U7506 : XOR2_X1 port map( A1 => n29489, A2 => n4761, Z => n8553);
   U7507 : XOR2_X1 port map( A1 => n10087, A2 => n28868, Z => n29489);
   U7514 : XOR2_X1 port map( A1 => n24635, A2 => n10146, Z => n17448);
   U7515 : NOR2_X2 port map( A1 => n7480, A2 => n7483, ZN => n24635);
   U7518 : NAND2_X2 port map( A1 => n13341, A2 => n28356, ZN => n28355);
   U7519 : NAND2_X1 port map( A1 => n26325, A2 => n1318, ZN => n26927);
   U7521 : XOR2_X1 port map( A1 => n7694, A2 => n7693, Z => n29543);
   U7531 : XOR2_X1 port map( A1 => n8714, A2 => n8265, Z => n8713);
   U7534 : XOR2_X1 port map( A1 => n6513, A2 => n9385, Z => n9564);
   U7549 : NOR2_X1 port map( A1 => n29792, A2 => n20549, ZN => n31232);
   U7557 : NAND2_X2 port map( A1 => n11466, A2 => n22783, ZN => n8226);
   U7569 : OAI21_X1 port map( A1 => n22558, A2 => n9630, B => n29495, ZN => 
                           n29494);
   U7570 : INV_X2 port map( I => n994, ZN => n29495);
   U7576 : INV_X1 port map( I => n32957, ZN => n29497);
   U7577 : INV_X2 port map( I => n15365, ZN => n29498);
   U7579 : OR2_X1 port map( A1 => n596, A2 => n14290, Z => n14562);
   U7583 : XOR2_X1 port map( A1 => n14727, A2 => n25549, Z => n31093);
   U7593 : NAND2_X2 port map( A1 => n13633, A2 => n13632, ZN => n14727);
   U7617 : NAND2_X2 port map( A1 => n2394, A2 => n2393, ZN => n22102);
   U7677 : NAND2_X1 port map( A1 => n14661, A2 => n29213, ZN => n19889);
   U7680 : NAND2_X1 port map( A1 => n12042, A2 => n32875, ZN => n24863);
   U7700 : XOR2_X1 port map( A1 => n16886, A2 => n16887, Z => n23156);
   U7711 : OR2_X1 port map( A1 => n9411, A2 => n30668, Z => n7488);
   U7722 : NAND2_X2 port map( A1 => n30856, A2 => n9803, ZN => n20715);
   U7739 : NOR2_X2 port map( A1 => n6533, A2 => n28429, ZN => n16736);
   U7744 : NAND2_X2 port map( A1 => n30483, A2 => n21216, ZN => n6533);
   U7745 : NAND2_X2 port map( A1 => n30139, A2 => n30138, ZN => n20536);
   U7749 : NAND2_X2 port map( A1 => n32075, A2 => n31734, ZN => n21866);
   U7756 : NAND2_X2 port map( A1 => n5743, A2 => n29508, ZN => n29507);
   U7759 : NOR2_X1 port map( A1 => n30666, A2 => n14803, ZN => n29510);
   U7763 : OAI21_X2 port map( A1 => n28510, A2 => n11240, B => n29509, ZN => 
                           n17580);
   U7764 : NAND2_X1 port map( A1 => n10673, A2 => n499, ZN => n29509);
   U7787 : NAND2_X2 port map( A1 => n9123, A2 => n31573, ZN => n4704);
   U7821 : XOR2_X1 port map( A1 => n23504, A2 => n23164, Z => n14370);
   U7828 : NAND2_X1 port map( A1 => n31815, A2 => n21289, ZN => n21291);
   U7837 : NOR2_X1 port map( A1 => n5273, A2 => n17814, ZN => n4204);
   U7841 : NAND2_X1 port map( A1 => n27320, A2 => n27321, ZN => n29517);
   U7847 : NAND2_X2 port map( A1 => n17579, A2 => n16388, ZN => n29518);
   U7862 : XOR2_X1 port map( A1 => n22896, A2 => n23126, Z => n14154);
   U7867 : NAND2_X2 port map( A1 => n30705, A2 => n20163, ZN => n20720);
   U7876 : OR2_X1 port map( A1 => n17405, A2 => n16996, Z => n11508);
   U7877 : OAI21_X2 port map( A1 => n23158, A2 => n22914, B => n29522, ZN => 
                           n14613);
   U7879 : NOR2_X2 port map( A1 => n8943, A2 => n6382, ZN => n29522);
   U7880 : NOR2_X2 port map( A1 => n1350, A2 => n15434, ZN => n29586);
   U7888 : NOR2_X2 port map( A1 => n9962, A2 => n27501, ZN => n15283);
   U7891 : NOR2_X1 port map( A1 => n29714, A2 => n8314, ZN => n13770);
   U7895 : BUF_X2 port map( I => n19049, Z => n29525);
   U7896 : NOR3_X2 port map( A1 => n8378, A2 => n12925, A3 => n21430, ZN => 
                           n7666);
   U7899 : NAND2_X2 port map( A1 => n24461, A2 => n29526, ZN => n31656);
   U7901 : NAND3_X2 port map( A1 => n27118, A2 => n1223, A3 => n18219, ZN => 
                           n29526);
   U7903 : NAND2_X2 port map( A1 => n29527, A2 => n30938, ZN => n16831);
   U7911 : XOR2_X1 port map( A1 => n19476, A2 => n19575, Z => n11093);
   U7915 : OR2_X1 port map( A1 => n29213, A2 => n14661, Z => n4938);
   U7916 : XOR2_X1 port map( A1 => n24826, A2 => n7879, Z => n29534);
   U7920 : XOR2_X1 port map( A1 => n12413, A2 => n19490, Z => n9528);
   U7921 : XOR2_X1 port map( A1 => n19746, A2 => n12442, Z => n19490);
   U7936 : XOR2_X1 port map( A1 => n24090, A2 => n29531, Z => n28816);
   U7940 : XOR2_X1 port map( A1 => n24419, A2 => n29639, Z => n29531);
   U7943 : OAI21_X2 port map( A1 => n15673, A2 => n15672, B => n29532, ZN => 
                           n10371);
   U7956 : NAND2_X2 port map( A1 => n30953, A2 => n25874, ZN => n14737);
   U7958 : OAI22_X1 port map( A1 => n790, A2 => n25900, B1 => n25867, B2 => 
                           n27118, ZN => n25899);
   U7970 : XOR2_X1 port map( A1 => n24807, A2 => n28939, Z => n24439);
   U7974 : AOI22_X1 port map( A1 => n4417, A2 => n25743, B1 => n9414, B2 => 
                           n4416, ZN => n29572);
   U7975 : XOR2_X1 port map( A1 => n29534, A2 => n33927, Z => n26125);
   U7986 : XOR2_X1 port map( A1 => n30767, A2 => n7071, Z => n7825);
   U7987 : XOR2_X1 port map( A1 => n29536, A2 => n22303, Z => n21927);
   U7989 : NAND2_X2 port map( A1 => n21589, A2 => n21588, ZN => n22303);
   U7990 : INV_X2 port map( I => n13553, ZN => n29536);
   U7997 : AOI22_X2 port map( A1 => n23850, A2 => n32477, B1 => n23847, B2 => 
                           n23809, ZN => n3239);
   U7998 : INV_X2 port map( I => n29537, ZN => n10435);
   U8002 : XNOR2_X1 port map( A1 => n26854, A2 => n2064, ZN => n29537);
   U8009 : XOR2_X1 port map( A1 => n29538, A2 => n24824, Z => n31598);
   U8019 : CLKBUF_X12 port map( I => n10248, Z => n29539);
   U8030 : NOR2_X2 port map( A1 => n709, A2 => n31953, ZN => n14794);
   U8032 : INV_X4 port map( I => n10435, ZN => n15278);
   U8040 : OR2_X1 port map( A1 => n33981, A2 => n21832, Z => n10401);
   U8063 : NAND3_X1 port map( A1 => n15146, A2 => n1063, A3 => n1185, ZN => 
                           n9886);
   U8064 : OAI21_X1 port map( A1 => n17497, A2 => n30099, B => n5781, ZN => 
                           n15929);
   U8066 : NOR2_X2 port map( A1 => n6610, A2 => n20209, ZN => n30099);
   U8074 : NOR2_X2 port map( A1 => n12433, A2 => n23753, ZN => n6363);
   U8090 : NAND3_X1 port map( A1 => n31924, A2 => n29013, A3 => n4744, ZN => 
                           n26958);
   U8096 : XOR2_X1 port map( A1 => n2142, A2 => n17040, Z => n2143);
   U8098 : XOR2_X1 port map( A1 => n6386, A2 => n17052, Z => n17040);
   U8101 : NAND2_X2 port map( A1 => n8453, A2 => n164, ZN => n7667);
   U8133 : XOR2_X1 port map( A1 => n14136, A2 => n51, Z => n3847);
   U8140 : XOR2_X1 port map( A1 => n29545, A2 => n24699, Z => n25385);
   U8146 : OAI21_X1 port map( A1 => n13526, A2 => n18794, B => n18793, ZN => 
                           n9887);
   U8152 : NOR2_X2 port map( A1 => n1898, A2 => n29548, ZN => n1897);
   U8169 : XOR2_X1 port map( A1 => n19568, A2 => n10552, Z => n29550);
   U8173 : NAND3_X1 port map( A1 => n4916, A2 => n22651, A3 => n14253, ZN => 
                           n29551);
   U8176 : NAND2_X2 port map( A1 => n30988, A2 => n11948, ZN => n7226);
   U8184 : XOR2_X1 port map( A1 => n27226, A2 => n29554, Z => n10402);
   U8188 : XOR2_X1 port map( A1 => n1971, A2 => n1905, Z => n29554);
   U8193 : NOR2_X1 port map( A1 => n20162, A2 => n20161, ZN => n29725);
   U8194 : NOR2_X2 port map( A1 => n18666, A2 => n29555, ZN => n19308);
   U8195 : OAI22_X1 port map( A1 => n2523, A2 => n18866, B1 => n18665, B2 => 
                           n711, ZN => n29555);
   U8199 : NAND2_X2 port map( A1 => n1008, A2 => n10699, ZN => n21932);
   U8202 : AOI22_X2 port map( A1 => n5252, A2 => n1265, B1 => n4777, B2 => 
                           n26612, ZN => n4776);
   U8204 : NAND2_X2 port map( A1 => n4780, A2 => n4779, ZN => n4778);
   U8205 : NAND2_X2 port map( A1 => n29557, A2 => n17718, ZN => n30538);
   U8223 : XOR2_X1 port map( A1 => n22109, A2 => n22111, Z => n4797);
   U8231 : XOR2_X1 port map( A1 => n29559, A2 => n27243, Z => n31611);
   U8232 : XOR2_X1 port map( A1 => n23262, A2 => n25049, Z => n29559);
   U8245 : NOR2_X1 port map( A1 => n19972, A2 => n20444, ZN => n29560);
   U8250 : NAND2_X1 port map( A1 => n10132, A2 => n23821, ZN => n29561);
   U8251 : NAND2_X2 port map( A1 => n29562, A2 => n30641, ZN => n30640);
   U8263 : XOR2_X1 port map( A1 => n20769, A2 => n1340, Z => n20687);
   U8269 : NAND2_X2 port map( A1 => n29563, A2 => n22436, ZN => n8365);
   U8276 : XOR2_X1 port map( A1 => n20839, A2 => n28813, Z => n8855);
   U8277 : NAND3_X2 port map( A1 => n29899, A2 => n20500, A3 => n16759, ZN => 
                           n20839);
   U8278 : AOI22_X1 port map( A1 => n10229, A2 => n19167, B1 => n25985, B2 => 
                           n10228, ZN => n9711);
   U8284 : INV_X2 port map( I => n24339, ZN => n24163);
   U8285 : NAND3_X2 port map( A1 => n8720, A2 => n8719, A3 => n23780, ZN => 
                           n24339);
   U8323 : XOR2_X1 port map( A1 => n1044, A2 => n31138, Z => n14223);
   U8326 : XOR2_X1 port map( A1 => n29572, A2 => n1192, Z => Ciphertext(156));
   U8327 : NAND2_X2 port map( A1 => n25846, A2 => n25844, ZN => n27162);
   U8332 : NAND2_X2 port map( A1 => n25838, A2 => n7143, ZN => n25846);
   U8342 : NAND2_X1 port map( A1 => n21132, A2 => n21442, ZN => n29573);
   U8370 : XOR2_X1 port map( A1 => n4949, A2 => n30463, Z => n18048);
   U8382 : XOR2_X1 port map( A1 => n2308, A2 => n22096, Z => n22166);
   U8393 : OAI21_X1 port map( A1 => n31144, A2 => n22377, B => n31143, ZN => 
                           n13535);
   U8398 : NAND3_X2 port map( A1 => n11139, A2 => n11140, A3 => n20254, ZN => 
                           n12459);
   U8399 : AOI21_X2 port map( A1 => n25901, A2 => n25904, B => n29578, ZN => 
                           n26569);
   U8400 : NAND2_X2 port map( A1 => n28455, A2 => n25902, ZN => n29578);
   U8402 : XOR2_X1 port map( A1 => n9781, A2 => n23264, Z => n23311);
   U8424 : OAI22_X2 port map( A1 => n18917, A2 => n18916, B1 => n13200, B2 => 
                           n19119, ZN => n29581);
   U8427 : XOR2_X1 port map( A1 => n9121, A2 => n29582, Z => n9120);
   U8429 : XOR2_X1 port map( A1 => n17705, A2 => n29475, Z => n29582);
   U8440 : NOR2_X2 port map( A1 => n29586, A2 => n16070, ZN => n28802);
   U8442 : INV_X4 port map( I => n4834, ZN => n23085);
   U8446 : NAND2_X1 port map( A1 => n5673, A2 => n12593, ZN => n5672);
   U8447 : INV_X4 port map( I => n23832, ZN => n29965);
   U8450 : OAI21_X2 port map( A1 => n22448, A2 => n1297, B => n27886, ZN => 
                           n14402);
   U8455 : XOR2_X1 port map( A1 => n24492, A2 => n29588, Z => n10841);
   U8459 : XOR2_X1 port map( A1 => n28258, A2 => n12, Z => n29588);
   U8468 : NOR2_X1 port map( A1 => n11915, A2 => n8074, ZN => n29743);
   U8474 : XOR2_X1 port map( A1 => n19544, A2 => n19431, Z => n18083);
   U8477 : NAND3_X1 port map( A1 => n21316, A2 => n20330, A3 => n8115, ZN => 
                           n16048);
   U8524 : INV_X2 port map( I => n10187, ZN => n30360);
   U8526 : XOR2_X1 port map( A1 => n29600, A2 => n15415, Z => Ciphertext(17));
   U8528 : AOI22_X1 port map( A1 => n24961, A2 => n28662, B1 => n24958, B2 => 
                           n24959, ZN => n29600);
   U8532 : OAI22_X2 port map( A1 => n9842, A2 => n21335, B1 => n21337, B2 => 
                           n21336, ZN => n8140);
   U8557 : BUF_X4 port map( I => n29268, Z => n4991);
   U8566 : NOR2_X2 port map( A1 => n9900, A2 => n9899, ZN => n29606);
   U8578 : XOR2_X1 port map( A1 => n23192, A2 => n23462, Z => n29719);
   U8579 : NAND2_X2 port map( A1 => n27008, A2 => n29607, ZN => n9280);
   U8582 : OAI21_X2 port map( A1 => n28456, A2 => n28019, B => n905, ZN => 
                           n29607);
   U8590 : NAND2_X1 port map( A1 => n817, A2 => n20595, ZN => n20598);
   U8595 : AOI22_X2 port map( A1 => n1297, A2 => n15763, B1 => n22570, B2 => 
                           n18073, ZN => n29608);
   U8597 : NOR2_X2 port map( A1 => n17348, A2 => n27635, ZN => n21696);
   U8608 : XOR2_X1 port map( A1 => n4260, A2 => n8116, Z => n21224);
   U8620 : NOR3_X1 port map( A1 => n19322, A2 => n19274, A3 => n30894, ZN => 
                           n6023);
   U8622 : INV_X1 port map( I => n10075, ZN => n12419);
   U8624 : XOR2_X1 port map( A1 => n10075, A2 => n29609, Z => n22003);
   U8629 : INV_X1 port map( I => n25098, ZN => n29609);
   U8631 : NAND2_X2 port map( A1 => n6766, A2 => n6764, ZN => n10075);
   U8643 : OR2_X2 port map( A1 => n2019, A2 => n28245, Z => n10264);
   U8661 : OAI22_X2 port map( A1 => n21843, A2 => n338, B1 => n21841, B2 => 
                           n27937, ZN => n14595);
   U8674 : NAND2_X1 port map( A1 => n4259, A2 => n18767, ZN => n18377);
   U8683 : INV_X2 port map( I => n29330, ZN => n10376);
   U8684 : NAND2_X2 port map( A1 => n4709, A2 => n4706, ZN => n2600);
   U8691 : OAI21_X2 port map( A1 => n19843, A2 => n7609, B => n29615, ZN => 
                           n15169);
   U8720 : XOR2_X1 port map( A1 => n22078, A2 => n22059, Z => n22284);
   U8732 : NAND2_X2 port map( A1 => n9545, A2 => n27445, ZN => n13473);
   U8743 : XOR2_X1 port map( A1 => n29618, A2 => n19713, Z => n9760);
   U8744 : XOR2_X1 port map( A1 => n19711, A2 => n25998, Z => n29618);
   U8751 : NOR2_X1 port map( A1 => n27910, A2 => n386, ZN => n15405);
   U8764 : OR2_X1 port map( A1 => n9759, A2 => n5287, Z => n5267);
   U8772 : NAND3_X1 port map( A1 => n22670, A2 => n858, A3 => n994, ZN => 
                           n29620);
   U8779 : NAND2_X1 port map( A1 => n18089, A2 => n8100, ZN => n8783);
   U8792 : INV_X2 port map( I => n16209, ZN => n18976);
   U8830 : XOR2_X1 port map( A1 => n29828, A2 => n20671, Z => n29624);
   U8877 : XOR2_X1 port map( A1 => n24116, A2 => n25990, Z => n30774);
   U8883 : INV_X2 port map( I => n15633, ZN => n725);
   U8884 : NAND2_X2 port map( A1 => n15636, A2 => n28894, ZN => n15633);
   U8898 : OR2_X1 port map( A1 => n10899, A2 => n10900, Z => n18118);
   U8901 : INV_X2 port map( I => n11172, ZN => n29629);
   U8924 : BUF_X4 port map( I => n4646, Z => n38);
   U8930 : INV_X2 port map( I => n29631, ZN => n12974);
   U8937 : NAND2_X1 port map( A1 => n3673, A2 => n4041, ZN => n4040);
   U8938 : XOR2_X1 port map( A1 => n14385, A2 => n24602, Z => n8987);
   U8939 : NAND2_X2 port map( A1 => n8989, A2 => n8988, ZN => n24602);
   U8940 : NAND2_X2 port map( A1 => n23046, A2 => n23045, ZN => n23047);
   U8949 : XOR2_X1 port map( A1 => n24755, A2 => n12754, Z => n18001);
   U8960 : NAND2_X2 port map( A1 => n17587, A2 => n8114, ZN => n24755);
   U8984 : NAND2_X1 port map( A1 => n25736, A2 => n10285, ZN => n8555);
   U8991 : NOR2_X1 port map( A1 => n31325, A2 => n27007, ZN => n10972);
   U9014 : XOR2_X1 port map( A1 => n13716, A2 => n29633, Z => n20657);
   U9019 : XOR2_X1 port map( A1 => n27643, A2 => n26647, Z => n29633);
   U9030 : OAI22_X2 port map( A1 => n834, A2 => n1214, B1 => n32590, B2 => 
                           n33155, ZN => n1620);
   U9032 : BUF_X4 port map( I => n13646, Z => n29769);
   U9035 : NOR2_X1 port map( A1 => n22899, A2 => n31325, ZN => n27410);
   U9037 : NOR2_X1 port map( A1 => n15947, A2 => n15946, ZN => n29706);
   U9038 : INV_X2 port map( I => n14238, ZN => n18242);
   U9042 : NAND2_X2 port map( A1 => n7049, A2 => n7050, ZN => n31085);
   U9050 : XOR2_X1 port map( A1 => n15083, A2 => n29636, Z => n27766);
   U9055 : XOR2_X1 port map( A1 => n3009, A2 => n24833, Z => n29636);
   U9063 : NAND2_X1 port map( A1 => n23984, A2 => n1233, ZN => n31553);
   U9086 : XOR2_X1 port map( A1 => n29638, A2 => n15427, Z => n15425);
   U9091 : NOR2_X1 port map( A1 => n29213, A2 => n14661, ZN => n31442);
   U9092 : XOR2_X1 port map( A1 => n22237, A2 => n1716, Z => n85);
   U9094 : XOR2_X1 port map( A1 => n22294, A2 => n18189, Z => n22237);
   U9100 : XOR2_X1 port map( A1 => n4400, A2 => n11219, Z => n6720);
   U9116 : NAND2_X1 port map( A1 => n24210, A2 => n29785, ZN => n2944);
   U9117 : NAND2_X2 port map( A1 => n7261, A2 => n23582, ZN => n24210);
   U9124 : NAND2_X1 port map( A1 => n3094, A2 => n3096, ZN => n20189);
   U9125 : AND2_X2 port map( A1 => n11333, A2 => n26551, Z => n19845);
   U9129 : INV_X2 port map( I => n29642, ZN => n596);
   U9136 : NAND2_X2 port map( A1 => n31074, A2 => n8910, ZN => n8909);
   U9148 : NOR2_X2 port map( A1 => n21573, A2 => n33992, ZN => n21627);
   U9154 : XOR2_X1 port map( A1 => n12714, A2 => n29643, Z => n16886);
   U9160 : XOR2_X1 port map( A1 => n29042, A2 => n2616, Z => n20794);
   U9161 : NAND2_X2 port map( A1 => n30942, A2 => n2610, ZN => n2616);
   U9162 : NOR2_X1 port map( A1 => n28455, A2 => n11045, ZN => n1522);
   U9165 : BUF_X2 port map( I => n19668, Z => n29644);
   U9166 : AOI22_X2 port map( A1 => n30854, A2 => n11912, B1 => n5480, B2 => 
                           n6842, ZN => n9842);
   U9175 : XOR2_X1 port map( A1 => n4884, A2 => n29645, Z => n4881);
   U9178 : XOR2_X1 port map( A1 => n4883, A2 => n28859, Z => n29645);
   U9179 : XOR2_X1 port map( A1 => n29646, A2 => n5207, Z => n6039);
   U9182 : XOR2_X1 port map( A1 => n14593, A2 => n5206, Z => n29646);
   U9185 : XOR2_X1 port map( A1 => n20920, A2 => n20892, Z => n20972);
   U9193 : OAI22_X2 port map( A1 => n9435, A2 => n6675, B1 => n17202, B2 => 
                           n22861, ZN => n23519);
   U9195 : NAND2_X1 port map( A1 => n30637, A2 => n28064, ZN => n17878);
   U9202 : NAND2_X2 port map( A1 => n20188, A2 => n20190, ZN => n30637);
   U9220 : XOR2_X1 port map( A1 => n9303, A2 => n4858, Z => n20974);
   U9232 : INV_X2 port map( I => n29650, ZN => n15467);
   U9235 : XOR2_X1 port map( A1 => n27135, A2 => n1445, Z => n29650);
   U9239 : NOR2_X2 port map( A1 => n32800, A2 => n15371, ZN => n21652);
   U9241 : XOR2_X1 port map( A1 => n22269, A2 => n31913, Z => n27106);
   U9242 : XOR2_X1 port map( A1 => n21945, A2 => n26193, Z => n22269);
   U9243 : XOR2_X1 port map( A1 => n8571, A2 => n30943, Z => n31857);
   U9247 : NOR2_X1 port map( A1 => n20258, A2 => n29603, ZN => n29651);
   U9249 : XOR2_X1 port map( A1 => n6609, A2 => n29653, Z => n30905);
   U9255 : XOR2_X1 port map( A1 => n30540, A2 => n16479, Z => n23552);
   U9257 : NAND2_X2 port map( A1 => n28113, A2 => n4928, ZN => n30540);
   U9265 : INV_X2 port map( I => n21846, ZN => n29654);
   U9267 : NOR2_X1 port map( A1 => n29118, A2 => n1180, ZN => n2869);
   U9281 : XOR2_X1 port map( A1 => n19664, A2 => n29657, Z => n19901);
   U9287 : XOR2_X1 port map( A1 => n19659, A2 => n19660, Z => n29657);
   U9295 : XOR2_X1 port map( A1 => n29660, A2 => n23264, Z => n23265);
   U9301 : XOR2_X1 port map( A1 => n29661, A2 => n19305, Z => n19307);
   U9325 : AND2_X1 port map( A1 => n11333, A2 => n6693, Z => n15072);
   U9332 : NOR2_X1 port map( A1 => n29663, A2 => n29662, ZN => n26611);
   U9333 : NOR2_X1 port map( A1 => n26198, A2 => n24956, ZN => n29662);
   U9352 : INV_X2 port map( I => n29666, ZN => n19418);
   U9354 : XNOR2_X1 port map( A1 => n5487, A2 => n11591, ZN => n29666);
   U9355 : INV_X2 port map( I => n10871, ZN => n903);
   U9359 : INV_X2 port map( I => n8438, ZN => n17590);
   U9361 : XOR2_X1 port map( A1 => n10707, A2 => n27766, Z => n8438);
   U9362 : OR2_X1 port map( A1 => n20120, A2 => n16595, Z => n6223);
   U9364 : INV_X2 port map( I => n29667, ZN => n20278);
   U9375 : BUF_X4 port map( I => n20990, Z => n31584);
   U9377 : XOR2_X1 port map( A1 => n24747, A2 => n29670, Z => n31849);
   U9378 : NAND2_X2 port map( A1 => n3902, A2 => n15224, ZN => n24747);
   U9381 : NOR2_X2 port map( A1 => n4521, A2 => n4522, ZN => n12414);
   U9382 : OAI22_X2 port map( A1 => n3624, A2 => n1163, B1 => n29671, B2 => 
                           n13348, ZN => n9352);
   U9383 : AOI22_X2 port map( A1 => n12408, A2 => n822, B1 => n3626, B2 => 
                           n3790, ZN => n29671);
   U9392 : NOR2_X2 port map( A1 => n28862, A2 => n28863, ZN => n14623);
   U9397 : XOR2_X1 port map( A1 => n12330, A2 => n14518, Z => n14517);
   U9398 : INV_X2 port map( I => n29673, ZN => n12408);
   U9402 : XOR2_X1 port map( A1 => n12411, A2 => n12409, Z => n29673);
   U9408 : XOR2_X1 port map( A1 => n3109, A2 => n29675, Z => n29674);
   U9415 : NAND2_X2 port map( A1 => n26291, A2 => n29225, ZN => n31504);
   U9420 : NOR2_X2 port map( A1 => n5966, A2 => n26615, ZN => n6016);
   U9421 : AND2_X1 port map( A1 => n12471, A2 => n23085, Z => n13839);
   U9426 : NAND2_X2 port map( A1 => n31139, A2 => n34018, ZN => n5485);
   U9428 : NOR2_X2 port map( A1 => n6794, A2 => n6793, ZN => n6763);
   U9448 : INV_X4 port map( I => n29679, ZN => n8178);
   U9449 : OAI22_X2 port map( A1 => n155, A2 => n1933, B1 => n15681, B2 => 
                           n15683, ZN => n29679);
   U9451 : XOR2_X1 port map( A1 => n29680, A2 => n5421, Z => n5441);
   U9454 : XOR2_X1 port map( A1 => n22180, A2 => n2763, Z => n29680);
   U9456 : NOR2_X2 port map( A1 => n9510, A2 => n9509, ZN => n9508);
   U9462 : XOR2_X1 port map( A1 => n13606, A2 => n13457, Z => n20806);
   U9464 : AOI22_X2 port map( A1 => n12030, A2 => n8186, B1 => n11951, B2 => 
                           n1082, ZN => n29681);
   U9475 : NAND2_X1 port map( A1 => n29682, A2 => n23851, ZN => n4106);
   U9491 : AOI21_X2 port map( A1 => n12209, A2 => n29380, B => n992, ZN => 
                           n13894);
   U9507 : NAND2_X2 port map( A1 => n30966, A2 => n4268, ZN => n6169);
   U9512 : XOR2_X1 port map( A1 => n1344, A2 => n20996, Z => n20911);
   U9518 : AOI22_X2 port map( A1 => n13548, A2 => n18892, B1 => n18792, B2 => 
                           n8376, ZN => n5456);
   U9534 : XOR2_X1 port map( A1 => n12258, A2 => n29687, Z => n5500);
   U9536 : XOR2_X1 port map( A1 => n30048, A2 => n5348, Z => n12258);
   U9537 : INV_X2 port map( I => n29688, ZN => n9390);
   U9541 : XOR2_X1 port map( A1 => n7887, A2 => n29689, Z => n30600);
   U9542 : XOR2_X1 port map( A1 => n9629, A2 => n9292, Z => n2363);
   U9545 : AOI22_X2 port map( A1 => n1768, A2 => n19236, B1 => n1766, B2 => 
                           n1767, ZN => n9292);
   U9558 : NAND2_X1 port map( A1 => n21412, A2 => n11513, ZN => n21113);
   U9568 : XOR2_X1 port map( A1 => n29696, A2 => n29447, Z => n575);
   U9579 : XOR2_X1 port map( A1 => n19444, A2 => n26534, Z => n29696);
   U9606 : NAND2_X2 port map( A1 => n19928, A2 => n19929, ZN => n16606);
   U9624 : INV_X2 port map( I => n4107, ZN => n9218);
   U9628 : XOR2_X1 port map( A1 => n13644, A2 => n17837, Z => n4107);
   U9637 : NAND2_X2 port map( A1 => n4456, A2 => n28364, ZN => n23273);
   U9653 : XOR2_X1 port map( A1 => n13347, A2 => n23333, Z => n23440);
   U9661 : AOI22_X2 port map( A1 => n22574, A2 => n9959, B1 => n16503, B2 => 
                           n22926, ZN => n9647);
   U9664 : NAND2_X2 port map( A1 => n29699, A2 => n26713, ZN => n24328);
   U9674 : XOR2_X1 port map( A1 => n6229, A2 => n14817, Z => n29702);
   U9677 : OAI22_X2 port map( A1 => n16013, A2 => n21488, B1 => n16736, B2 => 
                           n16012, ZN => n22044);
   U9686 : XOR2_X1 port map( A1 => n8810, A2 => n8811, Z => n29704);
   U9705 : XOR2_X1 port map( A1 => n23242, A2 => n29707, Z => n450);
   U9707 : INV_X1 port map( I => n16598, ZN => n29707);
   U9734 : XOR2_X1 port map( A1 => n28552, A2 => n23264, Z => n29709);
   U9740 : AND2_X1 port map( A1 => n23840, A2 => n739, Z => n23493);
   U9742 : XOR2_X1 port map( A1 => n30057, A2 => n7874, Z => n31248);
   U9744 : INV_X2 port map( I => n22251, ZN => n6435);
   U9751 : NAND2_X2 port map( A1 => n29711, A2 => n21399, ZN => n21628);
   U9758 : XOR2_X1 port map( A1 => n7796, A2 => n24632, Z => n24754);
   U9761 : INV_X2 port map( I => n29712, ZN => n11805);
   U9762 : XNOR2_X1 port map( A1 => n7998, A2 => n11806, ZN => n29712);
   U9764 : XOR2_X1 port map( A1 => n33633, A2 => n16138, Z => n29989);
   U9772 : NOR2_X2 port map( A1 => n28915, A2 => n17960, ZN => n29714);
   U9779 : OAI22_X2 port map( A1 => n21343, A2 => n5141, B1 => n9073, B2 => 
                           n21341, ZN => n29717);
   U9782 : OAI21_X2 port map( A1 => n30681, A2 => n27574, B => n15032, ZN => 
                           n30410);
   U9792 : BUF_X2 port map( I => n28951, Z => n29718);
   U9803 : XOR2_X1 port map( A1 => n33492, A2 => n12454, Z => n6687);
   U9806 : NOR2_X2 port map( A1 => n31785, A2 => n15973, ZN => n27922);
   U9807 : AND2_X1 port map( A1 => n17963, A2 => n10327, Z => n1521);
   U9813 : AND2_X1 port map( A1 => n8857, A2 => n19960, Z => n29841);
   U9821 : OAI22_X2 port map( A1 => n9191, A2 => n17985, B1 => n30313, B2 => 
                           n18035, ZN => n21264);
   U9834 : XOR2_X1 port map( A1 => n29720, A2 => n12628, Z => n10475);
   U9842 : OAI22_X2 port map( A1 => n1008, A2 => n21708, B1 => n21709, B2 => 
                           n30440, ZN => n29721);
   U9852 : NAND2_X2 port map( A1 => n30688, A2 => n29722, ZN => n9107);
   U9857 : NOR2_X1 port map( A1 => n11916, A2 => n15467, ZN => n29922);
   U9867 : XOR2_X1 port map( A1 => n29723, A2 => n25071, Z => Ciphertext(43));
   U9874 : NOR2_X2 port map( A1 => n29725, A2 => n29724, ZN => n10949);
   U9876 : AND2_X1 port map( A1 => n432, A2 => n5016, Z => n5017);
   U9878 : NAND2_X2 port map( A1 => n31136, A2 => n26431, ZN => n432);
   U9894 : NAND2_X2 port map( A1 => n29727, A2 => n12379, ZN => n13346);
   U9908 : NOR2_X2 port map( A1 => n12296, A2 => n12297, ZN => n11454);
   U9914 : AOI21_X2 port map( A1 => n6864, A2 => n1826, B => n6263, ZN => 
                           n29729);
   U9915 : NAND2_X2 port map( A1 => n24152, A2 => n5317, ZN => n27259);
   U9925 : NAND2_X1 port map( A1 => n3204, A2 => n18359, ZN => n29731);
   U9926 : XOR2_X1 port map( A1 => n29732, A2 => n16507, Z => Ciphertext(22));
   U9930 : NAND2_X1 port map( A1 => n16021, A2 => n26275, ZN => n29732);
   U9933 : XOR2_X1 port map( A1 => n29733, A2 => n4004, Z => n4243);
   U9934 : XOR2_X1 port map( A1 => n30774, A2 => n5425, Z => n29733);
   U9942 : XOR2_X1 port map( A1 => n1342, A2 => n20861, Z => n6465);
   U9978 : NOR2_X2 port map( A1 => n15991, A2 => n18839, ZN => n19389);
   U9986 : NOR2_X2 port map( A1 => n729, A2 => n19853, ZN => n19854);
   U9997 : NAND3_X1 port map( A1 => n16389, A2 => n16466, A3 => n16572, ZN => 
                           n29738);
   U10023 : NAND2_X2 port map( A1 => n2360, A2 => n30140, ZN => n7256);
   U10031 : OR2_X1 port map( A1 => n11814, A2 => n12037, Z => n30227);
   U10043 : BUF_X4 port map( I => n28885, Z => n30010);
   U10045 : NAND2_X1 port map( A1 => n28736, A2 => n7554, ZN => n6816);
   U10087 : XOR2_X1 port map( A1 => n20717, A2 => n31526, Z => n20785);
   U10094 : NAND2_X1 port map( A1 => n15298, A2 => n26109, ZN => n29741);
   U10123 : NAND3_X2 port map( A1 => n2337, A2 => n8753, A3 => n396, ZN => 
                           n31051);
   U10131 : NOR2_X2 port map( A1 => n2795, A2 => n28183, ZN => n31408);
   U10151 : NAND2_X2 port map( A1 => n887, A2 => n24805, ZN => n1646);
   U10189 : NAND2_X2 port map( A1 => n29751, A2 => n16948, ZN => n18576);
   U10204 : NAND2_X2 port map( A1 => n29148, A2 => n31404, ZN => n21945);
   U10258 : AOI21_X1 port map( A1 => n1074, A2 => n27183, B => n32867, ZN => 
                           n15855);
   U10266 : NAND2_X2 port map( A1 => n22974, A2 => n22973, ZN => n7004);
   U10273 : NAND2_X1 port map( A1 => n29755, A2 => n3931, ZN => n8305);
   U10274 : NAND2_X1 port map( A1 => n12804, A2 => n8813, ZN => n29755);
   U10275 : NAND2_X2 port map( A1 => n14176, A2 => n20466, ZN => n21018);
   U10280 : INV_X2 port map( I => n16451, ZN => n753);
   U10309 : OAI21_X1 port map( A1 => n26753, A2 => n25773, B => n25788, ZN => 
                           n25777);
   U10311 : NAND2_X2 port map( A1 => n14703, A2 => n11200, ZN => n17566);
   U10320 : NAND2_X1 port map( A1 => n21165, A2 => n4755, ZN => n7063);
   U10321 : NOR2_X2 port map( A1 => n3308, A2 => n3307, ZN => n3350);
   U10333 : NAND2_X2 port map( A1 => n29934, A2 => n29759, ZN => n24094);
   U10334 : NAND3_X1 port map( A1 => n15803, A2 => n23939, A3 => n12080, ZN => 
                           n29759);
   U10343 : XOR2_X1 port map( A1 => n19439, A2 => n19440, Z => n9004);
   U10365 : XOR2_X1 port map( A1 => n8283, A2 => n9760, Z => n9759);
   U10368 : OAI21_X2 port map( A1 => n8084, A2 => n7544, B => n29761, ZN => 
                           n7357);
   U10371 : NAND2_X2 port map( A1 => n22890, A2 => n16501, ZN => n29761);
   U10374 : XOR2_X1 port map( A1 => n22157, A2 => n33437, Z => n22213);
   U10382 : XOR2_X1 port map( A1 => n24503, A2 => n29762, Z => n16510);
   U10396 : NAND2_X2 port map( A1 => n3556, A2 => n8769, ZN => n30450);
   U10397 : XOR2_X1 port map( A1 => n29765, A2 => n24833, Z => Ciphertext(6));
   U10398 : NAND4_X2 port map( A1 => n24348, A2 => n24349, A3 => n24930, A4 => 
                           n24350, ZN => n29765);
   U10401 : NAND2_X2 port map( A1 => n14579, A2 => n26793, ZN => n25796);
   U10413 : NOR2_X2 port map( A1 => n31016, A2 => n29396, ZN => n31015);
   U10415 : INV_X4 port map( I => n11904, ZN => n15682);
   U10416 : AOI21_X2 port map( A1 => n17566, A2 => n5041, B => n28945, ZN => 
                           n26874);
   U10426 : OAI21_X2 port map( A1 => n21668, A2 => n11991, B => n21674, ZN => 
                           n5996);
   U10438 : OAI21_X2 port map( A1 => n30512, A2 => n17963, B => n17894, ZN => 
                           n17475);
   U10439 : NAND2_X2 port map( A1 => n29771, A2 => n33480, ZN => n17894);
   U10446 : NOR2_X1 port map( A1 => n16194, A2 => n31379, ZN => n16195);
   U10457 : XOR2_X1 port map( A1 => Plaintext(144), A2 => Key(144), Z => n29776
                           );
   U10458 : XOR2_X1 port map( A1 => n6702, A2 => n29778, Z => n6700);
   U10459 : XOR2_X1 port map( A1 => n13644, A2 => n20801, Z => n29778);
   U10485 : NOR3_X2 port map( A1 => n2582, A2 => n4017, A3 => n1181, ZN => 
                           n16353);
   U10490 : NOR2_X1 port map( A1 => n30727, A2 => n29978, ZN => n6786);
   U10503 : NAND2_X2 port map( A1 => n21698, A2 => n21699, ZN => n3704);
   U10522 : XOR2_X1 port map( A1 => n24766, A2 => n29787, Z => n13511);
   U10523 : XOR2_X1 port map( A1 => n30290, A2 => n3294, Z => n29787);
   U10525 : XOR2_X1 port map( A1 => n24393, A2 => n12493, Z => n24829);
   U10529 : NAND3_X2 port map( A1 => n31208, A2 => n13576, A3 => n31209, ZN => 
                           n29788);
   U10531 : XOR2_X1 port map( A1 => n2489, A2 => n265, Z => n5020);
   U10551 : OR2_X1 port map( A1 => n12615, A2 => n23841, Z => n31691);
   U10552 : OAI21_X2 port map( A1 => n29791, A2 => n8990, B => n2113, ZN => 
                           n2112);
   U10557 : XOR2_X1 port map( A1 => n23230, A2 => n16073, Z => n23427);
   U10559 : NAND3_X2 port map( A1 => n7412, A2 => n26705, A3 => n22717, ZN => 
                           n23230);
   U10568 : XOR2_X1 port map( A1 => n29536, A2 => n27185, Z => n28868);
   U10572 : NAND2_X2 port map( A1 => n1544, A2 => n1543, ZN => n27185);
   U10586 : AOI21_X2 port map( A1 => n18386, A2 => n3836, B => n18385, ZN => 
                           n5118);
   U10598 : NAND2_X2 port map( A1 => n20624, A2 => n20622, ZN => n29814);
   U10599 : XOR2_X1 port map( A1 => n30997, A2 => n21958, Z => n26340);
   U10612 : AND2_X1 port map( A1 => n15394, A2 => n13969, Z => n18172);
   U10628 : XOR2_X1 port map( A1 => n29800, A2 => n23509, Z => n28870);
   U10630 : XOR2_X1 port map( A1 => n8916, A2 => n8915, Z => n29800);
   U10633 : XOR2_X1 port map( A1 => n2665, A2 => n2668, Z => n25141);
   U10638 : OR2_X1 port map( A1 => n28731, A2 => n27958, Z => n28009);
   U10642 : INV_X2 port map( I => n29803, ZN => n29270);
   U10643 : XOR2_X1 port map( A1 => n6762, A2 => n6760, Z => n29803);
   U10652 : NAND3_X2 port map( A1 => n7580, A2 => n7579, A3 => n29804, ZN => 
                           n20605);
   U10653 : OR2_X1 port map( A1 => n16243, A2 => n20109, Z => n29804);
   U10664 : NAND2_X1 port map( A1 => n28263, A2 => n8553, ZN => n26046);
   U10666 : XOR2_X1 port map( A1 => n5462, A2 => n16642, Z => n9231);
   U10670 : INV_X2 port map( I => n21356, ZN => n5395);
   U10672 : NAND2_X1 port map( A1 => n9106, A2 => n9151, ZN => n28001);
   U10673 : XOR2_X1 port map( A1 => n4465, A2 => n4464, Z => n4224);
   U10678 : XOR2_X1 port map( A1 => n6445, A2 => n29969, Z => n29807);
   U10679 : NOR2_X2 port map( A1 => n4279, A2 => n29808, ZN => n19048);
   U10681 : XOR2_X1 port map( A1 => n29809, A2 => n6185, Z => n27352);
   U10695 : XOR2_X1 port map( A1 => n20822, A2 => n20842, Z => n21000);
   U10704 : XOR2_X1 port map( A1 => n29813, A2 => n29812, Z => n9929);
   U10707 : XOR2_X1 port map( A1 => n14404, A2 => n19443, Z => n29812);
   U10709 : XOR2_X1 port map( A1 => n19538, A2 => n9928, Z => n29813);
   U10724 : NAND2_X1 port map( A1 => n17597, A2 => n17598, ZN => n9836);
   U10728 : XOR2_X1 port map( A1 => n4087, A2 => n18121, Z => n22457);
   U10753 : AND2_X1 port map( A1 => n10199, A2 => n3013, Z => n30067);
   U10754 : NAND2_X2 port map( A1 => n10970, A2 => n10971, ZN => n23200);
   U10763 : XOR2_X1 port map( A1 => n22021, A2 => n21952, Z => n21984);
   U10777 : NOR2_X2 port map( A1 => n23623, A2 => n23622, ZN => n24816);
   U10792 : NAND2_X2 port map( A1 => n29818, A2 => n29817, ZN => n7363);
   U10799 : XOR2_X1 port map( A1 => n29820, A2 => n960, Z => Ciphertext(131));
   U10801 : AOI22_X1 port map( A1 => n10959, A2 => n691, B1 => n3639, B2 => 
                           n30285, ZN => n29820);
   U10804 : AOI22_X1 port map( A1 => n15429, A2 => n27142, B1 => n13809, B2 => 
                           n15888, ZN => n29821);
   U10813 : NOR2_X2 port map( A1 => n29070, A2 => n10641, ZN => n12762);
   U10823 : OAI22_X2 port map( A1 => n10321, A2 => n29444, B1 => n10322, B2 => 
                           n10323, ZN => n10332);
   U10836 : NAND2_X1 port map( A1 => n13561, A2 => n22648, ZN => n8427);
   U10849 : XOR2_X1 port map( A1 => n26842, A2 => n29825, Z => n3536);
   U10851 : XOR2_X1 port map( A1 => n9267, A2 => n28606, Z => n29825);
   U10852 : OR2_X1 port map( A1 => n30506, A2 => n28450, Z => n14525);
   U10855 : OR2_X1 port map( A1 => n21669, A2 => n21604, Z => n29827);
   U10859 : XOR2_X1 port map( A1 => n21881, A2 => n21880, Z => n22565);
   U10880 : XOR2_X1 port map( A1 => n22264, A2 => n13612, Z => n22023);
   U10881 : NOR2_X2 port map( A1 => n30965, A2 => n13613, ZN => n22264);
   U10884 : NAND2_X2 port map( A1 => n13355, A2 => n11295, ZN => n15117);
   U10891 : INV_X2 port map( I => n29829, ZN => n11983);
   U10895 : NOR2_X2 port map( A1 => n27307, A2 => n13587, ZN => n29829);
   U10902 : AND2_X1 port map( A1 => n16249, A2 => n18510, Z => n17623);
   U10908 : AND2_X1 port map( A1 => n8758, A2 => n15318, Z => n16406);
   U10911 : NOR2_X2 port map( A1 => n25670, A2 => n27173, ZN => n14780);
   U10916 : NOR2_X1 port map( A1 => n9582, A2 => n9584, ZN => n29830);
   U10923 : INV_X2 port map( I => n8189, ZN => n29832);
   U10926 : NAND2_X2 port map( A1 => n16606, A2 => n20565, ZN => n13253);
   U10930 : NOR2_X1 port map( A1 => n10409, A2 => n23768, ZN => n29834);
   U10935 : AOI22_X2 port map( A1 => n20234, A2 => n12263, B1 => n8942, B2 => 
                           n4647, ZN => n29835);
   U10940 : NAND3_X2 port map( A1 => n3546, A2 => n3545, A3 => n29836, ZN => 
                           n7731);
   U10943 : NOR2_X2 port map( A1 => n4164, A2 => n29837, ZN => n16356);
   U10945 : OAI21_X2 port map( A1 => n15682, A2 => n23804, B => n12248, ZN => 
                           n29837);
   U10949 : XOR2_X1 port map( A1 => n23451, A2 => n23265, Z => n23270);
   U10952 : OAI21_X2 port map( A1 => n29841, A2 => n26774, B => n16154, ZN => 
                           n3293);
   U10971 : NAND2_X1 port map( A1 => n29843, A2 => n26527, ZN => n30054);
   U10978 : OAI21_X2 port map( A1 => n7245, A2 => n7244, B => n29844, ZN => 
                           n7242);
   U11000 : NOR2_X2 port map( A1 => n13525, A2 => n4916, ZN => n4918);
   U11002 : NAND2_X2 port map( A1 => n29847, A2 => n29846, ZN => n5492);
   U11005 : NAND2_X2 port map( A1 => n27294, A2 => n32106, ZN => n29847);
   U11019 : NOR2_X1 port map( A1 => n26635, A2 => n28701, ZN => n29849);
   U11022 : XOR2_X1 port map( A1 => n20693, A2 => n29851, Z => n29850);
   U11043 : OR2_X1 port map( A1 => n16781, A2 => n13905, Z => n28670);
   U11047 : NOR2_X2 port map( A1 => n4774, A2 => n12981, ZN => n24133);
   U11055 : XOR2_X1 port map( A1 => n31709, A2 => n9020, Z => n27485);
   U11059 : XOR2_X1 port map( A1 => n29855, A2 => n19440, Z => n10780);
   U11060 : XOR2_X1 port map( A1 => n34119, A2 => n11867, Z => n19440);
   U11062 : XOR2_X1 port map( A1 => n10783, A2 => n29856, Z => n29855);
   U11064 : INV_X2 port map( I => n1372, ZN => n29856);
   U11071 : NOR2_X1 port map( A1 => n10680, A2 => n29451, ZN => n8260);
   U11108 : NAND2_X1 port map( A1 => n11898, A2 => n24611, ZN => n24362);
   U11117 : INV_X2 port map( I => n5572, ZN => n30048);
   U11119 : NAND3_X2 port map( A1 => n5351, A2 => n5349, A3 => n5350, ZN => 
                           n5572);
   U11122 : OAI22_X2 port map( A1 => n10752, A2 => n8443, B1 => n6263, B2 => 
                           n6200, ZN => n16050);
   U11124 : INV_X2 port map( I => n5187, ZN => n10752);
   U11131 : XOR2_X1 port map( A1 => n9573, A2 => n9571, Z => n6458);
   U11134 : XOR2_X1 port map( A1 => n14289, A2 => n1590, Z => n29858);
   U11160 : XOR2_X1 port map( A1 => n24543, A2 => n24542, Z => n30029);
   U11168 : BUF_X2 port map( I => n28232, Z => n29864);
   U11169 : NAND2_X1 port map( A1 => n29865, A2 => n1101, ZN => n30295);
   U11170 : XOR2_X1 port map( A1 => n5278, A2 => n22877, Z => n23924);
   U11172 : AND2_X1 port map( A1 => n29296, A2 => n20569, Z => n29867);
   U11176 : NAND2_X2 port map( A1 => n7218, A2 => n2237, ZN => n14280);
   U11177 : NAND2_X2 port map( A1 => n7549, A2 => n31319, ZN => n7218);
   U11188 : INV_X2 port map( I => n16603, ZN => n23840);
   U11189 : NAND2_X1 port map( A1 => n23887, A2 => n32611, ZN => n23491);
   U11193 : BUF_X2 port map( I => n16332, Z => n29868);
   U11211 : INV_X2 port map( I => n20992, ZN => n29870);
   U11222 : XOR2_X1 port map( A1 => n4861, A2 => n4859, Z => n4862);
   U11224 : NAND2_X2 port map( A1 => n7240, A2 => n7241, ZN => n21958);
   U11226 : XOR2_X1 port map( A1 => n4894, A2 => n29873, Z => n4014);
   U11227 : XOR2_X1 port map( A1 => n7530, A2 => n1366, Z => n29873);
   U11231 : NOR2_X1 port map( A1 => n12347, A2 => n14983, ZN => n29875);
   U11245 : OAI21_X2 port map( A1 => n5553, A2 => n16532, B => n33196, ZN => 
                           n29877);
   U11255 : NOR2_X2 port map( A1 => n8337, A2 => n8164, ZN => n29878);
   U11274 : XOR2_X1 port map( A1 => n23256, A2 => n29880, Z => n5278);
   U11276 : XOR2_X1 port map( A1 => n5277, A2 => n23536, Z => n29880);
   U11280 : OAI21_X2 port map( A1 => n17289, A2 => n28638, B => n32057, ZN => 
                           n28951);
   U11281 : AND2_X1 port map( A1 => n9170, A2 => n29868, Z => n22391);
   U11296 : AND2_X1 port map( A1 => n14083, A2 => n20120, Z => n19965);
   U11302 : XNOR2_X1 port map( A1 => n20723, A2 => n506, ZN => n30265);
   U11305 : NAND2_X2 port map( A1 => n29888, A2 => n3475, ZN => n27886);
   U11306 : NAND2_X2 port map( A1 => n22446, A2 => n18073, ZN => n29888);
   U11310 : NOR2_X1 port map( A1 => n18957, A2 => n29769, ZN => n18114);
   U11311 : OAI21_X2 port map( A1 => n13949, A2 => n30648, B => n13945, ZN => 
                           n13646);
   U11341 : NOR2_X2 port map( A1 => n8270, A2 => n10955, ZN => n23638);
   U11342 : XNOR2_X1 port map( A1 => n10262, A2 => n19462, ZN => n30137);
   U11363 : AOI21_X2 port map( A1 => n20506, A2 => n17531, B => n10057, ZN => 
                           n20511);
   U11364 : AOI21_X1 port map( A1 => n20392, A2 => n9252, B => n1158, ZN => 
                           n20393);
   U11367 : XOR2_X1 port map( A1 => n29895, A2 => n9593, Z => n9592);
   U11374 : XOR2_X1 port map( A1 => n22322, A2 => n29896, Z => n29895);
   U11384 : NAND2_X1 port map( A1 => n15377, A2 => n15375, ZN => n7884);
   U11411 : AOI22_X2 port map( A1 => n7446, A2 => n33882, B1 => n7430, B2 => 
                           n12933, ZN => n26202);
   U11415 : XOR2_X1 port map( A1 => n16897, A2 => n8630, Z => n9474);
   U11418 : NOR2_X2 port map( A1 => n7144, A2 => n14864, ZN => n21700);
   U11419 : INV_X2 port map( I => n27070, ZN => n817);
   U11420 : OAI21_X2 port map( A1 => n10440, A2 => n10394, B => n19809, ZN => 
                           n27070);
   U11428 : INV_X2 port map( I => n14845, ZN => n26410);
   U11436 : NAND2_X2 port map( A1 => n24094, A2 => n18077, ZN => n5160);
   U11447 : AOI21_X2 port map( A1 => n7238, A2 => n27842, B => n29900, ZN => 
                           n21390);
   U11449 : INV_X1 port map( I => n21220, ZN => n29901);
   U11454 : NAND2_X2 port map( A1 => n31021, A2 => n2770, ZN => n3009);
   U11457 : BUF_X2 port map( I => n21248, Z => n29903);
   U11470 : OAI21_X2 port map( A1 => n13840, A2 => n13841, B => n17608, ZN => 
                           n29904);
   U11488 : XOR2_X1 port map( A1 => n15862, A2 => n15860, Z => n25394);
   U11489 : XOR2_X1 port map( A1 => n22294, A2 => n28162, Z => n22322);
   U11503 : XOR2_X1 port map( A1 => n29907, A2 => n10877, Z => n26971);
   U11506 : XOR2_X1 port map( A1 => n20838, A2 => n27014, Z => n29907);
   U11511 : AND2_X1 port map( A1 => n7901, A2 => n10868, Z => n29089);
   U11519 : NAND2_X2 port map( A1 => n29909, A2 => n18524, ZN => n19143);
   U11521 : OAI21_X2 port map( A1 => n18521, A2 => n18522, B => n18849, ZN => 
                           n29909);
   U11530 : NAND2_X2 port map( A1 => n31356, A2 => n18926, ZN => n18928);
   U11547 : XOR2_X1 port map( A1 => n4219, A2 => n11481, Z => n22250);
   U11553 : XOR2_X1 port map( A1 => n10923, A2 => n24524, Z => n29912);
   U11554 : INV_X2 port map( I => n29913, ZN => n19177);
   U11556 : NAND2_X2 port map( A1 => n29769, A2 => n19120, ZN => n29913);
   U11562 : INV_X4 port map( I => n29914, ZN => n5781);
   U11563 : INV_X4 port map( I => n14248, ZN => n31012);
   U11581 : INV_X2 port map( I => n26677, ZN => n4337);
   U11586 : NAND2_X1 port map( A1 => n30025, A2 => n14062, ZN => n84);
   U11595 : XOR2_X1 port map( A1 => n31005, A2 => n26125, Z => n16939);
   U11596 : XOR2_X1 port map( A1 => n12801, A2 => n29442, Z => n30229);
   U11597 : XOR2_X1 port map( A1 => n19473, A2 => n27781, Z => n12801);
   U11598 : NAND2_X2 port map( A1 => n29915, A2 => n8013, ZN => n19749);
   U11599 : NAND2_X2 port map( A1 => n28883, A2 => n30412, ZN => n29915);
   U11602 : INV_X2 port map( I => n29916, ZN => n28087);
   U11611 : INV_X2 port map( I => n29919, ZN => n29278);
   U11637 : NAND2_X2 port map( A1 => n9113, A2 => n29921, ZN => n2180);
   U11642 : NAND2_X1 port map( A1 => n9110, A2 => n9111, ZN => n29921);
   U11646 : XOR2_X1 port map( A1 => n24593, A2 => n24644, Z => n9121);
   U11651 : AND2_X1 port map( A1 => n4274, A2 => n28737, Z => n9817);
   U11661 : INV_X4 port map( I => n28087, ZN => n20100);
   U11663 : XOR2_X1 port map( A1 => n30321, A2 => n23247, Z => n23478);
   U11668 : INV_X2 port map( I => n7935, ZN => n24156);
   U11708 : XOR2_X1 port map( A1 => n24369, A2 => n29930, Z => n24447);
   U11709 : XOR2_X1 port map( A1 => n24687, A2 => n28918, Z => n29930);
   U11714 : AOI22_X1 port map( A1 => n12077, A2 => n1362, B1 => n14210, B2 => 
                           n10286, ZN => n3946);
   U11720 : OAI21_X2 port map( A1 => n29932, A2 => n29931, B => n21811, ZN => 
                           n16477);
   U11721 : NOR2_X2 port map( A1 => n1132, A2 => n15772, ZN => n29932);
   U11722 : NAND2_X1 port map( A1 => n33474, A2 => n12358, ZN => n17169);
   U11723 : NAND3_X2 port map( A1 => n24011, A2 => n12143, A3 => n24012, ZN => 
                           n15988);
   U11732 : NAND3_X1 port map( A1 => n5901, A2 => n964, A3 => n314, ZN => 
                           n24997);
   U11756 : XOR2_X1 port map( A1 => n6731, A2 => n13951, Z => n30093);
   U11758 : NOR2_X2 port map( A1 => n5161, A2 => n5389, ZN => n24622);
   U11762 : OAI21_X2 port map( A1 => n33745, A2 => n179, B => n7690, ZN => 
                           n29933);
   U11763 : XOR2_X1 port map( A1 => n23387, A2 => n23333, Z => n23504);
   U11765 : OAI21_X2 port map( A1 => n22888, A2 => n22889, B => n1561, ZN => 
                           n23333);
   U11767 : AND2_X1 port map( A1 => n30763, A2 => n28471, Z => n3443);
   U11777 : OAI21_X2 port map( A1 => n29937, A2 => n5730, B => n5758, ZN => 
                           n14849);
   U11781 : BUF_X2 port map( I => n20519, Z => n29938);
   U11784 : INV_X1 port map( I => n1357, ZN => n30971);
   U11786 : NAND2_X1 port map( A1 => n21664, A2 => n8323, ZN => n3016);
   U11792 : AND2_X1 port map( A1 => n13896, A2 => n27143, Z => n29002);
   U11826 : NAND2_X1 port map( A1 => n32081, A2 => n14676, ZN => n22402);
   U11835 : XOR2_X1 port map( A1 => n2073, A2 => n2075, Z => n2072);
   U11849 : AOI21_X2 port map( A1 => n14705, A2 => n14706, B => n18743, ZN => 
                           n18435);
   U11850 : AND2_X1 port map( A1 => n3486, A2 => n20155, Z => n3529);
   U11851 : XOR2_X1 port map( A1 => n14132, A2 => n20813, Z => n6081);
   U11852 : NOR2_X2 port map( A1 => n9418, A2 => n10715, ZN => n14132);
   U11862 : OAI22_X2 port map( A1 => n890, A2 => n24325, B1 => n29141, B2 => 
                           n24327, ZN => n23982);
   U11865 : NAND2_X1 port map( A1 => n15907, A2 => n7460, ZN => n30036);
   U11869 : NOR2_X2 port map( A1 => n20951, A2 => n29946, ZN => n21876);
   U11871 : OAI22_X2 port map( A1 => n20947, A2 => n13194, B1 => n21313, B2 => 
                           n20949, ZN => n29946);
   U11883 : OAI21_X2 port map( A1 => n12276, A2 => n2741, B => n12277, ZN => 
                           n30628);
   U11900 : XOR2_X1 port map( A1 => n10598, A2 => n29951, Z => n26933);
   U11908 : OR3_X2 port map( A1 => n27134, A2 => n24970, A3 => n3843, Z => n699
                           );
   U11914 : INV_X4 port map( I => n29952, ZN => n6985);
   U11925 : XOR2_X1 port map( A1 => n22246, A2 => n29953, Z => n26214);
   U11929 : XOR2_X1 port map( A1 => n21923, A2 => n29954, Z => n29953);
   U11936 : INV_X1 port map( I => n25091, ZN => n29954);
   U11944 : XOR2_X1 port map( A1 => n13477, A2 => n2818, Z => n29955);
   U11951 : NOR2_X2 port map( A1 => n33675, A2 => n4208, ZN => n22886);
   U11966 : XNOR2_X1 port map( A1 => n14120, A2 => n19580, ZN => n19406);
   U11970 : NAND2_X2 port map( A1 => n6602, A2 => n6603, ZN => n19580);
   U11973 : AND2_X1 port map( A1 => n3147, A2 => n3077, Z => n10938);
   U11978 : AND2_X1 port map( A1 => n9285, A2 => n28203, Z => n9286);
   U11979 : NAND2_X2 port map( A1 => n7312, A2 => n10339, ZN => n9285);
   U11990 : INV_X2 port map( I => n9313, ZN => n2491);
   U11991 : NAND2_X2 port map( A1 => n21125, A2 => n21678, ZN => n9313);
   U11999 : INV_X2 port map( I => n29960, ZN => n26114);
   U12001 : XOR2_X1 port map( A1 => n13235, A2 => n13234, Z => n29960);
   U12005 : AOI21_X2 port map( A1 => n13109, A2 => n32459, B => n33544, ZN => 
                           n5389);
   U12032 : XOR2_X1 port map( A1 => n12310, A2 => n29970, Z => n29969);
   U12033 : NAND3_X2 port map( A1 => n11991, A2 => n21673, A3 => n918, ZN => 
                           n5995);
   U12041 : INV_X2 port map( I => n25859, ZN => n10897);
   U12047 : NAND2_X2 port map( A1 => n13051, A2 => n13053, ZN => n25859);
   U12051 : XOR2_X1 port map( A1 => n10535, A2 => n16690, Z => n23122);
   U12052 : NAND2_X2 port map( A1 => n1471, A2 => n4936, ZN => n10535);
   U12053 : INV_X2 port map( I => n4378, ZN => n9578);
   U12055 : AND2_X1 port map( A1 => n19104, A2 => n18923, Z => n27616);
   U12056 : XOR2_X1 port map( A1 => n27352, A2 => n24470, Z => n24471);
   U12065 : AOI22_X2 port map( A1 => n8086, A2 => n8165, B1 => n13268, B2 => 
                           n24213, ZN => n31086);
   U12082 : INV_X2 port map( I => n32747, ZN => n29972);
   U12099 : NAND2_X2 port map( A1 => n30088, A2 => n11919, ZN => n14498);
   U12108 : OAI21_X2 port map( A1 => n26067, A2 => n13210, B => n29973, ZN => 
                           n13001);
   U12109 : NAND2_X2 port map( A1 => n13210, A2 => n12708, ZN => n29973);
   U12113 : NAND2_X1 port map( A1 => n4378, A2 => n9064, ZN => n26333);
   U12154 : NAND2_X2 port map( A1 => n349, A2 => n26971, ZN => n21219);
   U12164 : AND2_X1 port map( A1 => n1299, A2 => n16647, Z => n15449);
   U12176 : NAND2_X2 port map( A1 => n29975, A2 => n31612, ZN => n21860);
   U12187 : NOR2_X1 port map( A1 => n9133, A2 => n8632, ZN => n29978);
   U12216 : XOR2_X1 port map( A1 => n22249, A2 => n22160, Z => n2349);
   U12221 : OAI22_X2 port map( A1 => n2352, A2 => n21861, B1 => n2351, B2 => 
                           n3756, ZN => n22160);
   U12228 : NAND2_X2 port map( A1 => n6099, A2 => n1109, ZN => n26937);
   U12256 : XOR2_X1 port map( A1 => n13305, A2 => n471, Z => n11507);
   U12279 : XOR2_X1 port map( A1 => n22114, A2 => n22096, Z => n22171);
   U12288 : NAND3_X2 port map( A1 => n27569, A2 => n18147, A3 => n27764, ZN => 
                           n4289);
   U12292 : NAND2_X1 port map( A1 => n19035, A2 => n13796, ZN => n26817);
   U12296 : NAND2_X2 port map( A1 => n6170, A2 => n6172, ZN => n13796);
   U12299 : XOR2_X1 port map( A1 => n31373, A2 => n16128, Z => n24528);
   U12334 : XOR2_X1 port map( A1 => n29986, A2 => n19752, Z => n3967);
   U12336 : INV_X2 port map( I => n29987, ZN => n4677);
   U12340 : XOR2_X1 port map( A1 => Plaintext(53), A2 => Key(53), Z => n29987);
   U12341 : NAND2_X1 port map( A1 => n31799, A2 => n26818, ZN => n18322);
   U12344 : XOR2_X1 port map( A1 => n34082, A2 => n19644, Z => n29988);
   U12357 : XOR2_X1 port map( A1 => n29989, A2 => n19669, Z => n19671);
   U12361 : XOR2_X1 port map( A1 => n27395, A2 => n19783, Z => n19505);
   U12365 : OAI21_X2 port map( A1 => n17242, A2 => n32618, B => n17241, ZN => 
                           n16452);
   U12366 : NAND2_X1 port map( A1 => n30656, A2 => n10173, ZN => n25604);
   U12370 : XOR2_X1 port map( A1 => n5429, A2 => n24519, Z => n678);
   U12391 : OR2_X1 port map( A1 => n31360, A2 => n13483, Z => n8805);
   U12393 : XNOR2_X1 port map( A1 => n8785, A2 => n1410, ZN => n31749);
   U12403 : AOI21_X1 port map( A1 => n16648, A2 => n11820, B => n26912, ZN => 
                           n30568);
   U12413 : AOI22_X2 port map( A1 => n19940, A2 => n13994, B1 => n19941, B2 => 
                           n16637, ZN => n26278);
   U12415 : XOR2_X1 port map( A1 => n17552, A2 => n11661, Z => n11660);
   U12431 : XOR2_X1 port map( A1 => n5324, A2 => n16852, Z => n27192);
   U12432 : NAND2_X1 port map( A1 => n20013, A2 => n31046, ZN => n16261);
   U12442 : XOR2_X1 port map( A1 => n2608, A2 => n2607, Z => n20098);
   U12443 : OAI21_X2 port map( A1 => n30004, A2 => n30003, B => n1030, ZN => 
                           n11617);
   U12447 : XOR2_X1 port map( A1 => n19483, A2 => n19599, Z => n19681);
   U12452 : OAI21_X2 port map( A1 => n18391, A2 => n18390, B => n18389, ZN => 
                           n19101);
   U12454 : XOR2_X1 port map( A1 => n26623, A2 => n30007, Z => n7572);
   U12458 : NAND2_X2 port map( A1 => n11336, A2 => n11489, ZN => n26623);
   U12463 : NAND2_X2 port map( A1 => n26543, A2 => n10850, ZN => n10847);
   U12469 : XOR2_X1 port map( A1 => n3030, A2 => n22274, Z => n2477);
   U12478 : AND2_X1 port map( A1 => n22364, A2 => n22588, Z => n30507);
   U12479 : OAI21_X2 port map( A1 => n26015, A2 => n25303, B => n18059, ZN => 
                           n11111);
   U12480 : XOR2_X1 port map( A1 => n13743, A2 => n30011, Z => n17886);
   U12483 : XOR2_X1 port map( A1 => n13741, A2 => n13742, Z => n30011);
   U12484 : AOI22_X1 port map( A1 => n2130, A2 => n28849, B1 => n22981, B2 => 
                           n1280, ZN => n17893);
   U12485 : XOR2_X1 port map( A1 => n32623, A2 => n25881, Z => n17753);
   U12489 : OR2_X1 port map( A1 => n23777, A2 => n23778, Z => n8720);
   U12501 : NAND2_X1 port map( A1 => n16725, A2 => n1048, ZN => n30012);
   U12506 : NOR2_X1 port map( A1 => n5657, A2 => n26317, ZN => n6232);
   U12509 : BUF_X2 port map( I => n8919, Z => n30014);
   U12512 : INV_X2 port map( I => n5003, ZN => n7394);
   U12515 : AND2_X1 port map( A1 => n19422, A2 => n12704, Z => n30015);
   U12520 : AOI22_X2 port map( A1 => n21091, A2 => n21687, B1 => n29286, B2 => 
                           n26513, ZN => n29148);
   U12525 : XOR2_X1 port map( A1 => n31088, A2 => n29009, Z => n31087);
   U12527 : BUF_X4 port map( I => n25700, Z => n146);
   U12538 : XOR2_X1 port map( A1 => n27976, A2 => n30016, Z => n14456);
   U12551 : OR2_X1 port map( A1 => n22332, A2 => n468, Z => n13369);
   U12556 : XOR2_X1 port map( A1 => n20792, A2 => n30018, Z => n20449);
   U12566 : INV_X2 port map( I => n30020, ZN => n10465);
   U12568 : XOR2_X1 port map( A1 => n16324, A2 => n10466, Z => n30020);
   U12577 : NAND2_X2 port map( A1 => n31793, A2 => n30021, ZN => n6595);
   U12579 : OAI22_X2 port map( A1 => n30522, A2 => n30983, B1 => n765, B2 => 
                           n16783, ZN => n30021);
   U12583 : OAI21_X2 port map( A1 => n18618, A2 => n10080, B => n10964, ZN => 
                           n10977);
   U12591 : NOR2_X2 port map( A1 => n9403, A2 => n20472, ZN => n31532);
   U12600 : OAI22_X1 port map( A1 => n25464, A2 => n25467, B1 => n25463, B2 => 
                           n25473, ZN => n28302);
   U12602 : NAND2_X2 port map( A1 => n19056, A2 => n6022, ZN => n2075);
   U12627 : OAI21_X2 port map( A1 => n26047, A2 => n28495, B => n852, ZN => 
                           n9244);
   U12640 : NAND2_X1 port map( A1 => n25715, A2 => n25714, ZN => n14352);
   U12651 : XOR2_X1 port map( A1 => n23516, A2 => n16382, Z => n16259);
   U12654 : INV_X2 port map( I => n30032, ZN => n26049);
   U12655 : XOR2_X1 port map( A1 => Plaintext(188), A2 => Key(188), Z => n30032
                           );
   U12656 : AND2_X1 port map( A1 => n17298, A2 => n17514, Z => n30222);
   U12660 : NAND2_X2 port map( A1 => n12977, A2 => n12975, ZN => n19049);
   U12670 : NAND3_X2 port map( A1 => n30036, A2 => n30072, A3 => n9381, ZN => 
                           n27105);
   U12702 : NAND2_X2 port map( A1 => n26742, A2 => n12533, ZN => n30039);
   U12709 : NAND2_X1 port map( A1 => n20464, A2 => n30728, ZN => n20466);
   U12713 : INV_X2 port map( I => n21860, ZN => n5628);
   U12719 : INV_X2 port map( I => n30042, ZN => n15623);
   U12735 : OAI22_X2 port map( A1 => n27318, A2 => n8107, B1 => n8108, B2 => 
                           n18089, ZN => n20188);
   U12736 : XOR2_X1 port map( A1 => Plaintext(43), A2 => Key(43), Z => n16585);
   U12744 : XNOR2_X1 port map( A1 => n14819, A2 => n23419, ZN => n30317);
   U12753 : OAI21_X2 port map( A1 => n7429, A2 => n22342, B => n26173, ZN => 
                           n30044);
   U12761 : NAND2_X1 port map( A1 => n20411, A2 => n29356, ZN => n20047);
   U12766 : INV_X2 port map( I => n21049, ZN => n30045);
   U12774 : OAI21_X2 port map( A1 => n11444, A2 => n11280, B => n11474, ZN => 
                           n19312);
   U12784 : OAI21_X2 port map( A1 => n3092, A2 => n3091, B => n31226, ZN => 
                           n6022);
   U12785 : NAND2_X1 port map( A1 => n28913, A2 => n26594, ZN => n30192);
   U12792 : NAND2_X1 port map( A1 => n13905, A2 => n6662, ZN => n28672);
   U12793 : XOR2_X1 port map( A1 => n13817, A2 => n9373, Z => n30049);
   U12797 : NAND2_X2 port map( A1 => n12563, A2 => n13693, ZN => n20328);
   U12799 : OR2_X1 port map( A1 => n29629, A2 => n29334, Z => n4968);
   U12801 : OAI21_X2 port map( A1 => n11633, A2 => n12332, B => n30054, ZN => 
                           n17697);
   U12805 : NOR2_X1 port map( A1 => n32055, A2 => n4378, ZN => n4054);
   U12809 : NAND2_X2 port map( A1 => n12542, A2 => n28155, ZN => n22078);
   U12815 : INV_X2 port map( I => n24996, ZN => n713);
   U12819 : INV_X1 port map( I => n19571, ZN => n30058);
   U12820 : NAND3_X2 port map( A1 => n10369, A2 => n20051, A3 => n11216, ZN => 
                           n21047);
   U12831 : BUF_X2 port map( I => n23579, Z => n30059);
   U12834 : OAI21_X2 port map( A1 => n29375, A2 => n30060, B => n8835, ZN => 
                           n3166);
   U12846 : NAND2_X2 port map( A1 => n30062, A2 => n7199, ZN => n19661);
   U12850 : OAI21_X2 port map( A1 => n16463, A2 => n13619, B => n13618, ZN => 
                           n23171);
   U12851 : XOR2_X1 port map( A1 => n30063, A2 => n16691, Z => Ciphertext(34));
   U12856 : INV_X2 port map( I => n10303, ZN => n22551);
   U12867 : NAND2_X2 port map( A1 => n24187, A2 => n24188, ZN => n15536);
   U12871 : OAI21_X2 port map( A1 => n12326, A2 => n14529, B => n798, ZN => 
                           n24187);
   U12880 : XOR2_X1 port map( A1 => n22269, A2 => n8061, Z => n8060);
   U12888 : XOR2_X1 port map( A1 => n19741, A2 => n19708, Z => n17010);
   U12896 : BUF_X2 port map( I => n6407, Z => n252);
   U12909 : NAND2_X2 port map( A1 => n5627, A2 => n34008, ZN => n23896);
   U12944 : XOR2_X1 port map( A1 => n30074, A2 => n26436, Z => n8373);
   U12952 : INV_X2 port map( I => n30076, ZN => n15719);
   U12958 : XOR2_X1 port map( A1 => n17570, A2 => n17572, Z => n30076);
   U12962 : XOR2_X1 port map( A1 => n23355, A2 => n23395, Z => n11324);
   U12971 : XOR2_X1 port map( A1 => n1044, A2 => n19780, Z => n19495);
   U12983 : INV_X2 port map( I => n30078, ZN => n11521);
   U12984 : XOR2_X1 port map( A1 => n11522, A2 => n11524, Z => n30078);
   U12989 : AOI21_X2 port map( A1 => n14500, A2 => n32054, B => n26768, ZN => 
                           n17369);
   U13012 : NAND2_X2 port map( A1 => n388, A2 => n387, ZN => n25473);
   U13014 : NAND2_X2 port map( A1 => n30080, A2 => n10329, ZN => n4732);
   U13015 : XOR2_X1 port map( A1 => n8762, A2 => n16497, Z => n30596);
   U13016 : NAND2_X2 port map( A1 => n7584, A2 => n30142, ZN => n8762);
   U13024 : NAND2_X2 port map( A1 => n21207, A2 => n30081, ZN => n14691);
   U13033 : NAND2_X2 port map( A1 => n30082, A2 => n9496, ZN => n25723);
   U13041 : NAND3_X2 port map( A1 => n27359, A2 => n25702, A3 => n27127, ZN => 
                           n30082);
   U13049 : NAND2_X2 port map( A1 => n10281, A2 => n24014, ZN => n11883);
   U13052 : XOR2_X1 port map( A1 => n13511, A2 => n13513, Z => n13567);
   U13055 : NAND2_X2 port map( A1 => n4734, A2 => n23065, ZN => n10644);
   U13067 : OAI22_X2 port map( A1 => n2152, A2 => n26918, B1 => n10472, B2 => 
                           n19152, ZN => n19644);
   U13070 : XOR2_X1 port map( A1 => n2330, A2 => n17213, Z => n11434);
   U13071 : XOR2_X1 port map( A1 => n2331, A2 => n1916, Z => n2330);
   U13075 : XOR2_X1 port map( A1 => n19493, A2 => n14223, Z => n14222);
   U13078 : XOR2_X1 port map( A1 => n19632, A2 => n33749, Z => n19493);
   U13083 : XOR2_X1 port map( A1 => n982, A2 => n5211, Z => n23402);
   U13084 : OR2_X1 port map( A1 => n23755, A2 => n6705, Z => n15400);
   U13088 : XOR2_X1 port map( A1 => n3932, A2 => n30188, Z => n29213);
   U13090 : XOR2_X1 port map( A1 => n30912, A2 => n3777, Z => n5097);
   U13096 : AOI22_X2 port map( A1 => n10627, A2 => n24237, B1 => n24131, B2 => 
                           n24130, ZN => n30084);
   U13100 : OAI22_X2 port map( A1 => n3866, A2 => n3867, B1 => n6568, B2 => 
                           n10096, ZN => n25975);
   U13120 : NOR2_X1 port map( A1 => n20630, A2 => n31471, ZN => n20383);
   U13121 : OAI22_X2 port map( A1 => n4230, A2 => n32618, B1 => n10695, B2 => 
                           n9139, ZN => n31471);
   U13125 : NAND2_X2 port map( A1 => n6580, A2 => n28459, ZN => n5879);
   U13135 : INV_X4 port map( I => n16453, ZN => n14233);
   U13138 : NOR2_X2 port map( A1 => n32935, A2 => n29329, ZN => n22840);
   U13139 : NAND2_X1 port map( A1 => n30085, A2 => n11465, ZN => n11464);
   U13142 : OAI21_X1 port map( A1 => n5911, A2 => n4261, B => n28812, ZN => 
                           n30085);
   U13144 : INV_X2 port map( I => n30086, ZN => n17316);
   U13145 : XNOR2_X1 port map( A1 => Plaintext(86), A2 => Key(86), ZN => n30086
                           );
   U13147 : XOR2_X1 port map( A1 => n13645, A2 => n28889, Z => n30679);
   U13152 : AOI22_X2 port map( A1 => n15716, A2 => n21496, B1 => n21601, B2 => 
                           n25975, ZN => n21602);
   U13159 : XOR2_X1 port map( A1 => n6462, A2 => n30087, Z => n31660);
   U13172 : AOI22_X2 port map( A1 => n5852, A2 => n4550, B1 => n14117, B2 => 
                           n18493, ZN => n30088);
   U13178 : AOI21_X1 port map( A1 => n14498, A2 => n18988, B => n19089, ZN => 
                           n18900);
   U13185 : XOR2_X1 port map( A1 => n22195, A2 => n17244, Z => n14301);
   U13188 : XOR2_X1 port map( A1 => n22255, A2 => n22014, Z => n22195);
   U13191 : NAND2_X2 port map( A1 => n30090, A2 => n31814, ZN => n3157);
   U13201 : INV_X2 port map( I => n29328, ZN => n1280);
   U13203 : OAI22_X1 port map( A1 => n12551, A2 => n12520, B1 => n3222, B2 => 
                           n24249, ZN => n8204);
   U13205 : INV_X2 port map( I => n24250, ZN => n3222);
   U13217 : NOR2_X1 port map( A1 => n28183, A2 => n33848, ZN => n16159);
   U13221 : XOR2_X1 port map( A1 => n11251, A2 => n30093, Z => n31128);
   U13222 : INV_X2 port map( I => n30094, ZN => n15559);
   U13223 : XOR2_X1 port map( A1 => n16178, A2 => n20691, Z => n3010);
   U13227 : XOR2_X1 port map( A1 => n20802, A2 => n20690, Z => n16178);
   U13229 : NAND2_X2 port map( A1 => n9460, A2 => n22774, ZN => n22778);
   U13232 : OAI22_X2 port map( A1 => n19078, A2 => n19283, B1 => n28721, B2 => 
                           n31254, ZN => n28638);
   U13245 : AOI21_X2 port map( A1 => n27023, A2 => n16327, B => n27560, ZN => 
                           n16796);
   U13246 : NOR3_X2 port map( A1 => n3214, A2 => n30096, A3 => n24108, ZN => 
                           n3504);
   U13249 : NAND2_X1 port map( A1 => n4069, A2 => n29305, ZN => n12568);
   U13253 : XOR2_X1 port map( A1 => n20820, A2 => n20851, Z => n20966);
   U13255 : XOR2_X1 port map( A1 => n12610, A2 => n6974, Z => n19343);
   U13256 : NOR2_X2 port map( A1 => n30097, A2 => n2930, ZN => n2929);
   U13257 : NOR2_X2 port map( A1 => n13585, A2 => n20084, ZN => n30097);
   U13261 : NAND2_X2 port map( A1 => n12640, A2 => n12641, ZN => n13872);
   U13263 : XOR2_X1 port map( A1 => n22016, A2 => n10963, Z => n30098);
   U13265 : XOR2_X1 port map( A1 => n9468, A2 => n12800, Z => n6688);
   U13272 : XOR2_X1 port map( A1 => n12675, A2 => n25560, Z => n6103);
   U13273 : OAI21_X2 port map( A1 => n6105, A2 => n6106, B => n6104, ZN => 
                           n12675);
   U13280 : XOR2_X1 port map( A1 => n10150, A2 => n27866, Z => n10291);
   U13292 : XOR2_X1 port map( A1 => n30137, A2 => n30102, Z => n568);
   U13294 : XOR2_X1 port map( A1 => n19476, A2 => n7741, Z => n30102);
   U13297 : OAI21_X2 port map( A1 => n29976, A2 => n16752, B => n25143, ZN => 
                           n25168);
   U13304 : NOR2_X2 port map( A1 => n8760, A2 => n23721, ZN => n23722);
   U13308 : XOR2_X1 port map( A1 => n28730, A2 => n2825, Z => n2824);
   U13313 : XOR2_X1 port map( A1 => n30107, A2 => n5166, Z => n12584);
   U13320 : NAND2_X1 port map( A1 => n7515, A2 => n25214, ZN => n15339);
   U13322 : XOR2_X1 port map( A1 => n19579, A2 => n30109, Z => n7939);
   U13326 : XOR2_X1 port map( A1 => n19737, A2 => n1367, Z => n30109);
   U13331 : XOR2_X1 port map( A1 => n24399, A2 => n29348, Z => n13358);
   U13334 : NAND2_X2 port map( A1 => n30110, A2 => n24319, ZN => n14789);
   U13349 : XOR2_X1 port map( A1 => n22066, A2 => n21986, Z => n61);
   U13353 : XOR2_X1 port map( A1 => n22157, A2 => n22225, Z => n22066);
   U13357 : XOR2_X1 port map( A1 => n11660, A2 => n30111, Z => n12467);
   U13360 : XOR2_X1 port map( A1 => n19444, A2 => n11663, Z => n30111);
   U13368 : NAND2_X1 port map( A1 => n14016, A2 => n5820, ZN => n30888);
   U13372 : XOR2_X1 port map( A1 => n13436, A2 => n30644, Z => n637);
   U13378 : NOR3_X2 port map( A1 => n7857, A2 => n26667, A3 => n26739, ZN => 
                           n30578);
   U13386 : NAND3_X2 port map( A1 => n7488, A2 => n14024, A3 => n30112, ZN => 
                           n14600);
   U13391 : OAI21_X1 port map( A1 => n18843, A2 => n5700, B => n4927, ZN => 
                           n4507);
   U13392 : NAND2_X2 port map( A1 => n30115, A2 => n30114, ZN => n13579);
   U13393 : INV_X2 port map( I => n24110, ZN => n889);
   U13405 : BUF_X2 port map( I => n469, Z => n30116);
   U13427 : AND2_X1 port map( A1 => n7320, A2 => n414, Z => n2705);
   U13429 : AND2_X1 port map( A1 => n25480, A2 => n25482, Z => n30117);
   U13435 : NAND2_X1 port map( A1 => n3181, A2 => n29043, ZN => n27934);
   U13472 : NAND2_X2 port map( A1 => n30122, A2 => n26568, ZN => n4208);
   U13497 : NOR2_X2 port map( A1 => n25229, A2 => n18059, ZN => n11409);
   U13500 : AOI21_X1 port map( A1 => n9832, A2 => n9833, B => n8087, ZN => 
                           n30236);
   U13501 : OAI22_X2 port map( A1 => n18784, A2 => n34141, B1 => n6777, B2 => 
                           n18785, ZN => n13963);
   U13503 : NAND2_X2 port map( A1 => n8395, A2 => n13254, ZN => n18784);
   U13523 : INV_X2 port map( I => n30125, ZN => n11516);
   U13528 : XOR2_X1 port map( A1 => n30127, A2 => n8920, Z => n30126);
   U13537 : BUF_X2 port map( I => n21816, Z => n30129);
   U13551 : NAND2_X2 port map( A1 => n8378, A2 => n21430, ZN => n11299);
   U13555 : OR2_X1 port map( A1 => n11516, A2 => n29139, Z => n23859);
   U13568 : XOR2_X1 port map( A1 => n6904, A2 => n30135, Z => n6886);
   U13570 : XOR2_X1 port map( A1 => n22138, A2 => n30906, Z => n30135);
   U13572 : XOR2_X1 port map( A1 => n30136, A2 => n14885, Z => Ciphertext(109))
                           ;
   U13573 : AOI22_X1 port map( A1 => n25492, A2 => n25464, B1 => n25460, B2 => 
                           n25459, ZN => n30136);
   U13586 : NAND2_X2 port map( A1 => n13001, A2 => n13002, ZN => n14337);
   U13591 : INV_X2 port map( I => n25557, ZN => n15134);
   U13599 : XOR2_X1 port map( A1 => n21003, A2 => n21038, Z => n6895);
   U13600 : NAND2_X2 port map( A1 => n12365, A2 => n12364, ZN => n21038);
   U13603 : OR2_X1 port map( A1 => n4054, A2 => n9580, Z => n8199);
   U13614 : NAND3_X2 port map( A1 => n24166, A2 => n31416, A3 => n24165, ZN => 
                           n28830);
   U13615 : AOI22_X2 port map( A1 => n25657, A2 => n25664, B1 => n7083, B2 => 
                           n25666, ZN => n25668);
   U13616 : INV_X2 port map( I => n20344, ZN => n30139);
   U13622 : XNOR2_X1 port map( A1 => n24638, A2 => n25208, ZN => n30607);
   U13628 : XOR2_X1 port map( A1 => n28762, A2 => n17898, Z => n22004);
   U13630 : NAND2_X1 port map( A1 => n6841, A2 => n6840, ZN => n30140);
   U13635 : NOR2_X2 port map( A1 => n28361, A2 => n18994, ZN => n19058);
   U13636 : NAND2_X2 port map( A1 => n31856, A2 => n94, ZN => n18994);
   U13649 : XOR2_X1 port map( A1 => n24540, A2 => n9681, Z => n2210);
   U13653 : AOI21_X2 port map( A1 => n782, A2 => n20535, B => n31250, ZN => 
                           n26082);
   U13672 : NAND2_X2 port map( A1 => n31244, A2 => n10825, ZN => n3550);
   U13674 : INV_X2 port map( I => n30143, ZN => n636);
   U13676 : XOR2_X1 port map( A1 => n1589, A2 => n1588, Z => n30143);
   U13677 : NAND2_X2 port map( A1 => n29307, A2 => n24171, ZN => n24191);
   U13687 : NOR2_X2 port map( A1 => n29307, A2 => n24171, ZN => n24273);
   U13706 : NAND2_X2 port map( A1 => n4683, A2 => n320, ZN => n6338);
   U13711 : NOR2_X2 port map( A1 => n30148, A2 => n8354, ZN => n8797);
   U13714 : XOR2_X1 port map( A1 => n30149, A2 => n9116, Z => n19788);
   U13715 : XOR2_X1 port map( A1 => n19785, A2 => n19786, Z => n30149);
   U13719 : OAI21_X2 port map( A1 => n16096, A2 => n29402, B => n751, ZN => 
                           n30151);
   U13728 : XNOR2_X1 port map( A1 => n32894, A2 => n25541, ZN => n30722);
   U13736 : XOR2_X1 port map( A1 => n9683, A2 => n5462, Z => n27957);
   U13742 : NAND2_X2 port map( A1 => n27159, A2 => n17310, ZN => n26459);
   U13751 : NAND2_X2 port map( A1 => n22845, A2 => n14882, ZN => n23287);
   U13759 : OAI22_X2 port map( A1 => n14232, A2 => n27577, B1 => n14133, B2 => 
                           n13720, ZN => n23956);
   U13762 : INV_X2 port map( I => n25657, ZN => n26322);
   U13771 : XOR2_X1 port map( A1 => n27952, A2 => n12954, Z => n23905);
   U13777 : NAND2_X2 port map( A1 => n795, A2 => n29307, ZN => n23991);
   U13779 : NAND2_X1 port map( A1 => n11960, A2 => n33813, ZN => n17562);
   U13780 : XOR2_X1 port map( A1 => n23389, A2 => n23444, Z => n23296);
   U13795 : XOR2_X1 port map( A1 => n8154, A2 => n30559, Z => n627);
   U13799 : XOR2_X1 port map( A1 => n14499, A2 => n29345, Z => n671);
   U13811 : XOR2_X1 port map( A1 => n27882, A2 => n27881, Z => n28343);
   U13821 : NAND2_X1 port map( A1 => n30458, A2 => n30157, ZN => n31065);
   U13822 : AOI22_X1 port map( A1 => n17845, A2 => n25606, B1 => n25612, B2 => 
                           n32856, ZN => n30157);
   U13836 : XOR2_X1 port map( A1 => n20794, A2 => n20706, Z => n20708);
   U13842 : XOR2_X1 port map( A1 => n2672, A2 => n30159, Z => n87);
   U13846 : XOR2_X1 port map( A1 => n2671, A2 => n19732, Z => n30159);
   U13847 : NAND2_X2 port map( A1 => n32866, A2 => n2234, ZN => n2654);
   U13855 : NAND3_X2 port map( A1 => n24115, A2 => n3213, A3 => n3212, ZN => 
                           n24116);
   U13860 : NOR2_X2 port map( A1 => n22724, A2 => n22723, ZN => n23103);
   U13864 : NAND2_X2 port map( A1 => n26324, A2 => n26178, ZN => n22724);
   U13865 : OR2_X1 port map( A1 => n7941, A2 => n5492, Z => n5112);
   U13890 : XOR2_X1 port map( A1 => n19539, A2 => n19384, Z => n19721);
   U13893 : NOR2_X2 port map( A1 => n18457, A2 => n18458, ZN => n19539);
   U13894 : NAND2_X2 port map( A1 => n2729, A2 => n30169, ZN => n13175);
   U13896 : OR2_X1 port map( A1 => n5889, A2 => n19108, Z => n12034);
   U13904 : NAND2_X2 port map( A1 => n5632, A2 => n9219, ZN => n24295);
   U13937 : XOR2_X1 port map( A1 => n2356, A2 => n21009, Z => n7016);
   U13938 : XOR2_X1 port map( A1 => n30173, A2 => n31869, Z => n686);
   U13940 : BUF_X4 port map( I => n17361, Z => n3506);
   U13944 : BUF_X2 port map( I => n18879, Z => n16588);
   U13945 : AOI21_X2 port map( A1 => n15827, A2 => n26726, B => n26725, ZN => 
                           n27472);
   U13946 : NAND2_X2 port map( A1 => n30174, A2 => n1763, ZN => n9629);
   U13949 : XOR2_X1 port map( A1 => n19376, A2 => n19377, Z => n16324);
   U13971 : NAND2_X2 port map( A1 => n30175, A2 => n18320, ZN => n8379);
   U13974 : XOR2_X1 port map( A1 => n30177, A2 => n30176, Z => n21266);
   U13976 : XOR2_X1 port map( A1 => n20889, A2 => n20850, Z => n30176);
   U13982 : XOR2_X1 port map( A1 => n20664, A2 => n20663, Z => n30177);
   U13983 : NAND2_X1 port map( A1 => n17543, A2 => n1101, ZN => n30198);
   U13985 : AOI21_X2 port map( A1 => n15286, A2 => n8558, B => n20136, ZN => 
                           n20139);
   U14014 : NOR2_X2 port map( A1 => n17698, A2 => n30180, ZN => n16519);
   U14015 : NOR3_X1 port map( A1 => n4248, A2 => n9518, A3 => n21311, ZN => 
                           n30180);
   U14024 : NAND2_X2 port map( A1 => n16435, A2 => n18481, ZN => n18604);
   U14030 : NAND2_X1 port map( A1 => n13669, A2 => n13668, ZN => n26713);
   U14045 : BUF_X2 port map( I => n3935, Z => n30183);
   U14058 : XOR2_X1 port map( A1 => n32255, A2 => n10075, Z => n1937);
   U14060 : XOR2_X1 port map( A1 => n1441, A2 => n29386, Z => n31184);
   U14061 : NAND2_X2 port map( A1 => n9954, A2 => n23031, ZN => n30442);
   U14065 : NAND3_X2 port map( A1 => n11700, A2 => n4082, A3 => n21137, ZN => 
                           n21496);
   U14069 : XOR2_X1 port map( A1 => n20552, A2 => n20752, Z => n10789);
   U14093 : INV_X2 port map( I => n30187, ZN => n31915);
   U14094 : NOR3_X2 port map( A1 => n28037, A2 => n32644, A3 => n924, ZN => 
                           n26411);
   U14098 : OAI21_X2 port map( A1 => n951, A2 => n17557, B => n12989, ZN => 
                           n26203);
   U14104 : INV_X2 port map( I => n26203, ZN => n13752);
   U14105 : NAND2_X2 port map( A1 => n12567, A2 => n12565, ZN => n30193);
   U14113 : XOR2_X1 port map( A1 => n19432, A2 => n19435, Z => n30188);
   U14121 : XOR2_X1 port map( A1 => n23501, A2 => n30189, Z => n5158);
   U14122 : XOR2_X1 port map( A1 => n11193, A2 => n5157, Z => n30189);
   U14124 : NAND2_X1 port map( A1 => n17439, A2 => n1329, ZN => n2833);
   U14129 : NOR2_X2 port map( A1 => n11621, A2 => n13308, ZN => n23946);
   U14130 : INV_X2 port map( I => n13764, ZN => n16853);
   U14133 : XOR2_X1 port map( A1 => n23505, A2 => n14492, Z => n30190);
   U14177 : INV_X2 port map( I => n1787, ZN => n2356);
   U14179 : NAND2_X2 port map( A1 => n15662, A2 => n30195, ZN => n20736);
   U14184 : OAI22_X2 port map( A1 => n32068, A2 => n20451, B1 => n20450, B2 => 
                           n5471, ZN => n30195);
   U14196 : XOR2_X1 port map( A1 => n20737, A2 => n20738, Z => n20739);
   U14206 : XOR2_X1 port map( A1 => n20964, A2 => n500, Z => n8701);
   U14207 : XOR2_X1 port map( A1 => n31950, A2 => n2789, Z => n20964);
   U14222 : OAI22_X2 port map( A1 => n5653, A2 => n19121, B1 => n1051, B2 => 
                           n19148, ZN => n31438);
   U14225 : OR2_X1 port map( A1 => n25665, A2 => n25664, Z => n25651);
   U14236 : AOI21_X2 port map( A1 => n25292, A2 => n5468, B => n7081, ZN => 
                           n11069);
   U14237 : NAND2_X2 port map( A1 => n30198, A2 => n23927, ZN => n15227);
   U14241 : XOR2_X1 port map( A1 => n19386, A2 => n1363, Z => n19168);
   U14245 : XOR2_X1 port map( A1 => n30199, A2 => n24991, Z => Ciphertext(25));
   U14249 : NAND2_X2 port map( A1 => n6768, A2 => n6767, ZN => n7879);
   U14271 : XOR2_X1 port map( A1 => n30203, A2 => n16010, Z => n27201);
   U14273 : XOR2_X1 port map( A1 => n7211, A2 => n12715, Z => n30203);
   U14274 : NOR2_X2 port map( A1 => n2158, A2 => n2156, ZN => n24805);
   U14280 : XOR2_X1 port map( A1 => n24743, A2 => n7838, Z => n7984);
   U14284 : NAND2_X2 port map( A1 => n26120, A2 => n27184, ZN => n24073);
   U14287 : NAND2_X1 port map( A1 => n15528, A2 => n24511, ZN => n30204);
   U14289 : OAI22_X2 port map( A1 => n17906, A2 => n14664, B1 => n28365, B2 => 
                           n16097, ZN => n10763);
   U14294 : OR2_X1 port map( A1 => n24315, A2 => n13232, Z => n16152);
   U14304 : NAND2_X2 port map( A1 => n4730, A2 => n30207, ZN => n9153);
   U14326 : INV_X2 port map( I => n32886, ZN => n25620);
   U14328 : XOR2_X1 port map( A1 => n17498, A2 => n6397, Z => n17499);
   U14340 : BUF_X2 port map( I => n23587, Z => n23588);
   U14345 : NOR2_X1 port map( A1 => n12049, A2 => n25617, ZN => n30497);
   U14349 : INV_X2 port map( I => n32887, ZN => n789);
   U14363 : INV_X4 port map( I => n20414, ZN => n1150);
   U14365 : OAI21_X2 port map( A1 => n32746, A2 => n14761, B => n873, ZN => 
                           n11510);
   U14371 : XOR2_X1 port map( A1 => n23218, A2 => n15742, Z => n13498);
   U14373 : AOI22_X2 port map( A1 => n10108, A2 => n26251, B1 => n10107, B2 => 
                           n850, ZN => n23218);
   U14379 : AOI21_X2 port map( A1 => n7361, A2 => n29141, B => n890, ZN => 
                           n9824);
   U14380 : OAI21_X2 port map( A1 => n23035, A2 => n23034, B => n13063, ZN => 
                           n12446);
   U14382 : XOR2_X1 port map( A1 => n30214, A2 => n7908, Z => n29230);
   U14403 : BUF_X2 port map( I => n10469, Z => n30318);
   U14406 : NAND2_X2 port map( A1 => n18279, A2 => n18278, ZN => n31451);
   U14409 : XOR2_X1 port map( A1 => n30216, A2 => n671, Z => n9932);
   U14411 : XOR2_X1 port map( A1 => n24450, A2 => n16738, Z => n30216);
   U14415 : NOR2_X2 port map( A1 => n31459, A2 => n31333, ZN => n30879);
   U14417 : XOR2_X1 port map( A1 => n20896, A2 => n30218, Z => n4756);
   U14419 : XOR2_X1 port map( A1 => n15275, A2 => n4758, Z => n30218);
   U14420 : XOR2_X1 port map( A1 => n30220, A2 => n31405, Z => n25762);
   U14425 : NAND3_X1 port map( A1 => n932, A2 => n28011, A3 => n7242, ZN => 
                           n17298);
   U14429 : NAND2_X2 port map( A1 => n8854, A2 => n25594, ZN => n25615);
   U14433 : XOR2_X1 port map( A1 => n23171, A2 => n16672, Z => n6091);
   U14438 : NOR2_X2 port map( A1 => n8079, A2 => n21793, ZN => n30223);
   U14441 : NOR2_X2 port map( A1 => n932, A2 => n7242, ZN => n10351);
   U14444 : NAND2_X2 port map( A1 => n9408, A2 => n9407, ZN => n30943);
   U14445 : XOR2_X1 port map( A1 => n225, A2 => n30224, Z => n17050);
   U14446 : XOR2_X1 port map( A1 => n4792, A2 => n4467, Z => n30224);
   U14447 : NAND3_X1 port map( A1 => n14562, A2 => n15160, A3 => n11915, ZN => 
                           n14561);
   U14448 : BUF_X2 port map( I => n33566, Z => n16459);
   U14464 : NAND2_X2 port map( A1 => n12849, A2 => n14455, ZN => n19744);
   U14467 : OAI21_X2 port map( A1 => n28385, A2 => n10093, B => n30225, ZN => 
                           n21463);
   U14469 : OAI21_X2 port map( A1 => n24052, A2 => n30595, B => n9973, ZN => 
                           n5968);
   U14478 : INV_X2 port map( I => n3519, ZN => n23532);
   U14479 : NAND2_X2 port map( A1 => n32253, A2 => n8379, ZN => n19215);
   U14480 : XOR2_X1 port map( A1 => n10130, A2 => n8609, Z => n412);
   U14481 : XOR2_X1 port map( A1 => n30380, A2 => n23536, Z => n10130);
   U14484 : INV_X2 port map( I => n17941, ZN => n12105);
   U14490 : BUF_X2 port map( I => n24335, Z => n30230);
   U14504 : XOR2_X1 port map( A1 => n26256, A2 => n30815, Z => n31467);
   U14513 : INV_X2 port map( I => n18994, ZN => n14893);
   U14515 : NAND2_X2 port map( A1 => n29330, A2 => n32887, ZN => n6915);
   U14517 : INV_X2 port map( I => n15955, ZN => n15956);
   U14519 : AOI21_X1 port map( A1 => n13528, A2 => n25555, B => n30232, ZN => 
                           n13527);
   U14522 : OAI22_X1 port map( A1 => n28759, A2 => n6391, B1 => n25555, B2 => 
                           n12864, ZN => n30232);
   U14526 : NOR2_X2 port map( A1 => n20087, A2 => n20086, ZN => n9115);
   U14528 : NOR2_X2 port map( A1 => n7182, A2 => n27954, ZN => n30233);
   U14533 : OR2_X1 port map( A1 => n24910, A2 => n24909, Z => n10754);
   U14536 : XOR2_X1 port map( A1 => n30235, A2 => n18019, Z => Ciphertext(178))
                           ;
   U14541 : NAND3_X1 port map( A1 => n27217, A2 => n18021, A3 => n18020, ZN => 
                           n30235);
   U14552 : INV_X1 port map( I => n30236, ZN => n2197);
   U14554 : XOR2_X1 port map( A1 => n17745, A2 => n16816, Z => n5601);
   U14562 : XOR2_X1 port map( A1 => n30237, A2 => n20966, Z => n17999);
   U14564 : XOR2_X1 port map( A1 => n13681, A2 => n33219, Z => n30237);
   U14567 : INV_X2 port map( I => n25855, ZN => n25858);
   U14569 : NAND2_X2 port map( A1 => n12697, A2 => n17627, ZN => n30293);
   U14595 : NAND2_X2 port map( A1 => n11899, A2 => n25756, ZN => n5292);
   U14596 : XOR2_X1 port map( A1 => n23166, A2 => n23199, Z => n3905);
   U14601 : XOR2_X1 port map( A1 => n23266, A2 => n11891, Z => n23199);
   U14635 : NAND2_X2 port map( A1 => n2045, A2 => n10358, ZN => n30248);
   U14636 : INV_X1 port map( I => n31560, ZN => n23601);
   U14637 : XOR2_X1 port map( A1 => n17128, A2 => n5244, Z => n8361);
   U14641 : XOR2_X1 port map( A1 => n29137, A2 => n4285, Z => n5244);
   U14652 : INV_X1 port map( I => n2861, ZN => n31629);
   U14659 : NAND2_X2 port map( A1 => n30779, A2 => n28754, ZN => n30389);
   U14660 : NOR2_X2 port map( A1 => n29224, A2 => n25678, ZN => n27173);
   U14661 : NOR2_X2 port map( A1 => n24438, A2 => n24437, ZN => n29224);
   U14665 : XOR2_X1 port map( A1 => n27868, A2 => n30250, Z => n28624);
   U14676 : XOR2_X1 port map( A1 => n19658, A2 => n27138, Z => n19659);
   U14691 : NAND2_X1 port map( A1 => n22455, A2 => n7965, ZN => n30833);
   U14699 : NAND2_X2 port map( A1 => n20429, A2 => n31533, ZN => n20594);
   U14700 : XOR2_X1 port map( A1 => n24762, A2 => n24626, Z => n8893);
   U14701 : INV_X2 port map( I => n8834, ZN => n30252);
   U14714 : AOI22_X2 port map( A1 => n6660, A2 => n33992, B1 => n16600, B2 => 
                           n21628, ZN => n21776);
   U14715 : INV_X2 port map( I => n21626, ZN => n16600);
   U14722 : NOR2_X2 port map( A1 => n31084, A2 => n31083, ZN => n27914);
   U14737 : AND2_X1 port map( A1 => n2317, A2 => n20376, Z => n2316);
   U14745 : NAND2_X2 port map( A1 => n9378, A2 => n8866, ZN => n2575);
   U14749 : XOR2_X1 port map( A1 => n30257, A2 => n5726, Z => n5725);
   U14755 : XOR2_X1 port map( A1 => n20693, A2 => n20776, Z => n12609);
   U14764 : NAND2_X2 port map( A1 => n20004, A2 => n20003, ZN => n20693);
   U14765 : NAND2_X2 port map( A1 => n24728, A2 => n30259, ZN => n14915);
   U14775 : NOR2_X1 port map( A1 => n146, A2 => n25763, ZN => n24715);
   U14779 : BUF_X4 port map( I => n20483, Z => n21306);
   U14787 : NAND2_X2 port map( A1 => n30262, A2 => n7027, ZN => n7197);
   U14788 : NAND2_X1 port map( A1 => n12174, A2 => n12173, ZN => n30262);
   U14798 : NOR2_X1 port map( A1 => n25607, A2 => n10504, ZN => n10501);
   U14810 : NAND2_X2 port map( A1 => n24716, A2 => n24717, ZN => n25818);
   U14815 : INV_X1 port map( I => n8243, ZN => n28308);
   U14816 : XNOR2_X1 port map( A1 => n2305, A2 => n30849, ZN => n8243);
   U14830 : XOR2_X1 port map( A1 => n17859, A2 => n12538, Z => n1538);
   U14836 : OR2_X1 port map( A1 => n23003, A2 => n23000, Z => n31225);
   U14840 : NAND2_X2 port map( A1 => n30342, A2 => n7815, ZN => n5863);
   U14848 : NAND2_X2 port map( A1 => n6369, A2 => n13043, ZN => n13638);
   U14859 : XOR2_X1 port map( A1 => n15776, A2 => n29441, Z => n30387);
   U14861 : XOR2_X1 port map( A1 => n17026, A2 => n30265, Z => n30713);
   U14871 : NAND2_X2 port map( A1 => n1882, A2 => n5944, ZN => n30506);
   U14876 : OAI21_X2 port map( A1 => n6661, A2 => n28671, B => n4026, ZN => 
                           n4025);
   U14878 : NAND2_X2 port map( A1 => n27426, A2 => n13943, ZN => n12616);
   U14902 : NAND2_X2 port map( A1 => n951, A2 => n5473, ZN => n31710);
   U14903 : NAND2_X2 port map( A1 => n13764, A2 => n12864, ZN => n17403);
   U14914 : OAI22_X2 port map( A1 => n18118, A2 => n9127, B1 => n4993, B2 => 
                           n16113, ZN => n9017);
   U14930 : INV_X2 port map( I => n19289, ZN => n745);
   U14935 : OAI21_X1 port map( A1 => n7397, A2 => n7836, B => n20628, ZN => 
                           n7396);
   U14966 : INV_X1 port map( I => n22598, ZN => n22595);
   U14969 : AOI22_X1 port map( A1 => n1521, A2 => n836, B1 => n1522, B2 => 
                           n25901, ZN => n26793);
   U14972 : AOI21_X1 port map( A1 => n24724, A2 => n29771, B => n836, ZN => 
                           n8299);
   U14977 : OR2_X1 port map( A1 => n22336, A2 => n22486, Z => n22416);
   U14991 : NAND2_X1 port map( A1 => n24104, A2 => n18077, ZN => n30459);
   U14993 : NAND3_X1 port map( A1 => n15770, A2 => n17717, A3 => n28136, ZN => 
                           n24585);
   U15015 : OAI22_X1 port map( A1 => n18828, A2 => n16782, B1 => n17231, B2 => 
                           n16915, ZN => n4279);
   U15016 : NAND3_X1 port map( A1 => n17053, A2 => n21767, A3 => n21520, ZN => 
                           n1648);
   U15023 : NOR2_X1 port map( A1 => n9127, A2 => n4993, ZN => n30269);
   U15024 : NOR2_X1 port map( A1 => n757, A2 => n23940, ZN => n13677);
   U15032 : INV_X1 port map( I => n24479, ZN => n31762);
   U15041 : NAND2_X1 port map( A1 => n24735, A2 => n9126, ZN => n13944);
   U15042 : BUF_X4 port map( I => n16315, Z => n13597);
   U15047 : INV_X1 port map( I => n19261, ZN => n28544);
   U15049 : NAND2_X1 port map( A1 => n21537, A2 => n8196, ZN => n22308);
   U15052 : NAND2_X1 port map( A1 => n5741, A2 => n29307, ZN => n30270);
   U15053 : NAND3_X1 port map( A1 => n24130, A2 => n32515, A3 => n974, ZN => 
                           n8005);
   U15054 : OAI21_X1 port map( A1 => n1858, A2 => n1861, B => n25227, ZN => 
                           n26380);
   U15055 : XOR2_X1 port map( A1 => n18388, A2 => Key(111), Z => n30271);
   U15056 : AND2_X1 port map( A1 => n4651, A2 => n4650, Z => n30272);
   U15058 : INV_X2 port map( I => Plaintext(111), ZN => n18388);
   U15064 : INV_X1 port map( I => n1227, ZN => n24648);
   U15068 : XNOR2_X1 port map( A1 => n16448, A2 => n13864, ZN => n30273);
   U15069 : INV_X2 port map( I => n31772, ZN => n31918);
   U15084 : INV_X2 port map( I => n21455, ZN => n780);
   U15102 : NAND2_X1 port map( A1 => n115, A2 => n34084, ZN => n22286);
   U15112 : CLKBUF_X12 port map( I => n23720, Z => n16620);
   U15121 : AND3_X1 port map( A1 => n17963, A2 => n11045, A3 => n25903, Z => 
                           n10792);
   U15125 : INV_X1 port map( I => n18655, ZN => n6118);
   U15128 : AND3_X2 port map( A1 => n25342, A2 => n25341, A3 => n25340, Z => 
                           n30276);
   U15130 : OAI21_X1 port map( A1 => n25712, A2 => n25711, B => n27208, ZN => 
                           n31403);
   U15134 : NAND2_X1 port map( A1 => n355, A2 => n6882, ZN => n3597);
   U15145 : AOI22_X1 port map( A1 => n11469, A2 => n965, B1 => n24960, B2 => 
                           n24948, ZN => n24950);
   U15147 : NAND2_X1 port map( A1 => n31564, A2 => n22871, ZN => n30638);
   U15155 : NAND2_X1 port map( A1 => n6338, A2 => n6337, ZN => n21315);
   U15160 : NAND2_X1 port map( A1 => n28037, A2 => n924, ZN => n2468);
   U15163 : NOR2_X1 port map( A1 => n924, A2 => n9678, ZN => n1553);
   U15164 : NOR2_X1 port map( A1 => n5883, A2 => n924, ZN => n26369);
   U15171 : NOR3_X1 port map( A1 => n21568, A2 => n30389, A3 => n21569, ZN => 
                           n21351);
   U15173 : OAI21_X1 port map( A1 => n14983, A2 => n21569, B => n30389, ZN => 
                           n3580);
   U15189 : NAND2_X1 port map( A1 => n837, A2 => n967, ZN => n13464);
   U15195 : NOR2_X1 port map( A1 => n29269, A2 => n23681, ZN => n8535);
   U15202 : NAND2_X1 port map( A1 => n22314, A2 => n22549, ZN => n22315);
   U15213 : XOR2_X1 port map( A1 => n9868, A2 => n30278, Z => n30277);
   U15214 : XNOR2_X1 port map( A1 => n24774, A2 => n1948, ZN => n30278);
   U15220 : NOR2_X1 port map( A1 => n9127, A2 => n4993, ZN => n28223);
   U15222 : INV_X2 port map( I => n25707, ZN => n25708);
   U15225 : NAND2_X1 port map( A1 => n27864, A2 => n27863, ZN => n24020);
   U15241 : INV_X1 port map( I => n24133, ZN => n27864);
   U15243 : AND2_X1 port map( A1 => n24052, A2 => n29157, Z => n31424);
   U15244 : INV_X2 port map( I => n17133, ZN => n23872);
   U15245 : AND3_X2 port map( A1 => n23695, A2 => n18182, A3 => n17133, Z => 
                           n31396);
   U15248 : INV_X2 port map( I => n22824, ZN => n723);
   U15254 : NAND2_X1 port map( A1 => n24913, A2 => n27248, ZN => n8278);
   U15266 : NOR2_X1 port map( A1 => n14686, A2 => n15852, ZN => n5689);
   U15282 : INV_X2 port map( I => n14686, ZN => n15039);
   U15283 : OAI21_X1 port map( A1 => n25760, A2 => n33976, B => n25712, ZN => 
                           n24438);
   U15287 : NAND3_X1 port map( A1 => n8902, A2 => n749, A3 => n1204, ZN => 
                           n1946);
   U15297 : NAND2_X2 port map( A1 => n2997, A2 => n30855, ZN => n30279);
   U15298 : NOR2_X2 port map( A1 => n2999, A2 => n2998, ZN => n2997);
   U15312 : NAND2_X1 port map( A1 => n28691, A2 => n32176, ZN => n11436);
   U15316 : INV_X2 port map( I => n21300, ZN => n6082);
   U15317 : OAI21_X1 port map( A1 => n20791, A2 => n20790, B => n6082, ZN => 
                           n3973);
   U15320 : NAND2_X1 port map( A1 => n1808, A2 => n7581, ZN => n24132);
   U15331 : NAND2_X1 port map( A1 => n10135, A2 => n1332, ZN => n30342);
   U15332 : NAND2_X1 port map( A1 => n25343, A2 => n25344, ZN => n14244);
   U15348 : CLKBUF_X4 port map( I => n25855, Z => n14199);
   U15349 : NOR2_X1 port map( A1 => n14681, A2 => n21704, ZN => n21595);
   U15353 : INV_X2 port map( I => n14681, ZN => n21705);
   U15361 : NOR2_X1 port map( A1 => n21816, A2 => n1137, ZN => n6626);
   U15362 : NAND2_X1 port map( A1 => n21816, A2 => n31958, ZN => n21818);
   U15364 : NAND2_X1 port map( A1 => n254, A2 => n3019, ZN => n24881);
   U15372 : NAND2_X1 port map( A1 => n9953, A2 => n10354, ZN => n22406);
   U15373 : INV_X1 port map( I => n10354, ZN => n1000);
   U15380 : NAND2_X1 port map( A1 => n25604, A2 => n27057, ZN => n28775);
   U15384 : NAND2_X1 port map( A1 => n16633, A2 => n16239, ZN => n15442);
   U15386 : INV_X2 port map( I => n17721, ZN => n23867);
   U15390 : INV_X1 port map( I => n23025, ZN => n23653);
   U15418 : INV_X1 port map( I => n11931, ZN => n831);
   U15448 : NAND2_X1 port map( A1 => n22377, A2 => n17936, ZN => n28225);
   U15454 : NOR2_X1 port map( A1 => n11931, A2 => n10174, ZN => n25606);
   U15462 : AOI21_X1 port map( A1 => n10497, A2 => n25713, B => n10393, ZN => 
                           n11511);
   U15470 : NAND3_X2 port map( A1 => n12399, A2 => n9736, A3 => n26069, ZN => 
                           n29131);
   U15473 : NOR2_X1 port map( A1 => n12541, A2 => n2958, ZN => n10419);
   U15474 : NAND2_X1 port map( A1 => n20525, A2 => n2958, ZN => n2957);
   U15494 : CLKBUF_X4 port map( I => n5988, Z => n5926);
   U15498 : AOI21_X1 port map( A1 => n26887, A2 => n22808, B => n26886, ZN => 
                           n26885);
   U15505 : NAND2_X1 port map( A1 => n34089, A2 => n13989, ZN => n21181);
   U15508 : INV_X1 port map( I => n13989, ZN => n17467);
   U15517 : INV_X2 port map( I => n8168, ZN => n221);
   U15518 : NAND2_X1 port map( A1 => n9342, A2 => n24031, ZN => n24142);
   U15522 : NAND2_X1 port map( A1 => n26479, A2 => n8079, ZN => n6619);
   U15527 : OAI21_X1 port map( A1 => n21479, A2 => n21711, B => n21496, ZN => 
                           n21480);
   U15531 : AOI21_X1 port map( A1 => n28623, A2 => n16985, B => n12374, ZN => 
                           n16984);
   U15537 : NOR2_X1 port map( A1 => n16984, A2 => n16983, ZN => n16982);
   U15538 : NAND2_X1 port map( A1 => n11943, A2 => n651, ZN => n9772);
   U15549 : INV_X1 port map( I => n23916, ZN => n23920);
   U15550 : NAND2_X1 port map( A1 => n13326, A2 => n24985, ZN => n14269);
   U15555 : NAND3_X1 port map( A1 => n907, A2 => n10206, A3 => n856, ZN => 
                           n13892);
   U15556 : INV_X1 port map( I => n907, ZN => n10907);
   U15558 : INV_X1 port map( I => n14865, ZN => n714);
   U15569 : NAND2_X2 port map( A1 => n2000, A2 => n2001, ZN => n30288);
   U15572 : INV_X1 port map( I => n2795, ZN => n11587);
   U15581 : INV_X1 port map( I => n3718, ZN => n24211);
   U15582 : NAND2_X1 port map( A1 => n17426, A2 => n3718, ZN => n7060);
   U15585 : OAI21_X1 port map( A1 => n11132, A2 => n25339, B => n10569, ZN => 
                           n25338);
   U15586 : OR2_X2 port map( A1 => n10569, A2 => n14788, Z => n3430);
   U15594 : NOR2_X1 port map( A1 => n16066, A2 => n4151, ZN => n17069);
   U15595 : INV_X2 port map( I => n16066, ZN => n24285);
   U15597 : NAND2_X1 port map( A1 => n21805, A2 => n17077, ZN => n10689);
   U15601 : NAND2_X1 port map( A1 => n19220, A2 => n30995, ZN => n18475);
   U15602 : NOR2_X1 port map( A1 => n19220, A2 => n30995, ZN => n31757);
   U15603 : AND2_X1 port map( A1 => n4025, A2 => n27341, Z => n30289);
   U15610 : AOI21_X1 port map( A1 => n12485, A2 => n10822, B => n25066, ZN => 
                           n31206);
   U15612 : NAND2_X1 port map( A1 => n13622, A2 => n30584, ZN => n22745);
   U15618 : OAI21_X1 port map( A1 => n5864, A2 => n5865, B => n16809, ZN => 
                           n30961);
   U15620 : NOR2_X2 port map( A1 => n16815, A2 => n26966, ZN => n30290);
   U15624 : NOR2_X1 port map( A1 => n11298, A2 => n4184, ZN => n18088);
   U15625 : OAI21_X1 port map( A1 => n32652, A2 => n2092, B => n25120, ZN => 
                           n16611);
   U15631 : NAND2_X1 port map( A1 => n25121, A2 => n2092, ZN => n14867);
   U15644 : NAND2_X1 port map( A1 => n25412, A2 => n25405, ZN => n25299);
   U15646 : NAND3_X1 port map( A1 => n32602, A2 => n10955, A3 => n843, ZN => 
                           n9225);
   U15647 : INV_X2 port map( I => n10955, ZN => n17694);
   U15648 : BUF_X2 port map( I => n23639, Z => n14078);
   U15651 : NAND2_X1 port map( A1 => n23735, A2 => n23765, ZN => n30296);
   U15652 : NAND3_X1 port map( A1 => n24213, A2 => n24210, A3 => n24209, ZN => 
                           n23987);
   U15656 : NAND2_X1 port map( A1 => n22622, A2 => n22497, ZN => n22628);
   U15681 : NOR2_X1 port map( A1 => n8576, A2 => n20029, ZN => n30474);
   U15686 : OAI22_X1 port map( A1 => n14793, A2 => n14747, B1 => n20155, B2 => 
                           n3486, ZN => n5347);
   U15693 : NAND2_X1 port map( A1 => n16812, A2 => n27808, ZN => n6671);
   U15698 : OR2_X1 port map( A1 => n25429, A2 => n17948, Z => n25415);
   U15703 : INV_X1 port map( I => n27189, ZN => n25745);
   U15708 : CLKBUF_X12 port map( I => Key(185), Z => n25493);
   U15724 : NAND2_X2 port map( A1 => n11439, A2 => n11440, ZN => n30301);
   U15738 : XNOR2_X1 port map( A1 => n23371, A2 => n23530, ZN => n23249);
   U15743 : OAI21_X2 port map( A1 => n14247, A2 => n14245, B => n14243, ZN => 
                           n30302);
   U15746 : CLKBUF_X4 port map( I => n14577, Z => n1647);
   U15757 : OAI21_X2 port map( A1 => n18959, A2 => n4622, B => n4619, ZN => 
                           n30305);
   U15775 : NAND3_X1 port map( A1 => n21433, A2 => n4683, A3 => n5049, ZN => 
                           n8603);
   U15786 : NAND2_X1 port map( A1 => n11438, A2 => n29157, ZN => n11236);
   U15805 : NAND2_X1 port map( A1 => n8057, A2 => n28451, ZN => n20301);
   U15806 : INV_X1 port map( I => n20301, ZN => n6559);
   U15820 : OAI22_X1 port map( A1 => n24909, A2 => n10099, B1 => n24911, B2 => 
                           n24910, ZN => n24916);
   U15822 : NAND2_X1 port map( A1 => n30816, A2 => n4097, ZN => n31202);
   U15852 : NAND2_X1 port map( A1 => n21308, A2 => n16180, ZN => n21309);
   U15853 : NOR3_X1 port map( A1 => n21307, A2 => n21443, A3 => n21306, ZN => 
                           n21230);
   U15857 : NAND2_X1 port map( A1 => n19290, A2 => n27726, ZN => n3204);
   U15865 : NAND2_X1 port map( A1 => n4580, A2 => n16486, ZN => n22905);
   U15871 : NAND2_X1 port map( A1 => n9522, A2 => n24148, ZN => n2153);
   U15872 : NOR2_X1 port map( A1 => n24881, A2 => n30279, ZN => n27062);
   U15881 : OAI21_X1 port map( A1 => n5631, A2 => n9219, B => n4286, ZN => 
                           n10103);
   U15884 : INV_X1 port map( I => n19654, ZN => n30766);
   U15894 : AOI22_X1 port map( A1 => n7813, A2 => n7811, B1 => n5863, B2 => 
                           n21870, ZN => n10493);
   U15907 : AOI22_X2 port map( A1 => n31284, A2 => n34098, B1 => n21495, B2 => 
                           n1014, ZN => n30309);
   U15908 : AOI22_X1 port map( A1 => n31284, A2 => n34098, B1 => n21495, B2 => 
                           n1014, ZN => n22080);
   U15919 : NAND2_X1 port map( A1 => n10847, A2 => n29628, ZN => n11616);
   U15926 : NOR2_X1 port map( A1 => n14133, A2 => n12287, ZN => n30991);
   U15938 : NAND2_X1 port map( A1 => n21504, A2 => n21749, ZN => n11585);
   U15947 : INV_X1 port map( I => n30033, ZN => n21690);
   U15949 : INV_X2 port map( I => n16528, ZN => n25405);
   U15956 : NOR2_X1 port map( A1 => n10112, A2 => n29866, ZN => n4522);
   U15957 : XOR2_X1 port map( A1 => n4228, A2 => n7477, Z => n30311);
   U15958 : NAND2_X1 port map( A1 => n25277, A2 => n25276, ZN => n25271);
   U15976 : NOR2_X1 port map( A1 => n25780, A2 => n12611, ZN => n25774);
   U15989 : XNOR2_X1 port map( A1 => n18095, A2 => n16820, ZN => n30313);
   U15994 : NAND3_X1 port map( A1 => n6111, A2 => n13624, A3 => n30285, ZN => 
                           n10035);
   U15997 : NOR2_X1 port map( A1 => n7004, A2 => n13191, ZN => n2712);
   U15999 : CLKBUF_X4 port map( I => n11722, Z => n11370);
   U16013 : OAI21_X1 port map( A1 => n17726, A2 => n8045, B => n30252, ZN => 
                           n9382);
   U16020 : NOR2_X1 port map( A1 => n7083, A2 => n25653, ZN => n25645);
   U16021 : NAND2_X1 port map( A1 => n7083, A2 => n25659, ZN => n25644);
   U16029 : AOI21_X1 port map( A1 => n7083, A2 => n25653, B => n25657, ZN => 
                           n11211);
   U16045 : AND3_X1 port map( A1 => n25403, A2 => n30308, A3 => n25295, Z => 
                           n11259);
   U16047 : INV_X1 port map( I => n3405, ZN => n30316);
   U16052 : INV_X1 port map( I => n10469, ZN => n14940);
   U16055 : INV_X2 port map( I => n25334, ZN => n25390);
   U16058 : OR2_X1 port map( A1 => n17133, A2 => n8694, Z => n23640);
   U16085 : OR2_X1 port map( A1 => n29658, A2 => n15519, Z => n13466);
   U16086 : NAND2_X1 port map( A1 => n26322, A2 => n7083, ZN => n6497);
   U16087 : INV_X1 port map( I => n9517, ZN => n19515);
   U16090 : OAI22_X1 port map( A1 => n8950, A2 => n7373, B1 => n7370, B2 => 
                           n7369, ZN => n6526);
   U16097 : INV_X1 port map( I => n22063, ZN => n1128);
   U16103 : NOR2_X1 port map( A1 => n9041, A2 => n9042, ZN => n30322);
   U16122 : INV_X2 port map( I => n23833, ZN => n17726);
   U16131 : NAND2_X1 port map( A1 => n25317, A2 => n31407, ZN => n25315);
   U16138 : INV_X2 port map( I => n8606, ZN => n19357);
   U16151 : NAND2_X1 port map( A1 => n7312, A2 => n10339, ZN => n30326);
   U16152 : NOR2_X1 port map( A1 => n13279, A2 => n18581, ZN => n8627);
   U16153 : NAND2_X1 port map( A1 => n490, A2 => n18581, ZN => n18583);
   U16156 : NAND2_X1 port map( A1 => n18581, A2 => n31821, ZN => n31820);
   U16158 : INV_X1 port map( I => n14770, ZN => n24346);
   U16170 : NAND2_X1 port map( A1 => n6075, A2 => n4755, ZN => n30666);
   U16171 : INV_X2 port map( I => n4755, ZN => n30784);
   U16180 : NOR2_X1 port map( A1 => n30473, A2 => n24025, ZN => n30328);
   U16182 : OAI21_X1 port map( A1 => n16406, A2 => n1573, B => n32760, ZN => 
                           n25033);
   U16184 : NAND2_X2 port map( A1 => n2394, A2 => n2393, ZN => n30329);
   U16206 : INV_X1 port map( I => n25666, ZN => n25660);
   U16215 : NOR2_X2 port map( A1 => n22820, A2 => n22819, ZN => n23120);
   U16228 : NOR2_X1 port map( A1 => n7273, A2 => n7371, ZN => n16833);
   U16230 : AOI22_X1 port map( A1 => n7339, A2 => n7371, B1 => n14737, B2 => 
                           n16973, ZN => n30740);
   U16231 : OAI21_X1 port map( A1 => n7371, A2 => n32059, B => n3489, ZN => 
                           n7370);
   U16232 : INV_X2 port map( I => n28839, ZN => n899);
   U16240 : AND2_X2 port map( A1 => n23035, A2 => n28839, Z => n17740);
   U16241 : NAND2_X1 port map( A1 => n26261, A2 => n3469, ZN => n30332);
   U16253 : NAND3_X1 port map( A1 => n27785, A2 => n20575, A3 => n31968, ZN => 
                           n8143);
   U16259 : AOI22_X1 port map( A1 => n22509, A2 => n15601, B1 => n987, B2 => 
                           n22508, ZN => n6503);
   U16262 : NOR2_X1 port map( A1 => n987, A2 => n22955, ZN => n6300);
   U16267 : AOI21_X1 port map( A1 => n13532, A2 => n967, B => n9858, ZN => 
                           n9857);
   U16273 : NAND2_X1 port map( A1 => n26566, A2 => n20577, ZN => n20244);
   U16290 : INV_X2 port map( I => n27021, ZN => n7968);
   U16291 : OR3_X2 port map( A1 => n29306, A2 => n24171, A3 => n3483, Z => 
                           n15781);
   U16292 : NOR2_X1 port map( A1 => n1181, A2 => n339, ZN => n11080);
   U16293 : OR2_X2 port map( A1 => n30059, A2 => n28069, Z => n23600);
   U16295 : INV_X1 port map( I => n15077, ZN => n19961);
   U16298 : AND2_X1 port map( A1 => n15077, A2 => n5870, Z => n5871);
   U16299 : NAND2_X1 port map( A1 => n8062, A2 => n4897, ZN => n4999);
   U16332 : INV_X1 port map( I => n11707, ZN => n328);
   U16346 : NOR2_X1 port map( A1 => n10943, A2 => n31254, ZN => n26037);
   U16355 : INV_X1 port map( I => n10943, ZN => n11876);
   U16358 : NOR2_X1 port map( A1 => n13129, A2 => n28942, ZN => n13066);
   U16376 : INV_X1 port map( I => n10579, ZN => n3152);
   U16377 : AND2_X2 port map( A1 => n4036, A2 => n11599, Z => n18812);
   U16383 : OR2_X2 port map( A1 => n4036, A2 => n11599, Z => n2733);
   U16384 : AOI22_X1 port map( A1 => n18450, A2 => n17477, B1 => n18677, B2 => 
                           n18662, ZN => n28943);
   U16391 : AOI21_X1 port map( A1 => n17478, A2 => n18660, B => n18677, ZN => 
                           n31427);
   U16396 : NAND2_X1 port map( A1 => n20635, A2 => n4693, ZN => n30970);
   U16398 : AOI21_X1 port map( A1 => n28408, A2 => n22949, B => n805, ZN => 
                           n6802);
   U16400 : NOR2_X1 port map( A1 => n28555, A2 => n31129, ZN => n17483);
   U16403 : NAND2_X2 port map( A1 => n6950, A2 => n6952, ZN => n8870);
   U16405 : AND2_X1 port map( A1 => n31324, A2 => n19049, Z => n12927);
   U16406 : NAND2_X2 port map( A1 => n13752, A2 => n14859, ZN => n31324);
   U16408 : INV_X2 port map( I => n13363, ZN => n18581);
   U16412 : XOR2_X1 port map( A1 => Plaintext(153), A2 => Key(153), Z => n13363
                           );
   U16413 : XOR2_X1 port map( A1 => n5503, A2 => n5875, Z => n31576);
   U16415 : XNOR2_X1 port map( A1 => n22123, A2 => n13564, ZN => n5875);
   U16419 : NAND2_X2 port map( A1 => n14815, A2 => n14572, ZN => n20124);
   U16420 : NAND2_X1 port map( A1 => n31127, A2 => n31126, ZN => n11706);
   U16424 : XNOR2_X1 port map( A1 => n12868, A2 => n13236, ZN => n1227);
   U16445 : XOR2_X1 port map( A1 => n14682, A2 => n26575, Z => n30338);
   U16447 : XOR2_X1 port map( A1 => n32050, A2 => n30339, Z => n6833);
   U16448 : XOR2_X1 port map( A1 => n23294, A2 => n25815, Z => n30339);
   U16449 : OAI21_X2 port map( A1 => n17414, A2 => n30340, B => n10848, ZN => 
                           n28967);
   U16453 : NAND2_X2 port map( A1 => n12449, A2 => n30341, ZN => n23388);
   U16455 : AOI22_X1 port map( A1 => n11210, A2 => n22961, B1 => n13396, B2 => 
                           n22962, ZN => n30341);
   U16456 : XNOR2_X1 port map( A1 => n21964, A2 => n2894, ZN => n21951);
   U16459 : OAI21_X2 port map( A1 => n26899, A2 => n10346, B => n10343, ZN => 
                           n2894);
   U16473 : AOI21_X2 port map( A1 => n28306, A2 => n8760, B => n30344, ZN => 
                           n10500);
   U16478 : NOR2_X2 port map( A1 => n5759, A2 => n23920, ZN => n30344);
   U16479 : INV_X2 port map( I => n30345, ZN => n30731);
   U16483 : XOR2_X1 port map( A1 => n4136, A2 => n28446, Z => n30345);
   U16486 : XOR2_X1 port map( A1 => n20781, A2 => n20783, Z => n3117);
   U16494 : NAND2_X1 port map( A1 => n7485, A2 => n24312, ZN => n30348);
   U16499 : XOR2_X1 port map( A1 => n20746, A2 => n20993, Z => n9815);
   U16500 : NAND3_X1 port map( A1 => n10243, A2 => n10244, A3 => n11895, ZN => 
                           n30349);
   U16503 : XOR2_X1 port map( A1 => n22255, A2 => n30571, Z => n7160);
   U16525 : NAND2_X1 port map( A1 => n14174, A2 => n4518, ZN => n16265);
   U16537 : NAND2_X2 port map( A1 => n19450, A2 => n18089, ZN => n3310);
   U16543 : OAI21_X1 port map( A1 => n30353, A2 => n15746, B => n22690, ZN => 
                           n3451);
   U16548 : NOR2_X1 port map( A1 => n1122, A2 => n31931, ZN => n30353);
   U16556 : NAND2_X2 port map( A1 => n1641, A2 => n26224, ZN => n30354);
   U16559 : OAI21_X2 port map( A1 => n30357, A2 => n30356, B => n12947, ZN => 
                           n20344);
   U16562 : OR2_X1 port map( A1 => n18151, A2 => n15295, Z => n25637);
   U16563 : XOR2_X1 port map( A1 => n16158, A2 => n18109, Z => n19552);
   U16564 : AOI22_X2 port map( A1 => n2124, A2 => n28276, B1 => n30602, B2 => 
                           n2123, ZN => n18109);
   U16567 : NOR2_X1 port map( A1 => n515, A2 => n10433, ZN => n4382);
   U16573 : NAND2_X2 port map( A1 => n8897, A2 => n16797, ZN => n14588);
   U16584 : AND2_X1 port map( A1 => n31408, A2 => n19971, Z => n31514);
   U16586 : NOR2_X1 port map( A1 => n33809, A2 => n27491, ZN => n30475);
   U16597 : NOR2_X2 port map( A1 => n8062, A2 => n14490, ZN => n24176);
   U16598 : AND2_X2 port map( A1 => n18655, A2 => n32358, Z => n18894);
   U16601 : BUF_X4 port map( I => n7600, Z => n30602);
   U16604 : NAND2_X2 port map( A1 => n21637, A2 => n21633, ZN => n12792);
   U16605 : OAI21_X2 port map( A1 => n5978, A2 => n21244, B => n17803, ZN => 
                           n21637);
   U16606 : BUF_X2 port map( I => n19991, Z => n30366);
   U16608 : OAI21_X1 port map( A1 => n29438, A2 => n23045, B => n6553, ZN => 
                           n29114);
   U16611 : XOR2_X1 port map( A1 => n24551, A2 => n30367, Z => n26754);
   U16613 : XOR2_X1 port map( A1 => n24620, A2 => n16662, Z => n30367);
   U16621 : INV_X1 port map( I => n8275, ZN => n902);
   U16623 : XOR2_X1 port map( A1 => n21927, A2 => n30368, Z => n4859);
   U16626 : XOR2_X1 port map( A1 => n10006, A2 => n8356, Z => n30368);
   U16634 : XOR2_X1 port map( A1 => n13661, A2 => n30370, Z => n31098);
   U16635 : XOR2_X1 port map( A1 => n14613, A2 => n24999, Z => n30370);
   U16648 : NAND3_X1 port map( A1 => n29958, A2 => n1577, A3 => n8334, ZN => 
                           n14516);
   U16659 : AOI22_X2 port map( A1 => n29383, A2 => n31653, B1 => n21744, B2 => 
                           n17021, ZN => n17692);
   U16690 : INV_X2 port map( I => n17679, ZN => n31493);
   U16691 : NAND2_X2 port map( A1 => n17680, A2 => n17681, ZN => n17679);
   U16698 : INV_X2 port map( I => n20818, ZN => n31526);
   U16703 : NOR2_X2 port map( A1 => n20246, A2 => n20245, ZN => n20818);
   U16704 : NOR2_X2 port map( A1 => n17685, A2 => n16282, ZN => n21604);
   U16716 : XOR2_X1 port map( A1 => n21937, A2 => n11819, Z => n8596);
   U16719 : XOR2_X1 port map( A1 => n22189, A2 => n22055, Z => n21937);
   U16726 : OAI21_X1 port map( A1 => n7197, A2 => n31970, B => n825, ZN => 
                           n17593);
   U16728 : NAND2_X2 port map( A1 => n4025, A2 => n27341, ZN => n13601);
   U16730 : AOI21_X2 port map( A1 => n30379, A2 => n2574, B => n32248, ZN => 
                           n27973);
   U16737 : XOR2_X1 port map( A1 => n8761, A2 => n30381, Z => n29209);
   U16738 : XOR2_X1 port map( A1 => n23536, A2 => n23189, Z => n30381);
   U16743 : XOR2_X1 port map( A1 => n30382, A2 => n31534, Z => n14576);
   U16747 : XOR2_X1 port map( A1 => n19653, A2 => n18051, Z => n30382);
   U16753 : XOR2_X1 port map( A1 => n30385, A2 => n8249, Z => n8813);
   U16754 : XOR2_X1 port map( A1 => n20654, A2 => n30045, Z => n30385);
   U16755 : NAND2_X2 port map( A1 => n3962, A2 => n13107, ZN => n5748);
   U16762 : NOR2_X2 port map( A1 => n30442, A2 => n773, ZN => n31273);
   U16765 : XOR2_X1 port map( A1 => n29244, A2 => n8972, Z => n6957);
   U16768 : XOR2_X1 port map( A1 => n6081, A2 => n30240, Z => n8972);
   U16781 : NAND2_X2 port map( A1 => n8245, A2 => n30386, ZN => n8168);
   U16783 : INV_X2 port map( I => n30387, ZN => n6344);
   U16784 : NAND2_X2 port map( A1 => n15599, A2 => n15597, ZN => n10174);
   U16800 : INV_X2 port map( I => n30390, ZN => n15424);
   U16808 : INV_X2 port map( I => n7811, ZN => n27685);
   U16810 : NAND2_X2 port map( A1 => n4208, A2 => n12619, ZN => n22964);
   U16812 : NAND2_X2 port map( A1 => n7610, A2 => n28681, ZN => n12619);
   U16814 : XOR2_X1 port map( A1 => n10870, A2 => n24652, Z => n24653);
   U16826 : OAI21_X2 port map( A1 => n2604, A2 => n2605, B => n30391, ZN => 
                           n3286);
   U16829 : OAI21_X2 port map( A1 => n2602, A2 => n2603, B => n29207, ZN => 
                           n30391);
   U16833 : OAI21_X2 port map( A1 => n10735, A2 => n30441, B => n11552, ZN => 
                           n10935);
   U16835 : XOR2_X1 port map( A1 => n23473, A2 => n770, Z => n6094);
   U16840 : XOR2_X1 port map( A1 => n1302, A2 => n22256, Z => n4136);
   U16844 : XOR2_X1 port map( A1 => n29898, A2 => n12459, Z => n14875);
   U16847 : NAND2_X2 port map( A1 => n30394, A2 => n10160, ZN => n11789);
   U16848 : XOR2_X1 port map( A1 => n28730, A2 => n30495, Z => n11128);
   U16856 : XOR2_X1 port map( A1 => n5127, A2 => n15236, Z => n2362);
   U16860 : NAND2_X2 port map( A1 => n8692, A2 => n19204, ZN => n5127);
   U16865 : INV_X2 port map( I => n30047, ZN => n25467);
   U16874 : INV_X2 port map( I => n25883, ZN => n25872);
   U16882 : NOR3_X1 port map( A1 => n30401, A2 => n19013, A3 => n19009, ZN => 
                           n19014);
   U16886 : XOR2_X1 port map( A1 => n24478, A2 => n24516, Z => n24806);
   U16888 : NAND2_X2 port map( A1 => n24166, A2 => n24165, ZN => n24516);
   U16895 : NAND3_X1 port map( A1 => n6497, A2 => n25643, A3 => n25658, ZN => 
                           n26745);
   U16908 : XOR2_X1 port map( A1 => n30402, A2 => n1604, Z => n22224);
   U16911 : AOI22_X2 port map( A1 => n5488, A2 => n67, B1 => n2574, B2 => n1632
                           , ZN => n30403);
   U16939 : NAND2_X2 port map( A1 => n12746, A2 => n21423, ZN => n5978);
   U16940 : XOR2_X1 port map( A1 => n1338, A2 => n20843, Z => n20674);
   U16958 : XOR2_X1 port map( A1 => n8359, A2 => n28162, Z => n8358);
   U16973 : INV_X1 port map( I => n7672, ZN => n30973);
   U16976 : AOI22_X1 port map( A1 => n12928, A2 => n27743, B1 => n13925, B2 => 
                           n12927, ZN => n13002);
   U16979 : NAND2_X2 port map( A1 => n19046, A2 => n19041, ZN => n27743);
   U16988 : XOR2_X1 port map( A1 => n16076, A2 => n30041, Z => n23407);
   U17002 : XOR2_X1 port map( A1 => n2592, A2 => n2590, Z => n2589);
   U17005 : BUF_X2 port map( I => n31658, Z => n30412);
   U17030 : NAND2_X2 port map( A1 => n30417, A2 => n3508, ZN => n7603);
   U17037 : XOR2_X1 port map( A1 => n30418, A2 => n24937, Z => Ciphertext(11));
   U17038 : NAND2_X1 port map( A1 => n7787, A2 => n31348, ZN => n30418);
   U17049 : NOR2_X2 port map( A1 => n7430, A2 => n12363, ZN => n26268);
   U17055 : XOR2_X1 port map( A1 => n23383, A2 => n30420, Z => n27673);
   U17056 : XOR2_X1 port map( A1 => n26426, A2 => n23536, Z => n30420);
   U17070 : NOR2_X2 port map( A1 => n30423, A2 => n25634, ZN => n26581);
   U17073 : NOR2_X2 port map( A1 => n11090, A2 => n3405, ZN => n25632);
   U17099 : XOR2_X1 port map( A1 => n30309, A2 => n32885, Z => n22039);
   U17100 : OAI21_X1 port map( A1 => n9472, A2 => n21870, B => n5385, ZN => 
                           n5384);
   U17106 : INV_X2 port map( I => n27655, ZN => n2795);
   U17107 : XOR2_X1 port map( A1 => n2796, A2 => n19687, Z => n27655);
   U17113 : XOR2_X1 port map( A1 => n7630, A2 => n7675, Z => n30427);
   U17117 : NAND2_X2 port map( A1 => n8995, A2 => n30428, ZN => n8997);
   U17118 : AND2_X1 port map( A1 => n10063, A2 => n8996, Z => n30428);
   U17123 : NAND2_X2 port map( A1 => n30429, A2 => n22822, ZN => n9185);
   U17125 : NAND2_X1 port map( A1 => n16203, A2 => n16202, ZN => n30429);
   U17126 : NOR3_X1 port map( A1 => n21872, A2 => n9472, A3 => n7811, ZN => 
                           n4220);
   U17143 : AOI21_X2 port map( A1 => n20247, A2 => n20248, B => n17732, ZN => 
                           n20717);
   U17145 : XOR2_X1 port map( A1 => n1468, A2 => n1466, Z => n25150);
   U17180 : XOR2_X1 port map( A1 => n23419, A2 => n14819, Z => n11290);
   U17183 : NAND2_X2 port map( A1 => n31096, A2 => n14147, ZN => n17941);
   U17191 : XOR2_X1 port map( A1 => n30439, A2 => n16253, Z => Ciphertext(117))
                           ;
   U17194 : NOR2_X1 port map( A1 => n25511, A2 => n1945, ZN => n30439);
   U17195 : INV_X2 port map( I => n21655, ZN => n30441);
   U17203 : XOR2_X1 port map( A1 => n27545, A2 => n8306, Z => n24812);
   U17216 : INV_X2 port map( I => n30444, ZN => n26606);
   U17219 : XOR2_X1 port map( A1 => n3303, A2 => n3304, Z => n30444);
   U17220 : INV_X2 port map( I => n30445, ZN => n11272);
   U17226 : BUF_X2 port map( I => n15360, Z => n31554);
   U17227 : NAND2_X2 port map( A1 => n30446, A2 => n15745, ZN => n9303);
   U17236 : NAND2_X2 port map( A1 => n25581, A2 => n1082, ZN => n15287);
   U17238 : OAI22_X2 port map( A1 => n16413, A2 => n25707, B1 => n25621, B2 => 
                           n11944, ZN => n25581);
   U17239 : AOI21_X2 port map( A1 => n30641, A2 => n30448, B => n22644, ZN => 
                           n27867);
   U17241 : BUF_X4 port map( I => n3989, Z => n31080);
   U17249 : NAND2_X2 port map( A1 => n26990, A2 => n7360, ZN => n7358);
   U17284 : XOR2_X1 port map( A1 => n5509, A2 => n30453, Z => n23157);
   U17287 : XOR2_X1 port map( A1 => n5508, A2 => n29291, Z => n30453);
   U17307 : AND2_X1 port map( A1 => n16022, A2 => n14045, Z => n28491);
   U17317 : XOR2_X1 port map( A1 => n7234, A2 => n7235, Z => n7453);
   U17318 : NAND2_X1 port map( A1 => n5704, A2 => n15716, ZN => n17333);
   U17327 : AOI21_X1 port map( A1 => n25611, A2 => n27262, B => n27528, ZN => 
                           n30458);
   U17331 : OAI22_X1 port map( A1 => n710, A2 => n3157, B1 => n28261, B2 => 
                           n30130, ZN => n1964);
   U17332 : NOR2_X2 port map( A1 => n6398, A2 => n16924, ZN => n28261);
   U17342 : NAND2_X2 port map( A1 => n28307, A2 => n30515, ZN => n23974);
   U17352 : XOR2_X1 port map( A1 => n14935, A2 => n30462, Z => n5432);
   U17355 : XOR2_X1 port map( A1 => n14937, A2 => n7829, Z => n30462);
   U17356 : NOR2_X2 port map( A1 => n1312, A2 => n21466, ZN => n21465);
   U17360 : XOR2_X1 port map( A1 => n5630, A2 => n5629, Z => n30463);
   U17364 : XOR2_X1 port map( A1 => n21026, A2 => n2525, Z => n2524);
   U17365 : OR2_X2 port map( A1 => n16440, A2 => n15559, Z => n9073);
   U17366 : NAND2_X1 port map( A1 => n31309, A2 => n11208, ZN => n21708);
   U17369 : XOR2_X1 port map( A1 => n30465, A2 => n12260, Z => n29254);
   U17371 : XOR2_X1 port map( A1 => n11062, A2 => n30466, Z => n30465);
   U17375 : INV_X1 port map( I => n19748, ZN => n30466);
   U17382 : OAI21_X2 port map( A1 => n28757, A2 => n18609, B => n18608, ZN => 
                           n30467);
   U17384 : NOR2_X2 port map( A1 => n31309, A2 => n21655, ZN => n21797);
   U17385 : NAND2_X2 port map( A1 => n30469, A2 => n7733, ZN => n19332);
   U17389 : NAND2_X2 port map( A1 => n2391, A2 => n20156, ZN => n5470);
   U17393 : NAND2_X2 port map( A1 => n31275, A2 => n5373, ZN => n30470);
   U17396 : XOR2_X1 port map( A1 => n1644, A2 => n1642, Z => n23668);
   U17406 : NAND2_X2 port map( A1 => n26956, A2 => n9046, ZN => n14194);
   U17409 : XOR2_X1 port map( A1 => n22150, A2 => n9208, Z => n9207);
   U17415 : NAND2_X1 port map( A1 => n30731, A2 => n11805, ZN => n22544);
   U17423 : XOR2_X1 port map( A1 => n24786, A2 => n24776, Z => n24518);
   U17425 : NOR2_X2 port map( A1 => n30475, A2 => n30474, ZN => n20433);
   U17428 : NAND2_X2 port map( A1 => n15074, A2 => n15073, ZN => n19703);
   U17437 : NAND2_X1 port map( A1 => n21847, A2 => n30291, ZN => n30479);
   U17439 : NAND2_X2 port map( A1 => n30480, A2 => n8459, ZN => n9809);
   U17440 : OAI21_X2 port map( A1 => n29405, A2 => n26298, B => n1016, ZN => 
                           n30480);
   U17454 : XOR2_X1 port map( A1 => n20832, A2 => n8997, Z => n18180);
   U17461 : OAI22_X1 port map( A1 => n966, A2 => n25214, B1 => n5578, B2 => 
                           n16509, ZN => n25223);
   U17467 : NOR2_X2 port map( A1 => n26528, A2 => n18259, ZN => n25214);
   U17469 : BUF_X2 port map( I => n5511, Z => n30482);
   U17472 : NOR2_X1 port map( A1 => n8334, A2 => n1577, ZN => n11210);
   U17474 : XOR2_X1 port map( A1 => n6052, A2 => n6054, Z => n16757);
   U17475 : AOI22_X2 port map( A1 => n8856, A2 => n21214, B1 => n15428, B2 => 
                           n21372, ZN => n30483);
   U17481 : XOR2_X1 port map( A1 => n30486, A2 => n2889, Z => n30861);
   U17490 : BUF_X2 port map( I => n4219, Z => n30489);
   U17505 : XOR2_X1 port map( A1 => n23272, A2 => n5399, Z => n23334);
   U17508 : AOI21_X2 port map( A1 => n18073, A2 => n9456, B => n29222, ZN => 
                           n16260);
   U17514 : XOR2_X1 port map( A1 => n30493, A2 => n30290, Z => n24369);
   U17517 : OAI21_X2 port map( A1 => n11637, A2 => n20575, B => n20571, ZN => 
                           n5590);
   U17518 : OR2_X1 port map( A1 => n1877, A2 => n14436, Z => n27605);
   U17521 : NAND2_X2 port map( A1 => n28235, A2 => n11079, ZN => n30505);
   U17530 : AOI21_X1 port map( A1 => n25692, A2 => n25691, B => n30494, ZN => 
                           n30521);
   U17534 : AOI21_X1 port map( A1 => n2017, A2 => n2016, B => n26447, ZN => 
                           n30494);
   U17539 : OAI22_X1 port map( A1 => n30497, A2 => n17845, B1 => n25618, B2 => 
                           n10174, ZN => n17844);
   U17540 : INV_X2 port map( I => n30498, ZN => n490);
   U17542 : XOR2_X1 port map( A1 => Plaintext(151), A2 => Key(151), Z => n30498
                           );
   U17545 : XOR2_X1 port map( A1 => n19544, A2 => n19545, Z => n13441);
   U17553 : BUF_X2 port map( I => n23066, Z => n30502);
   U17568 : NAND2_X1 port map( A1 => n10812, A2 => n30508, ZN => n23965);
   U17575 : OR2_X1 port map( A1 => n31155, A2 => n11754, Z => n30508);
   U17592 : OAI21_X2 port map( A1 => n30511, A2 => n21514, B => n30243, ZN => 
                           n31404);
   U17593 : XOR2_X1 port map( A1 => n30513, A2 => n29082, Z => n28640);
   U17595 : XOR2_X1 port map( A1 => n27875, A2 => n11897, Z => n30513);
   U17608 : XOR2_X1 port map( A1 => n32564, A2 => n30306, Z => n15822);
   U17610 : NAND2_X2 port map( A1 => n21525, A2 => n21524, ZN => n22306);
   U17614 : XOR2_X1 port map( A1 => n20808, A2 => n20645, Z => n30514);
   U17630 : XOR2_X1 port map( A1 => n24756, A2 => n30517, Z => n1466);
   U17632 : XOR2_X1 port map( A1 => n30358, A2 => n30069, Z => n30517);
   U17641 : NOR2_X1 port map( A1 => n15283, A2 => n9934, ZN => n9847);
   U17648 : NAND2_X1 port map( A1 => n33928, A2 => n28934, ZN => n28349);
   U17650 : XOR2_X1 port map( A1 => n30521, A2 => n25694, Z => Ciphertext(148))
                           ;
   U17654 : AOI22_X2 port map( A1 => n27565, A2 => n12254, B1 => n29232, B2 => 
                           n12256, ZN => n8040);
   U17656 : XOR2_X1 port map( A1 => n17775, A2 => n23218, Z => n23399);
   U17660 : INV_X1 port map( I => n7503, ZN => n30586);
   U17664 : AND2_X1 port map( A1 => n29270, A2 => n14398, Z => n6759);
   U17667 : XOR2_X1 port map( A1 => n15710, A2 => n16253, Z => n30524);
   U17686 : AOI22_X1 port map( A1 => n14434, A2 => n1206, B1 => n690, B2 => 
                           n25916, ZN => n14433);
   U17693 : XOR2_X1 port map( A1 => n27841, A2 => n30069, Z => n24418);
   U17708 : INV_X2 port map( I => n30526, ZN => n17963);
   U17710 : XOR2_X1 port map( A1 => n17703, A2 => n29450, Z => n26597);
   U17721 : INV_X2 port map( I => n1994, ZN => n16138);
   U17723 : NOR2_X2 port map( A1 => n11770, A2 => n13859, ZN => n11769);
   U17729 : XOR2_X1 port map( A1 => n16831, A2 => n3629, Z => n20894);
   U17736 : XNOR2_X1 port map( A1 => n21946, A2 => n10370, ZN => n30575);
   U17744 : AOI21_X2 port map( A1 => n16883, A2 => n20220, B => n30530, ZN => 
                           n14428);
   U17770 : XOR2_X1 port map( A1 => n2854, A2 => n30317, Z => n30535);
   U17772 : XOR2_X1 port map( A1 => n30536, A2 => n4719, Z => n17903);
   U17773 : XOR2_X1 port map( A1 => n24797, A2 => n12239, Z => n30536);
   U17776 : XOR2_X1 port map( A1 => n18024, A2 => n18025, Z => n11677);
   U17789 : NAND2_X2 port map( A1 => n30537, A2 => n29406, ZN => n3773);
   U17793 : NOR2_X2 port map( A1 => n30538, A2 => n17584, ZN => n30537);
   U17795 : AOI21_X2 port map( A1 => n6876, A2 => n23032, B => n31273, ZN => 
                           n14610);
   U17806 : XOR2_X1 port map( A1 => n14103, A2 => n30541, Z => n23639);
   U17815 : XOR2_X1 port map( A1 => n23446, A2 => n11667, Z => n30541);
   U17820 : XOR2_X1 port map( A1 => n4797, A2 => n30542, Z => n9750);
   U17823 : XOR2_X1 port map( A1 => n22110, A2 => n13437, Z => n30542);
   U17832 : XOR2_X1 port map( A1 => n20856, A2 => n20785, Z => n9040);
   U17833 : INV_X1 port map( I => n29263, ZN => n1122);
   U17836 : XOR2_X1 port map( A1 => n27792, A2 => n5126, Z => n29263);
   U17850 : XOR2_X1 port map( A1 => n16893, A2 => n22264, Z => n6058);
   U17852 : OAI21_X2 port map( A1 => n30546, A2 => n28911, B => n4602, ZN => 
                           n20569);
   U17859 : XOR2_X1 port map( A1 => n23113, A2 => n13123, Z => n30547);
   U17861 : OAI21_X2 port map( A1 => n276, A2 => n517, B => n21777, ZN => 
                           n30548);
   U17868 : XOR2_X1 port map( A1 => n22198, A2 => n22197, Z => n14755);
   U17870 : BUF_X2 port map( I => n21592, Z => n30549);
   U17878 : XOR2_X1 port map( A1 => n32881, A2 => n28005, Z => n30550);
   U17883 : OAI22_X2 port map( A1 => n1908, A2 => n31374, B1 => n30552, B2 => 
                           n30551, ZN => n5647);
   U17888 : XOR2_X1 port map( A1 => n13321, A2 => n5742, Z => n23471);
   U17890 : NAND2_X2 port map( A1 => n10849, A2 => n31454, ZN => n30553);
   U17896 : BUF_X2 port map( I => n27097, Z => n30554);
   U17899 : XOR2_X1 port map( A1 => n30556, A2 => n5980, Z => n5979);
   U17910 : XOR2_X1 port map( A1 => n28315, A2 => n30557, Z => n30556);
   U17918 : NAND2_X2 port map( A1 => n14774, A2 => n14776, ZN => n28934);
   U17926 : XOR2_X1 port map( A1 => n26094, A2 => n16700, Z => n30559);
   U17927 : NOR2_X2 port map( A1 => n9133, A2 => n31040, ZN => n21152);
   U17934 : INV_X2 port map( I => n30563, ZN => n16738);
   U17940 : NAND2_X1 port map( A1 => n5991, A2 => n28825, ZN => n30564);
   U17947 : XOR2_X1 port map( A1 => n23355, A2 => n31554, Z => n30565);
   U17953 : XOR2_X1 port map( A1 => n19473, A2 => n32267, Z => n9577);
   U17954 : NAND2_X1 port map( A1 => n29424, A2 => n26803, ZN => n30658);
   U17957 : NAND2_X1 port map( A1 => n9990, A2 => n10098, ZN => n30587);
   U17962 : OAI21_X2 port map( A1 => n30569, A2 => n30568, B => n11992, ZN => 
                           n9982);
   U17963 : AOI22_X1 port map( A1 => n6825, A2 => n14922, B1 => n13273, B2 => 
                           n9162, ZN => n6824);
   U17973 : NAND2_X2 port map( A1 => n8743, A2 => n25109, ZN => n25128);
   U17980 : NAND2_X2 port map( A1 => n18205, A2 => n6228, ZN => n20835);
   U17984 : NAND2_X1 port map( A1 => n25944, A2 => n8253, ZN => n11597);
   U17985 : INV_X2 port map( I => n30570, ZN => n1736);
   U17997 : NAND2_X2 port map( A1 => n7550, A2 => n7551, ZN => n8770);
   U17999 : XOR2_X1 port map( A1 => n19668, A2 => n253, Z => n4883);
   U18001 : AOI21_X2 port map( A1 => n10073, A2 => n28104, B => n14757, ZN => 
                           n19668);
   U18008 : XOR2_X1 port map( A1 => n16727, A2 => n6488, Z => n19660);
   U18018 : OR2_X1 port map( A1 => n20109, A2 => n28183, Z => n30614);
   U18022 : XOR2_X1 port map( A1 => n10917, A2 => n30574, Z => n10916);
   U18023 : XOR2_X1 port map( A1 => n31750, A2 => n9434, Z => n30574);
   U18034 : XOR2_X1 port map( A1 => n10154, A2 => n30575, Z => n28589);
   U18040 : NAND2_X1 port map( A1 => n31306, A2 => n5477, ZN => n15193);
   U18044 : INV_X1 port map( I => n9107, ZN => n23096);
   U18068 : NOR2_X1 port map( A1 => n12973, A2 => n21241, ZN => n11405);
   U18071 : INV_X1 port map( I => n21330, ZN => n12973);
   U18082 : XOR2_X1 port map( A1 => n20778, A2 => n13725, Z => n13724);
   U18087 : NOR2_X2 port map( A1 => n19172, A2 => n19078, ZN => n11875);
   U18092 : NAND2_X2 port map( A1 => n1376, A2 => n10943, ZN => n19172);
   U18106 : XOR2_X1 port map( A1 => n20925, A2 => n20927, Z => n7032);
   U18112 : XOR2_X1 port map( A1 => n2520, A2 => n31394, Z => n23126);
   U18116 : NAND2_X2 port map( A1 => n18160, A2 => n18162, ZN => n30995);
   U18126 : NOR3_X1 port map( A1 => n25026, A2 => n25025, A3 => n25024, ZN => 
                           n31320);
   U18128 : XOR2_X1 port map( A1 => n24424, A2 => n4720, Z => n4719);
   U18134 : XOR2_X1 port map( A1 => n7731, A2 => n24440, Z => n24424);
   U18136 : XOR2_X1 port map( A1 => n30583, A2 => n25038, Z => Ciphertext(37));
   U18142 : NOR2_X2 port map( A1 => n24008, A2 => n10033, ZN => n26027);
   U18147 : NAND2_X2 port map( A1 => n31163, A2 => n27679, ZN => n27676);
   U18149 : NOR2_X1 port map( A1 => n14133, A2 => n29203, ZN => n14529);
   U18150 : NAND3_X1 port map( A1 => n7302, A2 => n7299, A3 => n7298, ZN => 
                           Ciphertext(72));
   U18157 : NAND2_X2 port map( A1 => n1172, A2 => n7573, ZN => n19850);
   U18176 : OAI21_X2 port map( A1 => n7001, A2 => n26088, B => n2271, ZN => 
                           n6996);
   U18178 : XOR2_X1 port map( A1 => n13198, A2 => n29457, Z => n27868);
   U18187 : OAI21_X2 port map( A1 => n31938, A2 => n14513, B => n16099, ZN => 
                           n1776);
   U18188 : NOR2_X2 port map( A1 => n15038, A2 => n976, ZN => n14513);
   U18211 : OAI22_X1 port map( A1 => n898, A2 => n23066, B1 => n849, B2 => 
                           n4067, ZN => n4477);
   U18222 : INV_X2 port map( I => n30592, ZN => n12120);
   U18224 : XOR2_X1 port map( A1 => n18280, A2 => Key(64), Z => n30592);
   U18232 : INV_X2 port map( I => n30593, ZN => n6444);
   U18241 : NAND2_X2 port map( A1 => n5945, A2 => n29044, ZN => n6488);
   U18242 : BUF_X2 port map( I => n14123, Z => n30595);
   U18245 : XOR2_X1 port map( A1 => n30596, A2 => n23507, Z => n31429);
   U18256 : XOR2_X1 port map( A1 => n30597, A2 => n4186, Z => n11749);
   U18257 : XOR2_X1 port map( A1 => n11748, A2 => n21944, Z => n30597);
   U18260 : NAND2_X2 port map( A1 => n23627, A2 => n23626, ZN => n24479);
   U18264 : XOR2_X1 port map( A1 => n22302, A2 => n10292, Z => n7289);
   U18271 : NAND2_X2 port map( A1 => n2338, A2 => n31051, ZN => n10292);
   U18272 : XOR2_X1 port map( A1 => n7363, A2 => n23332, Z => n23383);
   U18275 : OAI22_X2 port map( A1 => n30598, A2 => n9066, B1 => n24199, B2 => 
                           n12574, ZN => n24764);
   U18282 : XOR2_X1 port map( A1 => n30601, A2 => n30600, Z => n26551);
   U18286 : XOR2_X1 port map( A1 => n13842, A2 => n19447, Z => n30601);
   U18307 : XOR2_X1 port map( A1 => n23162, A2 => n6169, Z => n1796);
   U18314 : NAND3_X2 port map( A1 => n30608, A2 => n28158, A3 => n28159, ZN => 
                           n22149);
   U18326 : XOR2_X1 port map( A1 => n30610, A2 => n5107, Z => n5106);
   U18336 : XOR2_X1 port map( A1 => n33572, A2 => n5109, Z => n30610);
   U18344 : INV_X1 port map( I => n16109, ZN => n31167);
   U18359 : NOR2_X2 port map( A1 => n5308, A2 => n7546, ZN => n24046);
   U18367 : NAND2_X2 port map( A1 => n30615, A2 => n25149, ZN => n25151);
   U18380 : XOR2_X1 port map( A1 => n5336, A2 => n6604, Z => n10932);
   U18383 : NAND2_X1 port map( A1 => n26237, A2 => n820, ZN => n9232);
   U18385 : AND2_X2 port map( A1 => n18186, A2 => n16417, Z => n18370);
   U18391 : NOR2_X1 port map( A1 => n31823, A2 => n20045, ZN => n30617);
   U18397 : NAND2_X2 port map( A1 => n30618, A2 => n39, ZN => n23368);
   U18398 : OAI21_X2 port map( A1 => n10885, A2 => n16236, B => n22900, ZN => 
                           n30618);
   U18433 : NAND3_X2 port map( A1 => n29335, A2 => n28472, A3 => n28473, ZN => 
                           n31181);
   U18434 : NAND3_X2 port map( A1 => n30623, A2 => n13161, A3 => n30622, ZN => 
                           n13651);
   U18445 : XOR2_X1 port map( A1 => n19546, A2 => n19591, Z => n3285);
   U18450 : NAND2_X1 port map( A1 => n18184, A2 => n28232, ZN => n9205);
   U18451 : NAND2_X2 port map( A1 => n30624, A2 => n2908, ZN => n20445);
   U18453 : OR2_X2 port map( A1 => n4735, A2 => n31287, Z => n2538);
   U18454 : NAND2_X2 port map( A1 => n11069, A2 => n3430, ZN => n5533);
   U18455 : NOR2_X2 port map( A1 => n29353, A2 => n30625, ZN => n10302);
   U18460 : NAND2_X1 port map( A1 => n5640, A2 => n33594, ZN => n22338);
   U18464 : NAND2_X2 port map( A1 => n30626, A2 => n4872, ZN => n24544);
   U18471 : OR3_X1 port map( A1 => n2958, A2 => n868, A3 => n8374, Z => n28353)
                           ;
   U18476 : NOR2_X1 port map( A1 => n15564, A2 => n11912, ZN => n30627);
   U18485 : OAI22_X2 port map( A1 => n31149, A2 => n25561, B1 => n25562, B2 => 
                           n25331, ZN => n25523);
   U18495 : NAND3_X2 port map( A1 => n6645, A2 => n6643, A3 => n14171, ZN => 
                           n20267);
   U18515 : XOR2_X1 port map( A1 => n13084, A2 => n13085, Z => n16913);
   U18528 : XOR2_X1 port map( A1 => n20924, A2 => n20885, Z => n14899);
   U18532 : NAND2_X2 port map( A1 => n28452, A2 => n28454, ZN => n14436);
   U18542 : AOI21_X2 port map( A1 => n14076, A2 => n4262, B => n8784, ZN => 
                           n30634);
   U18547 : XOR2_X1 port map( A1 => n30635, A2 => n4401, Z => n564);
   U18553 : INV_X2 port map( I => n10915, ZN => n30636);
   U18558 : AND2_X1 port map( A1 => n20479, A2 => n11637, Z => n28226);
   U18563 : AOI21_X1 port map( A1 => n22872, A2 => n15718, B => n30638, ZN => 
                           n30800);
   U18568 : XOR2_X1 port map( A1 => n22218, A2 => n1131, Z => n1716);
   U18577 : NAND2_X2 port map( A1 => n21292, A2 => n21291, ZN => n6669);
   U18586 : XOR2_X1 port map( A1 => n16150, A2 => n13435, Z => n30644);
   U18588 : NOR2_X2 port map( A1 => n30645, A2 => n29084, ZN => n8337);
   U18589 : NAND2_X2 port map( A1 => n30940, A2 => n517, ZN => n30645);
   U18592 : NAND2_X1 port map( A1 => n3203, A2 => n30677, ZN => n26207);
   U18600 : NAND2_X2 port map( A1 => n3001, A2 => n3003, ZN => n3203);
   U18620 : AOI22_X2 port map( A1 => n31990, A2 => n31175, B1 => n23788, B2 => 
                           n15272, ZN => n30649);
   U18629 : NAND2_X1 port map( A1 => n1134, A2 => n30652, ZN => n12995);
   U18642 : OAI21_X2 port map( A1 => n31934, A2 => n13127, B => n22444, ZN => 
                           n22878);
   U18646 : XOR2_X1 port map( A1 => n30653, A2 => n16030, Z => n3686);
   U18647 : XOR2_X1 port map( A1 => n6094, A2 => n17628, Z => n30653);
   U18656 : XOR2_X1 port map( A1 => n19636, A2 => n19635, Z => n19640);
   U18658 : XOR2_X1 port map( A1 => n22317, A2 => n156, Z => n21924);
   U18659 : NOR2_X2 port map( A1 => n21562, A2 => n21561, ZN => n156);
   U18668 : XOR2_X1 port map( A1 => n4574, A2 => n4572, Z => n24726);
   U18671 : INV_X4 port map( I => n11521, ZN => n13747);
   U18675 : INV_X1 port map( I => n27262, ZN => n17845);
   U18685 : NAND2_X2 port map( A1 => n18192, A2 => n25585, ZN => n27262);
   U18695 : INV_X2 port map( I => n16847, ZN => n30663);
   U18698 : OR2_X1 port map( A1 => n30663, A2 => n2581, Z => n30936);
   U18699 : INV_X1 port map( I => n22312, ZN => n31203);
   U18700 : INV_X2 port map( I => n18397, ZN => n18687);
   U18703 : XOR2_X1 port map( A1 => n18396, A2 => Key(183), Z => n18397);
   U18704 : XOR2_X1 port map( A1 => n19667, A2 => n19666, Z => n17689);
   U18710 : XOR2_X1 port map( A1 => n12048, A2 => n5462, Z => n19667);
   U18713 : XOR2_X1 port map( A1 => n26530, A2 => n21007, Z => n30664);
   U18719 : NAND2_X2 port map( A1 => n30824, A2 => n12465, ZN => n28580);
   U18729 : INV_X2 port map( I => n14600, ZN => n9293);
   U18735 : AOI22_X2 port map( A1 => n22375, A2 => n9411, B1 => n25947, B2 => 
                           n22479, ZN => n23000);
   U18737 : INV_X2 port map( I => n9168, ZN => n30668);
   U18740 : NOR2_X1 port map( A1 => n31150, A2 => n28949, ZN => n30670);
   U18744 : XOR2_X1 port map( A1 => n28086, A2 => n6790, Z => n31040);
   U18751 : AOI21_X2 port map( A1 => n24712, A2 => n24711, B => n1077, ZN => 
                           n25678);
   U18765 : OAI22_X1 port map( A1 => n1028, A2 => n7774, B1 => n2237, B2 => 
                           n7218, ZN => n9693);
   U18766 : INV_X2 port map( I => n11089, ZN => n3405);
   U18783 : XOR2_X1 port map( A1 => n24749, A2 => n5525, Z => n30676);
   U18797 : NAND2_X2 port map( A1 => n27232, A2 => n23547, ZN => n24283);
   U18799 : INV_X4 port map( I => n31668, ZN => n1351);
   U18801 : NAND2_X2 port map( A1 => n7820, A2 => n28622, ZN => n31668);
   U18807 : NAND2_X1 port map( A1 => n30961, A2 => n5866, ZN => n30777);
   U18808 : XOR2_X1 port map( A1 => n30679, A2 => n18932, Z => n26815);
   U18810 : NAND2_X2 port map( A1 => n14084, A2 => n19968, ZN => n20384);
   U18811 : NOR2_X2 port map( A1 => n13770, A2 => n27878, ZN => n30681);
   U18819 : BUF_X2 port map( I => n31324, Z => n30682);
   U18826 : XOR2_X1 port map( A1 => n15516, A2 => n20691, Z => n8682);
   U18832 : OAI22_X1 port map( A1 => n20332, A2 => n28390, B1 => n20549, B2 => 
                           n11710, ZN => n11709);
   U18833 : XOR2_X1 port map( A1 => n15329, A2 => n16506, Z => n10443);
   U18835 : NAND2_X2 port map( A1 => n12908, A2 => n12909, ZN => n15329);
   U18836 : INV_X2 port map( I => n7012, ZN => n14251);
   U18840 : XOR2_X1 port map( A1 => n11889, A2 => n29312, Z => n14820);
   U18841 : NAND2_X2 port map( A1 => n19311, A2 => n19312, ZN => n11889);
   U18842 : XOR2_X1 port map( A1 => n15236, A2 => n19668, Z => n13863);
   U18845 : AOI21_X2 port map( A1 => n12798, A2 => n10452, B => n10451, ZN => 
                           n15236);
   U18846 : XOR2_X1 port map( A1 => n28121, A2 => n30685, Z => n3106);
   U18851 : XOR2_X1 port map( A1 => n10081, A2 => n29205, Z => n30685);
   U18853 : NOR2_X2 port map( A1 => n10828, A2 => n1377, ZN => n19309);
   U18854 : INV_X2 port map( I => n19308, ZN => n1377);
   U18866 : NOR3_X1 port map( A1 => n33722, A2 => n23813, A3 => n8166, ZN => 
                           n30687);
   U18898 : XOR2_X1 port map( A1 => n7677, A2 => n19712, Z => n9517);
   U18901 : NAND3_X2 port map( A1 => n2585, A2 => n8672, A3 => n2587, ZN => 
                           n19712);
   U18902 : XOR2_X1 port map( A1 => n23270, A2 => n23269, Z => n31034);
   U18904 : INV_X2 port map( I => n12287, ZN => n13720);
   U18912 : XOR2_X1 port map( A1 => n47, A2 => n12288, Z => n12287);
   U18916 : NAND2_X2 port map( A1 => n21804, A2 => n11231, ZN => n115);
   U18922 : NAND2_X2 port map( A1 => n12711, A2 => n12712, ZN => n21804);
   U18923 : INV_X2 port map( I => n30690, ZN => n31911);
   U18931 : NAND3_X2 port map( A1 => n21119, A2 => n7913, A3 => n21118, ZN => 
                           n30690);
   U18933 : XOR2_X1 port map( A1 => n30691, A2 => n9911, Z => n31839);
   U18935 : XOR2_X1 port map( A1 => n11271, A2 => n22287, Z => n30691);
   U18938 : OAI21_X2 port map( A1 => n30693, A2 => n30692, B => n16789, ZN => 
                           n30923);
   U18940 : XOR2_X1 port map( A1 => n23297, A2 => n1825, Z => n23119);
   U18950 : AND2_X1 port map( A1 => n3251, A2 => n31012, Z => n14314);
   U18951 : NAND2_X2 port map( A1 => n2186, A2 => n30695, ZN => n2864);
   U18963 : XOR2_X1 port map( A1 => n7256, A2 => n30540, Z => n24540);
   U18970 : OAI21_X2 port map( A1 => n30698, A2 => n30697, B => n31012, ZN => 
                           n12977);
   U18972 : OAI21_X2 port map( A1 => n30700, A2 => n30699, B => n13968, ZN => 
                           n14983);
   U18979 : NOR2_X1 port map( A1 => n3042, A2 => n31201, ZN => n3045);
   U18981 : XOR2_X1 port map( A1 => n6792, A2 => n30702, Z => n7368);
   U18982 : XOR2_X1 port map( A1 => n7870, A2 => n13181, Z => n30702);
   U19002 : NAND2_X2 port map( A1 => n16552, A2 => n24056, ZN => n26374);
   U19004 : NAND2_X2 port map( A1 => n4483, A2 => n4481, ZN => n24056);
   U19009 : NAND2_X2 port map( A1 => n8482, A2 => n18294, ZN => n27921);
   U19010 : XNOR2_X1 port map( A1 => n2304, A2 => n21022, ZN => n30849);
   U19019 : XOR2_X1 port map( A1 => n23467, A2 => n9185, Z => n16200);
   U19020 : XOR2_X1 port map( A1 => n11862, A2 => n22205, Z => n22153);
   U19022 : OAI22_X2 port map( A1 => n10493, A2 => n28729, B1 => n5495, B2 => 
                           n10492, ZN => n22205);
   U19028 : AOI21_X2 port map( A1 => n6505, A2 => n30703, B => n9777, ZN => 
                           n5035);
   U19036 : NAND2_X2 port map( A1 => n30748, A2 => n28857, ZN => n30705);
   U19042 : XOR2_X1 port map( A1 => n20810, A2 => n20809, Z => n30706);
   U19046 : XOR2_X1 port map( A1 => n29140, A2 => n30707, Z => n1642);
   U19049 : XOR2_X1 port map( A1 => n3295, A2 => n9468, Z => n30707);
   U19052 : XOR2_X1 port map( A1 => n22154, A2 => n7685, Z => n7684);
   U19061 : NAND2_X1 port map( A1 => n3343, A2 => n743, ZN => n30710);
   U19062 : OR2_X2 port map( A1 => n7, A2 => n21970, Z => n22488);
   U19064 : XOR2_X1 port map( A1 => n8809, A2 => n30711, Z => n8806);
   U19069 : XOR2_X1 port map( A1 => n31138, A2 => n30712, Z => n30711);
   U19071 : INV_X2 port map( I => n30713, ZN => n21412);
   U19073 : XOR2_X1 port map( A1 => n22008, A2 => n30714, Z => n27160);
   U19076 : XOR2_X1 port map( A1 => n22288, A2 => n22006, Z => n30714);
   U19083 : NOR2_X2 port map( A1 => n30716, A2 => n17016, ZN => n30732);
   U19088 : NAND2_X2 port map( A1 => n24047, A2 => n8567, ZN => n30716);
   U19089 : OR2_X1 port map( A1 => n9073, A2 => n21428, Z => n17415);
   U19091 : NOR3_X2 port map( A1 => n6414, A2 => n14975, A3 => n14974, ZN => 
                           n30717);
   U19092 : AOI21_X1 port map( A1 => n1284, A2 => n6976, B => n30718, ZN => 
                           n2348);
   U19096 : INV_X2 port map( I => n980, ZN => n30720);
   U19104 : XOR2_X1 port map( A1 => n13208, A2 => n30721, Z => n21432);
   U19105 : XOR2_X1 port map( A1 => n20967, A2 => n30722, Z => n30721);
   U19106 : AOI21_X2 port map( A1 => n29398, A2 => n15505, B => n30760, ZN => 
                           n19273);
   U19107 : XOR2_X1 port map( A1 => n30723, A2 => n19687, Z => n5837);
   U19109 : XOR2_X1 port map( A1 => n5236, A2 => n19430, Z => n30723);
   U19110 : NOR3_X2 port map( A1 => n17211, A2 => n28214, A3 => n22705, ZN => 
                           n30724);
   U19112 : NAND2_X1 port map( A1 => n23640, A2 => n14078, ZN => n30725);
   U19118 : NAND2_X2 port map( A1 => n30931, A2 => n16684, ZN => n27317);
   U19121 : BUF_X2 port map( I => n31040, Z => n30727);
   U19127 : OR2_X1 port map( A1 => n32051, A2 => n5225, Z => n18352);
   U19146 : OAI22_X2 port map( A1 => n9741, A2 => n9740, B1 => n5764, B2 => 
                           n23788, ZN => n7581);
   U19158 : NAND3_X2 port map( A1 => n7324, A2 => n21519, A3 => n7323, ZN => 
                           n22028);
   U19168 : XOR2_X1 port map( A1 => n14742, A2 => n19503, Z => n17434);
   U19177 : BUF_X2 port map( I => n31882, Z => n30729);
   U19181 : NAND2_X2 port map( A1 => n15123, A2 => n6605, ZN => n22946);
   U19185 : OAI22_X2 port map( A1 => n12601, A2 => n28705, B1 => n12131, B2 => 
                           n12600, ZN => n19370);
   U19187 : INV_X1 port map( I => n30730, ZN => n8631);
   U19198 : NAND2_X2 port map( A1 => n31223, A2 => n6667, ZN => n339);
   U19199 : OAI21_X2 port map( A1 => n2409, A2 => n2408, B => n2407, ZN => 
                           n13762);
   U19206 : NAND2_X2 port map( A1 => n7798, A2 => n14945, ZN => n17837);
   U19208 : XOR2_X1 port map( A1 => n22085, A2 => n6462, Z => n17377);
   U19213 : AND2_X1 port map( A1 => n632, A2 => n10681, Z => n15763);
   U19216 : NAND3_X2 port map( A1 => n31963, A2 => n29078, A3 => n123, ZN => 
                           n26324);
   U19217 : AND2_X1 port map( A1 => n23843, A2 => n299, Z => n14088);
   U19220 : NAND2_X1 port map( A1 => n20339, A2 => n15169, ZN => n15042);
   U19238 : NAND2_X2 port map( A1 => n11090, A2 => n3405, ZN => n25565);
   U19250 : XOR2_X1 port map( A1 => n23342, A2 => n30733, Z => n23136);
   U19251 : NOR2_X1 port map( A1 => n1348, A2 => n19402, ZN => n26358);
   U19256 : XOR2_X1 port map( A1 => n30734, A2 => n31321, Z => n14726);
   U19266 : OAI21_X2 port map( A1 => n30737, A2 => n30736, B => n23864, ZN => 
                           n17183);
   U19288 : NOR2_X2 port map( A1 => n19023, A2 => n19020, ZN => n27726);
   U19292 : AOI21_X2 port map( A1 => n3429, A2 => n732, B => n2682, ZN => 
                           n19023);
   U19293 : XOR2_X1 port map( A1 => n9848, A2 => n24567, Z => n8575);
   U19298 : NOR2_X2 port map( A1 => n23404, A2 => n30741, ZN => n5505);
   U19299 : XOR2_X1 port map( A1 => n30742, A2 => n25880, Z => Ciphertext(182))
                           ;
   U19303 : OAI22_X1 port map( A1 => n5303, A2 => n25995, B1 => n5301, B2 => 
                           n5300, ZN => n30742);
   U19311 : XOR2_X1 port map( A1 => n30746, A2 => n16555, Z => Ciphertext(103))
                           ;
   U19321 : AND2_X1 port map( A1 => n3911, A2 => n22420, Z => n30758);
   U19334 : NAND3_X1 port map( A1 => n17087, A2 => n23764, A3 => n1101, ZN => 
                           n17088);
   U19340 : XOR2_X1 port map( A1 => n11062, A2 => n15297, Z => n1941);
   U19341 : NAND2_X1 port map( A1 => n7486, A2 => n28166, ZN => n20553);
   U19344 : AOI21_X2 port map( A1 => n27372, A2 => n29317, B => n30753, ZN => 
                           n26656);
   U19345 : NAND2_X2 port map( A1 => n30754, A2 => n28956, ZN => n24289);
   U19356 : INV_X2 port map( I => n12945, ZN => n1231);
   U19358 : NAND2_X2 port map( A1 => n7246, A2 => n27480, ZN => n12945);
   U19367 : XOR2_X1 port map( A1 => n30757, A2 => n19417, Z => n11591);
   U19372 : NOR2_X2 port map( A1 => n29156, A2 => n19884, ZN => n13840);
   U19377 : XOR2_X1 port map( A1 => n11545, A2 => n11543, Z => n20152);
   U19378 : BUF_X2 port map( I => n19268, Z => n30760);
   U19411 : XOR2_X1 port map( A1 => n112, A2 => n30766, Z => n30765);
   U19420 : XOR2_X1 port map( A1 => n15424, A2 => n23411, Z => n30767);
   U19428 : XOR2_X1 port map( A1 => n20753, A2 => n15557, Z => n15556);
   U19434 : OAI22_X1 port map( A1 => n19079, A2 => n34005, B1 => n19080, B2 => 
                           n948, ZN => n30768);
   U19437 : NAND3_X1 port map( A1 => n13286, A2 => n17624, A3 => n21338, ZN => 
                           n2242);
   U19441 : NAND2_X2 port map( A1 => n8489, A2 => n14326, ZN => n31254);
   U19444 : INV_X2 port map( I => n30770, ZN => n14458);
   U19464 : XOR2_X1 port map( A1 => n19736, A2 => n19654, Z => n7887);
   U19468 : NAND2_X2 port map( A1 => n10532, A2 => n4098, ZN => n11231);
   U19472 : XOR2_X1 port map( A1 => n5146, A2 => n30776, Z => n31747);
   U19473 : XOR2_X1 port map( A1 => n24741, A2 => n16381, Z => n30776);
   U19474 : XOR2_X1 port map( A1 => n30777, A2 => n24895, Z => Ciphertext(47));
   U19477 : XOR2_X1 port map( A1 => n1938, A2 => n1935, Z => n9870);
   U19480 : OR2_X2 port map( A1 => n26345, A2 => n4740, Z => n21173);
   U19483 : NAND2_X2 port map( A1 => n30780, A2 => n31694, ZN => n16804);
   U19485 : OAI22_X2 port map( A1 => n4142, A2 => n16812, B1 => n20044, B2 => 
                           n20045, ZN => n30780);
   U19510 : XOR2_X1 port map( A1 => n21996, A2 => n8356, Z => n15726);
   U19525 : XOR2_X1 port map( A1 => n11304, A2 => n20773, Z => n28621);
   U19528 : INV_X2 port map( I => n14383, ZN => n21358);
   U19535 : XOR2_X1 port map( A1 => n3010, A2 => n11530, Z => n14383);
   U19540 : NAND2_X2 port map( A1 => n31036, A2 => n10297, ZN => n19743);
   U19542 : NAND2_X1 port map( A1 => n1734, A2 => n1733, ZN => n30792);
   U19548 : XOR2_X1 port map( A1 => n22252, A2 => n21919, Z => n7686);
   U19550 : NAND2_X2 port map( A1 => n20089, A2 => n5405, ZN => n2271);
   U19551 : NAND2_X2 port map( A1 => n31046, A2 => n1161, ZN => n20089);
   U19558 : NAND4_X2 port map( A1 => n17756, A2 => n12758, A3 => n2619, A4 => 
                           n2618, ZN => n30942);
   U19565 : NAND3_X2 port map( A1 => n5581, A2 => n9597, A3 => n20407, ZN => 
                           n8728);
   U19570 : AND2_X1 port map( A1 => n30293, A2 => n29313, Z => n7529);
   U19592 : NAND2_X1 port map( A1 => n654, A2 => n23899, ZN => n23628);
   U19594 : NOR2_X2 port map( A1 => n31399, A2 => n30800, ZN => n1260);
   U19617 : XOR2_X1 port map( A1 => n30532, A2 => n17871, Z => n13661);
   U19623 : XOR2_X1 port map( A1 => n30807, A2 => n16002, Z => n4574);
   U19627 : XOR2_X1 port map( A1 => n30808, A2 => n25849, Z => Ciphertext(176))
                           ;
   U19631 : NAND2_X2 port map( A1 => n8628, A2 => n30810, ZN => n16748);
   U19632 : AOI22_X1 port map( A1 => n8627, A2 => n11123, B1 => n18541, B2 => 
                           n31821, ZN => n30810);
   U19646 : NOR2_X2 port map( A1 => n743, A2 => n11302, ZN => n5034);
   U19652 : INV_X1 port map( I => n31180, ZN => n5056);
   U19655 : AOI21_X1 port map( A1 => n12486, A2 => n28658, B => n31206, ZN => 
                           n31214);
   U19656 : XOR2_X1 port map( A1 => n8750, A2 => n29347, Z => n30815);
   U19658 : AND2_X1 port map( A1 => n25429, A2 => n17948, Z => n31142);
   U19667 : NAND2_X1 port map( A1 => n28353, A2 => n31563, ZN => n14394);
   U19676 : XOR2_X1 port map( A1 => n33509, A2 => n23239, Z => n31191);
   U19679 : NOR2_X1 port map( A1 => n28915, A2 => n8314, ZN => n26660);
   U19684 : INV_X2 port map( I => n22602, ZN => n8314);
   U19688 : XOR2_X1 port map( A1 => n15727, A2 => n26487, Z => n22602);
   U19701 : XOR2_X1 port map( A1 => n2375, A2 => n30818, Z => n31495);
   U19702 : XOR2_X1 port map( A1 => n30819, A2 => n11889, Z => n30818);
   U19706 : INV_X2 port map( I => n30820, ZN => n23807);
   U19707 : XOR2_X1 port map( A1 => n7616, A2 => n7614, Z => n30820);
   U19725 : OAI22_X2 port map( A1 => n14678, A2 => n18424, B1 => n17102, B2 => 
                           n14117, ZN => n19158);
   U19728 : XOR2_X1 port map( A1 => n30822, A2 => n15765, Z => n3987);
   U19746 : AND2_X1 port map( A1 => n7251, A2 => n4656, Z => n2646);
   U19751 : XOR2_X1 port map( A1 => n21036, A2 => n20842, Z => n11578);
   U19756 : NOR2_X2 port map( A1 => n12514, A2 => n20742, ZN => n21036);
   U19766 : AOI21_X1 port map( A1 => n19128, A2 => n7968, B => n31177, ZN => 
                           n12268);
   U19772 : NAND2_X2 port map( A1 => n79, A2 => n31942, ZN => n22831);
   U19776 : NOR2_X2 port map( A1 => n27455, A2 => n11922, ZN => n23646);
   U19788 : AND3_X1 port map( A1 => n23730, A2 => n23938, A3 => n12469, Z => 
                           n31028);
   U19794 : AOI21_X1 port map( A1 => n30828, A2 => n27265, B => n17181, ZN => 
                           n17178);
   U19816 : NOR2_X1 port map( A1 => n30326, A2 => n11394, ZN => n21123);
   U19823 : XOR2_X1 port map( A1 => n30830, A2 => n15307, Z => n23683);
   U19825 : XOR2_X1 port map( A1 => n23513, A2 => n23514, Z => n30830);
   U19828 : INV_X4 port map( I => n7552, ZN => n14005);
   U19832 : INV_X2 port map( I => n14851, ZN => n22238);
   U19833 : NAND2_X2 port map( A1 => n21765, A2 => n21764, ZN => n14851);
   U19848 : XOR2_X1 port map( A1 => n30837, A2 => n16655, Z => Ciphertext(19));
   U19857 : XOR2_X1 port map( A1 => n30840, A2 => n25648, Z => Ciphertext(140))
                           ;
   U19860 : AOI22_X1 port map( A1 => n26745, A2 => n25646, B1 => n25660, B2 => 
                           n25645, ZN => n30840);
   U19870 : XOR2_X1 port map( A1 => n24645, A2 => n4244, Z => n24482);
   U19886 : NAND2_X1 port map( A1 => n24977, A2 => n17684, ZN => n24892);
   U19891 : NOR2_X2 port map( A1 => n15169, A2 => n15043, ZN => n28504);
   U19894 : XOR2_X1 port map( A1 => n7772, A2 => n30843, Z => n9018);
   U19899 : BUF_X4 port map( I => n14396, Z => n30885);
   U19900 : AND2_X1 port map( A1 => n27748, A2 => n29688, Z => n13083);
   U19912 : XOR2_X1 port map( A1 => n30844, A2 => n7570, Z => n14702);
   U19917 : XOR2_X1 port map( A1 => n10169, A2 => n7569, Z => n30844);
   U19928 : XOR2_X1 port map( A1 => n33492, A2 => n24620, Z => n24766);
   U19932 : XOR2_X1 port map( A1 => n20692, A2 => n20769, Z => n11304);
   U19945 : XOR2_X1 port map( A1 => n30850, A2 => n5067, Z => n1487);
   U19949 : XOR2_X1 port map( A1 => n5100, A2 => n8997, Z => n30850);
   U19982 : NAND2_X2 port map( A1 => n27391, A2 => n6716, ZN => n6713);
   U19989 : XOR2_X1 port map( A1 => n15630, A2 => n5647, Z => n4672);
   U20005 : NAND2_X2 port map( A1 => n2997, A2 => n30855, ZN => n3229);
   U20006 : NOR2_X2 port map( A1 => n2996, A2 => n28519, ZN => n30855);
   U20014 : OAI21_X2 port map( A1 => n13083, A2 => n33714, B => n13157, ZN => 
                           n30857);
   U20038 : XOR2_X1 port map( A1 => n10539, A2 => n24846, Z => n24597);
   U20039 : OAI21_X2 port map( A1 => n2851, A2 => n2849, B => n2848, ZN => 
                           n24846);
   U20065 : XOR2_X1 port map( A1 => n9526, A2 => n19491, Z => n3980);
   U20066 : NAND2_X1 port map( A1 => n12270, A2 => n18983, ZN => n31177);
   U20074 : INV_X2 port map( I => n30861, ZN => n17522);
   U20075 : OAI21_X1 port map( A1 => n30863, A2 => n30862, B => n21368, ZN => 
                           n26504);
   U20087 : NOR2_X1 port map( A1 => n21367, A2 => n21391, ZN => n30862);
   U20090 : NAND2_X2 port map( A1 => n30957, A2 => n30959, ZN => n19245);
   U20091 : NAND3_X1 port map( A1 => n25121, A2 => n2092, A3 => n25120, ZN => 
                           n13667);
   U20093 : AOI22_X1 port map( A1 => n11518, A2 => n2209, B1 => n2208, B2 => 
                           n25670, ZN => n6469);
   U20095 : NAND2_X1 port map( A1 => n146, A2 => n9195, ZN => n30867);
   U20097 : NAND2_X1 port map( A1 => n30933, A2 => n30932, ZN => n31150);
   U20112 : NOR2_X2 port map( A1 => n30869, A2 => n29603, ZN => n15591);
   U20113 : NOR2_X2 port map( A1 => n9560, A2 => n6958, ZN => n31136);
   U20117 : NAND2_X2 port map( A1 => n8015, A2 => n8016, ZN => n2387);
   U20120 : XOR2_X1 port map( A1 => n23471, A2 => n23356, Z => n15712);
   U20124 : XOR2_X1 port map( A1 => n6886, A2 => n30871, Z => n16277);
   U20125 : XOR2_X1 port map( A1 => n16912, A2 => n16910, Z => n30871);
   U20126 : XOR2_X1 port map( A1 => n1261, A2 => n12491, Z => n9222);
   U20133 : NAND2_X1 port map( A1 => n30872, A2 => n16699, ZN => n8437);
   U20137 : NAND2_X1 port map( A1 => n19335, A2 => n2207, ZN => n30872);
   U20146 : OR2_X1 port map( A1 => n31532, A2 => n20471, Z => n30873);
   U20154 : NAND3_X2 port map( A1 => n5222, A2 => n5221, A3 => n12755, ZN => 
                           n19627);
   U20158 : INV_X2 port map( I => n13530, ZN => n24209);
   U20162 : XOR2_X1 port map( A1 => n15825, A2 => n22226, Z => n12495);
   U20174 : XNOR2_X1 port map( A1 => n10539, A2 => n24760, ZN => n24576);
   U20181 : NOR2_X1 port map( A1 => n10542, A2 => n30980, ZN => n30979);
   U20183 : NAND2_X1 port map( A1 => n29367, A2 => n30979, ZN => n3840);
   U20184 : NAND2_X1 port map( A1 => n20602, A2 => n15230, ZN => n20601);
   U20187 : OAI22_X2 port map( A1 => n21839, A2 => n21840, B1 => n13816, B2 => 
                           n21844, ZN => n14594);
   U20192 : XOR2_X1 port map( A1 => n14969, A2 => n22300, Z => n22008);
   U20201 : XOR2_X1 port map( A1 => n20799, A2 => n30880, Z => n31841);
   U20203 : XOR2_X1 port map( A1 => n20921, A2 => n30881, Z => n30880);
   U20204 : XOR2_X1 port map( A1 => n31043, A2 => n21018, Z => n2304);
   U20211 : NAND2_X2 port map( A1 => n27646, A2 => n5103, ZN => n31043);
   U20222 : NAND2_X2 port map( A1 => n31967, A2 => n28840, ZN => n11103);
   U20228 : INV_X2 port map( I => n2347, ZN => n5379);
   U20230 : XOR2_X1 port map( A1 => n29057, A2 => n616, Z => n2347);
   U20261 : XOR2_X1 port map( A1 => n17546, A2 => n30887, Z => n31875);
   U20262 : XOR2_X1 port map( A1 => n5211, A2 => n27613, Z => n30887);
   U20269 : AOI21_X2 port map( A1 => n10468, A2 => n30889, B => n32816, ZN => 
                           n9071);
   U20278 : NAND2_X2 port map( A1 => n327, A2 => n16334, ZN => n6649);
   U20280 : INV_X1 port map( I => n1694, ZN => n19771);
   U20294 : OR2_X1 port map( A1 => n26040, A2 => n3601, Z => n13087);
   U20298 : OR2_X1 port map( A1 => n20322, A2 => n20379, Z => n30892);
   U20311 : OR2_X1 port map( A1 => n20008, A2 => n20080, Z => n13771);
   U20312 : NAND2_X2 port map( A1 => n17183, A2 => n30898, ZN => n1931);
   U20318 : XOR2_X1 port map( A1 => n19662, A2 => n13099, Z => n30899);
   U20321 : XOR2_X1 port map( A1 => n30900, A2 => n13689, Z => n14621);
   U20323 : XOR2_X1 port map( A1 => n26794, A2 => n30993, Z => n30900);
   U20325 : XOR2_X1 port map( A1 => n22016, A2 => n4739, Z => n30901);
   U20334 : AOI21_X2 port map( A1 => n867, A2 => n10488, B => n31135, ZN => 
                           n10486);
   U20339 : XOR2_X1 port map( A1 => n2117, A2 => n25783, Z => n4567);
   U20340 : NAND2_X2 port map( A1 => n31297, A2 => n31872, ZN => n2117);
   U20363 : XOR2_X1 port map( A1 => n30749, A2 => n16690, Z => n26929);
   U20365 : INV_X2 port map( I => n30905, ZN => n20092);
   U20368 : BUF_X2 port map( I => n8392, Z => n30906);
   U20378 : XOR2_X1 port map( A1 => n13132, A2 => n13131, Z => n15401);
   U20399 : OAI21_X2 port map( A1 => n30914, A2 => n30913, B => n728, ZN => 
                           n28821);
   U20405 : INV_X2 port map( I => n21433, ZN => n30914);
   U20406 : NOR2_X1 port map( A1 => n31207, A2 => n25072, ZN => n5864);
   U20407 : NAND2_X1 port map( A1 => n33288, A2 => n5003, ZN => n30915);
   U20412 : NAND2_X1 port map( A1 => n11195, A2 => n858, ZN => n30989);
   U20423 : OR2_X1 port map( A1 => n25072, A2 => n32900, Z => n28655);
   U20437 : AOI21_X2 port map( A1 => n29394, A2 => n30727, B => n2941, ZN => 
                           n10769);
   U20440 : NAND3_X2 port map( A1 => n30919, A2 => n27618, A3 => n3149, ZN => 
                           n3093);
   U20454 : NAND2_X2 port map( A1 => n25966, A2 => n11988, ZN => n13353);
   U20464 : NAND3_X1 port map( A1 => n28734, A2 => n25312, A3 => n25322, ZN => 
                           n17105);
   U20481 : NAND2_X2 port map( A1 => n23679, A2 => n23680, ZN => n24652);
   U20482 : XOR2_X1 port map( A1 => n3322, A2 => n3319, Z => n3318);
   U20483 : XOR2_X1 port map( A1 => n27176, A2 => n23295, Z => n3322);
   U20485 : NOR2_X2 port map( A1 => n2272, A2 => n31215, ZN => n30978);
   U20490 : NAND2_X2 port map( A1 => n10769, A2 => n2719, ZN => n21816);
   U20508 : INV_X2 port map( I => n30926, ZN => n22425);
   U20509 : XOR2_X1 port map( A1 => n16000, A2 => n15999, Z => n30926);
   U20521 : XNOR2_X1 port map( A1 => n12442, A2 => n29030, ZN => n19584);
   U20529 : AOI22_X2 port map( A1 => n23962, A2 => n28410, B1 => n24046, B2 => 
                           n3506, ZN => n3508);
   U20538 : NAND2_X2 port map( A1 => n25442, A2 => n25439, ZN => n25437);
   U20563 : OAI21_X2 port map( A1 => n739, A2 => n23887, B => n23841, ZN => 
                           n8689);
   U20575 : NOR2_X2 port map( A1 => n11742, A2 => n13732, ZN => n16141);
   U20587 : NAND2_X2 port map( A1 => n21532, A2 => n30389, ZN => n17274);
   U20592 : XOR2_X1 port map( A1 => n21951, A2 => n16036, Z => n13436);
   U20606 : OR2_X1 port map( A1 => n12974, A2 => n23843, Z => n7524);
   U20612 : XOR2_X1 port map( A1 => n30380, A2 => n23233, Z => n23384);
   U20619 : NAND2_X2 port map( A1 => n11162, A2 => n23089, ZN => n23233);
   U20629 : NAND2_X2 port map( A1 => n27793, A2 => n23550, ZN => n24403);
   U20631 : NAND3_X1 port map( A1 => n24325, A2 => n24327, A3 => n29141, ZN => 
                           n24080);
   U20650 : AOI21_X2 port map( A1 => n30948, A2 => n25121, B => n25025, ZN => 
                           n16469);
   U20660 : AOI22_X2 port map( A1 => n15902, A2 => n8184, B1 => n16538, B2 => 
                           n18407, ZN => n27953);
   U20661 : OAI21_X2 port map( A1 => n13839, A2 => n22967, B => n13837, ZN => 
                           n23475);
   U20667 : NOR2_X2 port map( A1 => n9959, A2 => n10258, ZN => n9958);
   U20670 : XOR2_X1 port map( A1 => n26054, A2 => n22268, Z => n30951);
   U20690 : OR2_X1 port map( A1 => n16226, A2 => n20657, Z => n20662);
   U20691 : NAND2_X2 port map( A1 => n5448, A2 => n22806, ZN => n26724);
   U20697 : AOI22_X2 port map( A1 => n4931, A2 => n4932, B1 => n4930, B2 => 
                           n33904, ZN => n30953);
   U20699 : XOR2_X1 port map( A1 => n20955, A2 => n30954, Z => n587);
   U20703 : NAND2_X2 port map( A1 => n13276, A2 => n13275, ZN => n7229);
   U20707 : XOR2_X1 port map( A1 => n17400, A2 => n30955, Z => n28818);
   U20720 : NOR2_X2 port map( A1 => n31949, A2 => n30958, ZN => n30957);
   U20722 : INV_X2 port map( I => n18876, ZN => n30959);
   U20724 : OR2_X2 port map( A1 => n15721, A2 => n7865, Z => n4602);
   U20746 : XOR2_X1 port map( A1 => n12936, A2 => n12935, Z => n24360);
   U20750 : XOR2_X1 port map( A1 => n30964, A2 => n23188, Z => n10772);
   U20774 : XOR2_X1 port map( A1 => n24841, A2 => n26121, Z => n29072);
   U20782 : XOR2_X1 port map( A1 => n11651, A2 => n1084, Z => n24841);
   U20783 : OAI21_X1 port map( A1 => n30971, A2 => n20635, B => n30970, ZN => 
                           n1811);
   U20785 : NAND2_X1 port map( A1 => n15569, A2 => n3994, ZN => n7786);
   U20786 : OR2_X1 port map( A1 => n28702, A2 => n30973, Z => n5836);
   U20814 : INV_X2 port map( I => n843, ZN => n30980);
   U20815 : XOR2_X1 port map( A1 => n30981, A2 => n29467, Z => n31140);
   U20827 : XOR2_X1 port map( A1 => n16992, A2 => n13702, Z => n30981);
   U20831 : NOR2_X2 port map( A1 => n27555, A2 => n10030, ZN => n30982);
   U20832 : XOR2_X1 port map( A1 => n30985, A2 => n20719, Z => n26401);
   U20851 : XOR2_X1 port map( A1 => n5296, A2 => n6050, Z => n30986);
   U20860 : NOR2_X1 port map( A1 => n18098, A2 => n22394, ZN => n31144);
   U20861 : XOR2_X1 port map( A1 => n20757, A2 => n5210, Z => n5209);
   U20870 : XOR2_X1 port map( A1 => n23282, A2 => n32899, Z => n15432);
   U20871 : NAND2_X2 port map( A1 => n16630, A2 => n16789, ZN => n10413);
   U20877 : XOR2_X1 port map( A1 => n2192, A2 => n30992, Z => n509);
   U20887 : XOR2_X1 port map( A1 => n31477, A2 => n30993, Z => n30992);
   U20895 : INV_X2 port map( I => n30994, ZN => n9170);
   U20906 : NAND2_X2 port map( A1 => n29525, A2 => n13925, ZN => n18922);
   U20932 : XOR2_X1 port map( A1 => n1781, A2 => n1778, Z => n17683);
   U20940 : BUF_X2 port map( I => n22634, Z => n31001);
   U20941 : XOR2_X1 port map( A1 => n7646, A2 => n7644, Z => n12804);
   U20945 : NAND2_X2 port map( A1 => n29088, A2 => n424, ZN => n9439);
   U20948 : NAND3_X1 port map( A1 => n5494, A2 => n30832, A3 => n21872, ZN => 
                           n12604);
   U20952 : AND2_X1 port map( A1 => n22421, A2 => n22420, Z => n31006);
   U20967 : AOI21_X1 port map( A1 => n18822, A2 => n18701, B => n31012, ZN => 
                           n16395);
   U20969 : NAND2_X2 port map( A1 => n23663, A2 => n31015, ZN => n24632);
   U20971 : NOR2_X2 port map( A1 => n16442, A2 => n10899, ZN => n25893);
   U20974 : INV_X2 port map( I => n24096, ZN => n17404);
   U20979 : OAI21_X2 port map( A1 => n28303, A2 => n17490, B => n23649, ZN => 
                           n24096);
   U20996 : XOR2_X1 port map( A1 => n4059, A2 => n6707, Z => n6705);
   U21004 : INV_X4 port map( I => n26157, ZN => n3748);
   U21019 : NOR2_X1 port map( A1 => n19165, A2 => n4835, ZN => n31029);
   U21025 : INV_X2 port map( I => n27933, ZN => n468);
   U21026 : XOR2_X1 port map( A1 => n19642, A2 => n19163, Z => n6624);
   U21032 : AOI22_X2 port map( A1 => n31781, A2 => n21846, B1 => n21518, B2 => 
                           n7969, ZN => n31032);
   U21033 : XOR2_X1 port map( A1 => n15433, A2 => n15430, Z => n15514);
   U21041 : AND2_X1 port map( A1 => n16686, A2 => n29268, Z => n31524);
   U21048 : INV_X2 port map( I => n31034, ZN => n9828);
   U21049 : XOR2_X1 port map( A1 => n23516, A2 => n23254, Z => n9865);
   U21056 : OAI21_X2 port map( A1 => n12160, A2 => n2886, B => n12159, ZN => 
                           n31037);
   U21063 : NOR2_X2 port map( A1 => n29397, A2 => n7105, ZN => n31039);
   U21065 : OAI21_X1 port map( A1 => n9285, A2 => n31042, B => n31041, ZN => 
                           n11646);
   U21067 : INV_X2 port map( I => n31044, ZN => n20120);
   U21069 : XOR2_X1 port map( A1 => n19640, A2 => n14574, Z => n31044);
   U21076 : NOR2_X2 port map( A1 => n18658, A2 => n18657, ZN => n27807);
   U21079 : INV_X2 port map( I => n20011, ZN => n31046);
   U21088 : AND2_X1 port map( A1 => n5415, A2 => n819, Z => n31047);
   U21112 : XOR2_X1 port map( A1 => n7288, A2 => n34050, Z => n27699);
   U21114 : OAI22_X2 port map( A1 => n18344, A2 => n26181, B1 => n19052, B2 => 
                           n10015, ZN => n18345);
   U21147 : XOR2_X1 port map( A1 => n8113, A2 => n8110, Z => n18080);
   U21151 : NAND2_X1 port map( A1 => n17277, A2 => n13950, ZN => n24107);
   U21167 : NAND2_X1 port map( A1 => n25876, A2 => n25875, ZN => n25877);
   U21174 : OAI22_X1 port map( A1 => n22329, A2 => n1000, B1 => n22406, B2 => 
                           n30529, ZN => n13071);
   U21181 : XOR2_X1 port map( A1 => n5380, A2 => n31056, Z => n31055);
   U21187 : NAND2_X2 port map( A1 => n1146, A2 => n16639, ZN => n21433);
   U21195 : OAI22_X2 port map( A1 => n18841, A2 => n18840, B1 => n2148, B2 => 
                           n1181, ZN => n31882);
   U21198 : NOR2_X1 port map( A1 => n963, A2 => n14940, ZN => n6043);
   U21200 : NOR2_X1 port map( A1 => n18944, A2 => n7345, ZN => n8573);
   U21202 : INV_X2 port map( I => n25313, ZN => n1074);
   U21217 : NAND2_X2 port map( A1 => n25293, A2 => n25294, ZN => n25313);
   U21219 : AND2_X1 port map( A1 => n22523, A2 => n22605, Z => n29027);
   U21223 : XOR2_X1 port map( A1 => n31059, A2 => n20835, Z => n20895);
   U21224 : AOI21_X2 port map( A1 => n5413, A2 => n5416, B => n31976, ZN => 
                           n5414);
   U21236 : XOR2_X1 port map( A1 => n31731, A2 => n25457, Z => n19693);
   U21238 : NAND2_X2 port map( A1 => n16106, A2 => n19155, ZN => n31731);
   U21246 : XNOR2_X1 port map( A1 => n24646, A2 => n24231, ZN => n31312);
   U21254 : NAND2_X2 port map( A1 => n13985, A2 => n25302, ZN => n31060);
   U21260 : NAND2_X2 port map( A1 => n13768, A2 => n20556, ZN => n20520);
   U21263 : XOR2_X1 port map( A1 => n9135, A2 => n9136, Z => n10197);
   U21266 : XOR2_X1 port map( A1 => n8152, A2 => n24452, Z => n28896);
   U21267 : XOR2_X1 port map( A1 => n12283, A2 => n19737, Z => n2750);
   U21281 : NAND2_X2 port map( A1 => n21312, A2 => n21448, ZN => n21314);
   U21288 : NOR2_X2 port map( A1 => n17699, A2 => n16633, ZN => n21312);
   U21289 : XOR2_X1 port map( A1 => n18091, A2 => n31063, Z => n10944);
   U21290 : XOR2_X1 port map( A1 => n10084, A2 => n1423, Z => n31063);
   U21296 : XOR2_X1 port map( A1 => n31065, A2 => n25598, Z => Ciphertext(132))
                           ;
   U21297 : NAND2_X2 port map( A1 => n19031, A2 => n31066, ZN => n7971);
   U21305 : XOR2_X1 port map( A1 => n3235, A2 => n3233, Z => n24503);
   U21321 : NAND2_X1 port map( A1 => n26891, A2 => n27965, ZN => n2970);
   U21322 : NAND2_X1 port map( A1 => n23706, A2 => n499, ZN => n15266);
   U21326 : XOR2_X1 port map( A1 => n31070, A2 => n6086, Z => n8074);
   U21330 : INV_X2 port map( I => n24091, ZN => n10198);
   U21338 : NAND2_X2 port map( A1 => n1035, A2 => n19990, ZN => n13077);
   U21339 : XOR2_X1 port map( A1 => n20850, A2 => n16823, Z => n20853);
   U21341 : XOR2_X1 port map( A1 => n20963, A2 => n20904, Z => n20850);
   U21359 : NAND2_X2 port map( A1 => n919, A2 => n21687, ZN => n21686);
   U21370 : AOI22_X1 port map( A1 => n6043, A2 => n25995, B1 => n30318, B2 => 
                           n3489, ZN => n31075);
   U21386 : NAND2_X2 port map( A1 => n31077, A2 => n9975, ZN => n29157);
   U21387 : OAI21_X2 port map( A1 => n28210, A2 => n14973, B => n23784, ZN => 
                           n31077);
   U21400 : NAND2_X1 port map( A1 => n9485, A2 => n9483, ZN => n31078);
   U21410 : XOR2_X1 port map( A1 => n15438, A2 => n13793, Z => n13792);
   U21411 : OAI21_X2 port map( A1 => n24013, A2 => n10198, B => n24130, ZN => 
                           n7246);
   U21420 : XOR2_X1 port map( A1 => n31151, A2 => n27812, Z => n24883);
   U21422 : XOR2_X1 port map( A1 => n11775, A2 => n14442, Z => n31081);
   U21434 : XOR2_X1 port map( A1 => n4792, A2 => n4790, Z => n4791);
   U21447 : OAI22_X2 port map( A1 => n31086, A2 => n24322, B1 => n7059, B2 => 
                           n24213, ZN => n9468);
   U21448 : XOR2_X1 port map( A1 => n20765, A2 => n20764, Z => n3793);
   U21452 : XOR2_X1 port map( A1 => n31087, A2 => n14202, Z => n28750);
   U21468 : NAND2_X2 port map( A1 => n31091, A2 => n16088, ZN => n19046);
   U21473 : NAND2_X2 port map( A1 => n27709, A2 => n16086, ZN => n31091);
   U21474 : XOR2_X1 port map( A1 => n24569, A2 => n5358, Z => n31092);
   U21476 : INV_X1 port map( I => n23536, ZN => n1258);
   U21478 : XOR2_X1 port map( A1 => n20835, A2 => n17592, Z => n20771);
   U21490 : XOR2_X1 port map( A1 => n24662, A2 => n31093, Z => n12083);
   U21494 : INV_X1 port map( I => n25549, ZN => n31094);
   U21502 : NOR2_X2 port map( A1 => n4017, A2 => n10017, ZN => n19007);
   U21503 : BUF_X4 port map( I => n841, Z => n31096);
   U21507 : NOR2_X1 port map( A1 => n8946, A2 => n1826, ZN => n31097);
   U21510 : XOR2_X1 port map( A1 => n23384, A2 => n531, Z => n12738);
   U21511 : XOR2_X1 port map( A1 => n19463, A2 => n19445, Z => n19642);
   U21537 : INV_X2 port map( I => n31099, ZN => n18623);
   U21544 : AOI21_X1 port map( A1 => n25306, A2 => n18059, B => n692, ZN => 
                           n5792);
   U21567 : XOR2_X1 port map( A1 => n613, A2 => n10186, Z => n31100);
   U21570 : NAND2_X2 port map( A1 => n548, A2 => n32602, ZN => n23866);
   U21572 : INV_X2 port map( I => n31101, ZN => n515);
   U21590 : XOR2_X1 port map( A1 => n31104, A2 => n4427, Z => n31561);
   U21594 : XOR2_X1 port map( A1 => n21995, A2 => n22275, Z => n31104);
   U21620 : INV_X2 port map( I => n11248, ZN => n397);
   U21627 : NOR2_X2 port map( A1 => n31110, A2 => n31109, ZN => n25743);
   U21637 : XOR2_X1 port map( A1 => n19638, A2 => n19639, Z => n14574);
   U21644 : XOR2_X1 port map( A1 => n23286, A2 => n4047, Z => n1795);
   U21648 : NAND2_X2 port map( A1 => n13861, A2 => n17893, ZN => n4047);
   U21653 : OAI21_X2 port map( A1 => n3911, A2 => n18181, B => n9737, ZN => 
                           n28058);
   U21658 : NAND2_X2 port map( A1 => n21799, A2 => n12211, ZN => n21709);
   U21660 : XOR2_X1 port map( A1 => n2747, A2 => n27365, Z => n28430);
   U21664 : INV_X2 port map( I => n31114, ZN => n31909);
   U21668 : XOR2_X1 port map( A1 => n6895, A2 => n26087, Z => n31114);
   U21671 : XOR2_X1 port map( A1 => n1845, A2 => n1844, Z => n31116);
   U21672 : XOR2_X1 port map( A1 => n31117, A2 => n31756, Z => n7672);
   U21674 : XOR2_X1 port map( A1 => n20888, A2 => n5282, Z => n31117);
   U21676 : NAND2_X1 port map( A1 => n4714, A2 => n32619, ZN => n4715);
   U21686 : NOR2_X1 port map( A1 => n2720, A2 => n30129, ZN => n2948);
   U21687 : NOR2_X2 port map( A1 => n27406, A2 => n22479, ZN => n31145);
   U21707 : NOR2_X2 port map( A1 => n31118, A2 => n2178, ZN => n22216);
   U21726 : INV_X1 port map( I => n23052, ZN => n31120);
   U21735 : XOR2_X1 port map( A1 => n26145, A2 => n3318, Z => n31409);
   U21752 : XOR2_X1 port map( A1 => n23530, A2 => n1428, Z => n17353);
   U21760 : AOI21_X2 port map( A1 => n11048, A2 => n10896, B => n31758, ZN => 
                           n23530);
   U21772 : XOR2_X1 port map( A1 => n31123, A2 => n24820, Z => n24821);
   U21774 : XOR2_X1 port map( A1 => n27801, A2 => n24853, Z => n31123);
   U21787 : OAI22_X1 port map( A1 => n9655, A2 => n25194, B1 => n1071, B2 => 
                           n9247, ZN => n4767);
   U21788 : INV_X2 port map( I => n4770, ZN => n1071);
   U21793 : NAND2_X2 port map( A1 => n13267, A2 => n11786, ZN => n4770);
   U21797 : NAND2_X1 port map( A1 => n10071, A2 => n11441, ZN => n31124);
   U21814 : INV_X2 port map( I => n31128, ZN => n15189);
   U21823 : NOR2_X2 port map( A1 => n22870, A2 => n22869, ZN => n23439);
   U21844 : XOR2_X1 port map( A1 => n15543, A2 => n31132, Z => n25325);
   U21859 : XOR2_X1 port map( A1 => n14639, A2 => n25720, Z => n31133);
   U21864 : OAI21_X2 port map( A1 => n31784, A2 => n16501, B => n22890, ZN => 
                           n1563);
   U21866 : NAND3_X1 port map( A1 => n24911, A2 => n10099, A3 => n24910, ZN => 
                           n4898);
   U21876 : NOR3_X1 port map( A1 => n1032, A2 => n20379, A3 => n18078, ZN => 
                           n31135);
   U21878 : NAND2_X1 port map( A1 => n31137, A2 => n29385, ZN => n26696);
   U21881 : OAI21_X1 port map( A1 => n17712, A2 => n16516, B => n26547, ZN => 
                           n31137);
   U21883 : NAND2_X2 port map( A1 => n7281, A2 => n16009, ZN => n20624);
   U21890 : BUF_X2 port map( I => n19779, Z => n31138);
   U21894 : NAND3_X2 port map( A1 => n7396, A2 => n7395, A3 => n7834, ZN => 
                           n21037);
   U21895 : INV_X2 port map( I => n19002, ZN => n743);
   U21896 : NAND2_X2 port map( A1 => n6753, A2 => n9265, ZN => n19002);
   U21898 : XOR2_X1 port map( A1 => n27523, A2 => n26125, Z => n28119);
   U21899 : INV_X2 port map( I => n31140, ZN => n10955);
   U21915 : OAI21_X2 port map( A1 => n31145, A2 => n22482, B => n22480, ZN => 
                           n22824);
   U21931 : NOR2_X2 port map( A1 => n1353, A2 => n7280, ZN => n7397);
   U21933 : NAND2_X1 port map( A1 => n25877, A2 => n25709, ZN => n31146);
   U21939 : INV_X2 port map( I => n31147, ZN => n31579);
   U21942 : XNOR2_X1 port map( A1 => Plaintext(57), A2 => Key(57), ZN => n31147
                           );
   U21959 : NAND2_X2 port map( A1 => n11149, A2 => n11150, ZN => n15091);
   U21980 : NOR2_X2 port map( A1 => n6907, A2 => n9324, ZN => n9994);
   U21982 : XOR2_X1 port map( A1 => n24800, A2 => n26429, Z => n31151);
   U21983 : NAND2_X2 port map( A1 => n5119, A2 => n7995, ZN => n8800);
   U21984 : XOR2_X1 port map( A1 => n29728, A2 => n19769, Z => n2628);
   U21989 : NOR2_X2 port map( A1 => n3060, A2 => n3059, ZN => n19769);
   U22013 : XOR2_X1 port map( A1 => n8695, A2 => n27996, Z => n23341);
   U22016 : NOR2_X2 port map( A1 => n6676, A2 => n6677, ZN => n8695);
   U22018 : OR3_X1 port map( A1 => n11814, A2 => n14383, A3 => n3193, Z => 
                           n31583);
   U22019 : AOI21_X2 port map( A1 => n6108, A2 => n28423, B => n31157, ZN => 
                           n7292);
   U22027 : NOR2_X1 port map( A1 => n18973, A2 => n15502, ZN => n19227);
   U22035 : NAND2_X2 port map( A1 => n26627, A2 => n16713, ZN => n18973);
   U22039 : XOR2_X1 port map( A1 => n16319, A2 => n7511, Z => n24409);
   U22043 : NOR2_X2 port map( A1 => n23992, A2 => n28725, ZN => n16319);
   U22046 : BUF_X4 port map( I => n24789, Z => n31687);
   U22060 : XOR2_X1 port map( A1 => n31159, A2 => n14300, Z => Ciphertext(0));
   U22062 : AOI22_X1 port map( A1 => n6155, A2 => n6154, B1 => n8980, B2 => 
                           n10755, ZN => n31159);
   U22071 : OAI22_X2 port map( A1 => n29448, A2 => n15869, B1 => n15759, B2 => 
                           n18975, ZN => n19679);
   U22072 : XOR2_X1 port map( A1 => n22319, A2 => n22320, Z => n22324);
   U22088 : XOR2_X1 port map( A1 => n31527, A2 => n1695, Z => n13941);
   U22089 : INV_X2 port map( I => n5725, ZN => n31161);
   U22093 : NAND2_X2 port map( A1 => n3327, A2 => n31162, ZN => n22990);
   U22111 : XOR2_X1 port map( A1 => n3682, A2 => n22128, Z => n10889);
   U22112 : OAI21_X2 port map( A1 => n21487, A2 => n21488, B => n3685, ZN => 
                           n3682);
   U22128 : XOR2_X1 port map( A1 => n23306, A2 => n27252, Z => n2142);
   U22133 : XOR2_X1 port map( A1 => n343, A2 => n16322, Z => n22287);
   U22135 : XOR2_X1 port map( A1 => n7477, A2 => n22205, Z => n22313);
   U22148 : XOR2_X1 port map( A1 => n31168, A2 => n18166, Z => n20011);
   U22153 : XOR2_X1 port map( A1 => n18165, A2 => n19700, Z => n31168);
   U22161 : XOR2_X1 port map( A1 => n19485, A2 => n31169, Z => n19388);
   U22176 : XOR2_X1 port map( A1 => n2611, A2 => n27144, Z => n31169);
   U22180 : NAND2_X2 port map( A1 => n11287, A2 => n11310, ZN => n24158);
   U22181 : INV_X4 port map( I => n20375, ZN => n20361);
   U22194 : XOR2_X1 port map( A1 => n22259, A2 => n22261, Z => n18121);
   U22200 : XOR2_X1 port map( A1 => n22119, A2 => n22291, Z => n22259);
   U22202 : INV_X2 port map( I => n16042, ZN => n18539);
   U22207 : NAND2_X1 port map( A1 => n14156, A2 => n16042, ZN => n13787);
   U22222 : XOR2_X1 port map( A1 => Plaintext(135), A2 => Key(135), Z => n16042
                           );
   U22224 : NAND3_X1 port map( A1 => n15534, A2 => n28478, A3 => n33143, ZN => 
                           n11778);
   U22253 : XOR2_X1 port map( A1 => n19439, A2 => n15485, Z => n14459);
   U22257 : XOR2_X1 port map( A1 => n17554, A2 => n26530, Z => n6789);
   U22259 : NAND2_X1 port map( A1 => n18530, A2 => n18531, ZN => n18534);
   U22277 : OR2_X1 port map( A1 => n25316, A2 => n31178, Z => n17058);
   U22295 : OAI21_X2 port map( A1 => n22573, A2 => n1298, B => n31181, ZN => 
                           n10905);
   U22296 : OAI22_X2 port map( A1 => n22524, A2 => n1728, B1 => n901, B2 => 
                           n17960, ZN => n22605);
   U22304 : XOR2_X1 port map( A1 => n31182, A2 => n16690, Z => Ciphertext(30));
   U22308 : AOI21_X1 port map( A1 => n24250, A2 => n24251, B => n28553, ZN => 
                           n1513);
   U22312 : NAND2_X1 port map( A1 => n32902, A2 => n21374, ZN => n21377);
   U22314 : INV_X2 port map( I => n31184, ZN => n24874);
   U22319 : XOR2_X1 port map( A1 => n31186, A2 => n14754, Z => n11327);
   U22323 : XOR2_X1 port map( A1 => n22286, A2 => n11166, Z => n31186);
   U22329 : INV_X2 port map( I => n20872, ZN => n31189);
   U22332 : XOR2_X1 port map( A1 => n6327, A2 => n31190, Z => n6955);
   U22333 : XOR2_X1 port map( A1 => n21960, A2 => n31191, Z => n31190);
   U22341 : XOR2_X1 port map( A1 => n3982, A2 => n31194, Z => n14572);
   U22343 : XOR2_X1 port map( A1 => n17540, A2 => n17541, Z => n31194);
   U22347 : BUF_X2 port map( I => n8243, Z => n31195);
   U22351 : AOI22_X1 port map( A1 => n5638, A2 => n5043, B1 => n25223, B2 => 
                           n28358, ZN => n5243);
   U22353 : AND2_X1 port map( A1 => n16117, A2 => n1141, Z => n4496);
   U22367 : XOR2_X1 port map( A1 => n23341, A2 => n23340, Z => n31200);
   U22368 : XOR2_X1 port map( A1 => n17395, A2 => n31203, Z => n2104);
   U22371 : NAND2_X2 port map( A1 => n30744, A2 => n1430, ZN => n18187);
   U22373 : NAND2_X2 port map( A1 => n17900, A2 => n27067, ZN => n16076);
   U22382 : XOR2_X1 port map( A1 => n31205, A2 => n18898, Z => n27599);
   U22383 : XOR2_X1 port map( A1 => n19630, A2 => n4976, Z => n31205);
   U22386 : INV_X2 port map( I => n17906, ZN => n31208);
   U22395 : AOI22_X2 port map( A1 => n27975, A2 => n26160, B1 => n5400, B2 => 
                           n1265, ZN => n5399);
   U22399 : NAND2_X2 port map( A1 => n22977, A2 => n1484, ZN => n3600);
   U22411 : XOR2_X1 port map( A1 => n20715, A2 => n20926, Z => n20752);
   U22418 : NAND2_X2 port map( A1 => n12504, A2 => n31213, ZN => n12610);
   U22435 : XOR2_X1 port map( A1 => n31214, A2 => n25065, Z => Ciphertext(42));
   U22436 : NAND3_X2 port map( A1 => n22778, A2 => n22777, A3 => n22776, ZN => 
                           n23335);
   U22455 : NAND2_X1 port map( A1 => n24969, A2 => n3843, ZN => n13736);
   U22481 : NAND2_X2 port map( A1 => n10203, A2 => n19199, ZN => n19033);
   U22484 : NAND2_X2 port map( A1 => n22470, A2 => n4156, ZN => n22885);
   U22486 : INV_X2 port map( I => n11438, ZN => n24182);
   U22494 : AOI21_X1 port map( A1 => n21286, A2 => n21285, B => n21398, ZN => 
                           n27198);
   U22499 : XOR2_X1 port map( A1 => n14094, A2 => n19682, Z => n8921);
   U22504 : XOR2_X1 port map( A1 => n2261, A2 => n2554, Z => n31221);
   U22515 : NAND2_X1 port map( A1 => n21705, A2 => n21704, ZN => n21145);
   U22530 : NAND3_X1 port map( A1 => n24920, A2 => n15799, A3 => n15569, ZN => 
                           n24353);
   U22539 : XOR2_X1 port map( A1 => n29320, A2 => n24750, Z => n5525);
   U22541 : XOR2_X1 port map( A1 => n11562, A2 => n22189, Z => n11781);
   U22543 : NAND2_X2 port map( A1 => n12183, A2 => n16477, ZN => n22189);
   U22554 : OAI21_X2 port map( A1 => n7388, A2 => n21812, B => n5474, ZN => 
                           n11481);
   U22563 : XOR2_X1 port map( A1 => n20979, A2 => n31235, Z => n31234);
   U22579 : XOR2_X1 port map( A1 => n6706, A2 => n31703, Z => n31237);
   U22580 : XOR2_X1 port map( A1 => n16861, A2 => n17259, Z => n29101);
   U22581 : XOR2_X1 port map( A1 => n24676, A2 => n15161, Z => n15473);
   U22584 : NAND2_X2 port map( A1 => n31238, A2 => n13021, ZN => n20625);
   U22595 : OAI21_X2 port map( A1 => n9855, A2 => n27343, B => n19991, ZN => 
                           n31238);
   U22621 : NAND2_X2 port map( A1 => n31241, A2 => n13089, ZN => n20820);
   U22622 : OAI21_X2 port map( A1 => n10380, A2 => n19804, B => n2565, ZN => 
                           n31241);
   U22625 : NOR2_X2 port map( A1 => n2149, A2 => n2584, ZN => n18841);
   U22630 : NAND2_X1 port map( A1 => n19984, A2 => n11508, ZN => n31242);
   U22632 : XOR2_X1 port map( A1 => n1690, A2 => n31243, Z => n25345);
   U22638 : XOR2_X1 port map( A1 => n24626, A2 => n29346, Z => n31243);
   U22642 : XOR2_X1 port map( A1 => n15941, A2 => n16076, Z => n23505);
   U22645 : AOI21_X2 port map( A1 => n7882, A2 => n29118, B => n31246, ZN => 
                           n8908);
   U22651 : NAND2_X2 port map( A1 => n2448, A2 => n31247, ZN => n9919);
   U22652 : INV_X2 port map( I => n31248, ZN => n16966);
   U22667 : XOR2_X1 port map( A1 => n4013, A2 => n1128, Z => n31252);
   U22673 : XOR2_X1 port map( A1 => n4013, A2 => n9960, Z => n31253);
   U22695 : XOR2_X1 port map( A1 => n21950, A2 => n16692, Z => n22412);
   U22702 : XOR2_X1 port map( A1 => n1886, A2 => n31258, Z => n28260);
   U22709 : XOR2_X1 port map( A1 => n11012, A2 => n20749, Z => n31258);
   U22710 : XOR2_X1 port map( A1 => n24598, A2 => n24523, Z => n14918);
   U22711 : XOR2_X1 port map( A1 => n7574, A2 => n31259, Z => n24598);
   U22714 : INV_X2 port map( I => n24520, ZN => n31259);
   U22718 : BUF_X2 port map( I => n21122, Z => n31260);
   U22730 : OAI21_X2 port map( A1 => n15154, A2 => n31262, B => n12811, ZN => 
                           n21704);
   U22734 : NAND3_X2 port map( A1 => n21549, A2 => n21548, A3 => n21550, ZN => 
                           n22067);
   U22758 : OAI21_X2 port map( A1 => n17251, A2 => n15956, B => n31265, ZN => 
                           n31264);
   U22768 : NAND2_X2 port map( A1 => n14831, A2 => n15956, ZN => n31265);
   U22778 : OAI21_X1 port map( A1 => n12033, A2 => n22801, B => n26868, ZN => 
                           n12597);
   U22781 : NAND2_X2 port map( A1 => n20294, A2 => n20293, ZN => n20556);
   U22787 : XOR2_X1 port map( A1 => n12453, A2 => n19316, Z => n31828);
   U22788 : XOR2_X1 port map( A1 => n29030, A2 => n12048, Z => n12453);
   U22790 : XOR2_X1 port map( A1 => n20654, A2 => n28541, Z => n17973);
   U22811 : BUF_X2 port map( I => n11947, Z => n31268);
   U22822 : NAND2_X2 port map( A1 => n25968, A2 => n19115, ZN => n13330);
   U22829 : INV_X2 port map( I => n31272, ZN => n13255);
   U22832 : OR2_X1 port map( A1 => n22873, A2 => n22791, Z => n22872);
   U22835 : OAI22_X2 port map( A1 => n1664, A2 => n1663, B1 => n1661, B2 => 
                           n14253, ZN => n22873);
   U22866 : NAND3_X1 port map( A1 => n7924, A2 => n7926, A3 => n11571, ZN => 
                           n31281);
   U22870 : NOR2_X2 port map( A1 => n13482, A2 => n13481, ZN => n13477);
   U22894 : NAND2_X2 port map( A1 => n21550, A2 => n21494, ZN => n31284);
   U22906 : INV_X2 port map( I => n25144, ZN => n16751);
   U22909 : NAND2_X1 port map( A1 => n25144, A2 => n25145, ZN => n15330);
   U22911 : XOR2_X1 port map( A1 => n16719, A2 => n6452, Z => n25144);
   U22913 : NOR2_X2 port map( A1 => n10495, A2 => n31285, ZN => n10201);
   U22914 : AND2_X1 port map( A1 => n6696, A2 => n22944, Z => n31285);
   U22917 : OAI21_X2 port map( A1 => n31286, A2 => n20540, B => n26730, ZN => 
                           n26165);
   U22928 : INV_X2 port map( I => n31287, ZN => n634);
   U22930 : XNOR2_X1 port map( A1 => n22019, A2 => n8352, ZN => n31287);
   U22935 : OR2_X1 port map( A1 => n19203, A2 => n19291, Z => n31356);
   U22936 : NOR2_X2 port map( A1 => n1052, A2 => n19300, ZN => n19203);
   U22946 : XOR2_X1 port map( A1 => n28983, A2 => n20792, Z => n14647);
   U22956 : OAI21_X2 port map( A1 => n1572, A2 => n33548, B => n16538, ZN => 
                           n18403);
   U22957 : NAND2_X2 port map( A1 => n20625, A2 => n20623, ZN => n7280);
   U22959 : NAND2_X2 port map( A1 => n31292, A2 => n13397, ZN => n6679);
   U22963 : OAI21_X2 port map( A1 => n15477, A2 => n19935, B => n5371, ZN => 
                           n31292);
   U22988 : NAND2_X2 port map( A1 => n23109, A2 => n853, ZN => n23112);
   U22993 : XOR2_X1 port map( A1 => n31296, A2 => n8687, Z => n13272);
   U22997 : OR2_X1 port map( A1 => n12535, A2 => n861, Z => n21247);
   U22999 : NAND2_X1 port map( A1 => n7785, A2 => n7786, ZN => n31348);
   U23004 : XOR2_X1 port map( A1 => n2785, A2 => n2788, Z => n2784);
   U23021 : XOR2_X1 port map( A1 => n26754, A2 => n18188, Z => n679);
   U23031 : NOR2_X2 port map( A1 => n10444, A2 => n502, ZN => n9619);
   U23041 : XOR2_X1 port map( A1 => n20975, A2 => n16958, Z => n20887);
   U23048 : NAND2_X2 port map( A1 => n20311, A2 => n12902, ZN => n20975);
   U23057 : XOR2_X1 port map( A1 => n11504, A2 => n32981, Z => n14053);
   U23058 : NAND2_X2 port map( A1 => n23049, A2 => n23048, ZN => n11504);
   U23061 : XOR2_X1 port map( A1 => n11816, A2 => n31301, Z => n11833);
   U23063 : XOR2_X1 port map( A1 => n15950, A2 => n22265, Z => n31301);
   U23067 : NAND2_X2 port map( A1 => n23009, A2 => n23011, ZN => n6975);
   U23092 : AND2_X2 port map( A1 => n9753, A2 => n9750, Z => n22467);
   U23097 : XOR2_X1 port map( A1 => n22167, A2 => n16767, Z => n31303);
   U23098 : OR2_X1 port map( A1 => n18879, A2 => n8213, Z => n18441);
   U23106 : XNOR2_X1 port map( A1 => n30329, A2 => n21994, ZN => n21926);
   U23112 : NAND2_X2 port map( A1 => n21796, A2 => n21795, ZN => n21994);
   U23114 : NAND2_X2 port map( A1 => n25738, A2 => n27189, ZN => n4642);
   U23131 : OAI22_X2 port map( A1 => n18047, A2 => n9460, B1 => n15717, B2 => 
                           n27090, ZN => n12878);
   U23137 : OR2_X1 port map( A1 => n31960, A2 => n6442, Z => n26726);
   U23139 : OR2_X1 port map( A1 => n11932, A2 => n32606, Z => n16531);
   U23145 : OR2_X1 port map( A1 => n32414, A2 => n19128, Z => n31306);
   U23148 : NAND2_X2 port map( A1 => n28660, A2 => n5573, ZN => n28659);
   U23159 : XOR2_X1 port map( A1 => n1604, A2 => n31308, Z => n371);
   U23161 : INV_X1 port map( I => n25311, ZN => n31308);
   U23162 : NAND2_X2 port map( A1 => n1543, A2 => n1544, ZN => n1604);
   U23180 : NAND2_X2 port map( A1 => n27472, A2 => n15828, ZN => n22226);
   U23218 : XOR2_X1 port map( A1 => n24377, A2 => n31312, Z => n6293);
   U23223 : NOR2_X2 port map( A1 => n31798, A2 => n27752, ZN => n11330);
   U23225 : XOR2_X1 port map( A1 => n12980, A2 => n8992, Z => n4251);
   U23226 : AOI21_X2 port map( A1 => n21522, A2 => n21523, B => n21744, ZN => 
                           n21524);
   U23235 : INV_X4 port map( I => n31746, ZN => n4747);
   U23237 : NAND2_X2 port map( A1 => n3631, A2 => n3633, ZN => n15508);
   U23243 : NAND2_X1 port map( A1 => n23176, A2 => n28740, ZN => n31314);
   U23250 : XOR2_X1 port map( A1 => n31316, A2 => n17487, Z => n22679);
   U23253 : XOR2_X1 port map( A1 => n17486, A2 => n17485, Z => n31316);
   U23256 : XOR2_X1 port map( A1 => n32052, A2 => n21001, Z => n13336);
   U23264 : INV_X1 port map( I => n18540, ZN => n31821);
   U23267 : XOR2_X1 port map( A1 => n6808, A2 => n20678, Z => n7596);
   U23275 : XOR2_X1 port map( A1 => n20776, A2 => n12721, Z => n20678);
   U23276 : NOR2_X2 port map( A1 => n12864, A2 => n13764, ZN => n13811);
   U23277 : NAND2_X2 port map( A1 => n13555, A2 => n15156, ZN => n25546);
   U23278 : OR2_X1 port map( A1 => n14236, A2 => n6489, Z => n7476);
   U23281 : NAND2_X2 port map( A1 => n13690, A2 => n28138, ZN => n27996);
   U23285 : XNOR2_X1 port map( A1 => n20680, A2 => n20679, ZN => n31423);
   U23288 : OAI22_X2 port map( A1 => n17897, A2 => n17896, B1 => n28357, B2 => 
                           n2609, ZN => n20679);
   U23289 : INV_X2 port map( I => n6454, ZN => n22017);
   U23290 : OAI22_X2 port map( A1 => n28067, A2 => n28068, B1 => n4516, B2 => 
                           n28018, ZN => n6454);
   U23299 : AND2_X1 port map( A1 => n18540, A2 => n13363, Z => n18302);
   U23305 : NAND3_X2 port map( A1 => n4101, A2 => n24591, A3 => n25013, ZN => 
                           n14964);
   U23307 : XOR2_X1 port map( A1 => n3868, A2 => n23420, Z => n23359);
   U23316 : INV_X2 port map( I => n31318, ZN => n31920);
   U23321 : XOR2_X1 port map( A1 => n2044, A2 => n2043, Z => n31318);
   U23322 : NAND2_X1 port map( A1 => n25022, A2 => n13427, ZN => n2909);
   U23326 : NOR2_X2 port map( A1 => n1549, A2 => n31320, ZN => n25060);
   U23327 : XOR2_X1 port map( A1 => n13927, A2 => n13928, Z => n31321);
   U23344 : NOR2_X1 port map( A1 => n15133, A2 => n15132, ZN => n31323);
   U23347 : NAND2_X2 port map( A1 => n13279, A2 => n490, ZN => n12320);
   U23359 : NAND2_X1 port map( A1 => n9284, A2 => n14917, ZN => n12183);
   U23368 : OR2_X2 port map( A1 => n26733, A2 => n14082, Z => n20134);
   U23369 : NAND2_X1 port map( A1 => n31811, A2 => n20460, ZN => n20461);
   U23371 : INV_X2 port map( I => n17338, ZN => n25999);
   U23372 : OAI21_X2 port map( A1 => n17054, A2 => n18565, B => n17135, ZN => 
                           n17338);
   U23391 : NAND2_X2 port map( A1 => n13546, A2 => n13547, ZN => n17517);
   U23411 : NAND2_X1 port map( A1 => n31932, A2 => n17879, ZN => n31327);
   U23418 : XOR2_X1 port map( A1 => n9574, A2 => n6458, Z => n9436);
   U23420 : NAND2_X2 port map( A1 => n13285, A2 => n19892, ZN => n20228);
   U23421 : OAI21_X2 port map( A1 => n8147, A2 => n8146, B => n19891, ZN => 
                           n13285);
   U23441 : XOR2_X1 port map( A1 => n22172, A2 => n9129, Z => n15950);
   U23448 : OAI22_X2 port map( A1 => n28137, A2 => n21702, B1 => n11981, B2 => 
                           n32519, ZN => n22172);
   U23449 : OAI21_X2 port map( A1 => n31329, A2 => n11480, B => n12925, ZN => 
                           n7447);
   U23464 : XOR2_X1 port map( A1 => n31330, A2 => n1742, Z => n27819);
   U23475 : XOR2_X1 port map( A1 => n31331, A2 => n31336, Z => n31330);
   U23488 : INV_X1 port map( I => n15950, ZN => n31336);
   U23492 : OAI21_X1 port map( A1 => n17582, A2 => n17223, B => n31339, ZN => 
                           n14537);
   U23495 : XNOR2_X1 port map( A1 => n17090, A2 => n19573, ZN => n31387);
   U23499 : OAI21_X2 port map( A1 => n10405, A2 => n28613, B => n22876, ZN => 
                           n28364);
   U23508 : XOR2_X1 port map( A1 => n11636, A2 => n7889, Z => n14518);
   U23509 : NOR2_X2 port map( A1 => n28226, A2 => n11634, ZN => n11636);
   U23516 : NAND2_X2 port map( A1 => n31345, A2 => n31344, ZN => n9399);
   U23521 : XOR2_X1 port map( A1 => n31346, A2 => n9298, Z => n10258);
   U23528 : XOR2_X1 port map( A1 => n22271, A2 => n28575, Z => n28574);
   U23531 : NAND3_X1 port map( A1 => n16112, A2 => n12309, A3 => n25796, ZN => 
                           n25791);
   U23533 : XOR2_X1 port map( A1 => n7826, A2 => n31410, Z => n31529);
   U23536 : OR2_X1 port map( A1 => n26600, A2 => n19300, Z => n31350);
   U23550 : BUF_X2 port map( I => n8695, Z => n31354);
   U23552 : INV_X2 port map( I => n31357, ZN => n7915);
   U23560 : XOR2_X1 port map( A1 => n7916, A2 => n7917, Z => n31357);
   U23562 : XOR2_X1 port map( A1 => n13419, A2 => n24664, Z => n24814);
   U23566 : AOI21_X2 port map( A1 => n9367, A2 => n24061, B => n9366, ZN => 
                           n13419);
   U23569 : OAI21_X2 port map( A1 => n27466, A2 => n21871, B => n27596, ZN => 
                           n31359);
   U23571 : NAND2_X1 port map( A1 => n17255, A2 => n26249, ZN => n17062);
   U23605 : OR2_X1 port map( A1 => n15101, A2 => n12118, Z => n31365);
   U23607 : NOR2_X1 port map( A1 => n16453, A2 => n4016, ZN => n31366);
   U23608 : INV_X2 port map( I => n9468, ZN => n8491);
   U23612 : NAND2_X1 port map( A1 => n4806, A2 => n22905, ZN => n4805);
   U23614 : XOR2_X1 port map( A1 => n4791, A2 => n31367, Z => n23579);
   U23619 : XOR2_X1 port map( A1 => n31588, A2 => n4794, Z => n31367);
   U23620 : NAND2_X2 port map( A1 => n21085, A2 => n21170, ZN => n21354);
   U23624 : OAI21_X2 port map( A1 => n31369, A2 => n31368, B => n16819, ZN => 
                           n28073);
   U23626 : NOR2_X2 port map( A1 => n4259, A2 => n12074, ZN => n31368);
   U23627 : XOR2_X1 port map( A1 => n31370, A2 => n25519, Z => Ciphertext(119))
                           ;
   U23637 : NAND4_X2 port map( A1 => n4325, A2 => n16468, A3 => n18215, A4 => 
                           n25518, ZN => n31370);
   U23640 : XOR2_X1 port map( A1 => n17517, A2 => n5772, Z => n20897);
   U23645 : NAND2_X2 port map( A1 => n26082, A2 => n26296, ZN => n5772);
   U23649 : XOR2_X1 port map( A1 => n31371, A2 => n10024, Z => n10426);
   U23651 : XOR2_X1 port map( A1 => n19723, A2 => n15990, Z => n31371);
   U23652 : AND2_X1 port map( A1 => n9959, A2 => n11833, Z => n10310);
   U23660 : XOR2_X1 port map( A1 => n1259, A2 => n27708, Z => n8609);
   U23667 : NAND2_X2 port map( A1 => n31547, A2 => n5058, ZN => n27708);
   U23670 : XOR2_X1 port map( A1 => n20963, A2 => n20820, Z => n20888);
   U23672 : NAND2_X2 port map( A1 => n3835, A2 => n31372, ZN => n4450);
   U23676 : XOR2_X1 port map( A1 => n24528, A2 => n24529, Z => n16125);
   U23677 : INV_X2 port map( I => n24440, ZN => n31373);
   U23680 : BUF_X2 port map( I => n6500, Z => n31374);
   U23683 : NOR2_X1 port map( A1 => n16819, A2 => n31579, ZN => n18608);
   U23686 : XOR2_X1 port map( A1 => n17128, A2 => n17395, Z => n27135);
   U23689 : XOR2_X1 port map( A1 => n32537, A2 => n22192, Z => n12882);
   U23691 : XOR2_X1 port map( A1 => n6948, A2 => n29428, Z => n6093);
   U23702 : NOR2_X1 port map( A1 => n26445, A2 => n29302, ZN => n31379);
   U23721 : INV_X1 port map( I => n31532, ZN => n20476);
   U23723 : XOR2_X1 port map( A1 => n31380, A2 => n21930, Z => n9533);
   U23728 : NAND2_X1 port map( A1 => n9180, A2 => n25819, ZN => n31381);
   U23737 : NAND2_X2 port map( A1 => n3792, A2 => n29364, ZN => n13267);
   U23752 : AOI22_X2 port map( A1 => n31385, A2 => n12394, B1 => n5383, B2 => 
                           n4689, ZN => n22123);
   U23761 : NAND2_X1 port map( A1 => n26283, A2 => n12354, ZN => n31385);
   U23767 : XOR2_X1 port map( A1 => n13780, A2 => n31387, Z => n245);
   U23782 : NOR2_X1 port map( A1 => n20329, A2 => n31390, ZN => n31389);
   U23786 : NAND3_X1 port map( A1 => n15304, A2 => n12308, A3 => n12309, ZN => 
                           n28989);
   U23789 : INV_X2 port map( I => n5016, ZN => n31458);
   U23790 : INV_X2 port map( I => n9285, ZN => n14384);
   U23792 : XOR2_X1 port map( A1 => n17014, A2 => n17012, Z => n17015);
   U23800 : NAND2_X1 port map( A1 => n10419, A2 => n31393, ZN => n27738);
   U23811 : XOR2_X1 port map( A1 => n31395, A2 => n7866, Z => n7865);
   U23816 : NOR2_X2 port map( A1 => n31397, A2 => n78, ZN => n1471);
   U23820 : NOR2_X1 port map( A1 => n4935, A2 => n23110, ZN => n31397);
   U23829 : NOR2_X2 port map( A1 => n8425, A2 => n31398, ZN => n20425);
   U23850 : INV_X1 port map( I => n1260, ZN => n6905);
   U23869 : AOI21_X2 port map( A1 => n31400, A2 => n12140, B => n32397, ZN => 
                           n28439);
   U23871 : XOR2_X1 port map( A1 => n9353, A2 => n5268, Z => n12422);
   U23892 : BUF_X2 port map( I => n13622, Z => n31402);
   U23908 : NAND2_X1 port map( A1 => n26637, A2 => n12265, ZN => n12264);
   U23932 : XOR2_X1 port map( A1 => n12212, A2 => n19729, Z => n4631);
   U23934 : NAND2_X2 port map( A1 => n8717, A2 => n8716, ZN => n12212);
   U23935 : XOR2_X1 port map( A1 => n18042, A2 => n24379, Z => n31405);
   U23940 : NAND2_X2 port map( A1 => n10854, A2 => n31406, ZN => n19597);
   U23942 : NAND3_X1 port map( A1 => n25671, A2 => n25673, A3 => n25672, ZN => 
                           n31478);
   U23946 : XOR2_X1 port map( A1 => n16893, A2 => n14851, Z => n16896);
   U23947 : NOR2_X2 port map( A1 => n27753, A2 => n27754, ZN => n16893);
   U23952 : INV_X2 port map( I => n31409, ZN => n17133);
   U23957 : NAND2_X1 port map( A1 => n1387, A2 => n18994, ZN => n18943);
   U23971 : XOR2_X1 port map( A1 => n22033, A2 => n25801, Z => n22034);
   U23977 : NAND2_X2 port map( A1 => n16888, A2 => n16889, ZN => n22033);
   U23981 : AND2_X1 port map( A1 => n13921, A2 => n5480, Z => n11457);
   U24000 : XOR2_X1 port map( A1 => n19345, A2 => n5526, Z => n17575);
   U24006 : INV_X2 port map( I => n20371, ZN => n20533);
   U24010 : XOR2_X1 port map( A1 => n20853, A2 => n17957, Z => n21220);
   U24019 : AOI21_X1 port map( A1 => n2858, A2 => n5962, B => n4459, ZN => 
                           n3810);
   U24036 : NAND2_X2 port map( A1 => n18928, A2 => n18927, ZN => n31415);
   U24056 : NOR2_X1 port map( A1 => n11596, A2 => n21876, ZN => n14822);
   U24063 : NAND2_X1 port map( A1 => n31922, A2 => n20133, ZN => n19806);
   U24073 : NOR2_X1 port map( A1 => n7802, A2 => n14129, ZN => n13838);
   U24087 : NAND2_X2 port map( A1 => n13878, A2 => n28850, ZN => n24204);
   U24088 : NAND2_X2 port map( A1 => n10848, A2 => n32953, ZN => n31422);
   U24097 : XOR2_X1 port map( A1 => n31423, A2 => n20678, Z => n18025);
   U24109 : NAND3_X2 port map( A1 => n4717, A2 => n5561, A3 => n5560, ZN => 
                           n9319);
   U24116 : NOR3_X1 port map( A1 => n18884, A2 => n18660, A3 => n18888, ZN => 
                           n10537);
   U24126 : OAI21_X2 port map( A1 => n29379, A2 => n31424, B => n10381, ZN => 
                           n13205);
   U24145 : XOR2_X1 port map( A1 => n31426, A2 => n24795, Z => n12637);
   U24147 : XOR2_X1 port map( A1 => n10870, A2 => n4997, Z => n31426);
   U24150 : NAND2_X2 port map( A1 => n6362, A2 => n28943, ZN => n19265);
   U24151 : XOR2_X1 port map( A1 => n20899, A2 => n15275, Z => n21041);
   U24155 : XOR2_X1 port map( A1 => n23284, A2 => n31429, Z => n10525);
   U24159 : NAND2_X2 port map( A1 => n31689, A2 => n1668, ZN => n14392);
   U24207 : XOR2_X1 port map( A1 => n31432, A2 => n16551, Z => Ciphertext(190))
                           ;
   U24213 : NAND4_X2 port map( A1 => n25920, A2 => n25919, A3 => n25918, A4 => 
                           n25917, ZN => n31432);
   U24218 : XOR2_X1 port map( A1 => n28633, A2 => n22224, Z => n8275);
   U24240 : NOR2_X2 port map( A1 => n24265, A2 => n31096, ZN => n24230);
   U24253 : NAND2_X2 port map( A1 => n21405, A2 => n32069, ZN => n15807);
   U24279 : NOR2_X2 port map( A1 => n26220, A2 => n27329, ZN => n24141);
   U24290 : XOR2_X1 port map( A1 => n19550, A2 => n19661, Z => n19739);
   U24293 : NAND2_X2 port map( A1 => n3072, A2 => n6576, ZN => n19550);
   U24313 : XOR2_X1 port map( A1 => n14689, A2 => n1230, Z => n31440);
   U24314 : INV_X2 port map( I => n8327, ZN => n26733);
   U24317 : INV_X1 port map( I => n31564, ZN => n22915);
   U24338 : XOR2_X1 port map( A1 => n11868, A2 => n24442, Z => n14362);
   U24348 : INV_X2 port map( I => n31445, ZN => n29253);
   U24349 : XOR2_X1 port map( A1 => n8772, A2 => n8771, Z => n31445);
   U24386 : NAND2_X1 port map( A1 => n26284, A2 => n17626, ZN => n16411);
   U24389 : NAND3_X1 port map( A1 => n547, A2 => n24466, A3 => n12358, ZN => 
                           n3828);
   U24398 : BUF_X2 port map( I => n19629, Z => n31450);
   U24400 : XOR2_X1 port map( A1 => n24416, A2 => n7837, Z => n5146);
   U24410 : NAND3_X2 port map( A1 => n20406, A2 => n32061, A3 => n10849, ZN => 
                           n9597);
   U24421 : NAND2_X2 port map( A1 => n1913, A2 => n1910, ZN => n21655);
   U24451 : OAI22_X2 port map( A1 => n13262, A2 => n6392, B1 => n13261, B2 => 
                           n12658, ZN => n24180);
   U24463 : INV_X2 port map( I => n26785, ZN => n31457);
   U24465 : NAND2_X2 port map( A1 => n21472, A2 => n21471, ZN => n26785);
   U24476 : OAI21_X2 port map( A1 => n4585, A2 => n10849, B => n4586, ZN => 
                           n7954);
   U24481 : AND2_X1 port map( A1 => n564, A2 => n13510, Z => n12179);
   U24485 : NOR2_X1 port map( A1 => n2958, A2 => n31504, ZN => n15953);
   U24499 : NAND2_X1 port map( A1 => n28435, A2 => n31458, ZN => n8584);
   U24526 : OAI22_X1 port map( A1 => n23729, A2 => n23939, B1 => n23730, B2 => 
                           n23731, ZN => n26220);
   U24544 : INV_X4 port map( I => n32040, ZN => n21811);
   U24548 : NAND3_X1 port map( A1 => n29351, A2 => n15084, A3 => n17787, ZN => 
                           n12004);
   U24550 : XOR2_X1 port map( A1 => n1344, A2 => n1923, Z => n5067);
   U24552 : INV_X2 port map( I => n31467, ZN => n31914);
   U24555 : NAND2_X2 port map( A1 => n28350, A2 => n9214, ZN => n3205);
   U24559 : OAI21_X1 port map( A1 => n4415, A2 => n25736, B => n25739, ZN => 
                           n7038);
   U24561 : NAND2_X2 port map( A1 => n1601, A2 => n1600, ZN => n4415);
   U24584 : XOR2_X1 port map( A1 => n30304, A2 => n20872, Z => n26647);
   U24587 : INV_X2 port map( I => n15299, ZN => n15301);
   U24589 : OAI22_X2 port map( A1 => n15450, A2 => n13966, B1 => n15449, B2 => 
                           n15448, ZN => n15299);
   U24591 : NOR2_X2 port map( A1 => n31473, A2 => n28882, ZN => n7312);
   U24596 : NAND2_X1 port map( A1 => n21270, A2 => n11814, ZN => n31474);
   U24600 : XOR2_X1 port map( A1 => n24116, A2 => n17912, Z => n24574);
   U24603 : AOI21_X1 port map( A1 => n23940, A2 => n11933, B => n757, ZN => n98
                           );
   U24607 : OAI21_X1 port map( A1 => n16425, A2 => n24064, B => n25570, ZN => 
                           n27354);
   U24608 : NOR2_X2 port map( A1 => n28488, A2 => n10428, ZN => n16425);
   U24610 : XOR2_X1 port map( A1 => n31478, A2 => n16687, Z => Ciphertext(145))
                           ;
   U24618 : NAND2_X2 port map( A1 => n5886, A2 => n12264, ZN => n12611);
   U24624 : NAND2_X2 port map( A1 => n21180, A2 => n21179, ZN => n26439);
   U24633 : NOR2_X1 port map( A1 => n24729, A2 => n4490, ZN => n4492);
   U24635 : INV_X1 port map( I => n25762, ZN => n24729);
   U24636 : NAND3_X2 port map( A1 => n4713, A2 => n4710, A3 => n4711, ZN => 
                           n23292);
   U24637 : NOR2_X1 port map( A1 => n563, A2 => n9469, ZN => n7014);
   U24646 : NOR2_X1 port map( A1 => n18711, A2 => n11707, ZN => n18506);
   U24677 : NAND3_X1 port map( A1 => n6595, A2 => n17637, A3 => n33400, ZN => 
                           n25518);
   U24678 : NAND2_X2 port map( A1 => n13246, A2 => n13247, ZN => n19866);
   U24697 : XOR2_X1 port map( A1 => n210, A2 => n22231, Z => n31486);
   U24704 : NAND2_X2 port map( A1 => n31487, A2 => n13003, ZN => n15613);
   U24711 : OAI21_X2 port map( A1 => n13006, A2 => n22861, B => n22895, ZN => 
                           n31487);
   U24713 : NAND2_X1 port map( A1 => n23943, A2 => n3375, ZN => n27078);
   U24739 : NOR2_X2 port map( A1 => n32076, A2 => n21700, ZN => n28137);
   U24744 : XOR2_X1 port map( A1 => n31488, A2 => n32796, Z => Ciphertext(129))
                           ;
   U24747 : NOR2_X1 port map( A1 => n31489, A2 => n6114, ZN => n31488);
   U24750 : NAND2_X1 port map( A1 => n25696, A2 => n25695, ZN => n31490);
   U24765 : NOR2_X2 port map( A1 => n28278, A2 => n5170, ZN => n27704);
   U24780 : XOR2_X1 port map( A1 => n128, A2 => n19555, Z => n17559);
   U24783 : XNOR2_X1 port map( A1 => n9189, A2 => n28188, ZN => n31552);
   U24787 : XOR2_X1 port map( A1 => n20754, A2 => n13041, Z => n20889);
   U24794 : NAND2_X2 port map( A1 => n20399, A2 => n26216, ZN => n20754);
   U24824 : AND2_X1 port map( A1 => n12932, A2 => n14770, Z => n7767);
   U24826 : XOR2_X1 port map( A1 => n23296, A2 => n23206, Z => n8810);
   U24834 : AOI21_X2 port map( A1 => n18124, A2 => n17360, B => n31500, ZN => 
                           n19300);
   U24835 : OAI22_X2 port map( A1 => n17599, A2 => n18863, B1 => n15583, B2 => 
                           n17360, ZN => n31500);
   U24850 : NAND2_X2 port map( A1 => n13852, A2 => n16694, ZN => n19862);
   U24856 : NOR2_X1 port map( A1 => n11173, A2 => n14055, ZN => n5662);
   U24860 : NAND3_X1 port map( A1 => n5774, A2 => n5773, A3 => n24919, ZN => 
                           n439);
   U24864 : AOI21_X2 port map( A1 => n10808, A2 => n29963, B => n31503, ZN => 
                           n18321);
   U24870 : NOR2_X2 port map( A1 => n10315, A2 => n11146, ZN => n31505);
   U24888 : NAND2_X2 port map( A1 => n31675, A2 => n17443, ZN => n9403);
   U24896 : OAI21_X2 port map( A1 => n22881, A2 => n33395, B => n17463, ZN => 
                           n23534);
   U24910 : XNOR2_X1 port map( A1 => n19395, A2 => n17369, ZN => n19709);
   U24933 : NAND2_X2 port map( A1 => n13937, A2 => n13939, ZN => n19395);
   U24937 : OAI21_X1 port map( A1 => n406, A2 => n405, B => n25863, ZN => 
                           n27217);
   U24941 : NAND2_X2 port map( A1 => n26778, A2 => n16641, ZN => n4335);
   U24953 : XOR2_X1 port map( A1 => n31509, A2 => n24828, Z => n1851);
   U24957 : XOR2_X1 port map( A1 => n11612, A2 => n11610, Z => n8042);
   U24977 : INV_X4 port map( I => n22977, ZN => n31549);
   U24984 : XOR2_X1 port map( A1 => n14348, A2 => n31510, Z => n23567);
   U24989 : XOR2_X1 port map( A1 => n23184, A2 => n4003, Z => n31510);
   U24995 : NAND2_X2 port map( A1 => n9170, A2 => n22390, ZN => n22393);
   U24996 : XOR2_X1 port map( A1 => n12410, A2 => n31512, Z => n18200);
   U24998 : XOR2_X1 port map( A1 => n19740, A2 => n31513, Z => n31512);
   U25016 : XOR2_X1 port map( A1 => n14645, A2 => n31516, Z => n13556);
   U25017 : NAND2_X1 port map( A1 => n13468, A2 => n13467, ZN => n31516);
   U25046 : INV_X2 port map( I => n6544, ZN => n21854);
   U25047 : XOR2_X1 port map( A1 => n19509, A2 => n15844, Z => n19544);
   U25048 : INV_X2 port map( I => n4820, ZN => n23741);
   U25050 : NOR2_X2 port map( A1 => n28616, A2 => n31521, ZN => n16453);
   U25064 : XOR2_X1 port map( A1 => n23258, A2 => n29190, Z => n17549);
   U25082 : XOR2_X1 port map( A1 => n31525, A2 => n29400, Z => n26433);
   U25088 : XOR2_X1 port map( A1 => n1303, A2 => n3142, Z => n31525);
   U25089 : XOR2_X1 port map( A1 => n17551, A2 => n15064, Z => n19468);
   U25099 : NAND2_X2 port map( A1 => n18505, A2 => n18504, ZN => n17551);
   U25102 : XOR2_X1 port map( A1 => n1694, A2 => n19552, Z => n31527);
   U25116 : INV_X2 port map( I => n13507, ZN => n13921);
   U25130 : XOR2_X1 port map( A1 => n13504, A2 => n12749, Z => n13507);
   U25131 : NAND4_X2 port map( A1 => n28728, A2 => n31528, A3 => n3401, A4 => 
                           n17578, ZN => n24189);
   U25132 : XOR2_X1 port map( A1 => n3009, A2 => n20926, Z => n20691);
   U25133 : XOR2_X1 port map( A1 => n10949, A2 => n9706, Z => n8312);
   U25139 : XOR2_X1 port map( A1 => n13829, A2 => n31529, Z => n6209);
   U25146 : XOR2_X1 port map( A1 => n19655, A2 => n29426, Z => n31534);
   U25156 : XOR2_X1 port map( A1 => n27951, A2 => n13876, Z => n292);
   U25199 : INV_X2 port map( I => n19124, ZN => n16288);
   U25202 : NAND2_X2 port map( A1 => n26442, A2 => n10564, ZN => n19124);
   U25221 : XOR2_X1 port map( A1 => n8424, A2 => n11321, Z => n31538);
   U25247 : INV_X2 port map( I => n16588, ZN => n31542);
   U25262 : NAND2_X1 port map( A1 => n25243, A2 => n31545, ZN => n4552);
   U25271 : OAI21_X2 port map( A1 => n29421, A2 => n31548, B => n11399, ZN => 
                           n31547);
   U25285 : NAND2_X2 port map( A1 => n28205, A2 => n31902, ZN => n5696);
   U25291 : NOR2_X1 port map( A1 => n17338, A2 => n19124, ZN => n18963);
   U25297 : AOI21_X2 port map( A1 => n18106, A2 => n11745, B => n21055, ZN => 
                           n28396);
   U25298 : XOR2_X1 port map( A1 => n22185, A2 => n11458, Z => n22110);
   U25302 : NAND2_X2 port map( A1 => n13034, A2 => n13803, ZN => n22185);
   U25311 : XOR2_X1 port map( A1 => n20960, A2 => n7717, Z => n20962);
   U25315 : XOR2_X1 port map( A1 => n1560, A2 => n16733, Z => n24762);
   U25319 : OR2_X1 port map( A1 => n13382, A2 => n2547, Z => n7964);
   U25331 : NAND2_X2 port map( A1 => n26835, A2 => n26834, ZN => n10987);
   U25332 : NAND2_X2 port map( A1 => n4135, A2 => n23018, ZN => n22883);
   U25337 : XOR2_X1 port map( A1 => n22084, A2 => n22195, Z => n10462);
   U25341 : INV_X2 port map( I => n31561, ZN => n4425);
   U25342 : INV_X2 port map( I => n31562, ZN => n31921);
   U25346 : XOR2_X1 port map( A1 => n4222, A2 => n24855, Z => n31562);
   U25351 : NAND3_X2 port map( A1 => n18966, A2 => n18964, A3 => n18965, ZN => 
                           n19398);
   U25354 : NAND3_X2 port map( A1 => n13653, A2 => n21863, A3 => n12724, ZN => 
                           n9129);
   U25383 : NOR3_X2 port map( A1 => n12280, A2 => n12279, A3 => n1, ZN => 
                           n12276);
   U25401 : OAI21_X2 port map( A1 => n12416, A2 => n9377, B => n29325, ZN => 
                           n12781);
   U25409 : NOR2_X1 port map( A1 => n17462, A2 => n31566, ZN => n28778);
   U25415 : XOR2_X1 port map( A1 => n10077, A2 => n10079, Z => n31671);
   U25426 : OAI21_X1 port map( A1 => n25621, A2 => n25705, B => n31570, ZN => 
                           n31569);
   U25427 : XOR2_X1 port map( A1 => n31571, A2 => n24707, Z => Ciphertext(110))
                           ;
   U25435 : NOR2_X1 port map( A1 => n21243, A2 => n11912, ZN => n25942);
   U25438 : AOI21_X1 port map( A1 => n31614, A2 => n21147, B => n15149, ZN => 
                           n4293);
   U25439 : XOR2_X1 port map( A1 => n24746, A2 => n24681, Z => n24684);
   U25442 : NOR2_X2 port map( A1 => n6600, A2 => n16445, ZN => n22121);
   U25447 : NAND2_X2 port map( A1 => n17017, A2 => n26998, ZN => n22138);
   U25455 : XOR2_X1 port map( A1 => Plaintext(91), A2 => Key(91), Z => n31574);
   U25461 : NOR2_X2 port map( A1 => n28737, A2 => n398, ZN => n1889);
   U25466 : XNOR2_X1 port map( A1 => n7989, A2 => n7988, ZN => n26699);
   U25468 : XOR2_X1 port map( A1 => n3083, A2 => n12014, Z => n3082);
   U25472 : XOR2_X1 port map( A1 => n31575, A2 => n32025, Z => n28595);
   U25479 : AND2_X1 port map( A1 => n6593, A2 => n22955, Z => n26507);
   U25501 : NAND2_X2 port map( A1 => n28081, A2 => n32032, ZN => n13617);
   U25512 : NAND2_X2 port map( A1 => n1956, A2 => n1954, ZN => n28390);
   U25525 : NAND2_X1 port map( A1 => n25963, A2 => n22350, ZN => n13561);
   U25530 : NAND2_X1 port map( A1 => n3448, A2 => n3449, ZN => n3447);
   U25532 : NAND2_X2 port map( A1 => n31585, A2 => n20229, ZN => n20413);
   U25540 : XOR2_X1 port map( A1 => n19679, A2 => n19743, Z => n19680);
   U25560 : NAND2_X1 port map( A1 => n21414, A2 => n8657, ZN => n5758);
   U25561 : XOR2_X1 port map( A1 => n702, A2 => n24527, Z => n7937);
   U25577 : NAND2_X2 port map( A1 => n4985, A2 => n50, ZN => n702);
   U25584 : XOR2_X1 port map( A1 => n4732, A2 => n1262, Z => n31588);
   U25620 : XOR2_X1 port map( A1 => n4756, A2 => n4759, Z => n6684);
   U25621 : XOR2_X1 port map( A1 => n31590, A2 => n22147, Z => n26462);
   U25624 : XOR2_X1 port map( A1 => n19711, A2 => n19398, Z => n19462);
   U25625 : AOI22_X2 port map( A1 => n32028, A2 => n27127, B1 => n146, B2 => 
                           n7065, ZN => n31591);
   U25669 : OAI21_X2 port map( A1 => n15898, A2 => n1153, B => n8206, ZN => 
                           n10324);
   U25672 : XOR2_X1 port map( A1 => n20804, A2 => n21047, Z => n20552);
   U25682 : NAND2_X1 port map( A1 => n8506, A2 => n19143, ZN => n16790);
   U25683 : INV_X2 port map( I => n31594, ZN => n31916);
   U25688 : XOR2_X1 port map( A1 => n10536, A2 => n2164, Z => n31594);
   U25705 : XOR2_X1 port map( A1 => n31596, A2 => n23276, Z => n10536);
   U25714 : XOR2_X1 port map( A1 => n13287, A2 => n721, Z => n31596);
   U25716 : XOR2_X1 port map( A1 => n27633, A2 => n29350, Z => n22223);
   U25720 : INV_X2 port map( I => n22317, ZN => n31597);
   U25722 : XOR2_X1 port map( A1 => n31598, A2 => n3540, Z => n10430);
   U25733 : NAND3_X1 port map( A1 => n27658, A2 => n21365, A3 => n12756, ZN => 
                           n1688);
   U25748 : XOR2_X1 port map( A1 => n31599, A2 => n13033, Z => Ciphertext(161))
                           ;
   U25794 : XOR2_X1 port map( A1 => n22260, A2 => n21959, Z => n31606);
   U25796 : NAND3_X1 port map( A1 => n29390, A2 => n29508, A3 => n31607, ZN => 
                           n11854);
   U25797 : NAND2_X1 port map( A1 => n22659, A2 => n22926, ZN => n31607);
   U25800 : INV_X2 port map( I => n14983, ZN => n21568);
   U25808 : XOR2_X1 port map( A1 => n24596, A2 => n24634, Z => n23554);
   U25815 : XOR2_X1 port map( A1 => n24740, A2 => n12067, Z => n24745);
   U25818 : XOR2_X1 port map( A1 => n7731, A2 => n24370, Z => n24740);
   U25831 : XOR2_X1 port map( A1 => n8795, A2 => n31608, Z => n4134);
   U25838 : NAND2_X1 port map( A1 => n31617, A2 => n712, ZN => n1830);
   U25847 : OR2_X1 port map( A1 => n16421, A2 => n4145, Z => n31619);
   U25855 : INV_X2 port map( I => n31622, ZN => n23603);
   U25857 : XOR2_X1 port map( A1 => n22969, A2 => n5263, Z => n31622);
   U25860 : AOI22_X1 port map( A1 => n23643, A2 => n15732, B1 => n6759, B2 => 
                           n11888, ZN => n31623);
   U25866 : XOR2_X1 port map( A1 => n7363, A2 => n10201, Z => n23257);
   U25871 : XOR2_X1 port map( A1 => n32604, A2 => n3682, Z => n31626);
   U25873 : NAND3_X2 port map( A1 => n21811, A2 => n29864, A3 => n8140, ZN => 
                           n31627);
   U25876 : NAND2_X1 port map( A1 => n18582, A2 => n18584, ZN => n6207);
   U25877 : OR2_X1 port map( A1 => n22640, A2 => n31914, Z => n6242);
   U25886 : XOR2_X1 port map( A1 => n31630, A2 => n14217, Z => n14216);
   U25887 : XOR2_X1 port map( A1 => n1004, A2 => n13146, Z => n31630);
   U25892 : INV_X2 port map( I => n20635, ZN => n867);
   U25894 : XOR2_X1 port map( A1 => n13855, A2 => n13853, Z => n27698);
   U25901 : NAND2_X1 port map( A1 => n22816, A2 => n33675, ZN => n22818);
   U25914 : OAI21_X1 port map( A1 => n2576, A2 => n16023, B => n21763, ZN => 
                           n26522);
   U25915 : NAND2_X1 port map( A1 => n31635, A2 => n31634, ZN => n22360);
   U25920 : XOR2_X1 port map( A1 => n19500, A2 => n29343, Z => n31638);
   U25921 : NAND2_X1 port map( A1 => n14840, A2 => n2826, ZN => n14592);
   U25925 : XOR2_X1 port map( A1 => n1937, A2 => n1936, Z => n1935);
   U25934 : XOR2_X1 port map( A1 => n6091, A2 => n23443, Z => n6090);
   U25936 : NAND2_X2 port map( A1 => n11643, A2 => n11645, ZN => n22137);
   U25943 : XOR2_X1 port map( A1 => n27395, A2 => n31361, Z => n31642);
   U25944 : NAND3_X2 port map( A1 => n2245, A2 => n2247, A3 => n16651, ZN => 
                           n31643);
   U25949 : AOI21_X2 port map( A1 => n19994, A2 => n19846, B => n17882, ZN => 
                           n31644);
   U25952 : AND2_X1 port map( A1 => n16354, A2 => n19301, Z => n19030);
   U25953 : INV_X2 port map( I => n7971, ZN => n19737);
   U25954 : XOR2_X1 port map( A1 => n7971, A2 => n31646, Z => n101);
   U25955 : NAND2_X2 port map( A1 => n19094, A2 => n19095, ZN => n31658);
   U25964 : NAND2_X2 port map( A1 => n27630, A2 => n27631, ZN => n21681);
   U25987 : XOR2_X1 port map( A1 => n9103, A2 => n29445, Z => n27058);
   U25997 : XOR2_X1 port map( A1 => n31655, A2 => n5714, Z => n560);
   U26003 : AND2_X1 port map( A1 => n17341, A2 => n4274, Z => n31673);
   U26006 : OAI22_X1 port map( A1 => n26198, A2 => n24955, B1 => n965, B2 => 
                           n24947, ZN => n24941);
   U26012 : NOR2_X1 port map( A1 => n27610, A2 => n25057, ZN => n31661);
   U26013 : INV_X1 port map( I => n27609, ZN => n31662);
   U26016 : NAND2_X1 port map( A1 => n31663, A2 => n17409, ZN => n11962);
   U26033 : NAND2_X2 port map( A1 => n26851, A2 => n15158, ZN => n10048);
   U26043 : XOR2_X1 port map( A1 => n31666, A2 => n24802, Z => n27812);
   U26044 : XOR2_X1 port map( A1 => n24799, A2 => n2864, Z => n31666);
   U26046 : OR2_X1 port map( A1 => n28228, A2 => n7862, Z => n25102);
   U26047 : AOI21_X1 port map( A1 => n31667, A2 => n34167, B => n23910, ZN => 
                           n12775);
   U26054 : NAND2_X2 port map( A1 => n10713, A2 => n18479, ZN => n7462);
   U26057 : NAND2_X2 port map( A1 => n31670, A2 => n31669, ZN => n10713);
   U26062 : NAND2_X1 port map( A1 => n16326, A2 => n16325, ZN => n27900);
   U26067 : NAND2_X2 port map( A1 => n25542, A2 => n25557, ZN => n25555);
   U26069 : INV_X1 port map( I => n5587, ZN => n18680);
   U26073 : NOR2_X1 port map( A1 => n16805, A2 => n18660, ZN => n5587);
   U26075 : AOI21_X2 port map( A1 => n21169, A2 => n11678, B => n31674, ZN => 
                           n3001);
   U26076 : AOI21_X2 port map( A1 => n15843, A2 => n15842, B => n19282, ZN => 
                           n15844);
   U26082 : NAND2_X2 port map( A1 => n27900, A2 => n23978, ZN => n25973);
   U26083 : AOI22_X2 port map( A1 => n7997, A2 => n30692, B1 => n17442, B2 => 
                           n17441, ZN => n31675);
   U26087 : NAND2_X2 port map( A1 => n31676, A2 => n27992, ZN => n20335);
   U26094 : XOR2_X1 port map( A1 => n26279, A2 => n14791, Z => n14190);
   U26095 : NOR2_X2 port map( A1 => n19284, A2 => n10943, ZN => n28949);
   U26096 : NAND2_X1 port map( A1 => n19523, A2 => n31678, ZN => n19528);
   U26097 : NAND2_X1 port map( A1 => n15593, A2 => n19834, ZN => n31678);
   U26099 : XOR2_X1 port map( A1 => n2353, A2 => n17968, Z => n26996);
   U26102 : NOR2_X1 port map( A1 => n793, A2 => n719, ZN => n31679);
   U26107 : XOR2_X1 port map( A1 => n31043, A2 => n5101, Z => n5100);
   U26112 : XOR2_X1 port map( A1 => n24782, A2 => n27153, Z => n13086);
   U26113 : NOR3_X1 port map( A1 => n25546, A2 => n25557, A3 => n25542, ZN => 
                           n15132);
   U26117 : XOR2_X1 port map( A1 => n9327, A2 => n19689, Z => n9326);
   U26118 : XOR2_X1 port map( A1 => n19589, A2 => n19508, Z => n19689);
   U26124 : NOR3_X1 port map( A1 => n17306, A2 => n15425, A3 => n29063, ZN => 
                           n6849);
   U26126 : INV_X2 port map( I => n14911, ZN => n29063);
   U26136 : XNOR2_X1 port map( A1 => n23498, A2 => n23497, ZN => n31709);
   U26142 : OAI21_X2 port map( A1 => n18813, A2 => n17370, B => n31682, ZN => 
                           n8741);
   U26147 : BUF_X2 port map( I => n16811, Z => n31683);
   U26154 : OAI21_X2 port map( A1 => n2060, A2 => n3821, B => n31686, ZN => 
                           n1917);
   U26155 : AOI22_X2 port map( A1 => n534, A2 => n1326, B1 => n1, B2 => n16736,
                           ZN => n31686);
   U26160 : XOR2_X1 port map( A1 => n24636, A2 => n24832, Z => n24600);
   U26163 : OR2_X1 port map( A1 => n27419, A2 => n33675, Z => n22817);
   U26167 : NOR2_X1 port map( A1 => n12329, A2 => n32900, ZN => n25078);
   U26168 : OAI21_X2 port map( A1 => n6204, A2 => n28706, B => n24889, ZN => 
                           n14650);
   U26174 : NAND2_X2 port map( A1 => n31695, A2 => n31693, ZN => n19909);
   U26175 : NAND3_X1 port map( A1 => n4143, A2 => n16298, A3 => n4142, ZN => 
                           n31695);
   U26183 : NOR2_X1 port map( A1 => n8010, A2 => n8605, ZN => n16779);
   U26191 : XOR2_X1 port map( A1 => n19620, A2 => n31698, Z => n11545);
   U26193 : XOR2_X1 port map( A1 => n19619, A2 => n1173, Z => n31698);
   U26194 : AOI21_X2 port map( A1 => n26133, A2 => n2277, B => n31699, ZN => 
                           n2272);
   U26196 : OAI21_X2 port map( A1 => n26798, A2 => n28714, B => n3673, ZN => 
                           n31699);
   U26199 : XOR2_X1 port map( A1 => n10697, A2 => n23331, Z => n31703);
   U26202 : AOI22_X2 port map( A1 => n3113, A2 => n3112, B1 => n3111, B2 => 
                           n28573, ZN => n3340);
   U26205 : XOR2_X1 port map( A1 => n24521, A2 => n14920, Z => n31704);
   U26213 : XOR2_X1 port map( A1 => n31706, A2 => n31913, Z => n27792);
   U26220 : NAND2_X2 port map( A1 => n1256, A2 => n27219, ZN => n26716);
   U26221 : XOR2_X1 port map( A1 => n2900, A2 => n29463, Z => n26537);
   U26222 : XOR2_X1 port map( A1 => n22239, A2 => n22240, Z => n12898);
   U26229 : XOR2_X1 port map( A1 => n24489, A2 => n15744, Z => n15743);
   U26230 : INV_X2 port map( I => n24197, ZN => n27430);
   U26231 : NAND3_X2 port map( A1 => n26211, A2 => n23676, A3 => n23677, ZN => 
                           n24197);
   U26247 : OAI21_X1 port map( A1 => n15912, A2 => n11516, B => n29271, ZN => 
                           n8914);
   U26250 : NAND3_X2 port map( A1 => n31710, A2 => n18384, A3 => n17649, ZN => 
                           n3836);
   U26251 : NAND2_X2 port map( A1 => n18559, A2 => n18494, ZN => n11774);
   U26254 : XOR2_X1 port map( A1 => Plaintext(77), A2 => Key(77), Z => n18494);
   U26255 : BUF_X2 port map( I => n24847, Z => n31713);
   U26261 : NAND2_X2 port map( A1 => n31834, A2 => n31714, ZN => n20399);
   U26275 : NAND3_X1 port map( A1 => n24051, A2 => n14490, A3 => n4897, ZN => 
                           n305);
   U26279 : OAI22_X1 port map( A1 => n15857, A2 => n11998, B1 => n15855, B2 => 
                           n15854, ZN => n26295);
   U26281 : INV_X2 port map( I => n31716, ZN => n17516);
   U26284 : XOR2_X1 port map( A1 => Plaintext(126), A2 => Key(126), Z => n31716
                           );
   U26288 : NAND3_X2 port map( A1 => n31718, A2 => n24038, A3 => n24039, ZN => 
                           n24416);
   U26291 : XOR2_X1 port map( A1 => n24758, A2 => n31719, Z => n28968);
   U26292 : XOR2_X1 port map( A1 => n5539, A2 => n31720, Z => n31719);
   U26294 : INV_X1 port map( I => n16619, ZN => n31720);
   U26297 : OAI22_X2 port map( A1 => n19605, A2 => n29730, B1 => n2717, B2 => 
                           n19196, ZN => n1944);
   U26300 : NOR2_X2 port map( A1 => n3207, A2 => n19195, ZN => n19605);
   U26305 : INV_X2 port map( I => n736, ZN => n25539);
   U26314 : XOR2_X1 port map( A1 => n8617, A2 => n25156, Z => n610);
   U26321 : XOR2_X1 port map( A1 => n15130, A2 => n8762, Z => n27011);
   U26324 : NAND3_X2 port map( A1 => n28846, A2 => n7582, A3 => n22276, ZN => 
                           n15130);
   U26330 : XOR2_X1 port map( A1 => n27763, A2 => n23346, Z => n23498);
   U26335 : XOR2_X1 port map( A1 => n24405, A2 => n24404, Z => n31725);
   U26337 : INV_X2 port map( I => n8106, ZN => n31730);
   U26338 : AOI21_X2 port map( A1 => n31732, A2 => n21644, B => n3418, ZN => 
                           n22119);
   U26339 : NAND3_X2 port map( A1 => n29389, A2 => n31893, A3 => n5424, ZN => 
                           n5612);
   U26345 : AOI21_X2 port map( A1 => n31736, A2 => n29158, B => n3495, ZN => 
                           n7905);
   U26350 : NAND2_X2 port map( A1 => n31344, A2 => n9022, ZN => n31736);
   U26354 : XOR2_X1 port map( A1 => n31738, A2 => n31737, Z => n31787);
   U26355 : XOR2_X1 port map( A1 => n23277, A2 => n23234, Z => n31738);
   U26356 : OR2_X1 port map( A1 => n421, A2 => n6581, Z => n26204);
   U26373 : XOR2_X1 port map( A1 => n31739, A2 => n25908, Z => Ciphertext(187))
                           ;
   U26377 : OAI22_X1 port map( A1 => n7716, A2 => n25907, B1 => n25927, B2 => 
                           n690, ZN => n31739);
   U26378 : OAI22_X1 port map( A1 => n1094, A2 => n24044, B1 => n23602, B2 => 
                           n13412, ZN => n26966);
   U26388 : AOI22_X2 port map( A1 => n28491, A2 => n6453, B1 => n23111, B2 => 
                           n853, ZN => n5893);
   U26390 : NAND2_X2 port map( A1 => n28003, A2 => n9080, ZN => n16429);
   U26391 : NOR2_X1 port map( A1 => n11923, A2 => n6479, ZN => n7444);
   U26392 : XNOR2_X1 port map( A1 => n9185, A2 => n32861, ZN => n16382);
   U26394 : AND2_X1 port map( A1 => n5034, A2 => n28157, Z => n19238);
   U26399 : NOR2_X1 port map( A1 => n20052, A2 => n13327, ZN => n31745);
   U26403 : XOR2_X1 port map( A1 => n31747, A2 => n16125, Z => n3339);
   U26404 : NOR2_X2 port map( A1 => n31748, A2 => n15808, ZN => n11744);
   U26414 : XOR2_X1 port map( A1 => n8809, A2 => n31749, Z => n8302);
   U26416 : XOR2_X1 port map( A1 => n26230, A2 => n19755, Z => n8809);
   U26418 : NAND2_X2 port map( A1 => n20379, A2 => n6679, ZN => n11303);
   U26424 : AND2_X1 port map( A1 => n636, A2 => n1119, Z => n28902);
   U26426 : XOR2_X1 port map( A1 => n1590, A2 => n1587, Z => n1589);
   U26430 : OAI21_X1 port map( A1 => n31954, A2 => n2386, B => n423, ZN => 
                           n21644);
   U26434 : NAND2_X2 port map( A1 => n6629, A2 => n12163, ZN => n7555);
   U26440 : XOR2_X1 port map( A1 => n17554, A2 => n20836, Z => n20957);
   U26442 : OAI22_X2 port map( A1 => n20048, A2 => n20047, B1 => n20546, B2 => 
                           n28904, ZN => n20836);
   U26443 : XOR2_X1 port map( A1 => n31751, A2 => n15470, Z => n15092);
   U26446 : XOR2_X1 port map( A1 => n22222, A2 => n22049, Z => n9701);
   U26447 : XOR2_X1 port map( A1 => n21913, A2 => n31457, Z => n22049);
   U26449 : INV_X2 port map( I => n31753, ZN => n26040);
   U26450 : XOR2_X1 port map( A1 => Plaintext(25), A2 => Key(25), Z => n31753);
   U26451 : XOR2_X1 port map( A1 => n21481, A2 => n31105, Z => n31754);
   U26452 : AOI21_X2 port map( A1 => n26253, A2 => n13129, B => n3659, ZN => 
                           n3658);
   U26454 : XOR2_X1 port map( A1 => n2384, A2 => n5647, Z => n31756);
   U26456 : NAND2_X2 port map( A1 => n18405, A2 => n3051, ZN => n3060);
   U26458 : XOR2_X1 port map( A1 => n16838, A2 => n31761, Z => n188);
   U26459 : XOR2_X1 port map( A1 => n31762, A2 => n28898, Z => n31761);
   U26460 : NAND2_X1 port map( A1 => n31763, A2 => n9558, ZN => n26431);
   U26461 : NOR2_X1 port map( A1 => n26142, A2 => n5395, ZN => n31763);
   U26462 : XOR2_X1 port map( A1 => n10789, A2 => n10788, Z => n27732);
   U26466 : NAND2_X2 port map( A1 => n5645, A2 => n31767, ZN => n7345);
   U26467 : AOI22_X2 port map( A1 => n5644, A2 => n18571, B1 => n953, B2 => 
                           n485, ZN => n31767);
   U26468 : AOI22_X1 port map( A1 => n1757, A2 => n1758, B1 => n1756, B2 => 
                           n13023, ZN => n28116);
   U26469 : XOR2_X1 port map( A1 => n21041, A2 => n4021, Z => n31769);
   U26470 : XOR2_X1 port map( A1 => n31770, A2 => n6940, Z => n6938);
   U26471 : XOR2_X1 port map( A1 => n24692, A2 => n24376, Z => n31770);
   U26472 : XOR2_X1 port map( A1 => n22171, A2 => n17258, Z => n16861);
   U26473 : XOR2_X1 port map( A1 => n31771, A2 => n8020, Z => n17721);
   U26475 : NAND2_X1 port map( A1 => n9249, A2 => n9248, ZN => n9251);
   U26479 : XOR2_X1 port map( A1 => n1851, A2 => n6574, Z => n29228);
   U26480 : XOR2_X1 port map( A1 => n18398, A2 => Key(184), Z => n31773);
   U26484 : NOR2_X2 port map( A1 => n28836, A2 => n6530, ZN => n31776);
   U26486 : NAND2_X2 port map( A1 => n10656, A2 => n10655, ZN => n9076);
   U26490 : OAI21_X2 port map( A1 => n12029, A2 => n16484, B => n4518, ZN => 
                           n31777);
   U26491 : NOR2_X2 port map( A1 => n18266, A2 => n18265, ZN => n4858);
   U26492 : OAI22_X2 port map( A1 => n20426, A2 => n12421, B1 => n20428, B2 => 
                           n32747, ZN => n18265);
   U26493 : NAND2_X2 port map( A1 => n31780, A2 => n31778, ZN => n25136);
   U26495 : OAI21_X2 port map( A1 => n7969, A2 => n196, B => n31960, ZN => 
                           n31781);
   U26496 : BUF_X2 port map( I => n16267, Z => n31784);
   U26497 : INV_X2 port map( I => n4036, ZN => n10579);
   U26498 : XOR2_X1 port map( A1 => Plaintext(29), A2 => Key(29), Z => n4036);
   U26499 : AOI21_X2 port map( A1 => n25523, A2 => n27236, B => n31786, ZN => 
                           n25369);
   U26500 : INV_X2 port map( I => n13113, ZN => n16386);
   U26502 : INV_X2 port map( I => n31787, ZN => n23834);
   U26503 : OAI22_X1 port map( A1 => n25380, A2 => n25379, B1 => n25377, B2 => 
                           n30302, ZN => n27487);
   U26504 : AOI21_X1 port map( A1 => n18459, A2 => n956, B => n16854, ZN => 
                           n7163);
   U26505 : INV_X2 port map( I => n17261, ZN => n24265);
   U26506 : NAND2_X2 port map( A1 => n12774, A2 => n26967, ZN => n17261);
   U26508 : NOR2_X2 port map( A1 => n28974, A2 => n31790, ZN => n28782);
   U26509 : XOR2_X1 port map( A1 => n19660, A2 => n29341, Z => n26003);
   U26512 : INV_X2 port map( I => n22949, ZN => n31795);
   U26513 : NAND2_X2 port map( A1 => n6733, A2 => n19840, ZN => n20431);
   U26514 : INV_X2 port map( I => n31797, ZN => n26078);
   U26515 : NAND2_X1 port map( A1 => n26817, A2 => n14625, ZN => n31799);
   U26516 : XOR2_X1 port map( A1 => n31800, A2 => n19443, Z => n28216);
   U26517 : XOR2_X1 port map( A1 => n27444, A2 => n7057, Z => n31800);
   U26521 : XOR2_X1 port map( A1 => n24602, A2 => n31803, Z => n7535);
   U26522 : XOR2_X1 port map( A1 => n25991, A2 => n7828, Z => n31803);
   U26526 : NAND2_X2 port map( A1 => n5418, A2 => n4191, ZN => n26683);
   U26529 : XOR2_X1 port map( A1 => n19543, A2 => n19702, Z => n7375);
   U26530 : OAI22_X2 port map( A1 => n229, A2 => n15920, B1 => n15919, B2 => 
                           n16724, ZN => n31824);
   U26534 : OAI21_X2 port map( A1 => n2744, A2 => n32298, B => n14663, ZN => 
                           n31813);
   U26535 : OAI21_X2 port map( A1 => n18141, A2 => n20142, B => n1458, ZN => 
                           n31814);
   U26543 : INV_X2 port map( I => n31819, ZN => n18960);
   U26544 : NOR2_X2 port map( A1 => n4747, A2 => n12585, ZN => n31819);
   U26545 : NAND2_X2 port map( A1 => n6750, A2 => n6749, ZN => n15829);
   U26546 : NOR2_X2 port map( A1 => n31820, A2 => n29602, ZN => n448);
   U26547 : INV_X2 port map( I => n25892, ZN => n31822);
   U26548 : OAI21_X1 port map( A1 => n773, A2 => n22945, B => n31825, ZN => 
                           n8923);
   U26550 : NOR2_X1 port map( A1 => n16832, A2 => n18977, ZN => n5842);
   U26552 : XOR2_X1 port map( A1 => n19671, A2 => n17689, Z => n26738);
   U26553 : AOI22_X2 port map( A1 => n31827, A2 => n1055, B1 => n4749, B2 => 
                           n28478, ZN => n11777);
   U26554 : OAI21_X2 port map( A1 => n1175, A2 => n1051, B => n25961, ZN => 
                           n31827);
   U26558 : NOR2_X2 port map( A1 => n31830, A2 => n29094, ZN => n1474);
   U26559 : NOR2_X1 port map( A1 => n19601, A2 => n10860, ZN => n19614);
   U26561 : NAND2_X2 port map( A1 => n28844, A2 => n20182, ZN => n20775);
   U26562 : XOR2_X1 port map( A1 => n9586, A2 => n17538, Z => n3982);
   U26564 : XOR2_X1 port map( A1 => n13586, A2 => n4329, Z => n27152);
   U26567 : NOR2_X1 port map( A1 => n5786, A2 => n12885, ZN => n31833);
   U26571 : OAI21_X2 port map( A1 => n31836, A2 => n16184, B => n8539, ZN => 
                           n21498);
   U26572 : NOR2_X2 port map( A1 => n31030, A2 => n1333, ZN => n31836);
   U26573 : NAND2_X2 port map( A1 => n31923, A2 => n12610, ZN => n5602);
   U26575 : XOR2_X1 port map( A1 => n19409, A2 => n17551, Z => n19732);
   U26576 : INV_X2 port map( I => n31839, ZN => n9910);
   U26579 : AOI21_X2 port map( A1 => n26591, A2 => n18729, B => n31980, ZN => 
                           n25971);
   U26580 : NOR2_X2 port map( A1 => n13616, A2 => n13615, ZN => n13614);
   U26583 : NOR2_X1 port map( A1 => n17669, A2 => n23087, ZN => n17668);
   U26586 : XOR2_X1 port map( A1 => n9674, A2 => n31841, Z => n28607);
   U26587 : XOR2_X1 port map( A1 => n22171, A2 => n16027, Z => n27312);
   U26588 : XOR2_X1 port map( A1 => n6689, A2 => n6686, Z => n10248);
   U26590 : XOR2_X1 port map( A1 => n22113, A2 => n22196, Z => n22289);
   U26591 : BUF_X2 port map( I => n3504, Z => n31843);
   U26592 : XOR2_X1 port map( A1 => n31844, A2 => n5846, Z => n5844);
   U26594 : XOR2_X1 port map( A1 => n19470, A2 => n27607, Z => n5925);
   U26599 : XOR2_X1 port map( A1 => n31849, A2 => n24539, Z => n29277);
   U26603 : NAND2_X2 port map( A1 => n3045, A2 => n3047, ZN => n22227);
   U26607 : XOR2_X1 port map( A1 => n3209, A2 => n2661, Z => n31852);
   U26608 : NAND2_X2 port map( A1 => n3211, A2 => n31853, ZN => n21779);
   U26612 : AOI22_X2 port map( A1 => n14828, A2 => n16915, B1 => n18464, B2 => 
                           n18489, ZN => n31856);
   U26613 : NAND3_X2 port map( A1 => n1772, A2 => n26979, A3 => n615, ZN => 
                           n29137);
   U26616 : NAND2_X2 port map( A1 => n13850, A2 => n12228, ZN => n13041);
   U26619 : XOR2_X1 port map( A1 => n23333, A2 => n1260, Z => n23128);
   U26620 : OAI21_X1 port map( A1 => n964, A2 => n713, B => n7941, ZN => n5903)
                           ;
   U26621 : XOR2_X1 port map( A1 => n12258, A2 => n29832, Z => n26920);
   U26622 : OAI21_X2 port map( A1 => n4497, A2 => n4496, B => n26152, ZN => 
                           n12211);
   U26623 : XOR2_X1 port map( A1 => n14407, A2 => n13299, Z => n4572);
   U26624 : NOR2_X2 port map( A1 => n18699, A2 => n22, ZN => n18833);
   U26625 : INV_X1 port map( I => n15139, ZN => n18699);
   U26626 : XOR2_X1 port map( A1 => n18388, A2 => Key(111), Z => n15139);
   U26627 : XOR2_X1 port map( A1 => n22284, A2 => n22003, Z => n1762);
   U26628 : BUF_X2 port map( I => n24616, Z => n31866);
   U26631 : XOR2_X1 port map( A1 => n9092, A2 => n9093, Z => n31869);
   U26632 : NAND3_X2 port map( A1 => n14838, A2 => n24344, A3 => n24342, ZN => 
                           n24531);
   U26636 : NAND2_X2 port map( A1 => n9561, A2 => n24084, ZN => n24137);
   U26637 : NAND2_X2 port map( A1 => n3170, A2 => n3172, ZN => n7772);
   U26638 : NAND2_X1 port map( A1 => n17535, A2 => n11957, ZN => n24730);
   U26639 : AND2_X1 port map( A1 => n23717, A2 => n10967, Z => n23682);
   U26640 : NAND2_X2 port map( A1 => n3845, A2 => n23999, ZN => n24533);
   U26642 : XOR2_X1 port map( A1 => n5194, A2 => n31875, Z => n27883);
   U26644 : AOI21_X1 port map( A1 => n25044, A2 => n31876, B => n25062, ZN => 
                           n8258);
   U26645 : NAND2_X1 port map( A1 => n25058, A2 => n25057, ZN => n31876);
   U26646 : OAI21_X1 port map( A1 => n3229, A2 => n2983, B => n14865, ZN => 
                           n2264);
   U26647 : NOR2_X1 port map( A1 => n20276, A2 => n14187, ZN => n20277);
   U26648 : XOR2_X1 port map( A1 => n6421, A2 => n31880, Z => n25146);
   U26649 : XOR2_X1 port map( A1 => n24840, A2 => n29417, Z => n31880);
   U26654 : OAI21_X2 port map( A1 => n11693, A2 => n17843, B => n31885, ZN => 
                           n18658);
   U26655 : NAND2_X2 port map( A1 => n17843, A2 => n18446, ZN => n31885);
   U26657 : XOR2_X1 port map( A1 => n5184, A2 => n29412, Z => n31887);
   U26658 : NAND2_X1 port map( A1 => n31888, A2 => n16083, ZN => n2729);
   U26659 : NOR2_X1 port map( A1 => n23620, A2 => n30360, ZN => n31888);
   U26660 : XOR2_X1 port map( A1 => n20802, A2 => n25266, Z => n7595);
   U26661 : OAI22_X2 port map( A1 => n9587, A2 => n9588, B1 => n20075, B2 => 
                           n20360, ZN => n20802);
   U26662 : BUF_X2 port map( I => n10312, Z => n31891);
   U26664 : XOR2_X1 port map( A1 => n28753, A2 => n23518, Z => n31892);
   U26665 : NOR2_X1 port map( A1 => n21848, A2 => n30291, ZN => n12852);
   U26666 : AOI21_X2 port map( A1 => n5611, A2 => n1216, B => n31895, ZN => 
                           n28304);
   U26667 : AOI21_X2 port map( A1 => n8031, A2 => n7577, B => n31898, ZN => 
                           n7157);
   U26669 : XOR2_X1 port map( A1 => n24573, A2 => n25991, Z => n31899);
   U26673 : XOR2_X1 port map( A1 => n26540, A2 => n24402, Z => n31901);
   U26677 : NAND2_X1 port map( A1 => n7334, A2 => n32859, ZN => n31904);
   U26680 : XOR2_X1 port map( A1 => n26075, A2 => n4771, Z => n392);
   U26681 : XOR2_X1 port map( A1 => n20849, A2 => n6857, Z => n4771);
   U26682 : XOR2_X1 port map( A1 => n19577, A2 => n19578, Z => n4465);
   U26683 : INV_X2 port map( I => n19958, ZN => n27808);
   U26684 : INV_X1 port map( I => n26088, ZN => n20090);
   U26686 : INV_X2 port map( I => n26194, ZN => n505);
   U26688 : NOR2_X2 port map( A1 => n13314, A2 => n13310, ZN => n21122);
   U26689 : NAND2_X2 port map( A1 => n27249, A2 => n28549, ZN => n28232);
   U26690 : XNOR2_X1 port map( A1 => n22067, A2 => n16482, ZN => n31912);
   U26691 : XNOR2_X1 port map( A1 => n6771, A2 => n10935, ZN => n31913);
   U26692 : INV_X2 port map( I => n3536, ZN => n22491);
   U26694 : INV_X1 port map( I => n9953, ZN => n11804);
   U26695 : INV_X1 port map( I => n6407, ZN => n22362);
   U4340 : AND2_X1 port map( A1 => n27077, A2 => n30010, Z => n1490);
   U1051 : INV_X2 port map( I => n21704, ZN => n26782);
   U1695 : NAND2_X2 port map( A1 => n10323, A2 => n15434, ZN => n7961);
   U5747 : AOI21_X2 port map( A1 => n8022, A2 => n1271, B => n12220, ZN => 
                           n9918);
   U14047 : INV_X4 port map( I => n20052, ZN => n19949);
   U3960 : BUF_X4 port map( I => n7251, Z => n29223);
   U1145 : INV_X2 port map( I => n13712, ZN => n26735);
   U1873 : INV_X2 port map( I => n26699, ZN => n29200);
   U5133 : INV_X2 port map( I => n4289, ZN => n20575);
   U5403 : INV_X2 port map( I => n17237, ZN => n20570);
   U1119 : INV_X2 port map( I => n11063, ZN => n15002);
   U15357 : NOR2_X2 port map( A1 => n4665, A2 => n4664, ZN => n4329);
   U3390 : INV_X2 port map( I => n18487, ZN => n26520);
   U15563 : NAND3_X2 port map( A1 => n23828, A2 => n23953, A3 => n13281, ZN => 
                           n4824);
   U7038 : INV_X2 port map( I => n9871, ZN => n22503);
   U5912 : NAND2_X2 port map( A1 => n29365, A2 => n19826, ZN => n30748);
   U8233 : NAND2_X2 port map( A1 => n21107, A2 => n10546, ZN => n21510);
   U2384 : NAND3_X2 port map( A1 => n20949, A2 => n5822, A3 => n29062, ZN => 
                           n20950);
   U867 : BUF_X4 port map( I => n17201, Z => n29222);
   U14806 : OR2_X2 port map( A1 => n6407, A2 => n11805, Z => n12869);
   U121 : NAND3_X2 port map( A1 => n11306, A2 => n25565, A3 => n11900, ZN => 
                           n2018);
   U54 : INV_X2 port map( I => n25686, ZN => n29243);
   U2203 : INV_X2 port map( I => n21761, ZN => n21847);
   U23123 : NAND3_X2 port map( A1 => n20178, A2 => n20179, A3 => n33301, ZN => 
                           n20182);
   U3531 : INV_X2 port map( I => n10170, ZN => n25695);
   U1425 : NAND2_X2 port map( A1 => n18035, A2 => n10679, ZN => n26848);
   U10624 : INV_X2 port map( I => n24235, ZN => n10627);
   U4438 : INV_X4 port map( I => n561, ZN => n1083);
   U11379 : OR2_X2 port map( A1 => n21350, A2 => n30389, Z => n21571);
   U17315 : AOI21_X2 port map( A1 => n14473, A2 => n16943, B => n4891, ZN => 
                           n27446);
   U21045 : NAND2_X2 port map( A1 => n981, A2 => n8217, ZN => n16943);
   U6595 : NOR2_X2 port map( A1 => n31108, A2 => n19052, ZN => n3092);
   U1587 : BUF_X4 port map( I => n25185, Z => n15641);
   U17991 : BUF_X4 port map( I => n10292, Z => n30571);
   U4868 : NOR3_X2 port map( A1 => n2296, A2 => n34046, A3 => n1322, ZN => 
                           n2339);
   U21491 : INV_X2 port map( I => n19244, ZN => n14698);
   U3667 : NAND2_X2 port map( A1 => n30010, A2 => n4202, ZN => n19244);
   U4859 : NAND2_X2 port map( A1 => n1322, A2 => n34046, ZN => n21830);
   U14769 : INV_X2 port map( I => n24147, ZN => n24120);
   U2978 : NAND2_X2 port map( A1 => n19234, A2 => n29003, ZN => n8119);
   U5167 : OR2_X1 port map( A1 => n8933, A2 => n4881, Z => n11785);
   U1690 : NAND2_X2 port map( A1 => n13920, A2 => n26881, ZN => n9364);
   U4967 : INV_X4 port map( I => n19249, ZN => n16274);
   U6141 : INV_X2 port map( I => n470, ZN => n31670);
   U26023 : AND2_X2 port map( A1 => n2207, A2 => n15411, Z => n12316);
   U1603 : INV_X2 port map( I => n16122, ZN => n27909);
   U13418 : NOR2_X2 port map( A1 => n7673, A2 => n1333, ZN => n26997);
   U5917 : NOR2_X2 port map( A1 => n2606, A2 => n16630, ZN => n20060);
   U15425 : BUF_X4 port map( I => n16453, Z => n7557);
   U14180 : NAND2_X2 port map( A1 => n16374, A2 => n9352, ZN => n10231);
   U23171 : NOR2_X2 port map( A1 => n9895, A2 => n8331, ZN => n22048);
   U3316 : INV_X2 port map( I => n10285, ZN => n25739);
   U16585 : INV_X4 port map( I => n13413, ZN => n23756);
   U150 : BUF_X2 port map( I => n18242, Z => n30512);
   U3433 : INV_X2 port map( I => n7280, ZN => n7279);
   U3187 : NAND2_X2 port map( A1 => n7195, A2 => n9663, ZN => n9664);
   U10260 : NAND2_X2 port map( A1 => n7044, A2 => n26777, ZN => n21214);
   U3464 : NAND2_X2 port map( A1 => n15179, A2 => n24254, ZN => n13378);
   U6410 : AOI21_X2 port map( A1 => n31765, A2 => n33139, B => n17139, ZN => 
                           n2741);
   U2405 : OAI21_X2 port map( A1 => n12113, A2 => n10085, B => n30512, ZN => 
                           n14579);
   U4135 : NAND2_X2 port map( A1 => n7486, A2 => n16374, ZN => n28167);
   U23081 : NOR2_X2 port map( A1 => n27336, A2 => n15026, ZN => n21612);
   U6334 : INV_X4 port map( I => n22599, ZN => n9580);
   U6036 : BUF_X2 port map( I => n27698, Z => n29339);
   U2902 : NAND2_X2 port map( A1 => n3077, A2 => n30191, ZN => n24270);
   U4665 : INV_X2 port map( I => n25615, ZN => n1202);
   U12698 : OAI22_X2 port map( A1 => n3779, A2 => n18511, B1 => n12327, B2 => 
                           n11380, ZN => n17130);
   U7845 : NOR2_X2 port map( A1 => n29518, A2 => n12094, ZN => n29138);
   U3069 : OAI21_X2 port map( A1 => n22866, A2 => n23068, B => n10641, ZN => 
                           n12529);
   U15717 : NOR2_X2 port map( A1 => n18791, A2 => n13548, ZN => n9511);
   U14677 : NAND2_X2 port map( A1 => n21702, A2 => n33833, ZN => n6764);
   U299 : AOI21_X2 port map( A1 => n11236, A2 => n32176, B => n10381, ZN => 
                           n3678);
   U3269 : NAND2_X2 port map( A1 => n28338, A2 => n25756, ZN => n25875);
   U3048 : BUF_X4 port map( I => n15715, Z => n5471);
   U44 : INV_X2 port map( I => n32063, ZN => n26198);
   U2804 : INV_X2 port map( I => n25897, ZN => n27118);
   U15211 : AOI21_X2 port map( A1 => n26185, A2 => n14463, B => n33103, ZN => 
                           n30625);
   U9307 : NOR2_X2 port map( A1 => n22747, A2 => n1278, ZN => n12220);
   U11090 : NAND2_X1 port map( A1 => n15007, A2 => n1125, ZN => n9451);
   U7167 : NOR2_X2 port map( A1 => n1703, A2 => n32452, ZN => n21161);
   U2078 : INV_X4 port map( I => n23085, ZN => n17639);
   U3302 : INV_X4 port map( I => n25620, ZN => n8186);
   U14727 : NAND2_X2 port map( A1 => n28081, A2 => n32032, ZN => n27113);
   U18939 : INV_X4 port map( I => n29200, ZN => n30692);
   U1670 : BUF_X4 port map( I => n14564, Z => n4468);
   U1323 : NAND2_X2 port map( A1 => n19063, A2 => n19108, ZN => n19365);
   U265 : BUF_X2 port map( I => n10170, Z => n4146);
   U1579 : AOI22_X2 port map( A1 => n9668, A2 => n9667, B1 => n11098, B2 => 
                           n1182, ZN => n10481);
   U8820 : INV_X4 port map( I => n470, ZN => n14213);
   U807 : INV_X2 port map( I => n7024, ZN => n16225);
   U5354 : OAI21_X2 port map( A1 => n13127, A2 => n31934, B => n22444, ZN => 
                           n17462);
   U1040 : INV_X2 port map( I => n156, ZN => n13371);
   U4484 : AND2_X1 port map( A1 => n18037, A2 => n8964, Z => n22536);
   U1800 : INV_X2 port map( I => n19423, ZN => n4942);
   U2549 : BUF_X2 port map( I => n24682, Z => n27385);
   U1217 : BUF_X4 port map( I => n12211, Z => n1008);
   U5227 : INV_X2 port map( I => n29272, ZN => n980);
   U800 : NAND3_X2 port map( A1 => n31506, A2 => n22488, A3 => n22489, ZN => 
                           n10832);
   U2279 : INV_X2 port map( I => n713, ZN => n314);
   U639 : OAI21_X2 port map( A1 => n10895, A2 => n22900, B => n3830, ZN => 
                           n31758);
   U4046 : INV_X4 port map( I => n17184, ZN => n957);
   U14889 : NOR2_X2 port map( A1 => n23085, A2 => n23087, ZN => n22967);
   U5182 : NAND2_X2 port map( A1 => n16435, A2 => n18602, ZN => n15909);
   U17651 : NOR2_X2 port map( A1 => n10085, A2 => n7963, ZN => n25839);
   U4881 : INV_X4 port map( I => n9220, ZN => n12143);
   U6555 : AOI21_X2 port map( A1 => n12912, A2 => n12911, B => n810, ZN => 
                           n26595);
   U8503 : NAND2_X2 port map( A1 => n4639, A2 => n19883, ZN => n4638);
   U26384 : NAND2_X2 port map( A1 => n12257, A2 => n24873, ZN => n8777);
   U1360 : NOR2_X2 port map( A1 => n21839, A2 => n27937, ZN => n13030);
   U4400 : BUF_X4 port map( I => n33146, Z => n3468);
   U4761 : AND2_X1 port map( A1 => n28329, A2 => n9430, Z => n10045);
   U21161 : OAI21_X1 port map( A1 => n12831, A2 => n12707, B => n18922, ZN => 
                           n12830);
   U1809 : AND2_X2 port map( A1 => n2499, A2 => n12379, Z => n20079);
   U7587 : INV_X2 port map( I => n15146, ZN => n18892);
   U20711 : INV_X2 port map( I => n11677, ZN => n12037);
   U6718 : NOR2_X2 port map( A1 => n22666, A2 => n22664, ZN => n26406);
   U3993 : INV_X2 port map( I => n12044, ZN => n21406);
   U2725 : INV_X2 port map( I => n25295, ZN => n25398);
   U3686 : INV_X2 port map( I => n25429, ZN => n25453);
   U2727 : NAND2_X2 port map( A1 => n25295, A2 => n25397, ZN => n27586);
   U3437 : INV_X2 port map( I => n16534, ZN => n842);
   U10878 : NAND3_X2 port map( A1 => n13251, A2 => n1108, A3 => n1109, ZN => 
                           n16928);
   U943 : NAND2_X2 port map( A1 => n3567, A2 => n30529, ZN => n11202);
   U2930 : INV_X2 port map( I => n31965, ZN => n1017);
   U24696 : INV_X2 port map( I => n20614, ZN => n20392);
   U20610 : INV_X2 port map( I => n18873, ZN => n11460);
   U207 : INV_X2 port map( I => n6286, ZN => n1239);
   U11504 : NAND2_X2 port map( A1 => n28860, A2 => n28635, ZN => n26682);
   U6767 : OAI22_X2 port map( A1 => n27415, A2 => n16149, B1 => n22664, B2 => 
                           n16567, ZN => n28860);
   U5310 : NOR2_X2 port map( A1 => n23949, A2 => n11676, ZN => n11708);
   U4052 : AND2_X1 port map( A1 => n12211, A2 => n30690, Z => n31335);
   U8815 : NAND2_X2 port map( A1 => n15956, A2 => n13738, ZN => n18463);
   U5046 : INV_X2 port map( I => n9375, ZN => n23576);
   U6079 : NAND2_X2 port map( A1 => n10126, A2 => n10127, ZN => n6504);
   U4373 : NAND2_X2 port map( A1 => n25142, A2 => n25184, ZN => n25170);
   U15083 : INV_X4 port map( I => n13693, ZN => n125);
   U25336 : NAND3_X2 port map( A1 => n14973, A2 => n23785, A3 => n23903, ZN => 
                           n23710);
   U22375 : AOI21_X2 port map( A1 => n10700, A2 => n19115, B => n25968, ZN => 
                           n15143);
   U12873 : NAND2_X1 port map( A1 => n16904, A2 => n17405, ZN => n30064);
   U12242 : INV_X1 port map( I => n16904, ZN => n29981);
   U6760 : NAND2_X2 port map( A1 => n33761, A2 => n9427, ZN => n9426);
   U3799 : NAND2_X2 port map( A1 => n22364, A2 => n1125, ZN => n3970);
   U3349 : NOR2_X2 port map( A1 => n13796, A2 => n32253, ZN => n29962);
   U15551 : INV_X2 port map( I => n17361, ZN => n13950);
   U10530 : NOR2_X2 port map( A1 => n10667, A2 => n10666, ZN => n6490);
   U7411 : NOR2_X2 port map( A1 => n29218, A2 => n30360, ZN => n26241);
   U16285 : OAI22_X2 port map( A1 => n5266, A2 => n18743, B1 => n18744, B2 => 
                           n18745, ZN => n27261);
   U869 : INV_X2 port map( I => n575, ZN => n1170);
   U6762 : NOR2_X2 port map( A1 => n16432, A2 => n11930, ZN => n1669);
   U254 : INV_X2 port map( I => n24308, ZN => n27739);
   U281 : AOI21_X2 port map( A1 => n24230, A2 => n24228, B => n30696, ZN => 
                           n30695);
   U1191 : INV_X2 port map( I => n21044, ZN => n8284);
   U10844 : OAI21_X2 port map( A1 => n6148, A2 => n26609, B => n26608, ZN => 
                           n26607);
   U15376 : AOI21_X2 port map( A1 => n28900, A2 => n3487, B => n28899, ZN => 
                           n8285);
   U3869 : INV_X2 port map( I => n8084, ZN => n27537);
   U9191 : NOR2_X2 port map( A1 => n17288, A2 => n17287, ZN => n17286);
   U4878 : INV_X2 port map( I => n32108, ZN => n16403);
   U4448 : BUF_X4 port map( I => n25112, Z => n25235);
   U977 : INV_X2 port map( I => n9737, ZN => n31344);
   U6479 : INV_X4 port map( I => n12966, ZN => n20427);
   U1458 : OAI21_X2 port map( A1 => n11655, A2 => n27828, B => n1331, ZN => 
                           n30972);
   U17361 : INV_X4 port map( I => n11820, ZN => n15964);
   U48 : INV_X1 port map( I => n10285, ZN => n27164);
   U12754 : AOI21_X2 port map( A1 => n6951, A2 => n32559, B => n26827, ZN => 
                           n6950);
   U1904 : INV_X2 port map( I => n19215, ZN => n31503);
   U1288 : NAND2_X2 port map( A1 => n15027, A2 => n20463, ZN => n11035);
   U19235 : INV_X2 port map( I => n12866, ZN => n21733);
   U10119 : NOR3_X2 port map( A1 => n16358, A2 => n5269, A3 => n18705, ZN => 
                           n10833);
   U3671 : NAND2_X2 port map( A1 => n21579, A2 => n6669, ZN => n21659);
   U5990 : INV_X1 port map( I => n16855, ZN => n1183);
   U7369 : NAND2_X2 port map( A1 => n17675, A2 => n9749, ZN => n4639);
   U8788 : NOR2_X2 port map( A1 => n5269, A2 => n18746, ZN => n5266);
   U6865 : INV_X2 port map( I => n26415, ZN => n23794);
   U18021 : NAND2_X1 port map( A1 => n7067, A2 => n969, ZN => n7069);
   U6855 : INV_X2 port map( I => n9153, ZN => n10052);
   U4808 : INV_X4 port map( I => n11923, ZN => n739);
   U4669 : NAND2_X2 port map( A1 => n18983, A2 => n27021, ZN => n18965);
   U9972 : INV_X2 port map( I => n19436, ZN => n3417);
   U15096 : NOR2_X2 port map( A1 => n7081, A2 => n25339, ZN => n25233);
   U12100 : NAND2_X1 port map( A1 => n18887, A2 => n10326, ZN => n6362);
   U11820 : NAND2_X2 port map( A1 => n12625, A2 => n31742, ZN => n9728);
   U5745 : AOI21_X2 port map( A1 => n7946, A2 => n29325, B => n27589, ZN => 
                           n7945);
   U5909 : OAI21_X2 port map( A1 => n11832, A2 => n15052, B => n14913, ZN => 
                           n11831);
   U1993 : NAND2_X2 port map( A1 => n19265, A2 => n18973, ZN => n26469);
   U2762 : NAND2_X2 port map( A1 => n24609, A2 => n28815, ZN => n15232);
   U4982 : BUF_X2 port map( I => n19583, Z => n27240);
   U2387 : BUF_X4 port map( I => n14002, Z => n4135);
   U2455 : NAND3_X1 port map( A1 => n16582, A2 => n16583, A3 => n7871, ZN => 
                           n26877);
   U2991 : INV_X2 port map( I => n12561, ZN => n919);
   U7098 : OR2_X1 port map( A1 => n28904, A2 => n20545, Z => n29356);
   U3375 : NOR2_X2 port map( A1 => n23766, A2 => n23736, ZN => n28637);
   U462 : OR2_X2 port map( A1 => n5736, A2 => n9828, Z => n29372);
   U1104 : NAND2_X2 port map( A1 => n26573, A2 => n26513, ZN => n31400);
   U25118 : OAI21_X1 port map( A1 => n14251, A2 => n32830, B => n22350, ZN => 
                           n22650);
   U6 : NAND2_X2 port map( A1 => n2962, A2 => n5839, ZN => n25732);
   U7766 : AOI21_X2 port map( A1 => n14491, A2 => n14703, B => n28945, ZN => 
                           n3257);
   U3368 : INV_X2 port map( I => n13862, ZN => n1299);
   U4430 : INV_X1 port map( I => n18059, ZN => n25227);
   U6126 : INV_X4 port map( I => n9561, ZN => n14913);
   U6798 : BUF_X4 port map( I => n9107, Z => n30365);
   U4281 : BUF_X2 port map( I => Key(157), Z => n16525);
   U4292 : BUF_X2 port map( I => Key(36), Z => n16497);
   U18780 : NAND2_X1 port map( A1 => n16607, A2 => n25120, ZN => n30673);
   U370 : NAND2_X2 port map( A1 => n31531, A2 => n4124, ZN => n2114);
   U6558 : INV_X4 port map( I => n15522, ZN => n11745);
   U3541 : OAI21_X2 port map( A1 => n14699, A2 => n14698, B => n19245, ZN => 
                           n14697);
   U6203 : NAND3_X2 port map( A1 => n1057, A2 => n3928, A3 => n3927, ZN => 
                           n5155);
   U7331 : INV_X2 port map( I => n20413, ZN => n933);
   U610 : INV_X2 port map( I => n12878, ZN => n13321);
   U5973 : INV_X2 port map( I => n18859, ZN => n1057);
   U2969 : AOI21_X2 port map( A1 => n16308, A2 => n14556, B => n1022, ZN => 
                           n20249);
   U11643 : NAND2_X2 port map( A1 => n28899, A2 => n20362, ZN => n20364);
   U8355 : INV_X2 port map( I => n599, ZN => n21324);
   U15762 : OR2_X2 port map( A1 => n23587, A2 => n23130, Z => n8145);
   U4048 : AND2_X1 port map( A1 => n17184, A2 => n17030, Z => n18850);
   U3258 : NAND2_X2 port map( A1 => n33909, A2 => n6961, ZN => n9413);
   U23948 : NAND2_X2 port map( A1 => n26573, A2 => n21687, ZN => n12562);
   U16155 : NOR2_X2 port map( A1 => n12320, A2 => n18581, ZN => n30560);
   U7043 : INV_X4 port map( I => n7831, ZN => n4525);
   U8273 : NOR2_X2 port map( A1 => n8197, A2 => n154, ZN => n15931);
   U3438 : OAI22_X2 port map( A1 => n773, A2 => n9954, B1 => n22945, B2 => n850
                           , ZN => n26253);
   U2133 : NOR2_X1 port map( A1 => n30619, A2 => n4220, ZN => n12753);
   U237 : INV_X2 port map( I => n25890, ZN => n7689);
   U5090 : NAND2_X2 port map( A1 => n18078, A2 => n6679, ZN => n1469);
   U15596 : INV_X2 port map( I => n21240, ZN => n2239);
   U25834 : OAI21_X2 port map( A1 => n17791, A2 => n20278, B => n17790, ZN => 
                           n28829);
   U23973 : NAND2_X2 port map( A1 => n18169, A2 => n33312, ZN => n18168);
   U10497 : NAND4_X2 port map( A1 => n25768, A2 => n25770, A3 => n29168, A4 => 
                           n25769, ZN => n26571);
   U2442 : NOR2_X2 port map( A1 => n14752, A2 => n24915, ZN => n24905);
   U12077 : INV_X4 port map( I => n8790, ZN => n1009);
   U15791 : INV_X1 port map( I => n6969, ZN => n6968);
   U3830 : BUF_X2 port map( I => n20423, Z => n4647);
   U11981 : INV_X2 port map( I => n18960, ZN => n18959);
   U1121 : INV_X2 port map( I => n32606, ZN => n22608);
   U1989 : BUF_X2 port map( I => n2983, Z => n42);
   U5322 : NOR2_X2 port map( A1 => n9797, A2 => n11943, ZN => n11078);
   U1140 : OAI21_X2 port map( A1 => n27991, A2 => n21627, B => n16601, ZN => 
                           n28712);
   U2964 : NAND2_X2 port map( A1 => n1287, A2 => n15644, ZN => n30703);
   U619 : OAI21_X2 port map( A1 => n17064, A2 => n11929, B => n22830, ZN => 
                           n18056);
   U24244 : NAND2_X2 port map( A1 => n18472, A2 => n22, ZN => n18389);
   U2096 : INV_X2 port map( I => n18696, ZN => n12951);
   U5806 : INV_X2 port map( I => n10438, ZN => n16306);
   U24840 : OAI21_X2 port map( A1 => n21419, A2 => n4381, B => n21117, ZN => 
                           n21119);
   U3708 : BUF_X4 port map( I => n10974, Z => n29047);
   U21216 : NAND2_X2 port map( A1 => n14576, A2 => n14815, ZN => n19966);
   U7017 : NAND2_X2 port map( A1 => n680, A2 => n24610, ZN => n3013);
   U14 : INV_X2 port map( I => n24927, ZN => n24933);
   U21764 : INV_X2 port map( I => n18648, ZN => n17114);
   U2366 : BUF_X2 port map( I => n18186, Z => n10964);
   U18311 : NOR2_X2 port map( A1 => n31428, A2 => n17477, ZN => n18886);
   U4217 : OR2_X1 port map( A1 => n6555, A2 => n14770, Z => n9148);
   U972 : INV_X2 port map( I => n9789, ZN => n10288);
   U24634 : NAND2_X2 port map( A1 => n20025, A2 => n16461, ZN => n20026);
   U667 : OAI21_X2 port map( A1 => n22722, A2 => n22908, B => n30447, ZN => 
                           n22556);
   U64 : INV_X2 port map( I => n16751, ZN => n16752);
   U2273 : INV_X2 port map( I => n4124, ZN => n22720);
   U4964 : INV_X2 port map( I => n11900, ZN => n25630);
   U4755 : NOR2_X2 port map( A1 => n28704, A2 => n5433, ZN => n19824);
   U13447 : AOI21_X2 port map( A1 => n7767, A2 => n29819, B => n30121, ZN => 
                           n8114);
   U2012 : INV_X4 port map( I => n1060, ZN => n31428);
   U22052 : INV_X2 port map( I => n19252, ZN => n28276);
   U23951 : INV_X2 port map( I => n17559, ZN => n19990);
   U759 : INV_X2 port map( I => n23086, ZN => n28948);
   U6654 : NAND2_X1 port map( A1 => n7319, A2 => n7318, ZN => n2706);
   U3382 : INV_X4 port map( I => n8100, ZN => n1172);
   U5454 : INV_X4 port map( I => n10845, ZN => n1039);
   U8396 : INV_X2 port map( I => n10351, ZN => n7719);
   U8817 : AOI21_X2 port map( A1 => n18515, A2 => n11918, B => n13663, ZN => 
                           n9211);
   U4063 : OR2_X1 port map( A1 => n22737, A2 => n2449, Z => n23030);
   U159 : NAND2_X2 port map( A1 => n9275, A2 => n24157, ZN => n24206);
   U3618 : NAND3_X2 port map( A1 => n32816, A2 => n21427, A3 => n33949, ZN => 
                           n14618);
   U5177 : AOI21_X2 port map( A1 => n19060, A2 => n9787, B => n1374, ZN => 
                           n2411);
   U8730 : NOR2_X2 port map( A1 => n18363, A2 => n18161, ZN => n18160);
   U1741 : NAND2_X2 port map( A1 => n29208, A2 => n20043, ZN => n11414);
   U10126 : NOR2_X2 port map( A1 => n6470, A2 => n785, ZN => n5122);
   U6257 : BUF_X4 port map( I => n6846, Z => n5119);
   U2188 : OAI21_X1 port map( A1 => n292, A2 => n12358, B => n30019, ZN => 
                           n24467);
   U10177 : NOR2_X2 port map( A1 => n9305, A2 => n5225, ZN => n9215);
   U6340 : INV_X2 port map( I => n8857, ZN => n6748);
   U14716 : NOR2_X1 port map( A1 => n6041, A2 => n6042, ZN => n3996);
   U13804 : INV_X2 port map( I => n27007, ZN => n22899);
   U1725 : OAI21_X2 port map( A1 => n16675, A2 => n31745, B => n29845, ZN => 
                           n4209);
   U3435 : OR2_X2 port map( A1 => n17306, A2 => n14911, Z => n25887);
   U4950 : INV_X2 port map( I => n20630, ZN => n20213);
   U2625 : OAI21_X2 port map( A1 => n801, A2 => n31179, B => n23640, ZN => 
                           n29570);
   U4224 : NAND2_X2 port map( A1 => n23956, A2 => n23824, ZN => n18044);
   U24872 : NAND2_X2 port map( A1 => n28869, A2 => n21430, ZN => n21331);
   U2072 : NAND2_X2 port map( A1 => n18618, A2 => n18779, ZN => n30686);
   U15153 : BUF_X4 port map( I => n22871, Z => n31861);
   U6098 : BUF_X2 port map( I => n18780, Z => n31095);
   U19953 : NOR2_X2 port map( A1 => n22339, A2 => n14145, ZN => n22786);
   U1477 : OAI21_X2 port map( A1 => n26554, A2 => n26553, B => n25960, ZN => 
                           n13705);
   U8759 : OAI22_X2 port map( A1 => n18606, A2 => n18607, B1 => n18605, B2 => 
                           n18604, ZN => n12768);
   U10143 : AOI21_X2 port map( A1 => n18493, A2 => n5677, B => n18324, ZN => 
                           n15071);
   U15790 : AOI21_X2 port map( A1 => n23082, A2 => n22885, B => n13592, ZN => 
                           n12450);
   U10828 : BUF_X2 port map( I => n23696, Z => n8217);
   U2484 : NAND3_X2 port map( A1 => n2715, A2 => n2716, A3 => n16473, ZN => 
                           n2719);
   U15767 : NAND3_X2 port map( A1 => n27103, A2 => n5757, A3 => n33571, ZN => 
                           n21886);
   U23588 : INV_X4 port map( I => n17767, ZN => n28502);
   U5270 : NAND2_X2 port map( A1 => n29462, A2 => n12310, ZN => n7839);
   U3241 : INV_X2 port map( I => n18983, ZN => n17339);
   U2798 : OAI22_X2 port map( A1 => n11299, A2 => n8453, B1 => n7430, B2 => 
                           n21328, ZN => n21334);
   U1681 : NAND2_X2 port map( A1 => n17688, A2 => n19901, ZN => n20109);
   U7614 : NOR2_X2 port map( A1 => n497, A2 => n18535, ZN => n18704);
   U8475 : INV_X2 port map( I => n20633, ZN => n2873);
   U16674 : NAND2_X1 port map( A1 => n8955, A2 => n8958, ZN => n27363);
   U816 : NAND2_X2 port map( A1 => n6027, A2 => n20066, ZN => n20094);
   U4820 : OAI22_X2 port map( A1 => n25943, A2 => n11814, B1 => n12037, B2 => 
                           n21358, ZN => n21359);
   U19642 : INV_X2 port map( I => n20120, ZN => n20019);
   U12950 : INV_X1 port map( I => n7896, ZN => n30075);
   U7588 : NOR2_X2 port map( A1 => n1060, A2 => n18660, ZN => n18887);
   U15481 : OAI21_X2 port map( A1 => n1051, A2 => n18919, B => n15534, ZN => 
                           n4622);
   U17232 : NAND3_X2 port map( A1 => n27814, A2 => n22981, A3 => n29329, ZN => 
                           n30447);
   U1784 : BUF_X4 port map( I => n21006, Z => n28262);
   U175 : INV_X2 port map( I => n9962, ZN => n1246);
   U20199 : INV_X2 port map( I => n5226, ZN => n24221);
   U1227 : NAND2_X2 port map( A1 => n29676, A2 => n20392, ZN => n28900);
   U942 : INV_X4 port map( I => n12585, ZN => n1051);
   U2833 : OAI22_X2 port map( A1 => n13913, A2 => n32951, B1 => n13219, B2 => 
                           n4210, ZN => n13541);
   U8138 : NAND2_X1 port map( A1 => n17734, A2 => n1132, ZN => n11536);
   U14017 : OAI21_X2 port map( A1 => n30181, A2 => n18292, B => n18290, ZN => 
                           n8482);
   U12534 : OAI21_X2 port map( A1 => n30931, A2 => n17790, B => n20562, ZN => 
                           n3352);
   U5649 : INV_X2 port map( I => n17201, ZN => n809);
   U23 : INV_X2 port map( I => n5942, ZN => n6092);
   U6646 : NOR2_X2 port map( A1 => n32005, A2 => n6597, ZN => n6920);
   U69 : INV_X2 port map( I => n25437, ZN => n11640);
   U22948 : OAI22_X2 port map( A1 => n22817, A2 => n33968, B1 => n13597, B2 => 
                           n22818, ZN => n22819);
   U1537 : OAI21_X2 port map( A1 => n16011, A2 => n20359, B => n30793, ZN => 
                           n2319);
   U6623 : INV_X4 port map( I => n19220, ZN => n9787);
   U1868 : NAND2_X2 port map( A1 => n31161, A2 => n9563, ZN => n11872);
   U5709 : INV_X2 port map( I => n548, ZN => n15272);
   U912 : INV_X2 port map( I => n14760, ZN => n1374);
   U1069 : NAND2_X2 port map( A1 => n10456, A2 => n2300, ZN => n2299);
   U79 : INV_X2 port map( I => n25378, ZN => n750);
   U20376 : NOR2_X2 port map( A1 => n8403, A2 => n8402, ZN => n27972);
   U6875 : NAND2_X2 port map( A1 => n6247, A2 => n893, ZN => n11589);
   U11866 : OAI21_X2 port map( A1 => n11971, A2 => n16307, B => n8259, ZN => 
                           n19929);
   U1235 : NAND2_X2 port map( A1 => n1158, A2 => n20614, ZN => n28603);
   U2040 : INV_X2 port map( I => n4734, ZN => n22826);
   U3448 : OAI21_X2 port map( A1 => n2923, A2 => n24057, B => n27592, ZN => 
                           n2922);
   U2298 : INV_X2 port map( I => n19849, ZN => n9563);
   U8584 : INV_X2 port map( I => n11198, ZN => n6970);
   U6116 : NOR2_X2 port map( A1 => n33990, A2 => n2847, ZN => n2851);
   U9011 : INV_X2 port map( I => n10183, ZN => n10202);
   U15564 : INV_X4 port map( I => n23828, ZN => n23669);
   U3188 : BUF_X2 port map( I => n7195, Z => n31498);
   U2858 : OAI22_X2 port map( A1 => n25113, A2 => n16632, B1 => n14895, B2 => 
                           n18132, ZN => n27575);
   U6285 : INV_X2 port map( I => n22737, ZN => n850);
   U4835 : INV_X1 port map( I => n21248, ZN => n22521);
   U5152 : NAND2_X2 port map( A1 => n12585, A2 => n25959, ZN => n18958);
   U14032 : NOR2_X2 port map( A1 => n32018, A2 => n28320, ZN => n30182);
   U2226 : INV_X4 port map( I => n1931, ZN => n16651);
   U4378 : INV_X2 port map( I => n14797, ZN => n26608);
   U660 : NOR2_X2 port map( A1 => n9377, A2 => n23017, ZN => n14797);
   U7461 : NAND2_X2 port map( A1 => n10453, A2 => n19050, ZN => n10452);
   U1050 : INV_X2 port map( I => n21706, ZN => n1316);
   U25795 : NAND2_X2 port map( A1 => n28802, A2 => n3425, ZN => n3424);
   U8132 : INV_X2 port map( I => n51, ZN => n848);
   U15119 : INV_X2 port map( I => n9980, ZN => n16933);
   U4962 : NOR2_X2 port map( A1 => n13074, A2 => n34115, ZN => n9615);
   U10548 : OAI22_X2 port map( A1 => n4961, A2 => n26580, B1 => n4960, B2 => 
                           n15068, ZN => n4959);
   U15438 : AOI21_X2 port map( A1 => n7830, A2 => n33641, B => n14563, ZN => 
                           n7206);
   U13433 : NAND2_X2 port map( A1 => n2514, A2 => n862, ZN => n2513);
   U16640 : AOI21_X2 port map( A1 => n18539, A2 => n18537, B => n14651, ZN => 
                           n5457);
   U9115 : NOR2_X2 port map( A1 => n30724, A2 => n17604, ZN => n30142);
   U50 : INV_X2 port map( I => n25901, ZN => n7143);
   U22526 : NOR2_X2 port map( A1 => n6298, A2 => n6666, ZN => n31223);
   U7000 : INV_X2 port map( I => n17673, ZN => n25403);
   U5213 : INV_X2 port map( I => n25479, ZN => n25486);
   U18060 : NAND2_X2 port map( A1 => n13407, A2 => n4381, ZN => n7118);
   U11455 : NAND2_X2 port map( A1 => n7206, A2 => n7205, ZN => n7204);
   U3329 : INV_X2 port map( I => n10226, ZN => n10513);
   U13637 : INV_X4 port map( I => n9133, ZN => n10113);
   U16375 : AOI21_X2 port map( A1 => n21580, A2 => n5795, B => n3467, ZN => 
                           n7349);
   U880 : INV_X2 port map( I => n17303, ZN => n31506);
   U8800 : NAND2_X2 port map( A1 => n34013, A2 => n4071, ZN => n10105);
   U687 : INV_X2 port map( I => n6681, ZN => n15874);
   U10948 : NAND2_X1 port map( A1 => n24449, A2 => n1079, ZN => n11696);
   U8537 : OAI21_X2 port map( A1 => n8294, A2 => n8295, B => n19863, ZN => 
                           n2674);
   U1297 : NOR2_X2 port map( A1 => n21705, A2 => n21704, ZN => n21794);
   U7188 : INV_X4 port map( I => n21322, ZN => n15015);
   U582 : INV_X2 port map( I => n28343, ZN => n31810);
   U9423 : CLKBUF_X4 port map( I => n580, Z => n29676);
   U3544 : INV_X2 port map( I => n31954, ZN => n1007);
   U324 : AOI21_X2 port map( A1 => n24263, A2 => n15974, B => n1239, ZN => 
                           n31785);
   U7498 : NOR2_X2 port map( A1 => n10229, A2 => n33335, ZN => n10857);
   U6299 : BUF_X4 port map( I => n20133, Z => n16637);
   U4350 : AND2_X1 port map( A1 => n29928, A2 => n11986, Z => n7851);
   U24657 : NAND3_X2 port map( A1 => n9688, A2 => n13920, A3 => n1154, ZN => 
                           n20180);
   U7025 : INV_X2 port map( I => n25621, ZN => n25752);
   U11478 : AOI22_X2 port map( A1 => n1374, A2 => n29146, B1 => n31757, B2 => 
                           n16185, ZN => n31213);
   U20791 : NAND2_X2 port map( A1 => n22811, A2 => n22810, ZN => n16028);
   U6602 : OAI21_X2 port map( A1 => n11228, A2 => n7183, B => n15595, ZN => 
                           n31148);
   U15127 : INV_X2 port map( I => n19310, ZN => n14178);
   U10065 : NAND2_X2 port map( A1 => n10229, A2 => n25985, ZN => n10352);
   U8016 : BUF_X2 port map( I => n15502, Z => n31726);
   U2408 : NAND2_X2 port map( A1 => n33146, A2 => n21721, ZN => n21580);
   U6571 : INV_X2 port map( I => n17369, ZN => n16081);
   U1998 : OAI22_X2 port map( A1 => n18615, A2 => n31115, B1 => n18029, B2 => 
                           n16948, ZN => n31459);
   U13224 : OAI22_X2 port map( A1 => n1469, A2 => n20379, B1 => n2904, B2 => 
                           n2203, ZN => n26907);
   U1712 : NAND2_X2 port map( A1 => n2879, A2 => n868, ZN => n31393);
   U318 : NAND2_X2 port map( A1 => n10427, A2 => n9946, ZN => n28488);
   U3411 : NOR2_X2 port map( A1 => n27697, A2 => n20595, ZN => n20258);
   U10831 : INV_X4 port map( I => n906, ZN => n30641);
   U26249 : AOI22_X2 port map( A1 => n4867, A2 => n24926, B1 => n24921, B2 => 
                           n15569, ZN => n29127);
   U4380 : INV_X2 port map( I => n8622, ZN => n13934);
   U11863 : OR2_X1 port map( A1 => n8244, A2 => n2927, Z => n2934);
   U6249 : NAND2_X2 port map( A1 => n19267, A2 => n18974, ZN => n13831);
   U1977 : NOR2_X2 port map( A1 => n26417, A2 => n8141, ZN => n19032);
   U21417 : NAND2_X2 port map( A1 => n28130, A2 => n8137, ZN => n29211);
   U2050 : INV_X2 port map( I => n27779, ZN => n25169);
   U2465 : OAI21_X2 port map( A1 => n3842, A2 => n1567, B => n2909, ZN => 
                           n27779);
   U6787 : NAND2_X2 port map( A1 => n11268, A2 => n10031, ZN => n27556);
   U14331 : AOI22_X2 port map( A1 => n3407, A2 => n16694, B1 => n12061, B2 => 
                           n1360, ZN => n15965);
   U7360 : NAND2_X2 port map( A1 => n17456, A2 => n11350, ZN => n11408);
   U5993 : AOI21_X2 port map( A1 => n20125, A2 => n20124, B => n20123, ZN => 
                           n20126);
   U6321 : NAND2_X2 port map( A1 => n1926, A2 => n17891, ZN => n17890);
   U21763 : INV_X2 port map( I => n18392, ZN => n15888);
   U24 : BUF_X2 port map( I => n17927, Z => n29085);
   U1762 : OAI21_X1 port map( A1 => n14426, A2 => n33069, B => n8193, ZN => 
                           n14425);
   U7396 : NAND2_X2 port map( A1 => n19993, A2 => n1040, ZN => n2288);
   U4161 : BUF_X2 port map( I => n17261, Z => n28436);
   U482 : NOR2_X2 port map( A1 => n4991, A2 => n23828, ZN => n13196);
   U20913 : AOI21_X2 port map( A1 => n14864, A2 => n21877, B => n28059, ZN => 
                           n15315);
   U694 : INV_X4 port map( I => n21070, ZN => n21430);
   U7543 : NOR2_X2 port map( A1 => n5456, A2 => n1185, ZN => n6793);
   U6567 : NOR2_X2 port map( A1 => n21583, A2 => n21781, ZN => n8164);
   U2089 : AOI22_X2 port map( A1 => n21711, A2 => n727, B1 => n862, B2 => 
                           n21710, ZN => n6514);
   U10422 : NAND2_X2 port map( A1 => n24224, A2 => n10687, ZN => n28467);
   U1511 : INV_X2 port map( I => n3351, ZN => n20789);
   U5430 : BUF_X4 port map( I => n2566, Z => n2565);
   U8407 : NAND2_X2 port map( A1 => n20486, A2 => n20485, ZN => n20252);
   U6476 : OAI21_X2 port map( A1 => n11445, A2 => n10848, B => n10074, ZN => 
                           n30552);
   U14925 : INV_X2 port map( I => n11676, ZN => n30359);
   U2368 : NOR2_X2 port map( A1 => n15371, A2 => n7868, ZN => n17354);
   U1495 : CLKBUF_X4 port map( I => n16239, Z => n5822);
   U3041 : NAND2_X2 port map( A1 => n8219, A2 => n561, ZN => n9612);
   U6530 : NAND3_X2 port map( A1 => n27715, A2 => n17711, A3 => n11264, ZN => 
                           n10152);
   U1739 : OAI21_X2 port map( A1 => n27541, A2 => n27542, B => n15110, ZN => 
                           n31173);
   U2002 : NOR2_X2 port map( A1 => n15789, A2 => n13554, ZN => n30648);
   U2505 : NOR2_X2 port map( A1 => n27, A2 => n23691, ZN => n28688);
   U5114 : INV_X2 port map( I => n6556, ZN => n17640);
   U1369 : NAND2_X2 port map( A1 => n27715, A2 => n19947, ZN => n27714);
   U7427 : INV_X2 port map( I => n5433, ZN => n10444);
   U3262 : NAND2_X2 port map( A1 => n26158, A2 => n26157, ZN => n24063);
   U4172 : INV_X4 port map( I => n14849, ZN => n1137);
   U9497 : AOI21_X2 port map( A1 => n32079, A2 => n14848, B => n33842, ZN => 
                           n6698);
   U15611 : INV_X1 port map( I => n32647, ZN => n21413);
   U5007 : BUF_X4 port map( I => n19122, Z => n15534);
   U45 : INV_X4 port map( I => n25276, ZN => n25278);
   U2576 : AOI22_X2 port map( A1 => n22837, A2 => n10360, B1 => n22835, B2 => 
                           n22836, ZN => n4231);
   U18297 : INV_X2 port map( I => n19484, ZN => n27607);
   U17842 : INV_X4 port map( I => n3748, ZN => n16443);
   U2468 : NOR2_X2 port map( A1 => n3085, A2 => n384, ZN => n11105);
   U1723 : INV_X2 port map( I => n20335, ZN => n20546);
   U6943 : BUF_X2 port map( I => n5317, Z => n29866);
   U15945 : AOI22_X2 port map( A1 => n6770, A2 => n24191, B1 => n28726, B2 => 
                           n6769, ZN => n6768);
   U4557 : AOI21_X2 port map( A1 => n1155, A2 => n33721, B => n32941, ZN => 
                           n29692);
   U4261 : BUF_X4 port map( I => n13719, Z => n13663);
   U9493 : OAI21_X2 port map( A1 => n16953, A2 => n16952, B => n18079, ZN => 
                           n7703);
   U10706 : NAND2_X2 port map( A1 => n15272, A2 => n23638, ZN => n8799);
   U1525 : INV_X2 port map( I => n20670, ZN => n21046);
   U6500 : INV_X4 port map( I => n20607, ZN => n15217);
   U17368 : NAND3_X2 port map( A1 => n17808, A2 => n29603, A3 => n17809, ZN => 
                           n15745);
   U1980 : AOI21_X2 port map( A1 => n16485, A2 => n13685, B => n947, ZN => 
                           n9078);
   U1421 : INV_X2 port map( I => n17711, ZN => n942);
   U2933 : OAI21_X2 port map( A1 => n33097, A2 => n1098, B => n4538, ZN => 
                           n17923);
   U7094 : AND2_X1 port map( A1 => n13936, A2 => n31650, Z => n29353);
   U5028 : BUF_X2 port map( I => n23683, Z => n23864);
   U6974 : BUF_X4 port map( I => n24180, Z => n5913);
   U15167 : NOR2_X1 port map( A1 => n2069, A2 => n9788, ZN => n28700);
   U12883 : BUF_X4 port map( I => n14339, Z => n30065);
   U15671 : NAND2_X2 port map( A1 => n6962, A2 => n4373, ZN => n13583);
   U973 : BUF_X4 port map( I => n22411, Z => n31551);
   U502 : INV_X2 port map( I => n23770, ZN => n27910);
   U599 : INV_X2 port map( I => n23508, ZN => n1259);
   U871 : INV_X2 port map( I => n9370, ZN => n29232);
   U19191 : NOR2_X2 port map( A1 => n14027, A2 => n8582, ZN => n13572);
   U425 : NAND2_X2 port map( A1 => n12817, A2 => n23752, ZN => n12816);
   U74 : BUF_X2 port map( I => n25490, Z => n4183);
   U3547 : OAI21_X2 port map( A1 => n20594, A2 => n29603, B => n20599, ZN => 
                           n31401);
   U6443 : NAND2_X2 port map( A1 => n27697, A2 => n27070, ZN => n20599);
   U1276 : NAND2_X2 port map( A1 => n28379, A2 => n744, ZN => n19136);
   U1103 : INV_X2 port map( I => n30506, ZN => n1326);
   U14412 : NOR2_X2 port map( A1 => n19122, A2 => n30879, ZN => n26550);
   U224 : OAI21_X2 port map( A1 => n1634, A2 => n8004, B => n4458, ZN => n8003)
                           ;
   U15426 : AOI22_X2 port map( A1 => n1820, A2 => n992, B1 => n17394, B2 => 
                           n22583, ZN => n1486);
   U17000 : NAND3_X2 port map( A1 => n161, A2 => n1036, A3 => n27345, ZN => 
                           n3272);
   U5271 : INV_X2 port map( I => n12310, ZN => n5135);
   U15075 : NAND2_X2 port map( A1 => n24057, A2 => n31918, ZN => n24496);
   U24626 : AOI21_X2 port map( A1 => n26567, A2 => n28471, B => n741, ZN => 
                           n20001);
   U2425 : NOR2_X2 port map( A1 => n14384, A2 => n32384, ZN => n11644);
   U3175 : NAND2_X2 port map( A1 => n12715, A2 => n23318, ZN => n3281);
   U20445 : INV_X4 port map( I => n29335, ZN => n15322);
   U5109 : AND2_X1 port map( A1 => n23692, A2 => n13147, Z => n31239);
   U5453 : INV_X2 port map( I => n17405, ZN => n19819);
   U11065 : NAND2_X1 port map( A1 => n9030, A2 => n9032, ZN => n30119);
   U4623 : OAI21_X2 port map( A1 => n14461, A2 => n1316, B => n21613, ZN => 
                           n6253);
   U372 : BUF_X2 port map( I => n8178, Z => n29977);
   U9471 : INV_X2 port map( I => n29854, ZN => n26474);
   U19205 : INV_X1 port map( I => n30731, ZN => n6257);
   U15476 : NAND2_X2 port map( A1 => n786, A2 => n10858, ZN => n10574);
   U3150 : NAND2_X2 port map( A1 => n20155, A2 => n10059, ZN => n2089);
   U776 : NOR2_X2 port map( A1 => n28101, A2 => n29957, ZN => n28035);
   U8748 : NOR2_X2 port map( A1 => n15018, A2 => n1185, ZN => n18161);
   U2602 : NAND2_X2 port map( A1 => n15682, A2 => n23860, ZN => n11158);
   U19615 : INV_X4 port map( I => n9390, ZN => n15394);
   U3695 : NOR2_X2 port map( A1 => n18617, A2 => n18616, ZN => n16418);
   U4377 : INV_X2 port map( I => n25007, ZN => n1205);
   U12141 : NAND2_X2 port map( A1 => n11270, A2 => n33039, ZN => n10247);
   U26161 : INV_X2 port map( I => n24785, ZN => n1085);
   U1479 : NAND2_X2 port map( A1 => n31004, A2 => n9439, ZN => n31003);
   U8086 : INV_X1 port map( I => n16306, ZN => n22621);
   U13175 : INV_X4 port map( I => n2256, ZN => n22780);
   U147 : NAND2_X2 port map( A1 => n18154, A2 => n25114, ZN => n16024);
   U480 : INV_X1 port map( I => n2021, ZN => n14497);
   U2648 : INV_X4 port map( I => n33069, ZN => n19181);
   U3895 : INV_X2 port map( I => n27931, ZN => n5335);
   U8724 : NAND3_X2 port map( A1 => n22624, A2 => n22623, A3 => n2538, ZN => 
                           n26393);
   U5388 : INV_X2 port map( I => n22098, ZN => n22260);
   U19442 : INV_X2 port map( I => n22072, ZN => n27837);
   U8085 : INV_X2 port map( I => n2547, ZN => n994);
   U439 : INV_X4 port map( I => n22534, ZN => n1120);
   U3579 : BUF_X4 port map( I => n5625, Z => n4643);
   U5524 : INV_X2 port map( I => n7195, ZN => n927);
   U3894 : BUF_X4 port map( I => n17967, Z => n27345);
   U1493 : INV_X2 port map( I => n12804, ZN => n21223);
   U17223 : INV_X2 port map( I => n16011, ZN => n27426);
   U10129 : OAI21_X2 port map( A1 => n9215, A2 => n18518, B => n18672, ZN => 
                           n9304);
   U1419 : INV_X2 port map( I => n21109, ZN => n17438);
   U5979 : INV_X4 port map( I => n14454, ZN => n3080);
   U1542 : BUF_X2 port map( I => n19289, Z => n28528);
   U6599 : NOR2_X2 port map( A1 => n19357, A2 => n19229, ZN => n19354);
   U5139 : NOR2_X2 port map( A1 => n5962, A2 => n28825, ZN => n29928);
   U8258 : AOI21_X2 port map( A1 => n15220, A2 => n15219, B => n32799, ZN => 
                           n15358);
   U15782 : AOI21_X2 port map( A1 => n4371, A2 => n10947, B => n13747, ZN => 
                           n4370);
   U4607 : INV_X2 port map( I => n19947, ZN => n11264);
   U2938 : BUF_X2 port map( I => n26363, Z => n31072);
   U13167 : NAND2_X2 port map( A1 => n28528, A2 => n10124, ZN => n19076);
   U3010 : OAI21_X1 port map( A1 => n23688, A2 => n17181, B => n25987, ZN => 
                           n23689);
   U1034 : BUF_X2 port map( I => n4034, Z => n27850);
   U834 : NAND2_X2 port map( A1 => n11161, A2 => n22669, ZN => n2311);
   U4196 : OR2_X1 port map( A1 => n24466, A2 => n292, Z => n26281);
   U15271 : NOR2_X2 port map( A1 => n776, A2 => n14686, ZN => n28071);
   U15622 : NAND2_X2 port map( A1 => n2577, A2 => n347, ZN => n30291);
   U4752 : BUF_X4 port map( I => n596, Z => n28287);
   U21006 : INV_X2 port map( I => n19637, ZN => n15063);
   U2639 : INV_X4 port map( I => n17895, ZN => n844);
   U6995 : NOR2_X2 port map( A1 => n24973, A2 => n17118, ZN => n17782);
   U2513 : AOI21_X2 port map( A1 => n10589, A2 => n22919, B => n10588, ZN => 
                           n10760);
   U7426 : INV_X4 port map( I => n12168, ZN => n8927);
   U656 : NOR2_X2 port map( A1 => n28314, A2 => n3614, ZN => n12728);
   U7069 : BUF_X2 port map( I => Key(177), Z => n25436);
   U6929 : INV_X2 port map( I => n23109, ZN => n1264);
   U3623 : OR2_X1 port map( A1 => n19915, A2 => n31671, Z => n28208);
   U22197 : NOR2_X2 port map( A1 => n818, A2 => n20411, ZN => n28268);
   U17087 : OAI21_X2 port map( A1 => n18953, A2 => n18952, B => n28935, ZN => 
                           n11336);
   U4516 : NAND2_X2 port map( A1 => n20468, A2 => n14138, ZN => n6536);
   U8029 : NAND2_X2 port map( A1 => n27737, A2 => n30066, ZN => n15919);
   U6780 : NAND2_X2 port map( A1 => n12952, A2 => n16432, ZN => n27737);
   U10699 : NAND2_X1 port map( A1 => n14497, A2 => n14496, ZN => n2036);
   U18957 : NAND2_X2 port map( A1 => n19927, A2 => n30554, ZN => n19928);
   U9877 : OAI21_X2 port map( A1 => n6970, A2 => n19926, B => n13591, ZN => 
                           n19927);
   U4317 : BUF_X2 port map( I => Key(47), Z => n25195);
   U6807 : INV_X2 port map( I => n24243, ZN => n24337);
   U10231 : CLKBUF_X2 port map( I => Key(159), Z => n25881);
   U7842 : NAND2_X1 port map( A1 => n12020, A2 => n313, ZN => n12858);
   U2907 : NAND2_X2 port map( A1 => n20335, A2 => n30130, ZN => n20411);
   U2062 : NAND2_X2 port map( A1 => n489, A2 => n4194, ZN => n17321);
   U13793 : NOR2_X2 port map( A1 => n15434, A2 => n2843, ZN => n17993);
   U10085 : INV_X4 port map( I => n29146, ZN => n1179);
   U4762 : NAND2_X2 port map( A1 => n24167, A2 => n24279, ZN => n11121);
   U7848 : NOR2_X2 port map( A1 => n23778, A2 => n23775, ZN => n5438);
   U6295 : INV_X2 port map( I => n19406, ZN => n31755);
   U18497 : INV_X2 port map( I => n14138, ZN => n742);
   U5298 : NAND2_X2 port map( A1 => n20059, A2 => n224, ZN => n12696);
   U21970 : INV_X4 port map( I => n12707, ZN => n13210);
   U1238 : NOR2_X1 port map( A1 => n12354, A2 => n12394, ZN => n30619);
   U1157 : INV_X2 port map( I => n21743, ZN => n31654);
   U689 : INV_X2 port map( I => n16129, ZN => n16906);
   U2145 : BUF_X2 port map( I => n12707, Z => n12249);
   U3034 : AND2_X2 port map( A1 => n26114, A2 => n10772, Z => n23809);
   U2975 : OR2_X2 port map( A1 => n5975, A2 => n625, Z => n22364);
   U14485 : INV_X2 port map( I => n10390, ZN => n4568);
   U13486 : AOI22_X2 port map( A1 => n34005, A2 => n30932, B1 => n13475, B2 => 
                           n29715, ZN => n15486);
   U1558 : NAND2_X2 port map( A1 => n8689, A2 => n17234, ZN => n32);
   U1163 : INV_X1 port map( I => n6842, ZN => n21075);
   U14037 : OAI21_X2 port map( A1 => n13428, A2 => n24780, B => n3080, ZN => 
                           n3079);
   U9144 : OAI21_X1 port map( A1 => n29743, A2 => n12654, B => n29742, ZN => 
                           n7207);
   U25183 : NAND3_X2 port map( A1 => n27589, A2 => n13778, A3 => n6149, ZN => 
                           n23021);
   U845 : OAI21_X2 port map( A1 => n28902, A2 => n22280, B => n22379, ZN => 
                           n261);
   U6376 : NAND2_X2 port map( A1 => n20089, A2 => n2229, ZN => n11120);
   U12927 : OR2_X1 port map( A1 => n23805, A2 => n2752, Z => n2004);
   U2181 : OAI21_X2 port map( A1 => n2945, A2 => n13268, B => n2943, ZN => 
                           n15303);
   U3750 : INV_X4 port map( I => n14392, ZN => n4113);
   U5417 : NAND3_X2 port map( A1 => n33301, A2 => n13300, A3 => n20310, ZN => 
                           n13563);
   U6914 : INV_X4 port map( I => n29785, ZN => n24213);
   U4420 : OR2_X1 port map( A1 => n32903, A2 => n16144, Z => n2675);
   U5718 : INV_X2 port map( I => n10193, ZN => n1098);
   U15562 : NAND3_X1 port map( A1 => n23616, A2 => n33260, A3 => n23828, ZN => 
                           n9998);
   U13954 : INV_X4 port map( I => n3601, ZN => n18893);
   U9950 : INV_X2 port map( I => n17456, ZN => n16579);
   U2131 : NOR2_X2 port map( A1 => n15246, A2 => n15247, ZN => n13302);
   U2083 : INV_X4 port map( I => n2019, ZN => n29658);
   U7336 : BUF_X2 port map( I => n12375, Z => n6553);
   U2683 : NOR2_X2 port map( A1 => n10264, A2 => n959, ZN => n8309);
   U674 : INV_X2 port map( I => n8490, ZN => n11215);
   U4586 : NAND2_X2 port map( A1 => n12836, A2 => n34054, ZN => n6014);
   U2718 : BUF_X4 port map( I => n10657, Z => n7007);
   U1893 : NAND3_X2 port map( A1 => n26288, A2 => n29118, A3 => n19256, ZN => 
                           n18526);
   U755 : INV_X2 port map( I => n33007, ZN => n13474);
   U14915 : NAND3_X2 port map( A1 => n14106, A2 => n14107, A3 => n9221, ZN => 
                           n20503);
   U18411 : NAND2_X2 port map( A1 => n19457, A2 => n33631, ZN => n7708);
   U3931 : NAND2_X2 port map( A1 => n33007, A2 => n33115, ZN => n30364);
   U15166 : AOI21_X2 port map( A1 => n24191, A2 => n795, B => n28726, ZN => 
                           n24172);
   U2326 : NOR2_X2 port map( A1 => n27678, A2 => n1257, ZN => n23308);
   U6771 : NOR2_X2 port map( A1 => n22664, A2 => n22576, ZN => n22454);
   U10367 : INV_X2 port map( I => n25513, ZN => n1204);
   U1532 : INV_X4 port map( I => n13160, ZN => n19137);
   U974 : INV_X4 port map( I => n22640, ZN => n29626);
   U4107 : INV_X1 port map( I => n10673, ZN => n23782);
   U2350 : INV_X4 port map( I => n12039, ZN => n1213);
   U15575 : AOI21_X2 port map( A1 => n16443, A2 => n24148, B => n9946, ZN => 
                           n8962);
   U10964 : NAND2_X2 port map( A1 => n22843, A2 => n28330, ZN => n5680);
   U1833 : INV_X2 port map( I => n31408, ZN => n19969);
   U25333 : NOR2_X2 port map( A1 => n1257, A2 => n10142, ZN => n23698);
   U2610 : BUF_X2 port map( I => n25115, Z => n14495);
   U710 : INV_X2 port map( I => n16315, ZN => n15852);
   U448 : NAND2_X2 port map( A1 => n18098, A2 => n27122, ZN => n9620);
   U2775 : BUF_X4 port map( I => n24680, Z => n25561);
   U470 : INV_X2 port map( I => n34125, ZN => n1287);
   U16260 : AND2_X1 port map( A1 => n5035, A2 => n987, Z => n22509);
   U854 : INV_X2 port map( I => n502, ZN => n13061);
   U20478 : NAND2_X2 port map( A1 => n7792, A2 => n33403, ZN => n30924);
   U13010 : OR2_X2 port map( A1 => n18146, A2 => n24031, Z => n24143);
   U15492 : OAI21_X2 port map( A1 => n16443, A2 => n5335, B => n29655, ZN => 
                           n9521);
   U15043 : BUF_X4 port map( I => n25409, Z => n419);
   U289 : NAND2_X2 port map( A1 => n9824, A2 => n9823, ZN => n9825);
   U566 : NOR2_X2 port map( A1 => n8525, A2 => n23819, ZN => n10749);
   U20909 : NOR2_X2 port map( A1 => n21410, A2 => n16473, ZN => n2941);
   U2255 : OAI21_X2 port map( A1 => n24067, A2 => n32036, B => n7503, ZN => 
                           n10827);
   U248 : BUF_X4 port map( I => n6911, Z => n27501);
   U7250 : AOI21_X2 port map( A1 => n20566, A2 => n16515, B => n12263, ZN => 
                           n8941);
   U7371 : INV_X2 port map( I => n19601, ZN => n13591);
   U20282 : INV_X2 port map( I => n27958, ZN => n489);
   U4181 : INV_X2 port map( I => n16077, ZN => n709);
   U3851 : OAI21_X2 port map( A1 => n9261, A2 => n9262, B => n29269, ZN => 
                           n27756);
   U25014 : NAND2_X2 port map( A1 => n621, A2 => n22557, ZN => n22071);
   U4289 : BUF_X2 port map( I => Key(43), Z => n25190);
   U16549 : INV_X2 port map( I => n19969, ZN => n30612);
   U10864 : INV_X2 port map( I => n13814, ZN => n17188);
   U12011 : INV_X4 port map( I => n11940, ZN => n29963);
   U1909 : AOI21_X2 port map( A1 => n880, A2 => n879, B => n15396, ZN => n15395
                           );
   U15465 : AND2_X2 port map( A1 => n29124, A2 => n14587, Z => n27159);
   U2641 : AOI21_X2 port map( A1 => n22438, A2 => n12236, B => n17007, ZN => 
                           n17006);
   U2616 : NAND3_X2 port map( A1 => n26459, A2 => n33544, A3 => n30459, ZN => 
                           n14371);
   U21563 : INV_X2 port map( I => n19844, ZN => n19923);
   U8316 : OR2_X2 port map( A1 => n34151, A2 => n30387, Z => n19888);
   U5868 : INV_X2 port map( I => n20519, ZN => n20517);
   U9048 : NOR2_X2 port map( A1 => n15665, A2 => n20056, ZN => n17573);
   U5448 : NAND2_X2 port map( A1 => n12398, A2 => n71, ZN => n6405);
   U14931 : INV_X2 port map( I => n13040, ZN => n28726);
   U7640 : INV_X2 port map( I => n14159, ZN => n18853);
   U2541 : NAND3_X1 port map( A1 => n5217, A2 => n26587, A3 => n14280, ZN => 
                           n5216);
   U3592 : NOR2_X2 port map( A1 => n7218, A2 => n8770, ZN => n20304);
   U4723 : NAND2_X2 port map( A1 => n20150, A2 => n20152, ZN => n19915);
   U5111 : INV_X1 port map( I => n17590, ZN => n21373);
   U5914 : INV_X2 port map( I => n29688, ZN => n820);
   U6151 : NAND2_X2 port map( A1 => n18496, A2 => n10043, ZN => n8824);
   U12195 : INV_X1 port map( I => n24527, ZN => n16253);
   U1519 : INV_X4 port map( I => n31970, ZN => n763);
   U2980 : NOR2_X2 port map( A1 => n25980, A2 => n397, ZN => n8775);
   U12914 : NAND2_X1 port map( A1 => n26858, A2 => n26856, ZN => n21956);
   U6319 : BUF_X2 port map( I => n12452, Z => n28923);
   U2688 : NAND2_X2 port map( A1 => n18159, A2 => n29070, ZN => n17873);
   U18708 : NAND2_X2 port map( A1 => n10142, A2 => n33216, ZN => n27679);
   U14996 : INV_X2 port map( I => n17717, ZN => n11556);
   U5754 : INV_X2 port map( I => n23695, ZN => n27163);
   U16071 : NAND2_X2 port map( A1 => n26900, A2 => n27457, ZN => n2221);
   U3089 : INV_X2 port map( I => n13670, ZN => n28017);
   U3844 : OAI21_X2 port map( A1 => n5745, A2 => n14119, B => n8273, ZN => 
                           n27377);
   U7927 : NOR2_X2 port map( A1 => n17739, A2 => n32500, ZN => n2222);
   U274 : INV_X2 port map( I => n29323, ZN => n8273);
   U7525 : INV_X2 port map( I => n18988, ZN => n19087);
   U5617 : NAND2_X2 port map( A1 => n5135, A2 => n5380, ZN => n30008);
   U2086 : INV_X1 port map( I => n18677, ZN => n30558);
   U2095 : NAND2_X2 port map( A1 => n15371, A2 => n31511, ZN => n28973);
   U12155 : NAND2_X2 port map( A1 => n18495, A2 => n28987, ZN => n6026);
   U5994 : INV_X2 port map( I => n18847, ZN => n18731);
   U18265 : OAI21_X2 port map( A1 => n16461, A2 => n1042, B => n6109, ZN => 
                           n6108);
   U4802 : NAND2_X2 port map( A1 => n2713, A2 => n7004, ZN => n22838);
   U535 : NOR2_X1 port map( A1 => n8082, A2 => n26780, ZN => n8081);
   U20256 : NOR2_X2 port map( A1 => n16189, A2 => n10686, ZN => n15154);
   U2818 : INV_X4 port map( I => n563, ZN => n11961);
   U5961 : BUF_X2 port map( I => n20445, Z => n31768);
   U2287 : INV_X4 port map( I => n4373, ZN => n5966);
   U1669 : NAND2_X2 port map( A1 => n13341, A2 => n6098, ZN => n13340);
   U4976 : NOR2_X2 port map( A1 => n53, A2 => n7280, ZN => n16882);
   U17887 : NAND3_X2 port map( A1 => n26333, A2 => n9579, A3 => n16432, ZN => 
                           n31689);
   U7993 : AOI22_X1 port map( A1 => n17184, A2 => n18593, B1 => n18594, B2 => 
                           n18849, ZN => n18598);
   U25251 : NAND2_X2 port map( A1 => n9275, A2 => n32349, ZN => n31543);
   U2192 : CLKBUF_X12 port map( I => n2956, Z => n29011);
   U3792 : NOR2_X2 port map( A1 => n23017, A2 => n23018, ZN => n12416);
   U16079 : INV_X2 port map( I => n10420, ZN => n25890);
   U6200 : INV_X4 port map( I => n23807, ZN => n14664);
   U5148 : AOI22_X2 port map( A1 => n10732, A2 => n16906, B1 => n21212, B2 => 
                           n21211, ZN => n29503);
   U7134 : INV_X2 port map( I => n21721, ZN => n1133);
   U539 : NAND3_X2 port map( A1 => n187, A2 => n17773, A3 => n185, ZN => n15677
                           );
   U11795 : INV_X2 port map( I => n11408, ZN => n3407);
   U1524 : NAND2_X2 port map( A1 => n18913, A2 => n7995, ZN => n19100);
   U5991 : BUF_X4 port map( I => n16855, Z => n6597);
   U22960 : AOI21_X2 port map( A1 => n16132, A2 => n1150, B => n14710, ZN => 
                           n20416);
   U7550 : OAI21_X2 port map( A1 => n9090, A2 => n18633, B => n18711, ZN => 
                           n2987);
   U5432 : OAI21_X2 port map( A1 => n215, A2 => n33763, B => n214, ZN => n23623
                           );
   U18436 : NAND2_X1 port map( A1 => n12391, A2 => n12392, ZN => n30623);
   U4855 : CLKBUF_X4 port map( I => n20467, Z => n26567);
   U14940 : INV_X2 port map( I => n11705, ZN => n25348);
   U10967 : NAND2_X2 port map( A1 => n22843, A2 => n33016, ZN => n11467);
   U15097 : OAI21_X2 port map( A1 => n1243, A2 => n23991, B => n23990, ZN => 
                           n23992);
   U3338 : AOI22_X2 port map( A1 => n10853, A2 => n33822, B1 => n10857, B2 => 
                           n25985, ZN => n31406);
   U927 : INV_X4 port map( I => n13295, ZN => n19229);
   U15784 : NAND2_X2 port map( A1 => n26544, A2 => n12143, ZN => n31421);
   U24134 : OAI21_X2 port map( A1 => n18226, A2 => n18848, B => n18849, ZN => 
                           n18224);
   U3176 : AOI21_X1 port map( A1 => n12781, A2 => n12099, B => n23318, ZN => 
                           n12716);
   U3419 : NOR2_X1 port map( A1 => n401, A2 => n8573, ZN => n9123);
   U1547 : INV_X2 port map( I => n11103, ZN => n30882);
   U16111 : INV_X2 port map( I => n10291, ZN => n8270);
   U11093 : NOR2_X2 port map( A1 => n30375, A2 => n19724, ZN => n2927);
   U6525 : INV_X4 port map( I => n21237, ZN => n21453);
   U11283 : NAND2_X1 port map( A1 => n27317, A2 => n27316, ZN => n30454);
   U2807 : NAND2_X2 port map( A1 => n15833, A2 => n29938, ZN => n15832);
   U141 : NOR2_X2 port map( A1 => n10178, A2 => n10177, ZN => n10176);
   U26133 : OAI22_X2 port map( A1 => n29035, A2 => n29034, B1 => n6580, B2 => 
                           n729, ZN => n11493);
   U6393 : NAND2_X2 port map( A1 => n6611, A2 => n11624, ZN => n13021);
   U15117 : NAND2_X2 port map( A1 => n13037, A2 => n13035, ZN => n19319);
   U4376 : OAI21_X2 port map( A1 => n15189, A2 => n20155, B => n11959, ZN => 
                           n27111);
   U2812 : INV_X2 port map( I => n13510, ZN => n16346);
   U1665 : NAND3_X2 port map( A1 => n29365, A2 => n17672, A3 => n14731, ZN => 
                           n30938);
   U7114 : NAND2_X2 port map( A1 => n21632, A2 => n21871, ZN => n4689);
   U11935 : INV_X4 port map( I => n6344, ZN => n3989);
   U13567 : OR2_X2 port map( A1 => n25695, A2 => n25628, Z => n13641);
   U21245 : NOR2_X1 port map( A1 => n28098, A2 => n18194, ZN => n18192);
   U598 : INV_X2 port map( I => n21849, ZN => n21763);
   U6353 : BUF_X4 port map( I => n31922, Z => n16461);
   U17036 : INV_X1 port map( I => n2655, ZN => n27378);
   U2135 : NAND2_X1 port map( A1 => n12441, A2 => n7063, ZN => n30562);
   U21030 : NAND2_X2 port map( A1 => n32940, A2 => n295, ZN => n15344);
   U12508 : OR2_X2 port map( A1 => n13941, A2 => n1696, Z => n19450);
   U17412 : OR2_X2 port map( A1 => n30282, A2 => n6394, Z => n4675);
   U1752 : AOI21_X2 port map( A1 => n15383, A2 => n20066, B => n30771, ZN => 
                           n17346);
   U2600 : NOR2_X2 port map( A1 => n15682, A2 => n23860, ZN => n15681);
   U17076 : NOR2_X2 port map( A1 => n27387, A2 => n13045, ZN => n13043);
   U17077 : NOR2_X2 port map( A1 => n15364, A2 => n3891, ZN => n27387);
   U11396 : INV_X4 port map( I => n21630, ZN => n2217);
   U1956 : NOR2_X2 port map( A1 => n9345, A2 => n9344, ZN => n9343);
   U6237 : NAND2_X2 port map( A1 => n18767, A2 => n4624, ZN => n17905);
   U4616 : NOR2_X1 port map( A1 => n28494, A2 => n11938, ZN => n12787);
   U19587 : NOR2_X1 port map( A1 => n14264, A2 => n14261, ZN => n30798);
   U2617 : NOR2_X2 port map( A1 => n6599, A2 => n914, ZN => n11797);
   U1538 : INV_X2 port map( I => n17586, ZN => n17004);
   U3754 : INV_X2 port map( I => n18575, ZN => n10043);
   U25902 : NOR2_X2 port map( A1 => n19063, A2 => n19108, ZN => n19110);
   U3779 : OR2_X1 port map( A1 => n20219, A2 => n9014, Z => n583);
   U12728 : INV_X4 port map( I => n1835, ZN => n18633);
   U4883 : BUF_X2 port map( I => n9220, Z => n7779);
   U9693 : NAND3_X2 port map( A1 => n26499, A2 => n22828, A3 => n28327, ZN => 
                           n26501);
   U17097 : NAND2_X2 port map( A1 => n6082, A2 => n12654, ZN => n14560);
   U1324 : INV_X2 port map( I => n18187, ZN => n18185);
   U13276 : INV_X2 port map( I => n23057, ZN => n31566);
   U24688 : NAND2_X2 port map( A1 => n384, A2 => n20338, ZN => n20340);
   U6363 : INV_X2 port map( I => n22119, ZN => n22092);
   U3859 : OAI21_X2 port map( A1 => n6285, A2 => n8290, B => n14420, ZN => 
                           n27695);
   U10029 : NAND2_X2 port map( A1 => n18988, A2 => n6510, ZN => n18899);
   U7254 : INV_X4 port map( I => n30879, ZN => n18919);
   U16238 : NOR2_X2 port map( A1 => n33022, A2 => n23034, ZN => n16919);
   U1411 : AOI22_X2 port map( A1 => n13680, A2 => n922, B1 => n28886, B2 => 
                           n13582, ZN => n16085);
   U6822 : INV_X4 port map( I => n4568, ZN => n26167);
   U21313 : INV_X4 port map( I => n24114, ZN => n17068);
   U4832 : AOI22_X2 port map( A1 => n18413, A2 => n18845, B1 => n18730, B2 => 
                           n18412, ZN => n30336);
   U23716 : AOI21_X1 port map( A1 => n20244, A2 => n20312, B => n936, ZN => 
                           n20245);
   U7844 : INV_X2 port map( I => n29303, ZN => n21396);
   U8726 : AOI21_X1 port map( A1 => n32009, A2 => n5677, B => n5676, ZN => 
                           n9840);
   U4555 : OAI22_X2 port map( A1 => n1290, A2 => n6478, B1 => n33320, B2 => 
                           n22588, ZN => n22438);
   U11797 : INV_X2 port map( I => n13610, ZN => n13609);
   U15013 : INV_X2 port map( I => n7809, ZN => n24260);
   U14744 : NAND2_X1 port map( A1 => n16921, A2 => n28415, ZN => n16920);
   U3129 : BUF_X2 port map( I => n13320, Z => n25967);
   U2660 : NAND2_X2 port map( A1 => n205, A2 => n204, ZN => n20204);
   U17965 : NAND2_X2 port map( A1 => n22478, A2 => n900, ZN => n6956);
   U1185 : NOR3_X2 port map( A1 => n31220, A2 => n517, A3 => n29084, ZN => 
                           n15885);
   U12980 : NAND2_X1 port map( A1 => n2070, A2 => n9146, ZN => n2069);
   U20432 : NOR2_X1 port map( A1 => n4067, A2 => n1281, ZN => n11058);
   U3953 : OR2_X1 port map( A1 => n8622, A2 => n3843, Z => n29050);
   U3877 : NAND2_X2 port map( A1 => n10031, A2 => n22876, ZN => n14667);
   U6166 : NOR2_X2 port map( A1 => n29239, A2 => n31428, ZN => n28933);
   U2621 : INV_X2 port map( I => n19195, ZN => n19606);
   U5458 : INV_X2 port map( I => n9759, ZN => n16193);
   U635 : INV_X4 port map( I => n510, ZN => n10686);
   U6610 : INV_X2 port map( I => n7680, ZN => n1379);
   U13315 : AND2_X2 port map( A1 => n20615, A2 => n9252, Z => n20362);
   U14493 : OAI21_X2 port map( A1 => n4339, A2 => n23103, B => n3600, ZN => 
                           n12790);
   U21037 : AOI21_X2 port map( A1 => n905, A2 => n1116, B => n12632, ZN => 
                           n13104);
   U8508 : NAND3_X2 port map( A1 => n7737, A2 => n11408, A3 => n32296, ZN => 
                           n7736);
   U16201 : INV_X2 port map( I => n28697, ZN => n3570);
   U12957 : INV_X2 port map( I => n11068, ZN => n20008);
   U2281 : OAI21_X2 port map( A1 => n17223, A2 => n12837, B => n15108, ZN => 
                           n8823);
   U26328 : NOR2_X2 port map( A1 => n22396, A2 => n22398, ZN => n5304);
   U17397 : NOR2_X2 port map( A1 => n33915, A2 => n6345, ZN => n11990);
   U11903 : NAND2_X2 port map( A1 => n15267, A2 => n12168, ZN => n3941);
   U49 : INV_X2 port map( I => n31407, ZN => n27183);
   U8786 : NAND2_X2 port map( A1 => n16538, A2 => n1189, ZN => n14614);
   U1410 : NAND3_X1 port map( A1 => n14943, A2 => n15400, A3 => n27455, ZN => 
                           n14942);
   U7641 : INV_X4 port map( I => n24328, ZN => n890);
   U3095 : NOR2_X2 port map( A1 => n26912, A2 => n16648, ZN => n15979);
   U5470 : AOI21_X2 port map( A1 => n18953, A2 => n17445, B => n18952, ZN => 
                           n18924);
   U14583 : NAND2_X2 port map( A1 => n14173, A2 => n19875, ZN => n20290);
   U5472 : AOI21_X2 port map( A1 => n19356, A2 => n6516, B => n19359, ZN => 
                           n14709);
   U1748 : NAND2_X1 port map( A1 => n29202, A2 => n29201, ZN => n20171);
   U23504 : NAND2_X2 port map( A1 => n33659, A2 => n23559, ZN => n16083);
   U13400 : INV_X4 port map( I => n27390, ZN => n17185);
   U1182 : INV_X4 port map( I => n21259, ZN => n28257);
   U20370 : OR2_X1 port map( A1 => n30010, A2 => n27970, Z => n7282);
   U551 : INV_X4 port map( I => n31220, ZN => n17021);
   U22594 : OAI22_X1 port map( A1 => n11156, A2 => n25916, B1 => n11155, B2 => 
                           n1206, ZN => n28331);
   U6751 : OAI21_X2 port map( A1 => n10310, A2 => n9958, B => n22574, ZN => 
                           n5453);
   U15796 : NAND2_X2 port map( A1 => n4385, A2 => n28806, ZN => n4384);
   U10093 : INV_X4 port map( I => n14812, ZN => n16916);
   U3426 : OR3_X1 port map( A1 => n1127, A2 => n9630, A3 => n3392, Z => n2548);
   U12826 : INV_X2 port map( I => n7672, ZN => n17341);
   U16264 : INV_X2 port map( I => n987, ZN => n27298);
   U6615 : AOI21_X2 port map( A1 => n29454, A2 => n1009, B => n2339, ZN => 
                           n2338);
   U8489 : INV_X2 port map( I => n20463, ZN => n16518);
   U3147 : BUF_X2 port map( I => n21210, Z => n16512);
   U7738 : INV_X2 port map( I => n5897, ZN => n1081);
   U4683 : INV_X2 port map( I => n10775, ZN => n26725);
   U12040 : NAND2_X2 port map( A1 => n5033, A2 => n946, ZN => n1767);
   U3643 : OR2_X1 port map( A1 => n8444, A2 => n17117, Z => n24878);
   U3812 : BUF_X2 port map( I => n8700, Z => n8010);
   U1664 : NOR2_X2 port map( A1 => n17263, A2 => n13154, ZN => n26375);
   U20496 : NAND2_X2 port map( A1 => n10389, A2 => n17186, ZN => n27994);
   U2421 : NAND2_X2 port map( A1 => n13884, A2 => n28203, ZN => n31859);
   U22350 : CLKBUF_X4 port map( I => n24254, Z => n28296);
   U3488 : NAND2_X2 port map( A1 => n33889, A2 => n33147, ZN => n2715);
   U8457 : NAND2_X2 port map( A1 => n1150, A2 => n16684, ZN => n1635);
   U7602 : AOI21_X2 port map( A1 => n18633, A2 => n1439, B => n17516, ZN => 
                           n15811);
   U10686 : NAND2_X1 port map( A1 => n16832, A2 => n1603, ZN => n1602);
   U16889 : INV_X2 port map( I => n13147, ZN => n23611);
   U13694 : INV_X2 port map( I => n19699, ZN => n19619);
   U14071 : OAI21_X2 port map( A1 => n732, A2 => n27228, B => n16318, ZN => 
                           n3112);
   U14352 : AOI21_X2 port map( A1 => n21645, A2 => n861, B => n27073, ZN => 
                           n27754);
   U290 : NAND2_X2 port map( A1 => n31419, A2 => n31421, ZN => n30509);
   U1826 : NAND2_X1 port map( A1 => n7462, A2 => n26320, ZN => n26956);
   U11035 : NAND2_X2 port map( A1 => n7066, A2 => n32678, ZN => n27486);
   U15623 : INV_X4 port map( I => n16458, ZN => n851);
   U223 : NAND2_X2 port map( A1 => n16704, A2 => n25561, ZN => n30561);
   U1492 : BUF_X4 port map( I => n34156, Z => n31030);
   U7215 : BUF_X4 port map( I => n20882, Z => n21163);
   U633 : NOR2_X2 port map( A1 => n8967, A2 => n22956, ZN => n28495);
   U8970 : OAI21_X2 port map( A1 => n32911, A2 => n5202, B => n25114, ZN => 
                           n9050);
   U4073 : AOI21_X2 port map( A1 => n24074, A2 => n24073, B => n27038, ZN => 
                           n9068);
   U17337 : INV_X2 port map( I => n27211, ZN => n27458);
   U6901 : INV_X2 port map( I => n17150, ZN => n893);
   U1814 : INV_X2 port map( I => n13327, ZN => n29338);
   U10582 : NOR2_X2 port map( A1 => n16443, A2 => n32178, ZN => n10397);
   U5496 : OAI21_X2 port map( A1 => n4518, A2 => n21078, B => n28502, ZN => 
                           n28501);
   U20099 : INV_X2 port map( I => n10337, ZN => n11814);
   U294 : NOR3_X1 port map( A1 => n30715, A2 => n1550, A3 => n28410, ZN => 
                           n3214);
   U311 : BUF_X4 port map( I => n15227, Z => n11200);
   U24479 : NAND3_X2 port map( A1 => n19962, A2 => n28767, A3 => n6748, ZN => 
                           n9978);
   U2668 : NAND2_X2 port map( A1 => n8593, A2 => n22642, ZN => n8332);
   U1122 : NOR2_X2 port map( A1 => n9721, A2 => n17841, ZN => n16189);
   U10383 : NAND2_X2 port map( A1 => n9807, A2 => n1079, ZN => n9806);
   U3801 : INV_X4 port map( I => n19332, ZN => n7732);
   U3181 : INV_X1 port map( I => n23925, ZN => n23763);
   U20730 : INV_X4 port map( I => n11744, ZN => n18923);
   U1085 : OAI21_X2 port map( A1 => n21187, A2 => n5239, B => n5238, ZN => 
                           n26413);
   U14426 : INV_X4 port map( I => n25889, ZN => n14805);
   U4980 : INV_X1 port map( I => n25865, ZN => n12266);
   U8947 : OAI22_X2 port map( A1 => n12164, A2 => n32911, B1 => n9936, B2 => 
                           n12165, ZN => n6629);
   U15009 : NAND2_X1 port map( A1 => n30283, A2 => n14759, ZN => n14758);
   U15008 : NOR2_X1 port map( A1 => n16100, A2 => n7203, ZN => n14759);
   U3821 : NAND3_X2 port map( A1 => n20872, A2 => n12902, A3 => n20311, ZN => 
                           n3402);
   U853 : NAND2_X2 port map( A1 => n16009, A2 => n14281, ZN => n14283);
   U3540 : INV_X4 port map( I => n19315, ZN => n2081);
   U3863 : OAI21_X2 port map( A1 => n7529, A2 => n7528, B => n22986, ZN => 
                           n29060);
   U1720 : NOR2_X2 port map( A1 => n18137, A2 => n20910, ZN => n18136);
   U14880 : OAI21_X1 port map( A1 => n3862, A2 => n23608, B => n3861, ZN => 
                           n23610);
   U16820 : AOI22_X2 port map( A1 => n7643, A2 => n10845, B1 => n19338, B2 => 
                           n5707, ZN => n7327);
   U4605 : AOI21_X2 port map( A1 => n25453, A2 => n17948, B => n11640, ZN => 
                           n25454);
   U7255 : INV_X2 port map( I => n18919, ZN => n18621);
   U1083 : BUF_X4 port map( I => n7753, Z => n230);
   U440 : NAND2_X1 port map( A1 => n29360, A2 => n22636, ZN => n15611);
   U2435 : AOI21_X2 port map( A1 => n10113, A2 => n21149, B => n2738, ZN => 
                           n8727);
   U748 : NAND2_X2 port map( A1 => n20200, A2 => n1789, ZN => n205);
   U6915 : OR2_X2 port map( A1 => n22591, A2 => n31549, Z => n11873);
   U5680 : INV_X4 port map( I => n13343, ZN => n794);
   U813 : OR2_X2 port map( A1 => n22656, A2 => n17899, Z => n13318);
   U1611 : CLKBUF_X4 port map( I => n18768, Z => n28757);
   U3809 : INV_X4 port map( I => n1736, ZN => n1329);
   U8606 : BUF_X2 port map( I => n9201, Z => n2166);
   U1589 : NAND2_X2 port map( A1 => n5535, A2 => n25337, ZN => n5534);
   U1266 : BUF_X4 port map( I => n6255, Z => n26471);
   U17386 : NAND2_X1 port map( A1 => n12192, A2 => n12193, ZN => n30469);
   U5010 : BUF_X2 port map( I => n12763, Z => n29323);
   U8011 : NAND2_X2 port map( A1 => n22522, A2 => n27638, ZN => n10389);
   U3055 : INV_X1 port map( I => n17503, ZN => n22752);
   U1552 : OAI22_X2 port map( A1 => n3313, A2 => n18106, B1 => n9191, B2 => 
                           n10571, ZN => n3312);
   U11365 : OAI22_X2 port map( A1 => n26904, A2 => n8825, B1 => n11276, B2 => 
                           n21818, ZN => n6699);
   U7018 : INV_X2 port map( I => n24874, ZN => n17787);
   U10749 : INV_X1 port map( I => n17579, ZN => n10498);
   U15377 : NAND2_X2 port map( A1 => n11892, A2 => n10354, ZN => n5140);
   U592 : INV_X4 port map( I => n21651, ZN => n15371);
   U8728 : NOR2_X2 port map( A1 => n22795, A2 => n33007, ZN => n13120);
   U8364 : OAI22_X2 port map( A1 => n18859, A2 => n18543, B1 => n18854, B2 => 
                           n18855, ZN => n18417);
   U3058 : AOI21_X2 port map( A1 => n14231, A2 => n1633, B => n1887, ZN => 
                           n1524);
   U5751 : BUF_X4 port map( I => n15329, Z => n27875);
   U3385 : NAND3_X1 port map( A1 => n13981, A2 => n11096, A3 => n13982, ZN => 
                           n31090);
   U166 : NAND2_X2 port map( A1 => n23982, A2 => n24246, ZN => n13633);
   U6968 : NAND2_X2 port map( A1 => n24325, A2 => n24328, ZN => n24246);
   U18955 : NAND2_X2 port map( A1 => n19844, A2 => n10086, ZN => n7309);
   U21506 : NOR2_X2 port map( A1 => n31097, A2 => n19923, ZN => n4648);
   U9883 : OAI21_X2 port map( A1 => n16029, A2 => n16346, B => n940, ZN => 
                           n2492);
   U2675 : NAND2_X2 port map( A1 => n1874, A2 => n16323, ZN => n9807);
   U14139 : INV_X2 port map( I => n21532, ZN => n30678);
   U4852 : NAND2_X2 port map( A1 => n27738, A2 => n12540, ZN => n5059);
   U261 : INV_X1 port map( I => n29268, ZN => n13291);
   U23826 : INV_X2 port map( I => n17143, ZN => n18701);
   U1397 : NOR2_X1 port map( A1 => n31906, A2 => n26774, ZN => n5869);
   U12156 : NAND2_X1 port map( A1 => n8860, A2 => n28056, ZN => n12192);
   U1899 : NOR2_X2 port map( A1 => n11075, A2 => n28345, ZN => n30743);
   U15092 : NAND2_X1 port map( A1 => n14209, A2 => n16231, ZN => n8122);
   U17244 : NOR2_X2 port map( A1 => n12221, A2 => n423, ZN => n6447);
   U10772 : INV_X2 port map( I => n9328, ZN => n3241);
   U1897 : NOR2_X2 port map( A1 => n747, A2 => n30288, ZN => n16973);
   U11423 : OAI21_X2 port map( A1 => n18106, A2 => n18035, B => n7723, ZN => 
                           n7722);
   U22287 : OAI21_X1 port map( A1 => n1132, A2 => n21811, B => n31627, ZN => 
                           n11167);
   U2867 : NAND3_X2 port map( A1 => n434, A2 => n14449, A3 => n433, ZN => 
                           n30199);
   U8113 : INV_X2 port map( I => n22225, ZN => n10650);
   U14089 : NOR2_X1 port map( A1 => n24329, A2 => n24328, ZN => n30186);
   U4930 : NAND2_X1 port map( A1 => n28261, A2 => n20546, ZN => n20547);
   U3145 : AOI21_X2 port map( A1 => n15611, A2 => n16240, B => n15609, ZN => 
                           n15608);
   U2945 : NAND2_X2 port map( A1 => n2877, A2 => n23055, ZN => n4845);
   U16746 : INV_X2 port map( I => n14619, ZN => n14745);
   U21720 : AOI22_X2 port map( A1 => n31120, A2 => n17483, B1 => n17482, B2 => 
                           n772, ZN => n9747);
   U19305 : NOR2_X2 port map( A1 => n31722, A2 => n28691, ZN => n9973);
   U10648 : OAI21_X2 port map( A1 => n13879, A2 => n17612, B => n30980, ZN => 
                           n13878);
   U13153 : NAND3_X2 port map( A1 => n16261, A2 => n16262, A3 => n2229, ZN => 
                           n16747);
   U4453 : BUF_X2 port map( I => n2256, Z => n27694);
   U4569 : NAND2_X2 port map( A1 => n28840, A2 => n15169, ZN => n20430);
   U1948 : INV_X2 port map( I => n30663, ZN => n30937);
   U4584 : AND2_X1 port map( A1 => n15057, A2 => n10708, Z => n14644);
   U10286 : INV_X4 port map( I => n6985, ZN => n13592);
   U96 : OR2_X2 port map( A1 => n8542, A2 => n13050, Z => n25874);
   U17725 : BUF_X4 port map( I => n639, Z => n30529);
   U1115 : INV_X2 port map( I => n14594, ZN => n30115);
   U18692 : NAND2_X1 port map( A1 => n30661, A2 => n30660, ZN => n13707);
   U11739 : NOR2_X1 port map( A1 => n7872, A2 => n20615, ZN => n6797);
   U2037 : OAI22_X2 port map( A1 => n8739, A2 => n18815, B1 => n18639, B2 => 
                           n9118, ZN => n4843);
   U5088 : INV_X1 port map( I => n10757, ZN => n12281);
   U6796 : NOR2_X2 port map( A1 => n708, A2 => n28160, ZN => n10138);
   U15401 : OAI21_X1 port map( A1 => n23042, A2 => n17930, B => n808, ZN => 
                           n13121);
   U11350 : INV_X2 port map( I => n21496, ZN => n21713);
   U12524 : INV_X1 port map( I => n11513, ZN => n14483);
   U14874 : NAND2_X1 port map( A1 => n21483, A2 => n1327, ZN => n21484);
   U20853 : NAND2_X1 port map( A1 => n21427, A2 => n33215, ZN => n14598);
   U3256 : NAND3_X2 port map( A1 => n1492, A2 => n1382, A3 => n19205, ZN => 
                           n1491);
   U9702 : INV_X4 port map( I => n29314, ZN => n22992);
   U10870 : NOR2_X1 port map( A1 => n28141, A2 => n15885, ZN => n31889);
   U264 : CLKBUF_X4 port map( I => n17037, Z => n16957);
   U212 : BUF_X4 port map( I => n25382, Z => n31149);
   U71 : INV_X4 port map( I => n25546, ZN => n12864);
   U2516 : NAND2_X2 port map( A1 => n11895, A2 => n22435, ZN => n2522);
   U18827 : NOR2_X2 port map( A1 => n6176, A2 => n2217, ZN => n8274);
   U17240 : INV_X4 port map( I => n10724, ZN => n30448);
   U1636 : INV_X4 port map( I => n14213, ZN => n1182);
   U768 : BUF_X4 port map( I => n4084, Z => n29648);
   U345 : NAND2_X2 port map( A1 => n28745, A2 => n28744, ZN => n4481);
   U3612 : INV_X1 port map( I => n7880, ZN => n31509);
   U1554 : NAND2_X1 port map( A1 => n30471, A2 => n15898, ZN => n26720);
   U3854 : INV_X2 port map( I => n25, ZN => n17955);
   U1688 : BUF_X2 port map( I => n20401, Z => n27785);
   U1150 : BUF_X4 port map( I => n29258, Z => n2551);
   U14873 : INV_X2 port map( I => n18198, ZN => n12290);
   U5860 : OR2_X1 port map( A1 => n26881, A2 => n13300, Z => n13562);
   U7184 : INV_X4 port map( I => n505, ZN => n5239);
   U7900 : INV_X4 port map( I => n7915, ZN => n8547);
   U8482 : INV_X4 port map( I => n27504, ZN => n29258);
   U7235 : OR2_X1 port map( A1 => n8314, A2 => n17960, Z => n29424);
   U5312 : INV_X2 port map( I => n31810, ZN => n16271);
   U8070 : INV_X2 port map( I => n22589, ZN => n22584);
   U22583 : INV_X4 port map( I => n28329, ZN => n2023);
   U1883 : CLKBUF_X4 port map( I => n15960, Z => n400);
   U4772 : NAND2_X1 port map( A1 => n5494, A2 => n30832, ZN => n12788);
   U1526 : NAND3_X1 port map( A1 => n17270, A2 => n26800, A3 => n16762, ZN => 
                           n29899);
   U6189 : NAND2_X2 port map( A1 => n15211, A2 => n14159, ZN => n28438);
   U6230 : NAND2_X2 port map( A1 => n1057, A2 => n18721, ZN => n6203);
   U21203 : INV_X2 port map( I => n16570, ZN => n14034);
   U10975 : NOR2_X2 port map( A1 => n16927, A2 => n22760, ZN => n16926);
   U5445 : NAND2_X1 port map( A1 => n9173, A2 => n20143, ZN => n7820);
   U4186 : BUF_X2 port map( I => n8277, Z => n28091);
   U14680 : AOI21_X2 port map( A1 => n11013, A2 => n20052, B => n3769, ZN => 
                           n6931);
   U3287 : BUF_X4 port map( I => n18028, Z => n27801);
   U485 : INV_X4 port map( I => n11895, ZN => n1298);
   U352 : NAND2_X2 port map( A1 => n8058, A2 => n18077, ZN => n13109);
   U16168 : OR2_X1 port map( A1 => n30988, A2 => n17271, Z => n17272);
   U10696 : NOR2_X2 port map( A1 => n8654, A2 => n11653, ZN => n3983);
   U7156 : NAND3_X2 port map( A1 => n21192, A2 => n26542, A3 => n33949, ZN => 
                           n8046);
   U2104 : NAND2_X2 port map( A1 => n20520, A2 => n5460, ZN => n73);
   U9351 : NOR2_X2 port map( A1 => n14157, A2 => n7179, ZN => n14773);
   U1659 : NOR2_X1 port map( A1 => n29409, A2 => n19792, ZN => n30572);
   U10000 : NAND2_X2 port map( A1 => n18667, A2 => n26518, ZN => n8211);
   U967 : AOI21_X2 port map( A1 => n909, A2 => n22427, B => n22537, ZN => 
                           n14388);
   U4427 : AOI22_X1 port map( A1 => n17802, A2 => n6476, B1 => n17801, B2 => 
                           n16868, ZN => n17800);
   U8111 : INV_X1 port map( I => n13553, ZN => n1004);
   U7434 : INV_X4 port map( I => n12408, ZN => n3790);
   U5650 : OAI21_X2 port map( A1 => n22635, A2 => n22640, B => n4511, ZN => 
                           n4510);
   U15070 : NAND3_X2 port map( A1 => n1243, A2 => n24193, A3 => n31918, ZN => 
                           n23990);
   U8769 : AOI21_X2 port map( A1 => n26036, A2 => n8273, B => n26397, ZN => 
                           n27391);
   U6984 : BUF_X2 port map( I => n8480, Z => n27211);
   U13505 : NOR2_X1 port map( A1 => n30124, A2 => n2764, ZN => n31021);
   U5753 : NAND2_X2 port map( A1 => n17568, A2 => n17567, ZN => n22961);
   U11507 : INV_X1 port map( I => n29908, ZN => n565);
   U8612 : NAND2_X2 port map( A1 => n26751, A2 => n8237, ZN => n8717);
   U7441 : NAND2_X2 port map( A1 => n18668, A2 => n18669, ZN => n8237);
   U5080 : INV_X2 port map( I => n3723, ZN => n15798);
   U16250 : NAND2_X1 port map( A1 => n31968, A2 => n17236, ZN => n7035);
   U516 : INV_X2 port map( I => n22121, ZN => n1305);
   U6746 : AOI21_X2 port map( A1 => n26347, A2 => n22425, B => n14728, ZN => 
                           n22603);
   U829 : NAND2_X2 port map( A1 => n16665, A2 => n28915, ZN => n26347);
   U4041 : BUF_X2 port map( I => n10303, Z => n22546);
   U20479 : NOR2_X1 port map( A1 => n28614, A2 => n31174, ZN => n7440);
   U2413 : NOR2_X2 port map( A1 => n4318, A2 => n15550, ZN => n13052);
   U1813 : INV_X2 port map( I => n871, ZN => n7460);
   U5023 : NOR2_X2 port map( A1 => n23930, A2 => n29269, ZN => n23538);
   U13660 : NAND2_X2 port map( A1 => n17726, A2 => n8834, ZN => n31560);
   U19562 : AND2_X2 port map( A1 => n8386, A2 => n32051, Z => n18878);
   U708 : INV_X2 port map( I => n12315, ZN => n22807);
   U6636 : NAND2_X2 port map( A1 => n18760, A2 => n18759, ZN => n15281);
   U4085 : NAND2_X2 port map( A1 => n6249, A2 => n6248, ZN => n23594);
   U15979 : NAND2_X2 port map( A1 => n11232, A2 => n17832, ZN => n7651);
   U10893 : INV_X2 port map( I => n8786, ZN => n8415);
   U8953 : NAND2_X2 port map( A1 => n16024, A2 => n32911, ZN => n9936);
   U11201 : OR2_X2 port map( A1 => n22599, A2 => n16432, Z => n22510);
   U23068 : NOR2_X2 port map( A1 => n4113, A2 => n27090, ZN => n22775);
   U1966 : CLKBUF_X4 port map( I => n19206, Z => n4202);
   U6838 : OAI21_X2 port map( A1 => n22993, A2 => n22992, B => n30388, ZN => 
                           n22997);
   U5653 : BUF_X4 port map( I => n22978, Z => n8990);
   U8603 : NAND3_X2 port map( A1 => n26384, A2 => n17880, A3 => n26383, ZN => 
                           n26589);
   U25107 : NAND2_X2 port map( A1 => n22563, A2 => n14034, ZN => n22564);
   U15040 : AOI21_X2 port map( A1 => n27314, A2 => n15084, B => n24983, ZN => 
                           n15223);
   U1848 : NAND2_X2 port map( A1 => n23940, A2 => n26965, ZN => n13678);
   U153 : INV_X2 port map( I => n24436, ZN => n718);
   U1484 : AOI22_X2 port map( A1 => n1490, A2 => n27970, B1 => n19242, B2 => 
                           n1494, ZN => n26293);
   U12836 : AND2_X1 port map( A1 => n13354, A2 => n33789, Z => n26836);
   U15827 : INV_X2 port map( I => n20310, ZN => n1154);
   U1004 : INV_X4 port map( I => n22435, ZN => n31636);
   U16891 : INV_X2 port map( I => n7463, ZN => n11235);
   U5715 : INV_X1 port map( I => n522, ZN => n29336);
   U11050 : NOR2_X2 port map( A1 => n26628, A2 => n13677, ZN => n27044);
   U473 : INV_X2 port map( I => n18098, ZN => n22474);
   U4240 : BUF_X4 port map( I => n15411, Z => n1883);
   U15295 : NAND3_X1 port map( A1 => n17742, A2 => n17743, A3 => n17741, ZN => 
                           n30583);
   U18159 : NOR3_X2 port map( A1 => n31007, A2 => n21642, A3 => n32613, ZN => 
                           n12274);
   U14981 : NAND2_X2 port map( A1 => n25399, A2 => n1700, ZN => n25402);
   U24680 : NOR2_X2 port map( A1 => n20563, A2 => n17329, ZN => n20285);
   U14095 : NOR2_X2 port map( A1 => n32788, A2 => n15137, ZN => n7437);
   U53 : NOR2_X2 port map( A1 => n15531, A2 => n15530, ZN => n15529);
   U11126 : NAND2_X2 port map( A1 => n7398, A2 => n10630, ZN => n6455);
   U12629 : NAND2_X1 port map( A1 => n26808, A2 => n15971, ZN => n9166);
   U6549 : INV_X2 port map( I => n20008, ZN => n1359);
   U6062 : NAND2_X2 port map( A1 => n10897, A2 => n14915, ZN => n15546);
   U23220 : NAND2_X1 port map( A1 => n15418, A2 => n15416, ZN => n28444);
   U655 : INV_X4 port map( I => n758, ZN => n23104);
   U11520 : OAI21_X2 port map( A1 => n15632, A2 => n12027, B => n31826, ZN => 
                           n15631);
   U14770 : OAI22_X2 port map( A1 => n25470, A2 => n25490, B1 => n25479, B2 => 
                           n25487, ZN => n25492);
   U3783 : INV_X2 port map( I => n27741, ZN => n7873);
   U6286 : INV_X2 port map( I => n18261, ZN => n23100);
   U14868 : NAND2_X2 port map( A1 => n25479, A2 => n25488, ZN => n25463);
   U1934 : NOR2_X2 port map( A1 => n19267, A2 => n19268, ZN => n2098);
   U417 : NAND2_X2 port map( A1 => n27163, A2 => n23872, ZN => n31528);
   U1435 : BUF_X2 port map( I => n21442, Z => n16180);
   U9691 : NAND2_X2 port map( A1 => n17939, A2 => n32457, ZN => n3211);
   U8339 : OAI21_X2 port map( A1 => n31729, A2 => n29574, B => n29573, ZN => 
                           n17939);
   U24760 : OAI21_X1 port map( A1 => n17200, A2 => n17199, B => n25467, ZN => 
                           n31492);
   U4259 : INV_X4 port map( I => n5225, ZN => n16466);
   U16121 : NAND2_X1 port map( A1 => n2052, A2 => n19782, ZN => n19791);
   U5460 : INV_X2 port map( I => n20010, ZN => n1167);
   U22924 : BUF_X4 port map( I => n14624, Z => n28386);
   U3604 : INV_X2 port map( I => n23300, ZN => n23414);
   U6876 : NAND2_X2 port map( A1 => n4408, A2 => n976, ZN => n5417);
   U17074 : NOR3_X2 port map( A1 => n28625, A2 => n30793, A3 => n27386, ZN => 
                           n4980);
   U3281 : NOR3_X2 port map( A1 => n9817, A2 => n1019, A3 => n9816, ZN => 
                           n29221);
   U16610 : INV_X2 port map( I => n14156, ZN => n18637);
   U9000 : BUF_X2 port map( I => n15777, Z => n11716);
   U10988 : NOR2_X2 port map( A1 => n29242, A2 => n28680, ZN => n22988);
   U24731 : NAND3_X2 port map( A1 => n15468, A2 => n33154, A3 => n28899, ZN => 
                           n20619);
   U3090 : INV_X2 port map( I => n15123, ZN => n23033);
   U24127 : BUF_X4 port map( I => n20103, Z => n28600);
   U1505 : CLKBUF_X4 port map( I => n19101, Z => n6511);
   U18259 : AOI21_X2 port map( A1 => n1246, A2 => n24311, B => n7481, ZN => 
                           n7480);
   U10887 : OAI22_X1 port map( A1 => n6035, A2 => n3202, B1 => n3201, B2 => 
                           n1107, ZN => n3200);
   U10427 : NAND3_X1 port map( A1 => n29116, A2 => n30047, A3 => n25462, ZN => 
                           n25458);
   U14911 : NAND2_X2 port map( A1 => n31883, A2 => n24154, ZN => n5367);
   U857 : NOR2_X2 port map( A1 => n2471, A2 => n22926, ZN => n9335);
   U6707 : INV_X4 port map( I => n16732, ZN => n956);
   U7652 : INV_X4 port map( I => n18131, ZN => n18815);
   U20835 : NAND2_X2 port map( A1 => n15638, A2 => n33730, ZN => n12847);
   U846 : INV_X4 port map( I => n19998, ZN => n7609);
   U26365 : OAI22_X2 port map( A1 => n19147, A2 => n15534, B1 => n1175, B2 => 
                           n1055, ZN => n5654);
   U1781 : INV_X1 port map( I => n20886, ZN => n29169);
   U22629 : INV_X2 port map( I => n19267, ZN => n15869);
   U6282 : INV_X1 port map( I => n22848, ZN => n15976);
   U3261 : BUF_X4 port map( I => n25894, Z => n4993);
   U2077 : CLKBUF_X4 port map( I => n6039, Z => n1125);
   U4465 : CLKBUF_X4 port map( I => n13232, Z => n2744);
   U6738 : NAND2_X2 port map( A1 => n23104, A2 => n23103, ZN => n26161);
   U4764 : NAND2_X2 port map( A1 => n24067, A2 => n10033, ZN => n3216);
   U21348 : NAND3_X2 port map( A1 => n28435, A2 => n27619, A3 => n27336, ZN => 
                           n31886);
   U17378 : AOI21_X2 port map( A1 => n17260, A2 => n71, B => n12398, ZN => 
                           n16977);
   U2697 : AND2_X2 port map( A1 => n16275, A2 => n515, Z => n21320);
   U15270 : INV_X2 port map( I => n32358, ZN => n6119);
   U15544 : BUF_X4 port map( I => n11570, Z => n15054);
   U8860 : BUF_X2 port map( I => Key(32), Z => n25428);
   U3968 : INV_X4 port map( I => n13905, ZN => n23760);
   U4233 : BUF_X2 port map( I => n14255, Z => n27577);
   U4266 : INV_X1 port map( I => n23827, ZN => n26775);
   U4706 : NAND2_X1 port map( A1 => n7756, A2 => n28257, ZN => n27245);
   U6077 : INV_X2 port map( I => n18892, ZN => n29683);
   U22274 : INV_X4 port map( I => n839, ZN => n24154);
   U3153 : OAI21_X2 port map( A1 => n19248, A2 => n3535, B => n19247, ZN => 
                           n19251);
   U9823 : NAND2_X2 port map( A1 => n7307, A2 => n19844, ZN => n3061);
   U6180 : NOR2_X1 port map( A1 => n23712, A2 => n17234, ZN => n14778);
   U3507 : BUF_X2 port map( I => n25696, Z => n16609);
   U15156 : NAND3_X1 port map( A1 => n1555, A2 => n9258, A3 => n27462, ZN => 
                           n30779);
   U16574 : NAND3_X2 port map( A1 => n22686, A2 => n33964, A3 => n22685, ZN => 
                           n31902);
   U1067 : AOI21_X2 port map( A1 => n11713, A2 => n17445, B => n8192, ZN => 
                           n11178);
   U17214 : NOR3_X2 port map( A1 => n32831, A2 => n13703, A3 => n13525, ZN => 
                           n6216);
   U22560 : NAND2_X2 port map( A1 => n20484, A2 => n31009, ZN => n28324);
   U10139 : AOI22_X2 port map( A1 => n18470, A2 => n18007, B1 => n18469, B2 => 
                           n18006, ZN => n18473);
   U13278 : AOI21_X2 port map( A1 => n13730, A2 => n31826, B => n6520, ZN => 
                           n3888);
   U12586 : NOR2_X1 port map( A1 => n15041, A2 => n12843, ZN => n3035);
   U84 : NAND2_X2 port map( A1 => n11696, A2 => n11697, ZN => n11695);
   U21458 : OAI21_X2 port map( A1 => n13036, A2 => n32143, B => n29602, ZN => 
                           n13035);
   U14192 : INV_X2 port map( I => n11516, ZN => n13521);
   U7833 : NOR2_X2 port map( A1 => n26282, A2 => n18033, ZN => n18032);
   U3594 : NAND2_X2 port map( A1 => n8770, A2 => n7218, ZN => n20576);
   U14799 : NAND3_X2 port map( A1 => n7803, A2 => n8033, A3 => n8107, ZN => 
                           n7550);
   U5904 : INV_X2 port map( I => n31906, ZN => n19960);
   U14044 : NAND2_X2 port map( A1 => n16834, A2 => n26542, ZN => n27016);
   U11557 : OAI21_X2 port map( A1 => n21426, A2 => n13286, B => n14168, ZN => 
                           n16834);
   U15050 : INV_X2 port map( I => n26724, ZN => n17828);
   U8987 : INV_X2 port map( I => n2023, ZN => n26416);
   U888 : OAI21_X2 port map( A1 => n25, A2 => n22621, B => n995, ZN => n22624);
   U11040 : OAI21_X2 port map( A1 => n22024, A2 => n16170, B => n2258, ZN => 
                           n2257);
   U4370 : AOI22_X2 port map( A1 => n11924, A2 => n29180, B1 => n21531, B2 => 
                           n8886, ZN => n31244);
   U5894 : BUF_X2 port map( I => n19601, Z => n19914);
   U5652 : BUF_X2 port map( I => n7012, Z => n26884);
   U4045 : NOR2_X2 port map( A1 => n18846, A2 => n17184, ZN => n18413);
   U2215 : BUF_X4 port map( I => n16209, Z => n100);
   U6086 : NAND2_X1 port map( A1 => n6287, A2 => n10651, ZN => n4520);
   U1203 : NAND2_X2 port map( A1 => n8941, A2 => n28126, ZN => n8940);
   U542 : OAI21_X2 port map( A1 => n21794, A2 => n21792, B => n30549, ZN => 
                           n11560);
   U25504 : NAND3_X1 port map( A1 => n24701, A2 => n11366, A3 => n25406, ZN => 
                           n24704);
   U10366 : NAND2_X1 port map( A1 => n6824, A2 => n6822, ZN => n8743);
   U3012 : INV_X4 port map( I => n15278, ZN => n8817);
   U11232 : CLKBUF_X4 port map( I => n19744, Z => n29876);
   U22907 : OAI21_X2 port map( A1 => n25160, A2 => n32553, B => n25159, ZN => 
                           n25163);
   U18993 : AOI22_X2 port map( A1 => n25173, A2 => n7765, B1 => n8929, B2 => 
                           n25158, ZN => n25159);
   U1110 : AOI22_X2 port map( A1 => n19421, A2 => n29156, B1 => n19420, B2 => 
                           n19868, ZN => n12705);
   U11167 : NAND2_X1 port map( A1 => n29863, A2 => n5937, ZN => n5935);
   U15136 : OAI22_X2 port map( A1 => n11706, A2 => n22690, B1 => n8944, B2 => 
                           n32194, ZN => n6943);
   U16965 : NAND2_X2 port map( A1 => n355, A2 => n22690, ZN => n8944);
   U10991 : NAND2_X2 port map( A1 => n6371, A2 => n6370, ZN => n6369);
   U663 : AOI21_X2 port map( A1 => n26868, A2 => n14188, B => n30904, ZN => 
                           n6371);
   U20735 : INV_X2 port map( I => n11765, ZN => n11923);
   U9840 : NOR2_X2 port map( A1 => n29774, A2 => n20627, ZN => n7836);
   U5267 : INV_X2 port map( I => n15063, ZN => n27275);
   U16179 : OAI21_X2 port map( A1 => n7765, A2 => n25175, B => n25174, ZN => 
                           n25177);
   U10158 : OAI21_X1 port map( A1 => n882, A2 => n14213, B => n12663, ZN => 
                           n9046);
   U19699 : BUF_X4 port map( I => n27807, Z => n30817);
   U4071 : NAND2_X2 port map( A1 => n15068, A2 => n13601, ZN => n23995);
   U14839 : NOR2_X2 port map( A1 => n32890, A2 => n23807, ZN => n13578);
   U18599 : AOI22_X2 port map( A1 => n9316, A2 => n27077, B1 => n9315, B2 => 
                           n27818, ZN => n9314);
   U359 : BUF_X4 port map( I => n13472, Z => n7068);
   U15977 : NAND2_X2 port map( A1 => n27367, A2 => n11232, ZN => n26679);
   U22597 : NAND2_X2 port map( A1 => n8862, A2 => n950, ZN => n19329);
   U24851 : AOI22_X2 port map( A1 => n21190, A2 => n21189, B1 => n33649, B2 => 
                           n21321, ZN => n21191);
   U17638 : AOI21_X2 port map( A1 => n18366, A2 => n18367, B => n13254, ZN => 
                           n27509);
   U5703 : BUF_X2 port map( I => n15617, Z => n2471);
   U22925 : INV_X2 port map( I => n14605, ZN => n17382);
   U3917 : BUF_X4 port map( I => n21693, Z => n27635);
   U4904 : BUF_X4 port map( I => n18310, Z => n14651);
   U6391 : OAI21_X2 port map( A1 => n6954, A2 => n6953, B => n1168, ZN => n6952
                           );
   U14473 : AND2_X2 port map( A1 => n11707, A2 => n16462, Z => n18634);
   U9767 : NOR2_X1 port map( A1 => n16176, A2 => n782, ZN => n5735);
   U15621 : NAND2_X2 port map( A1 => n16611, A2 => n25149, ZN => n6204);
   U16070 : NAND2_X2 port map( A1 => n26900, A2 => n27457, ZN => n30320);
   U1388 : OAI21_X1 port map( A1 => n8348, A2 => n8349, B => n9270, ZN => n6945
                           );
   U2073 : INV_X2 port map( I => n31773, ZN => n8756);
   U1620 : NAND2_X1 port map( A1 => n29995, A2 => n29994, ZN => n29993);
   U12381 : NAND2_X1 port map( A1 => n20259, A2 => n817, ZN => n29995);
   U541 : INV_X1 port map( I => n4281, ZN => n23593);
   U11735 : INV_X2 port map( I => n20328, ZN => n11808);
   U21396 : NAND2_X2 port map( A1 => n17993, A2 => n1350, ZN => n17992);
   U6447 : BUF_X4 port map( I => n19260, Z => n28379);
   U11933 : CLKBUF_X4 port map( I => n15476, Z => n15381);
   U16750 : AOI21_X2 port map( A1 => n13597, A2 => n30960, B => n33675, ZN => 
                           n5620);
   U16956 : INV_X2 port map( I => n21317, ZN => n27367);
   U7298 : NOR2_X2 port map( A1 => n33302, A2 => n32477, ZN => n3240);
   U4822 : NAND2_X2 port map( A1 => n17512, A2 => n28324, ZN => n17511);
   U21713 : INV_X2 port map( I => n17916, ZN => n22610);
   U2353 : NOR2_X1 port map( A1 => n23058, A2 => n17462, ZN => n28783);
   U9126 : NAND2_X1 port map( A1 => n12568, A2 => n23896, ZN => n3950);
   U6990 : NAND2_X1 port map( A1 => n5140, A2 => n10216, ZN => n10388);
   U453 : INV_X2 port map( I => n32926, ZN => n15853);
   U15964 : NAND2_X1 port map( A1 => n19803, A2 => n20006, ZN => n27196);
   U8995 : NOR2_X2 port map( A1 => n33120, A2 => n25697, ZN => n3774);
   U556 : NOR2_X2 port map( A1 => n13597, A2 => n15851, ZN => n13619);
   U5584 : NOR2_X1 port map( A1 => n23595, A2 => n11567, ZN => n16969);
   U5151 : INV_X2 port map( I => n16625, ZN => n941);
   U22755 : AOI22_X1 port map( A1 => n17464, A2 => n30234, B1 => n22879, B2 => 
                           n22880, ZN => n17463);
   U17330 : NAND2_X2 port map( A1 => n2225, A2 => n7287, ZN => n27457);
   U94 : OR2_X2 port map( A1 => n1215, A2 => n25260, Z => n6280);
   U12095 : NAND2_X1 port map( A1 => n6207, A2 => n11122, ZN => n8628);
   U14752 : NAND2_X2 port map( A1 => n23791, A2 => n14460, ZN => n9522);
   U3613 : OR2_X1 port map( A1 => n13693, A2 => n20329, Z => n20551);
   U1338 : NAND3_X1 port map( A1 => n7386, A2 => n6309, A3 => n13291, ZN => 
                           n6308);
   U184 : OR2_X2 port map( A1 => n18151, A2 => n18150, Z => n25591);
   U122 : AOI21_X2 port map( A1 => n6551, A2 => n25332, B => n15880, ZN => 
                           n31786);
   U198 : INV_X1 port map( I => n15528, ZN => n25411);
   U4156 : OAI21_X2 port map( A1 => n13578, A2 => n6132, B => n31208, ZN => 
                           n6131);
   U1874 : INV_X1 port map( I => n16, ZN => n29656);
   U11432 : OAI22_X2 port map( A1 => n1785, A2 => n1329, B1 => n32248, B2 => 
                           n21061, ZN => n1456);
   U9703 : NAND2_X1 port map( A1 => n31350, A2 => n19291, ZN => n31349);
   U5752 : NAND2_X1 port map( A1 => n31871, A2 => n10344, ZN => n10343);
   U360 : INV_X2 port map( I => n31437, ZN => n1274);
   U9347 : OAI22_X2 port map( A1 => n4812, A2 => n22467, B1 => n14376, B2 => 
                           n28865, ZN => n4811);
   U613 : NAND2_X1 port map( A1 => n13316, A2 => n13315, ZN => n13314);
   U19960 : NOR2_X1 port map( A1 => n30852, A2 => n12747, ZN => n5248);
   U15076 : CLKBUF_X8 port map( I => n30978, Z => n30769);
   U8615 : CLKBUF_X4 port map( I => n706, Z => n25980);
   U3155 : CLKBUF_X4 port map( I => n16333, Z => n9797);
   U7655 : BUF_X2 port map( I => Key(35), Z => n25131);
   U22987 : INV_X2 port map( I => n14798, ZN => n17313);
   U4239 : INV_X4 port map( I => n1385, ZN => n1047);
   U11580 : NOR2_X1 port map( A1 => n28648, A2 => n986, ZN => n26688);
   U10973 : NAND3_X2 port map( A1 => n13597, A2 => n23093, A3 => n15039, ZN => 
                           n23094);
   U1530 : INV_X4 port map( I => n9191, ZN => n18106);
   U5450 : INV_X4 port map( I => n20100, ZN => n937);
   U1282 : AOI21_X2 port map( A1 => n15551, A2 => n16980, B => n16979, ZN => 
                           n16978);
   U3177 : NOR2_X2 port map( A1 => n4205, A2 => n4204, ZN => n5270);
   U2703 : BUF_X2 port map( I => n20939, Z => n21357);
   U17911 : NOR2_X1 port map( A1 => n5342, A2 => n27383, ZN => n30984);
   U7553 : NAND2_X2 port map( A1 => n18289, A2 => n18288, ZN => n18290);
   U8413 : INV_X2 port map( I => n21085, ZN => n11948);
   U1614 : NAND2_X2 port map( A1 => n73, A2 => n14876, ZN => n31878);
   U19347 : NAND2_X1 port map( A1 => n23613, A2 => n29839, ZN => n30754);
   U6874 : BUF_X2 port map( I => n29273, Z => n31796);
   U21118 : NAND2_X2 port map( A1 => n17466, A2 => n32242, ZN => n12912);
   U9500 : NOR2_X2 port map( A1 => n9206, A2 => n9204, ZN => n5474);
   U11984 : BUF_X2 port map( I => n4314, Z => n3727);
   U21314 : NAND2_X1 port map( A1 => n17563, A2 => n17562, ZN => n17561);
   U10847 : INV_X4 port map( I => n5381, ZN => n9223);
   U18711 : NAND2_X2 port map( A1 => n31007, A2 => n7553, ZN => n21554);
   U7148 : INV_X2 port map( I => n17316, ZN => n180);
   U5636 : OAI22_X2 port map( A1 => n6225, A2 => n10529, B1 => n24216, B2 => 
                           n24109, ZN => n10531);
   U68 : NAND2_X1 port map( A1 => n27099, A2 => n9050, ZN => n27731);
   U5084 : INV_X2 port map( I => n18539, ZN => n14346);
   U377 : NAND2_X2 port map( A1 => n26950, A2 => n8178, ZN => n27826);
   U3780 : OAI21_X2 port map( A1 => n20097, A2 => n1041, B => n8182, ZN => 
                           n8181);
   U1295 : INV_X2 port map( I => n26363, ZN => n28471);
   U20140 : OR2_X2 port map( A1 => n20208, A2 => n20207, Z => n10460);
   U21244 : NAND3_X1 port map( A1 => n19948, A2 => n20068, A3 => n20067, ZN => 
                           n16084);
   U7846 : NOR2_X2 port map( A1 => n23947, A2 => n29198, ZN => n6272);
   U10957 : INV_X2 port map( I => n23088, ZN => n14602);
   U11700 : NAND2_X1 port map( A1 => n20159, A2 => n20333, ZN => n12150);
   U20901 : OAI21_X1 port map( A1 => n909, A2 => n5597, B => n14388, ZN => 
                           n14387);
   U4577 : AND3_X1 port map( A1 => n10845, A2 => n34103, A3 => n6532, Z => 
                           n10846);
   U19901 : NAND2_X2 port map( A1 => n3180, A2 => n12886, ZN => n9540);
   U1638 : NAND2_X2 port map( A1 => n8454, A2 => n29867, ZN => n11760);
   U18580 : NAND2_X2 port map( A1 => n30640, A2 => n30639, ZN => n22424);
   U10566 : OR2_X1 port map( A1 => n9789, A2 => n11100, Z => n17853);
   U1183 : INV_X2 port map( I => n20803, ZN => n1343);
   U21309 : AOI21_X2 port map( A1 => n22483, A2 => n9910, B => n29158, ZN => 
                           n15835);
   U1880 : INV_X2 port map( I => n19395, ZN => n19740);
   U20218 : NOR3_X2 port map( A1 => n15591, A2 => n15590, A3 => n20497, ZN => 
                           n4061);
   U11185 : OAI21_X1 port map( A1 => n22549, A2 => n27416, B => n22315, ZN => 
                           n22326);
   U2948 : INV_X4 port map( I => n11970, ZN => n950);
   U9365 : NAND2_X2 port map( A1 => n12334, A2 => n17960, ZN => n12333);
   U4083 : INV_X1 port map( I => n24251, ZN => n1092);
   U3242 : INV_X2 port map( I => n17439, ZN => n21222);
   U20810 : BUF_X2 port map( I => n20657, Z => n21079);
   U3781 : INV_X1 port map( I => n20097, ZN => n20061);
   U14397 : NOR2_X1 port map( A1 => n31514, A2 => n2906, ZN => n30624);
   U21302 : INV_X1 port map( I => n18167, ZN => n17730);
   U14672 : NOR2_X1 port map( A1 => n2023, A2 => n23794, ZN => n30251);
   U14366 : NAND3_X2 port map( A1 => n31072, A2 => n28626, A3 => n28316, ZN => 
                           n3465);
   U14999 : NOR2_X1 port map( A1 => n25593, A2 => n13763, ZN => n8246);
   U10138 : OAI21_X2 port map( A1 => n18815, A2 => n18515, B => n9211, ZN => 
                           n8478);
   U8776 : INV_X4 port map( I => n18761, ZN => n18288);
   U24628 : AOI22_X2 port map( A1 => n20160, A2 => n20002, B1 => n742, B2 => 
                           n31072, ZN => n20003);
   U21284 : NAND2_X1 port map( A1 => n15490, A2 => n26965, ZN => n13669);
   U16414 : NAND2_X2 port map( A1 => n32012, A2 => n10629, ZN => n27294);
   U20599 : NOR2_X1 port map( A1 => n10381, A2 => n11435, ZN => n11437);
   U679 : NOR2_X2 port map( A1 => n22529, A2 => n28661, ZN => n28660);
   U11248 : INV_X2 port map( I => n10946, ZN => n4228);
   U3102 : NAND2_X2 port map( A1 => n21378, A2 => n26798, ZN => n13621);
   U1618 : NOR2_X2 port map( A1 => n18805, A2 => n18806, ZN => n18807);
   U409 : NAND2_X2 port map( A1 => n23684, A2 => n28091, ZN => n26529);
   U5882 : BUF_X2 port map( I => n9322, Z => n30755);
   U15593 : NAND2_X2 port map( A1 => n18383, A2 => n18515, ZN => n4206);
   U1251 : AOI21_X2 port map( A1 => n15053, A2 => n20243, B => n26232, ZN => 
                           n20246);
   U18867 : NAND2_X1 port map( A1 => n10886, A2 => n8433, ZN => n11179);
   U25792 : INV_X2 port map( I => n30231, ZN => n28801);
   U9903 : NOR2_X2 port map( A1 => n2391, A2 => n4215, ZN => n10683);
   U3114 : INV_X1 port map( I => n23087, ZN => n26243);
   U3113 : INV_X1 port map( I => n20037, ZN => n28826);
   U5143 : INV_X4 port map( I => n14559, ZN => n1358);
   U10904 : NAND2_X1 port map( A1 => n13914, A2 => n3162, ZN => n3161);
   U20382 : NOR2_X2 port map( A1 => n10964, A2 => n10966, ZN => n10965);
   U3441 : OAI22_X2 port map( A1 => n19365, A2 => n27921, B1 => n19109, B2 => 
                           n5907, ZN => n7185);
   U471 : AND2_X2 port map( A1 => n13413, A2 => n27883, Z => n23650);
   U18475 : NOR2_X2 port map( A1 => n5248, A2 => n30627, ZN => n28139);
   U14398 : NOR2_X1 port map( A1 => n30318, A2 => n7272, ZN => n7271);
   U16031 : INV_X1 port map( I => n34108, ZN => n11182);
   U14732 : NAND2_X1 port map( A1 => n27432, A2 => n27431, ZN => n28652);
   U11807 : INV_X1 port map( I => n17494, ZN => n24617);
   U13772 : NOR2_X2 port map( A1 => n30155, A2 => n20141, ZN => n15592);
   U17578 : OR2_X2 port map( A1 => n6681, A2 => n16756, Z => n21285);
   U2069 : INV_X1 port map( I => n34110, ZN => n30697);
   U22658 : INV_X2 port map( I => n3503, ZN => n28338);
   U14407 : NOR2_X1 port map( A1 => n10651, A2 => n24061, ZN => n10653);
   U5330 : NAND2_X1 port map( A1 => n1890, A2 => n30867, ZN => n4095);
   U6243 : INV_X2 port map( I => n26550, ZN => n16592);
   U9660 : NOR2_X2 port map( A1 => n833, A2 => n24667, ZN => n28246);
   U685 : INV_X1 port map( I => n21253, ZN => n17437);
   U7283 : INV_X1 port map( I => n17829, ZN => n21252);
   U17043 : INV_X2 port map( I => n25582, ZN => n27637);
   U3975 : BUF_X2 port map( I => n5306, Z => n2539);
   U4053 : CLKBUF_X4 port map( I => n29470, Z => n29305);
   U14738 : NOR2_X1 port map( A1 => n29018, A2 => n2847, ZN => n28281);
   U16287 : NAND2_X2 port map( A1 => n19124, A2 => n27021, ZN => n12270);
   U4609 : CLKBUF_X4 port map( I => n19796, Z => n20052);
   U13428 : NAND3_X1 port map( A1 => n15280, A2 => n22838, A3 => n13191, ZN => 
                           n30853);
   U1621 : OAI21_X1 port map( A1 => n13760, A2 => n33301, B => n29983, ZN => 
                           n4535);
   U9597 : NOR2_X1 port map( A1 => n12372, A2 => n21121, ZN => n12371);
   U18197 : INV_X2 port map( I => n31918, ZN => n27592);
   U15265 : INV_X1 port map( I => n11707, ZN => n27142);
   U13160 : INV_X1 port map( I => n1577, ZN => n1581);
   U7359 : AOI22_X2 port map( A1 => n870, A2 => n26368, B1 => n16811, B2 => 
                           n20044, ZN => n15198);
   U428 : NAND3_X2 port map( A1 => n17726, A2 => n16424, A3 => n11960, ZN => 
                           n23835);
   U650 : AOI21_X2 port map( A1 => n31712, A2 => n22701, B => n23081, ZN => 
                           n22704);
   U16686 : NAND3_X2 port map( A1 => n30831, A2 => n25600, A3 => n25602, ZN => 
                           n27308);
   U4676 : CLKBUF_X4 port map( I => n17431, Z => n27560);
   U23919 : INV_X4 port map( I => n16933, ZN => n21251);
   U9290 : INV_X2 port map( I => n6359, ZN => n29659);
   U12823 : NOR2_X1 port map( A1 => n15098, A2 => n23575, ZN => n15097);
   U4170 : AOI21_X2 port map( A1 => n21686, A2 => n21551, B => n861, ZN => 
                           n9493);
   U1656 : AOI21_X2 port map( A1 => n12699, A2 => n11999, B => n12651, ZN => 
                           n12650);
   U17431 : NOR2_X2 port map( A1 => n9549, A2 => n8422, ZN => n18369);
   U13658 : NOR2_X2 port map( A1 => n32087, A2 => n17132, ZN => n27008);
   U1176 : CLKBUF_X4 port map( I => n12561, Z => n26573);
   U11634 : NAND2_X1 port map( A1 => n20223, A2 => n2203, ZN => n2206);
   U9612 : NOR2_X1 port map( A1 => n5332, A2 => n29768, ZN => n30426);
   U5420 : INV_X2 port map( I => n12342, ZN => n1024);
   U1196 : BUF_X2 port map( I => n7294, Z => n28983);
   U8576 : NAND2_X2 port map( A1 => n14589, A2 => n8611, ZN => n13571);
   U4099 : INV_X1 port map( I => n7188, ZN => n12932);
   U930 : NAND2_X2 port map( A1 => n16570, A2 => n16556, ZN => n22560);
   U22823 : INV_X2 port map( I => n34156, ZN => n7673);
   U21992 : AOI21_X2 port map( A1 => n32378, A2 => n22474, B => n28225, ZN => 
                           n17935);
   U19914 : INV_X2 port map( I => n11637, ZN => n27901);
   U12833 : NOR2_X1 port map( A1 => n26837, A2 => n26836, ZN => n26835);
   U19689 : INV_X1 port map( I => n9549, ZN => n18782);
   U11867 : NOR2_X1 port map( A1 => n19897, A2 => n33743, ZN => n15259);
   U2092 : BUF_X2 port map( I => n17405, Z => n71);
   U7868 : INV_X2 port map( I => n23759, ZN => n6662);
   U10640 : NOR2_X2 port map( A1 => n22478, A2 => n32378, ZN => n21968);
   U9172 : NOR2_X2 port map( A1 => n7088, A2 => n2561, ZN => n13402);
   U22916 : INV_X2 port map( I => n14572, ZN => n16595);
   U8533 : NAND2_X1 port map( A1 => n26376, A2 => n12892, ZN => n12891);
   U13509 : AOI21_X1 port map( A1 => n2766, A2 => n2767, B => n31156, ZN => 
                           n30124);
   U14990 : OAI21_X2 port map( A1 => n10658, A2 => n17093, B => n4041, ZN => 
                           n21180);
   U6361 : INV_X1 port map( I => n6569, ZN => n1131);
   U25352 : NAND2_X2 port map( A1 => n23796, A2 => n14193, ZN => n23803);
   U3984 : AOI21_X1 port map( A1 => n19109, A2 => n6566, B => n6565, ZN => 
                           n6564);
   U1074 : NOR3_X2 port map( A1 => n3168, A2 => n5017, A3 => n1325, ZN => 
                           n29737);
   U18582 : NOR2_X2 port map( A1 => n7990, A2 => n28701, ZN => n9560);
   U4142 : BUF_X2 port map( I => n17204, Z => n6297);
   U7227 : AOI22_X2 port map( A1 => n20397, A2 => n7577, B1 => n20396, B2 => 
                           n20395, ZN => n26216);
   U22434 : OR2_X1 port map( A1 => n18187, A2 => n10080, Z => n437);
   U534 : AOI21_X1 port map( A1 => n12853, A2 => n13490, B => n12852, ZN => 
                           n12855);
   U19905 : NOR2_X2 port map( A1 => n27899, A2 => n10117, ZN => n10116);
   U23534 : OAI21_X2 port map( A1 => n8824, A2 => n8948, B => n8823, ZN => 
                           n8822);
   U886 : OAI21_X2 port map( A1 => n18985, A2 => n18984, B => n15378, ZN => 
                           n18986);
   U14077 : OAI21_X1 port map( A1 => n14667, A2 => n802, B => n22761, ZN => 
                           n12907);
   U7322 : INV_X4 port map( I => n17157, ZN => n23878);
   U12897 : INV_X4 port map( I => n15467, ZN => n17394);
   U4147 : INV_X4 port map( I => n8965, ZN => n909);
   U24153 : NAND2_X2 port map( A1 => n179, A2 => n21438, ZN => n20330);
   U20022 : NOR2_X1 port map( A1 => n30858, A2 => n25084, ZN => n25087);
   U5343 : INV_X2 port map( I => n13969, ZN => n13157);
   U23543 : NOR2_X2 port map( A1 => n28993, A2 => n31351, ZN => n7403);
   U3940 : NAND2_X2 port map( A1 => n7238, A2 => n349, ZN => n11153);
   U4745 : BUF_X2 port map( I => n21428, Z => n26542);
   U25326 : INV_X1 port map( I => n22143, ZN => n3041);
   U2613 : INV_X2 port map( I => n23942, ZN => n757);
   U16233 : NOR2_X1 port map( A1 => n7344, A2 => n7343, ZN => n29106);
   U1518 : INV_X2 port map( I => n16309, ZN => n21867);
   U8963 : OAI21_X2 port map( A1 => n5897, A2 => n17787, B => n15084, ZN => 
                           n16387);
   U4730 : NOR2_X1 port map( A1 => n21415, A2 => n21416, ZN => n27010);
   U1969 : NAND2_X2 port map( A1 => n948, A2 => n19078, ZN => n31539);
   U17809 : AOI22_X2 port map( A1 => n18525, A2 => n19256, B1 => n26969, B2 => 
                           n33608, ZN => n18527);
   U14353 : NAND2_X1 port map( A1 => n4774, A2 => n3421, ZN => n12576);
   U6009 : BUF_X2 port map( I => Key(115), Z => n16472);
   U4300 : BUF_X2 port map( I => Key(66), Z => n24623);
   U4311 : BUF_X2 port map( I => Key(145), Z => n16680);
   U7658 : BUF_X2 port map( I => Key(98), Z => n25208);
   U7061 : CLKBUF_X2 port map( I => Key(111), Z => n25610);
   U7671 : BUF_X2 port map( I => Key(97), Z => n24991);
   U10222 : BUF_X2 port map( I => Key(175), Z => n16381);
   U4909 : CLKBUF_X2 port map( I => Key(144), Z => n16575);
   U7663 : BUF_X2 port map( I => Key(106), Z => n16602);
   U10251 : BUF_X2 port map( I => Key(92), Z => n16671);
   U8861 : BUF_X2 port map( I => Key(19), Z => n25071);
   U4280 : CLKBUF_X2 port map( I => Key(33), Z => n25722);
   U16647 : CLKBUF_X2 port map( I => n494, Z => n30371);
   U6150 : CLKBUF_X4 port map( I => n18429, Z => n18510);
   U10203 : INV_X1 port map( I => n16561, ZN => n1394);
   U10198 : INV_X1 port map( I => n24804, ZN => n1410);
   U508 : INV_X1 port map( I => n25476, ZN => n1404);
   U5528 : CLKBUF_X4 port map( I => n18357, Z => n18797);
   U3412 : CLKBUF_X4 port map( I => n16596, Z => n1430);
   U15934 : BUF_X2 port map( I => n18777, Z => n12863);
   U25448 : INV_X1 port map( I => n31574, ZN => n28231);
   U21786 : CLKBUF_X4 port map( I => n18392, Z => n18711);
   U12235 : CLKBUF_X2 port map( I => n18498, Z => n16435);
   U8812 : INV_X2 port map( I => n17813, ZN => n5677);
   U6094 : CLKBUF_X2 port map( I => n16249, Z => n29514);
   U15066 : CLKBUF_X4 port map( I => n17558, Z => n5327);
   U12168 : OAI21_X1 port map( A1 => n18428, A2 => n18832, B => n18698, ZN => 
                           n17254);
   U3577 : INV_X1 port map( I => n489, ZN => n958);
   U16380 : INV_X1 port map( I => n19295, ZN => n15859);
   U12092 : NAND2_X1 port map( A1 => n10640, A2 => n10639, ZN => n7285);
   U12096 : INV_X1 port map( I => n3986, ZN => n3985);
   U1568 : CLKBUF_X4 port map( I => n2692, Z => n26603);
   U10044 : INV_X2 port map( I => n31254, ZN => n1376);
   U5168 : BUF_X2 port map( I => n9553, Z => n3535);
   U12701 : INV_X2 port map( I => n30039, ZN => n5610);
   U1550 : CLKBUF_X2 port map( I => n19149, Z => n25961);
   U15279 : CLKBUF_X4 port map( I => n19335, Z => n8212);
   U10070 : INV_X1 port map( I => n11477, ZN => n19326);
   U5014 : CLKBUF_X2 port map( I => n4392, Z => n29093);
   U3278 : BUF_X2 port map( I => n6763, Z => n28157);
   U24058 : INV_X2 port map( I => n16801, ZN => n11444);
   U7775 : NOR2_X1 port map( A1 => n19228, A2 => n19357, ZN => n13389);
   U2698 : OAI21_X1 port map( A1 => n1049, A2 => n7687, B => n11477, ZN => 
                           n11113);
   U23186 : AOI21_X1 port map( A1 => n2582, A2 => n30937, B => n19053, ZN => 
                           n8433);
   U1912 : INV_X1 port map( I => n19323, ZN => n31618);
   U17052 : NOR2_X1 port map( A1 => n18971, A2 => n1177, ZN => n6024);
   U17184 : OAI21_X1 port map( A1 => n27420, A2 => n29245, B => n19263, ZN => 
                           n9237);
   U15100 : AND2_X1 port map( A1 => n18753, A2 => n17339, Z => n12271);
   U3417 : INV_X1 port map( I => n19013, ZN => n19010);
   U25845 : NOR2_X1 port map( A1 => n19067, A2 => n31618, ZN => n3133);
   U8257 : NAND2_X1 port map( A1 => n30936, A2 => n9839, ZN => n2583);
   U3480 : NAND2_X1 port map( A1 => n4594, A2 => n34040, ZN => n415);
   U12847 : NAND2_X1 port map( A1 => n2598, A2 => n6795, ZN => n30062);
   U24473 : NAND3_X1 port map( A1 => n19352, A2 => n19351, A3 => n19350, ZN => 
                           n19353);
   U4969 : CLKBUF_X4 port map( I => n253, Z => n28601);
   U23579 : BUF_X2 port map( I => n19672, Z => n31361);
   U7818 : CLKBUF_X4 port map( I => n30193, Z => n29515);
   U24480 : INV_X1 port map( I => n19550, ZN => n19379);
   U4854 : INV_X2 port map( I => n20064, ZN => n20096);
   U5463 : BUF_X2 port map( I => n20098, Z => n2606);
   U22086 : INV_X1 port map( I => n13941, ZN => n19849);
   U19175 : BUF_X2 port map( I => n13922, Z => n28704);
   U4520 : AND2_X1 port map( A1 => n31951, A2 => n10860, Z => n20153);
   U841 : INV_X1 port map( I => n8421, ZN => n20032);
   U26148 : CLKBUF_X2 port map( I => n4577, Z => n31684);
   U1371 : NOR2_X1 port map( A1 => n33419, A2 => n16346, ZN => n27787);
   U4610 : CLKBUF_X2 port map( I => n19419, Z => n19886);
   U5459 : INV_X1 port map( I => n27748, ZN => n4441);
   U1803 : CLKBUF_X4 port map( I => n26733, Z => n30375);
   U6430 : CLKBUF_X4 port map( I => n27748, Z => n26130);
   U1417 : INV_X2 port map( I => n26733, ZN => n27938);
   U6017 : CLKBUF_X1 port map( I => n17559, Z => n29944);
   U3952 : CLKBUF_X2 port map( I => n12241, Z => n27624);
   U9880 : NAND2_X1 port map( A1 => n9031, A2 => n27938, ZN => n9030);
   U9911 : NOR2_X1 port map( A1 => n9748, A2 => n4163, ZN => n4162);
   U7356 : NAND2_X1 port map( A1 => n12119, A2 => n18126, ZN => n1681);
   U19159 : INV_X1 port map( I => n5470, ZN => n27788);
   U1347 : NAND2_X1 port map( A1 => n9149, A2 => n19840, ZN => n27764);
   U6031 : BUF_X2 port map( I => n871, Z => n31103);
   U11817 : NAND2_X1 port map( A1 => n6223, A2 => n6221, ZN => n19898);
   U16217 : INV_X1 port map( I => n570, ZN => n20095);
   U11898 : INV_X1 port map( I => n19888, ZN => n4972);
   U25900 : CLKBUF_X4 port map( I => n34153, Z => n28876);
   U11858 : NAND2_X1 port map( A1 => n19798, A2 => n29040, ZN => n6645);
   U9870 : OAI21_X1 port map( A1 => n19990, A2 => n1035, B => n9661, ZN => 
                           n9660);
   U21584 : NAND2_X1 port map( A1 => n7461, A2 => n7460, ZN => n28153);
   U5977 : NAND2_X1 port map( A1 => n20094, A2 => n12669, ZN => n10926);
   U16811 : NAND2_X1 port map( A1 => n19828, A2 => n4587, ZN => n28209);
   U26295 : CLKBUF_X4 port map( I => n7102, Z => n31721);
   U21600 : NAND2_X1 port map( A1 => n31106, A2 => n28767, ZN => n27279);
   U15592 : OR2_X1 port map( A1 => n4637, A2 => n4636, Z => n4635);
   U21598 : INV_X2 port map( I => n6444, ZN => n20078);
   U21583 : NAND2_X1 port map( A1 => n28154, A2 => n28153, ZN => n1976);
   U24325 : NAND2_X1 port map( A1 => n31443, A2 => n20154, ZN => n26543);
   U24412 : CLKBUF_X2 port map( I => n31668, Z => n31454);
   U5863 : NOR2_X1 port map( A1 => n17497, A2 => n26585, ZN => n17693);
   U6303 : CLKBUF_X4 port map( I => n20560, Z => n16684);
   U15346 : BUF_X1 port map( I => n9403, Z => n31156);
   U10545 : INV_X1 port map( I => n28390, ZN => n29792);
   U4416 : CLKBUF_X4 port map( I => n28064, Z => n27755);
   U8467 : CLKBUF_X4 port map( I => n20371, Z => n15898);
   U4897 : AOI21_X1 port map( A1 => n27846, A2 => n12351, B => n12832, ZN => 
                           n2903);
   U1706 : CLKBUF_X4 port map( I => n17544, Z => n28812);
   U5436 : CLKBUF_X4 port map( I => n16515, Z => n28085);
   U13991 : AND2_X1 port map( A1 => n20395, A2 => n7292, Z => n7290);
   U18155 : NAND2_X1 port map( A1 => n31811, A2 => n20606, ZN => n20610);
   U8036 : OR2_X1 port map( A1 => n15282, A2 => n3944, Z => n17531);
   U7187 : CLKBUF_X2 port map( I => n12563, Z => n26343);
   U15776 : INV_X2 port map( I => n9352, ZN => n13768);
   U8463 : INV_X2 port map( I => n20529, ZN => n1155);
   U15811 : INV_X1 port map( I => n20288, ZN => n4964);
   U22262 : NOR2_X1 port map( A1 => n17425, A2 => n266, ZN => n17424);
   U18863 : INV_X1 port map( I => n14683, ZN => n20251);
   U8890 : CLKBUF_X2 port map( I => n8903, Z => n29628);
   U1667 : INV_X1 port map( I => n12227, ZN => n12226);
   U8452 : INV_X1 port map( I => n20604, ZN => n3751);
   U22416 : OAI21_X1 port map( A1 => n1349, A2 => n1351, B => n11312, ZN => 
                           n31211);
   U9805 : NAND2_X1 port map( A1 => n13537, A2 => n9688, ZN => n13760);
   U11638 : NOR2_X1 port map( A1 => n3746, A2 => n17322, ZN => n4241);
   U1206 : OAI21_X1 port map( A1 => n13090, A2 => n20494, B => n20493, ZN => 
                           n13089);
   U11711 : NOR2_X1 port map( A1 => n27020, A2 => n6797, ZN => n8325);
   U2313 : NAND2_X1 port map( A1 => n120, A2 => n20199, ZN => n1788);
   U11725 : NAND2_X1 port map( A1 => n20321, A2 => n1032, ZN => n10063);
   U16452 : INV_X1 port map( I => n4586, ZN => n30340);
   U21631 : NAND2_X1 port map( A1 => n31112, A2 => n31111, ZN => n20177);
   U5930 : NAND2_X1 port map( A1 => n30464, A2 => n15951, ZN => n8959);
   U11622 : NAND2_X1 port map( A1 => n2206, A2 => n2204, ZN => n12479);
   U1344 : NAND2_X1 port map( A1 => n15257, A2 => n15256, ZN => n19910);
   U11690 : INV_X1 port map( I => n7978, ZN => n20580);
   U728 : OAI21_X1 port map( A1 => n20230, A2 => n20562, B => n3352, ZN => 
                           n20233);
   U18510 : AOI21_X1 port map( A1 => n30632, A2 => n20493, B => n17318, ZN => 
                           n16858);
   U9244 : NAND2_X1 port map( A1 => n29651, A2 => n26089, ZN => n30446);
   U22344 : CLKBUF_X2 port map( I => n20900, Z => n28295);
   U17282 : OAI21_X1 port map( A1 => n16758, A2 => n20505, B => n20504, ZN => 
                           n13092);
   U1852 : CLKBUF_X4 port map( I => n6857, Z => n15);
   U11275 : INV_X1 port map( I => n29652, ZN => n20804);
   U4201 : CLKBUF_X2 port map( I => n20913, Z => n3799);
   U3140 : CLKBUF_X4 port map( I => n7330, Z => n25969);
   U26653 : CLKBUF_X2 port map( I => n20924, Z => n31884);
   U1192 : INV_X1 port map( I => n4680, ZN => n28897);
   U22845 : CLKBUF_X2 port map( I => n12748, Z => n31277);
   U4805 : INV_X1 port map( I => n20648, ZN => n26692);
   U1184 : INV_X1 port map( I => n12618, ZN => n28584);
   U1199 : NAND2_X1 port map( A1 => n2649, A2 => n17554, ZN => n2648);
   U22328 : NAND2_X1 port map( A1 => n31189, A2 => n31188, ZN => n3403);
   U23585 : INV_X1 port map( I => n31423, ZN => n20979);
   U5883 : NAND2_X1 port map( A1 => n30083, A2 => n8579, ZN => n8578);
   U23503 : INV_X2 port map( I => n17218, ZN => n16072);
   U1481 : BUF_X2 port map( I => n11733, Z => n29207);
   U7072 : CLKBUF_X2 port map( I => n21184, Z => n17466);
   U2723 : CLKBUF_X4 port map( I => n21070, Z => n164);
   U5849 : INV_X1 port map( I => n9351, ZN => n9405);
   U4792 : CLKBUF_X2 port map( I => n21454, Z => n27912);
   U5879 : CLKBUF_X4 port map( I => n4755, Z => n30988);
   U7286 : CLKBUF_X2 port map( I => n17829, Z => n28037);
   U2502 : CLKBUF_X4 port map( I => n21232, Z => n16526);
   U3387 : CLKBUF_X4 port map( I => n11942, Z => n7430);
   U7214 : INV_X2 port map( I => n16512, ZN => n922);
   U5499 : CLKBUF_X4 port map( I => n21330, Z => n8378);
   U5146 : INV_X2 port map( I => n16906, ZN => n21209);
   U7152 : INV_X1 port map( I => n6192, ZN => n11487);
   U24777 : INV_X1 port map( I => n21202, ZN => n20791);
   U3996 : OR2_X1 port map( A1 => n12044, A2 => n31114, Z => n21114);
   U7208 : CLKBUF_X4 port map( I => n515, Z => n4381);
   U5529 : INV_X2 port map( I => n13255, ZN => n21211);
   U21131 : INV_X1 port map( I => n21297, ZN => n15335);
   U20884 : NOR2_X1 port map( A1 => n922, A2 => n13582, ZN => n13581);
   U26457 : CLKBUF_X2 port map( I => n505, Z => n31760);
   U2195 : CLKBUF_X4 port map( I => n10558, Z => n4683);
   U18974 : NAND2_X1 port map( A1 => n20705, A2 => n12756, ZN => n30699);
   U4716 : INV_X1 port map( I => n3889, ZN => n21077);
   U8340 : INV_X1 port map( I => n21398, ZN => n16755);
   U17350 : CLKBUF_X2 port map( I => n21253, Z => n27462);
   U3043 : CLKBUF_X4 port map( I => n11063, Z => n9721);
   U15576 : INV_X1 port map( I => n8041, ZN => n6826);
   U11442 : NAND2_X1 port map( A1 => n6743, A2 => n13896, ZN => n6501);
   U16200 : NAND2_X1 port map( A1 => n7757, A2 => n21259, ZN => n27246);
   U1316 : NAND2_X1 port map( A1 => n30654, A2 => n21093, ZN => n4919);
   U15982 : NOR2_X1 port map( A1 => n12348, A2 => n12017, ZN => n1687);
   U4701 : OR2_X1 port map( A1 => n21176, A2 => n21175, Z => n26468);
   U9655 : NOR2_X1 port map( A1 => n12243, A2 => n1331, ZN => n10093);
   U7953 : NAND2_X1 port map( A1 => n12507, A2 => n10730, ZN => n26302);
   U18990 : NAND2_X1 port map( A1 => n8267, A2 => n21147, ZN => n12018);
   U2874 : BUF_X2 port map( I => n9472, Z => n28729);
   U11368 : NAND2_X1 port map( A1 => n11152, A2 => n17217, ZN => n11149);
   U13769 : CLKBUF_X2 port map( I => n21738, Z => n30154);
   U9586 : INV_X1 port map( I => n2575, ZN => n21848);
   U2109 : CLKBUF_X4 port map( I => n13113, Z => n338);
   U1152 : NAND2_X1 port map( A1 => n21315, A2 => n8011, ZN => n9397);
   U8317 : INV_X2 port map( I => n21573, ZN => n6660);
   U3669 : OR2_X1 port map( A1 => n5795, A2 => n6669, Z => n21660);
   U5568 : INV_X1 port map( I => n21235, ZN => n4607);
   U3915 : CLKBUF_X2 port map( I => n8313, Z => n28895);
   U3037 : INV_X1 port map( I => n7182, ZN => n917);
   U1764 : INV_X2 port map( I => n16987, ZN => n4234);
   U1031 : CLKBUF_X2 port map( I => n4356, Z => n28387);
   U3401 : CLKBUF_X4 port map( I => n8790, Z => n396);
   U6613 : BUF_X1 port map( I => n21761, Z => n26443);
   U4176 : CLKBUF_X4 port map( I => n6669, Z => n6483);
   U22307 : NAND4_X1 port map( A1 => n13148, A2 => n13150, A3 => n13151, A4 => 
                           n13152, ZN => n21786);
   U7247 : AND2_X1 port map( A1 => n21779, A2 => n21743, Z => n29434);
   U608 : INV_X2 port map( I => n21592, ZN => n21793);
   U2944 : CLKBUF_X4 port map( I => n3539, Z => n276);
   U10651 : INV_X2 port map( I => n31085, ZN => n1136);
   U15183 : CLKBUF_X4 port map( I => n5016, Z => n27619);
   U6556 : NAND2_X1 port map( A1 => n1327, A2 => n21707, ZN => n5788);
   U3934 : INV_X1 port map( I => n21649, ZN => n16013);
   U13927 : NOR2_X1 port map( A1 => n1535, A2 => n21749, ZN => n1534);
   U1211 : AOI21_X1 port map( A1 => n21649, A2 => n21648, B => n31765, ZN => 
                           n28432);
   U21519 : OAI21_X1 port map( A1 => n21683, A2 => n26443, B => n14870, ZN => 
                           n14869);
   U23265 : NAND2_X1 port map( A1 => n1316, A2 => n1319, ZN => n15413);
   U17466 : NAND2_X1 port map( A1 => n913, A2 => n9286, ZN => n21125);
   U2288 : NAND2_X1 port map( A1 => n14730, A2 => n16165, ZN => n27759);
   U14838 : NOR2_X1 port map( A1 => n3048, A2 => n31202, ZN => n31201);
   U10425 : CLKBUF_X2 port map( I => n11458, Z => n26562);
   U21710 : NAND2_X1 port map( A1 => n12994, A2 => n12995, ZN => n31118);
   U1734 : INV_X1 port map( I => n28432, ZN => n28431);
   U18387 : NAND2_X1 port map( A1 => n30616, A2 => n26163, ZN => n275);
   U893 : INV_X2 port map( I => n21913, ZN => n28162);
   U12886 : INV_X2 port map( I => n26875, ZN => n8269);
   U25966 : CLKBUF_X2 port map( I => n22149, Z => n28926);
   U15748 : INV_X2 port map( I => n16893, ZN => n26957);
   U889 : CLKBUF_X4 port map( I => n22232, Z => n28730);
   U14920 : INV_X1 port map( I => n7545, ZN => n8359);
   U4971 : INV_X2 port map( I => n11166, ZN => n22239);
   U11220 : INV_X1 port map( I => n22144, ZN => n9311);
   U14293 : CLKBUF_X2 port map( I => n22367, Z => n30205);
   U22162 : INV_X2 port map( I => n28263, ZN => n629);
   U22049 : OR2_X1 port map( A1 => n9757, A2 => n31692, Z => n16986);
   U3950 : CLKBUF_X2 port map( I => n16710, Z => n9022);
   U6768 : INV_X2 port map( I => n628, ZN => n12496);
   U6688 : INV_X2 port map( I => n31914, ZN => n22637);
   U5804 : CLKBUF_X2 port map( I => n9871, Z => n8131);
   U5708 : BUF_X4 port map( I => n14514, Z => n10354);
   U11207 : CLKBUF_X2 port map( I => n21971, Z => n22489);
   U4474 : AND2_X1 port map( A1 => n9064, A2 => n32055, Z => n13079);
   U2471 : OR2_X1 port map( A1 => n8505, A2 => n6955, Z => n22475);
   U5781 : CLKBUF_X4 port map( I => n635, Z => n22557);
   U2839 : INV_X1 port map( I => n16986, ZN => n26367);
   U4568 : BUF_X2 port map( I => n5657, Z => n27959);
   U5645 : NAND2_X1 port map( A1 => n8912, A2 => n29903, ZN => n8911);
   U6343 : INV_X1 port map( I => n22683, ZN => n22686);
   U13805 : INV_X2 port map( I => n2858, ZN => n22647);
   U960 : NAND2_X1 port map( A1 => n22434, A2 => n701, ZN => n10243);
   U24655 : AOI21_X1 port map( A1 => n250, A2 => n5648, B => n1292, ZN => 
                           n31485);
   U9812 : INV_X1 port map( I => n22657, ZN => n31267);
   U2744 : INV_X1 port map( I => n30529, ZN => n11926);
   U903 : AOI21_X1 port map( A1 => n32007, A2 => n26046, B => n17394, ZN => 
                           n29758);
   U5669 : INV_X2 port map( I => n16647, ZN => n1001);
   U24078 : NAND2_X1 port map( A1 => n28592, A2 => n22595, ZN => n28681);
   U14388 : OAI21_X1 port map( A1 => n32042, A2 => n4560, B => n16334, ZN => 
                           n30215);
   U23023 : NAND2_X1 port map( A1 => n10654, A2 => n13525, ZN => n18062);
   U11051 : NOR2_X1 port map( A1 => n11615, A2 => n17631, ZN => n11614);
   U9960 : OAI21_X1 port map( A1 => n29736, A2 => n12840, B => n22648, ZN => 
                           n27307);
   U19955 : OAI21_X1 port map( A1 => n15322, A2 => n11895, B => n31636, ZN => 
                           n10071);
   U6952 : NAND2_X1 port map( A1 => n11243, A2 => n11245, ZN => n26925);
   U16957 : NAND2_X1 port map( A1 => n9108, A2 => n995, ZN => n6685);
   U4526 : INV_X2 port map( I => n9224, ZN => n13129);
   U11672 : INV_X1 port map( I => n31854, ZN => n22849);
   U19382 : NAND2_X1 port map( A1 => n22360, A2 => n1298, ZN => n30762);
   U3088 : BUF_X2 port map( I => n15243, Z => n27612);
   U4422 : BUF_X2 port map( I => n6798, Z => n28853);
   U5155 : CLKBUF_X2 port map( I => n22909, Z => n29328);
   U22235 : INV_X2 port map( I => n23053, ZN => n28277);
   U3436 : NAND2_X1 port map( A1 => n13129, A2 => n22945, ZN => n31825);
   U1750 : INV_X2 port map( I => n13191, ZN => n14420);
   U777 : CLKBUF_X4 port map( I => n5696, Z => n3163);
   U744 : CLKBUF_X4 port map( I => n14126, Z => n28680);
   U5352 : INV_X2 port map( I => n28942, ZN => n773);
   U6255 : OAI21_X1 port map( A1 => n6782, A2 => n26251, B => n6942, ZN => 
                           n10107);
   U11027 : NOR2_X1 port map( A1 => n14977, A2 => n31867, ZN => n7528);
   U21941 : CLKBUF_X2 port map( I => n22824, Z => n28214);
   U4451 : BUF_X2 port map( I => n16297, Z => n28330);
   U6268 : INV_X4 port map( I => n33675, ZN => n15851);
   U5013 : CLKBUF_X4 port map( I => n31637, Z => n29325);
   U10956 : OAI21_X1 port map( A1 => n22813, A2 => n4937, B => n17099, ZN => 
                           n4936);
   U18838 : INV_X1 port map( I => n11383, ZN => n22853);
   U2506 : NOR2_X1 port map( A1 => n32091, A2 => n22919, ZN => n2775);
   U13339 : NAND2_X1 port map( A1 => n1746, A2 => n1745, ZN => n4155);
   U8039 : NAND2_X1 port map( A1 => n27263, A2 => n26312, ZN => n26960);
   U4374 : INV_X1 port map( I => n27988, ZN => n27987);
   U2221 : INV_X1 port map( I => n22792, ZN => n29967);
   U23505 : NAND2_X1 port map( A1 => n4487, A2 => n4486, ZN => n28487);
   U11882 : NOR2_X1 port map( A1 => n30968, A2 => n30967, ZN => n30966);
   U10907 : NAND2_X1 port map( A1 => n2078, A2 => n2076, ZN => n5058);
   U10889 : NAND2_X1 port map( A1 => n3778, A2 => n13778, ZN => n13275);
   U2119 : CLKBUF_X2 port map( I => n5399, Z => n26915);
   U11644 : INV_X1 port map( I => n23461, ZN => n30274);
   U4326 : NAND2_X1 port map( A1 => n26311, A2 => n26590, ZN => n27701);
   U596 : INV_X1 port map( I => n23460, ZN => n2862);
   U10817 : INV_X1 port map( I => n663, ZN => n23853);
   U469 : CLKBUF_X4 port map( I => n22617, Z => n27455);
   U580 : CLKBUF_X4 port map( I => n17015, Z => n14974);
   U3504 : BUF_X4 port map( I => n22936, Z => n23778);
   U15236 : CLKBUF_X4 port map( I => n665, Z => n4069);
   U2441 : CLKBUF_X4 port map( I => n661, Z => n6869);
   U15391 : BUF_X2 port map( I => n23025, Z => n23775);
   U3503 : CLKBUF_X2 port map( I => n8838, Z => n313);
   U4810 : INV_X2 port map( I => n23575, ZN => n23939);
   U17418 : CLKBUF_X4 port map( I => n16534, Z => n27474);
   U483 : CLKBUF_X2 port map( I => n23719, Z => n16186);
   U18798 : INV_X2 port map( I => n8251, ZN => n11240);
   U4234 : BUF_X4 port map( I => n15399, Z => n1099);
   U5276 : NAND2_X1 port map( A1 => n23575, A2 => n15722, ZN => n12469);
   U578 : INV_X1 port map( I => n14133, ZN => n1255);
   U445 : NAND2_X1 port map( A1 => n23923, A2 => n11192, ZN => n17543);
   U262 : INV_X2 port map( I => n8270, ZN => n10145);
   U16796 : NAND2_X1 port map( A1 => n979, A2 => n14473, ZN => n17618);
   U3684 : CLKBUF_X4 port map( I => n15711, Z => n25987);
   U15843 : NAND2_X1 port map( A1 => n23653, A2 => n23746, ZN => n23777);
   U8874 : NAND2_X1 port map( A1 => n16186, A2 => n6869, ZN => n8372);
   U6879 : INV_X2 port map( I => n11240, ZN => n16388);
   U15293 : OR2_X1 port map( A1 => n23899, A2 => n32711, Z => n23704);
   U22620 : INV_X2 port map( I => n15623, ZN => n16343);
   U16075 : CLKBUF_X4 port map( I => n23945, Z => n27219);
   U16018 : NOR2_X1 port map( A1 => n12848, A2 => n8045, ZN => n27049);
   U14330 : NAND2_X1 port map( A1 => n16212, A2 => n16211, ZN => n28698);
   U17524 : NAND2_X1 port map( A1 => n7141, A2 => n7139, ZN => n23565);
   U6846 : NAND2_X1 port map( A1 => n17950, A2 => n17949, ZN => n3919);
   U21070 : AOI21_X1 port map( A1 => n23955, A2 => n15616, B => n23824, ZN => 
                           n14014);
   U6140 : AOI21_X1 port map( A1 => n18054, A2 => n9225, B => n28855, ZN => 
                           n24001);
   U13749 : AND2_X1 port map( A1 => n23353, A2 => n17088, Z => n29124);
   U9132 : OAI21_X1 port map( A1 => n12433, A2 => n978, B => n15351, ZN => 
                           n17490);
   U10764 : NAND2_X1 port map( A1 => n12592, A2 => n7781, ZN => n7780);
   U6159 : AND2_X1 port map( A1 => n16947, A2 => n7524, Z => n14907);
   U2325 : NAND2_X1 port map( A1 => n23308, A2 => n12603, ZN => n12602);
   U186 : INV_X2 port map( I => n24201, ZN => n738);
   U15711 : NOR2_X1 port map( A1 => n12974, A2 => n5373, ZN => n7407);
   U21849 : NAND2_X1 port map( A1 => n845, A2 => n8914, ZN => n3014);
   U4094 : INV_X1 port map( I => n10384, ZN => n7169);
   U10688 : NAND2_X1 port map( A1 => n13138, A2 => n13136, ZN => n8380);
   U5544 : CLKBUF_X2 port map( I => n24240, Z => n31862);
   U2791 : CLKBUF_X2 port map( I => n13623, Z => n11255);
   U12841 : CLKBUF_X2 port map( I => n6286, Z => n30061);
   U20942 : BUF_X2 port map( I => n3421, Z => n31002);
   U3204 : BUF_X2 port map( I => n9919, Z => n2444);
   U246 : INV_X2 port map( I => n24309, ZN => n28040);
   U3656 : INV_X1 port map( I => n15227, ZN => n24051);
   U10587 : NAND2_X1 port map( A1 => n23608, A2 => n794, ZN => n3861);
   U5489 : CLKBUF_X1 port map( I => n9146, Z => n29819);
   U15888 : CLKBUF_X4 port map( I => n24053, Z => n10381);
   U258 : CLKBUF_X4 port map( I => n11438, Z => n28691);
   U7758 : NAND2_X1 port map( A1 => n5914, A2 => n13260, ZN => n3255);
   U12931 : CLKBUF_X4 port map( I => n16643, Z => n8086);
   U3549 : AOI21_X1 port map( A1 => n7099, A2 => n24246, B => n28538, ZN => 
                           n7098);
   U10561 : INV_X1 port map( I => n14052, ZN => n8263);
   U17209 : NAND2_X1 port map( A1 => n13239, A2 => n13109, ZN => n13238);
   U15427 : AND3_X1 port map( A1 => n6773, A2 => n7729, A3 => n7727, Z => 
                           n27157);
   U11409 : OAI21_X1 port map( A1 => n17566, A2 => n33182, B => n305, ZN => 
                           n5000);
   U8546 : NAND2_X1 port map( A1 => n2398, A2 => n2400, ZN => n29924);
   U3025 : CLKBUF_X4 port map( I => n9300, Z => n4997);
   U17062 : NAND3_X1 port map( A1 => n24502, A2 => n24500, A3 => n24501, ZN => 
                           n30822);
   U277 : CLKBUF_X4 port map( I => n9708, Z => n29320);
   U13307 : CLKBUF_X2 port map( I => n5762, Z => n30104);
   U3379 : BUF_X2 port map( I => n24359, Z => n13050);
   U4059 : INV_X1 port map( I => n9120, ZN => n12676);
   U3645 : BUF_X2 port map( I => n17117, Z => n15046);
   U15256 : BUF_X4 port map( I => n24368, Z => n25707);
   U4038 : CLKBUF_X2 port map( I => n678, Z => n28958);
   U4055 : BUF_X2 port map( I => n25188, Z => n28591);
   U3221 : BUF_X2 port map( I => n25242, Z => n25977);
   U14574 : CLKBUF_X2 port map( I => n29278, Z => n30241);
   U25820 : INV_X2 port map( I => n24974, ZN => n28815);
   U23584 : CLKBUF_X4 port map( I => n25150, Z => n16293);
   U5260 : CLKBUF_X4 port map( I => n16659, Z => n29334);
   U156 : CLKBUF_X4 port map( I => n13427, Z => n1567);
   U4037 : CLKBUF_X2 port map( I => n25200, Z => n26432);
   U23995 : INV_X2 port map( I => n32652, ZN => n25025);
   U1946 : NOR2_X1 port map( A1 => n32872, A2 => n2642, ZN => n27757);
   U8943 : NAND2_X1 port map( A1 => n25868, A2 => n11716, ZN => n10066);
   U14510 : NOR2_X1 port map( A1 => n10890, A2 => n32760, ZN => n11082);
   U3586 : NAND2_X1 port map( A1 => n836, A2 => n11045, ZN => n24723);
   U16312 : NAND2_X1 port map( A1 => n10454, A2 => n25566, ZN => n27269);
   U5320 : NOR2_X1 port map( A1 => n30877, A2 => n30876, ZN => n31109);
   U21630 : NAND2_X1 port map( A1 => n3955, A2 => n24413, ZN => n31110);
   U7042 : CLKBUF_X4 port map( I => n17637, Z => n30935);
   U4309 : BUF_X2 port map( I => Key(69), Z => n25911);
   U8859 : BUF_X2 port map( I => Key(183), Z => n16672);
   U7666 : BUF_X2 port map( I => Key(75), Z => n25364);
   U4296 : CLKBUF_X2 port map( I => Key(110), Z => n25274);
   U6005 : BUF_X2 port map( I => Key(121), Z => n25091);
   U2282 : CLKBUF_X2 port map( I => Key(51), Z => n23239);
   U10244 : CLKBUF_X2 port map( I => Key(18), Z => n16464);
   U4285 : BUF_X2 port map( I => Key(7), Z => n24999);
   U4649 : BUF_X2 port map( I => Key(72), Z => n24804);
   U6122 : CLKBUF_X2 port map( I => n18860, Z => n31417);
   U24564 : INV_X1 port map( I => n19718, ZN => n25104);
   U12211 : CLKBUF_X2 port map( I => n18773, Z => n16522);
   U2065 : CLKBUF_X2 port map( I => n18228, Z => n30472);
   U1048 : CLKBUF_X4 port map( I => n18884, Z => n10669);
   U10121 : NOR2_X1 port map( A1 => n18653, A2 => n31542, ZN => n10640);
   U10102 : OAI21_X1 port map( A1 => n18796, A2 => n18795, B => n18799, ZN => 
                           n3986);
   U16024 : NAND2_X1 port map( A1 => n10220, A2 => n31972, ZN => n8645);
   U6064 : BUF_X2 port map( I => n18257, Z => n29715);
   U24266 : AND2_X1 port map( A1 => n19322, A2 => n19274, Z => n18415);
   U21526 : CLKBUF_X1 port map( I => n19224, Z => n28147);
   U6236 : CLKBUF_X1 port map( I => n19053, Z => n31108);
   U3021 : CLKBUF_X2 port map( I => n19149, Z => n25960);
   U20331 : CLKBUF_X4 port map( I => n2971, Z => n27965);
   U3969 : BUF_X2 port map( I => n27242, Z => n26350);
   U5004 : CLKBUF_X2 port map( I => n18626, Z => n28478);
   U3133 : OAI21_X1 port map( A1 => n32790, A2 => n19137, B => n744, ZN => 
                           n4594);
   U24444 : NAND2_X1 port map( A1 => n19189, A2 => n19257, ZN => n19190);
   U4992 : NAND2_X1 port map( A1 => n5082, A2 => n4405, ZN => n5083);
   U9910 : CLKBUF_X2 port map( I => n18109, Z => n29728);
   U11956 : NOR2_X1 port map( A1 => n3073, A2 => n6575, ZN => n3072);
   U4957 : CLKBUF_X2 port map( I => n29254, Z => n29013);
   U6033 : BUF_X2 port map( I => n18199, Z => n28183);
   U1867 : CLKBUF_X4 port map( I => n27808, Z => n31823);
   U4216 : INV_X2 port map( I => n17495, ZN => n939);
   U19604 : NOR2_X1 port map( A1 => n8616, A2 => n19451, ZN => n9379);
   U24583 : NAND2_X1 port map( A1 => n1168, A2 => n10340, ZN => n19823);
   U17250 : NAND2_X1 port map( A1 => n27938, A2 => n13994, ZN => n19805);
   U1831 : BUF_X2 port map( I => n20113, Z => n31715);
   U7390 : INV_X2 port map( I => n15192, ZN => n6644);
   U5985 : CLKBUF_X4 port map( I => n27070, Z => n29603);
   U3941 : CLKBUF_X2 port map( I => n20614, Z => n28527);
   U5394 : CLKBUF_X2 port map( I => n20634, Z => n2203);
   U3939 : INV_X2 port map( I => n20634, ZN => n20379);
   U3492 : CLKBUF_X2 port map( I => n816, Z => n420);
   U5936 : NAND2_X1 port map( A1 => n20258, A2 => n29603, ZN => n29994);
   U2847 : CLKBUF_X4 port map( I => n10717, Z => n1863);
   U5942 : BUF_X2 port map( I => n4460, Z => n30793);
   U1644 : NOR2_X1 port map( A1 => n20442, A2 => n1032, ZN => n30952);
   U4492 : NAND2_X1 port map( A1 => n1032, A2 => n18078, ZN => n28135);
   U1730 : CLKBUF_X4 port map( I => n9831, Z => n9688);
   U26483 : OAI21_X1 port map( A1 => n4964, A2 => n31776, B => n20174, ZN => 
                           n27611);
   U4060 : BUF_X2 port map( I => n8625, Z => n5141);
   U2085 : CLKBUF_X2 port map( I => n601, Z => n67);
   U5872 : CLKBUF_X2 port map( I => n21168, Z => n31874);
   U1497 : CLKBUF_X1 port map( I => n27503, Z => n27773);
   U2729 : BUF_X4 port map( I => n16784, Z => n28642);
   U4190 : CLKBUF_X4 port map( I => n18110, Z => n6408);
   U5856 : NAND2_X2 port map( A1 => n810, A2 => n27773, ZN => n21366);
   U1149 : NOR2_X1 port map( A1 => n21267, A2 => n31965, ZN => n28922);
   U8230 : NOR2_X1 port map( A1 => n12756, A2 => n810, ZN => n12017);
   U4734 : OAI21_X1 port map( A1 => n21138, A2 => n1553, B => n9699, ZN => 
                           n28754);
   U1254 : INV_X2 port map( I => n26622, ZN => n21755);
   U9651 : INV_X1 port map( I => n26494, ZN => n21153);
   U4675 : CLKBUF_X2 port map( I => n13442, Z => n26163);
   U14975 : CLKBUF_X2 port map( I => n21849, Z => n13490);
   U5827 : CLKBUF_X2 port map( I => n21573, Z => n29552);
   U4166 : CLKBUF_X2 port map( I => n15863, Z => n3821);
   U4171 : BUF_X2 port map( I => n12866, Z => n15655);
   U998 : NAND2_X1 port map( A1 => n5383, A2 => n5494, ZN => n12391);
   U22461 : NAND2_X1 port map( A1 => n7182, A2 => n196, ZN => n5850);
   U9582 : INV_X2 port map( I => n4097, ZN => n16165);
   U5552 : INV_X1 port map( I => n4356, ZN => n21560);
   U18339 : NAND2_X1 port map( A1 => n30978, A2 => n11301, ZN => n3680);
   U14323 : NOR2_X1 port map( A1 => n7476, A2 => n21854, ZN => n27065);
   U21579 : BUF_X2 port map( I => n6442, Z => n31102);
   U15941 : INV_X1 port map( I => n21749, ZN => n1532);
   U8120 : OAI22_X1 port map( A1 => n16723, A2 => n1134, B1 => n21283, B2 => 
                           n1312, ZN => n16722);
   U18390 : NAND2_X1 port map( A1 => n21839, A2 => n21685, ZN => n30616);
   U21177 : NAND2_X1 port map( A1 => n21591, A2 => n3756, ZN => n15846);
   U11964 : INV_X1 port map( I => n21717, ZN => n26732);
   U21734 : NAND2_X1 port map( A1 => n21247, A2 => n31121, ZN => n27753);
   U3892 : CLKBUF_X4 port map( I => n9129, Z => n343);
   U14540 : INV_X1 port map( I => n12789, ZN => n13146);
   U5716 : INV_X2 port map( I => n32753, ZN => n29951);
   U4547 : CLKBUF_X2 port map( I => n17151, Z => n27415);
   U9436 : INV_X2 port map( I => n16627, ZN => n22434);
   U16980 : CLKBUF_X1 port map( I => n10183, Z => n30405);
   U2967 : INV_X2 port map( I => n22926, ZN => n22657);
   U762 : BUF_X2 port map( I => n29287, Z => n16334);
   U3173 : INV_X2 port map( I => n4425, ZN => n12043);
   U4498 : NAND2_X1 port map( A1 => n33283, A2 => n994, ZN => n27495);
   U16505 : OAI21_X1 port map( A1 => n22434, A2 => n11895, B => n28473, ZN => 
                           n14329);
   U25077 : NOR2_X1 port map( A1 => n22550, A2 => n15260, ZN => n22392);
   U6298 : NAND3_X1 port map( A1 => n15322, A2 => n11895, A3 => n22435, ZN => 
                           n12688);
   U4527 : NAND3_X1 port map( A1 => n22200, A2 => n8519, A3 => n31636, ZN => 
                           n3384);
   U3565 : BUF_X4 port map( I => n15501, Z => n29070);
   U7168 : BUF_X2 port map( I => n28942, Z => n26251);
   U6955 : BUF_X2 port map( I => n6874, Z => n3657);
   U697 : BUF_X2 port map( I => n23065, Z => n4067);
   U6795 : BUF_X2 port map( I => n15123, Z => n28313);
   U20492 : CLKBUF_X1 port map( I => n31854, Z => n30925);
   U4065 : CLKBUF_X1 port map( I => n2449, Z => n30455);
   U5644 : BUF_X2 port map( I => n15324, Z => n26526);
   U6837 : OAI21_X1 port map( A1 => n23096, A2 => n22786, B => n18261, ZN => 
                           n3297);
   U2272 : CLKBUF_X1 port map( I => n4124, Z => n28849);
   U10961 : NOR2_X1 port map( A1 => n22781, A2 => n29173, ZN => n11741);
   U2990 : AOI21_X1 port map( A1 => n28348, A2 => n28349, B => n22720, ZN => 
                           n5345);
   U14187 : NAND2_X1 port map( A1 => n13004, A2 => n28853, ZN => n13003);
   U24011 : BUF_X1 port map( I => n27175, Z => n23238);
   U16177 : BUF_X2 port map( I => n23171, Z => n27243);
   U584 : CLKBUF_X4 port map( I => n23916, Z => n23721);
   U3223 : BUF_X2 port map( I => n29270, Z => n354);
   U6217 : INV_X1 port map( I => n29271, ZN => n895);
   U4470 : CLKBUF_X2 port map( I => n14031, Z => n28273);
   U6880 : OAI21_X1 port map( A1 => n11821, A2 => n8408, B => n10142, ZN => 
                           n13224);
   U410 : BUF_X2 port map( I => n17872, Z => n6392);
   U332 : OAI21_X1 port map( A1 => n31071, A2 => n13600, B => n32520, ZN => 
                           n31872);
   U13696 : CLKBUF_X1 port map( I => n24096, Z => n30146);
   U9539 : OR2_X1 port map( A1 => n24177, A2 => n15720, Z => n14052);
   U5520 : NAND2_X1 port map( A1 => n1092, A2 => n31342, ZN => n31341);
   U25164 : AOI21_X1 port map( A1 => n15537, A2 => n15899, B => n28726, ZN => 
                           n28725);
   U5465 : NAND2_X1 port map( A1 => n31341, A2 => n29949, ZN => n28522);
   U2526 : CLKBUF_X2 port map( I => n9353, Z => n30358);
   U15900 : AND2_X1 port map( A1 => n25628, A2 => n17523, Z => n12926);
   U9006 : OR2_X1 port map( A1 => n17641, A2 => n34169, Z => n25566);
   U2960 : CLKBUF_X1 port map( I => n25277, Z => n298);
   U13184 : AOI21_X1 port map( A1 => n1205, A2 => n42, B => n2264, ZN => n2263)
                           ;
   U8145 : NOR2_X1 port map( A1 => n18034, A2 => n28923, ZN => n18033);
   U5395 : INV_X2 port map( I => n20227, ZN => n3972);
   U20867 : INV_X2 port map( I => n4119, ZN => n21200);
   U6301 : INV_X2 port map( I => n19779, ZN => n19434);
   U105 : NOR2_X2 port map( A1 => n24725, A2 => n12699, ZN => n12651);
   U11678 : OAI21_X2 port map( A1 => n4468, A2 => n8998, B => n12516, ZN => 
                           n12515);
   U6471 : INV_X2 port map( I => n20385, ZN => n12514);
   U15300 : BUF_X4 port map( I => n24823, Z => n4240);
   U5953 : BUF_X4 port map( I => n17820, Z => n3388);
   U15203 : INV_X4 port map( I => n5889, ZN => n19063);
   U8492 : INV_X4 port map( I => n20384, ZN => n8998);
   U634 : AOI21_X2 port map( A1 => n21374, A2 => n4145, B => n32452, ZN => 
                           n21141);
   U641 : AOI22_X2 port map( A1 => n27410, A2 => n27409, B1 => n17212, B2 => 
                           n29635, ZN => n7584);
   U9905 : OAI21_X2 port map( A1 => n939, A2 => n16489, B => n4938, ZN => 
                           n19438);
   U2684 : BUF_X4 port map( I => n25973, Z => n25974);
   U16038 : BUF_X4 port map( I => n15212, Z => n31263);
   U3098 : AOI21_X2 port map( A1 => n24317, A2 => n14112, B => n2913, ZN => 
                           n9892);
   U6590 : NOR2_X2 port map( A1 => n19259, A2 => n28379, ZN => n6342);
   U594 : BUF_X4 port map( I => n17929, Z => n26582);
   U3414 : NAND3_X2 port map( A1 => n31381, A2 => n25821, A3 => n18246, ZN => 
                           n8345);
   U21542 : NOR2_X2 port map( A1 => n3183, A2 => n31824, ZN => n22740);
   U19079 : NAND2_X1 port map( A1 => n17578, A2 => n23874, ZN => n23875);
   U17316 : NAND3_X2 port map( A1 => n2128, A2 => n3006, A3 => n1934, ZN => 
                           n30837);
   U3866 : INV_X4 port map( I => n31824, ZN => n29173);
   U21587 : OAI21_X2 port map( A1 => n831, A2 => n27262, B => n25607, ZN => 
                           n25600);
   U6619 : NOR2_X1 port map( A1 => n4494, A2 => n27539, ZN => n26152);
   U8607 : INV_X4 port map( I => n19926, ZN => n20149);
   U16275 : OAI21_X2 port map( A1 => n24152, A2 => n24154, B => n27259, ZN => 
                           n24066);
   U8432 : NOR2_X2 port map( A1 => n29583, A2 => n6216, ZN => n30122);
   U4158 : NOR2_X1 port map( A1 => n300, A2 => n13263, ZN => n13262);
   U5519 : INV_X2 port map( I => n29087, ZN => n18571);
   U17233 : INV_X1 port map( I => n27428, ZN => n12006);
   U6147 : NOR2_X1 port map( A1 => n18639, A2 => n18815, ZN => n18383);
   U21163 : NAND2_X1 port map( A1 => n18633, A2 => n18710, ZN => n16295);
   U10456 : INV_X1 port map( I => n29776, ZN => n27958);
   U22552 : INV_X1 port map( I => n28321, ZN => n14926);
   U8805 : INV_X2 port map( I => n18737, ZN => n17360);
   U984 : INV_X1 port map( I => n18862, ZN => n18738);
   U26412 : NOR2_X1 port map( A1 => n15811, A2 => n27142, ZN => n31748);
   U3453 : CLKBUF_X2 port map( I => n495, Z => n46);
   U1639 : BUF_X2 port map( I => n18874, Z => n16538);
   U987 : NOR2_X1 port map( A1 => n1659, A2 => n5700, ZN => n18400);
   U7471 : INV_X1 port map( I => n26249, ZN => n18018);
   U5185 : INV_X1 port map( I => n962, ZN => n6891);
   U5120 : INV_X1 port map( I => n18586, ZN => n17166);
   U6722 : INV_X1 port map( I => n13719, ZN => n8739);
   U7649 : BUF_X2 port map( I => n10664, Z => n5269);
   U6703 : INV_X1 port map( I => n18756, ZN => n18602);
   U7650 : INV_X1 port map( I => n18580, ZN => n17419);
   U6711 : INV_X2 port map( I => n18722, ZN => n18727);
   U12190 : OR2_X1 port map( A1 => n490, A2 => n18723, Z => n18584);
   U975 : NOR2_X1 port map( A1 => n29182, A2 => n18727, ZN => n11164);
   U6701 : INV_X1 port map( I => n7216, ZN => n1853);
   U6668 : INV_X2 port map( I => n15873, ZN => n1059);
   U24350 : NOR2_X1 port map( A1 => n28675, A2 => n18687, ZN => n18691);
   U1009 : INV_X1 port map( I => n15519, ZN => n959);
   U20742 : NOR2_X1 port map( A1 => n18559, A2 => n18623, ZN => n18328);
   U7624 : NAND2_X1 port map( A1 => n882, A2 => n11097, ZN => n12876);
   U23918 : NOR2_X1 port map( A1 => n882, A2 => n30472, ZN => n17422);
   U15509 : NOR2_X1 port map( A1 => n3954, A2 => n8386, ZN => n18653);
   U22518 : NOR2_X1 port map( A1 => n18815, A2 => n13663, ZN => n18816);
   U8806 : INV_X2 port map( I => n15902, ZN => n18875);
   U10184 : NAND2_X1 port map( A1 => n18710, A2 => n18711, ZN => n11270);
   U10751 : NOR2_X1 port map( A1 => n15888, A2 => n32337, ZN => n17190);
   U12165 : NAND2_X1 port map( A1 => n16393, A2 => n13663, ZN => n8735);
   U10165 : INV_X1 port map( I => n15211, ZN => n18856);
   U5522 : INV_X2 port map( I => n18743, ZN => n16358);
   U24363 : NAND2_X1 port map( A1 => n18288, A2 => n27940, ZN => n18760);
   U7616 : INV_X2 port map( I => n18774, ZN => n18556);
   U10208 : INV_X1 port map( I => n16249, ZN => n1186);
   U8823 : NAND2_X1 port map( A1 => n18849, A2 => n18845, ZN => n6312);
   U5967 : NOR2_X1 port map( A1 => n5834, A2 => n18681, ZN => n4926);
   U14717 : INV_X1 port map( I => n16915, ZN => n6256);
   U4901 : INV_X1 port map( I => n490, ZN => n11123);
   U1608 : INV_X1 port map( I => n488, ZN => n1185);
   U1822 : NOR2_X1 port map( A1 => n14651, A2 => n18638, ZN => n14344);
   U12151 : INV_X1 port map( I => n9667, ZN => n3018);
   U16367 : AND2_X1 port map( A1 => n15966, A2 => n17030, Z => n18733);
   U2830 : INV_X1 port map( I => n13445, ZN => n18511);
   U16157 : INV_X1 port map( I => n18581, ZN => n18726);
   U3389 : INV_X1 port map( I => n18487, ZN => n18829);
   U2809 : OR2_X1 port map( A1 => n15216, A2 => n15347, Z => n18579);
   U7551 : NAND2_X1 port map( A1 => n18288, A2 => n33472, ZN => n18603);
   U5029 : NOR3_X1 port map( A1 => n18881, A2 => n18880, A3 => n16588, ZN => 
                           n10637);
   U2836 : NAND2_X1 port map( A1 => n180, A2 => n18493, ZN => n18326);
   U8773 : NAND2_X1 port map( A1 => n5269, A2 => n18746, ZN => n14705);
   U6156 : INV_X1 port map( I => n18579, ZN => n6873);
   U15658 : NAND2_X1 port map( A1 => n4259, A2 => n31579, ZN => n18277);
   U20416 : NAND2_X1 port map( A1 => n11164, A2 => n12320, ZN => n11023);
   U14039 : NAND2_X1 port map( A1 => n951, A2 => n8570, ZN => n5646);
   U12608 : NOR2_X1 port map( A1 => n15902, A2 => n10181, ZN => n1710);
   U26256 : NOR2_X1 port map( A1 => n16393, A2 => n18815, ZN => n6393);
   U1622 : INV_X1 port map( I => n28438, ZN => n18578);
   U2006 : INV_X1 port map( I => n18604, ZN => n30181);
   U19820 : NOR2_X1 port map( A1 => n10964, A2 => n12120, ZN => n15136);
   U7438 : NOR2_X1 port map( A1 => n31972, A2 => n28675, ZN => n13860);
   U14734 : NAND2_X1 port map( A1 => n1059, A2 => n9651, ZN => n30255);
   U7645 : INV_X2 port map( I => n16474, ZN => n17465);
   U4891 : NOR2_X1 port map( A1 => n13014, A2 => n13013, ZN => n18921);
   U8781 : INV_X1 port map( I => n18880, ZN => n18112);
   U10168 : NOR2_X1 port map( A1 => n16564, A2 => n18770, ZN => n18495);
   U3167 : NAND2_X1 port map( A1 => n18617, A2 => n16948, ZN => n2042);
   U4650 : INV_X1 port map( I => n26040, ZN => n732);
   U24291 : INV_X1 port map( I => n18563, ZN => n18464);
   U12401 : AND2_X1 port map( A1 => n18874, A2 => n27311, Z => n14658);
   U8813 : INV_X1 port map( I => n34139, ZN => n18566);
   U23513 : OAI21_X1 port map( A1 => n18880, A2 => n16572, B => n16588, ZN => 
                           n16109);
   U22172 : NOR2_X1 port map( A1 => n31972, A2 => n10283, ZN => n18399);
   U6168 : AOI22_X1 port map( A1 => n18543, A2 => n18854, B1 => n18307, B2 => 
                           n18853, ZN => n18308);
   U5971 : NOR2_X1 port map( A1 => n2042, A2 => n17224, ZN => n6298);
   U21153 : OAI21_X1 port map( A1 => n18553, A2 => n15694, B => n28548, ZN => 
                           n15693);
   U992 : OAI22_X1 port map( A1 => n3436, A2 => n1853, B1 => n3437, B2 => n956,
                           ZN => n17131);
   U20188 : AOI21_X1 port map( A1 => n31724, A2 => n6119, B => n17843, ZN => 
                           n18447);
   U950 : NOR2_X1 port map( A1 => n13548, A2 => n26810, ZN => n10125);
   U6191 : NOR2_X1 port map( A1 => n18496, A2 => n10043, ZN => n6666);
   U18796 : NOR2_X1 port map( A1 => n18880, A2 => n16466, ZN => n15984);
   U1617 : INV_X1 port map( I => n6138, ZN => n26680);
   U1596 : NAND2_X1 port map( A1 => n11097, A2 => n14213, ZN => n26320);
   U24225 : NAND2_X1 port map( A1 => n7454, A2 => n13514, ZN => n18362);
   U2049 : NOR2_X1 port map( A1 => n18643, A2 => n16766, ZN => n31369);
   U20825 : NAND2_X1 port map( A1 => n18817, A2 => n18714, ZN => n16088);
   U24326 : NOR2_X1 port map( A1 => n18584, A2 => n29602, ZN => n18585);
   U12130 : NAND2_X1 port map( A1 => n10565, A2 => n18574, ZN => n10564);
   U10120 : AOI22_X1 port map( A1 => n6393, A2 => n829, B1 => n18515, B2 => 
                           n7977, ZN => n4114);
   U20817 : NOR3_X1 port map( A1 => n13566, A2 => n18633, A3 => n1439, ZN => 
                           n13565);
   U14729 : NAND2_X1 port map( A1 => n16867, A2 => n30255, ZN => n11470);
   U24307 : NAND2_X1 port map( A1 => n33783, A2 => n18633, ZN => n18508);
   U6208 : AOI22_X1 port map( A1 => n10095, A2 => n18812, B1 => n18893, B2 => 
                           n27228, ZN => n27618);
   U3460 : INV_X2 port map( I => n29223, ZN => n1046);
   U10132 : NAND3_X1 port map( A1 => n18516, A2 => n1572, A3 => n33548, ZN => 
                           n14660);
   U2007 : INV_X1 port map( I => n18939, ZN => n30958);
   U4241 : BUF_X2 port map( I => n16748, Z => n13390);
   U2535 : INV_X2 port map( I => n16047, ZN => n19088);
   U5495 : INV_X1 port map( I => n13673, ZN => n19120);
   U24384 : INV_X1 port map( I => n19006, ZN => n18876);
   U4603 : INV_X1 port map( I => n19325, ZN => n19105);
   U6184 : NAND2_X1 port map( A1 => n19267, A2 => n19265, ZN => n19225);
   U12364 : NAND2_X1 port map( A1 => n11477, A2 => n10714, ZN => n19183);
   U1986 : INV_X1 port map( I => n8800, ZN => n31152);
   U6233 : NAND2_X1 port map( A1 => n5760, A2 => n18988, ZN => n5761);
   U8685 : INV_X1 port map( I => n19089, ZN => n6510);
   U21808 : INV_X1 port map( I => n19115, ZN => n13329);
   U1147 : BUF_X2 port map( I => n14198, Z => n6516);
   U934 : INV_X2 port map( I => n29757, ZN => n1180);
   U5009 : INV_X2 port map( I => n19285, ZN => n19078);
   U5498 : INV_X2 port map( I => n10974, ZN => n10203);
   U5479 : INV_X1 port map( I => n19199, ZN => n19093);
   U15405 : INV_X1 port map( I => n19049, ZN => n949);
   U3967 : INV_X1 port map( I => n19167, ZN => n824);
   U14584 : INV_X1 port map( I => n10714, ZN => n1049);
   U5955 : INV_X1 port map( I => n2692, ZN => n2901);
   U21867 : INV_X1 port map( I => n28197, ZN => n15239);
   U3180 : INV_X1 port map( I => n19104, ZN => n944);
   U14351 : INV_X1 port map( I => n8379, ZN => n1054);
   U920 : INV_X1 port map( I => n8141, ZN => n17386);
   U8697 : INV_X1 port map( I => n19265, ZN => n2101);
   U1938 : INV_X2 port map( I => n29769, ZN => n19179);
   U15846 : NAND2_X1 port map( A1 => n25968, A2 => n8787, ZN => n19114);
   U12085 : INV_X1 port map( I => n19274, ZN => n19321);
   U10014 : NAND2_X1 port map( A1 => n19248, A2 => n1050, ZN => n5082);
   U6229 : NAND2_X1 port map( A1 => n949, A2 => n19048, ZN => n12708);
   U21162 : OAI21_X1 port map( A1 => n27743, A2 => n29525, B => n12500, ZN => 
                           n12831);
   U6620 : NAND2_X1 port map( A1 => n19158, A2 => n14811, ZN => n19112);
   U21465 : NOR2_X1 port map( A1 => n19357, A2 => n14624, ZN => n16749);
   U8681 : NOR2_X1 port map( A1 => n13390, A2 => n19228, ZN => n18068);
   U1950 : NAND2_X1 port map( A1 => n26891, A2 => n10700, ZN => n13226);
   U2999 : INV_X1 port map( I => n19101, ZN => n19009);
   U9339 : NOR2_X1 port map( A1 => n880, A2 => n950, ZN => n2039);
   U22149 : OR2_X1 port map( A1 => n4747, A2 => n30879, Z => n5653);
   U7485 : NOR2_X1 port map( A1 => n17445, A2 => n7995, ZN => n11714);
   U12017 : INV_X1 port map( I => n19100, ZN => n11715);
   U20393 : OAI21_X1 port map( A1 => n26830, A2 => n6516, B => n19228, ZN => 
                           n16768);
   U21360 : CLKBUF_X2 port map( I => n26969, Z => n31074);
   U25977 : BUF_X2 port map( I => n19104, Z => n28935);
   U21560 : NAND2_X1 port map( A1 => n1380, A2 => n19222, ZN => n12468);
   U5238 : NAND2_X1 port map( A1 => n19318, A2 => n19319, ZN => n19317);
   U17411 : NAND3_X1 port map( A1 => n19040, A2 => n19049, A3 => n19042, ZN => 
                           n18135);
   U4999 : INV_X1 port map( I => n1807, ZN => n5656);
   U7475 : INV_X2 port map( I => n2935, ZN => n1766);
   U8673 : INV_X2 port map( I => n19301, ZN => n19291);
   U26347 : INV_X2 port map( I => n19180, ZN => n784);
   U21453 : NOR2_X1 port map( A1 => n18997, A2 => n18996, ZN => n12937);
   U1502 : CLKBUF_X2 port map( I => n8024, Z => n27818);
   U12308 : INV_X2 port map( I => n5491, ZN => n17370);
   U3709 : NAND2_X1 port map( A1 => n29047, A2 => n26417, ZN => n5877);
   U8708 : NOR2_X1 port map( A1 => n11940, A2 => n8379, ZN => n1764);
   U24129 : INV_X1 port map( I => n19212, ZN => n1373);
   U5940 : INV_X1 port map( I => n2799, ZN => n3207);
   U21428 : INV_X1 port map( I => n19178, ZN => n18957);
   U6202 : INV_X1 port map( I => n19156, ZN => n27587);
   U8712 : INV_X1 port map( I => n15411, ZN => n8742);
   U8017 : NAND2_X1 port map( A1 => n31726, A2 => n19265, ZN => n28447);
   U4619 : INV_X1 port map( I => n7197, ZN => n19152);
   U8627 : INV_X1 port map( I => n8024, ZN => n19242);
   U1521 : INV_X2 port map( I => n11203, ZN => n827);
   U8252 : OR2_X1 port map( A1 => n30879, A2 => n31746, Z => n19148);
   U8747 : NAND2_X1 port map( A1 => n19267, A2 => n19268, ZN => n19270);
   U16817 : AOI21_X1 port map( A1 => n19113, A2 => n19112, B => n27587, ZN => 
                           n27353);
   U1804 : CLKBUF_X2 port map( I => n19220, Z => n4);
   U3553 : NAND2_X1 port map( A1 => n1052, A2 => n26600, ZN => n4658);
   U26139 : OAI21_X1 port map( A1 => n19112, A2 => n12549, B => n19113, ZN => 
                           n26250);
   U21716 : NAND2_X1 port map( A1 => n19179, A2 => n18957, ZN => n11955);
   U1469 : AOI21_X1 port map( A1 => n19103, A2 => n19100, B => n17445, ZN => 
                           n27076);
   U4019 : NOR2_X1 port map( A1 => n4066, A2 => n19158, ZN => n18970);
   U1922 : NAND2_X1 port map( A1 => n4835, A2 => n30817, ZN => n18967);
   U10718 : NAND2_X1 port map( A1 => n19032, A2 => n10203, ZN => n18788);
   U5183 : NAND3_X1 port map( A1 => n19060, A2 => n9787, A3 => n1179, ZN => 
                           n2410);
   U12451 : NOR2_X1 port map( A1 => n19101, A2 => n11744, ZN => n18952);
   U12009 : INV_X1 port map( I => n19085, ZN => n18926);
   U7454 : NOR2_X1 port map( A1 => n6343, A2 => n6342, ZN => n9238);
   U7463 : NAND3_X1 port map( A1 => n12468, A2 => n12505, A3 => n1378, ZN => 
                           n12504);
   U7497 : INV_X1 port map( I => n9885, ZN => n12815);
   U8338 : INV_X1 port map( I => n13219, ZN => n26355);
   U9980 : AOI21_X1 port map( A1 => n19217, A2 => n29, B => n827, ZN => n6578);
   U5005 : INV_X1 port map( I => n18958, ZN => n4749);
   U8641 : NAND3_X1 port map( A1 => n14148, A2 => n19088, A3 => n12807, ZN => 
                           n18991);
   U5933 : NOR2_X1 port map( A1 => n14233, A2 => n11203, ZN => n18999);
   U15432 : OAI22_X1 port map( A1 => n19090, A2 => n1047, B1 => n19091, B2 => 
                           n5760, ZN => n17556);
   U8878 : OAI21_X1 port map( A1 => n16768, A2 => n16769, B => n18440, ZN => 
                           n17997);
   U9984 : NAND2_X1 port map( A1 => n9078, A2 => n2970, ZN => n8828);
   U22767 : NAND2_X1 port map( A1 => n8233, A2 => n19124, ZN => n18955);
   U7472 : INV_X1 port map( I => n31658, ZN => n15910);
   U8706 : INV_X1 port map( I => n18974, ZN => n1048);
   U938 : NAND2_X1 port map( A1 => n7134, A2 => n743, ZN => n19039);
   U5199 : NAND2_X1 port map( A1 => n947, A2 => n14312, ZN => n6446);
   U6587 : NAND2_X1 port map( A1 => n950, A2 => n7732, ZN => n15396);
   U3340 : NAND2_X1 port map( A1 => n1378, A2 => n16185, ZN => n379);
   U5487 : INV_X1 port map( I => n19262, ZN => n19140);
   U4945 : NOR2_X1 port map( A1 => n5118, A2 => n7995, ZN => n18953);
   U901 : INV_X1 port map( I => n27743, ZN => n17238);
   U1944 : NAND2_X1 port map( A1 => n1630, A2 => n33608, ZN => n2703);
   U8644 : NAND2_X1 port map( A1 => n2177, A2 => n19143, ZN => n1631);
   U1507 : NOR2_X1 port map( A1 => n15534, A2 => n4747, ZN => n26553);
   U9994 : OAI22_X1 port map( A1 => n19133, A2 => n15050, B1 => n19132, B2 => 
                           n1050, ZN => n15126);
   U22684 : AOI21_X1 port map( A1 => n7557, A2 => n12502, B => n27941, ZN => 
                           n13449);
   U5467 : AOI22_X1 port map( A1 => n6142, A2 => n1054, B1 => n1373, B2 => 
                           n29963, ZN => n4191);
   U11316 : OAI21_X1 port map( A1 => n19179, A2 => n19181, B => n13200, ZN => 
                           n18917);
   U6272 : NOR2_X1 port map( A1 => n11000, A2 => n19315, ZN => n18230);
   U15640 : OAI21_X1 port map( A1 => n32451, A2 => n19036, B => n12850, ZN => 
                           n12849);
   U5214 : NOR2_X1 port map( A1 => n19038, A2 => n31139, ZN => n7749);
   U890 : NAND2_X1 port map( A1 => n29378, A2 => n827, ZN => n18938);
   U3160 : OAI22_X1 port map( A1 => n19154, A2 => n950, B1 => n8862, B2 => n879
                           , ZN => n13072);
   U10027 : NAND2_X1 port map( A1 => n16068, A2 => n7968, ZN => n17319);
   U2534 : NAND2_X1 port map( A1 => n19309, A2 => n14178, ZN => n2519);
   U26143 : AOI22_X1 port map( A1 => n4102, A2 => n26417, B1 => n30412, B2 => 
                           n19032, ZN => n29044);
   U5244 : NAND2_X1 port map( A1 => n15845, A2 => n19281, ZN => n15843);
   U21190 : OAI21_X1 port map( A1 => n15628, A2 => n32908, B => n28386, ZN => 
                           n15627);
   U8632 : OAI21_X1 port map( A1 => n7201, A2 => n7200, B => n33581, ZN => 
                           n7199);
   U18140 : OAI21_X1 port map( A1 => n19291, A2 => n29223, B => n13957, ZN => 
                           n18927);
   U21730 : NOR2_X1 port map( A1 => n11875, A2 => n28175, ZN => n14355);
   U8633 : NOR2_X1 port map( A1 => n14030, A2 => n5812, ZN => n4386);
   U7505 : NAND2_X1 port map( A1 => n19315, A2 => n31970, ZN => n19151);
   U8648 : INV_X1 port map( I => n1494, ZN => n1492);
   U12420 : NAND2_X1 port map( A1 => n18477, A2 => n14760, ZN => n18381);
   U1512 : NAND2_X1 port map( A1 => n1883, A2 => n16699, ZN => n12813);
   U24469 : NOR2_X1 port map( A1 => n827, A2 => n7557, ZN => n19349);
   U12144 : OAI21_X1 port map( A1 => n19260, A2 => n744, B => n16740, ZN => 
                           n16741);
   U8422 : NAND2_X1 port map( A1 => n19177, A2 => n19178, ZN => n29580);
   U21486 : OAI21_X1 port map( A1 => n1883, A2 => n12815, B => n12813, ZN => 
                           n18813);
   U21017 : OAI21_X1 port map( A1 => n17527, A2 => n31029, B => n26518, ZN => 
                           n11295);
   U1921 : NAND2_X1 port map( A1 => n10013, A2 => n2582, ZN => n19056);
   U1456 : NAND3_X1 port map( A1 => n9441, A2 => n9442, A3 => n1180, ZN => 
                           n16797);
   U5160 : INV_X1 port map( I => n19676, ZN => n1369);
   U10240 : BUF_X2 port map( I => Key(60), Z => n25598);
   U15524 : AOI22_X1 port map( A1 => n19139, A2 => n28379, B1 => n19140, B2 => 
                           n16876, ZN => n16875);
   U6288 : AOI21_X1 port map( A1 => n18982, A2 => n13685, B => n17508, ZN => 
                           n17507);
   U4983 : NAND2_X1 port map( A1 => n26289, A2 => n26288, ZN => n8897);
   U9970 : NOR2_X1 port map( A1 => n17528, A2 => n17526, ZN => n13355);
   U1451 : CLKBUF_X2 port map( I => n19710, Z => n25998);
   U13057 : NAND2_X1 port map( A1 => n2126, A2 => n2125, ZN => n16158);
   U3091 : INV_X1 port map( I => n19768, ZN => n1363);
   U24436 : INV_X1 port map( I => n19136, ZN => n19142);
   U9765 : INV_X1 port map( I => n9629, ZN => n1368);
   U18921 : INV_X1 port map( I => n13480, ZN => n7826);
   U1885 : INV_X1 port map( I => n31882, ZN => n31057);
   U4949 : NOR3_X1 port map( A1 => n1984, A2 => n5606, A3 => n5608, ZN => n5605
                           );
   U20879 : INV_X1 port map( I => n30411, ZN => n19498);
   U18294 : INV_X1 port map( I => n14094, ZN => n19566);
   U12519 : BUF_X2 port map( I => n14120, Z => n26794);
   U1891 : CLKBUF_X2 port map( I => n6387, Z => n30212);
   U6569 : INV_X1 port map( I => n14214, ZN => n19375);
   U2821 : INV_X1 port map( I => n13645, ZN => n19479);
   U5273 : INV_X1 port map( I => n19780, ZN => n30712);
   U6322 : INV_X1 port map( I => n19568, ZN => n2375);
   U6269 : INV_X1 port map( I => n12610, ZN => n29046);
   U22847 : BUF_X2 port map( I => n29130, Z => n31279);
   U877 : INV_X1 port map( I => n19378, ZN => n1173);
   U15123 : BUF_X2 port map( I => Key(20), Z => n16581);
   U3254 : OAI22_X1 port map( A1 => n7438, A2 => n12532, B1 => n7437, B2 => 
                           n7436, ZN => n27144);
   U1442 : INV_X1 port map( I => n25266, ZN => n26000);
   U2103 : CLKBUF_X2 port map( I => n16158, Z => n29890);
   U24031 : INV_X1 port map( I => n31414, ZN => n31908);
   U16319 : INV_X1 port map( I => n4883, ZN => n14766);
   U1881 : INV_X1 port map( I => n24487, ZN => n30993);
   U10319 : INV_X1 port map( I => n26551, ZN => n219);
   U11937 : INV_X1 port map( I => n15189, ZN => n2780);
   U6314 : INV_X1 port map( I => n11333, ZN => n1040);
   U8527 : INV_X2 port map( I => n8443, ZN => n6864);
   U13579 : INV_X1 port map( I => n568, ZN => n1043);
   U25215 : INV_X1 port map( I => n31538, ZN => n31906);
   U7417 : NAND2_X1 port map( A1 => n1043, A2 => n16694, ZN => n7923);
   U9946 : INV_X1 port map( I => n14576, ZN => n20119);
   U21561 : NOR2_X1 port map( A1 => n20099, A2 => n29216, ZN => n13978);
   U14087 : INV_X1 port map( I => n9469, ZN => n12045);
   U11876 : INV_X2 port map( I => n20113, ZN => n20044);
   U8517 : NAND2_X1 port map( A1 => n6611, A2 => n19991, ZN => n17136);
   U849 : INV_X2 port map( I => n18089, ZN => n8107);
   U2753 : BUF_X2 port map( I => n19857, Z => n28645);
   U12114 : NAND2_X1 port map( A1 => n8816, A2 => n29250, ZN => n19933);
   U2760 : INV_X2 port map( I => n19857, ZN => n20068);
   U13413 : INV_X1 port map( I => n2499, ZN => n20076);
   U862 : INV_X2 port map( I => n11913, ZN => n19986);
   U14698 : INV_X2 port map( I => n17575, ZN => n20056);
   U20330 : INV_X1 port map( I => n10863, ZN => n13327);
   U19734 : INV_X1 port map( I => n578, ZN => n1165);
   U7403 : INV_X1 port map( I => n31453, ZN => n20043);
   U1438 : INV_X1 port map( I => n1043, ZN => n28684);
   U19246 : INV_X2 port map( I => n8684, ZN => n17882);
   U2905 : BUF_X2 port map( I => n19885, Z => n224);
   U4606 : INV_X2 port map( I => n14761, ZN => n17260);
   U820 : INV_X1 port map( I => n19991, ZN => n11624);
   U1416 : OAI22_X1 port map( A1 => n11350, A2 => n28684, B1 => n7920, B2 => 
                           n1360, ZN => n18003);
   U5300 : NAND2_X1 port map( A1 => n19845, A2 => n16681, ZN => n1878);
   U11927 : NAND2_X1 port map( A1 => n29013, A2 => n502, ZN => n15736);
   U20999 : OAI21_X1 port map( A1 => n20136, A2 => n19834, B => n15174, ZN => 
                           n12634);
   U10277 : INV_X1 port map( I => n9201, ZN => n26547);
   U21536 : NOR2_X1 port map( A1 => n16092, A2 => n19966, ZN => n15258);
   U2685 : NAND2_X1 port map( A1 => n12682, A2 => n1169, ZN => n28012);
   U11036 : NAND2_X1 port map( A1 => n31468, A2 => n16154, ZN => n29853);
   U23549 : NAND2_X1 port map( A1 => n9876, A2 => n8301, ZN => n20081);
   U6408 : NOR2_X1 port map( A1 => n17260, A2 => n1699, ZN => n15247);
   U1832 : INV_X1 port map( I => n20124, ZN => n16155);
   U19845 : INV_X2 port map( I => n28704, ZN => n10340);
   U2866 : INV_X2 port map( I => n20056, ZN => n19883);
   U6375 : BUF_X2 port map( I => n8857, Z => n431);
   U836 : INV_X1 port map( I => n20155, ZN => n14747);
   U9951 : INV_X2 port map( I => n14457, ZN => n5707);
   U1776 : INV_X1 port map( I => n32745, ZN => n15551);
   U8562 : INV_X1 port map( I => n12045, ZN => n19856);
   U5286 : NAND2_X1 port map( A1 => n11521, A2 => n10947, ZN => n28218);
   U26411 : INV_X1 port map( I => n29250, ZN => n570);
   U3035 : OR2_X1 port map( A1 => n10059, A2 => n9690, Z => n19974);
   U22765 : INV_X2 port map( I => n20135, ZN => n15286);
   U4232 : INV_X1 port map( I => n32807, ZN => n19451);
   U5456 : INV_X1 port map( I => n11959, ZN => n8611);
   U1436 : INV_X1 port map( I => n16595, ZN => n20020);
   U1828 : INV_X2 port map( I => n27808, ZN => n4142);
   U11427 : NAND2_X1 port map( A1 => n16625, A2 => n29252, ZN => n11593);
   U26138 : BUF_X2 port map( I => n19936, Z => n29040);
   U9916 : INV_X2 port map( I => n15381, ZN => n14976);
   U7421 : INV_X2 port map( I => n31448, ZN => n20066);
   U2520 : NAND2_X1 port map( A1 => n19724, A2 => n567, ZN => n9031);
   U14899 : INV_X1 port map( I => n16298, ZN => n31694);
   U17922 : AOI21_X1 port map( A1 => n13327, A2 => n584, B => n16489, ZN => 
                           n14801);
   U1847 : NOR2_X1 port map( A1 => n6532, A2 => n10845, ZN => n19338);
   U10882 : OAI22_X1 port map( A1 => n2089, A2 => n3486, B1 => n19974, B2 => 
                           n15189, ZN => n27604);
   U1797 : NOR3_X1 port map( A1 => n19808, A2 => n16491, A3 => n15278, ZN => 
                           n11902);
   U24641 : OAI22_X1 port map( A1 => n20085, A2 => n20084, B1 => n16664, B2 => 
                           n9876, ZN => n20086);
   U17717 : AOI22_X1 port map( A1 => n940, A2 => n4233, B1 => n4215, B2 => 
                           n20157, ZN => n4230);
   U10752 : NOR2_X1 port map( A1 => n20061, A2 => n27832, ZN => n20062);
   U20890 : NOR2_X1 port map( A1 => n20068, A2 => n20067, ZN => n20069);
   U12490 : OAI22_X1 port map( A1 => n19926, A2 => n13591, B1 => n19614, B2 => 
                           n27097, ZN => n19623);
   U17450 : NAND3_X1 port map( A1 => n9033, A2 => n19806, A3 => n30375, ZN => 
                           n9032);
   U1364 : OAI21_X1 port map( A1 => n16966, A2 => n28600, B => n1699, ZN => 
                           n20104);
   U7368 : NAND2_X1 port map( A1 => n19951, A2 => n12045, ZN => n2845);
   U15514 : NAND2_X1 port map( A1 => n18003, A2 => n27624, ZN => n4167);
   U21123 : AOI22_X1 port map( A1 => n28852, A2 => n375, B1 => n15192, B2 => 
                           n19874, ZN => n31048);
   U1413 : NOR2_X1 port map( A1 => n27715, A2 => n28645, ZN => n17712);
   U19196 : NAND2_X1 port map( A1 => n33419, A2 => n20156, ZN => n8591);
   U20359 : OAI21_X1 port map( A1 => n17714, A2 => n17713, B => n19451, ZN => 
                           n10925);
   U24643 : NOR2_X1 port map( A1 => n14083, A2 => n20120, ZN => n20121);
   U8563 : NOR2_X1 port map( A1 => n12657, A2 => n149, ZN => n10768);
   U3898 : INV_X1 port map( I => n6027, ZN => n30845);
   U2122 : AOI21_X1 port map( A1 => n20056, A2 => n11958, B => n15665, ZN => 
                           n4637);
   U1350 : NOR2_X1 port map( A1 => n19824, A2 => n15306, ZN => n8431);
   U1843 : NAND2_X1 port map( A1 => n14644, A2 => n20000, ZN => n30790);
   U4518 : AND2_X1 port map( A1 => n11198, A2 => n31951, Z => n17156);
   U21986 : OAI21_X1 port map( A1 => n11521, A2 => n28219, B => n28218, ZN => 
                           n19843);
   U1390 : NOR2_X1 port map( A1 => n20099, A2 => n28087, ZN => n9855);
   U16569 : NAND2_X1 port map( A1 => n19969, A2 => n19970, ZN => n2908);
   U18847 : NOR2_X1 port map( A1 => n1164, A2 => n16694, ZN => n8295);
   U832 : INV_X1 port map( I => n16154, ZN => n19840);
   U12300 : OAI21_X1 port map( A1 => n783, A2 => n20147, B => n4602, ZN => 
                           n4443);
   U23500 : NAND2_X1 port map( A1 => n27597, A2 => n11961, ZN => n17365);
   U1395 : NOR2_X1 port map( A1 => n2694, A2 => n19995, ZN => n26238);
   U5156 : INV_X1 port map( I => n3989, ZN => n14927);
   U10981 : INV_X1 port map( I => n1358, ZN => n29845);
   U26176 : NAND2_X1 port map( A1 => n28208, A2 => n28209, ZN => n5549);
   U1787 : AOI21_X1 port map( A1 => n20081, A2 => n13585, B => n32780, ZN => 
                           n20087);
   U8531 : AOI22_X1 port map( A1 => n9450, A2 => n33743, B1 => n16155, B2 => 
                           n20120, ZN => n9449);
   U14741 : INV_X1 port map( I => n11872, ZN => n27318);
   U6527 : NAND2_X1 port map( A1 => n4233, A2 => n20043, ZN => n13611);
   U20260 : NOR2_X1 port map( A1 => n29208, A2 => n17389, ZN => n10695);
   U20064 : NOR2_X1 port map( A1 => n10272, A2 => n16694, ZN => n10271);
   U5889 : NOR2_X1 port map( A1 => n12337, A2 => n14210, ZN => n20144);
   U6554 : INV_X1 port map( I => n17882, ZN => n19943);
   U2712 : NOR2_X1 port map( A1 => n31993, A2 => n8216, ZN => n14134);
   U15109 : NOR2_X1 port map( A1 => n1362, A2 => n18142, ZN => n18141);
   U21472 : NAND2_X1 port map( A1 => n14334, A2 => n16595, ZN => n20125);
   U19704 : AND2_X1 port map( A1 => n6275, A2 => n8933, Z => n4855);
   U21034 : INV_X1 port map( I => n20076, ZN => n16059);
   U25903 : NAND2_X1 port map( A1 => n149, A2 => n29040, ZN => n28880);
   U7413 : INV_X1 port map( I => n822, ZN => n1438);
   U5288 : NOR2_X1 port map( A1 => n4215, A2 => n940, ZN => n10556);
   U22551 : INV_X1 port map( I => n33714, ZN => n5598);
   U6519 : AOI21_X1 port map( A1 => n20144, A2 => n20143, B => n12851, ZN => 
                           n2495);
   U8265 : NOR3_X1 port map( A1 => n16059, A2 => n12379, A3 => n6444, ZN => 
                           n12832);
   U26088 : OAI21_X1 port map( A1 => n31697, A2 => n29284, B => n31715, ZN => 
                           n31676);
   U24393 : OAI21_X1 port map( A1 => n20036, A2 => n8775, B => n29187, ZN => 
                           n28622);
   U21275 : OAI21_X1 port map( A1 => n19932, A2 => n31103, B => n579, ZN => 
                           n14799);
   U9887 : AOI22_X1 port map( A1 => n10465, A2 => n20077, B1 => n20079, B2 => 
                           n20078, ZN => n12598);
   U15158 : OAI21_X1 port map( A1 => n4972, A2 => n7014, B => n19853, ZN => 
                           n13283);
   U17724 : NAND3_X1 port map( A1 => n6611, A2 => n28876, A3 => n30366, ZN => 
                           n15850);
   U6401 : NAND2_X1 port map( A1 => n19878, A2 => n20096, ZN => n8183);
   U6522 : NAND3_X1 port map( A1 => n13583, A2 => n6960, A3 => n12168, ZN => 
                           n4498);
   U1740 : NAND2_X1 port map( A1 => n20065, A2 => n2606, ZN => n30922);
   U11814 : OAI22_X1 port map( A1 => n12696, A2 => n821, B1 => n20059, B2 => 
                           n19886, ZN => n2146);
   U1351 : NAND2_X1 port map( A1 => n3366, A2 => n13585, ZN => n13772);
   U12313 : NOR2_X1 port map( A1 => n1458, A2 => n14210, ZN => n2549);
   U17681 : OAI21_X1 port map( A1 => n2933, A2 => n9875, B => n1167, ZN => 
                           n27517);
   U1377 : NAND2_X1 port map( A1 => n10340, A2 => n17670, ZN => n28912);
   U22852 : NAND2_X1 port map( A1 => n31280, A2 => n15381, ZN => n13397);
   U1837 : NAND2_X1 port map( A1 => n19438, A2 => n1358, ZN => n11);
   U3893 : NAND3_X1 port map( A1 => n8783, A2 => n8782, A3 => n17967, ZN => 
                           n20190);
   U1335 : OAI21_X1 port map( A1 => n32000, A2 => n14622, B => n29656, ZN => 
                           n13955);
   U6377 : NAND2_X1 port map( A1 => n20063, A2 => n20062, ZN => n15310);
   U6392 : NAND3_X1 port map( A1 => n27829, A2 => n27830, A3 => n20135, ZN => 
                           n31585);
   U2259 : NAND2_X1 port map( A1 => n18949, A2 => n7609, ZN => n15436);
   U5140 : OAI21_X1 port map( A1 => n2534, A2 => n8443, B => n6200, ZN => 
                           n16951);
   U3360 : NAND2_X1 port map( A1 => n2845, A2 => n31080, ZN => n13284);
   U16560 : NAND2_X1 port map( A1 => n20026, A2 => n6109, ZN => n30356);
   U21215 : NOR2_X1 port map( A1 => n19867, A2 => n19868, ZN => n12987);
   U6420 : OAI21_X1 port map( A1 => n13157, A2 => n783, B => n330, ZN => n19832
                           );
   U1365 : OAI22_X1 port map( A1 => n3593, A2 => n20053, B1 => n11893, B2 => 
                           n15665, ZN => n3592);
   U1726 : INV_X2 port map( I => n20560, ZN => n20562);
   U12098 : INV_X2 port map( I => n20632, ZN => n15162);
   U24889 : NAND2_X1 port map( A1 => n3940, A2 => n3941, ZN => n28696);
   U5429 : BUF_X2 port map( I => n14720, Z => n11086);
   U6486 : INV_X2 port map( I => n31969, ZN => n20360);
   U18405 : INV_X1 port map( I => n20404, ZN => n2237);
   U4204 : INV_X1 port map( I => n20339, ZN => n20590);
   U20929 : NAND2_X1 port map( A1 => n20430, A2 => n20590, ZN => n16133);
   U2897 : NAND2_X1 port map( A1 => n20158, A2 => n30130, ZN => n10614);
   U9605 : INV_X2 port map( I => n16606, ZN => n20563);
   U15862 : INV_X1 port map( I => n29763, ZN => n20524);
   U3203 : NOR2_X1 port map( A1 => n11086, A2 => n12966, ZN => n20263);
   U12462 : INV_X2 port map( I => n10847, ZN => n10849);
   U23084 : NOR2_X1 port map( A1 => n20371, A2 => n15027, ZN => n20205);
   U1280 : NAND2_X1 port map( A1 => n5471, A2 => n20374, ZN => n1774);
   U2166 : INV_X2 port map( I => n2821, ZN => n14731);
   U20413 : INV_X1 port map( I => n15169, ZN => n20591);
   U9827 : INV_X2 port map( I => n20361, ZN => n1789);
   U1284 : NAND2_X1 port map( A1 => n1150, A2 => n20562, ZN => n27316);
   U7308 : INV_X1 port map( I => n2843, ZN => n16070);
   U21108 : NAND2_X1 port map( A1 => n19864, A2 => n20360, ZN => n13247);
   U7348 : CLKBUF_X2 port map( I => n20582, Z => n26232);
   U5103 : INV_X2 port map( I => n6679, ZN => n1032);
   U4927 : INV_X2 port map( I => n28261, ZN => n818);
   U7335 : INV_X1 port map( I => n9025, ZN => n935);
   U21603 : NAND2_X1 port map( A1 => n20602, A2 => n6996, ZN => n12184);
   U7736 : INV_X1 port map( I => n8870, ZN => n11312);
   U19661 : INV_X1 port map( I => n14187, ZN => n9484);
   U1256 : INV_X1 port map( I => n20329, ZN => n1149);
   U17294 : INV_X2 port map( I => n20615, ZN => n27741);
   U11626 : INV_X1 port map( I => n26881, ZN => n13537);
   U1265 : INV_X1 port map( I => n9831, ZN => n13538);
   U15861 : INV_X1 port map( I => n4460, ZN => n20358);
   U12773 : INV_X1 port map( I => n20467, ZN => n20160);
   U3119 : INV_X2 port map( I => n4254, ZN => n20487);
   U1294 : INV_X1 port map( I => n7218, ZN => n1034);
   U10575 : INV_X1 port map( I => n28390, ZN => n6475);
   U2899 : INV_X2 port map( I => n30130, ZN => n710);
   U3587 : AOI22_X1 port map( A1 => n29453, A2 => n31504, B1 => n20524, B2 => 
                           n33222, ZN => n8794);
   U17626 : INV_X2 port map( I => n32504, ZN => n30987);
   U4206 : INV_X1 port map( I => n935, ZN => n1030);
   U17975 : NAND2_X1 port map( A1 => n20450, A2 => n14179, ZN => n12227);
   U774 : BUF_X4 port map( I => n10847, Z => n10848);
   U2314 : NOR2_X1 port map( A1 => n20202, A2 => n20361, ZN => n120);
   U11738 : NOR2_X1 port map( A1 => n12169, A2 => n2879, ZN => n20235);
   U1705 : INV_X1 port map( I => n14436, ZN => n1151);
   U783 : INV_X1 port map( I => n33515, ZN => n1152);
   U9781 : INV_X1 port map( I => n20327, ZN => n11809);
   U7285 : INV_X1 port map( I => n3944, ZN => n17866);
   U11868 : NAND2_X1 port map( A1 => n1357, A2 => n20635, ZN => n20442);
   U21098 : NAND2_X1 port map( A1 => n16182, A2 => n15230, ZN => n3644);
   U4886 : BUF_X2 port map( I => n20374, Z => n27887);
   U7317 : INV_X1 port map( I => n17236, ZN => n4807);
   U24692 : NOR2_X1 port map( A1 => n20381, A2 => n30594, ZN => n20382);
   U6457 : INV_X1 port map( I => n16452, ZN => n20510);
   U1241 : NAND2_X1 port map( A1 => n20428, A2 => n20427, ZN => n4856);
   U13218 : NAND2_X1 port map( A1 => n8870, A2 => n31668, ZN => n26424);
   U7297 : BUF_X2 port map( I => n16606, Z => n13589);
   U22958 : NOR2_X1 port map( A1 => n1150, A2 => n20413, ZN => n14710);
   U4862 : INV_X1 port map( I => n15230, ZN => n20603);
   U4263 : NOR2_X1 port map( A1 => n1349, A2 => n20447, ZN => n30003);
   U6498 : NOR2_X1 port map( A1 => n28812, A2 => n14049, ZN => n20221);
   U3773 : INV_X1 port map( I => n12563, ZN => n9854);
   U1293 : INV_X1 port map( I => n30763, ZN => n28316);
   U3410 : INV_X1 port map( I => n27697, ZN => n20497);
   U8404 : INV_X2 port map( I => n20489, ZN => n20484);
   U16246 : INV_X2 port map( I => n31968, ZN => n11637);
   U2359 : INV_X1 port map( I => n11303, ZN => n12010);
   U743 : INV_X1 port map( I => n20401, ZN => n20571);
   U5440 : NOR2_X1 port map( A1 => n7577, A2 => n20395, ZN => n20462);
   U1698 : INV_X1 port map( I => n20471, ZN => n931);
   U13916 : NAND2_X1 port map( A1 => n20317, A2 => n32504, ZN => n2965);
   U5442 : INV_X1 port map( I => n20447, ZN => n781);
   U7391 : NAND2_X1 port map( A1 => n3944, A2 => n15282, ZN => n1465);
   U2555 : NAND2_X1 port map( A1 => n17866, A2 => n1355, ZN => n15713);
   U26568 : NAND2_X1 port map( A1 => n32033, A2 => n8031, ZN => n31834);
   U21395 : NAND2_X1 port map( A1 => n14369, A2 => n20507, ZN => n17652);
   U2126 : INV_X1 port map( I => n30931, ZN => n30413);
   U17304 : NOR2_X1 port map( A1 => n5275, A2 => n10106, ZN => n27442);
   U7275 : NOR2_X1 port map( A1 => n1150, A2 => n20562, ZN => n5952);
   U14016 : NAND2_X1 port map( A1 => n20194, A2 => n27755, ZN => n3065);
   U23052 : NAND3_X1 port map( A1 => n28357, A2 => n31009, A3 => n20489, ZN => 
                           n14945);
   U735 : NAND2_X1 port map( A1 => n20412, A2 => n818, ZN => n3137);
   U13789 : NOR2_X1 port map( A1 => n14054, A2 => n2843, ZN => n17043);
   U7246 : OAI22_X1 port map( A1 => n19830, A2 => n20427, B1 => n28376, B2 => 
                           n14731, ZN => n9725);
   U1633 : AOI21_X1 port map( A1 => n20536, A2 => n20537, B => n20541, ZN => 
                           n11447);
   U16846 : NAND2_X1 port map( A1 => n15045, A2 => n20563, ZN => n16217);
   U1564 : NAND2_X1 port map( A1 => n13353, A2 => n28288, ZN => n5416);
   U22977 : NOR2_X1 port map( A1 => n28527, A2 => n7873, ZN => n14768);
   U20838 : NAND2_X1 port map( A1 => n19930, A2 => n13589, ZN => n16216);
   U6296 : NAND2_X1 port map( A1 => n27697, A2 => n31804, ZN => n26089);
   U21531 : NAND2_X1 port map( A1 => n8998, A2 => n20630, ZN => n14566);
   U19868 : AOI21_X1 port map( A1 => n20538, A2 => n760, B => n4071, ZN => 
                           n11446);
   U4843 : NAND2_X1 port map( A1 => n20382, A2 => n111, ZN => n26987);
   U11728 : INV_X1 port map( I => n13253, ZN => n8942);
   U18289 : OAI21_X1 port map( A1 => n30603, A2 => n16123, B => n16452, ZN => 
                           n28752);
   U5382 : INV_X1 port map( I => n16144, ZN => n930);
   U11718 : NOR2_X1 port map( A1 => n13253, A2 => n28085, ZN => n9776);
   U13369 : NAND2_X1 port map( A1 => n20235, A2 => n33530, ZN => n16488);
   U10454 : BUF_X2 port map( I => n29814, Z => n29774);
   U15324 : INV_X1 port map( I => n5781, ZN => n20493);
   U11653 : NAND2_X1 port map( A1 => n16882, A2 => n9014, ZN => n9288);
   U11687 : NAND2_X1 port map( A1 => n8650, A2 => n2879, ZN => n15954);
   U7904 : NOR2_X1 port map( A1 => n29363, A2 => n29528, ZN => n29527);
   U19041 : INV_X1 port map( I => n20224, ZN => n11712);
   U1549 : NAND2_X1 port map( A1 => n10848, A2 => n1349, ZN => n10074);
   U17889 : NAND2_X1 port map( A1 => n30553, A2 => n32061, ZN => n31444);
   U1841 : NOR2_X1 port map( A1 => n1151, A2 => n26587, ZN => n7707);
   U4856 : NAND2_X1 port map( A1 => n1149, A2 => n13693, ZN => n13325);
   U15901 : NOR2_X1 port map( A1 => n31072, A2 => n31961, ZN => n20002);
   U7556 : INV_X1 port map( I => n13867, ZN => n26257);
   U15237 : INV_X1 port map( I => n11453, ZN => n27386);
   U21606 : AOI21_X1 port map( A1 => n14368, A2 => n3944, B => n14369, ZN => 
                           n14367);
   U9385 : NAND3_X1 port map( A1 => n10231, A2 => n20520, A3 => n16218, ZN => 
                           n29672);
   U24627 : OAI21_X1 port map( A1 => n28626, A2 => n26567, B => n20001, ZN => 
                           n20004);
   U20924 : AOI21_X1 port map( A1 => n20325, A2 => n932, B => n16174, ZN => 
                           n16492);
   U9776 : OAI21_X1 port map( A1 => n20405, A2 => n10848, B => n11616, ZN => 
                           n11618);
   U12998 : AOI22_X1 port map( A1 => n3428, A2 => n29623, B1 => n1157, B2 => 
                           n17043, ZN => n30079);
   U21394 : OAI22_X1 port map( A1 => n17652, A2 => n20510, B1 => n20508, B2 => 
                           n20509, ZN => n16774);
   U1231 : NAND3_X1 port map( A1 => n28357, A2 => n20487, A3 => n20486, ZN => 
                           n17513);
   U8379 : OAI21_X1 port map( A1 => n12771, A2 => n12169, B => n15954, ZN => 
                           n8960);
   U21604 : NAND3_X1 port map( A1 => n7116, A2 => n1160, A3 => n16182, ZN => 
                           n14965);
   U11380 : AOI22_X1 port map( A1 => n5950, A2 => n20562, B1 => n933, B2 => 
                           n16684, ZN => n5949);
   U9753 : NAND2_X1 port map( A1 => n13353, A2 => n30878, ZN => n7054);
   U23085 : NAND3_X1 port map( A1 => n20533, A2 => n1153, A3 => n15027, ZN => 
                           n20353);
   U9750 : NOR2_X1 port map( A1 => n20252, A2 => n20484, ZN => n7479);
   U17404 : NAND3_X1 port map( A1 => n14566, A2 => n20631, A3 => n111, ZN => 
                           n14565);
   U7622 : AOI21_X1 port map( A1 => n15045, A2 => n13589, B => n9776, ZN => 
                           n9775);
   U1527 : NAND3_X1 port map( A1 => n30545, A2 => n30987, A3 => n7394, ZN => 
                           n2770);
   U20928 : NOR2_X1 port map( A1 => n20378, A2 => n5471, ZN => n16139);
   U20836 : NAND3_X1 port map( A1 => n20341, A2 => n20340, A3 => n26756, ZN => 
                           n12846);
   U1556 : INV_X1 port map( I => n7397, ZN => n20220);
   U1205 : NAND2_X1 port map( A1 => n16787, A2 => n14177, ZN => n14176);
   U9759 : OR2_X1 port map( A1 => n20341, A2 => n1347, Z => n14263);
   U11645 : OAI21_X1 port map( A1 => n14571, A2 => n14005, B => n15173, ZN => 
                           n6311);
   U23490 : AOI21_X1 port map( A1 => n31338, A2 => n3904, B => n20238, ZN => 
                           n9587);
   U6481 : AOI21_X1 port map( A1 => n20358, A2 => n28625, B => n31891, ZN => 
                           n2320);
   U7268 : OAI21_X1 port map( A1 => n3751, A2 => n3750, B => n15217, ZN => 
                           n20612);
   U9796 : NAND2_X1 port map( A1 => n14051, A2 => n14050, ZN => n31269);
   U1544 : NAND2_X1 port map( A1 => n31422, A2 => n31210, ZN => n30856);
   U1565 : NAND3_X1 port map( A1 => n266, A2 => n20268, A3 => n20492, ZN => 
                           n19954);
   U6473 : AOI21_X1 port map( A1 => n20440, A2 => n2565, B => n34155, ZN => 
                           n20441);
   U11747 : NAND2_X1 port map( A1 => n1159, A2 => n32201, ZN => n2619);
   U20528 : INV_X1 port map( I => n30929, ZN => n10489);
   U17456 : INV_X1 port map( I => n1344, ZN => n20832);
   U7239 : INV_X1 port map( I => n20698, ZN => n20783);
   U734 : NAND2_X1 port map( A1 => n20899, A2 => n20954, ZN => n4269);
   U11677 : NAND3_X1 port map( A1 => n817, A2 => n20499, A3 => n33116, ZN => 
                           n20500);
   U8408 : OAI21_X1 port map( A1 => n20451, A2 => n16139, B => n20452, ZN => 
                           n2318);
   U6497 : AOI21_X1 port map( A1 => n6530, A2 => n16174, B => n29938, ZN => 
                           n2250);
   U1562 : INV_X1 port map( I => n20963, ZN => n30013);
   U3813 : INV_X1 port map( I => n20729, ZN => n6548);
   U12816 : NOR2_X1 port map( A1 => n30552, A2 => n1909, ZN => n1908);
   U6469 : INV_X1 port map( I => n20849, ZN => n13602);
   U22770 : INV_X1 port map( I => n29898, ZN => n26255);
   U7237 : INV_X1 port map( I => n21043, ZN => n20586);
   U1187 : INV_X1 port map( I => n2198, ZN => n17659);
   U3398 : INV_X1 port map( I => n21016, ZN => n26575);
   U8368 : INV_X1 port map( I => n17423, ZN => n1341);
   U13935 : BUF_X2 port map( I => n1787, Z => n30171);
   U1194 : BUF_X2 port map( I => n16173, Z => n348);
   U1195 : BUF_X2 port map( I => n5572, Z => n28864);
   U8376 : INV_X1 port map( I => n20954, ZN => n4758);
   U717 : INV_X1 port map( I => n20961, ZN => n20183);
   U4200 : INV_X1 port map( I => n20726, ZN => n1338);
   U723 : INV_X1 port map( I => n20862, ZN => n1342);
   U11613 : INV_X1 port map( I => n20905, ZN => n5009);
   U5895 : CLKBUF_X2 port map( I => n20679, Z => n28822);
   U20594 : INV_X1 port map( I => n519, ZN => n924);
   U5477 : NAND2_X1 port map( A1 => n16652, A2 => n14556, ZN => n7756);
   U2223 : NAND2_X1 port map( A1 => n17313, A2 => n28714, ZN => n2230);
   U8343 : INV_X2 port map( I => n28642, ZN => n16785);
   U6459 : INV_X2 port map( I => n1337, ZN => n5883);
   U14875 : NAND2_X1 port map( A1 => n29460, A2 => n26407, ZN => n13130);
   U13964 : INV_X2 port map( I => n3193, ZN => n11967);
   U22158 : INV_X1 port map( I => n28260, ZN => n398);
   U6451 : INV_X1 port map( I => n15226, ZN => n21267);
   U24094 : INV_X1 port map( I => n28594, ZN => n21338);
   U8203 : INV_X2 port map( I => n17313, ZN => n3673);
   U7203 : INV_X2 port map( I => n515, ZN => n2822);
   U7205 : INV_X2 port map( I => n26712, ZN => n21434);
   U19491 : INV_X1 port map( I => n26345, ZN => n30783);
   U20843 : NAND2_X1 port map( A1 => n33498, A2 => n29062, ZN => n13101);
   U4947 : OR2_X1 port map( A1 => n5392, A2 => n8074, Z => n21402);
   U17672 : OAI21_X1 port map( A1 => n11187, A2 => n21189, B => n2822, ZN => 
                           n27515);
   U1663 : NAND2_X1 port map( A1 => n27939, A2 => n21328, ZN => n26326);
   U1133 : INV_X1 port map( I => n21152, ZN => n27689);
   U5551 : AOI21_X1 port map( A1 => n4381, A2 => n21322, B => n1145, ZN => 
                           n7122);
   U19988 : CLKBUF_X2 port map( I => n6855, Z => n30854);
   U2831 : INV_X2 port map( I => n14556, ZN => n921);
   U8602 : INV_X2 port map( I => n21165, ZN => n6075);
   U3005 : NAND2_X1 port map( A1 => n21160, A2 => n17305, ZN => n15428);
   U13744 : INV_X1 port map( I => n11272, ZN => n7822);
   U6462 : INV_X1 port map( I => n21412, ZN => n929);
   U6536 : INV_X1 port map( I => n34089, ZN => n27382);
   U12822 : INV_X2 port map( I => n28668, ZN => n18218);
   U6465 : INV_X2 port map( I => n27028, ZN => n17699);
   U5116 : INV_X1 port map( I => n21221, ZN => n6451);
   U657 : INV_X2 port map( I => n21403, ZN => n1335);
   U14559 : INV_X1 port map( I => n26971, ZN => n27842);
   U23300 : AND2_X1 port map( A1 => n8681, A2 => n17829, Z => n21138);
   U4195 : INV_X1 port map( I => n21233, ZN => n9699);
   U658 : INV_X1 port map( I => n12037, ZN => n1334);
   U5842 : INV_X1 port map( I => n16072, ZN => n21115);
   U15511 : NAND2_X1 port map( A1 => n14290, A2 => n21403, ZN => n21404);
   U3006 : NOR2_X1 port map( A1 => n34157, A2 => n31874, ZN => n21212);
   U690 : INV_X1 port map( I => n601, ZN => n925);
   U18123 : INV_X1 port map( I => n17271, ZN => n21353);
   U10925 : NAND2_X1 port map( A1 => n1018, A2 => n3193, ZN => n21169);
   U23460 : NOR2_X1 port map( A1 => n8490, A2 => n26407, ZN => n15968);
   U18565 : AOI21_X1 port map( A1 => n26014, A2 => n9699, B => n21138, ZN => 
                           n2464);
   U8236 : NAND2_X1 port map( A1 => n8604, A2 => n5049, ZN => n5048);
   U6458 : INV_X8 port map( I => n10533, ZN => n926);
   U8353 : INV_X1 port map( I => n17985, ZN => n21175);
   U24823 : NAND2_X1 port map( A1 => n921, A2 => n16652, ZN => n21052);
   U13105 : OAI21_X1 port map( A1 => n27075, A2 => n21085, B => n21173, ZN => 
                           n2176);
   U10182 : NAND2_X1 port map( A1 => n6075, A2 => n29750, ZN => n31170);
   U8298 : NAND2_X1 port map( A1 => n31909, A2 => n16072, ZN => n15220);
   U11569 : INV_X1 port map( I => n6451, ZN => n2574);
   U24882 : NOR2_X1 port map( A1 => n6408, A2 => n34157, ZN => n21383);
   U9773 : AND2_X1 port map( A1 => n15559, A2 => n28594, Z => n26829);
   U2239 : NAND2_X1 port map( A1 => n7430, A2 => n164, ZN => n21332);
   U22578 : INV_X1 port map( I => n29255, ZN => n21325);
   U22717 : NOR2_X1 port map( A1 => n21407, A2 => n4324, ZN => n14098);
   U17479 : NAND2_X1 port map( A1 => n30784, A2 => n27482, ZN => n3696);
   U628 : NOR2_X1 port map( A1 => n21163, A2 => n1148, ZN => n20881);
   U13168 : INV_X1 port map( I => n10787, ZN => n13194);
   U21129 : NOR2_X1 port map( A1 => n11966, A2 => n21369, ZN => n16313);
   U4791 : CLKBUF_X2 port map( I => n13255, Z => n28886);
   U5865 : CLKBUF_X2 port map( I => n10533, Z => n31826);
   U6514 : INV_X2 port map( I => n1146, ZN => n8011);
   U11523 : NAND2_X1 port map( A1 => n7122, A2 => n7121, ZN => n7120);
   U20944 : NAND2_X1 port map( A1 => n31003, A2 => n27912, ZN => n1982);
   U3146 : INV_X2 port map( I => n17624, ZN => n21192);
   U2568 : INV_X1 port map( I => n29460, ZN => n20676);
   U673 : INV_X1 port map( I => n29256, ZN => n779);
   U11560 : INV_X1 port map( I => n18035, ZN => n3717);
   U636 : INV_X2 port map( I => n1145, ZN => n21321);
   U6518 : INV_X1 port map( I => n17341, ZN => n1019);
   U6445 : INV_X1 port map( I => n21241, ZN => n8453);
   U1423 : NAND2_X1 port map( A1 => n3673, A2 => n7007, ZN => n3672);
   U16731 : NAND2_X1 port map( A1 => n67, A2 => n1632, ZN => n30379);
   U6134 : OR2_X1 port map( A1 => n9663, A2 => n8243, Z => n26021);
   U620 : NOR2_X1 port map( A1 => n32347, A2 => n11912, ZN => n21335);
   U19504 : INV_X1 port map( I => n9322, ZN => n17455);
   U3959 : INV_X1 port map( I => n17305, ZN => n12525);
   U8341 : INV_X1 port map( I => n21239, ZN => n21448);
   U8348 : INV_X1 port map( I => n21306, ZN => n29574);
   U1433 : NOR2_X1 port map( A1 => n6075, A2 => n21085, ZN => n31702);
   U18947 : NOR2_X1 port map( A1 => n31498, A2 => n13730, ZN => n30694);
   U20953 : OAI21_X1 port map( A1 => n21353, A2 => n30784, B => n27075, ZN => 
                           n21082);
   U8559 : NAND2_X1 port map( A1 => n21192, A2 => n21427, ZN => n30889);
   U15876 : NAND3_X1 port map( A1 => n13712, A2 => n21251, A3 => n20662, ZN => 
                           n28340);
   U2578 : NOR2_X1 port map( A1 => n9664, A2 => n926, ZN => n10527);
   U8303 : AOI21_X1 port map( A1 => n7690, A2 => n33745, B => n28641, ZN => 
                           n14722);
   U1100 : OAI21_X1 port map( A1 => n4119, A2 => n30755, B => n21408, ZN => 
                           n14998);
   U17655 : NOR3_X1 port map( A1 => n9518, A2 => n17699, A3 => n29062, ZN => 
                           n1967);
   U22732 : AOI21_X1 port map( A1 => n6584, A2 => n21408, B => n510, ZN => 
                           n31262);
   U22240 : NOR2_X1 port map( A1 => n26861, A2 => n11948, ZN => n21171);
   U5567 : OAI21_X1 port map( A1 => n11457, A2 => n21335, B => n21243, ZN => 
                           n11456);
   U1362 : INV_X1 port map( I => n21354, ZN => n2172);
   U10435 : NAND2_X1 port map( A1 => n31170, A2 => n21173, ZN => n27424);
   U22023 : NAND2_X1 port map( A1 => n8197, A2 => n1337, ZN => n9258);
   U10968 : NAND2_X1 port map( A1 => n29122, A2 => n6908, ZN => n6907);
   U8334 : NOR2_X1 port map( A1 => n21099, A2 => n21252, ZN => n7773);
   U1234 : OAI21_X1 port map( A1 => n4569, A2 => n2676, B => n33106, ZN => 
                           n2834);
   U14333 : NAND3_X1 port map( A1 => n15015, A2 => n599, A3 => n2822, ZN => 
                           n7913);
   U3588 : NOR2_X1 port map( A1 => n31909, A2 => n21406, ZN => n21298);
   U17293 : NAND2_X1 port map( A1 => n10148, A2 => n1020, ZN => n27440);
   U20402 : NOR2_X1 port map( A1 => n8011, A2 => n21434, ZN => n30913);
   U1132 : INV_X1 port map( I => n6908, ZN => n8957);
   U10147 : INV_X1 port map( I => n33641, ZN => n27230);
   U8282 : NOR2_X1 port map( A1 => n10730, A2 => n16459, ZN => n21619);
   U8240 : NOR2_X1 port map( A1 => n8378, A2 => n33882, ZN => n13975);
   U21409 : INV_X1 port map( I => n29062, ZN => n15444);
   U15184 : NOR2_X1 port map( A1 => n7690, A2 => n21223, ZN => n14273);
   U13766 : NOR2_X1 port map( A1 => n21322, A2 => n2822, ZN => n21323);
   U6532 : NAND2_X1 port map( A1 => n21082, A2 => n26861, ZN => n15961);
   U7146 : INV_X1 port map( I => n21619, ZN => n11265);
   U1285 : NOR2_X1 port map( A1 => n12746, A2 => n13921, ZN => n28074);
   U11471 : OAI21_X1 port map( A1 => n20795, A2 => n28287, B => n33641, ZN => 
                           n16046);
   U2695 : AOI22_X1 port map( A1 => n21320, A2 => n28017, B1 => n21323, B2 => 
                           n11187, ZN => n29799);
   U616 : AOI21_X1 port map( A1 => n21054, A2 => n5111, B => n14643, ZN => 
                           n10980);
   U1405 : NAND2_X1 port map( A1 => n5575, A2 => n21452, ZN => n9392);
   U9618 : NAND2_X1 port map( A1 => n21381, A2 => n21209, ZN => n10733);
   U8235 : OAI21_X1 port map( A1 => n13975, A2 => n21120, B => n12363, ZN => 
                           n12373);
   U24931 : NAND3_X1 port map( A1 => n21411, A2 => n34037, A3 => n11315, ZN => 
                           n28699);
   U1327 : NOR2_X1 port map( A1 => n16180, A2 => n21443, ZN => n31507);
   U1381 : AOI22_X1 port map( A1 => n31673, A2 => n18218, B1 => n8539, B2 => 
                           n1911, ZN => n1910);
   U22915 : NAND2_X1 port map( A1 => n21169, A2 => n10092, ZN => n28385);
   U20869 : AOI22_X1 port map( A1 => n12324, A2 => n21398, B1 => n3933, B2 => 
                           n12325, ZN => n21399);
   U11459 : OAI21_X1 port map( A1 => n30727, A2 => n10113, B => n8727, ZN => 
                           n7543);
   U4703 : NAND2_X1 port map( A1 => n26018, A2 => n20936, ZN => n28299);
   U9714 : NOR2_X1 port map( A1 => n8378, A2 => n7430, ZN => n11480);
   U9689 : NOR2_X1 port map( A1 => n7430, A2 => n12925, ZN => n7446);
   U9631 : OAI21_X1 port map( A1 => n14273, A2 => n21317, B => n15261, ZN => 
                           n14272);
   U23659 : NAND2_X1 port map( A1 => n15622, A2 => n779, ZN => n28526);
   U14613 : NOR2_X1 port map( A1 => n17011, A2 => n10527, ZN => n30246);
   U26419 : NAND3_X1 port map( A1 => n11456, A2 => n21069, A3 => n17666, ZN => 
                           n13442);
   U3468 : NAND2_X1 port map( A1 => n21447, A2 => n31730, ZN => n21824);
   U14883 : NAND2_X1 port map( A1 => n21264, A2 => n11745, ZN => n16851);
   U1112 : AOI21_X1 port map( A1 => n1329, A2 => n21109, B => n26167, ZN => 
                           n26166);
   U1300 : INV_X1 port map( I => n21738, ZN => n21864);
   U5830 : INV_X1 port map( I => n196, ZN => n14397);
   U17841 : OAI21_X1 port map( A1 => n29382, A2 => n30544, B => n21443, ZN => 
                           n31853);
   U9650 : OAI21_X1 port map( A1 => n11979, A2 => n12521, B => n32907, ZN => 
                           n21089);
   U9231 : OAI21_X1 port map( A1 => n28074, A2 => n25942, B => n32347, ZN => 
                           n6880);
   U2590 : NOR2_X1 port map( A1 => n6879, A2 => n6881, ZN => n6878);
   U24887 : AOI22_X1 port map( A1 => n21420, A2 => n21419, B1 => n33649, B2 => 
                           n21418, ZN => n21421);
   U2304 : NAND2_X1 port map( A1 => n6212, A2 => n16553, ZN => n21462);
   U25924 : NAND2_X1 port map( A1 => n3973, A2 => n16046, ZN => n8875);
   U21957 : INV_X2 port map( I => n15091, ZN => n1312);
   U20255 : AOI21_X1 port map( A1 => n21200, A2 => n10686, B => n9721, ZN => 
                           n16546);
   U562 : INV_X1 port map( I => n13652, ZN => n21736);
   U5402 : INV_X1 port map( I => n8457, ZN => n1016);
   U1212 : INV_X1 port map( I => n13884, ZN => n16157);
   U6383 : INV_X1 port map( I => n17716, ZN => n1321);
   U5811 : CLKBUF_X2 port map( I => n16222, Z => n8079);
   U2582 : BUF_X2 port map( I => n9999, Z => n2296);
   U1255 : INV_X2 port map( I => n31911, ZN => n30440);
   U5404 : INV_X2 port map( I => n13114, ZN => n1013);
   U1215 : INV_X2 port map( I => n10720, ZN => n861);
   U9305 : INV_X1 port map( I => n27954, ZN => n916);
   U17120 : INV_X1 port map( I => n27379, ZN => n21672);
   U4325 : INV_X2 port map( I => n17888, ZN => n11596);
   U15800 : AND2_X1 port map( A1 => n18208, A2 => n18206, Z => n27178);
   U25923 : INV_X1 port map( I => n8875, ZN => n21858);
   U1018 : INV_X2 port map( I => n30769, ZN => n11300);
   U18795 : INV_X1 port map( I => n30389, ZN => n30677);
   U1156 : INV_X1 port map( I => n21816, ZN => n912);
   U3365 : NOR2_X1 port map( A1 => n16157, A2 => n21122, ZN => n29784);
   U1269 : INV_X1 port map( I => n16023, ZN => n10254);
   U2573 : NAND2_X1 port map( A1 => n920, A2 => n21733, ZN => n185);
   U5558 : NAND2_X1 port map( A1 => n230, A2 => n21706, ZN => n6351);
   U10172 : OAI21_X1 port map( A1 => n11300, A2 => n17348, B => n32252, ZN => 
                           n4434);
   U1159 : NAND2_X1 port map( A1 => n21518, A2 => n916, ZN => n29690);
   U1166 : INV_X1 port map( I => n33766, ZN => n11276);
   U9550 : INV_X2 port map( I => n21730, ZN => n17773);
   U13969 : INV_X1 port map( I => n11756, ZN => n12711);
   U585 : NAND2_X1 port map( A1 => n1009, A2 => n21832, ZN => n15813);
   U1038 : INV_X1 port map( I => n31102, ZN => n26727);
   U9503 : AOI21_X1 port map( A1 => n16864, A2 => n16863, B => n31458, ZN => 
                           n16445);
   U8206 : NAND2_X1 port map( A1 => n31957, A2 => n2368, ZN => n14848);
   U11103 : INV_X1 port map( I => n3379, ZN => n10532);
   U3802 : NAND2_X1 port map( A1 => n1321, A2 => n3420, ZN => n31732);
   U1197 : INV_X1 port map( I => n21852, ZN => n8706);
   U15695 : INV_X1 port map( I => n32904, ZN => n862);
   U11344 : INV_X1 port map( I => n17274, ZN => n21535);
   U11872 : NOR2_X1 port map( A1 => n29947, A2 => n1008, ZN => n5342);
   U11831 : NOR2_X1 port map( A1 => n9590, A2 => n9591, ZN => n9589);
   U5589 : CLKBUF_X2 port map( I => n13652, Z => n28018);
   U20806 : NAND3_X1 port map( A1 => n6231, A2 => n3250, A3 => n29180, ZN => 
                           n31645);
   U11405 : INV_X1 port map( I => n32252, ZN => n3140);
   U8639 : INV_X1 port map( I => n31859, ZN => n31910);
   U4629 : OAI21_X1 port map( A1 => n727, A2 => n7592, B => n21496, ZN => n2514
                           );
   U16512 : INV_X1 port map( I => n14236, ZN => n1138);
   U4554 : INV_X1 port map( I => n9999, ZN => n11890);
   U18190 : AND2_X1 port map( A1 => n12866, A2 => n17431, Z => n21459);
   U1025 : AND2_X1 port map( A1 => n15863, A2 => n28429, Z => n534);
   U4389 : INV_X1 port map( I => n5170, ZN => n21625);
   U3675 : INV_X1 port map( I => n31309, ZN => n11499);
   U24911 : NAND2_X1 port map( A1 => n30885, A2 => n27635, ZN => n21529);
   U4657 : CLKBUF_X2 port map( I => n21767, Z => n28395);
   U5399 : BUF_X8 port map( I => n4029, Z => n3467);
   U17971 : OAI21_X1 port map( A1 => n1009, A2 => n33981, B => n11890, ZN => 
                           n6969);
   U1107 : NOR2_X1 port map( A1 => n432, A2 => n29302, ZN => n12028);
   U24859 : NAND3_X1 port map( A1 => n27560, A2 => n29854, A3 => n21730, ZN => 
                           n21277);
   U558 : NAND2_X1 port map( A1 => n10775, A2 => n21603, ZN => n5851);
   U4548 : NOR3_X1 port map( A1 => n11861, A2 => n31654, A3 => n21780, ZN => 
                           n28141);
   U1139 : NOR2_X1 port map( A1 => n5546, A2 => n6544, ZN => n4311);
   U4774 : AND2_X1 port map( A1 => n30832, A2 => n7811, Z => n27466);
   U4587 : OAI22_X1 port map( A1 => n28654, A2 => n1318, B1 => n21671, B2 => 
                           n918, ZN => n14541);
   U20737 : NOR2_X1 port map( A1 => n27596, A2 => n21632, ZN => n30962);
   U1013 : NOR2_X1 port map( A1 => n32519, A2 => n17887, ZN => n8403);
   U22943 : NAND2_X1 port map( A1 => n15838, A2 => n14681, ZN => n15837);
   U2580 : NOR2_X1 port map( A1 => n32865, A2 => n2296, ZN => n2298);
   U22469 : NAND3_X1 port map( A1 => n2217, A2 => n21628, A3 => n29322, ZN => 
                           n21574);
   U1127 : NAND2_X1 port map( A1 => n11861, A2 => n31317, ZN => n4212);
   U10778 : AOI21_X1 port map( A1 => n21535, A2 => n21566, B => n21351, ZN => 
                           n9884);
   U1086 : INV_X1 port map( I => n14595, ZN => n30114);
   U21522 : NAND2_X1 port map( A1 => n21581, A2 => n13133, ZN => n16723);
   U23870 : NOR2_X1 port map( A1 => n21571, A2 => n30678, ZN => n21572);
   U919 : OAI21_X1 port map( A1 => n17428, A2 => n21459, B => n21730, ZN => 
                           n13199);
   U24909 : NOR2_X1 port map( A1 => n21781, A2 => n31220, ZN => n21523);
   U1747 : NOR2_X1 port map( A1 => n7326, A2 => n11797, ZN => n7325);
   U11335 : INV_X1 port map( I => n11619, ZN => n13248);
   U532 : NOR2_X1 port map( A1 => n12275, A2 => n12274, ZN => n12273);
   U3901 : NAND2_X1 port map( A1 => n28824, A2 => n5309, ZN => n14948);
   U1124 : NAND2_X1 port map( A1 => n31711, A2 => n28018, ZN => n28067);
   U1782 : BUF_X2 port map( I => n14691, Z => n1);
   U1931 : NAND2_X1 port map( A1 => n17406, A2 => n21830, ZN => n21831);
   U17012 : NOR2_X1 port map( A1 => n6544, A2 => n6489, ZN => n4359);
   U9575 : NOR2_X1 port map( A1 => n21777, A2 => n21743, ZN => n21744);
   U2585 : AOI21_X1 port map( A1 => n10699, A2 => n30441, B => n30440, ZN => 
                           n26671);
   U1422 : INV_X1 port map( I => n16147, ZN => n21817);
   U5124 : INV_X1 port map( I => n26445, ZN => n1014);
   U6427 : INV_X1 port map( I => n28450, ZN => n864);
   U1063 : AND2_X1 port map( A1 => n21573, A2 => n29322, Z => n21607);
   U23153 : INV_X1 port map( I => n21832, ZN => n15242);
   U16913 : NOR2_X1 port map( A1 => n3539, A2 => n21781, ZN => n17019);
   U4390 : NOR2_X1 port map( A1 => n1135, A2 => n3468, ZN => n8230);
   U9583 : NOR2_X1 port map( A1 => n7553, A2 => n29234, ZN => n13500);
   U17358 : INV_X1 port map( I => n32519, ZN => n21701);
   U17590 : NOR2_X1 port map( A1 => n29084, A2 => n11861, ZN => n17018);
   U5094 : AOI22_X1 port map( A1 => n21794, A2 => n15838, B1 => n21793, B2 => 
                           n21792, ZN => n21795);
   U7065 : AOI21_X1 port map( A1 => n21666, A2 => n1312, B => n16577, ZN => 
                           n2178);
   U2935 : NAND3_X1 port map( A1 => n16194, A2 => n29302, A3 => n31458, ZN => 
                           n21548);
   U1054 : OAI21_X1 port map( A1 => n31335, A2 => n915, B => n11499, ZN => 
                           n11552);
   U21991 : OAI21_X1 port map( A1 => n27704, A2 => n32865, B => n1009, ZN => 
                           n4131);
   U14322 : NOR2_X1 port map( A1 => n27065, A2 => n1317, ZN => n16163);
   U8143 : NAND2_X1 port map( A1 => n5546, A2 => n1138, ZN => n2709);
   U2581 : AOI22_X1 port map( A1 => n2298, A2 => n21625, B1 => n2296, B2 => 
                           n396, ZN => n2297);
   U11391 : NAND2_X1 port map( A1 => n33146, A2 => n1133, ZN => n4262);
   U6381 : NAND2_X1 port map( A1 => n1647, A2 => n21520, ZN => n1770);
   U8142 : NAND2_X1 port map( A1 => n21852, A2 => n5546, ZN => n2710);
   U19647 : NAND2_X1 port map( A1 => n28729, A2 => n7813, ZN => n12605);
   U5817 : NAND3_X1 port map( A1 => n3467, A2 => n17077, A3 => n3468, ZN => 
                           n3469);
   U11298 : NAND2_X1 port map( A1 => n21701, A2 => n17887, ZN => n15316);
   U4658 : INV_X1 port map( I => n27704, ZN => n6967);
   U19852 : NAND2_X1 port map( A1 => n12751, A2 => n32076, ZN => n11448);
   U9520 : NAND2_X1 port map( A1 => n21657, A2 => n8886, ZN => n14829);
   U5606 : AOI21_X1 port map( A1 => n21566, A2 => n3315, B => n21570, ZN => 
                           n3314);
   U9543 : OAI21_X1 port map( A1 => n17019, A2 => n17018, B => n31220, ZN => 
                           n17017);
   U1066 : NAND2_X1 port map( A1 => n30548, A2 => n3588, ZN => n21525);
   U7059 : NAND2_X1 port map( A1 => n7366, A2 => n7365, ZN => n21680);
   U1033 : OAI22_X1 port map( A1 => n32071, A2 => n30549, B1 => n21594, B2 => 
                           n21595, ZN => n21597);
   U7083 : NAND2_X1 port map( A1 => n1326, A2 => n15864, ZN => n16012);
   U26464 : INV_X1 port map( I => n34084, ZN => n1531);
   U519 : OR2_X1 port map( A1 => n16796, A2 => n16192, Z => n3722);
   U3222 : INV_X1 port map( I => n8269, ZN => n1607);
   U20926 : OAI21_X1 port map( A1 => n1531, A2 => n21804, B => n11231, ZN => 
                           n30999);
   U9083 : AOI22_X1 port map( A1 => n29393, A2 => n3467, B1 => n1135, B2 => 
                           n4699, ZN => n13540);
   U22104 : NOR2_X1 port map( A1 => n21805, A2 => n3468, ZN => n21722);
   U15450 : AOI22_X1 port map( A1 => n26113, A2 => n16147, B1 => n6626, B2 => 
                           n1015, ZN => n4880);
   U5093 : BUF_X2 port map( I => n17697, Z => n4057);
   U15766 : NAND3_X1 port map( A1 => n27103, A2 => n5757, A3 => n33571, ZN => 
                           n30306);
   U15950 : BUF_X2 port map( I => n22249, Z => n2353);
   U11262 : INV_X1 port map( I => n8392, ZN => n1308);
   U1042 : INV_X1 port map( I => n22137, ZN => n6812);
   U11221 : NAND2_X1 port map( A1 => n910, A2 => n17362, ZN => n6206);
   U2271 : INV_X1 port map( I => n34078, ZN => n2308);
   U1605 : NAND2_X1 port map( A1 => n26875, A2 => n22047, ZN => n1609);
   U13604 : NAND2_X1 port map( A1 => n21945, A2 => n12594, ZN => n2777);
   U7028 : INV_X1 port map( I => n6771, ZN => n22128);
   U7618 : INV_X1 port map( I => n27767, ZN => n29501);
   U13520 : INV_X1 port map( I => n29693, ZN => n26942);
   U22737 : INV_X1 port map( I => n22302, ZN => n14125);
   U1024 : INV_X1 port map( I => n9809, ZN => n21959);
   U9481 : INV_X1 port map( I => n22294, ZN => n2554);
   U26198 : INV_X2 port map( I => n22681, ZN => n31701);
   U19066 : INV_X1 port map( I => n8452, ZN => n10680);
   U13958 : INV_X4 port map( I => n27004, ZN => n22330);
   U1253 : INV_X2 port map( I => n5640, ZN => n10724);
   U3848 : INV_X1 port map( I => n14307, ZN => n22578);
   U14614 : INV_X1 port map( I => n32081, ZN => n12530);
   U16897 : NAND2_X1 port map( A1 => n33466, A2 => n22647, ZN => n6187);
   U5631 : INV_X1 port map( I => n5657, ZN => n12733);
   U4836 : BUF_X2 port map( I => n21941, Z => n22645);
   U3296 : BUF_X2 port map( I => n22199, Z => n11895);
   U5800 : INV_X1 port map( I => n34162, ZN => n1119);
   U3928 : INV_X1 port map( I => n22332, ZN => n2417);
   U2741 : INV_X1 port map( I => n22625, ZN => n22497);
   U18662 : INV_X1 port map( I => n8099, ZN => n22547);
   U3076 : INV_X2 port map( I => n16567, ZN => n22666);
   U20732 : INV_X1 port map( I => n11749, ZN => n16558);
   U7048 : INV_X1 port map( I => n27897, ZN => n645);
   U6713 : INV_X1 port map( I => n10680, ZN => n9456);
   U1315 : INV_X2 port map( I => n10568, ZN => n14376);
   U15233 : INV_X2 port map( I => n22547, ZN => n22550);
   U8089 : INV_X1 port map( I => n21869, ZN => n22678);
   U9468 : INV_X1 port map( I => n8471, ZN => n22398);
   U13102 : INV_X2 port map( I => n29304, ZN => n905);
   U3489 : INV_X2 port map( I => n9515, ZN => n22574);
   U6687 : NOR2_X1 port map( A1 => n22681, A2 => n10354, ZN => n9802);
   U3705 : CLKBUF_X2 port map( I => n22414, Z => n137);
   U5381 : NOR2_X1 port map( A1 => n16567, A2 => n16149, ZN => n15805);
   U19539 : INV_X2 port map( I => n9234, ZN => n9370);
   U4112 : BUF_X2 port map( I => n637, Z => n14728);
   U9463 : INV_X2 port map( I => n9910, ZN => n3495);
   U23959 : INV_X2 port map( I => n634, ZN => n22626);
   U456 : INV_X2 port map( I => n12076, ZN => n900);
   U5798 : INV_X1 port map( I => n22597, ZN => n11930);
   U1529 : INV_X1 port map( I => n17879, ZN => n22667);
   U7757 : INV_X2 port map( I => n9959, ZN => n29508);
   U11205 : INV_X1 port map( I => n22452, ZN => n6658);
   U2047 : INV_X1 port map( I => n22340, ZN => n1300);
   U4924 : INV_X2 port map( I => n15089, ZN => n11874);
   U4369 : NAND2_X1 port map( A1 => n17147, A2 => n8965, ZN => n18038);
   U9399 : OAI21_X1 port map( A1 => n1290, A2 => n22588, B => n22584, ZN => 
                           n15007);
   U5643 : NAND3_X1 port map( A1 => n2417, A2 => n16334, A3 => n12733, ZN => 
                           n7053);
   U22682 : NAND2_X1 port map( A1 => n14376, A2 => n29304, ZN => n9751);
   U6705 : NOR3_X1 port map( A1 => n29261, A2 => n900, A3 => n22394, ZN => 
                           n13154);
   U9430 : NAND2_X1 port map( A1 => n9578, A2 => n22599, ZN => n9579);
   U5373 : OAI21_X1 port map( A1 => n22401, A2 => n27390, B => n32449, ZN => 
                           n6749);
   U4098 : INV_X1 port map( I => n637, ZN => n901);
   U5670 : NOR2_X1 port map( A1 => n1116, A2 => n22672, ZN => n12632);
   U7637 : NAND2_X1 port map( A1 => n9022, A2 => n10612, ZN => n11419);
   U8014 : NAND2_X1 port map( A1 => n10206, A2 => n856, ZN => n6709);
   U421 : NAND2_X1 port map( A1 => n22389, A2 => n33966, ZN => n17357);
   U866 : INV_X2 port map( I => n11932, ZN => n26173);
   U498 : INV_X1 port map( I => n5379, ZN => n904);
   U5787 : AOI21_X1 port map( A1 => n22574, A2 => n16503, B => n2471, ZN => 
                           n12888);
   U1443 : INV_X1 port map( I => n2538, ZN => n17123);
   U926 : NAND2_X1 port map( A1 => n22549, A2 => n30668, ZN => n25947);
   U468 : INV_X2 port map( I => n11920, ZN => n22478);
   U21999 : BUF_X2 port map( I => n11916, Z => n28669);
   U13576 : NAND2_X1 port map( A1 => n468, A2 => n33964, ZN => n22442);
   U15542 : INV_X1 port map( I => n33739, ZN => n708);
   U14853 : INV_X2 port map( I => n28378, ZN => n22483);
   U3170 : NAND2_X1 port map( A1 => n4425, A2 => n22636, ZN => n14478);
   U5803 : INV_X2 port map( I => n28825, ZN => n4459);
   U21847 : AND2_X1 port map( A1 => n22656, A2 => n17899, Z => n22583);
   U2749 : INV_X1 port map( I => n1127, ZN => n858);
   U8208 : NAND3_X1 port map( A1 => n1125, A2 => n22584, A3 => n1290, ZN => 
                           n29557);
   U4556 : BUF_X2 port map( I => n22580, Z => n26878);
   U826 : INV_X2 port map( I => n17764, ZN => n908);
   U15795 : INV_X1 port map( I => n9578, ZN => n13078);
   U19666 : NOR3_X1 port map( A1 => n16558, A2 => n31914, A3 => n22638, ZN => 
                           n15609);
   U7748 : OAI21_X1 port map( A1 => n15805, A2 => n22576, B => n26453, ZN => 
                           n27411);
   U18298 : AOI21_X1 port map( A1 => n16531, A2 => n22612, B => n855, ZN => 
                           n7464);
   U21751 : INV_X1 port map( I => n468, ZN => n22567);
   U918 : NAND2_X1 port map( A1 => n22666, A2 => n22577, ZN => n12439);
   U13026 : NAND2_X1 port map( A1 => n1300, A2 => n22622, ZN => n22623);
   U3057 : NAND3_X1 port map( A1 => n1633, A2 => n2697, A3 => n28568, ZN => 
                           n11376);
   U18055 : NOR2_X1 port map( A1 => n22505, A2 => n14728, ZN => n27574);
   U11112 : NOR2_X1 port map( A1 => n22646, A2 => n4459, ZN => n7850);
   U1713 : NAND2_X1 port map( A1 => n22537, A2 => n17147, ZN => n12698);
   U6305 : AOI21_X1 port map( A1 => n1842, A2 => n30668, B => n30669, ZN => 
                           n22482);
   U709 : NOR2_X1 port map( A1 => n16434, A2 => n8965, ZN => n16549);
   U11192 : NOR2_X1 port map( A1 => n22450, A2 => n17764, ZN => n2657);
   U7026 : INV_X1 port map( I => n31931, ZN => n22691);
   U6715 : NOR2_X1 port map( A1 => n15752, A2 => n16483, ZN => n14228);
   U21038 : NAND2_X1 port map( A1 => n22475, A2 => n22474, ZN => n17248);
   U5377 : AOI21_X1 port map( A1 => n17185, A2 => n10862, B => n8919, ZN => 
                           n2486);
   U20888 : NAND2_X1 port map( A1 => n8912, A2 => n17185, ZN => n13874);
   U9445 : NOR2_X1 port map( A1 => n16434, A2 => n22429, ZN => n9425);
   U835 : NOR3_X1 port map( A1 => n22330, A2 => n14376, A3 => n902, ZN => 
                           n29957);
   U8088 : NOR2_X1 port map( A1 => n1116, A2 => n905, ZN => n29541);
   U20828 : NAND2_X1 port map( A1 => n14231, A2 => n33966, ZN => n15450);
   U21257 : OAI21_X1 port map( A1 => n22576, A2 => n16567, B => n6658, ZN => 
                           n15379);
   U12887 : CLKBUF_X2 port map( I => n22599, Z => n30066);
   U874 : NOR2_X1 port map( A1 => n6401, A2 => n9653, ZN => n6432);
   U18640 : AOI21_X1 port map( A1 => n239, A2 => n7090, B => n16137, ZN => 
                           n2383);
   U4829 : NAND2_X1 port map( A1 => n22402, A2 => n9739, ZN => n13249);
   U767 : INV_X1 port map( I => n22634, ZN => n1291);
   U676 : NAND2_X1 port map( A1 => n5743, A2 => n9958, ZN => n22924);
   U8913 : OAI21_X1 port map( A1 => n17185, A2 => n26410, B => n32449, ZN => 
                           n26409);
   U4346 : INV_X1 port map( I => n29928, ZN => n5960);
   U2570 : NAND2_X1 port map( A1 => n2381, A2 => n7090, ZN => n30510);
   U7040 : INV_X1 port map( I => n22486, ZN => n1296);
   U11166 : INV_X1 port map( I => n7561, ZN => n7560);
   U25807 : NAND2_X1 port map( A1 => n1633, A2 => n17890, ZN => n15448);
   U848 : OAI22_X1 port map( A1 => n11928, A2 => n15379, B1 => n22454, B2 => 
                           n6658, ZN => n26799);
   U5683 : NAND2_X1 port map( A1 => n6956, A2 => n21963, ZN => n29632);
   U13557 : AOI21_X1 port map( A1 => n13525, A2 => n34058, B => n22651, ZN => 
                           n13524);
   U9336 : NAND2_X1 port map( A1 => n11161, A2 => n22670, ZN => n1579);
   U5771 : NAND3_X1 port map( A1 => n10907, A2 => n28669, A3 => n8801, ZN => 
                           n22459);
   U3064 : NAND2_X1 port map( A1 => n22388, A2 => n1633, ZN => n6063);
   U2750 : NAND2_X1 port map( A1 => n7239, A2 => n6072, ZN => n2408);
   U18502 : NAND3_X1 port map( A1 => n13534, A2 => n12072, A3 => n22478, ZN => 
                           n30631);
   U8912 : AOI21_X1 port map( A1 => n17185, A2 => n8912, B => n26409, ZN => 
                           n26408);
   U9341 : OAI21_X1 port map( A1 => n17960, A2 => n12335, B => n12333, ZN => 
                           n22011);
   U18868 : NOR2_X1 port map( A1 => n7851, A2 => n7850, ZN => n30688);
   U12067 : NAND2_X1 port map( A1 => n26813, A2 => n1658, ZN => n3670);
   U11159 : INV_X1 port map( I => n22633, ZN => n7400);
   U5372 : NAND3_X1 port map( A1 => n992, A2 => n1286, A3 => n10907, ZN => 
                           n13895);
   U15917 : INV_X2 port map( I => n23056, ZN => n31437);
   U8430 : NAND2_X1 port map( A1 => n4100, A2 => n4459, ZN => n5896);
   U5654 : INV_X1 port map( I => n22523, ZN => n28938);
   U12997 : OAI21_X1 port map( A1 => n29078, A2 => n17764, B => n26867, ZN => 
                           n4996);
   U6276 : NAND2_X1 port map( A1 => n13895, A2 => n13892, ZN => n4700);
   U778 : NAND2_X1 port map( A1 => n7802, A2 => n22968, ZN => n12471);
   U9291 : OAI21_X1 port map( A1 => n32055, A2 => n12952, B => n9580, ZN => 
                           n229);
   U792 : AOI22_X1 port map( A1 => n22594, A2 => n32831, B1 => n4918, B2 => 
                           n22651, ZN => n29598);
   U12930 : OAI21_X1 port map( A1 => n26065, A2 => n26862, B => n1117, ZN => 
                           n8667);
   U773 : INV_X2 port map( I => n22986, ZN => n29242);
   U11075 : OAI21_X1 port map( A1 => n5597, A2 => n1120, B => n2253, ZN => 
                           n2252);
   U18443 : NOR2_X1 port map( A1 => n22471, A2 => n31019, ZN => n17630);
   U23174 : NAND3_X1 port map( A1 => n10282, A2 => n10354, A3 => n31701, ZN => 
                           n22472);
   U12215 : BUF_X2 port map( I => n15299, Z => n11268);
   U21083 : INV_X2 port map( I => n28077, ZN => n641);
   U1023 : NAND2_X1 port map( A1 => n16501, A2 => n16267, ZN => n11018);
   U2373 : INV_X1 port map( I => n13129, ZN => n6782);
   U6924 : INV_X2 port map( I => n22786, ZN => n26667);
   U18461 : INV_X1 port map( I => n30868, ZN => n1112);
   U5065 : INV_X1 port map( I => n17462, ZN => n1269);
   U6260 : NOR2_X1 port map( A1 => n26251, A2 => n23031, ZN => n6876);
   U2636 : NAND2_X1 port map( A1 => n15301, A2 => n17855, ZN => n22761);
   U21994 : NOR2_X1 port map( A1 => n26667, A2 => n32510, ZN => n28648);
   U15370 : INV_X2 port map( I => n16280, ZN => n16976);
   U15232 : NOR2_X1 port map( A1 => n28313, A2 => n22894, ZN => n12377);
   U712 : INV_X2 port map( I => n641, ZN => n12259);
   U662 : BUF_X2 port map( I => n12701, Z => n3891);
   U15662 : BUF_X2 port map( I => n13063, Z => n28415);
   U3498 : CLKBUF_X2 port map( I => n22960, Z => n8334);
   U627 : INV_X2 port map( I => n22951, ZN => n28408);
   U24869 : INV_X2 port map( I => n31505, ZN => n2635);
   U17880 : NAND2_X1 port map( A1 => n28227, A2 => n31549, ZN => n5205);
   U12547 : INV_X1 port map( I => n3670, ZN => n22748);
   U8649 : INV_X2 port map( I => n29610, ZN => n15718);
   U4513 : INV_X1 port map( I => n22950, ZN => n2479);
   U732 : INV_X1 port map( I => n722, ZN => n31358);
   U17615 : INV_X1 port map( I => n7802, ZN => n22965);
   U14395 : INV_X1 port map( I => n23065, ZN => n898);
   U3479 : INV_X1 port map( I => n22885, ZN => n29958);
   U699 : NAND2_X1 port map( A1 => n22983, A2 => n8040, ZN => n28234);
   U2728 : NAND2_X1 port map( A1 => n28974, A2 => n22933, ZN => n2912);
   U5679 : NOR2_X1 port map( A1 => n22780, A2 => n29175, ZN => n29174);
   U2128 : NAND2_X1 port map( A1 => n22473, A2 => n27589, ZN => n7943);
   U10866 : BUF_X2 port map( I => n758, Z => n26612);
   U18597 : AOI22_X1 port map( A1 => n1278, A2 => n6975, B1 => n23010, B2 => 
                           n23014, ZN => n23016);
   U684 : OAI21_X1 port map( A1 => n27639, A2 => n23083, B => n26243, ZN => 
                           n30202);
   U670 : NAND2_X1 port map( A1 => n13778, A2 => n27580, ZN => n12417);
   U9780 : NAND2_X1 port map( A1 => n28328, A2 => n29314, ZN => n26499);
   U678 : NAND2_X1 port map( A1 => n22946, A2 => n23034, ZN => n5095);
   U672 : AOI21_X1 port map( A1 => n897, A2 => n15704, B => n10031, ZN => 
                           n11084);
   U6832 : OAI21_X1 port map( A1 => n23103, A2 => n23104, B => n3600, ZN => 
                           n5400);
   U739 : NOR2_X1 port map( A1 => n23107, A2 => n23106, ZN => n31455);
   U6812 : NAND2_X1 port map( A1 => n17211, A2 => n27719, ZN => n10895);
   U560 : INV_X2 port map( I => n10031, ZN => n983);
   U12893 : NOR2_X1 port map( A1 => n31358, A2 => n29384, ZN => n26222);
   U20900 : AOI21_X1 port map( A1 => n27798, A2 => n28680, B => n22988, ZN => 
                           n22993);
   U528 : NOR2_X1 port map( A1 => n28867, A2 => n9213, ZN => n15317);
   U3557 : NAND2_X1 port map( A1 => n14129, A2 => n22968, ZN => n23088);
   U5704 : NOR2_X1 port map( A1 => n12259, A2 => n27556, ZN => n27555);
   U9289 : INV_X1 port map( I => n22962, ZN => n23081);
   U2164 : NAND2_X1 port map( A1 => n22956, A2 => n987, ZN => n6592);
   U2816 : NOR3_X1 port map( A1 => n9293, A2 => n10031, A3 => n22876, ZN => 
                           n10030);
   U4115 : INV_X1 port map( I => n22399, ZN => n23043);
   U361 : INV_X1 port map( I => n22955, ZN => n852);
   U17164 : NAND2_X1 port map( A1 => n32119, A2 => n15851, ZN => n5618);
   U7917 : INV_X1 port map( I => n31937, ZN => n22866);
   U4515 : INV_X1 port map( I => n17161, ZN => n1265);
   U15674 : INV_X1 port map( I => n22919, ZN => n22880);
   U5336 : AND2_X1 port map( A1 => n15324, A2 => n22856, Z => n3296);
   U741 : INV_X2 port map( I => n28659, ZN => n14188);
   U3564 : INV_X1 port map( I => n15501, ZN => n989);
   U5341 : INV_X1 port map( I => n23070, ZN => n1277);
   U4452 : AND2_X1 port map( A1 => n6605, A2 => n22894, Z => n22769);
   U1181 : CLKBUF_X2 port map( I => n14045, Z => n16254);
   U15665 : NAND2_X1 port map( A1 => n23034, A2 => n13063, ZN => n22892);
   U2611 : NAND2_X1 port map( A1 => n23033, A2 => n22894, ZN => n23037);
   U6965 : INV_X1 port map( I => n23110, ZN => n6453);
   U14709 : NOR2_X1 port map( A1 => n6985, A2 => n23082, ZN => n13396);
   U546 : NAND3_X1 port map( A1 => n32868, A2 => n803, A3 => n14183, ZN => 
                           n4710);
   U23825 : NAND3_X1 port map( A1 => n1581, A2 => n22961, A3 => n8334, ZN => 
                           n13365);
   U14750 : NAND3_X1 port map( A1 => n18261, A2 => n986, A3 => n26667, ZN => 
                           n22789);
   U549 : OAI21_X1 port map( A1 => n4489, A2 => n23050, B => n25994, ZN => 
                           n4488);
   U2318 : NAND2_X1 port map( A1 => n853, A2 => n23108, ZN => n22614);
   U9271 : NAND2_X1 port map( A1 => n14797, A2 => n33382, ZN => n3851);
   U2372 : NAND3_X1 port map( A1 => n28659, A2 => n22982, A3 => n22983, ZN => 
                           n12702);
   U355 : NAND3_X1 port map( A1 => n6800, A2 => n22655, A3 => n28408, ZN => 
                           n22276);
   U14942 : AOI21_X1 port map( A1 => n22876, A2 => n10031, B => n11268, ZN => 
                           n15298);
   U15880 : NAND2_X1 port map( A1 => n898, A2 => n22826, ZN => n22863);
   U23053 : NAND3_X1 port map( A1 => n32868, A2 => n23158, A3 => n13751, ZN => 
                           n4713);
   U16748 : NAND2_X1 port map( A1 => n22738, A2 => n14610, ZN => n8381);
   U2583 : NOR3_X1 port map( A1 => n990, A2 => n1278, A3 => n4599, ZN => n4652)
                           ;
   U21258 : NOR2_X1 port map( A1 => n13159, A2 => n16078, ZN => n13635);
   U4506 : NOR2_X1 port map( A1 => n23079, A2 => n22885, ZN => n13411);
   U11008 : OAI21_X1 port map( A1 => n29242, A2 => n31867, B => n28328, ZN => 
                           n7744);
   U23542 : NOR2_X1 port map( A1 => n6592, A2 => n9778, ZN => n6591);
   U19423 : NOR2_X1 port map( A1 => n23111, A2 => n1264, ZN => n27835);
   U2269 : NAND2_X1 port map( A1 => n6012, A2 => n16022, ZN => n22725);
   U7928 : NAND2_X1 port map( A1 => n22760, A2 => n27612, ZN => n22410);
   U17430 : NAND2_X1 port map( A1 => n10360, A2 => n27389, ZN => n6370);
   U21543 : NOR2_X1 port map( A1 => n31854, A2 => n22780, ZN => n22739);
   U25150 : NOR2_X1 port map( A1 => n28867, A2 => n23101, ZN => n22842);
   U20488 : NAND2_X1 port map( A1 => n18240, A2 => n22774, ZN => n11204);
   U6919 : OAI21_X1 port map( A1 => n22762, A2 => n28314, B => n12726, ZN => 
                           n14680);
   U10869 : AOI21_X1 port map( A1 => n22698, A2 => n30960, B => n5689, ZN => 
                           n22699);
   U10953 : NAND2_X1 port map( A1 => n4805, A2 => n29648, ZN => n4804);
   U642 : NAND2_X1 port map( A1 => n28071, A2 => n22964, ZN => n3692);
   U13006 : NOR2_X1 port map( A1 => n28867, A2 => n985, ZN => n30168);
   U8698 : NOR2_X1 port map( A1 => n30488, A2 => n31455, ZN => n4174);
   U17761 : NAND2_X1 port map( A1 => n32088, A2 => n26526, ZN => n14769);
   U9446 : OAI21_X1 port map( A1 => n6149, A2 => n29325, B => n33382, ZN => 
                           n6148);
   U3266 : NOR2_X1 port map( A1 => n16142, A2 => n16236, ZN => n16993);
   U2589 : NOR2_X1 port map( A1 => n27798, A2 => n22986, ZN => n22864);
   U12020 : NAND2_X1 port map( A1 => n27090, A2 => n29967, ZN => n16514);
   U625 : CLKBUF_X2 port map( I => n31942, Z => n3999);
   U520 : INV_X1 port map( I => n5620, ZN => n5055);
   U2342 : NAND2_X1 port map( A1 => n23045, A2 => n22795, ZN => n15580);
   U10913 : NAND2_X1 port map( A1 => n7047, A2 => n5178, ZN => n5182);
   U17891 : OR2_X1 port map( A1 => n4599, A2 => n14540, Z => n14212);
   U5749 : OAI21_X1 port map( A1 => n26507, A2 => n22901, B => n15601, ZN => 
                           n18177);
   U9238 : NAND3_X1 port map( A1 => n802, A2 => n10031, A3 => n9293, ZN => 
                           n11108);
   U326 : OAI22_X1 port map( A1 => n12762, A2 => n32089, B1 => n22866, B2 => 
                           n1277, ZN => n4268);
   U9256 : NAND2_X1 port map( A1 => n22981, A2 => n2130, ZN => n2111);
   U6918 : NOR2_X1 port map( A1 => n30365, A2 => n28649, ZN => n3174);
   U16007 : NAND2_X1 port map( A1 => n4649, A2 => n990, ZN => n4650);
   U626 : OAI21_X1 port map( A1 => n29430, A2 => n29477, B => n27589, ZN => 
                           n7724);
   U9252 : NAND2_X1 port map( A1 => n8084, A2 => n26373, ZN => n7356);
   U640 : AOI22_X1 port map( A1 => n23064, A2 => n30437, B1 => n10643, B2 => 
                           n1275, ZN => n30080);
   U20254 : NAND3_X1 port map( A1 => n13916, A2 => n22914, A3 => n12071, ZN => 
                           n15341);
   U18113 : NOR2_X1 port map( A1 => n8149, A2 => n8150, ZN => n31394);
   U7777 : OAI21_X1 port map( A1 => n17639, A2 => n28948, B => n6236, ZN => 
                           n26274);
   U26320 : BUF_X2 port map( I => n15341, Z => n29190);
   U5620 : NAND2_X1 port map( A1 => n14623, A2 => n11873, ZN => n30741);
   U7776 : OAI21_X1 port map( A1 => n14192, A2 => n6236, B => n26274, ZN => 
                           n11162);
   U1273 : BUF_X2 port map( I => n23453, Z => n438);
   U15079 : INV_X1 port map( I => n30532, ZN => n23461);
   U22465 : INV_X1 port map( I => n23273, ZN => n23503);
   U3603 : INV_X1 port map( I => n23489, ZN => n13216);
   U4004 : INV_X1 port map( I => n17871, ZN => n23462);
   U19931 : NAND2_X1 port map( A1 => n29160, A2 => n1260, ZN => n3408);
   U16062 : NAND2_X1 port map( A1 => n26900, A2 => n27457, ZN => n30319);
   U5750 : CLKBUF_X2 port map( I => n6386, Z => n3739);
   U5049 : INV_X1 port map( I => n23439, ZN => n23413);
   U600 : INV_X1 port map( I => n13347, ZN => n27220);
   U589 : INV_X1 port map( I => n23936, ZN => n30949);
   U24264 : INV_X1 port map( I => n28611, ZN => n14297);
   U9219 : INV_X1 port map( I => n17812, ZN => n23951);
   U9678 : INV_X1 port map( I => n29704, ZN => n28069);
   U23439 : INV_X1 port map( I => n15917, ZN => n23578);
   U3607 : INV_X2 port map( I => n10213, ZN => n801);
   U11171 : INV_X1 port map( I => n23765, ZN => n29865);
   U5696 : INV_X1 port map( I => n30949, ZN => n17181);
   U4656 : CLKBUF_X2 port map( I => n13361, Z => n29185);
   U13110 : INV_X2 port map( I => n23735, ZN => n1489);
   U26258 : INV_X1 port map( I => n29139, ZN => n29271);
   U5596 : CLKBUF_X2 port map( I => n6474, Z => n31179);
   U10829 : BUF_X2 port map( I => n23886, Z => n17234);
   U17601 : INV_X1 port map( I => n9796, ZN => n10279);
   U2871 : INV_X2 port map( I => n23201, ZN => n4177);
   U21008 : INV_X1 port map( I => n28069, ZN => n8045);
   U14135 : INV_X1 port map( I => n3169, ZN => n8838);
   U14960 : INV_X1 port map( I => n23951, ZN => n14473);
   U19037 : INV_X1 port map( I => n16563, ZN => n23759);
   U4625 : OR2_X1 port map( A1 => n17285, A2 => n17352, Z => n23906);
   U25858 : INV_X1 port map( I => n28847, ZN => n548);
   U1857 : INV_X1 port map( I => n23586, ZN => n23910);
   U9217 : INV_X1 port map( I => n23754, ZN => n12433);
   U23116 : INV_X1 port map( I => n16961, ZN => n23945);
   U309 : INV_X1 port map( I => n29270, ZN => n979);
   U17142 : INV_X1 port map( I => n14255, ZN => n14164);
   U282 : INV_X1 port map( I => n23745, ZN => n11567);
   U19149 : INV_X2 port map( I => n16333, ZN => n8544);
   U5036 : AND2_X1 port map( A1 => n2450, A2 => n23706, Z => n2460);
   U3606 : INV_X1 port map( I => n499, ZN => n10217);
   U3536 : NOR3_X1 port map( A1 => n14473, A2 => n8217, A3 => n979, ZN => 
                           n16862);
   U23772 : AOI21_X1 port map( A1 => n981, A2 => n354, B => n11888, ZN => 
                           n17616);
   U19360 : NAND2_X1 port map( A1 => n10213, A2 => n23871, ZN => n23694);
   U6850 : NAND2_X1 port map( A1 => n2460, A2 => n23782, ZN => n9278);
   U21773 : NOR2_X1 port map( A1 => n10217, A2 => n756, ZN => n12094);
   U6894 : INV_X2 port map( I => n23786, ZN => n23903);
   U22127 : AOI21_X1 port map( A1 => n27678, A2 => n1257, B => n844, ZN => 
                           n31163);
   U1916 : INV_X1 port map( I => n23611, ZN => n769);
   U5610 : BUF_X2 port map( I => n9430, Z => n31890);
   U400 : INV_X2 port map( I => n6474, ZN => n28367);
   U16638 : NAND2_X1 port map( A1 => n23765, A2 => n23764, ZN => n23923);
   U5832 : CLKBUF_X2 port map( I => n23755, Z => n28222);
   U15327 : INV_X2 port map( I => n1099, ZN => n978);
   U4222 : BUF_X2 port map( I => n23764, Z => n28676);
   U273 : INV_X2 port map( I => n23756, ZN => n23749);
   U23685 : INV_X2 port map( I => n28266, ZN => n23891);
   U5332 : INV_X1 port map( I => n12974, ZN => n17872);
   U11142 : INV_X1 port map( I => n26641, ZN => n6394);
   U292 : INV_X1 port map( I => n23764, ZN => n16337);
   U16578 : NAND2_X1 port map( A1 => n5373, A2 => n299, ZN => n5372);
   U6176 : INV_X1 port map( I => n23755, ZN => n23726);
   U7341 : INV_X1 port map( I => n32711, ZN => n23897);
   U1464 : INV_X1 port map( I => n27, ZN => n23798);
   U15458 : INV_X1 port map( I => n31796, ZN => n1254);
   U4493 : INV_X1 port map( I => n17245, ZN => n7073);
   U561 : NOR2_X1 port map( A1 => n27678, A2 => n8655, ZN => n8654);
   U13176 : CLKBUF_X2 port map( I => n23742, Z => n30089);
   U3039 : NOR2_X1 port map( A1 => n31916, A2 => n29268, ZN => n7140);
   U464 : INV_X1 port map( I => n9172, ZN => n3687);
   U9596 : AOI21_X1 port map( A1 => n29240, A2 => n33337, B => n23841, ZN => 
                           n17950);
   U1595 : INV_X1 port map( I => n30282, ZN => n5163);
   U23877 : NOR2_X1 port map( A1 => n893, A2 => n30059, ZN => n23660);
   U6177 : NOR2_X1 port map( A1 => n23778, A2 => n8547, ZN => n15658);
   U13682 : NAND2_X1 port map( A1 => n7005, A2 => n23910, ZN => n1641);
   U6897 : OAI21_X1 port map( A1 => n980, A2 => n23885, B => n9278, ZN => n9277
                           );
   U6193 : NOR2_X1 port map( A1 => n23855, A2 => n4177, ZN => n2233);
   U8486 : NAND2_X1 port map( A1 => n2023, A2 => n23793, ZN => n23569);
   U366 : INV_X1 port map( I => n23753, ZN => n26397);
   U25144 : NAND2_X1 port map( A1 => n31938, A2 => n976, ZN => n22833);
   U386 : NAND2_X1 port map( A1 => n16343, A2 => n16496, ZN => n26185);
   U22389 : NAND2_X1 port map( A1 => n31435, A2 => n26114, ZN => n31209);
   U9389 : NOR2_X1 port map( A1 => n12722, A2 => n23611, ZN => n26465);
   U5031 : INV_X1 port map( I => n11708, ZN => n23811);
   U18430 : INV_X1 port map( I => n23877, ZN => n30621);
   U550 : BUF_X2 port map( I => n14974, Z => n28210);
   U15352 : NAND2_X1 port map( A1 => n5372, A2 => n27474, ZN => n4340);
   U19677 : NOR2_X1 port map( A1 => n4319, A2 => n11968, ZN => n17612);
   U253 : INV_X1 port map( I => n23672, ZN => n144);
   U6878 : OAI21_X1 port map( A1 => n11923, A2 => n23888, B => n6479, ZN => 
                           n11673);
   U488 : AOI21_X1 port map( A1 => n30295, A2 => n30296, B => n28676, ZN => 
                           n30294);
   U13380 : NOR2_X1 port map( A1 => n23704, A2 => n32308, ZN => n17922);
   U5714 : NOR2_X1 port map( A1 => n11050, A2 => n23708, ZN => n23880);
   U22780 : NOR2_X1 port map( A1 => n28266, A2 => n18133, ZN => n23895);
   U9156 : AOI21_X1 port map( A1 => n7073, A2 => n1256, B => n1253, ZN => n3371
                           );
   U20319 : NAND2_X1 port map( A1 => n29218, A2 => n10187, ZN => n23558);
   U484 : NOR2_X1 port map( A1 => n23891, A2 => n23892, ZN => n30527);
   U15323 : INV_X1 port map( I => n23578, ZN => n11096);
   U3038 : INV_X1 port map( I => n31916, ZN => n3481);
   U4242 : INV_X1 port map( I => n10279, ZN => n23787);
   U5608 : BUF_X2 port map( I => n17157, Z => n14973);
   U26617 : INV_X1 port map( I => n23765, ZN => n17087);
   U6862 : NAND2_X1 port map( A1 => n14325, A2 => n23806, ZN => n23805);
   U2778 : INV_X1 port map( I => n1098, ZN => n27615);
   U4793 : CLKBUF_X2 port map( I => n893, Z => n5357);
   U16972 : NAND2_X1 port map( A1 => n23600, A2 => n6247, ZN => n27369);
   U26172 : NAND2_X1 port map( A1 => n11673, A2 => n23841, ZN => n31690);
   U13770 : NAND2_X1 port map( A1 => n10213, A2 => n6474, ZN => n3401);
   U25334 : OAI21_X1 port map( A1 => n6414, A2 => n16238, B => n23906, ZN => 
                           n23707);
   U10760 : INV_X1 port map( I => n23805, ZN => n9900);
   U16717 : NOR2_X1 port map( A1 => n23895, A2 => n29068, ZN => n5555);
   U446 : NOR2_X1 port map( A1 => n28855, A2 => n3687, ZN => n9645);
   U6909 : OAI21_X1 port map( A1 => n12528, A2 => n23782, B => n11240, ZN => 
                           n12527);
   U25318 : NAND3_X1 port map( A1 => n23884, A2 => n756, A3 => n33936, ZN => 
                           n23635);
   U6890 : NOR2_X1 port map( A1 => n23953, A2 => n3481, ZN => n7383);
   U16991 : NAND2_X1 port map( A1 => n12658, A2 => n667, ZN => n30409);
   U449 : AOI22_X1 port map( A1 => n9002, A2 => n11621, B1 => n10753, B2 => 
                           n30359, ZN => n30169);
   U5297 : OAI21_X1 port map( A1 => n17750, A2 => n23773, B => n23778, ZN => 
                           n8719);
   U5702 : NOR2_X1 port map( A1 => n23866, A2 => n843, ZN => n24000);
   U19527 : NAND2_X1 port map( A1 => n31179, A2 => n23871, ZN => n28728);
   U16718 : NAND2_X1 port map( A1 => n32434, A2 => n28266, ZN => n5556);
   U6911 : OAI21_X1 port map( A1 => n23953, A2 => n31601, B => n29372, ZN => 
                           n23564);
   U25345 : NAND2_X1 port map( A1 => n23776, A2 => n8547, ZN => n23747);
   U13808 : AOI21_X1 port map( A1 => n3480, A2 => n16686, B => n23953, ZN => 
                           n28534);
   U24612 : INV_X1 port map( I => n14513, ZN => n31479);
   U6888 : NOR2_X1 port map( A1 => n29372, A2 => n4991, ZN => n26837);
   U415 : NAND2_X1 port map( A1 => n9382, A2 => n313, ZN => n27811);
   U25323 : NAND2_X1 port map( A1 => n23656, A2 => n23746, ZN => n23657);
   U420 : OAI21_X1 port map( A1 => n16969, A2 => n29474, B => n23741, ZN => 
                           n29795);
   U6905 : OAI21_X1 port map( A1 => n15659, A2 => n15658, B => n16271, ZN => 
                           n31058);
   U15194 : OAI21_X1 port map( A1 => n29269, A2 => n10993, B => n23681, ZN => 
                           n14124);
   U3500 : AOI22_X1 port map( A1 => n15272, A2 => n10143, B1 => n4319, B2 => 
                           n23638, ZN => n28850);
   U14941 : OAI21_X1 port map( A1 => n23947, A2 => n13308, B => n29294, ZN => 
                           n1528);
   U22047 : AOI21_X1 port map( A1 => n23493, A2 => n29240, B => n31158, ZN => 
                           n11492);
   U23589 : NAND2_X1 port map( A1 => n28503, A2 => n23654, ZN => n23658);
   U21432 : NAND2_X1 port map( A1 => n8836, A2 => n5357, ZN => n31082);
   U12619 : OAI21_X1 port map( A1 => n23697, A2 => n11943, B => n9772, ZN => 
                           n30028);
   U7816 : NOR2_X1 port map( A1 => n23896, A2 => n27615, ZN => n10480);
   U15428 : OR2_X1 port map( A1 => n23856, A2 => n25996, Z => n9214);
   U6854 : NAND2_X1 port map( A1 => n23704, A2 => n34008, ZN => n4539);
   U6861 : NAND3_X1 port map( A1 => n7073, A2 => n1253, A3 => n16677, ZN => 
                           n7074);
   U26068 : AOI21_X1 port map( A1 => n23593, A2 => n23891, B => n23892, ZN => 
                           n6723);
   U12616 : NAND2_X1 port map( A1 => n30028, A2 => n33924, ZN => n9770);
   U3263 : NOR2_X1 port map( A1 => n10019, A2 => n10020, ZN => n29699);
   U340 : NAND2_X1 port map( A1 => n1920, A2 => n31890, ZN => n14047);
   U24501 : NOR2_X1 port map( A1 => n28637, A2 => n16118, ZN => n4483);
   U4089 : NOR2_X1 port map( A1 => n12722, A2 => n769, ZN => n24331);
   U18096 : INV_X1 port map( I => n30505, ZN => n1090);
   U2017 : INV_X1 port map( I => n24315, ZN => n797);
   U5280 : INV_X2 port map( I => n24014, ZN => n974);
   U210 : INV_X1 port map( I => n12374, ZN => n1245);
   U15615 : NAND2_X1 port map( A1 => n24159, A2 => n29157, ZN => n9977);
   U3331 : BUF_X2 port map( I => n10226, Z => n9275);
   U21919 : INV_X1 port map( I => n12356, ZN => n23970);
   U8247 : NOR2_X1 port map( A1 => n3667, A2 => n29561, ZN => n5199);
   U14704 : INV_X2 port map( I => n3077, ZN => n3148);
   U283 : NAND2_X1 port map( A1 => n4655, A2 => n17261, ZN => n24228);
   U5877 : INV_X2 port map( I => n26387, ZN => n13343);
   U8802 : INV_X1 port map( I => n24207, ZN => n24157);
   U22219 : INV_X2 port map( I => n13175, ZN => n1244);
   U8767 : INV_X2 port map( I => n6713, ZN => n737);
   U6973 : INV_X2 port map( I => n7465, ZN => n793);
   U6834 : INV_X1 port map( I => n24164, ZN => n14840);
   U26170 : NOR2_X1 port map( A1 => n11503, A2 => n9616, ZN => n1550);
   U226 : INV_X1 port map( I => n4655, ZN => n16621);
   U201 : INV_X1 port map( I => n24087, ZN => n24139);
   U227 : INV_X2 port map( I => n13223, ZN => n24251);
   U197 : INV_X1 port map( I => n24141, ZN => n7203);
   U12982 : INV_X1 port map( I => n6555, ZN => n9146);
   U7907 : NAND2_X1 port map( A1 => n24052, A2 => n24053, ZN => n9976);
   U301 : INV_X1 port map( I => n24240, ZN => n29043);
   U200 : INV_X1 port map( I => n24218, ZN => n1240);
   U12733 : INV_X1 port map( I => n23748, ZN => n15096);
   U4781 : INV_X1 port map( I => n24180, ZN => n13260);
   U22429 : INV_X1 port map( I => n16215, ZN => n796);
   U13827 : NAND2_X1 port map( A1 => n33763, A2 => n24216, ZN => n5098);
   U3086 : INV_X1 port map( I => n3421, ZN => n24134);
   U1970 : INV_X1 port map( I => n6319, ZN => n24013);
   U3838 : NOR2_X1 port map( A1 => n24114, A2 => n24283, ZN => n23961);
   U21617 : NAND2_X1 port map( A1 => n16621, A2 => n28694, ZN => n17940);
   U220 : INV_X1 port map( I => n16868, ZN => n972);
   U11016 : NOR2_X1 port map( A1 => n27104, A2 => n3077, ZN => n29848);
   U6940 : NOR2_X1 port map( A1 => n30289, A2 => n15068, ZN => n31071);
   U17734 : NAND2_X1 port map( A1 => n7546, A2 => n24221, ZN => n11535);
   U2068 : NAND2_X1 port map( A1 => n6003, A2 => n12356, ZN => n5437);
   U9138 : NAND2_X1 port map( A1 => n32917, A2 => n23970, ZN => n26674);
   U4111 : BUF_X2 port map( I => n5199, Z => n29141);
   U6114 : NAND2_X1 port map( A1 => n9323, A2 => n8178, ZN => n2247);
   U14628 : INV_X1 port map( I => n33832, ZN => n14542);
   U1757 : BUF_X2 port map( I => n3718, Z => n8);
   U4215 : CLKBUF_X2 port map( I => n17426, Z => n8165);
   U9102 : NAND2_X1 port map( A1 => n24052, A2 => n24185, ZN => n24123);
   U14723 : INV_X2 port map( I => n24052, ZN => n11463);
   U271 : INV_X1 port map( I => n29307, ZN => n24272);
   U6951 : NAND2_X1 port map( A1 => n24230, A2 => n31355, ZN => n14861);
   U2802 : INV_X1 port map( I => n14195, ZN => n14443);
   U18877 : INV_X1 port map( I => n2558, ZN => n7150);
   U6108 : NOR2_X1 port map( A1 => n2744, A2 => n31377, ZN => n13170);
   U374 : INV_X1 port map( I => n1808, ZN => n24237);
   U10162 : INV_X1 port map( I => n29157, ZN => n29748);
   U2784 : INV_X1 port map( I => n9616, ZN => n5308);
   U13027 : OAI21_X1 port map( A1 => n4118, A2 => n4775, B => n24134, ZN => 
                           n17860);
   U193 : NAND2_X1 port map( A1 => n10188, A2 => n13260, ZN => n17943);
   U25398 : NAND3_X1 port map( A1 => n24118, A2 => n24223, A3 => n24225, ZN => 
                           n24119);
   U15765 : NAND2_X1 port map( A1 => n792, A2 => n27104, ZN => n2798);
   U17015 : NAND2_X1 port map( A1 => n27661, A2 => n1240, ZN => n6251);
   U18960 : NOR2_X1 port map( A1 => n24092, A2 => n31096, ZN => n30696);
   U10574 : NAND2_X1 port map( A1 => n26027, A2 => n4024, ZN => n3217);
   U2115 : NOR2_X1 port map( A1 => n24292, A2 => n32936, ZN => n24294);
   U9057 : INV_X1 port map( I => n13378, ZN => n3603);
   U12857 : NOR2_X1 port map( A1 => n891, A2 => n33597, ZN => n23962);
   U1991 : INV_X1 port map( I => n24005, ZN => n3903);
   U2446 : NOR2_X1 port map( A1 => n32917, A2 => n17404, ZN => n23701);
   U152 : INV_X1 port map( I => n24206, ZN => n24009);
   U11014 : OAI21_X1 port map( A1 => n10938, A2 => n29848, B => n24268, ZN => 
                           n31297);
   U21830 : NAND2_X1 port map( A1 => n5631, A2 => n12143, ZN => n24297);
   U15608 : INV_X1 port map( I => n24159, ZN => n24124);
   U20738 : NAND2_X1 port map( A1 => n9892, A2 => n14336, ZN => n31868);
   U327 : NOR2_X1 port map( A1 => n12862, A2 => n27661, ZN => n27334);
   U9711 : NAND2_X1 port map( A1 => n7779, A2 => n10104, ZN => n28351);
   U3078 : NAND3_X1 port map( A1 => n24027, A2 => n28040, A3 => n31002, ZN => 
                           n24029);
   U15567 : NOR2_X1 port map( A1 => n27436, A2 => n6476, ZN => n11950);
   U5259 : OR2_X1 port map( A1 => n11535, A2 => n3506, Z => n11534);
   U5474 : NAND2_X1 port map( A1 => n24182, A2 => n31722, ZN => n17100);
   U10590 : NOR2_X1 port map( A1 => n17232, A2 => n3506, ZN => n17016);
   U13737 : NAND2_X1 port map( A1 => n26459, A2 => n24093, ZN => n29123);
   U3611 : INV_X1 port map( I => n24270, ZN => n11721);
   U9040 : OAI22_X1 port map( A1 => n7149, A2 => n15179, B1 => n14399, B2 => 
                           n29120, ZN => n6877);
   U10554 : AOI21_X1 port map( A1 => n11997, A2 => n12576, B => n28040, ZN => 
                           n10667);
   U288 : NAND2_X1 port map( A1 => n30348, A2 => n24313, ZN => n7483);
   U15675 : NAND2_X1 port map( A1 => n14861, A2 => n11743, ZN => n11742);
   U17877 : NAND2_X1 port map( A1 => n27550, A2 => n32465, ZN => n14724);
   U18410 : NAND3_X1 port map( A1 => n24091, A2 => n16535, A3 => n24234, ZN => 
                           n24655);
   U9621 : NAND2_X1 port map( A1 => n24052, A2 => n24159, ZN => n24183);
   U20110 : NAND2_X1 port map( A1 => n33763, A2 => n31497, ZN => n24109);
   U6146 : INV_X1 port map( I => n24220, ZN => n1094);
   U9079 : NAND2_X1 port map( A1 => n11463, A2 => n24053, ZN => n30726);
   U155 : INV_X1 port map( I => n24216, ZN => n24290);
   U13048 : INV_X1 port map( I => n11883, ZN => n24233);
   U7357 : AND2_X1 port map( A1 => n4286, A2 => n16052, Z => n29473);
   U214 : INV_X1 port map( I => n28827, ZN => n3219);
   U308 : NAND2_X1 port map( A1 => n28300, A2 => n891, ZN => n16683);
   U19081 : NOR2_X1 port map( A1 => n3506, A2 => n7546, ZN => n30715);
   U7798 : NAND3_X1 port map( A1 => n24185, A2 => n11463, A3 => n1088, ZN => 
                           n11461);
   U1551 : NOR2_X1 port map( A1 => n24118, A2 => n10118, ZN => n10117);
   U7771 : NAND3_X1 port map( A1 => n2847, A2 => n24163, A3 => n24002, ZN => 
                           n23988);
   U20755 : NAND2_X1 port map( A1 => n23995, A2 => n24270, ZN => n24385);
   U189 : NAND3_X1 port map( A1 => n6001, A2 => n26516, A3 => n17404, ZN => 
                           n17493);
   U19785 : OAI21_X1 port map( A1 => n31113, A2 => n24290, B => n11613, ZN => 
                           n30826);
   U5001 : NAND3_X1 port map( A1 => n33597, A2 => n7546, A3 => n24286, ZN => 
                           n5307);
   U18351 : NAND2_X1 port map( A1 => n24046, A2 => n13950, ZN => n17233);
   U23100 : NAND2_X1 port map( A1 => n24249, A2 => n24248, ZN => n15085);
   U284 : NAND2_X1 port map( A1 => n16683, A2 => n28409, ZN => n30417);
   U4996 : NOR3_X1 port map( A1 => n24202, A2 => n738, A3 => n27501, ZN => 
                           n12262);
   U8664 : AOI21_X1 port map( A1 => n31679, A2 => n23748, B => n1499, ZN => 
                           n1497);
   U10635 : NAND2_X1 port map( A1 => n24273, A2 => n31918, ZN => n11724);
   U19113 : NOR2_X1 port map( A1 => n30726, A2 => n1088, ZN => n26307);
   U10571 : OAI21_X1 port map( A1 => n11950, A2 => n3632, B => n28296, ZN => 
                           n3631);
   U291 : NOR2_X1 port map( A1 => n24107, A2 => n891, ZN => n30096);
   U9904 : NAND3_X1 port map( A1 => n2865, A2 => n27786, A3 => n31096, ZN => 
                           n2186);
   U5439 : NAND2_X1 port map( A1 => n31544, A2 => n31543, ZN => n9367);
   U6109 : AOI21_X1 port map( A1 => n12693, A2 => n12692, B => n32917, ZN => 
                           n12691);
   U15924 : NAND2_X1 port map( A1 => n8142, A2 => n5490, ZN => n24017);
   U18278 : AOI21_X1 port map( A1 => n31002, A2 => n12982, B => n28040, ZN => 
                           n30598);
   U11543 : NAND2_X1 port map( A1 => n5631, A2 => n24292, ZN => n12429);
   U5164 : INV_X1 port map( I => n12868, ZN => n2424);
   U13150 : NAND4_X1 port map( A1 => n24343, A2 => n24342, A3 => n24344, A4 => 
                           n24341, ZN => n31311);
   U143 : NOR2_X1 port map( A1 => n28590, A2 => n9066, ZN => n11042);
   U279 : NAND2_X1 port map( A1 => n14445, A2 => n14444, ZN => n31788);
   U3234 : BUF_X2 port map( I => n7679, Z => n356);
   U18973 : CLKBUF_X2 port map( I => n24544, Z => n27733);
   U1275 : INV_X2 port map( I => n5970, ZN => n9907);
   U10527 : INV_X1 port map( I => n24393, ZN => n8703);
   U5162 : BUF_X2 port map( I => n12868, Z => n28977);
   U13673 : NOR2_X1 port map( A1 => n16815, A2 => n26966, ZN => n3295);
   U2483 : INV_X1 port map( I => n24805, ZN => n14533);
   U4747 : NAND2_X1 port map( A1 => n2421, A2 => n2420, ZN => n17682);
   U5418 : CLKBUF_X2 port map( I => n24843, Z => n10870);
   U21378 : INV_X1 port map( I => n28119, ZN => n4886);
   U4984 : INV_X1 port map( I => n679, ZN => n25397);
   U19889 : INV_X1 port map( I => n9932, ZN => n10062);
   U12755 : INV_X1 port map( I => n25707, ZN => n31570);
   U2814 : INV_X1 port map( I => n25394, ZN => n13993);
   U15333 : BUF_X2 port map( I => n23668, Z => n25871);
   U5247 : INV_X2 port map( I => n16957, ZN => n9917);
   U112 : INV_X1 port map( I => n25536, ZN => n833);
   U14756 : BUF_X2 port map( I => n25111, Z => n25234);
   U8982 : INV_X1 port map( I => n25238, ZN => n6910);
   U115 : INV_X1 port map( I => n5020, ZN => n11987);
   U14347 : INV_X1 port map( I => n27072, ZN => n17655);
   U5957 : INV_X1 port map( I => n25699, ZN => n751);
   U22211 : INV_X1 port map( I => n24360, ZN => n13042);
   U235 : INV_X1 port map( I => n680, ZN => n24973);
   U88 : INV_X1 port map( I => n17240, ZN => n885);
   U2134 : INV_X2 port map( I => n17655, ZN => n25633);
   U5956 : NAND2_X1 port map( A1 => n25867, A2 => n14111, ZN => n10549);
   U2638 : INV_X1 port map( I => n10199, ZN => n17839);
   U5601 : INV_X2 port map( I => n8219, ZN => n1216);
   U20653 : NAND2_X1 port map( A1 => n1567, A2 => n2092, ZN => n30948);
   U4981 : INV_X1 port map( I => n15777, ZN => n25870);
   U4056 : INV_X1 port map( I => n13993, ZN => n11704);
   U2860 : NAND2_X1 port map( A1 => n16632, A2 => n1786, ZN => n27479);
   U128 : INV_X1 port map( I => n25766, ZN => n27359);
   U2509 : CLKBUF_X2 port map( I => n25699, Z => n28242);
   U6777 : INV_X1 port map( I => n15719, ZN => n24983);
   U8968 : NAND2_X1 port map( A1 => n11945, A2 => n15046, ZN => n24609);
   U188 : NOR2_X1 port map( A1 => n24361, A2 => n17118, ZN => n30907);
   U2813 : BUF_X2 port map( I => n18156, Z => n5202);
   U5612 : INV_X2 port map( I => n17963, ZN => n25901);
   U106 : INV_X2 port map( I => n29629, ZN => n14055);
   U25721 : INV_X1 port map( I => n25763, ZN => n25704);
   U80 : INV_X1 port map( I => n11957, ZN => n754);
   U14968 : INV_X1 port map( I => n18242, ZN => n836);
   U190 : NAND2_X1 port map( A1 => n25977, A2 => n11947, ZN => n25239);
   U13661 : INV_X1 port map( I => n8892, ZN => n25587);
   U19564 : INV_X1 port map( I => n28591, ZN => n13709);
   U3522 : INV_X1 port map( I => n29334, ZN => n8758);
   U23355 : INV_X1 port map( I => n14111, ZN => n16835);
   U2427 : INV_X1 port map( I => n29279, ZN => n717);
   U91 : INV_X2 port map( I => n25561, ZN => n15880);
   U4064 : INV_X1 port map( I => n25885, ZN => n884);
   U9001 : INV_X1 port map( I => n25760, ZN => n1080);
   U14842 : NAND2_X1 port map( A1 => n25013, A2 => n14020, ZN => n4814);
   U8487 : OAI21_X1 port map( A1 => n1221, A2 => n7689, B => n25892, ZN => 
                           n29594);
   U13398 : NAND2_X1 port map( A1 => n27651, A2 => n25019, ZN => n9402);
   U2010 : NOR2_X1 port map( A1 => n25636, A2 => n25713, ZN => n25639);
   U109 : NOR2_X1 port map( A1 => n7413, A2 => n25900, ZN => n10550);
   U15038 : OAI21_X1 port map( A1 => n16528, A2 => n25412, B => n419, ZN => 
                           n28279);
   U11003 : NAND3_X1 port map( A1 => n4968, A2 => n4967, A3 => n18264, ZN => 
                           n29846);
   U2004 : NOR2_X1 port map( A1 => n16850, A2 => n16957, ZN => n26873);
   U16046 : NAND2_X1 port map( A1 => n25398, A2 => n25397, ZN => n25399);
   U3747 : OAI21_X1 port map( A1 => n25900, A2 => n16835, B => n790, ZN => 
                           n15672);
   U16628 : NAND2_X1 port map( A1 => n25205, A2 => n27376, ZN => n27332);
   U4733 : NOR2_X1 port map( A1 => n9127, A2 => n16113, ZN => n11022);
   U15520 : INV_X1 port map( I => n5050, ZN => n7317);
   U20084 : NOR2_X1 port map( A1 => n31268, A2 => n25977, ZN => n10314);
   U15439 : NAND2_X1 port map( A1 => n17987, A2 => n25145, ZN => n25184);
   U162 : INV_X1 port map( I => n32760, ZN => n24873);
   U10450 : NAND2_X1 port map( A1 => n3013, A2 => n28815, ZN => n24877);
   U23913 : NAND2_X1 port map( A1 => n11716, A2 => n4993, ZN => n24310);
   U26494 : NAND2_X1 port map( A1 => n25133, A2 => n31779, ZN => n31778);
   U20372 : NOR2_X1 port map( A1 => n17839, A2 => n30907, ZN => n5115);
   U3301 : NOR2_X1 port map( A1 => n25620, A2 => n25708, ZN => n15354);
   U2290 : NOR2_X1 port map( A1 => n13464, A2 => n9862, ZN => n12522);
   U25606 : INV_X1 port map( I => n25339, ZN => n25337);
   U3293 : NAND2_X1 port map( A1 => n15255, A2 => n31945, ZN => n25531);
   U4433 : INV_X1 port map( I => n6939, ZN => n1082);
   U10875 : INV_X1 port map( I => n7350, ZN => n6850);
   U6999 : INV_X1 port map( I => n12247, ZN => n11106);
   U7729 : INV_X1 port map( I => n25587, ZN => n25388);
   U7022 : INV_X1 port map( I => n25229, ZN => n1215);
   U25885 : NOR2_X1 port map( A1 => n25562, A2 => n16783, ZN => n28866);
   U2371 : NOR2_X1 port map( A1 => n15964, A2 => n25531, ZN => n24633);
   U10436 : NOR2_X1 port map( A1 => n15646, A2 => n27314, ZN => n2999);
   U78 : NAND3_X1 port map( A1 => n29976, A2 => n25183, A3 => n1218, ZN => 
                           n14632);
   U13514 : NAND2_X1 port map( A1 => n16609, A2 => n755, ZN => n24430);
   U2852 : OAI21_X1 port map( A1 => n25199, A2 => n1786, B => n16632, ZN => 
                           n27990);
   U11238 : NOR2_X1 port map( A1 => n5791, A2 => n5793, ZN => n5570);
   U20208 : NAND2_X1 port map( A1 => n5387, A2 => n13349, ZN => n4232);
   U4016 : NAND2_X1 port map( A1 => n28564, A2 => n28562, ZN => n15883);
   U10297 : AOI21_X1 port map( A1 => n146, A2 => n9363, B => n7064, ZN => 
                           n25767);
   U2333 : NAND2_X1 port map( A1 => n25396, A2 => n11556, ZN => n25439);
   U114 : NAND2_X1 port map( A1 => n15550, A2 => n4318, ZN => n2182);
   U75 : NOR2_X1 port map( A1 => n689, A2 => n15013, ZN => n14539);
   U13045 : NOR2_X1 port map( A1 => n15785, A2 => n26873, ZN => n15783);
   U4386 : NOR2_X1 port map( A1 => n10550, A2 => n8470, ZN => n10547);
   U2745 : OAI22_X1 port map( A1 => n2456, A2 => n25234, B1 => n25235, B2 => 
                           n25187, ZN => n24570);
   U17416 : NAND2_X1 port map( A1 => n25523, A2 => n25522, ZN => n8442);
   U67 : OAI21_X1 port map( A1 => n25896, A2 => n16113, B => n13349, ZN => 
                           n24708);
   U15626 : NAND3_X1 port map( A1 => n17673, A2 => n14247, A3 => n25404, ZN => 
                           n25441);
   U9087 : AOI21_X1 port map( A1 => n11306, A2 => n25633, B => n27637, ZN => 
                           n12000);
   U10381 : OAI21_X1 port map( A1 => n12025, A2 => n17367, B => n25388, ZN => 
                           n11823);
   U23903 : AOI21_X1 port map( A1 => n24604, A2 => n15719, B => n27314, ZN => 
                           n17379);
   U6028 : OAI22_X1 port map( A1 => n8186, A2 => n11944, B1 => n17092, B2 => 
                           n6939, ZN => n15276);
   U10372 : NOR2_X1 port map( A1 => n4095, A2 => n7041, ZN => n11698);
   U10428 : NAND2_X1 port map( A1 => n12058, A2 => n16752, ZN => n11347);
   U2719 : AOI21_X1 port map( A1 => n14484, A2 => n32761, B => n11082, ZN => 
                           n11429);
   U12511 : NAND2_X1 port map( A1 => n1620, A2 => n25887, ZN => n25914);
   U7030 : INV_X1 port map( I => n2270, ZN => n15061);
   U8008 : INV_X1 port map( I => n10174, ZN => n10504);
   U15219 : INV_X1 port map( I => n25376, ZN => n25352);
   U9998 : INV_X2 port map( I => n1597, ZN => n25738);
   U14917 : NAND2_X1 port map( A1 => n25107, A2 => n11360, ZN => n7862);
   U4928 : INV_X1 port map( I => n25478, ZN => n25487);
   U2934 : CLKBUF_X2 port map( I => n7702, Z => n7701);
   U14791 : INV_X1 port map( I => n25795, ZN => n16111);
   U57 : NAND2_X1 port map( A1 => n16494, A2 => n13640, ZN => n13124);
   U17512 : INV_X2 port map( I => n16380, ZN => n1951);
   U1540 : INV_X1 port map( I => n25154, ZN => n25179);
   U10377 : INV_X1 port map( I => n25369, ZN => n25367);
   U24431 : INV_X1 port map( I => n14915, ZN => n25834);
   U8903 : OAI21_X1 port map( A1 => n3489, A2 => n2536, B => n32059, ZN => 
                           n8951);
   U1905 : NOR2_X1 port map( A1 => n30279, A2 => n25002, ZN => n15078);
   U15859 : NAND2_X1 port map( A1 => n25687, A2 => n25686, ZN => n2016);
   U7032 : NOR2_X1 port map( A1 => n5411, A2 => n7701, ZN => n14434);
   U23575 : INV_X1 port map( I => n31360, ZN => n25552);
   U13124 : NOR2_X1 port map( A1 => n14199, A2 => n25863, ZN => n13952);
   U15732 : NAND2_X1 port map( A1 => n8202, A2 => n4525, ZN => n4524);
   U21482 : INV_X1 port map( I => n25464, ZN => n17200);
   U4329 : CLKBUF_X1 port map( I => n25557, Z => n31647);
   U25689 : NAND2_X1 port map( A1 => n29116, A2 => n25476, ZN => n25474);
   U10322 : INV_X1 port map( I => n25738, ZN => n25748);
   U5548 : INV_X1 port map( I => n25863, ZN => n25854);
   U19 : INV_X1 port map( I => n24915, ZN => n6154);
   U7051 : INV_X1 port map( I => n25724, ZN => n25729);
   U3985 : INV_X1 port map( I => n13483, ZN => n14944);
   U4 : NAND4_X1 port map( A1 => n25914, A2 => n25922, A3 => n11019, A4 => 
                           n25913, ZN => n25918);
   U10329 : NAND2_X1 port map( A1 => n24351, A2 => n24927, ZN => n24349);
   U3 : NAND3_X1 port map( A1 => n25318, A2 => n17058, A3 => n17105, ZN => 
                           n27063);
   U7 : NOR2_X1 port map( A1 => n8639, A2 => n32398, ZN => n32270);
   U16 : INV_X1 port map( I => n13960, ZN => n25925);
   U17 : INV_X1 port map( I => n25106, ZN => n32857);
   U18 : BUF_X2 port map( I => n25820, Z => n11003);
   U20 : NOR2_X1 port map( A1 => n16112, A2 => n12611, ZN => n12395);
   U21 : NOR2_X1 port map( A1 => n25788, A2 => n25796, ZN => n25775);
   U22 : NAND2_X1 port map( A1 => n7586, A2 => n11360, ZN => n25093);
   U25 : NAND2_X1 port map( A1 => n24925, A2 => n15799, ZN => n24928);
   U26 : NAND2_X1 port map( A1 => n34109, A2 => n25247, ZN => n7924);
   U27 : AND2_X1 port map( A1 => n25387, A2 => n33876, Z => n32869);
   U28 : INV_X1 port map( I => n15323, ZN => n712);
   U29 : BUF_X2 port map( I => n5578, Z => n5043);
   U30 : INV_X1 port map( I => n24910, ZN => n24902);
   U31 : AOI21_X1 port map( A1 => n5810, A2 => n8186, B => n32992, ZN => n25731
                           );
   U32 : CLKBUF_X2 port map( I => n25285, Z => n28532);
   U33 : INV_X1 port map( I => n6595, ZN => n33399);
   U37 : INV_X1 port map( I => n24955, ZN => n1201);
   U38 : INV_X1 port map( I => n25820, ZN => n17642);
   U40 : NAND2_X1 port map( A1 => n32882, A2 => n10609, ZN => n33900);
   U42 : NOR2_X1 port map( A1 => n25818, A2 => n4450, ZN => n9182);
   U51 : OAI21_X2 port map( A1 => n32471, A2 => n32565, B => n25010, ZN => 
                           n25062);
   U55 : OR2_X1 port map( A1 => n24572, A2 => n24570, Z => n32882);
   U56 : INV_X1 port map( I => n24995, ZN => n5072);
   U59 : NAND2_X1 port map( A1 => n33632, A2 => n12968, ZN => n25845);
   U60 : NOR2_X1 port map( A1 => n32030, A2 => n14872, ZN => n32311);
   U61 : NAND3_X1 port map( A1 => n15051, A2 => n5659, A3 => n5755, ZN => 
                           n30928);
   U65 : AOI21_X1 port map( A1 => n25564, A2 => n3405, B => n25582, ZN => 
                           n32585);
   U66 : NAND2_X1 port map( A1 => n32570, A2 => n5292, ZN => n32135);
   U70 : AND2_X1 port map( A1 => n13985, A2 => n25306, Z => n32020);
   U72 : NOR2_X1 port map( A1 => n33074, A2 => n16566, ZN => n32626);
   U73 : NAND3_X1 port map( A1 => n27119, A2 => n16339, A3 => n25412, ZN => 
                           n33245);
   U76 : NAND2_X1 port map( A1 => n33599, A2 => n33598, ZN => n33632);
   U77 : CLKBUF_X2 port map( I => n7532, Z => n31946);
   U81 : NAND2_X1 port map( A1 => n6851, A2 => n12440, ZN => n2000);
   U82 : NAND2_X1 port map( A1 => n32828, A2 => n32761, ZN => n8776);
   U83 : NAND2_X1 port map( A1 => n11703, A2 => n25347, ZN => n30930);
   U85 : OAI21_X1 port map( A1 => n30372, A2 => n25329, B => n28958, ZN => 
                           n33880);
   U86 : OAI21_X1 port map( A1 => n14991, A2 => n12093, B => n30461, ZN => 
                           n32205);
   U87 : OAI21_X1 port map( A1 => n15555, A2 => n25893, B => n9127, ZN => 
                           n11020);
   U89 : AOI21_X1 port map( A1 => n25711, A2 => n24729, B => n4407, ZN => 
                           n27208);
   U92 : NOR2_X1 port map( A1 => n16783, A2 => n25561, ZN => n30983);
   U93 : NOR2_X1 port map( A1 => n1221, A2 => n547, ZN => n12160);
   U95 : NAND2_X1 port map( A1 => n25755, A2 => n28338, ZN => n25876);
   U97 : OR2_X1 port map( A1 => n28242, A2 => n25627, Z => n32032);
   U98 : AND2_X1 port map( A1 => n17240, A2 => n25012, Z => n11977);
   U99 : CLKBUF_X2 port map( I => n25582, Z => n27947);
   U102 : NAND2_X1 port map( A1 => n28110, A2 => n1211, ZN => n33002);
   U104 : NOR2_X1 port map( A1 => n765, A2 => n25331, ZN => n30522);
   U108 : AND2_X1 port map( A1 => n9195, A2 => n25700, Z => n32028);
   U110 : OR2_X1 port map( A1 => n317, A2 => n16783, Z => n32029);
   U113 : INV_X1 port map( I => n32878, ZN => n32761);
   U116 : AND2_X1 port map( A1 => n17240, A2 => n25014, Z => n14991);
   U120 : OR2_X1 port map( A1 => n24667, A2 => n16957, Z => n33962);
   U125 : INV_X1 port map( I => n33067, ZN => n33066);
   U126 : NAND2_X1 port map( A1 => n16276, A2 => n25183, ZN => n14630);
   U140 : NAND2_X1 port map( A1 => n16751, A2 => n17987, ZN => n14629);
   U142 : NOR2_X1 port map( A1 => n1567, A2 => n25121, ZN => n7771);
   U144 : NAND2_X1 port map( A1 => n25891, A2 => n25890, ZN => n30811);
   U146 : INV_X2 port map( I => n11045, ZN => n25902);
   U148 : BUF_X2 port map( I => n25883, Z => n15152);
   U149 : INV_X2 port map( I => n25409, ZN => n752);
   U154 : NOR2_X1 port map( A1 => n28338, A2 => n25755, ZN => n28110);
   U157 : NAND2_X1 port map( A1 => n25014, A2 => n11974, ZN => n24977);
   U160 : OR2_X1 port map( A1 => n10569, A2 => n4951, Z => n25289);
   U161 : INV_X1 port map( I => n31945, ZN => n16648);
   U165 : AOI21_X1 port map( A1 => n15459, A2 => n25697, B => n751, ZN => 
                           n15458);
   U169 : BUF_X2 port map( I => n25238, Z => n28136);
   U172 : CLKBUF_X2 port map( I => n17382, Z => n27314);
   U174 : CLKBUF_X1 port map( I => n25334, Z => n33460);
   U177 : CLKBUF_X1 port map( I => n16510, Z => n32884);
   U178 : AOI21_X1 port map( A1 => n31149, A2 => n16704, B => n25561, ZN => 
                           n33067);
   U179 : BUF_X2 port map( I => n25563, Z => n317);
   U180 : CLKBUF_X2 port map( I => n24436, Z => n33120);
   U183 : OR2_X1 port map( A1 => n6725, A2 => n27181, Z => n25584);
   U185 : NAND2_X1 port map( A1 => n25295, A2 => n16650, ZN => n25343);
   U187 : INV_X1 port map( I => n10569, ZN => n5468);
   U191 : BUF_X2 port map( I => n25022, Z => n25121);
   U199 : BUF_X2 port map( I => n14246, Z => n33919);
   U202 : INV_X1 port map( I => n24692, ZN => n14110);
   U215 : INV_X1 port map( I => n24547, ZN => n32575);
   U216 : BUF_X2 port map( I => n3253, Z => n30069);
   U217 : INV_X1 port map( I => n27115, ZN => n32346);
   U219 : OAI22_X1 port map( A1 => n17581, A2 => n3219, B1 => n15086, B2 => 
                           n15085, ZN => n32871);
   U221 : AOI21_X1 port map( A1 => n32470, A2 => n28827, B => n25974, ZN => 
                           n13217);
   U222 : NAND2_X1 port map( A1 => n891, A2 => n33935, ZN => n27397);
   U228 : NAND2_X1 port map( A1 => n33123, A2 => n6978, ZN => n6167);
   U229 : NAND3_X1 port map( A1 => n16651, A2 => n30061, A3 => n29977, ZN => 
                           n7729);
   U233 : AOI22_X1 port map( A1 => n2853, A2 => n24163, B1 => n24002, B2 => 
                           n16552, ZN => n2848);
   U234 : OAI21_X1 port map( A1 => n13659, A2 => n29473, B => n9219, ZN => 
                           n29605);
   U238 : AOI21_X1 port map( A1 => n24268, A2 => n11768, B => n12644, ZN => 
                           n11767);
   U239 : OAI22_X1 port map( A1 => n24235, A2 => n24237, B1 => n11883, B2 => 
                           n24234, ZN => n24239);
   U242 : AOI21_X1 port map( A1 => n7150, A2 => n15179, B => n9889, ZN => 
                           n12341);
   U243 : INV_X1 port map( I => n32444, ZN => n13659);
   U244 : NAND2_X1 port map( A1 => n24052, A2 => n14123, ZN => n24125);
   U247 : NAND2_X1 port map( A1 => n14386, A2 => n7962, ZN => n33951);
   U249 : NAND2_X1 port map( A1 => n5132, A2 => n32228, ZN => n5130);
   U252 : NAND3_X1 port map( A1 => n890, A2 => n29141, A3 => n7361, ZN => n7360
                           );
   U255 : OR2_X1 port map( A1 => n29634, A2 => n12374, Z => n12054);
   U256 : CLKBUF_X1 port map( I => n10987, Z => n28538);
   U257 : OAI21_X1 port map( A1 => n32552, A2 => n32551, B => n24213, ZN => 
                           n24007);
   U260 : NAND2_X1 port map( A1 => n10687, A2 => n13, ZN => n13974);
   U263 : NAND2_X1 port map( A1 => n24337, A2 => n33680, ZN => n1998);
   U266 : NOR2_X1 port map( A1 => n28300, A2 => n31985, ZN => n6105);
   U269 : NAND2_X1 port map( A1 => n24318, A2 => n2913, ZN => n26488);
   U270 : AOI21_X1 port map( A1 => n9946, A2 => n27931, B => n4019, ZN => n5708
                           );
   U272 : NAND2_X1 port map( A1 => n31377, A2 => n24317, ZN => n32166);
   U275 : NAND2_X1 port map( A1 => n24143, A2 => n27430, ZN => n33653);
   U280 : NOR2_X1 port map( A1 => n31355, A2 => n28694, ZN => n33872);
   U286 : OR2_X1 port map( A1 => n24141, A2 => n24084, Z => n16017);
   U293 : AOI22_X1 port map( A1 => n32062, A2 => n27739, B1 => n24133, B2 => 
                           n23714, ZN => n2939);
   U296 : NAND3_X1 port map( A1 => n32298, A2 => n14112, A3 => n2913, ZN => 
                           n33912);
   U298 : AOI21_X1 port map( A1 => n28410, A2 => n5308, B => n3506, ZN => 
                           n28409);
   U300 : NAND3_X1 port map( A1 => n9066, A2 => n12982, A3 => n27739, ZN => 
                           n16950);
   U305 : NAND2_X1 port map( A1 => n24161, A2 => n24123, ZN => n5969);
   U306 : NAND2_X1 port map( A1 => n31342, A2 => n24249, ZN => n32470);
   U307 : INV_X2 port map( I => n15179, ZN => n15876);
   U310 : NAND2_X1 port map( A1 => n24340, A2 => n24056, ZN => n4049);
   U314 : NOR2_X1 port map( A1 => n24309, A2 => n3421, ZN => n24135);
   U315 : INV_X1 port map( I => n24248, ZN => n31342);
   U321 : INV_X2 port map( I => n12143, ZN => n33444);
   U331 : BUF_X2 port map( I => n24164, Z => n2847);
   U333 : NAND3_X1 port map( A1 => n13984, A2 => n5913, A3 => n31096, ZN => 
                           n11743);
   U334 : AND2_X1 port map( A1 => n2539, A2 => n11503, Z => n31985);
   U336 : NAND2_X1 port map( A1 => n31497, A2 => n10530, ZN => n2529);
   U337 : OR2_X1 port map( A1 => n24254, A2 => n33532, Z => n7149);
   U338 : INV_X1 port map( I => n27430, ZN => n33655);
   U341 : NOR2_X1 port map( A1 => n24209, A2 => n24212, ZN => n32551);
   U343 : NAND2_X1 port map( A1 => n12644, A2 => n3148, ZN => n4961);
   U344 : NOR2_X1 port map( A1 => n24347, A2 => n3165, ZN => n30121);
   U346 : NAND2_X1 port map( A1 => n13334, A2 => n6713, ZN => n1500);
   U347 : INV_X2 port map( I => n26120, ZN => n2640);
   U349 : INV_X1 port map( I => n24053, ZN => n24185);
   U350 : INV_X2 port map( I => n2826, ZN => n24340);
   U351 : BUF_X2 port map( I => n6555, Z => n6581);
   U354 : OAI21_X1 port map( A1 => n24225, A2 => n10687, B => n24223, ZN => 
                           n32677);
   U358 : NAND2_X1 port map( A1 => n7991, A2 => n26415, ZN => n23997);
   U362 : NAND2_X1 port map( A1 => n4024, A2 => n24312, ZN => n29051);
   U364 : INV_X1 port map( I => n15720, ZN => n14703);
   U365 : NAND3_X1 port map( A1 => n15943, A2 => n23903, A3 => n15942, ZN => 
                           n29575);
   U367 : OAI21_X1 port map( A1 => n28688, A2 => n2233, B => n23544, ZN => 
                           n29052);
   U368 : AOI22_X1 port map( A1 => n9768, A2 => n9797, B1 => n23787, B2 => 
                           n9769, ZN => n32442);
   U378 : AND2_X1 port map( A1 => n23867, A2 => n17895, Z => n12090);
   U379 : OAI21_X1 port map( A1 => n9736, A2 => n976, B => n4408, ZN => n6041);
   U380 : NOR2_X1 port map( A1 => n29198, A2 => n33659, ZN => n33055);
   U381 : NOR2_X1 port map( A1 => n25987, A2 => n23575, ZN => n27329);
   U384 : NOR3_X1 port map( A1 => n2752, A2 => n23806, A3 => n28273, ZN => 
                           n9899);
   U385 : NOR2_X1 port map( A1 => n33828, A2 => n33827, ZN => n4374);
   U387 : NOR3_X1 port map( A1 => n32210, A2 => n7444, A3 => n32209, ZN => 
                           n31084);
   U392 : OAI21_X1 port map( A1 => n12070, A2 => n32522, B => n23897, ZN => 
                           n18117);
   U396 : NAND3_X1 port map( A1 => n8835, A2 => n31560, A3 => n23600, ZN => 
                           n6932);
   U397 : OAI21_X1 port map( A1 => n30621, A2 => n30620, B => n23878, ZN => 
                           n33370);
   U401 : AOI21_X1 port map( A1 => n30991, A2 => n23824, B => n27893, ZN => 
                           n24188);
   U402 : NAND2_X1 port map( A1 => n28016, A2 => n32209, ZN => n33043);
   U405 : NAND2_X1 port map( A1 => n33340, A2 => n3371, ZN => n32128);
   U416 : NAND2_X1 port map( A1 => n33005, A2 => n23576, ZN => n30803);
   U418 : NOR2_X1 port map( A1 => n11904, A2 => n23860, ZN => n12592);
   U419 : NOR3_X1 port map( A1 => n6662, A2 => n23756, A3 => n23760, ZN => 
                           n13903);
   U422 : OAI21_X1 port map( A1 => n6661, A2 => n15600, B => n17691, ZN => 
                           n32607);
   U423 : NAND2_X1 port map( A1 => n32986, A2 => n1920, ZN => n7777);
   U427 : AOI22_X1 port map( A1 => n15451, A2 => n33110, B1 => n2561, B2 => 
                           n2560, ZN => n33071);
   U431 : OAI21_X1 port map( A1 => n23634, A2 => n23633, B => n11240, ZN => 
                           n5227);
   U432 : AOI22_X1 port map( A1 => n16224, A2 => n23754, B1 => n28297, B2 => 
                           n23726, ZN => n33313);
   U433 : OR2_X1 port map( A1 => n4281, A2 => n707, Z => n31982);
   U434 : INV_X1 port map( I => n33867, ZN => n32425);
   U435 : AND2_X1 port map( A1 => n8270, A2 => n843, Z => n10143);
   U436 : INV_X1 port map( I => n16320, ZN => n23697);
   U437 : CLKBUF_X2 port map( I => n23588, Z => n33103);
   U443 : NOR2_X1 port map( A1 => n6414, A2 => n14975, ZN => n32801);
   U444 : INV_X1 port map( I => n14335, ZN => n23812);
   U450 : NOR2_X1 port map( A1 => n756, A2 => n29272, ZN => n10384);
   U454 : AND2_X1 port map( A1 => n14975, A2 => n14974, Z => n31981);
   U459 : NOR2_X1 port map( A1 => n4069, A2 => n34009, ZN => n32522);
   U460 : NOR2_X1 port map( A1 => n32610, A2 => n11923, ZN => n32609);
   U467 : NAND2_X1 port map( A1 => n17777, A2 => n980, ZN => n31759);
   U472 : OAI21_X1 port map( A1 => n27678, A2 => n1257, B => n32547, ZN => 
                           n11654);
   U474 : NOR2_X1 port map( A1 => n23897, A2 => n4069, ZN => n33096);
   U475 : NOR2_X1 port map( A1 => n32434, A2 => n32657, ZN => n7262);
   U478 : NAND2_X1 port map( A1 => n846, A2 => n13549, ZN => n33340);
   U481 : NAND2_X1 port map( A1 => n33670, A2 => n651, ZN => n23881);
   U486 : NOR2_X1 port map( A1 => n23775, A2 => n31810, ZN => n17750);
   U494 : NAND3_X1 port map( A1 => n26775, A2 => n16677, A3 => n17373, ZN => 
                           n32354);
   U495 : NAND2_X1 port map( A1 => n6247, A2 => n17726, ZN => n8836);
   U500 : OAI22_X1 port map( A1 => n8093, A2 => n33831, B1 => n23583, B2 => 
                           n27910, ZN => n33018);
   U501 : NOR2_X1 port map( A1 => n13905, A2 => n13413, ZN => n15600);
   U505 : NAND2_X1 port map( A1 => n23590, A2 => n6661, ZN => n17691);
   U507 : OR2_X1 port map( A1 => n23871, A2 => n6474, Z => n32004);
   U509 : BUF_X2 port map( I => n11923, Z => n33337);
   U510 : INV_X1 port map( I => n8838, ZN => n6247);
   U513 : INV_X1 port map( I => n32999, ZN => n2561);
   U518 : NAND2_X1 port map( A1 => n10279, A2 => n9375, ZN => n23882);
   U522 : NAND2_X1 port map( A1 => n33354, A2 => n32711, ZN => n5627);
   U525 : CLKBUF_X2 port map( I => n5736, Z => n33260);
   U526 : CLKBUF_X2 port map( I => n15865, Z => n14325);
   U527 : INV_X1 port map( I => n29472, ZN => n23824);
   U530 : BUF_X1 port map( I => n9939, Z => n33499);
   U531 : INV_X2 port map( I => n13998, ZN => n33789);
   U533 : NOR2_X1 port map( A1 => n14133, A2 => n32170, ZN => n23825);
   U536 : NAND2_X1 port map( A1 => n34036, A2 => n23767, ZN => n1610);
   U538 : NAND2_X1 port map( A1 => n13905, A2 => n26115, ZN => n16292);
   U544 : BUF_X2 port map( I => n23156, Z => n18204);
   U548 : BUF_X2 port map( I => n12974, Z => n12658);
   U555 : CLKBUF_X2 port map( I => n17857, Z => n25996);
   U563 : CLKBUF_X2 port map( I => n17812, Z => n3760);
   U567 : NAND2_X1 port map( A1 => n23867, A2 => n657, ZN => n10140);
   U573 : BUF_X2 port map( I => n23202, Z => n29217);
   U574 : INV_X1 port map( I => n23363, ZN => n8915);
   U575 : INV_X1 port map( I => n23496, ZN => n33111);
   U576 : INV_X1 port map( I => n23202, ZN => n10625);
   U579 : INV_X1 port map( I => n11504, ZN => n32214);
   U581 : NAND2_X1 port map( A1 => n1565, A2 => n1564, ZN => n27148);
   U587 : NAND2_X1 port map( A1 => n11741, A2 => n11740, ZN => n60);
   U591 : NAND2_X1 port map( A1 => n32513, A2 => n22863, ZN => n13918);
   U593 : NAND2_X1 port map( A1 => n33640, A2 => n5182, ZN => n33556);
   U595 : OAI21_X1 port map( A1 => n22838, A2 => n33596, B => n32827, ZN => 
                           n4871);
   U601 : NOR2_X1 port map( A1 => n6350, A2 => n29648, ZN => n32324);
   U602 : AND2_X1 port map( A1 => n5274, A2 => n10295, Z => n11538);
   U603 : NAND2_X1 port map( A1 => n2114, A2 => n8990, ZN => n2113);
   U604 : NOR2_X1 port map( A1 => n28689, A2 => n11059, ZN => n32513);
   U609 : NAND2_X1 port map( A1 => n29115, A2 => n17399, ZN => n4649);
   U611 : AOI22_X1 port map( A1 => n29329, A2 => n32935, B1 => n6433, B2 => 
                           n27814, ZN => n22721);
   U612 : CLKBUF_X2 port map( I => n1266, Z => n26373);
   U614 : NAND2_X1 port map( A1 => n4845, A2 => n28974, ZN => n4846);
   U617 : OAI21_X1 port map( A1 => n27212, A2 => n31936, B => n9293, ZN => 
                           n16879);
   U621 : NAND2_X1 port map( A1 => n32960, A2 => n32959, ZN => n29401);
   U623 : OAI21_X1 port map( A1 => n16975, A2 => n29391, B => n23026, ZN => 
                           n8853);
   U624 : NAND2_X1 port map( A1 => n27798, A2 => n15349, ZN => n33346);
   U643 : NAND2_X1 port map( A1 => n23090, A2 => n33968, ZN => n33932);
   U644 : AOI21_X1 port map( A1 => n22720, A2 => n31531, B => n32935, ZN => 
                           n27775);
   U645 : NAND2_X1 port map( A1 => n2712, A2 => n23106, ZN => n32827);
   U648 : OAI21_X1 port map( A1 => n11317, A2 => n33563, B => n33562, ZN => 
                           n22881);
   U649 : INV_X1 port map( I => n34017, ZN => n29427);
   U652 : OAI21_X1 port map( A1 => n33022, A2 => n30976, B => n32258, ZN => 
                           n22770);
   U653 : NOR2_X1 port map( A1 => n12181, A2 => n15317, ZN => n33510);
   U654 : AOI21_X1 port map( A1 => n32307, A2 => n23079, B => n6985, ZN => 
                           n32318);
   U665 : NAND2_X1 port map( A1 => n22769, A2 => n28415, ZN => n32580);
   U669 : OAI21_X1 port map( A1 => n4208, A2 => n23093, B => n776, ZN => n32964
                           );
   U671 : CLKBUF_X4 port map( I => n23087, Z => n6236);
   U677 : NAND2_X1 port map( A1 => n6149, A2 => n22473, ZN => n12418);
   U681 : NOR2_X1 port map( A1 => n22832, A2 => n23000, ZN => n22753);
   U682 : AND2_X1 port map( A1 => n6835, A2 => n6836, Z => n32868);
   U686 : INV_X1 port map( I => n22592, ZN => n22900);
   U688 : NOR2_X1 port map( A1 => n899, A2 => n30976, ZN => n32959);
   U691 : NAND2_X1 port map( A1 => n15935, A2 => n7047, ZN => n23479);
   U692 : CLKBUF_X2 port map( I => n22848, Z => n3184);
   U701 : NOR2_X1 port map( A1 => n30909, A2 => n28313, ZN => n15915);
   U702 : NAND2_X1 port map( A1 => n14183, A2 => n5915, ZN => n27296);
   U705 : NAND2_X1 port map( A1 => n22792, A2 => n27090, ZN => n32560);
   U706 : NAND3_X1 port map( A1 => n15389, A2 => n27090, A3 => n4113, ZN => 
                           n28178);
   U707 : AOI21_X1 port map( A1 => n11495, A2 => n32820, B => n1106, ZN => 
                           n33179);
   U711 : NOR2_X1 port map( A1 => n32842, A2 => n34017, ZN => n15362);
   U713 : INV_X1 port map( I => n5682, ZN => n30825);
   U714 : NAND2_X1 port map( A1 => n22894, A2 => n30909, ZN => n15190);
   U720 : NOR2_X1 port map( A1 => n12586, A2 => n28697, ZN => n22835);
   U721 : AOI21_X1 port map( A1 => n23055, A2 => n3007, B => n29107, ZN => 
                           n14417);
   U722 : NOR2_X1 port map( A1 => n32500, A2 => n23056, ZN => n32424);
   U726 : NAND3_X1 port map( A1 => n7181, A2 => n898, A3 => n4734, ZN => n26312
                           );
   U727 : NAND2_X1 port map( A1 => n26526, A2 => n33132, ZN => n22709);
   U729 : INV_X1 port map( I => n22832, ZN => n79);
   U731 : INV_X1 port map( I => n22960, ZN => n23082);
   U737 : AND2_X1 port map( A1 => n9963, A2 => n30868, Z => n32092);
   U740 : INV_X1 port map( I => n15456, ZN => n12727);
   U742 : INV_X2 port map( I => n5274, ZN => n11317);
   U745 : AND2_X1 port map( A1 => n10528, A2 => n6975, Z => n8022);
   U746 : CLKBUF_X2 port map( I => n27419, Z => n32119);
   U749 : INV_X2 port map( I => n22795, ZN => n23042);
   U750 : INV_X2 port map( I => n22798, ZN => n772);
   U753 : INV_X1 port map( I => n22957, ZN => n9778);
   U756 : NOR2_X1 port map( A1 => n4580, A2 => n16486, ZN => n13648);
   U757 : CLKBUF_X2 port map( I => n30293, Z => n27798);
   U758 : INV_X2 port map( I => n31325, ZN => n17211);
   U763 : BUF_X2 port map( I => n13762, Z => n6800);
   U764 : BUF_X2 port map( I => n6605, Z => n30909);
   U765 : NOR2_X1 port map( A1 => n22885, A2 => n1577, ZN => n22815);
   U766 : INV_X1 port map( I => n6799, ZN => n22950);
   U772 : INV_X2 port map( I => n30297, ZN => n1278);
   U779 : NAND3_X1 port map( A1 => n32192, A2 => n32191, A3 => n5769, ZN => 
                           n5573);
   U781 : NAND2_X1 port map( A1 => n22530, A2 => n22531, ZN => n12256);
   U784 : AND2_X1 port map( A1 => n22442, A2 => n28692, Z => n31934);
   U785 : NAND2_X1 port map( A1 => n9425, A2 => n22539, ZN => n4502);
   U787 : NOR3_X1 port map( A1 => n5597, A2 => n22534, A3 => n16434, ZN => 
                           n4503);
   U794 : AOI22_X1 port map( A1 => n30065, A2 => n22570, B1 => n1297, B2 => 
                           n18073, ZN => n33855);
   U798 : NAND2_X1 port map( A1 => n32194, A2 => n32193, ZN => n32192);
   U801 : OAI21_X1 port map( A1 => n33061, A2 => n22407, B => n32448, ZN => 
                           n29982);
   U805 : NAND2_X1 port map( A1 => n22530, A2 => n15643, ZN => n6505);
   U809 : INV_X1 port map( I => n22612, ZN => n32757);
   U811 : AOI21_X1 port map( A1 => n22671, A2 => n29371, B => n26098, ZN => 
                           n33262);
   U814 : NAND2_X1 port map( A1 => n2066, A2 => n22487, ZN => n32680);
   U817 : NOR2_X1 port map( A1 => n29078, A2 => n11917, ZN => n33502);
   U823 : AOI21_X1 port map( A1 => n11874, A2 => n16556, B => n16570, ZN => 
                           n33974);
   U831 : OAI22_X1 port map( A1 => n14137, A2 => n5743, B1 => n22658, B2 => 
                           n22659, ZN => n22366);
   U838 : AOI21_X1 port map( A1 => n27959, A2 => n2418, B => n11250, ZN => 
                           n33463);
   U840 : AND2_X1 port map( A1 => n22476, A2 => n22394, Z => n15103);
   U842 : INV_X1 port map( I => n33227, ZN => n3596);
   U851 : NAND2_X1 port map( A1 => n12899, A2 => n22586, ZN => n9452);
   U856 : NAND2_X1 port map( A1 => n29261, A2 => n11920, ZN => n21963);
   U858 : NOR2_X1 port map( A1 => n34035, A2 => n5597, ZN => n33061);
   U861 : INV_X1 port map( I => n15746, ZN => n32193);
   U864 : AOI21_X1 port map( A1 => n18038, A2 => n22427, B => n28170, ZN => 
                           n32446);
   U868 : OR2_X1 port map( A1 => n22476, A2 => n29101, Z => n12072);
   U870 : OR2_X1 port map( A1 => n22474, A2 => n22476, Z => n17247);
   U872 : INV_X2 port map( I => n29508, ZN => n33455);
   U881 : NOR2_X1 port map( A1 => n29078, A2 => n908, ZN => n32823);
   U883 : NOR3_X1 port map( A1 => n22636, A2 => n22640, A3 => n12043, ZN => 
                           n22731);
   U902 : NAND3_X1 port map( A1 => n16529, A2 => n22926, A3 => n22658, ZN => 
                           n33368);
   U905 : OAI21_X1 port map( A1 => n30334, A2 => n29461, B => n30065, ZN => 
                           n33982);
   U906 : NOR2_X1 port map( A1 => n14728, A2 => n16375, ZN => n12335);
   U909 : INV_X1 port map( I => n6976, ZN => n22343);
   U910 : BUF_X2 port map( I => n6976, Z => n239);
   U913 : INV_X1 port map( I => n26884, ZN => n32831);
   U936 : INV_X1 port map( I => n29288, ZN => n22558);
   U948 : INV_X2 port map( I => n22476, ZN => n22377);
   U952 : NAND2_X1 port map( A1 => n2858, A2 => n5961, ZN => n7848);
   U955 : INV_X1 port map( I => n14227, ZN => n32334);
   U956 : NAND2_X1 port map( A1 => n22644, A2 => n22645, ZN => n33026);
   U965 : NAND2_X1 port map( A1 => n22330, A2 => n1116, ZN => n11011);
   U966 : NOR2_X1 port map( A1 => n14728, A2 => n12338, ZN => n27878);
   U968 : NAND3_X1 port map( A1 => n6242, A2 => n6244, A3 => n22639, ZN => 
                           n32987);
   U969 : NAND2_X1 port map( A1 => n22332, A2 => n28692, ZN => n22569);
   U971 : NAND2_X1 port map( A1 => n14251, A2 => n32830, ZN => n12840);
   U978 : NAND3_X1 port map( A1 => n33628, A2 => n6186, A3 => n6187, ZN => 
                           n33619);
   U980 : INV_X1 port map( I => n9630, ZN => n33281);
   U981 : INV_X1 port map( I => n22367, ZN => n31964);
   U986 : AND2_X1 port map( A1 => n27933, A2 => n26317, Z => n22688);
   U988 : CLKBUF_X2 port map( I => n8420, Z => n327);
   U993 : BUF_X2 port map( I => n9515, Z => n5743);
   U996 : BUF_X2 port map( I => n22350, Z => n1294);
   U997 : NOR2_X1 port map( A1 => n33320, A2 => n8409, ZN => n32569);
   U999 : NAND2_X1 port map( A1 => n8131, A2 => n12496, ZN => n9272);
   U1002 : INV_X1 port map( I => n4916, ZN => n10654);
   U1010 : AOI21_X1 port map( A1 => n32797, A2 => n17076, B => n10354, ZN => 
                           n13070);
   U1012 : NOR2_X1 port map( A1 => n998, A2 => n1116, ZN => n28019);
   U1019 : INV_X1 port map( I => n31692, ZN => n10183);
   U1021 : INV_X1 port map( I => n5961, ZN => n5991);
   U1026 : INV_X2 port map( I => n1926, ZN => n16647);
   U1028 : INV_X1 port map( I => n22157, ZN => n33593);
   U1035 : INV_X1 port map( I => n8617, ZN => n22296);
   U1039 : BUF_X2 port map( I => n22160, Z => n4295);
   U1049 : INV_X1 port map( I => n16237, ZN => n1307);
   U1055 : INV_X1 port map( I => n22032, ZN => n32714);
   U1057 : INV_X1 port map( I => n22211, ZN => n33151);
   U1062 : INV_X1 port map( I => n29137, ZN => n34063);
   U1064 : INV_X1 port map( I => n22113, ZN => n31165);
   U1072 : INV_X1 port map( I => n22076, ZN => n21892);
   U1075 : INV_X1 port map( I => n22283, ZN => n1129);
   U1076 : NAND2_X1 port map( A1 => n11727, A2 => n21964, ZN => n11359);
   U1079 : INV_X1 port map( I => n22042, ZN => n34014);
   U1080 : INV_X1 port map( I => n21945, ZN => n32126);
   U1081 : NAND3_X1 port map( A1 => n21933, A2 => n21932, A3 => n28895, ZN => 
                           n6426);
   U1082 : NOR2_X1 port map( A1 => n15639, A2 => n33298, ZN => n10234);
   U1087 : NAND3_X1 port map( A1 => n33481, A2 => n6238, A3 => n6237, ZN => 
                           n33471);
   U1089 : NAND2_X1 port map( A1 => n5228, A2 => n26671, ZN => n31657);
   U1090 : NAND3_X1 port map( A1 => n28895, A2 => n30440, A3 => n10699, ZN => 
                           n32608);
   U1091 : NAND2_X1 port map( A1 => n15465, A2 => n32833, ZN => n32832);
   U1092 : AOI22_X1 port map( A1 => n13248, A2 => n21546, B1 => n17429, B2 => 
                           n21730, ZN => n7457);
   U1097 : AND2_X1 port map( A1 => n2643, A2 => n21704, Z => n32071);
   U1099 : OAI21_X1 port map( A1 => n31260, A2 => n32384, B => n8029, ZN => 
                           n27631);
   U1101 : NOR2_X1 port map( A1 => n21856, A2 => n13116, ZN => n2352);
   U1106 : AOI22_X1 port map( A1 => n16016, A2 => n276, B1 => n31220, B2 => 
                           n21778, ZN => n33676);
   U1108 : OAI21_X1 port map( A1 => n14641, A2 => n17078, B => n32282, ZN => 
                           n9686);
   U1117 : INV_X1 port map( I => n396, ZN => n32321);
   U1120 : OAI21_X1 port map( A1 => n17225, A2 => n17226, B => n423, ZN => 
                           n8077);
   U1126 : OAI21_X1 port map( A1 => n11644, A2 => n29784, B => n8029, ZN => 
                           n11643);
   U1128 : OAI21_X1 port map( A1 => n33520, A2 => n33519, B => n4331, ZN => 
                           n6766);
   U1129 : NOR2_X1 port map( A1 => n14642, A2 => n914, ZN => n28393);
   U1142 : AOI21_X1 port map( A1 => n12626, A2 => n11619, B => n26474, ZN => 
                           n16192);
   U1146 : NOR2_X1 port map( A1 => n915, A2 => n31911, ZN => n32325);
   U1151 : NAND2_X1 port map( A1 => n33242, A2 => n30769, ZN => n32497);
   U1153 : NOR2_X1 port map( A1 => n21652, A2 => n7553, ZN => n33031);
   U1158 : OR2_X1 port map( A1 => n21466, A2 => n31085, Z => n32073);
   U1160 : INV_X1 port map( I => n32208, ZN => n7366);
   U1161 : NAND2_X1 port map( A1 => n21741, A2 => n423, ZN => n33364);
   U1165 : NAND2_X1 port map( A1 => n21625, A2 => n32865, ZN => n32320);
   U1168 : NOR2_X1 port map( A1 => n2643, A2 => n14681, ZN => n21792);
   U1171 : INV_X1 port map( I => n32435, ZN => n29286);
   U1172 : INV_X1 port map( I => n912, ZN => n33842);
   U1177 : INV_X2 port map( I => n1013, ZN => n32499);
   U1180 : OAI21_X1 port map( A1 => n14384, A2 => n31042, B => n32384, ZN => 
                           n32208);
   U1188 : NAND2_X1 port map( A1 => n21512, A2 => n26622, ZN => n11719);
   U1190 : AND2_X1 port map( A1 => n21860, A2 => n3286, Z => n13116);
   U1202 : NOR2_X1 port map( A1 => n11596, A2 => n11981, ZN => n33520);
   U1207 : NAND2_X1 port map( A1 => n13114, A2 => n30885, ZN => n21586);
   U1209 : NAND2_X1 port map( A1 => n12221, A2 => n21719, ZN => n21490);
   U1214 : NAND3_X1 port map( A1 => n33481, A2 => n21713, A3 => n5704, ZN => 
                           n32994);
   U1216 : NAND2_X1 port map( A1 => n12866, A2 => n13872, ZN => n27023);
   U1218 : INV_X2 port map( I => n31956, ZN => n1015);
   U1219 : INV_X1 port map( I => n2386, ZN => n21489);
   U1220 : NOR2_X1 port map( A1 => n30769, A2 => n32252, ZN => n4432);
   U1221 : INV_X1 port map( I => n21604, ZN => n1318);
   U1222 : INV_X1 port map( I => n21512, ZN => n1327);
   U1223 : INV_X1 port map( I => n16954, ZN => n21585);
   U1225 : INV_X2 port map( I => n1313, ZN => n517);
   U1228 : INV_X1 port map( I => n33146, ZN => n33731);
   U1230 : NAND2_X1 port map( A1 => n2386, A2 => n31954, ZN => n21717);
   U1239 : BUF_X2 port map( I => n7592, Z => n33481);
   U1245 : INV_X1 port map( I => n31960, ZN => n32643);
   U1246 : CLKBUF_X1 port map( I => n5086, Z => n31953);
   U1248 : NAND2_X1 port map( A1 => n32800, A2 => n15371, ZN => n32372);
   U1249 : INV_X1 port map( I => n7592, ZN => n16441);
   U1250 : INV_X1 port map( I => n12211, ZN => n5228);
   U1252 : NAND2_X1 port map( A1 => n21264, A2 => n21263, ZN => n12640);
   U1258 : INV_X1 port map( I => n9472, ZN => n5494);
   U1260 : INV_X1 port map( I => n3203, ZN => n32505);
   U1262 : INV_X2 port map( I => n7868, ZN => n27532);
   U1263 : AND2_X1 port map( A1 => n21466, A2 => n1136, Z => n4842);
   U1264 : OAI21_X1 port map( A1 => n21222, A2 => n21109, B => n26166, ZN => 
                           n2570);
   U1268 : INV_X2 port map( I => n28099, ZN => n777);
   U1270 : INV_X2 port map( I => n11755, ZN => n7969);
   U1271 : NAND2_X1 port map( A1 => n33802, A2 => n2834, ZN => n5086);
   U1272 : NAND2_X1 port map( A1 => n32455, A2 => n32454, ZN => n21134);
   U1277 : NOR2_X1 port map( A1 => n16204, A2 => n33167, ZN => n17432);
   U1281 : NAND3_X1 port map( A1 => n33926, A2 => n21336, A3 => n33925, ZN => 
                           n5250);
   U1286 : NAND3_X1 port map( A1 => n33755, A2 => n4988, A3 => n4324, ZN => 
                           n4062);
   U1291 : NOR2_X1 port map( A1 => n11138, A2 => n21411, ZN => n2722);
   U1296 : OAI21_X1 port map( A1 => n21403, A2 => n596, B => n12654, ZN => 
                           n29742);
   U1301 : OAI21_X1 port map( A1 => n1867, A2 => n1868, B => n21353, ZN => 
                           n32330);
   U1309 : OR2_X1 port map( A1 => n9191, A2 => n12323, Z => n10573);
   U1312 : INV_X1 port map( I => n11299, ZN => n31329);
   U1313 : AOI22_X1 port map( A1 => n21099, A2 => n17437, B1 => n154, B2 => 
                           n21138, ZN => n21067);
   U1318 : OAI22_X1 port map( A1 => n29802, A2 => n21363, B1 => n21183, B2 => 
                           n21182, ZN => n17685);
   U1319 : INV_X1 port map( I => n13593, ZN => n8587);
   U1321 : NAND2_X1 port map( A1 => n31730, A2 => n31728, ZN => n18208);
   U1325 : AND2_X1 port map( A1 => n2738, A2 => n9133, Z => n29394);
   U1328 : INV_X1 port map( I => n32655, ZN => n34081);
   U1329 : OR2_X1 port map( A1 => n11967, A2 => n21358, Z => n10092);
   U1330 : NOR2_X1 port map( A1 => n4274, A2 => n17341, ZN => n5039);
   U1333 : NOR2_X1 port map( A1 => n32273, A2 => n8560, ZN => n32407);
   U1336 : OAI21_X1 port map( A1 => n31997, A2 => n5239, B => n32203, ZN => 
                           n32979);
   U1342 : NAND3_X1 port map( A1 => n2831, A2 => n2833, A3 => n26167, ZN => 
                           n33802);
   U1343 : NAND2_X1 port map( A1 => n33972, A2 => n13073, ZN => n13366);
   U1345 : NAND2_X1 port map( A1 => n2370, A2 => n21441, ZN => n32808);
   U1358 : OAI21_X1 port map( A1 => n1020, A2 => n7007, B => n3672, ZN => n7051
                           );
   U1359 : NOR2_X1 port map( A1 => n26167, A2 => n1329, ZN => n33113);
   U1361 : NOR3_X1 port map( A1 => n31965, A2 => n28642, A3 => n29460, ZN => 
                           n27608);
   U1368 : NAND2_X1 port map( A1 => n5480, A2 => n32347, ZN => n33925);
   U1370 : OAI21_X1 port map( A1 => n922, A2 => n13255, B => n6408, ZN => 
                           n16640);
   U1372 : NOR2_X1 port map( A1 => n32550, A2 => n1141, ZN => n4497);
   U1374 : NAND2_X1 port map( A1 => n32457, A2 => n32456, ZN => n32455);
   U1375 : NAND2_X1 port map( A1 => n5469, A2 => n26021, ZN => n33523);
   U1378 : NOR2_X1 port map( A1 => n4341, A2 => n30813, ZN => n17011);
   U1382 : OAI22_X1 port map( A1 => n810, A2 => n21365, B1 => n4076, B2 => 
                           n17466, ZN => n29678);
   U1383 : NOR2_X1 port map( A1 => n21251, A2 => n21078, ZN => n30050);
   U1385 : NOR2_X1 port map( A1 => n18106, A2 => n15522, ZN => n33647);
   U1386 : INV_X1 port map( I => n21443, ZN => n32457);
   U1387 : NAND2_X1 port map( A1 => n32777, A2 => n32776, ZN => n5018);
   U1389 : NAND2_X1 port map( A1 => n2241, A2 => n2242, ZN => n33735);
   U1392 : NAND2_X1 port map( A1 => n16180, A2 => n16526, ZN => n32456);
   U1394 : AND2_X1 port map( A1 => n11967, A2 => n21358, Z => n31674);
   U1396 : NAND2_X1 port map( A1 => n21381, A2 => n16906, ZN => n15985);
   U1401 : NAND2_X1 port map( A1 => n21078, A2 => n4518, ZN => n13401);
   U1403 : NAND2_X1 port map( A1 => n14074, A2 => n21406, ZN => n32322);
   U1408 : NAND2_X1 port map( A1 => n33741, A2 => n4324, ZN => n33171);
   U1418 : OR2_X1 port map( A1 => n5395, A2 => n8028, Z => n31997);
   U1420 : NAND2_X1 port map( A1 => n21452, A2 => n780, ZN => n29122);
   U1426 : BUF_X2 port map( I => n21438, Z => n33745);
   U1429 : NOR2_X1 port map( A1 => n21255, A2 => n28257, ZN => n33137);
   U1439 : NAND2_X1 port map( A1 => n33849, A2 => n32147, ZN => n4076);
   U1445 : NOR2_X1 port map( A1 => n33889, A2 => n33888, ZN => n33887);
   U1446 : NOR2_X1 port map( A1 => n17956, A2 => n349, ZN => n32350);
   U1447 : NAND2_X1 port map( A1 => n4337, A2 => n4971, ZN => n32203);
   U1448 : NOR3_X1 port map( A1 => n21163, A2 => n27170, A3 => n11734, ZN => 
                           n33350);
   U1450 : NOR2_X1 port map( A1 => n21219, A2 => n33496, ZN => n32273);
   U1455 : NOR2_X1 port map( A1 => n2738, A2 => n8924, ZN => n8937);
   U1457 : NAND2_X1 port map( A1 => n31909, A2 => n16668, ZN => n21407);
   U1459 : INV_X2 port map( I => n16633, ZN => n20949);
   U1460 : BUF_X2 port map( I => n3879, Z => n30813);
   U1461 : BUF_X2 port map( I => n21395, Z => n27955);
   U1468 : CLKBUF_X2 port map( I => n26677, Z => n34131);
   U1471 : INV_X1 port map( I => n3193, ZN => n32777);
   U1472 : BUF_X2 port map( I => n6493, Z => n34054);
   U1473 : NAND2_X1 port map( A1 => n6855, A2 => n32883, ZN => n32239);
   U1475 : OAI21_X1 port map( A1 => n349, A2 => n33496, B => n33495, ZN => 
                           n21146);
   U1476 : INV_X2 port map( I => n21452, ZN => n1143);
   U1478 : OR2_X1 port map( A1 => n34156, A2 => n28260, Z => n31989);
   U1487 : INV_X1 port map( I => n4145, ZN => n1703);
   U1488 : BUF_X2 port map( I => n9351, Z => n9186);
   U1489 : CLKBUF_X2 port map( I => n13723, Z => n32147);
   U1490 : NAND2_X1 port map( A1 => n13692, A2 => n21357, ZN => n33336);
   U1509 : INV_X1 port map( I => n29901, ZN => n33496);
   U1510 : BUF_X2 port map( I => n10599, Z => n33498);
   U1513 : BUF_X2 port map( I => n21258, Z => n16652);
   U1516 : BUF_X2 port map( I => n13195, Z => n10599);
   U1520 : OR2_X1 port map( A1 => n31290, A2 => n31291, Z => n32889);
   U1523 : INV_X1 port map( I => n20641, ZN => n20920);
   U1541 : CLKBUF_X2 port map( I => n4680, Z => n29918);
   U1545 : INV_X1 port map( I => n20970, ZN => n29879);
   U1546 : INV_X1 port map( I => n20786, ZN => n21024);
   U1553 : INV_X1 port map( I => n20928, ZN => n12559);
   U1555 : NOR2_X1 port map( A1 => n17317, A2 => n4980, ZN => n32230);
   U1570 : NAND2_X1 port map( A1 => n10105, A2 => n5735, ZN => n5734);
   U1572 : OAI22_X1 port map( A1 => n32033, A2 => n8031, B1 => n28799, B2 => 
                           n1356, ZN => n32249);
   U1573 : NAND3_X1 port map( A1 => n20302, A2 => n27600, A3 => n20360, ZN => 
                           n12553);
   U1575 : OR2_X1 port map( A1 => n14161, A2 => n20628, Z => n20387);
   U1576 : NOR2_X1 port map( A1 => n15898, A2 => n15027, ZN => n11840);
   U1577 : AND2_X1 port map( A1 => n20627, A2 => n9014, Z => n14571);
   U1581 : OR2_X1 port map( A1 => n20534, A2 => n28028, Z => n30728);
   U1582 : AND2_X1 port map( A1 => n33117, A2 => n14138, Z => n2145);
   U1588 : AND2_X1 port map( A1 => n33117, A2 => n20468, Z => n3227);
   U1591 : AOI22_X1 port map( A1 => n15638, A2 => n26756, B1 => n11017, B2 => 
                           n1347, ZN => n33052);
   U1593 : CLKBUF_X2 port map( I => n28011, Z => n34052);
   U1594 : NAND2_X1 port map( A1 => n32765, A2 => n31891, ZN => n32764);
   U1597 : NAND2_X1 port map( A1 => n20607, A2 => n7577, ZN => n33843);
   U1601 : NAND2_X1 port map( A1 => n20551, A2 => n10834, ZN => n12148);
   U1602 : NOR2_X1 port map( A1 => n20243, A2 => n26471, ZN => n32684);
   U1604 : NAND3_X1 port map( A1 => n32941, A2 => n32940, A3 => n32939, ZN => 
                           n29431);
   U1606 : NAND3_X1 port map( A1 => n31969, A2 => n20072, A3 => n20073, ZN => 
                           n3904);
   U1610 : NOR3_X1 port map( A1 => n15898, A2 => n16518, A3 => n20534, ZN => 
                           n184);
   U1615 : AND2_X1 port map( A1 => n33117, A2 => n20467, Z => n3463);
   U1619 : AND2_X1 port map( A1 => n16144, A2 => n11984, Z => n20194);
   U1628 : INV_X1 port map( I => n20608, ZN => n33397);
   U1641 : INV_X1 port map( I => n10312, ZN => n29553);
   U1643 : AND2_X1 port map( A1 => n20515, A2 => n7242, Z => n6121);
   U1649 : BUF_X2 port map( I => n30643, Z => n4071);
   U1653 : CLKBUF_X2 port map( I => n20632, Z => n111);
   U1657 : NAND2_X1 port map( A1 => n12421, A2 => n14719, ZN => n17672);
   U1660 : BUF_X2 port map( I => n30763, Z => n31961);
   U1662 : CLKBUF_X1 port map( I => n14545, Z => n29623);
   U1666 : INV_X1 port map( I => n31811, ZN => n33398);
   U1671 : NAND2_X1 port map( A1 => n28085, A2 => n20563, ZN => n33194);
   U1675 : NAND2_X1 port map( A1 => n20492, A2 => n26585, ZN => n33944);
   U1677 : NAND2_X1 port map( A1 => n3084, A2 => n20339, ZN => n12244);
   U1683 : NOR2_X1 port map( A1 => n25966, A2 => n20602, ZN => n32341);
   U1686 : NAND2_X1 port map( A1 => n9403, A2 => n20472, ZN => n34113);
   U1689 : NOR2_X1 port map( A1 => n12966, A2 => n12421, ZN => n33734);
   U1692 : AND2_X1 port map( A1 => n26566, A2 => n32989, Z => n31975);
   U1696 : INV_X1 port map( I => n30643, ZN => n10106);
   U1697 : INV_X1 port map( I => n3157, ZN => n33091);
   U1699 : NOR2_X1 port map( A1 => n16218, A2 => n7486, ZN => n33776);
   U1701 : INV_X1 port map( I => n20549, ZN => n31390);
   U1704 : BUF_X2 port map( I => n28840, Z => n33730);
   U1707 : OR2_X1 port map( A1 => n20613, A2 => n9252, Z => n7872);
   U1709 : NAND2_X1 port map( A1 => n28028, A2 => n32240, ZN => n11036);
   U1710 : NAND2_X1 port map( A1 => n20630, A2 => n31471, ZN => n15225);
   U1716 : OAI21_X1 port map( A1 => n939, A2 => n31442, B => n19949, ZN => 
                           n17496);
   U1717 : NAND2_X1 port map( A1 => n30845, A2 => n149, ZN => n34032);
   U1718 : NAND2_X1 port map( A1 => n32377, A2 => n19820, ZN => n11402);
   U1719 : NOR2_X1 port map( A1 => n32197, A2 => n29187, ZN => n2550);
   U1721 : OAI21_X1 port map( A1 => n31993, A2 => n11142, B => n29233, ZN => 
                           n11141);
   U1722 : NAND2_X1 port map( A1 => n11510, A2 => n12398, ZN => n32956);
   U1724 : OAI21_X1 port map( A1 => n31593, A2 => n16159, B => n20033, ZN => 
                           n33732);
   U1728 : NAND2_X1 port map( A1 => n34006, A2 => n16489, ZN => n3094);
   U1732 : OAI21_X1 port map( A1 => n4215, A2 => n16346, B => n34051, ZN => 
                           n17242);
   U1735 : OAI21_X1 port map( A1 => n19996, A2 => n19922, B => n4674, ZN => 
                           n4266);
   U1737 : NOR2_X1 port map( A1 => n19932, A2 => n8817, ZN => n10440);
   U1738 : NAND2_X1 port map( A1 => n13569, A2 => n19925, ZN => n32719);
   U1743 : AOI21_X1 port map( A1 => n431, A2 => n19840, B => n33504, ZN => 
                           n16924);
   U1746 : NAND2_X1 port map( A1 => n4215, A2 => n17243, ZN => n34051);
   U1751 : INV_X1 port map( I => n6961, ZN => n33148);
   U1753 : NOR3_X1 port map( A1 => n20135, A2 => n32141, A3 => n12682, ZN => 
                           n30155);
   U1754 : NAND2_X1 port map( A1 => n9619, A2 => n1168, ZN => n32674);
   U1755 : NOR2_X1 port map( A1 => n4371, A2 => n19998, ZN => n15366);
   U1756 : NOR2_X1 port map( A1 => n19854, A2 => n19855, ZN => n20070);
   U1758 : NAND2_X1 port map( A1 => n7309, A2 => n3090, ZN => n33439);
   U1761 : OAI21_X1 port map( A1 => n3989, A2 => n11961, B => n33627, ZN => 
                           n28459);
   U1763 : NOR2_X1 port map( A1 => n12075, A2 => n17495, ZN => n34006);
   U1765 : NOR2_X1 port map( A1 => n20020, A2 => n20120, ZN => n19812);
   U1768 : NAND2_X1 port map( A1 => n19898, A2 => n16092, ZN => n14712);
   U1769 : NAND2_X1 port map( A1 => n29853, A2 => n19961, ZN => n33504);
   U1770 : NOR2_X1 port map( A1 => n15192, A2 => n29040, ZN => n15477);
   U1773 : NAND2_X1 port map( A1 => n16977, A2 => n19920, ZN => n32792);
   U1775 : AOI21_X1 port map( A1 => n33264, A2 => n16848, B => n13583, ZN => 
                           n33553);
   U1778 : INV_X1 port map( I => n1826, ZN => n33526);
   U1785 : NOR2_X1 port map( A1 => n5966, A2 => n6962, ZN => n32479);
   U1786 : NAND3_X1 port map( A1 => n8259, A2 => n11199, A3 => n20154, ZN => 
                           n19621);
   U1789 : INV_X1 port map( I => n10286, ZN => n32197);
   U1790 : OAI21_X1 port map( A1 => n13348, A2 => n6444, B => n822, ZN => 
                           n33769);
   U1791 : NAND3_X1 port map( A1 => n7460, A2 => n16491, A3 => n7461, ZN => 
                           n1814);
   U1793 : NOR3_X1 port map( A1 => n19992, A2 => n19993, A3 => n1170, ZN => 
                           n33271);
   U1794 : INV_X1 port map( I => n26237, ZN => n33714);
   U1796 : OR2_X1 port map( A1 => n16625, A2 => n17127, Z => n8137);
   U1798 : AND2_X1 port map( A1 => n16595, A2 => n14815, Z => n9450);
   U1802 : AND2_X1 port map( A1 => n28293, A2 => n17882, Z => n31991);
   U1805 : NOR2_X1 port map( A1 => n28293, A2 => n16681, ZN => n19842);
   U1815 : AND2_X1 port map( A1 => n27748, A2 => n26237, Z => n11949);
   U1816 : OR2_X1 port map( A1 => n11720, A2 => n10934, Z => n14306);
   U1819 : NOR2_X1 port map( A1 => n6344, A2 => n29446, ZN => n19950);
   U1824 : CLKBUF_X2 port map( I => n6275, Z => n26615);
   U1825 : INV_X1 port map( I => n19966, ZN => n14575);
   U1827 : BUF_X2 port map( I => n19833, Z => n20136);
   U1834 : BUF_X2 port map( I => n11720, Z => n29187);
   U1838 : INV_X2 port map( I => n19938, ZN => n1161);
   U1840 : INV_X1 port map( I => n32915, ZN => n19885);
   U1842 : INV_X1 port map( I => n9161, ZN => n19616);
   U1846 : NAND2_X1 port map( A1 => n6022, A2 => n19056, ZN => n11867);
   U1850 : CLKBUF_X2 port map( I => n19778, Z => n28908);
   U1853 : INV_X1 port map( I => n24831, ZN => n32981);
   U1858 : INV_X1 port map( I => n19778, ZN => n33995);
   U1859 : OAI21_X1 port map( A1 => n17677, A2 => n17678, B => n31970, ZN => 
                           n33088);
   U1861 : OAI21_X1 port map( A1 => n28025, A2 => n18230, B => n763, ZN => 
                           n32431);
   U1863 : AOI22_X1 port map( A1 => n19119, A2 => n19181, B1 => n29769, B2 => 
                           n14424, ZN => n14423);
   U1866 : OR2_X1 port map( A1 => n28949, A2 => n19080, Z => n32057);
   U1870 : NOR2_X1 port map( A1 => n27965, A2 => n25967, ZN => n33825);
   U1872 : NAND2_X1 port map( A1 => n19074, A2 => n30760, ZN => n33852);
   U1884 : NAND2_X1 port map( A1 => n19311, A2 => n19312, ZN => n9683);
   U1888 : NOR2_X1 port map( A1 => n1807, A2 => n4643, ZN => n401);
   U1889 : NOR2_X1 port map( A1 => n26518, A2 => n11085, ZN => n11802);
   U1892 : CLKBUF_X1 port map( I => n29815, Z => n33635);
   U1894 : CLKBUF_X1 port map( I => n30894, Z => n33712);
   U1896 : AND2_X1 port map( A1 => n10472, A2 => n31970, Z => n32011);
   U1900 : NAND2_X1 port map( A1 => n4714, A2 => n9646, ZN => n16874);
   U1902 : AOI21_X1 port map( A1 => n11074, A2 => n3093, B => n2081, ZN => 
                           n28345);
   U1903 : NAND2_X1 port map( A1 => n33967, A2 => n4643, ZN => n30661);
   U1910 : AOI21_X1 port map( A1 => n826, A2 => n19290, B => n19288, ZN => 
                           n2717);
   U1911 : OAI21_X1 port map( A1 => n33143, A2 => n19147, B => n15534, ZN => 
                           n32293);
   U1914 : AND2_X1 port map( A1 => n7810, A2 => n19249, Z => n9648);
   U1915 : OAI21_X1 port map( A1 => n32653, A2 => n26037, B => n17311, ZN => 
                           n17819);
   U1918 : INV_X1 port map( I => n19348, ZN => n33232);
   U1919 : INV_X1 port map( I => n9677, ZN => n32219);
   U1924 : INV_X1 port map( I => n5625, ZN => n18977);
   U1925 : NOR2_X1 port map( A1 => n25960, A2 => n4747, ZN => n33671);
   U1927 : INV_X1 port map( I => n19308, ZN => n33718);
   U1928 : NOR2_X1 port map( A1 => n19102, A2 => n944, ZN => n8192);
   U1937 : INV_X1 port map( I => n18945, ZN => n33967);
   U1940 : INV_X1 port map( I => n28379, ZN => n32138);
   U1941 : NAND2_X1 port map( A1 => n19078, A2 => n30501, ZN => n30933);
   U1942 : INV_X1 port map( I => n19260, ZN => n32790);
   U1949 : INV_X1 port map( I => n31947, ZN => n27970);
   U1951 : BUF_X2 port map( I => n10228, Z => n10227);
   U1952 : NOR2_X1 port map( A1 => n18976, A2 => n14892, ZN => n18945);
   U1953 : NAND2_X1 port map( A1 => n764, A2 => n19167, ZN => n10353);
   U1958 : AOI22_X1 port map( A1 => n18641, A2 => n28238, B1 => n4259, B2 => 
                           n18642, ZN => n32121);
   U1959 : NOR2_X1 port map( A1 => n18974, A2 => n11322, ZN => n34031);
   U1963 : CLKBUF_X2 port map( I => n30865, Z => n31948);
   U1965 : INV_X2 port map( I => n18017, ZN => n1384);
   U1967 : AOI22_X1 port map( A1 => n18506, A2 => n9729, B1 => n18507, B2 => 
                           n1439, ZN => n33396);
   U1973 : BUF_X4 port map( I => n10953, Z => n2612);
   U1974 : NOR2_X1 port map( A1 => n18866, A2 => n711, ZN => n2507);
   U1976 : NOR2_X1 port map( A1 => n33528, A2 => n33559, ZN => n13112);
   U1979 : AND2_X1 port map( A1 => n18566, A2 => n18324, Z => n32009);
   U1983 : OAI21_X1 port map( A1 => n18702, A2 => n16352, B => n33736, ZN => 
                           n18431);
   U1984 : OAI21_X1 port map( A1 => n18866, A2 => n10283, B => n18871, ZN => 
                           n10220);
   U1985 : OAI21_X1 port map( A1 => n18112, A2 => n18672, B => n16572, ZN => 
                           n33324);
   U1988 : NOR2_X1 port map( A1 => n4259, A2 => n18768, ZN => n33799);
   U1992 : NAND2_X1 port map( A1 => n18510, A2 => n16352, ZN => n33736);
   U2009 : NOR2_X1 port map( A1 => n28009, A2 => n28010, ZN => n33559);
   U2013 : NAND2_X1 port map( A1 => n33997, A2 => n33999, ZN => n32763);
   U2015 : NAND2_X1 port map( A1 => n32411, A2 => n29309, ZN => n32410);
   U2016 : NOR2_X1 port map( A1 => n18603, A2 => n18602, ZN => n32491);
   U2019 : NAND3_X1 port map( A1 => n10043, A2 => n17255, A3 => n17223, ZN => 
                           n32294);
   U2021 : NAND3_X1 port map( A1 => n15108, A2 => n16881, A3 => n17255, ZN => 
                           n10561);
   U2022 : NAND2_X1 port map( A1 => n33999, A2 => n18672, ZN => n9289);
   U2023 : NOR2_X1 port map( A1 => n8400, A2 => n16614, ZN => n18859);
   U2027 : INV_X1 port map( I => n18228, ZN => n10903);
   U2032 : AND2_X1 port map( A1 => n29315, A2 => n18397, Z => n31986);
   U2039 : INV_X1 port map( I => n16995, ZN => n15406);
   U2046 : INV_X2 port map( I => n6860, ZN => n18854);
   U2054 : NOR2_X1 port map( A1 => n18702, A2 => n18510, ZN => n33792);
   U2055 : NOR2_X1 port map( A1 => n10325, A2 => n18677, ZN => n18679);
   U2057 : NAND2_X1 port map( A1 => n18738, A2 => n17166, ZN => n33207);
   U2063 : NAND2_X1 port map( A1 => n16287, A2 => n31417, ZN => n8860);
   U2066 : NAND2_X1 port map( A1 => n16372, A2 => n12863, ZN => n7497);
   U2067 : INV_X1 port map( I => n28245, ZN => n6359);
   U2074 : BUF_X2 port map( I => n18295, Z => n18324);
   U2079 : BUF_X2 port map( I => n18861, Z => n16287);
   U2080 : BUF_X2 port map( I => n34110, Z => n33093);
   U2084 : NAND2_X1 port map( A1 => n18006, A2 => n30271, ZN => n33040);
   U2088 : INV_X2 port map( I => n29309, ZN => n33989);
   U2093 : BUF_X2 port map( I => n32096, Z => n32798);
   U2094 : INV_X4 port map( I => n15716, ZN => n727);
   U2098 : NAND3_X1 port map( A1 => n18099, A2 => n15867, A3 => n6910, ZN => 
                           n28217);
   U2100 : NAND2_X2 port map( A1 => n22878, A2 => n23057, ZN => n22933);
   U2105 : NAND2_X2 port map( A1 => n27046, A2 => n25577, ZN => n33305);
   U2108 : NOR2_X2 port map( A1 => n123, A2 => n31327, ZN => n2656);
   U2112 : NAND3_X2 port map( A1 => n23177, A2 => n14350, A3 => n14756, ZN => 
                           n23178);
   U2118 : INV_X2 port map( I => n8778, ZN => n27150);
   U2120 : OAI22_X2 port map( A1 => n15284, A2 => n10472, B1 => n11072, B2 => 
                           n2081, ZN => n16909);
   U2130 : BUF_X4 port map( I => n24339, Z => n16552);
   U2132 : NAND3_X2 port map( A1 => n27833, A2 => n28917, A3 => n25609, ZN => 
                           n28156);
   U2136 : NAND2_X2 port map( A1 => n18261, A2 => n26739, ZN => n22860);
   U2137 : INV_X2 port map( I => n23746, ZN => n11392);
   U2139 : NOR2_X2 port map( A1 => n32855, A2 => n25615, ZN => n25607);
   U2141 : BUF_X2 port map( I => n23849, Z => n31435);
   U2144 : NOR2_X1 port map( A1 => n32301, A2 => n4607, ZN => n8653);
   U2147 : NAND2_X2 port map( A1 => n24262, A2 => n7809, ZN => n15974);
   U2152 : NOR2_X2 port map( A1 => n24104, A2 => n26750, ZN => n24102);
   U2153 : NOR2_X2 port map( A1 => n7093, A2 => n29566, ZN => n2853);
   U2155 : BUF_X4 port map( I => n2860, Z => n28957);
   U2156 : INV_X2 port map( I => n3181, ZN => n32186);
   U2158 : NOR2_X2 port map( A1 => n27651, A2 => n27461, ZN => n33643);
   U2159 : NAND2_X2 port map( A1 => n28181, A2 => n8140, ZN => n21460);
   U2160 : OR2_X2 port map( A1 => n4646, A2 => n31957, Z => n32079);
   U2163 : NAND2_X2 port map( A1 => n1015, A2 => n38, ZN => n8825);
   U2167 : INV_X4 port map( I => n28840, ZN => n26756);
   U2169 : INV_X2 port map( I => n25653, ZN => n734);
   U2172 : AND2_X2 port map( A1 => n30365, A2 => n22786, Z => n32088);
   U2173 : NAND3_X2 port map( A1 => n4436, A2 => n7810, A3 => n7680, ZN => 
                           n4591);
   U2175 : NAND2_X2 port map( A1 => n7093, A2 => n14839, ZN => n24344);
   U2182 : BUF_X2 port map( I => n7293, Z => n31957);
   U2189 : NAND2_X2 port map( A1 => n29634, A2 => n14619, ZN => n24153);
   U2190 : NAND2_X2 port map( A1 => n25452, A2 => n15212, ZN => n25430);
   U2191 : NAND2_X2 port map( A1 => n5820, A2 => n28957, ZN => n32712);
   U2194 : NAND3_X2 port map( A1 => n15580, A2 => n6553, A3 => n30364, ZN => 
                           n15579);
   U2196 : NOR2_X2 port map( A1 => n7116, A2 => n12184, ZN => n30148);
   U2197 : INV_X2 port map( I => n15051, ZN => n15060);
   U2199 : INV_X2 port map( I => n22033, ZN => n11727);
   U2204 : OAI22_X2 port map( A1 => n30934, A2 => n18567, B1 => n17316, B2 => 
                           n17813, ZN => n18423);
   U2206 : NAND2_X2 port map( A1 => n18423, A2 => n18493, ZN => n16806);
   U2207 : NAND2_X2 port map( A1 => n9620, A2 => n22377, ZN => n8176);
   U2208 : NAND2_X2 port map( A1 => n24251, A2 => n3220, ZN => n28827);
   U2209 : BUF_X4 port map( I => n23285, Z => n3868);
   U2212 : BUF_X4 port map( I => n12617, Z => n4774);
   U2213 : BUF_X2 port map( I => n15613, Z => n32975);
   U2214 : AND2_X1 port map( A1 => n9377, A2 => n23018, Z => n33862);
   U2216 : BUF_X2 port map( I => n31453, Z => n2391);
   U2217 : NOR2_X2 port map( A1 => n13712, A2 => n21251, ZN => n16204);
   U2219 : NAND2_X2 port map( A1 => n16387, A2 => n4216, ZN => n33044);
   U2220 : OAI21_X2 port map( A1 => n3731, A2 => n3732, B => n25236, ZN => 
                           n3730);
   U2222 : BUF_X2 port map( I => n32051, Z => n16389);
   U2224 : INV_X2 port map( I => n24269, ZN => n33891);
   U2225 : BUF_X2 port map( I => n8808, Z => n8301);
   U2227 : NOR2_X2 port map( A1 => n14752, A2 => n10099, ZN => n24904);
   U2228 : NAND2_X2 port map( A1 => n30252, A2 => n28069, ZN => n23750);
   U2229 : NAND2_X1 port map( A1 => n11597, A2 => n11596, ZN => n32739);
   U2235 : NOR3_X2 port map( A1 => n14463, A2 => n16496, A3 => n29965, ZN => 
                           n3445);
   U2236 : OAI21_X2 port map( A1 => n19165, A2 => n11085, B => n11444, ZN => 
                           n11474);
   U2238 : NOR2_X1 port map( A1 => n5304, A2 => n5305, ZN => n33385);
   U2240 : INV_X2 port map( I => n6402, ZN => n28200);
   U2244 : OAI21_X2 port map( A1 => n21434, A2 => n5049, B => n8010, ZN => 
                           n21074);
   U2248 : INV_X2 port map( I => n16809, ZN => n28658);
   U2249 : NOR2_X2 port map( A1 => n28408, A2 => n13762, ZN => n22861);
   U2250 : INV_X2 port map( I => n29213, ZN => n584);
   U2253 : NAND3_X1 port map( A1 => n32354, A2 => n7505, A3 => n7504, ZN => 
                           n24314);
   U2257 : OR2_X1 port map( A1 => n9159, A2 => n8602, Z => n25944);
   U2258 : BUF_X2 port map( I => n22579, Z => n16149);
   U2260 : AOI22_X2 port map( A1 => n1315, A2 => n33857, B1 => n8569, B2 => 
                           n5078, ZN => n5077);
   U2262 : NOR2_X2 port map( A1 => n34009, A2 => n34008, ZN => n6321);
   U2263 : OAI21_X2 port map( A1 => n33808, A2 => n29965, B => n28061, ZN => 
                           n33759);
   U2264 : NAND2_X2 port map( A1 => n1951, A2 => n25072, ZN => n10301);
   U2267 : NOR3_X1 port map( A1 => n33295, A2 => n30969, A3 => n24087, ZN => 
                           n14197);
   U2276 : NAND3_X1 port map( A1 => n2937, A2 => n8308, A3 => n23224, ZN => 
                           n2803);
   U2277 : INV_X1 port map( I => n23224, ZN => n26311);
   U2278 : CLKBUF_X4 port map( I => n20565, Z => n17329);
   U2280 : NOR2_X1 port map( A1 => n25681, A2 => n29243, ZN => n25682);
   U2289 : NAND2_X1 port map( A1 => n32879, A2 => n25675, ZN => n25681);
   U2296 : NAND2_X1 port map( A1 => n25002, A2 => n3229, ZN => n2266);
   U2297 : AOI21_X1 port map( A1 => n16127, A2 => n1134, B => n6074, ZN => 
                           n6678);
   U2306 : NAND2_X1 port map( A1 => n15217, A2 => n20608, ZN => n31714);
   U2310 : NOR2_X1 port map( A1 => n7290, A2 => n20608, ZN => n20186);
   U2311 : INV_X1 port map( I => n29815, ZN => n32951);
   U2312 : NAND2_X1 port map( A1 => n9646, A2 => n29815, ZN => n7575);
   U2319 : BUF_X2 port map( I => n28714, Z => n26133);
   U2320 : NOR2_X1 port map( A1 => n4041, A2 => n17313, ZN => n21158);
   U2322 : NAND2_X1 port map( A1 => n13579, A2 => n22033, ZN => n11728);
   U2328 : INV_X1 port map( I => n11205, ZN => n29927);
   U2332 : INV_X2 port map( I => n6593, ZN => n22956);
   U2335 : NOR2_X1 port map( A1 => n6593, A2 => n15601, ZN => n26047);
   U2344 : OAI21_X1 port map( A1 => n4918, A2 => n1294, B => n26884, ZN => 
                           n10611);
   U2346 : NAND2_X1 port map( A1 => n16964, A2 => n16963, ZN => n16962);
   U2347 : CLKBUF_X1 port map( I => n10285, Z => n28743);
   U2349 : AOI21_X1 port map( A1 => n22379, A2 => n33966, B => n636, ZN => 
                           n22380);
   U2351 : CLKBUF_X1 port map( I => n21079, Z => n32357);
   U2354 : NAND2_X1 port map( A1 => n11652, A2 => n11651, ZN => n8989);
   U2355 : NAND2_X1 port map( A1 => n28568, A2 => n857, ZN => n6062);
   U2356 : NAND2_X1 port map( A1 => n9028, A2 => n32583, ZN => n25176);
   U2361 : AOI21_X1 port map( A1 => n20112, A2 => n20113, B => n27808, ZN => 
                           n20116);
   U2362 : AOI22_X1 port map( A1 => n26787, A2 => n30230, B1 => n33624, B2 => 
                           n24337, ZN => n2401);
   U2365 : NOR2_X1 port map( A1 => n24244, A2 => n28374, ZN => n26787);
   U2369 : AOI22_X1 port map( A1 => n26367, A2 => n9370, B1 => n22503, B2 => 
                           n3332, ZN => n31162);
   U2375 : NOR2_X1 port map( A1 => n10202, A2 => n22503, ZN => n22404);
   U2376 : INV_X1 port map( I => n11898, ZN => n17781);
   U2378 : NOR3_X1 port map( A1 => n10931, A2 => n28131, A3 => n137, ZN => 
                           n2138);
   U2380 : AOI21_X1 port map( A1 => n30205, A2 => n11629, B => n28131, ZN => 
                           n16964);
   U2383 : OAI22_X1 port map( A1 => n14170, A2 => n25916, B1 => n25912, B2 => 
                           n25923, ZN => n14067);
   U2389 : AOI21_X1 port map( A1 => n1206, A2 => n25923, B => n690, ZN => 
                           n11156);
   U2392 : AOI21_X1 port map( A1 => n25909, A2 => n1206, B => n14067, ZN => 
                           n8394);
   U2393 : NAND2_X1 port map( A1 => n28743, A2 => n25743, ZN => n25734);
   U2398 : OAI22_X1 port map( A1 => n28743, A2 => n1597, B1 => n32863, B2 => 
                           n25746, ZN => n25750);
   U2399 : NOR2_X1 port map( A1 => n3019, A2 => n3229, ZN => n25005);
   U2400 : NAND2_X1 port map( A1 => n28639, A2 => n7862, ZN => n3208);
   U2401 : NOR2_X1 port map( A1 => n12861, A2 => n16688, ZN => n27662);
   U2402 : INV_X2 port map( I => n16688, ZN => n27661);
   U2403 : NAND2_X1 port map( A1 => n18204, A2 => n29498, ZN => n31266);
   U2409 : NAND2_X1 port map( A1 => n1086, A2 => n24220, ZN => n14445);
   U2410 : AOI21_X1 port map( A1 => n1086, A2 => n24220, B => n16688, ZN => 
                           n14447);
   U2411 : NAND2_X1 port map( A1 => n791, A2 => n24220, ZN => n12862);
   U2412 : NAND3_X1 port map( A1 => n25854, A2 => n14199, A3 => n10897, ZN => 
                           n15544);
   U2414 : INV_X1 port map( I => n21530, ZN => n33325);
   U2418 : OR2_X1 port map( A1 => n21530, A2 => n29980, Z => n31930);
   U2420 : NAND2_X1 port map( A1 => n15456, A2 => n3614, ZN => n22808);
   U2422 : NAND2_X1 port map( A1 => n15456, A2 => n12315, ZN => n15457);
   U2423 : NOR2_X1 port map( A1 => n1997, A2 => n1995, ZN => n24842);
   U2430 : INV_X2 port map( I => n700, ZN => n1223);
   U2433 : OAI21_X1 port map( A1 => n24249, A2 => n24248, B => n24250, ZN => 
                           n32976);
   U2434 : OAI22_X1 port map( A1 => n4070, A2 => n1182, B1 => n10713, B2 => 
                           n30472, ZN => n7493);
   U2437 : NAND2_X1 port map( A1 => n30651, A2 => n24207, ZN => n31160);
   U2445 : NAND2_X1 port map( A1 => n2427, A2 => n24030, ZN => n33963);
   U2450 : NAND2_X1 port map( A1 => n5611, A2 => n25236, ZN => n16400);
   U2451 : NAND2_X1 port map( A1 => n25236, A2 => n25234, ZN => n25133);
   U2458 : NOR2_X1 port map( A1 => n25875, A2 => n717, ZN => n13822);
   U2461 : CLKBUF_X1 port map( I => n7554, Z => n33702);
   U2466 : INV_X2 port map( I => n24150, ZN => n24317);
   U2469 : BUF_X1 port map( I => n25664, Z => n3883);
   U2470 : INV_X2 port map( I => n8370, ZN => n23892);
   U2472 : NOR2_X1 port map( A1 => n8370, A2 => n28266, ZN => n33827);
   U2474 : NAND2_X1 port map( A1 => n8370, A2 => n23894, ZN => n33829);
   U2475 : BUF_X2 port map( I => n8370, Z => n32434);
   U2476 : OAI22_X1 port map( A1 => n24737, A2 => n27162, B1 => n25836, B2 => 
                           n25860, ZN => n28887);
   U2477 : INV_X2 port map( I => n24909, ZN => n14752);
   U2478 : NAND2_X1 port map( A1 => n24205, A2 => n24204, ZN => n4519);
   U2479 : INV_X1 port map( I => n24205, ZN => n33549);
   U2481 : NAND2_X1 port map( A1 => n32328, A2 => n31160, ZN => n24205);
   U2486 : NAND2_X1 port map( A1 => n33543, A2 => n29056, ZN => n29520);
   U2487 : OAI21_X1 port map( A1 => n24260, A2 => n30280, B => n8248, ZN => 
                           n33543);
   U2489 : OAI21_X1 port map( A1 => n32872, A2 => n15641, B => n25184, ZN => 
                           n9192);
   U2490 : CLKBUF_X1 port map( I => n24779, Z => n32872);
   U2492 : NOR2_X1 port map( A1 => n24994, A2 => n5072, ZN => n26440);
   U2494 : NAND2_X1 port map( A1 => n24902, A2 => n10755, ZN => n24913);
   U2499 : INV_X1 port map( I => n10755, ZN => n24903);
   U2500 : AOI21_X1 port map( A1 => n16148, A2 => n22437, B => n14219, ZN => 
                           n4629);
   U2501 : INV_X1 port map( I => n3208, ZN => n32100);
   U2504 : AOI21_X1 port map( A1 => n26988, A2 => n6075, B => n30783, ZN => 
                           n2174);
   U2507 : NAND3_X1 port map( A1 => n5411, A2 => n11019, A3 => n1206, ZN => 
                           n25919);
   U2508 : OAI21_X1 port map( A1 => n6154, A2 => n14075, B => n24911, ZN => 
                           n8980);
   U2510 : INV_X1 port map( I => n9247, ZN => n25194);
   U2514 : NOR3_X1 port map( A1 => n32577, A2 => n27062, A3 => n14837, ZN => 
                           n8440);
   U2515 : NOR3_X1 port map( A1 => n15078, A2 => n15079, A3 => n42, ZN => 
                           n32577);
   U2525 : NAND2_X1 port map( A1 => n32611, A2 => n32609, ZN => n11670);
   U2527 : NAND2_X1 port map( A1 => n32531, A2 => n22944, ZN => n10108);
   U2531 : NOR2_X1 port map( A1 => n22944, A2 => n3657, ZN => n3659);
   U2532 : INV_X1 port map( I => n23171, ZN => n8068);
   U2533 : NOR2_X1 port map( A1 => n4193, A2 => n27668, ZN => n25097);
   U2536 : NAND2_X1 port map( A1 => n27668, A2 => n1203, ZN => n25088);
   U2539 : CLKBUF_X1 port map( I => n11360, Z => n27668);
   U2542 : NOR2_X1 port map( A1 => n24984, A2 => n14454, ZN => n16566);
   U2543 : OAI22_X1 port map( A1 => n24984, A2 => n3080, B1 => n1081, B2 => 
                           n27926, ZN => n17378);
   U2550 : NOR2_X1 port map( A1 => n24213, A2 => n26914, ZN => n342);
   U2551 : NAND2_X1 port map( A1 => n3376, A2 => n7831, ZN => n24988);
   U2552 : INV_X1 port map( I => n9963, ZN => n10296);
   U2556 : BUF_X2 port map( I => n9963, Z => n4750);
   U2557 : NAND3_X1 port map( A1 => n6713, A2 => n7891, A3 => n793, ZN => 
                           n24016);
   U2559 : NOR2_X1 port map( A1 => n8835, A2 => n23750, ZN => n23169);
   U2560 : NAND2_X1 port map( A1 => n15059, A2 => n15062, ZN => n15058);
   U2561 : AOI21_X1 port map( A1 => n5178, A2 => n23482, B => n22783, ZN => 
                           n5681);
   U2562 : AOI21_X1 port map( A1 => n25236, A2 => n25235, B => n1216, ZN => 
                           n4551);
   U2563 : NAND2_X1 port map( A1 => n25128, A2 => n15323, ZN => n25127);
   U2569 : AOI22_X1 port map( A1 => n18497, A2 => n19087, B1 => n19088, B2 => 
                           n28171, ZN => n18505);
   U2577 : NOR3_X1 port map( A1 => n33093, A2 => n14248, A3 => n33101, ZN => 
                           n29366);
   U2586 : BUF_X1 port map( I => n25228, Z => n28388);
   U2588 : CLKBUF_X4 port map( I => n11887, Z => n31807);
   U2591 : NOR3_X1 port map( A1 => n33583, A2 => n11887, A3 => n23942, ZN => 
                           n10020);
   U2592 : OR2_X1 port map( A1 => n3103, A2 => n16022, Z => n7626);
   U2598 : NAND2_X1 port map( A1 => n6491, A2 => n20517, ZN => n33240);
   U2601 : NAND2_X1 port map( A1 => n27267, A2 => n6336, ZN => n6334);
   U2603 : BUF_X2 port map( I => n3634, Z => n28239);
   U2604 : AND2_X1 port map( A1 => n15179, A2 => n2558, Z => n6772);
   U2605 : OAI21_X1 port map( A1 => n13560, A2 => n25587, B => n15964, ZN => 
                           n13559);
   U2606 : AOI21_X1 port map( A1 => n24631, A2 => n25587, B => n24633, ZN => 
                           n11824);
   U2612 : CLKBUF_X2 port map( I => n17306, Z => n31456);
   U2614 : NOR2_X1 port map( A1 => n28329, A2 => n26415, ZN => n2021);
   U2619 : NOR2_X1 port map( A1 => n2141, A2 => n24335, ZN => n33624);
   U2622 : INV_X1 port map( I => n16269, ZN => n910);
   U2629 : BUF_X2 port map( I => n16269, Z => n31105);
   U2633 : NAND3_X1 port map( A1 => n16269, A2 => n21680, A3 => n21681, ZN => 
                           n6570);
   U2635 : NAND2_X1 port map( A1 => n25229, A2 => n28388, ZN => n25261);
   U2643 : NOR3_X1 port map( A1 => n25227, A2 => n15705, A3 => n15738, ZN => 
                           n5532);
   U2647 : AOI21_X1 port map( A1 => n33900, A2 => n10608, B => n733, ZN => 
                           n10606);
   U2649 : NAND3_X1 port map( A1 => n733, A2 => n25278, A3 => n28532, ZN => 
                           n24590);
   U2652 : NAND2_X1 port map( A1 => n24262, A2 => n3205, ZN => n8248);
   U2654 : NAND2_X1 port map( A1 => n32859, A2 => n5713, ZN => n28639);
   U2656 : CLKBUF_X2 port map( I => n20994, Z => n28687);
   U2657 : INV_X1 port map( I => n20994, ZN => n1339);
   U2662 : NAND2_X1 port map( A1 => n28752, A2 => n17974, ZN => n20994);
   U2663 : NOR2_X1 port map( A1 => n14386, A2 => n24044, ZN => n14249);
   U2664 : NAND3_X1 port map( A1 => n25346, A2 => n24506, A3 => n753, ZN => 
                           n10330);
   U2665 : AOI22_X1 port map( A1 => n25732, A2 => n33386, B1 => n25730, B2 => 
                           n25731, ZN => n32508);
   U2667 : NAND2_X1 port map( A1 => n31941, A2 => n11704, ZN => n24588);
   U2680 : OAI21_X1 port map( A1 => n31941, A2 => n25392, B => n13993, ZN => 
                           n25442);
   U2686 : BUF_X2 port map( I => n28632, Z => n31229);
   U2689 : NOR2_X1 port map( A1 => n9181, A2 => n25820, ZN => n25807);
   U2691 : NAND2_X1 port map( A1 => n221, A2 => n13617, ZN => n25569);
   U2692 : INV_X1 port map( I => n13617, ZN => n6111);
   U2693 : NAND2_X1 port map( A1 => n13617, A2 => n691, ZN => n27046);
   U2696 : NAND2_X1 port map( A1 => n13617, A2 => n8168, ZN => n25568);
   U2701 : NAND2_X1 port map( A1 => n33894, A2 => n6319, ZN => n5089);
   U2705 : NOR2_X1 port map( A1 => n33894, A2 => n6319, ZN => n32526);
   U2706 : CLKBUF_X4 port map( I => n24471, Z => n25013);
   U2708 : NOR2_X1 port map( A1 => n419, A2 => n25405, ZN => n25328);
   U2710 : NAND2_X1 port map( A1 => n14810, A2 => n6402, ZN => n25124);
   U2711 : NAND3_X1 port map( A1 => n17872, A2 => n5373, A3 => n23901, ZN => 
                           n17995);
   U2713 : NAND2_X1 port map( A1 => n17149, A2 => n3898, ZN => n5136);
   U2721 : CLKBUF_X2 port map( I => n25369, Z => n30400);
   U2722 : NOR2_X1 port map( A1 => n13883, A2 => n13811, ZN => n25559);
   U2724 : BUF_X2 port map( I => n7925, Z => n34109);
   U2730 : INV_X1 port map( I => n7925, ZN => n3646);
   U2731 : OAI22_X1 port map( A1 => n6061, A2 => n2697, B1 => n6062, B2 => 
                           n16647, ZN => n33634);
   U2736 : NAND2_X1 port map( A1 => n1805, A2 => n16647, ZN => n6061);
   U2739 : NAND2_X1 port map( A1 => n31155, A2 => n30505, ZN => n31837);
   U2742 : NAND2_X1 port map( A1 => n1090, A2 => n31155, ZN => n10812);
   U2743 : BUF_X1 port map( I => n14531, Z => n32553);
   U2746 : NOR2_X1 port map( A1 => n25632, A2 => n29476, ZN => n30423);
   U2747 : NOR3_X1 port map( A1 => n30396, A2 => n10314, A3 => n14922, ZN => 
                           n26528);
   U2748 : OAI21_X1 port map( A1 => n33680, A2 => n33540, B => n24243, ZN => 
                           n23984);
   U2752 : NAND3_X1 port map( A1 => n29495, A2 => n1127, A3 => n22670, ZN => 
                           n33015);
   U2757 : INV_X1 port map( I => n23840, ZN => n32611);
   U2761 : OAI21_X1 port map( A1 => n13242, A2 => n23935, B => n15097, ZN => 
                           n14704);
   U2763 : NAND3_X1 port map( A1 => n13242, A2 => n23575, A3 => n17181, ZN => 
                           n33625);
   U2764 : OAI21_X1 port map( A1 => n31959, A2 => n23935, B => n13242, ZN => 
                           n28530);
   U2765 : NAND2_X1 port map( A1 => n31959, A2 => n13242, ZN => n15803);
   U2769 : INV_X1 port map( I => n4034, ZN => n1309);
   U2773 : NOR2_X1 port map( A1 => n1500, A2 => n24072, ZN => n1499);
   U2774 : BUF_X2 port map( I => n24072, Z => n27038);
   U2776 : AOI21_X1 port map( A1 => n25858, A2 => n14915, B => n25854, ZN => 
                           n24737);
   U2777 : NAND2_X1 port map( A1 => n25858, A2 => n25859, ZN => n25857);
   U2779 : NAND2_X1 port map( A1 => n13947, A2 => n13946, ZN => n13945);
   U2781 : INV_X1 port map( I => n11668, ZN => n29660);
   U2782 : NAND3_X1 port map( A1 => n23543, A2 => n23855, A3 => n14193, ZN => 
                           n23547);
   U2785 : NAND2_X1 port map( A1 => n5897, A2 => n17382, ZN => n24984);
   U2787 : INV_X1 port map( I => n17382, ZN => n13428);
   U2788 : NOR2_X1 port map( A1 => n25460, A2 => n25475, ZN => n32115);
   U2789 : CLKBUF_X2 port map( I => n25107, Z => n4193);
   U2792 : NOR2_X1 port map( A1 => n23857, A2 => n23201, ZN => n25951);
   U2795 : NOR2_X1 port map( A1 => n23201, A2 => n9152, ZN => n29178);
   U2797 : CLKBUF_X2 port map( I => n25859, Z => n13049);
   U2800 : AND2_X1 port map( A1 => n25513, A2 => n25517, Z => n25516);
   U2806 : OAI21_X1 port map( A1 => n25081, A2 => n30330, B => n32771, ZN => 
                           n16104);
   U2811 : AOI22_X1 port map( A1 => n1949, A2 => n30330, B1 => n1951, B2 => 
                           n16810, ZN => n32771);
   U2819 : AOI21_X1 port map( A1 => n25923, A2 => n25915, B => n11019, ZN => 
                           n14432);
   U2820 : CLKBUF_X4 port map( I => n13960, Z => n11019);
   U2828 : NOR2_X1 port map( A1 => n28694, A2 => n24004, ZN => n5912);
   U2829 : OAI21_X1 port map( A1 => n33871, A2 => n33872, B => n24004, ZN => 
                           n8001);
   U2832 : INV_X2 port map( I => n16273, ZN => n8929);
   U2834 : AOI22_X1 port map( A1 => n8207, A2 => n16273, B1 => n33851, B2 => 
                           n25174, ZN => n25180);
   U2835 : INV_X1 port map( I => n3220, ZN => n24069);
   U2837 : AOI21_X1 port map( A1 => n24249, A2 => n24248, B => n3220, ZN => 
                           n29949);
   U2843 : NAND2_X1 port map( A1 => n13223, A2 => n3220, ZN => n1511);
   U2844 : INV_X1 port map( I => n5043, ZN => n25211);
   U2851 : AOI21_X1 port map( A1 => n1186, A2 => n18701, B => n31012, ZN => 
                           n13947);
   U2854 : NAND3_X1 port map( A1 => n1186, A2 => n34110, A3 => n18701, ZN => 
                           n33412);
   U2861 : INV_X2 port map( I => n18701, ZN => n13554);
   U2862 : OAI22_X1 port map( A1 => n32100, A2 => n25090, B1 => n25094, B2 => 
                           n25089, ZN => n32529);
   U2863 : CLKBUF_X2 port map( I => n8678, Z => n26753);
   U2865 : NOR2_X1 port map( A1 => n8678, A2 => n25795, ZN => n25797);
   U2875 : AND2_X1 port map( A1 => n25317, A2 => n25313, Z => n25320);
   U2877 : NAND4_X1 port map( A1 => n693, A2 => n25070, A3 => n25069, A4 => 
                           n25068, ZN => n29723);
   U2878 : INV_X1 port map( I => n7198, ZN => n747);
   U2881 : OAI21_X1 port map( A1 => n32270, A2 => n34170, B => n24897, ZN => 
                           n33081);
   U2882 : CLKBUF_X2 port map( I => n16940, Z => n4024);
   U2884 : INV_X1 port map( I => n16940, ZN => n24311);
   U2886 : NAND3_X1 port map( A1 => n25744, A2 => n25739, A3 => n4415, ZN => 
                           n32279);
   U2887 : INV_X1 port map( I => n1506, ZN => n8235);
   U2888 : NAND2_X1 port map( A1 => n4778, A2 => n4776, ZN => n3589);
   U2890 : NOR3_X1 port map( A1 => n8258, A2 => n16377, A3 => n8257, ZN => 
                           n28486);
   U2891 : OR2_X1 port map( A1 => n25473, A2 => n30047, Z => n25460);
   U2893 : INV_X2 port map( I => n30584, ZN => n16501);
   U2895 : NAND2_X1 port map( A1 => n3909, A2 => n30584, ZN => n22744);
   U2904 : NOR2_X1 port map( A1 => n22953, A2 => n30584, ZN => n22327);
   U2911 : NAND2_X1 port map( A1 => n11105, A2 => n20591, ZN => n11104);
   U2912 : NAND2_X1 port map( A1 => n11255, A2 => n24327, ZN => n9823);
   U2913 : NAND3_X1 port map( A1 => n32510, A2 => n22855, A3 => n25979, ZN => 
                           n22859);
   U2914 : NOR2_X1 port map( A1 => n22709, A2 => n25979, ZN => n14162);
   U2927 : NAND3_X1 port map( A1 => n25979, A2 => n33132, A3 => n30365, ZN => 
                           n22857);
   U2931 : AOI21_X1 port map( A1 => n2480, A2 => n749, B => n32177, ZN => 
                           n25504);
   U2932 : CLKBUF_X2 port map( I => n6595, Z => n2480);
   U2937 : NAND2_X1 port map( A1 => n28427, A2 => n12471, ZN => n10361);
   U2940 : NAND2_X1 port map( A1 => n18084, A2 => n26390, ZN => n24709);
   U2941 : NOR2_X1 port map( A1 => n26390, A2 => n24310, ZN => n9016);
   U2942 : NAND2_X1 port map( A1 => n16609, A2 => n718, ZN => n25583);
   U2943 : INV_X1 port map( I => n16609, ZN => n13642);
   U2946 : NAND3_X1 port map( A1 => n27113, A2 => n6092, A3 => n5926, ZN => n36
                           );
   U2947 : CLKBUF_X4 port map( I => n5492, Z => n964);
   U2949 : NAND2_X1 port map( A1 => n13488, A2 => n19867, ZN => n28130);
   U2952 : NOR2_X1 port map( A1 => n16271, A2 => n33679, ZN => n33870);
   U2956 : NAND2_X1 port map( A1 => n5091, A2 => n5292, ZN => n24728);
   U2957 : INV_X1 port map( I => n10644, ZN => n23064);
   U2962 : NOR2_X1 port map( A1 => n714, A2 => n25006, ZN => n15079);
   U2963 : NOR2_X1 port map( A1 => n16519, A2 => n21662, ZN => n13213);
   U2966 : NOR2_X1 port map( A1 => n16519, A2 => n32898, ZN => n14730);
   U2968 : NAND3_X1 port map( A1 => n777, A2 => n21662, A3 => n16519, ZN => 
                           n27760);
   U2972 : AOI21_X1 port map( A1 => n7068, A2 => n24196, B => n28784, ZN => 
                           n2921);
   U2973 : NAND2_X1 port map( A1 => n25724, A2 => n16494, ZN => n25717);
   U2974 : OR2_X1 port map( A1 => n675, A2 => n24779, Z => n2727);
   U2982 : CLKBUF_X2 port map( I => n7940, Z => n3376);
   U2984 : NAND2_X1 port map( A1 => n25882, A2 => n5410, ZN => n33176);
   U2994 : CLKBUF_X2 port map( I => n17824, Z => n30396);
   U2995 : AOI21_X1 port map( A1 => n14922, A2 => n17824, B => n6034, ZN => 
                           n16169);
   U2997 : NAND2_X1 port map( A1 => n7515, A2 => n25221, ZN => n15462);
   U2998 : INV_X1 port map( I => n25221, ZN => n966);
   U3000 : NAND2_X1 port map( A1 => n15421, A2 => n22832, ZN => n23002);
   U3001 : OAI21_X1 port map( A1 => n22752, A2 => n15421, B => n16817, ZN => 
                           n22618);
   U3003 : AND2_X1 port map( A1 => n14873, A2 => n33155, Z => n32030);
   U3007 : NOR2_X1 port map( A1 => n13296, A2 => n13822, ZN => n33516);
   U3011 : OAI21_X1 port map( A1 => n10206, A2 => n28263, B => n6709, ZN => 
                           n6711);
   U3014 : OAI21_X1 port map( A1 => n22583, A2 => n10206, B => n28263, ZN => 
                           n10796);
   U3015 : NAND2_X1 port map( A1 => n33392, A2 => n6661, ZN => n30185);
   U3016 : NAND2_X1 port map( A1 => n16292, A2 => n23759, ZN => n33392);
   U3018 : NAND2_X1 port map( A1 => n31323, A2 => n32144, ZN => n32272);
   U3023 : AOI22_X1 port map( A1 => n25552, A2 => n13483, B1 => n33414, B2 => 
                           n13811, ZN => n32144);
   U3024 : OAI21_X1 port map( A1 => n16835, A2 => n700, B => n25900, ZN => 
                           n10756);
   U3033 : NAND3_X1 port map( A1 => n13366, A2 => n8657, A3 => n13367, ZN => 
                           n31734);
   U3042 : NAND2_X1 port map( A1 => n7831, A2 => n24995, ZN => n14208);
   U3046 : BUF_X2 port map( I => n14058, Z => n27750);
   U3047 : NAND2_X1 port map( A1 => n31907, A2 => n20507, ZN => n14683);
   U3049 : AND2_X1 port map( A1 => n3944, A2 => n31907, Z => n16123);
   U3051 : INV_X1 port map( I => n31907, ZN => n14369);
   U3054 : INV_X1 port map( I => n23456, ZN => n30843);
   U3059 : BUF_X2 port map( I => n23456, Z => n27481);
   U3061 : INV_X1 port map( I => n15425, ZN => n25865);
   U3062 : INV_X1 port map( I => n21012, ZN => n30487);
   U3063 : NAND2_X1 port map( A1 => n22772, A2 => n1106, ZN => n22773);
   U3066 : AND2_X1 port map( A1 => n24171, A2 => n3483, Z => n32041);
   U3067 : NAND2_X1 port map( A1 => n34149, A2 => n834, ZN => n12386);
   U3068 : INV_X1 port map( I => n834, ZN => n32591);
   U3070 : CLKBUF_X2 port map( I => n18911, Z => n33698);
   U3071 : NAND3_X1 port map( A1 => n34074, A2 => n29395, A3 => n22682, ZN => 
                           n3894);
   U3072 : NAND2_X1 port map( A1 => n22772, A2 => n28957, ZN => n22751);
   U3073 : NAND2_X1 port map( A1 => n3300, A2 => n25375, ZN => n25366);
   U3074 : NOR2_X1 port map( A1 => n25376, A2 => n25375, ZN => n14102);
   U3075 : NAND2_X1 port map( A1 => n21840, A2 => n16987, ZN => n21749);
   U3080 : NOR2_X1 port map( A1 => n32063, A2 => n24955, ZN => n24948);
   U3081 : CLKBUF_X4 port map( I => n24174, Z => n25900);
   U3084 : NAND2_X1 port map( A1 => n11899, A2 => n8307, ZN => n24710);
   U3085 : OAI21_X1 port map( A1 => n696, A2 => n1212, B => n11899, ZN => n4709
                           );
   U3092 : NOR2_X1 port map( A1 => n1202, A2 => n9982, ZN => n12049);
   U3093 : INV_X1 port map( I => n32906, ZN => n23152);
   U3094 : AOI22_X1 port map( A1 => n33176, A2 => n14737, B1 => n5407, B2 => 
                           n32059, ZN => n13902);
   U3096 : AND2_X1 port map( A1 => n16033, A2 => n17661, Z => n1933);
   U3097 : NAND2_X1 port map( A1 => n1100, A2 => n16033, ZN => n7781);
   U3099 : INV_X1 port map( I => n535, ZN => n16033);
   U3104 : INV_X1 port map( I => n16853, ZN => n28759);
   U3106 : NAND2_X1 port map( A1 => n5259, A2 => n12450, ZN => n12449);
   U3107 : INV_X1 port map( I => n23334, ZN => n31567);
   U3109 : NAND2_X1 port map( A1 => n30033, A2 => n8875, ZN => n21740);
   U3110 : CLKBUF_X4 port map( I => n24408, Z => n25756);
   U3121 : NOR2_X1 port map( A1 => n22546, A2 => n22550, ZN => n27406);
   U3122 : OAI21_X1 port map( A1 => n22546, A2 => n27402, B => n22550, ZN => 
                           n26855);
   U3123 : NOR3_X1 port map( A1 => n22546, A2 => n22549, A3 => n22547, ZN => 
                           n32943);
   U3128 : INV_X1 port map( I => n24275, ZN => n24196);
   U3130 : NOR2_X1 port map( A1 => n30129, A2 => n33766, ZN => n16229);
   U3134 : OAI21_X1 port map( A1 => n912, A2 => n33766, B => n1137, ZN => n2718
                           );
   U3136 : NAND2_X1 port map( A1 => n33766, A2 => n2368, ZN => n33841);
   U3137 : AOI21_X1 port map( A1 => n912, A2 => n33766, B => n38, ZN => n16231)
                           ;
   U3142 : NAND2_X1 port map( A1 => n25141, A2 => n25145, ZN => n2642);
   U3143 : CLKBUF_X2 port map( I => n25141, Z => n16276);
   U3151 : INV_X1 port map( I => n25141, ZN => n17987);
   U3154 : NAND2_X1 port map( A1 => n31915, A2 => n11850, ZN => n10470);
   U3158 : CLKBUF_X2 port map( I => n3874, Z => n29839);
   U3159 : NAND2_X1 port map( A1 => n27670, A2 => n22653, ZN => n3951);
   U3163 : AOI22_X1 port map( A1 => n16560, A2 => n22826, B1 => n23066, B2 => 
                           n7881, ZN => n22653);
   U3164 : NAND2_X1 port map( A1 => n23064, A2 => n28689, ZN => n27670);
   U3165 : INV_X2 port map( I => n19907, ZN => n20112);
   U3166 : NAND2_X1 port map( A1 => n16058, A2 => n21396, ZN => n27432);
   U3168 : NOR2_X1 port map( A1 => n12325, A2 => n21396, ZN => n12324);
   U3171 : NOR3_X1 port map( A1 => n21396, A2 => n27955, A3 => n21400, ZN => 
                           n32393);
   U3174 : NAND2_X1 port map( A1 => n15746, A2 => n16205, ZN => n3598);
   U3185 : NAND2_X1 port map( A1 => n22690, A2 => n15746, ZN => n32191);
   U3194 : NOR2_X1 port map( A1 => n22690, A2 => n15746, ZN => n30436);
   U3201 : NAND2_X1 port map( A1 => n15746, A2 => n30333, ZN => n31126);
   U3202 : NOR2_X1 port map( A1 => n25967, A2 => n10700, ZN => n15804);
   U3205 : NOR2_X1 port map( A1 => n32186, A2 => n7188, ZN => n9788);
   U3206 : NOR2_X1 port map( A1 => n3165, A2 => n32186, ZN => n34012);
   U3207 : INV_X1 port map( I => n12648, ZN => n32785);
   U3209 : CLKBUF_X2 port map( I => n9107, Z => n26739);
   U3211 : OR2_X1 port map( A1 => n4184, A2 => n13191, Z => n31052);
   U3212 : NAND2_X1 port map( A1 => n4184, A2 => n13191, ZN => n13995);
   U3213 : AND2_X1 port map( A1 => n2635, A2 => n4184, Z => n8290);
   U3214 : CLKBUF_X2 port map( I => n9708, Z => n29318);
   U3216 : CLKBUF_X2 port map( I => n16331, Z => n8347);
   U3217 : BUF_X2 port map( I => n21071, Z => n21426);
   U3218 : OR2_X1 port map( A1 => n17670, A2 => n5433, Z => n29357);
   U3219 : NAND2_X1 port map( A1 => n7081, A2 => n25232, ZN => n10570);
   U3220 : OR2_X1 port map( A1 => n339, A2 => n31217, Z => n18344);
   U3224 : NOR2_X1 port map( A1 => n32401, A2 => n339, ZN => n9839);
   U3228 : INV_X2 port map( I => n339, ZN => n19052);
   U3229 : AOI21_X1 port map( A1 => n32401, A2 => n339, B => n10015, ZN => 
                           n2148);
   U3230 : OAI21_X1 port map( A1 => n339, A2 => n10015, B => n10017, ZN => 
                           n31226);
   U3231 : OR3_X2 port map( A1 => n989, A2 => n12578, A3 => n13648, Z => n12577
                           );
   U3232 : INV_X1 port map( I => n33857, ZN => n33519);
   U3236 : NAND2_X1 port map( A1 => n18830, A2 => n16915, ZN => n3893);
   U3239 : AOI21_X1 port map( A1 => n18830, A2 => n9, B => n18829, ZN => n29808
                           );
   U3244 : INV_X1 port map( I => n3079, ZN => n32565);
   U3245 : NAND2_X1 port map( A1 => n10724, A2 => n906, ZN => n4315);
   U3246 : AOI22_X1 port map( A1 => n22643, A2 => n30448, B1 => n6297, B2 => 
                           n10724, ZN => n13461);
   U3247 : INV_X1 port map( I => n19470, ZN => n19561);
   U3249 : AND2_X1 port map( A1 => n11515, A2 => n30713, Z => n31180);
   U3255 : OAI21_X1 port map( A1 => n867, A2 => n1469, B => n20442, ZN => 
                           n30929);
   U3260 : NAND2_X1 port map( A1 => n19932, A2 => n8817, ZN => n1812);
   U3268 : NAND2_X1 port map( A1 => n11903, A2 => n2166, ZN => n2167);
   U3270 : NAND2_X1 port map( A1 => n2166, A2 => n28645, ZN => n28022);
   U3272 : OAI21_X1 port map( A1 => n2166, A2 => n20069, B => n27715, ZN => 
                           n6926);
   U3276 : INV_X1 port map( I => n32124, ZN => n297);
   U3282 : BUF_X2 port map( I => Key(57), Z => n25856);
   U3285 : NOR2_X1 port map( A1 => n5098, A2 => n24111, ZN => n10178);
   U3286 : NAND2_X1 port map( A1 => n13896, A2 => n16072, ZN => n14074);
   U3288 : OAI22_X1 port map( A1 => n4989, A2 => n4324, B1 => n13896, B2 => 
                           n32799, ZN => n30654);
   U3289 : CLKBUF_X4 port map( I => n24866, Z => n24667);
   U3292 : OAI22_X1 port map( A1 => n803, A2 => n27450, B1 => n23158, B2 => 
                           n14183, ZN => n27372);
   U3295 : OAI21_X1 port map( A1 => n3379, A2 => n11756, B => n31197, ZN => 
                           n13034);
   U3300 : NAND2_X1 port map( A1 => n31197, A2 => n28099, ZN => n21664);
   U3303 : OAI21_X1 port map( A1 => n15038, A2 => n16099, B => n31479, ZN => 
                           n5040);
   U3306 : BUF_X2 port map( I => n8926, Z => n8207);
   U3310 : NOR2_X1 port map( A1 => n25154, A2 => n8926, ZN => n25158);
   U3314 : INV_X1 port map( I => n8926, ZN => n25165);
   U3317 : NAND3_X1 port map( A1 => n15423, A2 => n23848, A3 => n26114, ZN => 
                           n6129);
   U3318 : INV_X1 port map( I => n30305, ZN => n19416);
   U3320 : INV_X1 port map( I => n24573, ZN => n11652);
   U3323 : NAND3_X1 port map( A1 => n24573, A2 => n14410, A3 => n14412, ZN => 
                           n8988);
   U3324 : CLKBUF_X2 port map( I => n21569, Z => n29806);
   U3327 : INV_X1 port map( I => n21569, ZN => n32506);
   U3330 : NAND2_X1 port map( A1 => n3203, A2 => n21569, ZN => n21491);
   U3333 : CLKBUF_X2 port map( I => n8622, Z => n33434);
   U3335 : NAND3_X1 port map( A1 => n21865, A2 => n30154, A3 => n28018, ZN => 
                           n21739);
   U3339 : AOI22_X1 port map( A1 => n26766, A2 => n8457, B1 => n21865, B2 => 
                           n21867, ZN => n4516);
   U3350 : NAND2_X1 port map( A1 => n21865, A2 => n21866, ZN => n16241);
   U3352 : NAND2_X1 port map( A1 => n32833, A2 => n21865, ZN => n31711);
   U3353 : NOR2_X1 port map( A1 => n21865, A2 => n21866, ZN => n31334);
   U3355 : INV_X2 port map( I => n21865, ZN => n15465);
   U3356 : CLKBUF_X2 port map( I => n22363, Z => n6478);
   U3357 : CLKBUF_X4 port map( I => n16052, Z => n5631);
   U3358 : INV_X2 port map( I => n16052, ZN => n5632);
   U3364 : NAND3_X1 port map( A1 => n4873, A2 => n23934, A3 => n11200, ZN => 
                           n4872);
   U3366 : NOR3_X1 port map( A1 => n33425, A2 => n28945, A3 => n11200, ZN => 
                           n32929);
   U3367 : NAND3_X1 port map( A1 => n27450, A2 => n32868, A3 => n803, ZN => 
                           n13914);
   U3372 : NOR2_X1 port map( A1 => n23051, A2 => n28277, ZN => n17482);
   U3378 : NOR2_X1 port map( A1 => n28277, A2 => n23051, ZN => n16054);
   U3381 : CLKBUF_X4 port map( I => n19418, Z => n19884);
   U3383 : NOR2_X1 port map( A1 => n19418, A2 => n19885, ZN => n13488);
   U3384 : CLKBUF_X4 port map( I => n2600, Z => n29330);
   U3388 : INV_X1 port map( I => n5268, ZN => n3146);
   U3397 : NOR3_X1 port map( A1 => n29634, A2 => n14619, A3 => n24154, ZN => 
                           n5613);
   U3399 : NOR2_X1 port map( A1 => n9062, A2 => n31471, ZN => n14568);
   U3407 : NAND2_X1 port map( A1 => n9062, A2 => n20630, ZN => n31469);
   U3408 : NOR3_X1 port map( A1 => n5335, A2 => n24148, A3 => n3748, ZN => 
                           n8543);
   U3409 : CLKBUF_X4 port map( I => n29279, Z => n33585);
   U3413 : NAND2_X1 port map( A1 => n25755, A2 => n29279, ZN => n32343);
   U3415 : NAND2_X1 port map( A1 => n31079, A2 => n30504, ZN => n30503);
   U3418 : NAND2_X1 port map( A1 => n15314, A2 => n15316, ZN => n30284);
   U3420 : NOR2_X1 port map( A1 => n23849, A2 => n26114, ZN => n23808);
   U3421 : AOI22_X1 port map( A1 => n12996, A2 => n100, B1 => n19057, B2 => 
                           n19058, ZN => n19059);
   U3425 : NAND2_X1 port map( A1 => n6718, A2 => n21719, ZN => n14717);
   U3427 : NAND2_X1 port map( A1 => n12221, A2 => n6718, ZN => n21741);
   U3429 : INV_X1 port map( I => n6718, ZN => n33083);
   U3431 : NAND2_X1 port map( A1 => n17227, A2 => n6718, ZN => n3420);
   U3444 : OR2_X1 port map( A1 => n13913, A2 => n29815, Z => n5223);
   U3452 : NAND2_X1 port map( A1 => n24960, A2 => n24896, ZN => n24939);
   U3456 : NOR2_X1 port map( A1 => n8420, A2 => n29287, ZN => n22683);
   U3458 : INV_X1 port map( I => n8420, ZN => n2418);
   U3459 : NAND2_X1 port map( A1 => n25012, A2 => n25015, ZN => n24591);
   U3466 : NOR2_X1 port map( A1 => n30145, A2 => n25015, ZN => n33757);
   U3469 : NOR2_X1 port map( A1 => n25015, A2 => n17240, ZN => n12093);
   U3471 : INV_X2 port map( I => n24975, ZN => n25015);
   U3472 : NOR2_X1 port map( A1 => n33648, A2 => n29387, ZN => n26389);
   U3473 : AOI21_X1 port map( A1 => n12657, A2 => n20066, B => n19874, ZN => 
                           n19798);
   U3476 : AOI21_X1 port map( A1 => n14976, A2 => n12657, B => n20066, ZN => 
                           n29905);
   U3478 : INV_X1 port map( I => n29258, ZN => n17053);
   U3482 : INV_X1 port map( I => n3147, ZN => n11768);
   U3484 : BUF_X2 port map( I => n3147, Z => n31228);
   U3491 : NAND2_X1 port map( A1 => n21072, A2 => n21428, ZN => n2241);
   U3495 : NAND2_X1 port map( A1 => n20009, A2 => n20008, ZN => n20085);
   U3496 : NAND3_X1 port map( A1 => n20009, A2 => n8301, A3 => n20008, ZN => 
                           n9338);
   U3499 : OR3_X2 port map( A1 => n20009, A2 => n20083, A3 => n11068, Z => 
                           n9339);
   U3501 : CLKBUF_X2 port map( I => n22457, Z => n16503);
   U3505 : INV_X2 port map( I => n12535, ZN => n26513);
   U3506 : INV_X1 port map( I => n12548, ZN => n18978);
   U3511 : NOR2_X1 port map( A1 => n16916, A2 => n12548, ZN => n6639);
   U3516 : NAND2_X1 port map( A1 => n12548, A2 => n14812, ZN => n19113);
   U3521 : CLKBUF_X1 port map( I => n17408, Z => n27984);
   U3523 : CLKBUF_X2 port map( I => n13694, Z => n27450);
   U3524 : NAND2_X1 port map( A1 => n1177, A2 => n32332, ZN => n32331);
   U3530 : INV_X2 port map( I => n1177, ZN => n32671);
   U3534 : AOI21_X1 port map( A1 => n19324, A2 => n19274, B => n1177, ZN => 
                           n19278);
   U3537 : OAI21_X1 port map( A1 => n29965, A2 => n23912, B => n23588, ZN => 
                           n16539);
   U3542 : OAI21_X1 port map( A1 => n16496, A2 => n34167, B => n29965, ZN => 
                           n28061);
   U3545 : NAND2_X1 port map( A1 => n16496, A2 => n29965, ZN => n26224);
   U3546 : INV_X2 port map( I => n20523, ZN => n17790);
   U3552 : NAND2_X1 port map( A1 => n30454, A2 => n20523, ZN => n28484);
   U3555 : NOR2_X1 port map( A1 => n16684, A2 => n20523, ZN => n20280);
   U3556 : OAI21_X1 port map( A1 => n16459, A2 => n31195, B => n31498, ZN => 
                           n2687);
   U3558 : OAI21_X1 port map( A1 => n16459, A2 => n926, B => n21077, ZN => 
                           n12506);
   U3561 : NAND2_X1 port map( A1 => n33523, A2 => n16459, ZN => n2569);
   U3562 : BUF_X2 port map( I => n16248, Z => n28904);
   U3568 : INV_X1 port map( I => n16248, ZN => n26182);
   U3575 : BUF_X2 port map( I => n18064, Z => n29216);
   U3576 : NAND2_X1 port map( A1 => n18064, A2 => n34122, ZN => n33570);
   U3580 : INV_X1 port map( I => n18064, ZN => n1035);
   U3591 : OR2_X1 port map( A1 => n10514, A2 => n18064, Z => n29022);
   U3595 : CLKBUF_X1 port map( I => n16215, Z => n10651);
   U3596 : INV_X1 port map( I => n16215, ZN => n29883);
   U3599 : AND2_X1 port map( A1 => n7935, A2 => n16215, Z => n9368);
   U3600 : NOR2_X1 port map( A1 => n16389, A2 => n28578, ZN => n18671);
   U3601 : NOR3_X1 port map( A1 => n16466, A2 => n16572, A3 => n16389, ZN => 
                           n10638);
   U3608 : NAND2_X1 port map( A1 => n31437, A2 => n23057, ZN => n2877);
   U3615 : INV_X2 port map( I => n14359, ZN => n1206);
   U3619 : NAND2_X1 port map( A1 => n14359, A2 => n7702, ZN => n25912);
   U3621 : CLKBUF_X2 port map( I => n24447, Z => n16413);
   U3622 : NAND2_X1 port map( A1 => n15116, A2 => n23742, ZN => n23583);
   U3630 : OAI21_X1 port map( A1 => n20460, A2 => n7852, B => n7292, ZN => 
                           n31898);
   U3631 : BUF_X2 port map( I => n7852, Z => n8031);
   U3636 : INV_X1 port map( I => n16175, ZN => n14968);
   U3640 : OAI21_X1 port map( A1 => n34115, A2 => n1216, B => n1083, ZN => 
                           n8120);
   U3653 : NOR2_X1 port map( A1 => n25234, A2 => n1083, ZN => n3731);
   U3655 : INV_X2 port map( I => n34167, ZN => n14463);
   U3658 : AOI21_X1 port map( A1 => n2507, A2 => n10283, B => n32409, ZN => 
                           n32541);
   U3664 : INV_X1 port map( I => n19967, ZN => n14334);
   U3668 : CLKBUF_X2 port map( I => n19967, Z => n16092);
   U3677 : INV_X1 port map( I => n16562, ZN => n32568);
   U3690 : NOR2_X1 port map( A1 => n32483, A2 => n16562, ZN => n2409);
   U3691 : INV_X1 port map( I => n16646, ZN => n19834);
   U3698 : NAND2_X1 port map( A1 => n19151, A2 => n11072, ZN => n2152);
   U3702 : NOR2_X1 port map( A1 => n6976, A2 => n5379, ZN => n30718);
   U3706 : NAND2_X1 port map( A1 => n6976, A2 => n5379, ZN => n2381);
   U3712 : NOR3_X1 port map( A1 => n2744, A2 => n24317, A3 => n26938, ZN => 
                           n33512);
   U3719 : NAND2_X1 port map( A1 => n26938, A2 => n13232, ZN => n14663);
   U3724 : NAND2_X1 port map( A1 => n26938, A2 => n32298, ZN => n2993);
   U3737 : AOI22_X1 port map( A1 => n24318, A2 => n26938, B1 => n2744, B2 => 
                           n24317, ZN => n24319);
   U3740 : NAND2_X1 port map( A1 => n6457, A2 => n11941, ZN => n3113);
   U3745 : INV_X2 port map( I => n11941, ZN => n16318);
   U3748 : NOR2_X1 port map( A1 => n33834, A2 => n14419, ZN => n29817);
   U3749 : INV_X1 port map( I => n7345, ZN => n945);
   U3751 : NAND2_X1 port map( A1 => n21627, A2 => n14095, ZN => n14153);
   U3752 : NOR2_X1 port map( A1 => n29322, A2 => n14095, ZN => n33459);
   U3756 : NOR2_X1 port map( A1 => n13773, A2 => n16333, ZN => n9714);
   U3757 : OAI21_X1 port map( A1 => n23881, A2 => n13773, B => n23882, ZN => 
                           n7170);
   U3758 : AOI22_X1 port map( A1 => n9714, A2 => n23787, B1 => n10619, B2 => 
                           n13773, ZN => n32942);
   U3760 : INV_X2 port map( I => n13773, ZN => n16320);
   U3763 : NAND2_X1 port map( A1 => n5915, A2 => n5696, ZN => n28970);
   U3765 : INV_X2 port map( I => n14365, ZN => n1355);
   U3766 : NOR2_X1 port map( A1 => n14365, A2 => n31907, ZN => n20435);
   U3767 : INV_X1 port map( I => n8625, ZN => n13286);
   U3770 : INV_X1 port map( I => n20518, ZN => n932);
   U3774 : CLKBUF_X2 port map( I => n20518, Z => n6530);
   U3776 : BUF_X2 port map( I => n21198, Z => n13896);
   U3777 : NOR2_X1 port map( A1 => n31161, A2 => n8100, ZN => n12297);
   U3784 : NOR2_X1 port map( A1 => n4359, A2 => n4356, ZN => n33746);
   U3785 : OAI21_X1 port map( A1 => n21855, A2 => n12229, B => n4356, ZN => 
                           n33664);
   U3786 : NAND2_X1 port map( A1 => n32642, A2 => n4356, ZN => n21823);
   U3788 : OAI21_X1 port map( A1 => n21853, A2 => n4356, B => n5546, ZN => 
                           n17748);
   U3791 : NAND2_X1 port map( A1 => n4184, A2 => n13558, ZN => n23107);
   U3793 : INV_X1 port map( I => n13558, ZN => n2713);
   U3796 : NAND2_X1 port map( A1 => n14131, A2 => n13558, ZN => n13386);
   U3798 : CLKBUF_X2 port map( I => n22127, Z => n28709);
   U3808 : INV_X1 port map( I => n22127, ZN => n26193);
   U3816 : NAND2_X1 port map( A1 => n16743, A2 => n16938, ZN => n33423);
   U3818 : NAND2_X1 port map( A1 => n10665, A2 => n18071, ZN => n18254);
   U3824 : OAI21_X1 port map( A1 => n17316, A2 => n34139, B => n33687, ZN => 
                           n12151);
   U3825 : AND2_X1 port map( A1 => n23862, A2 => n26290, Z => n9261);
   U3829 : NAND2_X1 port map( A1 => n23862, A2 => n23864, ZN => n33724);
   U3831 : INV_X1 port map( I => n15715, ZN => n20377);
   U3835 : NOR2_X1 port map( A1 => n14179, A2 => n15715, ZN => n9719);
   U3836 : OAI21_X1 port map( A1 => n1291, A2 => n26708, B => n15853, ZN => 
                           n7427);
   U3842 : OAI21_X1 port map( A1 => n26173, A2 => n26708, B => n29336, ZN => 
                           n33105);
   U3845 : NOR2_X1 port map( A1 => n26708, A2 => n26709, ZN => n34002);
   U3846 : NAND2_X1 port map( A1 => n22608, A2 => n26708, ZN => n32450);
   U3850 : INV_X2 port map( I => n32605, ZN => n26708);
   U3856 : BUF_X2 port map( I => n9292, Z => n4975);
   U3860 : INV_X1 port map( I => n14821, ZN => n20236);
   U3861 : BUF_X2 port map( I => n14821, Z => n7486);
   U3862 : INV_X1 port map( I => n19679, ZN => n17129);
   U3868 : NAND2_X1 port map( A1 => n5318, A2 => n29634, ZN => n16985);
   U3870 : CLKBUF_X2 port map( I => n5318, Z => n28833);
   U3871 : CLKBUF_X4 port map( I => n20521, Z => n16218);
   U3873 : NAND3_X1 port map( A1 => n15096, A2 => n737, A3 => n27038, ZN => 
                           n1837);
   U3878 : NAND2_X1 port map( A1 => n33019, A2 => n15096, ZN => n1496);
   U3879 : NAND3_X1 port map( A1 => n15096, A2 => n13334, A3 => n27184, ZN => 
                           n5129);
   U3882 : NAND2_X1 port map( A1 => n25757, A2 => n26056, ZN => n30259);
   U3888 : INV_X1 port map( I => n14682, ZN => n2649);
   U3896 : INV_X1 port map( I => n9287, ZN => n20628);
   U3903 : CLKBUF_X4 port map( I => n9287, Z => n9014);
   U3906 : INV_X1 port map( I => n2859, ZN => n31835);
   U3907 : BUF_X2 port map( I => n2859, Z => n2738);
   U3908 : NAND3_X1 port map( A1 => n5452, A2 => n4547, A3 => n16567, ZN => 
                           n31418);
   U3910 : OAI22_X1 port map( A1 => n5452, A2 => n6658, B1 => n22578, B2 => 
                           n29021, ZN => n5449);
   U3912 : AOI21_X1 port map( A1 => n5452, A2 => n22666, B => n22576, ZN => 
                           n5451);
   U3916 : CLKBUF_X4 port map( I => n22156, Z => n22664);
   U3920 : INV_X1 port map( I => n23899, ZN => n28914);
   U3924 : NAND2_X1 port map( A1 => n6985, A2 => n1577, ZN => n30945);
   U3925 : NOR2_X1 port map( A1 => n12593, A2 => n7778, ZN => n24293);
   U3926 : CLKBUF_X2 port map( I => n12593, Z => n26544);
   U3927 : NAND2_X1 port map( A1 => n12593, A2 => n7778, ZN => n32444);
   U3929 : INV_X1 port map( I => n4897, ZN => n15065);
   U3930 : NAND2_X1 port map( A1 => n15720, A2 => n4897, ZN => n15996);
   U3932 : NAND2_X1 port map( A1 => n23738, A2 => n23737, ZN => n23739);
   U3936 : INV_X1 port map( I => n21442, ZN => n6277);
   U3938 : INV_X1 port map( I => n23429, ZN => n29970);
   U3943 : NOR2_X1 port map( A1 => n27726, A2 => n745, ZN => n19287);
   U3945 : NAND2_X1 port map( A1 => n19288, A2 => n745, ZN => n9356);
   U3951 : INV_X1 port map( I => n19275, ZN => n19320);
   U3954 : NAND2_X1 port map( A1 => n19275, A2 => n19318, ZN => n33108);
   U3955 : NAND2_X1 port map( A1 => n27132, A2 => n19275, ZN => n18419);
   U3957 : NAND3_X1 port map( A1 => n808, A2 => n896, A3 => n22399, ZN => 
                           n15578);
   U3958 : NAND2_X1 port map( A1 => n32856, A2 => n25615, ZN => n28791);
   U3961 : NOR2_X1 port map( A1 => n5817, A2 => n30687, ZN => n30990);
   U3963 : NAND2_X1 port map( A1 => n2826, A2 => n24164, ZN => n17280);
   U3966 : NOR2_X1 port map( A1 => n14840, A2 => n2826, ZN => n14839);
   U3972 : NAND2_X1 port map( A1 => n4846, A2 => n4847, ZN => n32480);
   U3974 : NAND2_X1 port map( A1 => n12044, A2 => n27143, ZN => n21297);
   U3977 : CLKBUF_X4 port map( I => n12044, Z => n4324);
   U3979 : AND3_X1 port map( A1 => n21115, A2 => n12044, A3 => n21405, Z => 
                           n15466);
   U3986 : NOR2_X1 port map( A1 => n24221, A2 => n5306, ZN => n33935);
   U3987 : NOR3_X1 port map( A1 => n27077, A2 => n30010, A3 => n5789, ZN => 
                           n26164);
   U3991 : AND2_X1 port map( A1 => n29763, A2 => n8374, Z => n29453);
   U3994 : NOR2_X1 port map( A1 => n8374, A2 => n29763, ZN => n12541);
   U3995 : CLKBUF_X2 port map( I => n26724, Z => n30573);
   U3998 : INV_X2 port map( I => n22816, ZN => n23093);
   U3999 : NAND2_X1 port map( A1 => n22816, A2 => n27419, ZN => n12511);
   U4000 : NAND2_X1 port map( A1 => n14686, A2 => n22816, ZN => n22697);
   U4002 : INV_X1 port map( I => n14402, ZN => n32500);
   U4003 : BUF_X2 port map( I => n14402, Z => n29107);
   U4007 : INV_X2 port map( I => n22585, ZN => n1290);
   U4008 : NAND2_X1 port map( A1 => n6478, A2 => n22585, ZN => n7239);
   U4009 : BUF_X2 port map( I => n22585, Z => n32483);
   U4010 : CLKBUF_X2 port map( I => n7093, Z => n33990);
   U4011 : CLKBUF_X1 port map( I => n13586, Z => n33927);
   U4013 : NOR2_X1 port map( A1 => n17872, A2 => n14756, ZN => n7406);
   U4017 : INV_X2 port map( I => n20945, ZN => n810);
   U4018 : NOR2_X1 port map( A1 => n29240, A2 => n23713, ZN => n32210);
   U4026 : NOR2_X1 port map( A1 => n17234, A2 => n23713, ZN => n31696);
   U4027 : NAND2_X1 port map( A1 => n16615, A2 => n23735, ZN => n23738);
   U4028 : OAI21_X1 port map( A1 => n1489, A2 => n16121, B => n16615, ZN => 
                           n32931);
   U4031 : NOR2_X1 port map( A1 => n16615, A2 => n23735, ZN => n23351);
   U4040 : INV_X1 port map( I => n25119, ZN => n24884);
   U4042 : OR3_X1 port map( A1 => n25119, A2 => n18154, A3 => n27651, Z => 
                           n25021);
   U4047 : NOR2_X1 port map( A1 => n17879, A2 => n7965, ZN => n13143);
   U4054 : NAND2_X1 port map( A1 => n33032, A2 => n22791, ZN => n15390);
   U4057 : NAND2_X1 port map( A1 => n14770, A2 => n7188, ZN => n2070);
   U4061 : AOI21_X1 port map( A1 => n23621, A2 => n13176, B => n15977, ZN => 
                           n23622);
   U4062 : NOR2_X1 port map( A1 => n13330, A2 => n947, ZN => n14649);
   U4067 : NAND3_X1 port map( A1 => n16485, A2 => n13330, A3 => n13328, ZN => 
                           n13791);
   U4068 : INV_X1 port map( I => n13330, ZN => n17508);
   U4069 : NOR2_X1 port map( A1 => n13100, A2 => n17039, ZN => n9967);
   U4075 : CLKBUF_X2 port map( I => n33986, Z => n33822);
   U4081 : NOR2_X1 port map( A1 => n1056, A2 => n33986, ZN => n32218);
   U4082 : BUF_X2 port map( I => n1808, Z => n1634);
   U4084 : CLKBUF_X2 port map( I => n1808, Z => n32515);
   U4086 : OAI21_X1 port map( A1 => n1808, A2 => n32102, B => n16535, ZN => 
                           n2427);
   U4087 : CLKBUF_X2 port map( I => n5863, Z => n27596);
   U4088 : NOR2_X1 port map( A1 => n26169, A2 => n30231, ZN => n32233);
   U4091 : AND2_X1 port map( A1 => n7463, A2 => n30231, Z => n5821);
   U4092 : NOR2_X1 port map( A1 => n30643, A2 => n27105, ZN => n16176);
   U4095 : NAND2_X1 port map( A1 => n24275, A2 => n2654, ZN => n7067);
   U4096 : CLKBUF_X12 port map( I => n15077, Z => n8576);
   U4103 : XOR2_X1 port map( A1 => n10576, A2 => n17650, Z => n31922);
   U4108 : OR2_X2 port map( A1 => n12744, A2 => n17556, Z => n31923);
   U4110 : INV_X2 port map( I => n33665, ZN => n32930);
   U4114 : OR2_X1 port map( A1 => n502, A2 => n5433, Z => n31924);
   U4116 : INV_X2 port map( I => n20423, ZN => n20566);
   U4117 : OAI21_X1 port map( A1 => n28786, A2 => n1170, B => n33241, ZN => 
                           n32903);
   U4118 : OAI22_X2 port map( A1 => n31444, A2 => n15714, B1 => n20224, B2 => 
                           n1030, ZN => n1923);
   U4125 : AND2_X1 port map( A1 => n21239, A2 => n5822, Z => n31925);
   U4127 : AND2_X1 port map( A1 => n30769, A2 => n26337, Z => n31926);
   U4130 : OR2_X1 port map( A1 => n8875, A2 => n30033, Z => n31927);
   U4131 : INV_X1 port map( I => n21693, ZN => n11301);
   U4133 : INV_X1 port map( I => n27635, ZN => n33242);
   U4138 : INV_X2 port map( I => n7289, ZN => n34050);
   U4143 : XNOR2_X1 port map( A1 => n9536, A2 => n30018, ZN => n31928);
   U4145 : XNOR2_X1 port map( A1 => n14416, A2 => n15969, ZN => n31929);
   U4148 : INV_X1 port map( I => n26317, ZN => n11250);
   U4150 : INV_X4 port map( I => n28203, ZN => n8029);
   U4151 : XNOR2_X1 port map( A1 => n6543, A2 => n7152, ZN => n31931);
   U4153 : XOR2_X1 port map( A1 => n2309, A2 => n31303, Z => n31932);
   U4155 : INV_X1 port map( I => n9535, ZN => n22642);
   U4157 : CLKBUF_X4 port map( I => n9535, Z => n33594);
   U4159 : OR2_X2 port map( A1 => n22622, A2 => n22340, Z => n31933);
   U4162 : NOR2_X2 port map( A1 => n4396, A2 => n29288, ZN => n33283);
   U4164 : BUF_X4 port map( I => n23005, Z => n31942);
   U4167 : AND2_X1 port map( A1 => n27752, A2 => n30293, Z => n31935);
   U4177 : NAND2_X2 port map( A1 => n33126, A2 => n11382, ZN => n23391);
   U4180 : AND2_X1 port map( A1 => n10031, A2 => n15301, Z => n31936);
   U4183 : OR2_X2 port map( A1 => n13894, A2 => n4700, Z => n31937);
   U4184 : INV_X1 port map( I => n15722, ZN => n23935);
   U4191 : INV_X1 port map( I => n10463, ZN => n23918);
   U4192 : CLKBUF_X4 port map( I => n10463, Z => n8760);
   U4198 : BUF_X4 port map( I => n23586, Z => n16496);
   U4199 : AND2_X2 port map( A1 => n31915, A2 => n26641, Z => n31938);
   U4203 : INV_X2 port map( I => n24095, ZN => n24097);
   U4205 : INV_X2 port map( I => n24171, ZN => n24271);
   U4208 : INV_X4 port map( I => n29305, ZN => n32308);
   U4209 : XOR2_X1 port map( A1 => n27360, A2 => n24470, Z => n31939);
   U4212 : INV_X2 port map( I => n25412, ZN => n25406);
   U4223 : CLKBUF_X4 port map( I => n24511, Z => n25412);
   U4228 : AND2_X1 port map( A1 => n1080, A2 => n17120, Z => n31940);
   U4230 : NOR2_X1 port map( A1 => n16939, A2 => n25238, ZN => n31941);
   U4231 : INV_X2 port map( I => n25044, ZN => n27610);
   U4246 : NAND2_X1 port map( A1 => n22744, A2 => n1266, ZN => n9085);
   U4248 : OAI22_X1 port map( A1 => n22744, A2 => n7310, B1 => n11018, B2 => 
                           n1266, ZN => n30633);
   U4250 : NAND2_X1 port map( A1 => n18681, A2 => n5700, ZN => n19295);
   U4251 : OAI21_X1 port map( A1 => n18681, A2 => n18683, B => n29726, ZN => 
                           n7320);
   U4252 : NAND2_X1 port map( A1 => n25981, A2 => n18681, ZN => n29726);
   U4256 : INV_X2 port map( I => n18681, ZN => n15873);
   U4257 : OR2_X2 port map( A1 => n14534, A2 => n32628, Z => n6192);
   U4260 : AND2_X2 port map( A1 => n20468, A2 => n28471, Z => n17964);
   U4264 : BUF_X2 port map( I => n20468, Z => n28626);
   U4269 : NOR2_X1 port map( A1 => n12263, A2 => n17328, ZN => n19930);
   U4271 : NOR2_X1 port map( A1 => n13253, A2 => n17328, ZN => n31398);
   U4324 : INV_X1 port map( I => n17328, ZN => n3562);
   U4327 : NOR2_X1 port map( A1 => n20566, A2 => n17328, ZN => n28043);
   U4328 : AND2_X2 port map( A1 => n6531, A2 => n17328, Z => n15553);
   U4330 : AOI21_X1 port map( A1 => n9285, A2 => n12827, B => n31042, ZN => 
                           n8651);
   U4332 : NOR2_X1 port map( A1 => n9285, A2 => n12827, ZN => n31484);
   U4334 : NAND2_X1 port map( A1 => n21553, A2 => n12827, ZN => n21235);
   U4336 : NAND2_X1 port map( A1 => n9285, A2 => n12827, ZN => n31041);
   U4337 : CLKBUF_X4 port map( I => n7463, Z => n5820);
   U4343 : NOR2_X2 port map( A1 => n13474, A2 => n6553, ZN => n13142);
   U4351 : NAND2_X1 port map( A1 => n32619, A2 => n2612, ZN => n33795);
   U4354 : NAND2_X1 port map( A1 => n30033, A2 => n29523, ZN => n13115);
   U4355 : AOI21_X1 port map( A1 => n21859, A2 => n30033, B => n21858, ZN => 
                           n2351);
   U4358 : INV_X2 port map( I => n10953, ZN => n9646);
   U4360 : OR2_X2 port map( A1 => n31787, A2 => n17150, Z => n16091);
   U4364 : CLKBUF_X12 port map( I => n23005, Z => n31943);
   U4368 : AND2_X2 port map( A1 => n28014, A2 => n9753, Z => n22674);
   U4375 : OR3_X2 port map( A1 => n9737, A2 => n32078, A3 => n9910, Z => n22421
                           );
   U4387 : CLKBUF_X4 port map( I => n19456, Z => n5825);
   U4394 : INV_X2 port map( I => n19456, ZN => n19992);
   U4395 : AND2_X2 port map( A1 => n17930, A2 => n12375, Z => n9184);
   U4396 : OAI21_X1 port map( A1 => n25306, A2 => n18059, B => n1215, ZN => 
                           n27443);
   U4401 : INV_X1 port map( I => n23454, ZN => n23455);
   U4402 : AND3_X2 port map( A1 => n21350, A2 => n32505, A3 => n14983, Z => 
                           n3317);
   U4405 : NAND2_X1 port map( A1 => n21350, A2 => n30389, ZN => n16228);
   U4406 : NOR2_X1 port map( A1 => n8140, A2 => n28181, ZN => n2801);
   U4410 : INV_X2 port map( I => n5994, ZN => n22114);
   U4412 : NOR2_X2 port map( A1 => n30908, A2 => n10305, ZN => n10307);
   U4414 : NAND2_X1 port map( A1 => n31461, A2 => n24168, ZN => n34136);
   U4417 : AND2_X2 port map( A1 => n20561, A2 => n20413, Z => n5953);
   U4419 : NOR2_X1 port map( A1 => n33069, A2 => n784, ZN => n18916);
   U4421 : NOR2_X1 port map( A1 => n20119, A2 => n14815, ZN => n20122);
   U4425 : INV_X2 port map( I => n14815, ZN => n20021);
   U4426 : CLKBUF_X12 port map( I => n14815, Z => n8371);
   U4428 : AND2_X2 port map( A1 => n20561, A2 => n1636, Z => n5950);
   U4435 : INV_X2 port map( I => n20561, ZN => n30931);
   U4436 : INV_X1 port map( I => n30293, ZN => n22828);
   U4437 : OR2_X2 port map( A1 => n16603, A2 => n23144, Z => n23712);
   U4439 : CLKBUF_X12 port map( I => n652, Z => n27);
   U4440 : OR2_X2 port map( A1 => n7463, A2 => n12055, Z => n3901);
   U4441 : CLKBUF_X12 port map( I => n26317, Z => n28692);
   U4443 : OAI21_X1 port map( A1 => n9186, A2 => n424, B => n780, ZN => n9395);
   U4444 : NAND3_X1 port map( A1 => n29088, A2 => n6493, A3 => n424, ZN => 
                           n5687);
   U4447 : INV_X2 port map( I => n424, ZN => n6908);
   U4449 : INV_X1 port map( I => n23230, ZN => n12922);
   U4454 : NOR2_X1 port map( A1 => n24060, A2 => n30191, ZN => n26580);
   U4456 : NAND2_X1 port map( A1 => n3147, A2 => n30191, ZN => n14725);
   U4457 : AOI22_X1 port map( A1 => n20524, A2 => n2958, B1 => n868, B2 => 
                           n31504, ZN => n4398);
   U4458 : NAND2_X1 port map( A1 => n2879, A2 => n2958, ZN => n12771);
   U4459 : INV_X1 port map( I => n2958, ZN => n33225);
   U4460 : OR2_X2 port map( A1 => n28979, A2 => n26330, Z => n26709);
   U4461 : INV_X1 port map( I => n13762, ZN => n805);
   U4464 : AOI22_X1 port map( A1 => n22950, A2 => n22949, B1 => n22951, B2 => 
                           n13762, ZN => n17202);
   U4467 : CLKBUF_X12 port map( I => n13195, Z => n27028);
   U4469 : INV_X1 port map( I => n3395, ZN => n2763);
   U4476 : NAND2_X1 port map( A1 => n2913, A2 => n24315, ZN => n12005);
   U4477 : CLKBUF_X12 port map( I => n24315, Z => n31377);
   U4480 : NOR2_X1 port map( A1 => n31072, A2 => n33117, ZN => n20308);
   U4482 : NOR2_X1 port map( A1 => n742, A2 => n33117, ZN => n3226);
   U4489 : AND2_X2 port map( A1 => n33117, A2 => n26363, Z => n29432);
   U4490 : INV_X1 port map( I => n24254, ZN => n29120);
   U4494 : INV_X1 port map( I => n24747, ZN => n33058);
   U4495 : CLKBUF_X12 port map( I => n22873, Z => n18240);
   U4496 : NOR2_X1 port map( A1 => n4135, A2 => n9377, ZN => n33861);
   U4500 : BUF_X2 port map( I => n18575, Z => n15108);
   U4501 : INV_X2 port map( I => n21579, ZN => n21805);
   U4503 : OAI21_X1 port map( A1 => n32634, A2 => n19093, B => n8141, ZN => 
                           n8013);
   U4507 : OR3_X2 port map( A1 => n29047, A2 => n8141, A3 => n5813, Z => n27930
                           );
   U4509 : NAND2_X1 port map( A1 => n8141, A2 => n19095, ZN => n19097);
   U4510 : OAI22_X1 port map( A1 => n19977, A2 => n14761, B1 => n1699, B2 => 
                           n32745, ZN => n29548);
   U4511 : NAND2_X1 port map( A1 => n28011, A2 => n20519, ZN => n20288);
   U4512 : INV_X2 port map( I => n28011, ZN => n16174);
   U4519 : OAI21_X1 port map( A1 => n21466, A2 => n1134, B => n6678, ZN => 
                           n16889);
   U4521 : INV_X1 port map( I => n21466, ZN => n16577);
   U4524 : NAND2_X1 port map( A1 => n19165, A2 => n4835, ZN => n19153);
   U4530 : CLKBUF_X4 port map( I => n8396, Z => n7090);
   U4533 : INV_X1 port map( I => n8396, ZN => n22460);
   U4534 : NAND2_X1 port map( A1 => n17516, A2 => n1439, ZN => n18316);
   U4537 : INV_X2 port map( I => n17516, ZN => n18710);
   U4541 : BUF_X2 port map( I => n17516, Z => n33783);
   U4544 : INV_X2 port map( I => n29634, ZN => n24152);
   U4553 : AND2_X2 port map( A1 => n31787, A2 => n23833, Z => n29375);
   U4558 : OR2_X2 port map( A1 => n23925, A2 => n14585, Z => n11192);
   U4559 : BUF_X2 port map( I => n25589, Z => n31945);
   U4560 : CLKBUF_X12 port map( I => n25703, Z => n16323);
   U4561 : OR2_X2 port map( A1 => n15057, A2 => n10708, Z => n13650);
   U4564 : OAI21_X1 port map( A1 => n6003, A2 => n24095, B => n24015, ZN => 
                           n4393);
   U4566 : AND3_X2 port map( A1 => n14443, A2 => n6001, A3 => n24095, Z => 
                           n29396);
   U4567 : NOR2_X1 port map( A1 => n24095, A2 => n33868, ZN => n12312);
   U4571 : AOI21_X1 port map( A1 => n12452, A2 => n21463, B => n26439, ZN => 
                           n26325);
   U4574 : OAI21_X1 port map( A1 => n33810, A2 => n21604, B => n26439, ZN => 
                           n27454);
   U4588 : INV_X2 port map( I => n30894, ZN => n1177);
   U4592 : NAND2_X1 port map( A1 => n30894, A2 => n19274, ZN => n19323);
   U4593 : INV_X2 port map( I => n27419, ZN => n776);
   U4596 : OR2_X2 port map( A1 => n20148, A2 => n7865, Z => n29422);
   U4598 : INV_X1 port map( I => n17098, ZN => n16345);
   U4602 : NAND3_X1 port map( A1 => n24325, A2 => n24328, A3 => n10987, ZN => 
                           n26990);
   U4617 : NOR2_X1 port map( A1 => n2302, A2 => n30219, ZN => n2301);
   U4618 : NAND2_X1 port map( A1 => n28429, A2 => n14691, ZN => n21649);
   U4620 : NOR2_X1 port map( A1 => n14691, A2 => n28429, ZN => n2061);
   U4621 : CLKBUF_X12 port map( I => n28429, Z => n33139);
   U4622 : CLKBUF_X12 port map( I => n17779, Z => n17118);
   U4626 : INV_X1 port map( I => n17779, ZN => n24974);
   U4628 : AND2_X2 port map( A1 => n23746, A2 => n23603, Z => n15659);
   U4630 : NOR2_X1 port map( A1 => n11850, A2 => n31915, ZN => n29590);
   U4637 : NOR2_X1 port map( A1 => n6394, A2 => n11850, ZN => n32574);
   U4638 : NAND2_X1 port map( A1 => n4774, A2 => n12981, ZN => n24027);
   U4642 : INV_X1 port map( I => n12981, ZN => n12574);
   U4660 : CLKBUF_X12 port map( I => n12981, Z => n4118);
   U4661 : OR2_X2 port map( A1 => n23087, A2 => n23086, Z => n26242);
   U4663 : NAND3_X2 port map( A1 => n9915, A2 => n9916, A3 => n25390, ZN => 
                           n33064);
   U4666 : CLKBUF_X4 port map( I => n23197, Z => n23806);
   U4671 : CLKBUF_X12 port map( I => n30865, Z => n31947);
   U4672 : CLKBUF_X12 port map( I => n30865, Z => n31949);
   U4674 : INV_X1 port map( I => n13723, ZN => n20945);
   U4678 : BUF_X4 port map( I => n25988, Z => n31950);
   U4679 : INV_X1 port map( I => n11710, ZN => n20332);
   U4684 : OAI21_X1 port map( A1 => n6475, A2 => n31390, B => n11710, ZN => 
                           n8702);
   U4686 : NAND2_X1 port map( A1 => n7873, A2 => n20613, ZN => n28437);
   U4690 : NOR2_X1 port map( A1 => n14129, A2 => n22968, ZN => n22884);
   U4692 : INV_X1 port map( I => n14129, ZN => n17084);
   U4693 : AND2_X2 port map( A1 => n14129, A2 => n7802, Z => n27639);
   U4698 : INV_X2 port map( I => n12323, ZN => n28406);
   U4712 : AOI21_X1 port map( A1 => n3717, A2 => n12323, B => n30313, ZN => 
                           n21176);
   U4714 : NAND2_X1 port map( A1 => n12323, A2 => n595, ZN => n21055);
   U4717 : AOI21_X1 port map( A1 => n13386, A2 => n2638, B => n4184, ZN => 
                           n13384);
   U4719 : INV_X1 port map( I => n23741, ZN => n23769);
   U4721 : NOR2_X1 port map( A1 => n23741, A2 => n386, ZN => n8093);
   U4722 : AOI21_X1 port map( A1 => n23741, A2 => n17396, B => n30895, ZN => 
                           n33542);
   U4727 : AOI21_X1 port map( A1 => n23741, A2 => n23597, B => n23598, ZN => 
                           n14551);
   U4729 : NAND2_X1 port map( A1 => n23741, A2 => n30089, ZN => n2878);
   U4737 : NAND2_X1 port map( A1 => n27183, A2 => n25317, ZN => n1803);
   U4753 : INV_X1 port map( I => n25317, ZN => n31178);
   U4757 : AOI21_X1 port map( A1 => n977, A2 => n13773, B => n11943, ZN => 
                           n4514);
   U4759 : OAI22_X1 port map( A1 => n16320, A2 => n11943, B1 => n23882, B2 => 
                           n8544, ZN => n33535);
   U4765 : NAND2_X1 port map( A1 => n9714, A2 => n11943, ZN => n7167);
   U4770 : AOI21_X1 port map( A1 => n16320, A2 => n11943, B => n8544, ZN => 
                           n10620);
   U4773 : NAND2_X1 port map( A1 => n15261, A2 => n21438, ZN => n21440);
   U4775 : INV_X2 port map( I => n21438, ZN => n15589);
   U4780 : OR2_X2 port map( A1 => n29101, A2 => n15229, Z => n17936);
   U4785 : AOI22_X1 port map( A1 => n19030, A2 => n29223, B1 => n19300, B2 => 
                           n19029, ZN => n31066);
   U4786 : AOI22_X1 port map( A1 => n19085, A2 => n29223, B1 => n19084, B2 => 
                           n19300, ZN => n28237);
   U4794 : AND3_X2 port map( A1 => n20946, A2 => n10599, A3 => n10787, Z => 
                           n34159);
   U4797 : OR2_X2 port map( A1 => n20946, A2 => n13195, Z => n21313);
   U4801 : NAND2_X1 port map( A1 => n11086, A2 => n2821, ZN => n20261);
   U4809 : NAND2_X1 port map( A1 => n919, A2 => n28580, ZN => n26527);
   U4813 : NOR2_X1 port map( A1 => n28580, A2 => n12535, ZN => n32148);
   U4814 : NAND2_X1 port map( A1 => n28580, A2 => n10720, ZN => n32435);
   U4824 : INV_X1 port map( I => n28580, ZN => n21645);
   U4825 : INV_X1 port map( I => n12424, ZN => n21777);
   U4826 : CLKBUF_X12 port map( I => n12424, Z => n30940);
   U4828 : CLKBUF_X4 port map( I => n12424, Z => n11861);
   U4837 : CLKBUF_X12 port map( I => n24372, Z => n17833);
   U4838 : CLKBUF_X4 port map( I => n19829, Z => n31951);
   U4840 : NAND2_X1 port map( A1 => n23087, A2 => n4834, ZN => n28427);
   U4841 : CLKBUF_X12 port map( I => n12804, Z => n179);
   U4851 : INV_X1 port map( I => n20455, ZN => n20457);
   U4860 : NAND2_X1 port map( A1 => n20455, A2 => n15468, ZN => n14767);
   U4864 : INV_X1 port map( I => n17517, ZN => n33814);
   U4866 : NOR2_X1 port map( A1 => n23110, A2 => n3103, ZN => n22813);
   U4870 : NAND2_X1 port map( A1 => n853, A2 => n3103, ZN => n4935);
   U4872 : NAND2_X1 port map( A1 => n16022, A2 => n3103, ZN => n23108);
   U4874 : INV_X2 port map( I => n3103, ZN => n6012);
   U4875 : OAI21_X1 port map( A1 => n30168, A2 => n30167, B => n22999, ZN => 
                           n4305);
   U4876 : INV_X1 port map( I => n22999, ZN => n7220);
   U4877 : OR2_X2 port map( A1 => n9280, A2 => n22999, Z => n9213);
   U4880 : OAI21_X2 port map( A1 => n23101, A2 => n11956, B => n22999, ZN => 
                           n15935);
   U4882 : NAND2_X1 port map( A1 => n29883, A2 => n7935, ZN => n32328);
   U4884 : OR2_X2 port map( A1 => n18039, A2 => n26699, Z => n8182);
   U4885 : NAND2_X1 port map( A1 => n31129, A2 => n23051, ZN => n6102);
   U4887 : INV_X2 port map( I => n31129, ZN => n1108);
   U4888 : NAND2_X1 port map( A1 => n772, A2 => n31129, ZN => n1746);
   U4889 : AND2_X2 port map( A1 => n5962, A2 => n11986, Z => n8846);
   U4890 : INV_X2 port map( I => n32253, ZN => n14625);
   U4892 : NOR2_X1 port map( A1 => n7279, A2 => n20627, ZN => n8242);
   U4895 : OR2_X2 port map( A1 => n20627, A2 => n7280, Z => n17002);
   U4896 : BUF_X2 port map( I => n16954, Z => n8886);
   U4899 : NAND2_X1 port map( A1 => n16954, A2 => n15302, ZN => n27338);
   U4900 : NOR2_X1 port map( A1 => n28581, A2 => n16954, ZN => n31231);
   U4903 : NOR2_X1 port map( A1 => n14893, A2 => n5625, ZN => n12996);
   U4906 : NAND2_X1 port map( A1 => n19057, A2 => n5625, ZN => n18944);
   U4910 : CLKBUF_X4 port map( I => n5086, Z => n31954);
   U4913 : INV_X1 port map( I => n21891, ZN => n2082);
   U4922 : OR2_X2 port map( A1 => n31497, A2 => n24216, Z => n215);
   U4929 : INV_X1 port map( I => n31497, ZN => n24111);
   U4932 : NAND2_X1 port map( A1 => n13175, A2 => n31497, ZN => n13176);
   U4937 : NAND2_X1 port map( A1 => n22791, A2 => n14392, ZN => n31564);
   U4939 : NAND2_X1 port map( A1 => n22871, A2 => n22791, ZN => n22792);
   U4940 : INV_X1 port map( I => n7046, ZN => n4063);
   U4941 : INV_X1 port map( I => n27880, ZN => n621);
   U4944 : INV_X1 port map( I => n33288, ZN => n30425);
   U4946 : OAI21_X1 port map( A1 => n33288, A2 => n20317, B => n20471, ZN => 
                           n19402);
   U4951 : NAND3_X1 port map( A1 => n34113, A2 => n20471, A3 => n33288, ZN => 
                           n20248);
   U4952 : NAND2_X1 port map( A1 => n16144, A2 => n28064, ZN => n13599);
   U4956 : NAND3_X1 port map( A1 => n16144, A2 => n20531, A3 => n20529, ZN => 
                           n32840);
   U4960 : NOR2_X1 port map( A1 => n5274, A2 => n32967, ZN => n33344);
   U4961 : AOI21_X1 port map( A1 => n1112, A2 => n5274, B => n22931, ZN => 
                           n30875);
   U4966 : OAI21_X1 port map( A1 => n17297, A2 => n20324, B => n20515, ZN => 
                           n26576);
   U4968 : NAND2_X1 port map( A1 => n16174, A2 => n20515, ZN => n6491);
   U4970 : CLKBUF_X4 port map( I => n26750, Z => n33544);
   U4972 : NAND2_X1 port map( A1 => n1550, A2 => n24286, ZN => n24047);
   U4978 : CLKBUF_X12 port map( I => n24286, Z => n28300);
   U4985 : INV_X1 port map( I => n24286, ZN => n17277);
   U4993 : INV_X2 port map( I => n1130, ZN => n31706);
   U5002 : NAND2_X1 port map( A1 => n879, A2 => n19330, ZN => n19331);
   U5003 : INV_X1 port map( I => n17891, ZN => n22379);
   U5008 : CLKBUF_X12 port map( I => n17891, Z => n2697);
   U5012 : INV_X2 port map( I => n22361, ZN => n6149);
   U5015 : NOR2_X1 port map( A1 => n22361, A2 => n9575, ZN => n27580);
   U5018 : NOR2_X1 port map( A1 => n4135, A2 => n22361, ZN => n32692);
   U5019 : NOR2_X1 port map( A1 => n5119, A2 => n5118, ZN => n19013);
   U5021 : OAI21_X1 port map( A1 => n5118, A2 => n28929, B => n6511, ZN => 
                           n11489);
   U5024 : INV_X1 port map( I => n11720, ZN => n11911);
   U5025 : NOR2_X1 port map( A1 => n20507, A2 => n31907, ZN => n16167);
   U5026 : NAND2_X1 port map( A1 => n31907, A2 => n16452, ZN => n33501);
   U5027 : AOI21_X1 port map( A1 => n878, A2 => n5760, B => n14498, ZN => 
                           n18497);
   U5032 : NOR2_X1 port map( A1 => n19089, A2 => n14498, ZN => n15021);
   U5038 : INV_X2 port map( I => n14498, ZN => n1385);
   U5039 : NOR2_X1 port map( A1 => n26603, A2 => n32253, ZN => n6142);
   U5040 : NAND2_X1 port map( A1 => n15777, A2 => n9126, ZN => n27272);
   U5043 : OAI21_X1 port map( A1 => n16518, A2 => n28028, B => n32240, ZN => 
                           n20206);
   U5044 : NAND3_X1 port map( A1 => n1153, A2 => n20534, A3 => n28028, ZN => 
                           n18170);
   U5051 : INV_X2 port map( I => n28028, ZN => n8206);
   U5055 : AOI22_X1 port map( A1 => n17896, A2 => n31009, B1 => n28812, B2 => 
                           n4254, ZN => n2609);
   U5058 : NOR2_X1 port map( A1 => n19938, A2 => n16105, ZN => n32109);
   U5066 : NOR2_X2 port map( A1 => n28418, A2 => n28419, ZN => n12599);
   U5071 : AOI21_X1 port map( A1 => n16374, A2 => n16218, B => n15893, ZN => 
                           n13915);
   U5072 : NAND2_X1 port map( A1 => n16374, A2 => n20236, ZN => n14836);
   U5073 : NOR2_X1 port map( A1 => n13768, A2 => n16374, ZN => n15893);
   U5074 : OR2_X2 port map( A1 => n16374, A2 => n20555, Z => n32066);
   U5075 : INV_X1 port map( I => n9434, ZN => n28647);
   U5077 : NAND2_X1 port map( A1 => n9434, A2 => n29133, ZN => n9637);
   U5081 : AND2_X2 port map( A1 => n26848, A2 => n9744, Z => n7723);
   U5085 : OR2_X2 port map( A1 => n9744, A2 => n8899, Z => n21263);
   U5087 : NAND2_X1 port map( A1 => n34139, A2 => n18295, ZN => n12154);
   U5089 : INV_X2 port map( I => n17817, ZN => n19196);
   U5099 : NAND2_X1 port map( A1 => n6290, A2 => n11085, ZN => n19164);
   U5100 : NOR2_X1 port map( A1 => n1165, A2 => n5433, ZN => n11855);
   U5106 : BUF_X2 port map( I => n3007, Z => n28974);
   U5108 : INV_X2 port map( I => n3007, ZN => n17739);
   U5112 : OR2_X2 port map( A1 => n7965, A2 => n2655, Z => n26867);
   U5118 : CLKBUF_X12 port map( I => n7293, Z => n31956);
   U5119 : CLKBUF_X12 port map( I => n7293, Z => n31958);
   U5126 : NAND3_X1 port map( A1 => n14161, A2 => n20628, A3 => n53, ZN => 
                           n13172);
   U5127 : INV_X1 port map( I => n14161, ZN => n20629);
   U5132 : NOR2_X1 port map( A1 => n14005, A2 => n14161, ZN => n30022);
   U5136 : NAND2_X1 port map( A1 => n9616, A2 => n9625, ZN => n8567);
   U5138 : CLKBUF_X4 port map( I => n9616, Z => n891);
   U5141 : AOI21_X1 port map( A1 => n25088, A2 => n25083, B => n25082, ZN => 
                           n30858);
   U5142 : BUF_X1 port map( I => n24960, Z => n28662);
   U5144 : OAI21_X1 port map( A1 => n13273, A2 => n30396, B => n1213, ZN => 
                           n6822);
   U5150 : BUF_X1 port map( I => n3565, Z => n32678);
   U5154 : CLKBUF_X2 port map( I => n25188, Z => n12476);
   U5159 : CLKBUF_X1 port map( I => n24646, Z => n32759);
   U5163 : CLKBUF_X2 port map( I => n13695, Z => n33699);
   U5170 : CLKBUF_X2 port map( I => n24618, Z => n33348);
   U5179 : CLKBUF_X2 port map( I => n27922, Z => n33492);
   U5197 : INV_X1 port map( I => n13458, ZN => n32552);
   U5201 : CLKBUF_X2 port map( I => n24094, Z => n32459);
   U5205 : NOR2_X1 port map( A1 => n24263, A2 => n26950, ZN => n5936);
   U5207 : INV_X2 port map( I => n24210, ZN => n24322);
   U5208 : INV_X2 port map( I => n24008, ZN => n9962);
   U5209 : NAND2_X1 port map( A1 => n14038, A2 => n14039, ZN => n14037);
   U5210 : INV_X1 port map( I => n5627, ZN => n33104);
   U5211 : BUF_X2 port map( I => n23808, Z => n32477);
   U5212 : CLKBUF_X2 port map( I => n8408, Z => n33216);
   U5215 : INV_X1 port map( I => n23742, ZN => n34036);
   U5216 : BUF_X2 port map( I => n23775, Z => n33011);
   U5218 : CLKBUF_X2 port map( I => n29498, Z => n32657);
   U5219 : CLKBUF_X1 port map( I => n10279, Z => n33924);
   U5220 : INV_X2 port map( I => n662, ZN => n31959);
   U5225 : CLKBUF_X2 port map( I => n23389, Z => n32243);
   U5226 : NOR2_X1 port map( A1 => n5983, A2 => n11308, ZN => n26995);
   U5229 : BUF_X2 port map( I => n31937, Z => n33522);
   U5231 : OAI22_X1 port map( A1 => n3997, A2 => n7181, B1 => n22827, B2 => 
                           n11059, ZN => n4476);
   U5237 : AOI21_X1 port map( A1 => n28853, A2 => n28408, B => n2479, ZN => 
                           n32368);
   U5239 : BUF_X1 port map( I => n22880, Z => n33395);
   U5243 : NAND2_X1 port map( A1 => n22855, A2 => n28649, ZN => n32509);
   U5246 : OR2_X1 port map( A1 => n23057, A2 => n23056, Z => n32086);
   U5248 : BUF_X1 port map( I => n11983, Z => n34097);
   U5250 : NOR2_X1 port map( A1 => n6782, A2 => n22945, ZN => n33923);
   U5251 : NAND2_X1 port map( A1 => n31636, A2 => n16627, ZN => n31635);
   U5253 : NAND2_X1 port map( A1 => n33056, A2 => n10796, ZN => n29563);
   U5254 : INV_X1 port map( I => n22404, ZN => n33402);
   U5255 : NAND2_X1 port map( A1 => n16558, A2 => n22412, ZN => n15119);
   U5257 : NOR2_X1 port map( A1 => n22466, A2 => n998, ZN => n28101);
   U5258 : CLKBUF_X2 port map( I => n27122, Z => n32378);
   U5262 : CLKBUF_X2 port map( I => n7072, Z => n33966);
   U5266 : OR2_X1 port map( A1 => n14845, A2 => n16392, Z => n32080);
   U5269 : CLKBUF_X2 port map( I => n22318, Z => n32154);
   U5274 : CLKBUF_X4 port map( I => n7545, Z => n32537);
   U5275 : CLKBUF_X4 port map( I => n14953, Z => n2896);
   U5279 : INV_X1 port map( I => n33459, ZN => n32314);
   U5281 : INV_X1 port map( I => n26206, ZN => n32348);
   U5285 : NAND2_X1 port map( A1 => n3472, A2 => n17077, ZN => n34104);
   U5287 : CLKBUF_X1 port map( I => n914, Z => n33322);
   U5289 : NAND2_X1 port map( A1 => n31007, A2 => n32374, ZN => n32373);
   U5292 : NOR2_X1 port map( A1 => n21842, A2 => n30346, ZN => n33907);
   U5294 : INV_X1 port map( I => n338, ZN => n33908);
   U5296 : CLKBUF_X2 port map( I => n1652, Z => n32282);
   U5302 : CLKBUF_X4 port map( I => n27379, Z => n33810);
   U5305 : CLKBUF_X2 port map( I => n27336, Z => n34098);
   U5306 : CLKBUF_X2 port map( I => n16278, Z => n32642);
   U5313 : CLKBUF_X1 port map( I => n14864, Z => n33833);
   U5314 : BUF_X4 port map( I => n5830, Z => n31960);
   U5318 : AOI21_X1 port map( A1 => n27689, A2 => n21151, B => n27688, ZN => 
                           n26494);
   U5319 : OAI21_X1 port map( A1 => n21286, A2 => n32625, B => n21285, ZN => 
                           n32168);
   U5321 : CLKBUF_X2 port map( I => n21241, Z => n33882);
   U5323 : CLKBUF_X2 port map( I => n16668, Z => n33741);
   U5333 : NAND2_X1 port map( A1 => n21400, A2 => n15874, ZN => n32624);
   U5344 : CLKBUF_X2 port map( I => n4274, Z => n34037);
   U5345 : NOR2_X1 port map( A1 => n16473, A2 => n21152, ZN => n33979);
   U5346 : BUF_X2 port map( I => n599, Z => n33649);
   U5349 : CLKBUF_X2 port map( I => n8028, Z => n16629);
   U5350 : NOR2_X1 port map( A1 => n13573, A2 => n11635, ZN => n30083);
   U5351 : BUF_X1 port map( I => n6431, Z => n27375);
   U5355 : NOR2_X1 port map( A1 => n20277, A2 => n29453, ZN => n32304);
   U5356 : NAND2_X1 port map( A1 => n20231, A2 => n20413, ZN => n285);
   U5359 : OAI21_X1 port map( A1 => n20492, A2 => n14863, B => n33944, ZN => 
                           n30632);
   U5360 : NAND2_X1 port map( A1 => n26881, A2 => n20310, ZN => n9832);
   U5361 : CLKBUF_X2 port map( I => n20472, Z => n32201);
   U5362 : INV_X1 port map( I => n6536, ZN => n33341);
   U5363 : CLKBUF_X2 port map( I => n1351, Z => n32953);
   U5364 : CLKBUF_X2 port map( I => n20534, Z => n32329);
   U5365 : NAND2_X1 port map( A1 => n5781, A2 => n26585, ZN => n17425);
   U5366 : CLKBUF_X4 port map( I => n30637, Z => n33721);
   U5367 : CLKBUF_X2 port map( I => n20485, Z => n31009);
   U5368 : NAND2_X1 port map( A1 => n30017, A2 => n14281, ZN => n33136);
   U5371 : CLKBUF_X2 port map( I => n20138, Z => n32371);
   U5376 : CLKBUF_X2 port map( I => n17670, Z => n32559);
   U5379 : CLKBUF_X2 port map( I => n34119, Z => n33835);
   U5380 : NAND2_X1 port map( A1 => n10192, A2 => n11798, ZN => n33983);
   U5383 : BUF_X4 port map( I => n7492, Z => n10472);
   U5385 : CLKBUF_X2 port map( I => n14194, Z => n32485);
   U5386 : NAND2_X1 port map( A1 => n27941, A2 => n32805, ZN => n33230);
   U5389 : CLKBUF_X2 port map( I => n29781, Z => n32401);
   U5391 : BUF_X1 port map( I => n25971, Z => n34040);
   U5397 : BUF_X2 port map( I => n34107, Z => n32908);
   U5398 : CLKBUF_X1 port map( I => n4016, Z => n32805);
   U5400 : OAI22_X1 port map( A1 => n27641, A2 => n18629, B1 => n18628, B2 => 
                           n18627, ZN => n19149);
   U5406 : NOR2_X1 port map( A1 => n18885, A2 => n10669, ZN => n33255);
   U5407 : INV_X1 port map( I => n4733, ZN => n18622);
   U5408 : NAND2_X1 port map( A1 => n11123, A2 => n17419, ZN => n33421);
   U5409 : INV_X1 port map( I => n29514, ZN => n33101);
   U5410 : BUF_X2 port map( I => n18601, Z => n33472);
   U5414 : NOR2_X1 port map( A1 => n28686, A2 => n18228, ZN => n33309);
   U5416 : CLKBUF_X2 port map( I => n26980, Z => n32337);
   U5421 : NAND3_X1 port map( A1 => n32724, A2 => n28516, A3 => n28517, ZN => 
                           n32730);
   U5424 : AOI21_X1 port map( A1 => n25683, A2 => n25684, B => n25682, ZN => 
                           n16541);
   U5427 : NAND2_X1 port map( A1 => n14101, A2 => n16246, ZN => n32724);
   U5438 : NOR2_X1 port map( A1 => n33464, A2 => n25273, ZN => n14070);
   U5441 : OAI22_X1 port map( A1 => n25456, A2 => n33946, B1 => n25419, B2 => 
                           n25420, ZN => n30746);
   U5449 : AOI22_X1 port map( A1 => n25747, A2 => n25748, B1 => n25749, B2 => 
                           n25750, ZN => n31599);
   U5457 : OAI22_X1 port map( A1 => n10823, A2 => n1951, B1 => n10821, B2 => 
                           n1950, ZN => n32190);
   U5462 : INV_X1 port map( I => n25857, ZN => n406);
   U5473 : OAI22_X1 port map( A1 => n33702, A2 => n788, B1 => n25128, B2 => 
                           n33138, ZN => n6814);
   U5475 : NAND2_X1 port map( A1 => n25412, A2 => n33921, ZN => n9754);
   U5478 : CLKBUF_X2 port map( I => n31236, Z => n33414);
   U5483 : BUF_X2 port map( I => n16509, Z => n15359);
   U5485 : NOR2_X1 port map( A1 => n25583, A2 => n28242, ZN => n28098);
   U5488 : INV_X1 port map( I => n32427, ZN => n7768);
   U5494 : NAND2_X1 port map( A1 => n12386, A2 => n12369, ZN => n32825);
   U5497 : NAND2_X1 port map( A1 => n11994, A2 => n33199, ZN => n26400);
   U5505 : BUF_X1 port map( I => n25403, Z => n32920);
   U5510 : NOR2_X1 port map( A1 => n24730, A2 => n17120, ZN => n32556);
   U5517 : CLKBUF_X2 port map( I => n25865, Z => n33196);
   U5518 : INV_X2 port map( I => n33919, ZN => n31962);
   U5527 : CLKBUF_X2 port map( I => n17861, Z => n32659);
   U5530 : CLKBUF_X4 port map( I => n11372, Z => n33493);
   U5533 : BUF_X2 port map( I => n31783, Z => n33761);
   U5534 : INV_X1 port map( I => n6863, ZN => n32639);
   U5539 : CLKBUF_X2 port map( I => n14665, Z => n33574);
   U5541 : INV_X1 port map( I => n16045, ZN => n33375);
   U5543 : CLKBUF_X2 port map( I => n24760, Z => n33447);
   U5549 : CLKBUF_X2 port map( I => n30323, Z => n32660);
   U5557 : OAI21_X1 port map( A1 => n23701, A2 => n6003, B => n33727, ZN => 
                           n23702);
   U5560 : INV_X1 port map( I => n32677, ZN => n26851);
   U5561 : NAND2_X1 port map( A1 => n1240, A2 => n24219, ZN => n23625);
   U5571 : NAND2_X1 port map( A1 => n29567, A2 => n29566, ZN => n33853);
   U5574 : BUF_X1 port map( I => n14386, Z => n33470);
   U5575 : NAND2_X1 port map( A1 => n11200, A2 => n28945, ZN => n9687);
   U5577 : CLKBUF_X2 port map( I => n24159, Z => n32176);
   U5579 : CLKBUF_X2 port map( I => n15720, Z => n33425);
   U5585 : CLKBUF_X2 port map( I => n4286, Z => n32936);
   U5590 : CLKBUF_X2 port map( I => n33832, Z => n32102);
   U5593 : CLKBUF_X4 port map( I => n11041, Z => n9066);
   U5597 : INV_X1 port map( I => n2558, ZN => n33532);
   U5602 : INV_X2 port map( I => n24106, ZN => n24104);
   U5603 : INV_X2 port map( I => n8412, ZN => n795);
   U5604 : BUF_X4 port map( I => n11789, Z => n10687);
   U5616 : NAND2_X1 port map( A1 => n32336, A2 => n23749, ZN => n27340);
   U5618 : INV_X2 port map( I => n14080, ZN => n23884);
   U5622 : CLKBUF_X4 port map( I => n386, Z => n33867);
   U5624 : CLKBUF_X2 port map( I => n32711, Z => n33097);
   U5626 : NOR2_X1 port map( A1 => n23804, A2 => n14325, ZN => n33595);
   U5628 : CLKBUF_X2 port map( I => n23822, Z => n33110);
   U5630 : INV_X1 port map( I => n33679, ZN => n32973);
   U5635 : OAI21_X1 port map( A1 => n16496, A2 => n15623, B => n8145, ZN => 
                           n12777);
   U5642 : NOR2_X1 port map( A1 => n6247, A2 => n33812, ZN => n17563);
   U5646 : CLKBUF_X2 port map( I => n4892, Z => n33221);
   U5648 : BUF_X1 port map( I => n10213, Z => n26882);
   U5651 : CLKBUF_X2 port map( I => n23603, Z => n33679);
   U5655 : INV_X2 port map( I => n29498, ZN => n23894);
   U5656 : CLKBUF_X2 port map( I => n10673, Z => n33936);
   U5658 : BUF_X2 port map( I => n23931, Z => n10993);
   U5660 : CLKBUF_X2 port map( I => n7699, Z => n33345);
   U5661 : CLKBUF_X2 port map( I => n9796, Z => n33670);
   U5662 : INV_X1 port map( I => n23437, ZN => n32640);
   U5667 : INV_X1 port map( I => n4273, ZN => n32645);
   U5671 : INV_X1 port map( I => n23520, ZN => n32922);
   U5673 : CLKBUF_X2 port map( I => n23292, Z => n34047);
   U5676 : CLKBUF_X2 port map( I => n6373, Z => n28927);
   U5677 : CLKBUF_X2 port map( I => n31727, Z => n32516);
   U5682 : NAND3_X1 port map( A1 => n22804, A2 => n33596, A3 => n22805, ZN => 
                           n29818);
   U5686 : NAND2_X1 port map( A1 => n22756, A2 => n14977, ZN => n33347);
   U5687 : NAND2_X1 port map( A1 => n12742, A2 => n32368, ZN => n28846);
   U5688 : NAND2_X1 port map( A1 => n31795, A2 => n22951, ZN => n3201);
   U5689 : INV_X1 port map( I => n22694, ZN => n33360);
   U5691 : OAI21_X1 port map( A1 => n33923, A2 => n30455, B => n6942, ZN => 
                           n12443);
   U5693 : CLKBUF_X4 port map( I => n28934, Z => n32935);
   U5694 : OR2_X1 port map( A1 => n1577, A2 => n22885, Z => n5259);
   U5697 : NAND2_X1 port map( A1 => n22962, A2 => n29952, ZN => n30946);
   U5698 : CLKBUF_X2 port map( I => n14686, Z => n33968);
   U5707 : CLKBUF_X8 port map( I => n12619, Z => n33675);
   U5721 : BUF_X2 port map( I => n22990, Z => n31798);
   U5722 : BUF_X4 port map( I => n14201, Z => n33132);
   U5730 : INV_X2 port map( I => n22971, ZN => n23106);
   U5731 : AND2_X1 port map( A1 => n22957, A2 => n5035, Z => n32037);
   U5736 : CLKBUF_X4 port map( I => n28697, Z => n30904);
   U5737 : NAND2_X1 port map( A1 => n12097, A2 => n32080, ZN => n32104);
   U5738 : AOI21_X1 port map( A1 => n22571, A2 => n28473, B => n31636, ZN => 
                           n10904);
   U5739 : OAI21_X1 port map( A1 => n4100, A2 => n4459, B => n32344, ZN => 
                           n13983);
   U5744 : NAND2_X1 port map( A1 => n32406, A2 => n22663, ZN => n26404);
   U5755 : INV_X1 port map( I => n22372, ZN => n33180);
   U5756 : INV_X1 port map( I => n5766, ZN => n33456);
   U5762 : NAND2_X1 port map( A1 => n15812, A2 => n14228, ZN => n33948);
   U5765 : NAND2_X1 port map( A1 => n9546, A2 => n9547, ZN => n9545);
   U5769 : NAND2_X1 port map( A1 => n5960, A2 => n5963, ZN => n22607);
   U5770 : INV_X1 port map( I => n7848, ZN => n32344);
   U5775 : NAND2_X1 port map( A1 => n22380, A2 => n22388, ZN => n33753);
   U5778 : NOR2_X1 port map( A1 => n32217, A2 => n32216, ZN => n32215);
   U5780 : CLKBUF_X2 port map( I => n16558, Z => n29597);
   U5783 : CLKBUF_X2 port map( I => n22491, Z => n33750);
   U5785 : INV_X1 port map( I => n22600, ZN => n7633);
   U5786 : AOI22_X1 port map( A1 => n7490, A2 => n22359, B1 => n22551, B2 => 
                           n22391, ZN => n30112);
   U5790 : INV_X2 port map( I => n11917, ZN => n31963);
   U5793 : NAND2_X1 port map( A1 => n16434, A2 => n22429, ZN => n22408);
   U5794 : CLKBUF_X2 port map( I => n11892, Z => n34074);
   U5799 : BUF_X2 port map( I => n622, Z => n10282);
   U5807 : BUF_X2 port map( I => n11083, Z => n10612);
   U5812 : CLKBUF_X2 port map( I => n25963, Z => n34058);
   U5813 : INV_X1 port map( I => n30489, ZN => n32114);
   U5818 : BUF_X2 port map( I => n6569, Z => n32753);
   U5823 : CLKBUF_X4 port map( I => n22216, Z => n34150);
   U5826 : INV_X1 port map( I => n34016, ZN => n26351);
   U5828 : CLKBUF_X1 port map( I => n22145, Z => n33072);
   U5829 : INV_X1 port map( I => n22133, ZN => n32099);
   U5833 : INV_X1 port map( I => n10261, ZN => n3797);
   U5834 : INV_X1 port map( I => n11458, ZN => n33160);
   U5835 : NAND2_X1 port map( A1 => n28665, A2 => n10689, ZN => n33667);
   U5839 : NAND2_X1 port map( A1 => n33459, A2 => n29552, ZN => n607);
   U5843 : NAND2_X1 port map( A1 => n7947, A2 => n7949, ZN => n32149);
   U5848 : NAND2_X1 port map( A1 => n33908, A2 => n33907, ZN => n14738);
   U5850 : INV_X1 port map( I => n21622, ZN => n21623);
   U5855 : NAND2_X1 port map( A1 => n3048, A2 => n4097, ZN => n31871);
   U5861 : INV_X1 port map( I => n26386, ZN => n21683);
   U5864 : AND3_X1 port map( A1 => n21872, A2 => n30832, A3 => n21870, Z => 
                           n30963);
   U5867 : BUF_X2 port map( I => n13884, Z => n32384);
   U5869 : CLKBUF_X2 port map( I => n1313, Z => n31317);
   U5876 : CLKBUF_X4 port map( I => n11401, Z => n7553);
   U5878 : NAND2_X1 port map( A1 => n32223, A2 => n21188, ZN => n10134);
   U5881 : INV_X1 port map( I => n8323, ZN => n21663);
   U5887 : AOI22_X1 port map( A1 => n6826, A2 => n21252, B1 => n9699, B2 => 
                           n11792, ZN => n3924);
   U5888 : NAND2_X1 port map( A1 => n21059, A2 => n17984, ZN => n32521);
   U5893 : BUF_X4 port map( I => n29997, Z => n32252);
   U5900 : NAND2_X1 port map( A1 => n6198, A2 => n32001, ZN => n33826);
   U5902 : NAND2_X1 port map( A1 => n4341, A2 => n2689, ZN => n34130);
   U5905 : CLKBUF_X1 port map( I => n26622, Z => n32441);
   U5906 : OAI21_X1 port map( A1 => n8393, A2 => n33889, B => n33979, ZN => 
                           n12690);
   U5911 : NAND2_X1 port map( A1 => n32624, A2 => n12325, ZN => n16198);
   U5918 : NAND2_X1 port map( A1 => n31180, A2 => n17731, ZN => n32815);
   U5921 : AND2_X1 port map( A1 => n21253, A2 => n17829, Z => n11792);
   U5925 : OAI21_X1 port map( A1 => n32351, A2 => n32350, B => n31614, ZN => 
                           n17215);
   U5927 : NOR2_X1 port map( A1 => n33684, A2 => n33683, ZN => n33682);
   U5928 : NOR2_X1 port map( A1 => n21284, A2 => n16473, ZN => n7344);
   U5939 : NAND2_X1 port map( A1 => n34121, A2 => n30755, ZN => n27303);
   U5948 : BUF_X2 port map( I => n10787, Z => n9518);
   U5949 : INV_X1 port map( I => n32239, ZN => n13506);
   U5950 : BUF_X2 port map( I => n17144, Z => n31614);
   U5954 : BUF_X2 port map( I => n8813, Z => n7690);
   U5960 : CLKBUF_X2 port map( I => n21224, Z => n5595);
   U5965 : OR2_X1 port map( A1 => n15734, A2 => n15733, Z => n21362);
   U5966 : INV_X1 port map( I => n602, ZN => n33311);
   U5968 : CLKBUF_X4 port map( I => n8434, Z => n32452);
   U5970 : BUF_X4 port map( I => n21266, Z => n31965);
   U5976 : CLKBUF_X2 port map( I => n4858, Z => n32310);
   U5978 : CLKBUF_X2 port map( I => n20766, Z => n33969);
   U5980 : CLKBUF_X2 port map( I => n7653, Z => n32581);
   U5982 : INV_X1 port map( I => n20742, ZN => n20386);
   U5984 : CLKBUF_X2 port map( I => n20961, Z => n32749);
   U5986 : INV_X1 port map( I => n7294, ZN => n33234);
   U5987 : INV_X1 port map( I => n32996, ZN => n7800);
   U5989 : INV_X2 port map( I => n20913, ZN => n31966);
   U6013 : NOR2_X1 port map( A1 => n33899, A2 => n30952, ZN => n4909);
   U6018 : NOR2_X1 port map( A1 => n28135, A2 => n2203, ZN => n33899);
   U6026 : INV_X1 port map( I => n33944, ZN => n34155);
   U6032 : NAND2_X1 port map( A1 => n32277, A2 => n2237, ZN => n32276);
   U6034 : NAND2_X1 port map( A1 => n33341, A2 => n31961, ZN => n19454);
   U6037 : INV_X1 port map( I => n33193, ZN => n33192);
   U6039 : OAI21_X1 port map( A1 => n20216, A2 => n8998, B => n33639, ZN => 
                           n20218);
   U6040 : INV_X1 port map( I => n9808, ZN => n33307);
   U6047 : CLKBUF_X8 port map( I => n3086, Z => n31967);
   U6048 : CLKBUF_X8 port map( I => n29337, Z => n32504);
   U6049 : NOR2_X1 port map( A1 => n20193, A2 => n20192, ZN => n32939);
   U6050 : CLKBUF_X1 port map( I => n9352, Z => n34132);
   U6060 : INV_X1 port map( I => n31863, ZN => n33195);
   U6066 : INV_X4 port map( I => n30504, ZN => n31968);
   U6067 : CLKBUF_X2 port map( I => n20344, Z => n34013);
   U6070 : CLKBUF_X2 port map( I => n27697, Z => n33116);
   U6072 : BUF_X2 port map( I => n7292, Z => n31811);
   U6073 : NAND2_X1 port map( A1 => n34105, A2 => n14479, ZN => n29920);
   U6074 : AOI22_X1 port map( A1 => n30404, A2 => n1035, B1 => n19562, B2 => 
                           n11624, ZN => n33249);
   U6078 : CLKBUF_X2 port map( I => n20526, Z => n33222);
   U6081 : AND2_X1 port map( A1 => n29914, A2 => n17497, Z => n20438);
   U6084 : NAND2_X1 port map( A1 => n3790, A2 => n33769, ZN => n33768);
   U6089 : OAI21_X1 port map( A1 => n31988, A2 => n32371, B => n32416, ZN => 
                           n19839);
   U6097 : NAND2_X1 port map( A1 => n19528, A2 => n1617, ZN => n32740);
   U6099 : NAND2_X1 port map( A1 => n6929, A2 => n6930, ZN => n33896);
   U6101 : INV_X4 port map( I => n7762, ZN => n31969);
   U6106 : NAND2_X1 port map( A1 => n30614, A2 => n4201, ZN => n33037);
   U6111 : NOR2_X1 port map( A1 => n19939, A2 => n32109, ZN => n5694);
   U6113 : BUF_X2 port map( I => n20110, Z => n32408);
   U6115 : BUF_X1 port map( I => n13852, Z => n29233);
   U6118 : CLKBUF_X2 port map( I => n12008, Z => n34108);
   U6119 : BUF_X2 port map( I => n577, Z => n27832);
   U6131 : CLKBUF_X1 port map( I => n10426, Z => n32891);
   U6133 : BUF_X2 port map( I => n11630, Z => n33419);
   U6152 : BUF_X2 port map( I => n20108, Z => n16243);
   U6157 : CLKBUF_X2 port map( I => n7896, Z => n32184);
   U6161 : CLKBUF_X2 port map( I => n33339, Z => n32809);
   U6167 : INV_X1 port map( I => n19749, ZN => n32206);
   U6170 : BUF_X2 port map( I => n19494, Z => n207);
   U6171 : NAND2_X1 port map( A1 => n32758, A2 => n13494, ZN => n9080);
   U6172 : OAI21_X1 port map( A1 => n33825, A2 => n26350, B => n33824, ZN => 
                           n17509);
   U6174 : NAND2_X1 port map( A1 => n33231, A2 => n33230, ZN => n10741);
   U6175 : NAND2_X1 port map( A1 => n18360, A2 => n826, ZN => n32675);
   U6178 : NAND2_X1 port map( A1 => n32293, A2 => n32292, ZN => n13706);
   U6179 : NAND2_X1 port map( A1 => n29731, A2 => n29730, ZN => n32676);
   U6185 : NAND2_X1 port map( A1 => n27274, A2 => n27273, ZN => n33229);
   U6190 : NAND2_X1 port map( A1 => n17510, A2 => n26350, ZN => n33824);
   U6194 : INV_X1 port map( I => n19363, ZN => n32290);
   U6199 : CLKBUF_X2 port map( I => n30995, Z => n32788);
   U6206 : CLKBUF_X2 port map( I => n19262, Z => n33206);
   U6210 : OR2_X1 port map( A1 => n1883, A2 => n16699, Z => n9083);
   U6242 : NAND2_X1 port map( A1 => n8662, A2 => n19178, ZN => n33228);
   U6244 : AND2_X1 port map( A1 => n8379, A2 => n2902, Z => n32060);
   U6248 : CLKBUF_X2 port map( I => n19123, Z => n27033);
   U6252 : CLKBUF_X8 port map( I => n19314, Z => n31970);
   U6254 : INV_X2 port map( I => n19021, ZN => n19288);
   U6258 : NAND2_X1 port map( A1 => n15859, A2 => n30116, ZN => n32720);
   U6275 : NAND2_X1 port map( A1 => n18508, A2 => n18509, ZN => n32439);
   U6278 : OR2_X1 port map( A1 => n12648, A2 => n13016, Z => n13014);
   U6283 : NAND2_X1 port map( A1 => n33422, A2 => n33421, ZN => n27253);
   U6290 : NAND2_X1 port map( A1 => n29492, A2 => n18640, ZN => n8736);
   U6291 : NOR2_X1 port map( A1 => n9420, A2 => n14344, ZN => n32097);
   U6292 : AND2_X1 port map( A1 => n13554, A2 => n18510, Z => n32003);
   U6302 : NAND2_X1 port map( A1 => n13016, A2 => n32901, ZN => n32786);
   U6312 : INV_X1 port map( I => n18726, ZN => n33422);
   U6315 : INV_X1 port map( I => n17360, ZN => n33208);
   U6320 : INV_X4 port map( I => n8756, ZN => n31971);
   U6332 : INV_X1 port map( I => n14666, ZN => n18516);
   U6335 : CLKBUF_X2 port map( I => n11460, Z => n33548);
   U6338 : BUF_X2 port map( I => n18831, Z => n13846);
   U6342 : INV_X4 port map( I => n29315, ZN => n31972);
   U6344 : CLKBUF_X2 port map( I => n13445, Z => n33941);
   U6345 : INV_X1 port map( I => n25570, ZN => n32796);
   U6346 : INV_X1 port map( I => n25929, ZN => n32130);
   U6348 : CLKBUF_X2 port map( I => n17168, Z => n9);
   U6349 : CLKBUF_X1 port map( I => n493, Z => n171);
   U6360 : CLKBUF_X2 port map( I => n18862, Z => n33205);
   U6362 : INV_X1 port map( I => n24759, ZN => n33693);
   U6364 : NAND2_X1 port map( A1 => n10669, A2 => n18677, ZN => n10670);
   U6365 : INV_X1 port map( I => n16572, ZN => n33998);
   U6366 : CLKBUF_X2 port map( I => n18548, Z => n16122);
   U6367 : INV_X1 port map( I => n18707, ZN => n18535);
   U6373 : NAND2_X1 port map( A1 => n11097, A2 => n882, ZN => n4070);
   U6378 : INV_X2 port map( I => n12290, ZN => n3218);
   U6384 : CLKBUF_X2 port map( I => n9930, Z => n32358);
   U6387 : CLKBUF_X1 port map( I => n29182, Z => n32143);
   U6400 : NOR2_X1 port map( A1 => n8788, A2 => n18714, ZN => n6590);
   U6402 : CLKBUF_X2 port map( I => n18588, Z => n28056);
   U6405 : NAND2_X1 port map( A1 => n5269, A2 => n18705, ZN => n4043);
   U6406 : CLKBUF_X4 port map( I => n18373, Z => n18805);
   U6409 : NOR2_X1 port map( A1 => n18722, A2 => n18580, ZN => n12190);
   U6411 : NOR2_X1 port map( A1 => n33310, A2 => n33309, ZN => n9668);
   U6413 : INV_X1 port map( I => n12074, ZN => n18609);
   U6415 : NAND2_X1 port map( A1 => n18633, A2 => n15888, ZN => n15841);
   U6416 : NOR2_X1 port map( A1 => n11390, A2 => n14926, ZN => n18659);
   U6417 : CLKBUF_X1 port map( I => n18323, Z => n18492);
   U6424 : NOR2_X1 port map( A1 => n10844, A2 => n959, ZN => n4267);
   U6425 : NAND2_X1 port map( A1 => n9766, A2 => n18797, ZN => n18796);
   U6434 : NAND2_X1 port map( A1 => n13200, A2 => n19180, ZN => n7751);
   U6436 : AOI21_X1 port map( A1 => n31903, A2 => n18563, B => n6256, ZN => 
                           n18565);
   U6439 : AOI21_X1 port map( A1 => n33040, A2 => n18695, B => n16569, ZN => 
                           n18391);
   U6444 : OAI21_X1 port map( A1 => n18318, A2 => n18634, B => n18711, ZN => 
                           n30175);
   U6449 : NAND2_X1 port map( A1 => n19057, A2 => n18994, ZN => n32182);
   U6460 : NAND2_X1 port map( A1 => n32219, A2 => n32218, ZN => n10192);
   U6461 : NAND3_X1 port map( A1 => n19181, A2 => n19178, A3 => n29769, ZN => 
                           n13009);
   U6464 : NOR2_X1 port map( A1 => n3784, A2 => n879, ZN => n32758);
   U6474 : INV_X1 port map( I => n32622, ZN => n8303);
   U6477 : INV_X1 port map( I => n30781, ZN => n1056);
   U6480 : NAND2_X1 port map( A1 => n28276, A2 => n1630, ZN => n9442);
   U6482 : NAND2_X1 port map( A1 => n19076, A2 => n19288, ZN => n18360);
   U6483 : INV_X2 port map( I => n16093, ZN => n1052);
   U6484 : INV_X1 port map( I => n14892, ZN => n18995);
   U6487 : NOR2_X1 port map( A1 => n19091, A2 => n19088, ZN => n31174);
   U6494 : INV_X2 port map( I => n19258, ZN => n744);
   U6499 : NOR2_X1 port map( A1 => n19198, A2 => n26417, ZN => n13891);
   U6507 : INV_X1 port map( I => n19103, ZN => n11713);
   U6511 : NOR2_X1 port map( A1 => n32932, A2 => n7492, ZN => n17677);
   U6512 : AOI21_X1 port map( A1 => n14625, A2 => n8379, B => n2901, ZN => 
                           n12850);
   U6515 : CLKBUF_X2 port map( I => n14812, Z => n12549);
   U6521 : OAI21_X1 port map( A1 => n19148, A2 => n19147, B => n19150, ZN => 
                           n18267);
   U6526 : OAI22_X1 port map( A1 => n18475, A2 => n16185, B1 => n18901, B2 => 
                           n4, ZN => n18476);
   U6529 : NAND2_X1 port map( A1 => n6578, A2 => n6577, ZN => n6576);
   U6534 : INV_X1 port map( I => n19520, ZN => n10026);
   U6538 : INV_X1 port map( I => n6731, ZN => n11320);
   U6544 : NAND2_X1 port map( A1 => n14736, A2 => n14130, ZN => n14735);
   U6545 : CLKBUF_X2 port map( I => n14094, Z => n32286);
   U6550 : NOR2_X1 port map( A1 => n33712, A2 => n33389, ZN => n11581);
   U6553 : INV_X1 port map( I => n15787, ZN => n29090);
   U6557 : CLKBUF_X1 port map( I => n5150, Z => n32918);
   U6560 : INV_X1 port map( I => n26300, ZN => n19722);
   U6574 : INV_X1 port map( I => n19466, ZN => n17342);
   U6577 : INV_X1 port map( I => n19542, ZN => n32231);
   U6582 : INV_X1 port map( I => n2362, ZN => n12796);
   U6583 : INV_X1 port map( I => n31922, ZN => n8292);
   U6588 : NOR2_X1 port map( A1 => n13591, A2 => n11198, ZN => n19828);
   U6591 : INV_X1 port map( I => n19746, ZN => n30435);
   U6592 : INV_X1 port map( I => n11052, ZN => n2679);
   U6596 : NAND2_X1 port map( A1 => n34103, A2 => n6532, ZN => n13657);
   U6600 : NAND2_X1 port map( A1 => n20056, A2 => n32326, ZN => n14099);
   U6604 : NAND2_X1 port map( A1 => n32746, A2 => n32745, ZN => n19977);
   U6605 : NAND2_X1 port map( A1 => n19833, A2 => n1169, ZN => n15174);
   U6606 : INV_X1 port map( I => n579, ZN => n7461);
   U6609 : NOR2_X1 port map( A1 => n27491, A2 => n19961, ZN => n20128);
   U6612 : INV_X1 port map( I => n1361, ZN => n9749);
   U6614 : INV_X1 port map( I => n1169, ZN => n15593);
   U6616 : NOR2_X1 port map( A1 => n27808, A2 => n20113, ZN => n14729);
   U6628 : NOR2_X1 port map( A1 => n29216, A2 => n19990, ZN => n34106);
   U6629 : INV_X1 port map( I => n9106, ZN => n31106);
   U6631 : CLKBUF_X2 port map( I => n20108, Z => n33848);
   U6638 : NOR2_X1 port map( A1 => n20097, A2 => n1041, ZN => n30693);
   U6639 : INV_X1 port map( I => n20054, ZN => n11893);
   U6641 : CLKBUF_X4 port map( I => n14458, Z => n14281);
   U6642 : CLKBUF_X4 port map( I => n11333, Z => n28293);
   U6643 : NAND2_X1 port map( A1 => n20104, A2 => n873, ZN => n15177);
   U6649 : NOR3_X1 port map( A1 => n19724, A2 => n16461, A3 => n1042, ZN => 
                           n30357);
   U6652 : INV_X1 port map( I => n19885, ZN => n19799);
   U6655 : NAND2_X1 port map( A1 => n29153, A2 => n576, ZN => n9171);
   U6656 : CLKBUF_X4 port map( I => n16625, Z => n29156);
   U6659 : INV_X2 port map( I => n16694, ZN => n1360);
   U6660 : OAI21_X1 port map( A1 => n4674, A2 => n6200, B => n6263, ZN => n3090
                           );
   U6678 : CLKBUF_X4 port map( I => n18089, Z => n161);
   U6682 : NAND2_X1 port map( A1 => n33569, A2 => n17945, ZN => n32673);
   U6689 : NAND2_X1 port map( A1 => n9031, A2 => n1042, ZN => n19941);
   U6690 : OAI21_X1 port map( A1 => n27788, A2 => n27787, B => n20157, ZN => 
                           n30996);
   U6691 : NAND2_X1 port map( A1 => n28685, A2 => n28684, ZN => n28683);
   U6692 : AOI21_X1 port map( A1 => n938, A2 => n20052, B => n939, ZN => n6929)
                           ;
   U6694 : NAND2_X1 port map( A1 => n8181, A2 => n16630, ZN => n32775);
   U6700 : OAI21_X1 port map( A1 => n20053, A2 => n1361, B => n8616, ZN => 
                           n15312);
   U6709 : INV_X1 port map( I => n10752, ZN => n33525);
   U6710 : AOI21_X1 port map( A1 => n27714, A2 => n27716, B => n30355, ZN => 
                           n26784);
   U6731 : OAI21_X1 port map( A1 => n19950, A2 => n17363, B => n729, ZN => n14)
                           ;
   U6733 : NAND2_X1 port map( A1 => n295, A2 => n1155, ZN => n20337);
   U6734 : INV_X1 port map( I => n20267, ZN => n14863);
   U6742 : NAND2_X1 port map( A1 => n31242, A2 => n15551, ZN => n11505);
   U6747 : NOR2_X1 port map( A1 => n20607, A2 => n20460, ZN => n20396);
   U6749 : INV_X1 port map( I => n20410, ZN => n28128);
   U6754 : NAND2_X1 port map( A1 => n8903, A2 => n8870, ZN => n4586);
   U6755 : NAND2_X1 port map( A1 => n4807, A2 => n20571, ZN => n29077);
   U6756 : NOR2_X1 port map( A1 => n33091, A2 => n20545, ZN => n13629);
   U6757 : CLKBUF_X4 port map( I => n20503, Z => n28376);
   U6761 : NAND2_X1 port map( A1 => n7242, A2 => n20228, ZN => n20227);
   U6764 : INV_X1 port map( I => n19956, ZN => n10380);
   U6765 : NOR2_X1 port map( A1 => n20489, A2 => n33307, ZN => n17897);
   U6776 : NAND3_X1 port map( A1 => n26567, A2 => n3462, A3 => n741, ZN => 
                           n19453);
   U6778 : CLKBUF_X2 port map( I => n7280, Z => n32481);
   U6779 : AOI22_X1 port map( A1 => n20251, A2 => n20510, B1 => n20509, B2 => 
                           n20435, ZN => n17974);
   U6782 : NAND2_X1 port map( A1 => n5471, A2 => n14179, ZN => n20376);
   U6785 : INV_X1 port map( I => n9986, ZN => n5589);
   U6786 : OAI21_X1 port map( A1 => n20366, A2 => n7577, B => n33843, ZN => 
                           n20367);
   U6788 : NOR2_X1 port map( A1 => n17329, A2 => n6531, ZN => n9774);
   U6789 : INV_X2 port map( I => n15005, ZN => n1352);
   U6800 : INV_X2 port map( I => n31533, ZN => n30869);
   U6805 : NAND2_X1 port map( A1 => n13629, A2 => n20335, ZN => n13628);
   U6806 : NAND2_X1 port map( A1 => n20297, A2 => n14836, ZN => n14835);
   U6810 : NAND3_X1 port map( A1 => n3944, A2 => n17975, A3 => n1355, ZN => 
                           n14471);
   U6813 : NAND2_X1 port map( A1 => n16004, A2 => n13786, ZN => n13782);
   U6814 : INV_X1 port map( I => n20900, ZN => n29167);
   U6819 : OAI21_X1 port map( A1 => n11303, A2 => n1156, B => n6616, ZN => 
                           n20636);
   U6823 : NAND2_X1 port map( A1 => n19454, A2 => n19453, ZN => n3307);
   U6825 : INV_X1 port map( I => n12258, ZN => n31860);
   U6826 : AOI21_X1 port map( A1 => n29623, A2 => n1352, B => n20419, ZN => 
                           n20421);
   U6828 : NAND2_X1 port map( A1 => n5781, A2 => n17497, ZN => n19956);
   U6839 : CLKBUF_X1 port map( I => n21044, Z => n30240);
   U6840 : INV_X1 port map( I => n20860, ZN => n12671);
   U6843 : CLKBUF_X2 port map( I => n20680, Z => n31233);
   U6844 : CLKBUF_X4 port map( I => n13864, Z => n28315);
   U6845 : INV_X1 port map( I => n21025, ZN => n8138);
   U6849 : INV_X1 port map( I => n17440, ZN => n33085);
   U6851 : INV_X1 port map( I => n30492, ZN => n20855);
   U6853 : INV_X1 port map( I => n28981, ZN => n33892);
   U6858 : CLKBUF_X1 port map( I => n13189, Z => n28400);
   U6859 : INV_X2 port map( I => n16526, ZN => n31729);
   U6860 : NAND2_X1 port map( A1 => n12037, A2 => n21270, ZN => n27270);
   U6872 : NAND2_X1 port map( A1 => n2738, A2 => n9133, ZN => n8792);
   U6881 : INV_X2 port map( I => n28287, ZN => n14563);
   U6882 : INV_X1 port map( I => n21210, ZN => n16743);
   U6889 : NAND2_X1 port map( A1 => n1022, A2 => n33684, ZN => n7757);
   U6902 : NOR2_X1 port map( A1 => n21085, A2 => n4755, ZN => n29750);
   U6904 : CLKBUF_X2 port map( I => n13989, Z => n32242);
   U6913 : INV_X2 port map( I => n11814, ZN => n13692);
   U6916 : OAI21_X1 port map( A1 => n33106, A2 => n21109, B => n33705, ZN => 
                           n10922);
   U6920 : NAND3_X1 port map( A1 => n32357, A2 => n17767, A3 => n21078, ZN => 
                           n26018);
   U6921 : NAND2_X1 port map( A1 => n30646, A2 => n14721, ZN => n17101);
   U6922 : NAND2_X1 port map( A1 => n21379, A2 => n17313, ZN => n2275);
   U6925 : NAND2_X1 port map( A1 => n16668, A2 => n13896, ZN => n15219);
   U6927 : NOR2_X1 port map( A1 => n13896, A2 => n21115, ZN => n29001);
   U6930 : NOR2_X1 port map( A1 => n20879, A2 => n20880, ZN => n29739);
   U6933 : INV_X1 port map( I => n929, ZN => n33454);
   U6939 : INV_X1 port map( I => n11942, ZN => n21431);
   U6941 : NOR2_X1 port map( A1 => n20941, A2 => n16629, ZN => n32980);
   U6942 : NAND2_X1 port map( A1 => n13022, A2 => n32647, ZN => n16117);
   U6944 : NAND2_X1 port map( A1 => n20945, A2 => n27503, ZN => n21183);
   U6945 : CLKBUF_X4 port map( I => n17731, Z => n33972);
   U6946 : NAND2_X1 port map( A1 => n21129, A2 => n21443, ZN => n32454);
   U6948 : NOR2_X1 port map( A1 => n21109, A2 => n1632, ZN => n5488);
   U6950 : NAND2_X1 port map( A1 => n14230, A2 => n21440, ZN => n34083);
   U6956 : NAND2_X1 port map( A1 => n27303, A2 => n27305, ZN => n26903);
   U6961 : NOR2_X1 port map( A1 => n6584, A2 => n9721, ZN => n14997);
   U6962 : NAND2_X1 port map( A1 => n7845, A2 => n1333, ZN => n4179);
   U6963 : NOR2_X1 port map( A1 => n27193, A2 => n32239, ZN => n6879);
   U6970 : NOR2_X1 port map( A1 => n11487, A2 => n33682, ZN => n31848);
   U6971 : NOR2_X1 port map( A1 => n11215, A2 => n28922, ZN => n28921);
   U6975 : OAI22_X1 port map( A1 => n10149, A2 => n3673, B1 => n2275, B2 => 
                           n7007, ZN => n31215);
   U6976 : NAND2_X1 port map( A1 => n21411, A2 => n5039, ZN => n2721);
   U6980 : NOR2_X1 port map( A1 => n33417, A2 => n33418, ZN => n32116);
   U6983 : OR3_X1 port map( A1 => n4683, A2 => n16639, A3 => n29255, Z => 
                           n34158);
   U6985 : NOR2_X1 port map( A1 => n4517, A2 => n21251, ZN => n4284);
   U6987 : OAI21_X1 port map( A1 => n21259, A2 => n16652, B => n8757, ZN => 
                           n6568);
   U6989 : INV_X2 port map( I => n16519, ZN => n3048);
   U6991 : NOR2_X1 port map( A1 => n17348, A2 => n32252, ZN => n3703);
   U6993 : NOR2_X1 port map( A1 => n15302, A2 => n15296, ZN => n10875);
   U6994 : NOR2_X1 port map( A1 => n338, A2 => n4234, ZN => n4391);
   U6996 : INV_X2 port map( I => n16668, ZN => n4989);
   U6998 : OAI22_X1 port map( A1 => n21586, A2 => n32252, B1 => n3680, B2 => 
                           n26337, ZN => n29595);
   U7002 : NOR2_X1 port map( A1 => n21659, A2 => n8784, ZN => n4117);
   U7003 : NAND2_X1 port map( A1 => n29434, A2 => n517, ZN => n21747);
   U7004 : NOR2_X1 port map( A1 => n7969, A2 => n7182, ZN => n7183);
   U7008 : INV_X1 port map( I => n21687, ZN => n21514);
   U7010 : NOR2_X1 port map( A1 => n5546, A2 => n4356, ZN => n8705);
   U7012 : NAND2_X1 port map( A1 => n5546, A2 => n14236, ZN => n21622);
   U7019 : NAND3_X1 port map( A1 => n30479, A2 => n21850, A3 => n21763, ZN => 
                           n10968);
   U7020 : NAND2_X1 port map( A1 => n21585, A2 => n15302, ZN => n21234);
   U7024 : AOI21_X1 port map( A1 => n4391, A2 => n13816, B => n27816, ZN => 
                           n6076);
   U7035 : INV_X1 port map( I => n8753, ZN => n10456);
   U7039 : CLKBUF_X2 port map( I => n28762, Z => n33468);
   U7041 : NAND3_X1 port map( A1 => n32321, A2 => n21830, A3 => n32320, ZN => 
                           n34001);
   U7045 : CLKBUF_X1 port map( I => n21789, Z => n27543);
   U7049 : NOR2_X1 port map( A1 => n16796, A2 => n16192, ZN => n22126);
   U7052 : AOI21_X1 port map( A1 => n2217, A2 => n16600, B => n21772, ZN => 
                           n12328);
   U7055 : NAND3_X1 port map( A1 => n864, A2 => n15864, A3 => n12278, ZN => 
                           n12277);
   U7057 : INV_X1 port map( I => n10205, ZN => n30407);
   U7058 : CLKBUF_X2 port map( I => n22227, Z => n33509);
   U7063 : NAND3_X1 port map( A1 => n11657, A2 => n11656, A3 => n14829, ZN => 
                           n17898);
   U7068 : AOI21_X1 port map( A1 => n4311, A2 => n6489, B => n4310, ZN => 
                           n21624);
   U7070 : INV_X1 port map( I => n22000, ZN => n21875);
   U7073 : INV_X1 port map( I => n6571, ZN => n33707);
   U7078 : INV_X1 port map( I => n9267, ZN => n11422);
   U7079 : INV_X1 port map( I => n9914, ZN => n32696);
   U7091 : INV_X1 port map( I => n26933, ZN => n32155);
   U7097 : NAND2_X1 port map( A1 => n31701, A2 => n10282, ZN => n32797);
   U7099 : INV_X1 port map( I => n15260, ZN => n30669);
   U7100 : NOR2_X1 port map( A1 => n31001, A2 => n26708, ZN => n22342);
   U7101 : INV_X1 port map( I => n22487, ZN => n1288);
   U7104 : INV_X1 port map( I => n17204, ZN => n22644);
   U7108 : OAI21_X1 port map( A1 => n9910, A2 => n29158, B => n33237, ZN => 
                           n31838);
   U7110 : CLKBUF_X2 port map( I => n29263, Z => n355);
   U7111 : CLKBUF_X4 port map( I => n1805, Z => n1633);
   U7116 : NOR2_X1 port map( A1 => n1294, A2 => n14253, ZN => n22594);
   U7117 : INV_X1 port map( I => n22622, ZN => n995);
   U7121 : INV_X1 port map( I => n22491, ZN => n17302);
   U7125 : AOI21_X1 port map( A1 => n16745, A2 => n8919, B => n32080, ZN => 
                           n8918);
   U7126 : NOR2_X1 port map( A1 => n22660, A2 => n809, ZN => n30334);
   U7127 : CLKBUF_X1 port map( I => n17518, Z => n14493);
   U7130 : CLKBUF_X2 port map( I => n22332, Z => n33964);
   U7131 : CLKBUF_X4 port map( I => n8275, Z => n1116);
   U7133 : NAND2_X1 port map( A1 => n26098, A2 => n1127, ZN => n13193);
   U7137 : NAND2_X1 port map( A1 => n22460, A2 => n16137, ZN => n22344);
   U7138 : NAND2_X1 port map( A1 => n27880, A2 => n28312, ZN => n33945);
   U7145 : INV_X1 port map( I => n12952, ZN => n22511);
   U7150 : INV_X1 port map( I => n32448, ZN => n1720);
   U7151 : NAND2_X1 port map( A1 => n16884, A2 => n22336, ZN => n26813);
   U7158 : OAI22_X1 port map( A1 => n11419, A2 => n22420, B1 => n31345, B2 => 
                           n11420, ZN => n3934);
   U7164 : NAND2_X1 port map( A1 => n13524, A2 => n12840, ZN => n32518);
   U7169 : CLKBUF_X2 port map( I => n16332, Z => n27402);
   U7173 : OAI22_X1 port map( A1 => n32680, A2 => n11629, B1 => n30205, B2 => 
                           n15581, ZN => n2135);
   U7175 : INV_X1 port map( I => n10206, ZN => n8801);
   U7177 : NAND2_X1 port map( A1 => n32955, A2 => n29495, ZN => n1580);
   U7180 : AOI22_X1 port map( A1 => n22688, A2 => n22332, B1 => n2417, B2 => 
                           n12733, ZN => n27034);
   U7181 : INV_X2 port map( I => n636, ZN => n857);
   U7189 : NAND2_X1 port map( A1 => n32823, A2 => n31963, ZN => n27368);
   U7193 : NAND2_X1 port map( A1 => n22475, A2 => n22377, ZN => n31143);
   U7198 : INV_X2 port map( I => n10862, ZN => n8912);
   U7200 : CLKBUF_X2 port map( I => n30868, Z => n32967);
   U7206 : NAND3_X1 port map( A1 => n903, A2 => n30564, A3 => n7848, ZN => 
                           n29722);
   U7209 : INV_X1 port map( I => n2635, ZN => n11298);
   U7213 : INV_X1 port map( I => n31566, ZN => n33591);
   U7216 : OAI22_X1 port map( A1 => n30455, A2 => n9954, B1 => n773, B2 => 
                           n6782, ZN => n10280);
   U7218 : AOI22_X1 port map( A1 => n22651, A2 => n4916, B1 => n22433, B2 => 
                           n14251, ZN => n1661);
   U7231 : INV_X4 port map( I => n27090, ZN => n22774);
   U7232 : INV_X2 port map( I => n17147, ZN => n5597);
   U7233 : INV_X1 port map( I => n14978, ZN => n22756);
   U7236 : INV_X1 port map( I => n3296, ZN => n33388);
   U7238 : CLKBUF_X4 port map( I => n12729, Z => n28314);
   U7243 : NAND2_X1 port map( A1 => n32704, A2 => n15718, ZN => n18239);
   U7244 : NOR2_X1 port map( A1 => n4750, A2 => n30234, ZN => n11540);
   U7245 : NAND2_X1 port map( A1 => n31937, A2 => n15501, ZN => n6350);
   U7248 : NAND2_X1 port map( A1 => n7004, A2 => n22971, ZN => n22805);
   U7249 : NOR2_X1 port map( A1 => n23112, A2 => n23111, ZN => n32525);
   U7252 : INV_X1 port map( I => n2449, ZN => n23031);
   U7253 : NAND2_X1 port map( A1 => n641, A2 => n22876, ZN => n22766);
   U7258 : NAND2_X1 port map( A1 => n6800, A2 => n1107, ZN => n12742);
   U7260 : OAI21_X1 port map( A1 => n28408, A2 => n6799, B => n1107, ZN => 
                           n6035);
   U7262 : NOR2_X1 port map( A1 => n4750, A2 => n22919, ZN => n10588);
   U7266 : INV_X1 port map( I => n28934, ZN => n22908);
   U7269 : NAND2_X1 port map( A1 => n6874, A2 => n2449, ZN => n6942);
   U7271 : NAND2_X1 port map( A1 => n31225, A2 => n15421, ZN => n22383);
   U7277 : CLKBUF_X4 port map( I => n4208, Z => n30960);
   U7278 : AOI21_X1 port map( A1 => n30904, A2 => n28659, B => n10360, ZN => 
                           n5571);
   U7279 : INV_X1 port map( I => n23183, ZN => n23241);
   U7284 : CLKBUF_X2 port map( I => n23209, Z => n34100);
   U7291 : INV_X1 port map( I => n33971, ZN => n1263);
   U7292 : OAI22_X1 port map( A1 => n33996, A2 => n34097, B1 => n22938, B2 => 
                           n29173, ZN => n16922);
   U7296 : INV_X1 port map( I => n16998, ZN => n30362);
   U7299 : AOI22_X1 port map( A1 => n26195, A2 => n10296, B1 => n32092, B2 => 
                           n30234, ZN => n10759);
   U7305 : INV_X1 port map( I => n22867, ZN => n33811);
   U7307 : CLKBUF_X2 port map( I => n5512, Z => n33380);
   U7311 : NAND2_X1 port map( A1 => n8381, A2 => n5211, ZN => n10349);
   U7312 : OAI21_X1 port map( A1 => n28970, A2 => n32868, B => n3160, ZN => 
                           n3159);
   U7314 : INV_X1 port map( I => n11249, ZN => n32302);
   U7315 : INV_X1 port map( I => n4047, ZN => n13888);
   U7319 : INV_X1 port map( I => n23153, ZN => n33590);
   U7326 : NOR2_X1 port map( A1 => n23938, A2 => n662, ZN => n27266);
   U7327 : NOR2_X1 port map( A1 => n23951, A2 => n16431, ZN => n3759);
   U7329 : NOR2_X1 port map( A1 => n23691, A2 => n23857, ZN => n23570);
   U7330 : CLKBUF_X4 port map( I => n17285, Z => n14975);
   U7338 : NAND2_X1 port map( A1 => n27266, A2 => n23939, ZN => n33626);
   U7342 : INV_X1 port map( I => n23706, ZN => n33461);
   U7343 : INV_X1 port map( I => n10772, ZN => n9328);
   U7344 : OAI21_X1 port map( A1 => n23933, A2 => n29269, B => n23527, ZN => 
                           n13103);
   U7353 : BUF_X2 port map( I => n8270, Z => n32602);
   U7355 : INV_X1 port map( I => n12104, ZN => n33252);
   U7358 : NOR2_X1 port map( A1 => n11392, A2 => n23653, ZN => n6992);
   U7362 : NAND2_X1 port map( A1 => n23777, A2 => n23778, ZN => n32972);
   U7367 : NOR2_X1 port map( A1 => n23858, A2 => n2023, ZN => n1875);
   U7370 : INV_X1 port map( I => n651, ZN => n977);
   U7372 : INV_X1 port map( I => n16686, ZN => n1250);
   U7374 : NOR2_X1 port map( A1 => n4743, A2 => n23638, ZN => n18054);
   U7375 : INV_X2 port map( I => n18204, ZN => n28265);
   U7378 : NAND2_X1 port map( A1 => n23569, A2 => n23914, ZN => n32843);
   U7381 : AOI21_X1 port map( A1 => n13521, A2 => n29271, B => n23795, ZN => 
                           n16212);
   U7382 : INV_X1 port map( I => n32986, ZN => n23915);
   U7384 : OAI21_X1 port map( A1 => n23776, A2 => n31810, B => n23775, ZN => 
                           n23654);
   U7392 : NAND2_X1 port map( A1 => n1099, A2 => n23755, ZN => n14943);
   U7393 : NOR2_X1 port map( A1 => n11589, A2 => n16424, ZN => n33786);
   U7402 : CLKBUF_X1 port map( I => n666, Z => n28365);
   U7404 : CLKBUF_X4 port map( I => n10187, Z => n29198);
   U7410 : INV_X1 port map( I => n23867, ZN => n23637);
   U7412 : INV_X1 port map( I => n23906, ZN => n17288);
   U7415 : OAI22_X1 port map( A1 => n10384, A2 => n16388, B1 => n2460, B2 => 
                           n11240, ZN => n10382);
   U7420 : INV_X1 port map( I => n8547, ZN => n1252);
   U7428 : NOR2_X1 port map( A1 => n23826, A2 => n29839, ZN => n8472);
   U7431 : NAND2_X1 port map( A1 => n23939, A2 => n33499, ZN => n30828);
   U7433 : NAND2_X1 port map( A1 => n24095, A2 => n14195, ZN => n1619);
   U7442 : OAI21_X1 port map( A1 => n11708, A2 => n6272, B => n4111, ZN => 
                           n23671);
   U7444 : OAI22_X1 port map( A1 => n23760, A2 => n26115, B1 => n23759, B2 => 
                           n13905, ZN => n32336);
   U7445 : CLKBUF_X4 port map( I => n11516, Z => n1920);
   U7446 : INV_X1 port map( I => n29370, ZN => n33603);
   U7449 : NOR2_X1 port map( A1 => n23773, A2 => n23775, ZN => n16628);
   U7451 : NAND2_X1 port map( A1 => n23961, A2 => n13343, ZN => n6336);
   U7453 : CLKBUF_X4 port map( I => n10302, Z => n6001);
   U7456 : NAND2_X1 port map( A1 => n24204, A2 => n7935, ZN => n9202);
   U7459 : NAND2_X1 port map( A1 => n24114, A2 => n24283, ZN => n23549);
   U7466 : CLKBUF_X1 port map( I => n30191, Z => n32520);
   U7467 : NOR2_X1 port map( A1 => n13378, A2 => n2558, ZN => n4664);
   U7469 : INV_X2 port map( I => n6476, ZN => n24253);
   U7473 : NAND3_X1 port map( A1 => n8086, A2 => n24209, A3 => n8165, ZN => 
                           n17676);
   U7481 : AOI21_X1 port map( A1 => n24125, A2 => n24124, B => n24182, ZN => 
                           n24126);
   U7484 : OAI21_X1 port map( A1 => n24176, A2 => n11200, B => n17566, ZN => 
                           n24179);
   U7487 : INV_X1 port map( I => n24568, ZN => n30127);
   U7491 : NAND2_X1 port map( A1 => n3549, A2 => n16573, ZN => n2361);
   U7492 : NAND3_X1 port map( A1 => n13660, A2 => n11937, A3 => n24198, ZN => 
                           n32870);
   U7494 : NAND2_X1 port map( A1 => n11439, A2 => n11440, ZN => n24776);
   U7500 : INV_X1 port map( I => n18144, ZN => n33028);
   U7501 : CLKBUF_X2 port map( I => n24811, Z => n32814);
   U7502 : CLKBUF_X2 port map( I => n3694, Z => n32623);
   U7503 : INV_X1 port map( I => n8152, ZN => n24450);
   U7513 : INV_X1 port map( I => n24525, ZN => n33090);
   U7516 : NAND2_X1 port map( A1 => n4886, A2 => n32760, ZN => n10629);
   U7517 : NAND2_X1 port map( A1 => n5254, A2 => n11045, ZN => n5273);
   U7522 : INV_X1 port map( I => n15318, ZN => n29630);
   U7527 : INV_X1 port map( I => n25565, ZN => n6071);
   U7528 : INV_X1 port map( I => n10248, ZN => n13532);
   U7529 : NAND2_X1 port map( A1 => n32878, A2 => n4885, ZN => n10890);
   U7530 : INV_X1 port map( I => n25887, ZN => n5553);
   U7535 : NOR2_X1 port map( A1 => n25013, A2 => n24977, ZN => n6364);
   U7540 : CLKBUF_X2 port map( I => n4885, Z => n32106);
   U7541 : NAND2_X1 port map( A1 => n25582, A2 => n11900, ZN => n8712);
   U7544 : OAI22_X1 port map( A1 => n25411, A2 => n752, B1 => n25412, B2 => 
                           n11366, ZN => n1463);
   U7545 : CLKBUF_X2 port map( I => n11957, Z => n33976);
   U7546 : CLKBUF_X4 port map( I => n24181, Z => n25897);
   U7547 : NAND2_X1 port map( A1 => n32590, A2 => n25889, ZN => n32589);
   U7548 : INV_X1 port map( I => n24977, ZN => n14993);
   U7554 : NAND2_X1 port map( A1 => n25200, A2 => n12476, ZN => n17928);
   U7555 : NAND3_X1 port map( A1 => n1213, A2 => n25239, A3 => n14922, ZN => 
                           n31545);
   U7558 : INV_X1 port map( I => n28096, ZN => n25713);
   U7560 : INV_X1 port map( I => n17814, ZN => n25904);
   U7561 : NOR2_X1 port map( A1 => n25897, A2 => n9932, ZN => n10136);
   U7564 : NAND2_X1 port map( A1 => n27262, A2 => n10504, ZN => n30656);
   U7566 : OAI21_X1 port map( A1 => n32668, A2 => n32667, B => n7081, ZN => 
                           n28117);
   U7568 : AOI21_X1 port map( A1 => n25866, A2 => n25889, B => n1214, ZN => 
                           n6851);
   U7571 : BUF_X1 port map( I => n12676, Z => n33904);
   U7572 : NOR2_X1 port map( A1 => n27757, A2 => n27758, ZN => n33987);
   U7574 : CLKBUF_X2 port map( I => n25385, Z => n6551);
   U7578 : NAND2_X1 port map( A1 => n32825, A2 => n25866, ZN => n32312);
   U7580 : NAND3_X1 port map( A1 => n9495, A2 => n29331, A3 => n13640, ZN => 
                           n26992);
   U7591 : INV_X2 port map( I => n7554, ZN => n14810);
   U7594 : NAND2_X1 port map( A1 => n12864, A2 => n13483, ZN => n6391);
   U7597 : INV_X1 port map( I => n965, ZN => n24946);
   U7601 : INV_X1 port map( I => n1209, ZN => n33400);
   U7604 : NAND2_X1 port map( A1 => n13124, A2 => n789, ZN => n5786);
   U7608 : NOR2_X1 port map( A1 => n25127, A2 => n1075, ZN => n14638);
   U7612 : OAI22_X1 port map( A1 => n25272, A2 => n28532, B1 => n25271, B2 => 
                           n30281, ZN => n25273);
   U7615 : NAND2_X1 port map( A1 => n25041, A2 => n25052, ZN => n25048);
   U7619 : OAI21_X1 port map( A1 => n25041, A2 => n25029, B => n25060, ZN => 
                           n25035);
   U7620 : BUF_X2 port map( I => Key(6), Z => n25832);
   U7623 : AOI21_X1 port map( A1 => n5072, A2 => n24994, B => n964, ZN => 
                           n14318);
   U7627 : INV_X1 port map( I => n25418, ZN => n33946);
   U7629 : INV_X1 port map( I => n13684, ZN => n1076);
   U7634 : CLKBUF_X1 port map( I => Key(143), Z => n25801);
   U7635 : CLKBUF_X1 port map( I => Key(179), Z => n24937);
   U7639 : AOI21_X1 port map( A1 => n2265, A2 => n714, B => n2263, ZN => n2262)
                           ;
   U7648 : INV_X1 port map( I => n16525, ZN => n17914);
   U7651 : AND2_X1 port map( A1 => n15804, A2 => n13329, Z => n31973);
   U7675 : AND2_X2 port map( A1 => n11090, A2 => n11900, Z => n31974);
   U7678 : AND2_X1 port map( A1 => n32341, A2 => n20603, Z => n31976);
   U7681 : OR2_X1 port map( A1 => n24974, A2 => n11898, Z => n31977);
   U7682 : AND2_X2 port map( A1 => n29322, A2 => n14095, Z => n31978);
   U7686 : AND3_X2 port map( A1 => n32592, A2 => n32591, A3 => n32589, Z => 
                           n31979);
   U7687 : AND2_X2 port map( A1 => n29182, A2 => n18727, Z => n31980);
   U7689 : OR3_X1 port map( A1 => n9066, A2 => n12982, A3 => n24309, Z => 
                           n31983);
   U7691 : AND2_X1 port map( A1 => n1099, A2 => n27799, Z => n31984);
   U7694 : AND2_X2 port map( A1 => n29308, A2 => n29315, Z => n31987);
   U7695 : AND2_X1 port map( A1 => n20136, A2 => n19834, Z => n31988);
   U7696 : AND2_X1 port map( A1 => n3687, A2 => n32602, Z => n31990);
   U7698 : AND2_X1 port map( A1 => n19262, A2 => n19257, Z => n31992);
   U7702 : AND2_X2 port map( A1 => n16694, A2 => n19942, Z => n31993);
   U7703 : AND2_X1 port map( A1 => n25403, A2 => n16650, Z => n31994);
   U7704 : AND2_X1 port map( A1 => n6408, A2 => n16906, Z => n31995);
   U7705 : AND2_X1 port map( A1 => n7969, A2 => n31960, Z => n31996);
   U7709 : OR2_X1 port map( A1 => n14976, A2 => n149, Z => n31998);
   U7713 : AND2_X1 port map( A1 => n21251, A2 => n21249, Z => n31999);
   U7715 : AND2_X1 port map( A1 => n10947, A2 => n13747, Z => n32000);
   U7716 : OR2_X1 port map( A1 => n29574, A2 => n21303, Z => n32001);
   U7718 : AND2_X1 port map( A1 => n10295, A2 => n11317, Z => n32002);
   U7719 : OR2_X2 port map( A1 => n16732, A2 => n16854, Z => n32005);
   U7720 : OR2_X1 port map( A1 => n846, A2 => n16467, Z => n32006);
   U7723 : OR2_X1 port map( A1 => n28263, A2 => n907, Z => n32007);
   U7724 : OR2_X1 port map( A1 => n11392, A2 => n1252, Z => n32008);
   U7726 : AND2_X1 port map( A1 => n15421, A2 => n16078, Z => n32010);
   U7732 : OR2_X2 port map( A1 => n29334, A2 => n4886, Z => n32012);
   U7734 : AND2_X1 port map( A1 => n913, A2 => n13332, Z => n32013);
   U7735 : OR2_X2 port map( A1 => n3005, A2 => n8616, Z => n32014);
   U7742 : XNOR2_X1 port map( A1 => n23358, A2 => n25519, ZN => n32015);
   U7746 : OR2_X1 port map( A1 => n24125, A2 => n10381, Z => n32016);
   U7747 : AND3_X1 port map( A1 => n9934, A2 => n9962, A3 => n24201, Z => 
                           n32017);
   U7750 : AND2_X1 port map( A1 => n29314, A2 => n31867, Z => n32018);
   U7751 : AND2_X1 port map( A1 => n23881, A2 => n8544, Z => n32019);
   U7752 : OR2_X2 port map( A1 => n22491, A2 => n645, Z => n32021);
   U7753 : XNOR2_X1 port map( A1 => n33749, A2 => n1396, ZN => n32022);
   U7754 : AND2_X1 port map( A1 => n10252, A2 => n752, Z => n32023);
   U7755 : XNOR2_X1 port map( A1 => n14952, A2 => n24426, ZN => n32024);
   U7768 : XNOR2_X1 port map( A1 => n20786, A2 => n1393, ZN => n32025);
   U7769 : XNOR2_X1 port map( A1 => n14120, A2 => n16622, ZN => n32026);
   U7772 : XOR2_X1 port map( A1 => n29885, A2 => n16655, Z => n32027);
   U7773 : OR2_X1 port map( A1 => n2522, A2 => n15322, Z => n32031);
   U7774 : OR2_X2 port map( A1 => n7292, A2 => n20460, Z => n32033);
   U7779 : XNOR2_X1 port map( A1 => Plaintext(50), A2 => Key(50), ZN => n32034)
                           ;
   U7780 : AND2_X1 port map( A1 => n25966, A2 => n9115, Z => n32035);
   U7782 : AND2_X1 port map( A1 => n24201, A2 => n6911, Z => n32036);
   U7788 : AND2_X1 port map( A1 => n1567, A2 => n8210, Z => n32038);
   U7789 : OR2_X2 port map( A1 => n21532, A2 => n30389, Z => n32039);
   U7790 : OR2_X2 port map( A1 => n18221, A2 => n14487, Z => n32040);
   U7794 : INV_X2 port map( I => n9951, ZN => n985);
   U7797 : NOR2_X1 port map( A1 => n22332, A2 => n4330, ZN => n32042);
   U7799 : AND2_X1 port map( A1 => n30987, A2 => n32201, Z => n32043);
   U7801 : XNOR2_X1 port map( A1 => n19712, A2 => n25878, ZN => n32044);
   U7802 : AND2_X2 port map( A1 => n522, A2 => n7513, Z => n32045);
   U7804 : XNOR2_X1 port map( A1 => n19741, A2 => n24707, ZN => n32046);
   U7807 : XNOR2_X1 port map( A1 => n2073, A2 => n1393, ZN => n32047);
   U7809 : OR2_X1 port map( A1 => n22785, A2 => n3909, Z => n32048);
   U7814 : CLKBUF_X4 port map( I => n564, Z => n4215);
   U7817 : INV_X2 port map( I => n21812, ZN => n1132);
   U7819 : AND2_X1 port map( A1 => n24248, A2 => n28553, Z => n32049);
   U7822 : INV_X1 port map( I => n7292, ZN => n1356);
   U7823 : INV_X1 port map( I => n28945, ZN => n33182);
   U7824 : OR2_X2 port map( A1 => n30578, A2 => n33387, Z => n32050);
   U7826 : INV_X1 port map( I => n17316, ZN => n33688);
   U7827 : XOR2_X1 port map( A1 => Plaintext(6), A2 => Key(6), Z => n32051);
   U7830 : AND2_X2 port map( A1 => n30572, A2 => n27585, Z => n32052);
   U7834 : XNOR2_X1 port map( A1 => n19744, A2 => n19743, ZN => n32053);
   U7836 : OR2_X1 port map( A1 => n8212, A2 => n2207, Z => n32054);
   U7838 : CLKBUF_X4 port map( I => n18649, Z => n16474);
   U7840 : XOR2_X1 port map( A1 => n17284, A2 => n27268, Z => n32055);
   U7843 : AND2_X1 port map( A1 => n11444, A2 => n4835, Z => n32056);
   U7850 : XOR2_X1 port map( A1 => n11604, A2 => n1653, Z => n32058);
   U7852 : AND2_X2 port map( A1 => n2001, A2 => n2000, Z => n32059);
   U7853 : CLKBUF_X2 port map( I => n9320, Z => n26587);
   U7855 : INV_X1 port map( I => n19319, ZN => n33432);
   U7857 : OR2_X1 port map( A1 => n9025, A2 => n8870, Z => n32061);
   U7858 : AND2_X2 port map( A1 => n4775, A2 => n3421, Z => n32062);
   U7860 : OR2_X2 port map( A1 => n31656, A2 => n17295, Z => n32063);
   U7863 : OR2_X1 port map( A1 => n12548, A2 => n19156, Z => n32064);
   U7864 : INV_X1 port map( I => n34010, ZN => n29440);
   U7866 : NOR2_X1 port map( A1 => n10714, A2 => n9319, ZN => n34010);
   U7870 : XNOR2_X1 port map( A1 => n9141, A2 => n20792, ZN => n32065);
   U7871 : INV_X1 port map( I => n17144, ZN => n21218);
   U7872 : XNOR2_X1 port map( A1 => n20807, A2 => n20697, ZN => n32067);
   U7873 : INV_X1 port map( I => n11630, ZN => n17243);
   U7874 : NOR2_X1 port map( A1 => n20208, A2 => n20207, ZN => n32399);
   U7875 : INV_X1 port map( I => n16489, ZN => n938);
   U7881 : INV_X1 port map( I => n33856, ZN => n34154);
   U7883 : INV_X1 port map( I => n8813, ZN => n14721);
   U7892 : AND2_X2 port map( A1 => n12227, A2 => n20361, Z => n32068);
   U7893 : XNOR2_X1 port map( A1 => n20740, A2 => n20739, ZN => n32069);
   U7894 : INV_X1 port map( I => n21952, ZN => n32695);
   U7897 : XNOR2_X1 port map( A1 => n20862, A2 => n13357, ZN => n32070);
   U7905 : INV_X1 port map( I => n28254, ZN => n21257);
   U7909 : CLKBUF_X2 port map( I => n28254, Z => n33684);
   U7912 : INV_X1 port map( I => n21392, ZN => n21368);
   U7918 : XNOR2_X1 port map( A1 => n26785, A2 => n22220, ZN => n32072);
   U7919 : XNOR2_X1 port map( A1 => n13857, A2 => n13856, ZN => n32074);
   U7924 : AND2_X1 port map( A1 => n32815, A2 => n16117, Z => n32075);
   U7925 : INV_X2 port map( I => n13382, ZN => n1127);
   U7926 : OR2_X2 port map( A1 => n6765, A2 => n17888, Z => n32076);
   U7929 : XNOR2_X1 port map( A1 => n623, A2 => n22022, ZN => n32077);
   U7930 : XOR2_X1 port map( A1 => n33202, A2 => n3353, Z => n32078);
   U7931 : INV_X1 port map( I => n22148, ZN => n22221);
   U7932 : XNOR2_X1 port map( A1 => n6811, A2 => n6809, ZN => n32081);
   U7933 : XNOR2_X1 port map( A1 => n4589, A2 => n4590, ZN => n32082);
   U7937 : XNOR2_X1 port map( A1 => n22312, A2 => n21050, ZN => n32083);
   U7938 : AND2_X2 port map( A1 => n15314, A2 => n15316, Z => n32084);
   U7941 : INV_X1 port map( I => n10402, ZN => n28924);
   U7946 : INV_X1 port map( I => n26292, ZN => n33237);
   U7947 : INV_X1 port map( I => n25963, ZN => n32830);
   U7954 : XNOR2_X1 port map( A1 => n7623, A2 => n7622, ZN => n32085);
   U7955 : INV_X2 port map( I => n22425, ZN => n1728);
   U7959 : AND2_X1 port map( A1 => n28865, A2 => n22467, Z => n32087);
   U7961 : INV_X1 port map( I => n622, ZN => n11892);
   U7962 : AND2_X2 port map( A1 => n15806, A2 => n4580, Z => n32089);
   U7963 : NAND3_X1 port map( A1 => n22398, A2 => n708, A3 => n17853, ZN => 
                           n32090);
   U7964 : AND2_X1 port map( A1 => n30234, A2 => n30868, Z => n32091);
   U7967 : NAND2_X1 port map( A1 => n9798, A2 => n28608, ZN => n32093);
   U7968 : INV_X1 port map( I => n23886, ZN => n23889);
   U7969 : INV_X2 port map( I => n14540, ZN => n1271);
   U7971 : CLKBUF_X2 port map( I => n13704, Z => n13525);
   U7973 : AND3_X2 port map( A1 => n30651, A2 => n10226, A3 => n7935, Z => 
                           n32094);
   U7977 : CLKBUF_X1 port map( I => n24870, Z => n25152);
   U7978 : AND2_X1 port map( A1 => n24143, A2 => n24142, Z => n32095);
   U7979 : INV_X1 port map( I => n33235, ZN => n736);
   U7980 : INV_X1 port map( I => n24242, ZN => n33540);
   U7981 : XNOR2_X1 port map( A1 => n6898, A2 => n33359, ZN => n32096);
   U7984 : INV_X1 port map( I => n13232, ZN => n14112);
   U7985 : INV_X1 port map( I => n24719, ZN => n33155);
   U7991 : CLKBUF_X2 port map( I => n24719, Z => n25866);
   U7992 : INV_X1 port map( I => n31783, ZN => n25303);
   U8000 : XOR2_X1 port map( A1 => n1994, A2 => n19627, Z => n12413);
   U8003 : NAND2_X2 port map( A1 => n5223, A2 => n33719, ZN => n1994);
   U8007 : NAND2_X1 port map( A1 => n7310, A2 => n3909, ZN => n5832);
   U8010 : NAND2_X2 port map( A1 => n28083, A2 => n4221, ZN => n3909);
   U8012 : INV_X1 port map( I => n27728, ZN => n19464);
   U8013 : XNOR2_X1 port map( A1 => n3964, A2 => n19400, ZN => n27728);
   U8015 : NOR2_X2 port map( A1 => n14342, A2 => n32097, ZN => n14624);
   U8020 : OAI21_X2 port map( A1 => n32071, A2 => n30223, B => n21653, ZN => 
                           n30846);
   U8021 : XOR2_X1 port map( A1 => n8583, A2 => n12539, Z => n13455);
   U8023 : NAND2_X2 port map( A1 => n21410, A2 => n10113, ZN => n33886);
   U8024 : NAND2_X2 port map( A1 => n33888, A2 => n31835, ZN => n21410);
   U8026 : NAND3_X2 port map( A1 => n32706, A2 => n28206, A3 => n22651, ZN => 
                           n26568);
   U8028 : XOR2_X1 port map( A1 => n22136, A2 => n32098, Z => n32631);
   U8031 : XOR2_X1 port map( A1 => n22134, A2 => n32099, Z => n32098);
   U8034 : AOI21_X1 port map( A1 => n31904, A2 => n32101, B => n4193, ZN => 
                           n31216);
   U8035 : OR2_X1 port map( A1 => n7586, A2 => n5713, Z => n32101);
   U8037 : NAND2_X2 port map( A1 => n10922, A2 => n31677, ZN => n1313);
   U8042 : NOR2_X1 port map( A1 => n601, A2 => n1736, ZN => n33705);
   U8044 : XOR2_X1 port map( A1 => n3099, A2 => n32103, Z => n7119);
   U8045 : XOR2_X1 port map( A1 => n33892, A2 => n9464, Z => n32103);
   U8046 : XOR2_X1 port map( A1 => n9627, A2 => n20869, Z => n28981);
   U8050 : NAND2_X2 port map( A1 => n28733, A2 => n30197, ZN => n9627);
   U8051 : OR2_X1 port map( A1 => n20310, A2 => n7102, Z => n16004);
   U8052 : NAND2_X2 port map( A1 => n4079, A2 => n33724, ZN => n23684);
   U8053 : NAND2_X2 port map( A1 => n24292, A2 => n15520, ZN => n24011);
   U8054 : NAND2_X2 port map( A1 => n26529, A2 => n23685, ZN => n9219);
   U8058 : AOI21_X2 port map( A1 => n32104, A2 => n27094, B => n22335, ZN => 
                           n22999);
   U8060 : NOR2_X2 port map( A1 => n20378, A2 => n27887, ZN => n20323);
   U8062 : INV_X4 port map( I => n33817, ZN => n22876);
   U8068 : NAND2_X2 port map( A1 => n32105, A2 => n32090, ZN => n33817);
   U8071 : INV_X2 port map( I => n8601, ZN => n32105);
   U8072 : XOR2_X1 port map( A1 => n27289, A2 => n7129, Z => n9920);
   U8080 : INV_X2 port map( I => n32370, ZN => n27390);
   U8081 : XOR2_X1 port map( A1 => n5196, A2 => n31929, Z => n32370);
   U8082 : NOR2_X2 port map( A1 => n13903, A2 => n32107, ZN => n32462);
   U8087 : NOR3_X2 port map( A1 => n23749, A2 => n16781, A3 => n6661, ZN => 
                           n32107);
   U8094 : AOI22_X2 port map( A1 => n11022, A2 => n4993, B1 => n25896, B2 => 
                           n5387, ZN => n32132);
   U8099 : NOR2_X2 port map( A1 => n4993, A2 => n25870, ZN => n25896);
   U8100 : NAND2_X2 port map( A1 => n33044, A2 => n31946, ZN => n32859);
   U8102 : BUF_X2 port map( I => n32787, Z => n32108);
   U8105 : NAND2_X2 port map( A1 => n33321, A2 => n4131, ZN => n32255);
   U8108 : INV_X2 port map( I => n32109, ZN => n2229);
   U8109 : NOR2_X2 port map( A1 => n22557, A2 => n5379, ZN => n32496);
   U8114 : AOI22_X2 port map( A1 => n32110, A2 => n834, B1 => n1620, B2 => 
                           n12266, ZN => n25790);
   U8116 : NAND2_X2 port map( A1 => n12440, A2 => n25866, ZN => n32110);
   U8117 : XOR2_X1 port map( A1 => n14953, A2 => n14952, Z => n32124);
   U8118 : XOR2_X1 port map( A1 => n23469, A2 => n2854, Z => n9200);
   U8119 : NAND2_X2 port map( A1 => n30008, A2 => n7839, ZN => n2854);
   U8121 : NOR2_X2 port map( A1 => n927, A2 => n30813, ZN => n2370);
   U8122 : XOR2_X1 port map( A1 => n21023, A2 => n21025, Z => n6792);
   U8124 : XOR2_X1 port map( A1 => n13357, A2 => n5414, Z => n21023);
   U8125 : OAI22_X2 port map( A1 => n31964, A2 => n22487, B1 => n1289, B2 => 
                           n11629, ZN => n16884);
   U8127 : INV_X2 port map( I => n9617, ZN => n11629);
   U8129 : XOR2_X1 port map( A1 => n2144, A2 => n5353, Z => n9617);
   U8131 : XOR2_X1 port map( A1 => n2267, A2 => n28998, Z => n10657);
   U8135 : NAND3_X1 port map( A1 => n25793, A2 => n25792, A3 => n25791, ZN => 
                           n34070);
   U8136 : INV_X2 port map( I => n16486, ZN => n22865);
   U8137 : NOR3_X1 port map( A1 => n15382, A2 => n14905, A3 => n15476, ZN => 
                           n30771);
   U8139 : XOR2_X1 port map( A1 => n12972, A2 => n4992, Z => n5487);
   U8141 : NOR2_X2 port map( A1 => n1983, A2 => n5605, ZN => n4992);
   U8144 : XOR2_X1 port map( A1 => n4975, A2 => n12442, Z => n13908);
   U8147 : BUF_X2 port map( I => n29898, Z => n32111);
   U8148 : NOR2_X1 port map( A1 => n10987, A2 => n24326, ZN => n24329);
   U8149 : NAND2_X2 port map( A1 => n29811, A2 => n31090, ZN => n24326);
   U8150 : NAND2_X2 port map( A1 => n22353, A2 => n27638, ZN => n6750);
   U8154 : OAI22_X2 port map( A1 => n26410, A2 => n27390, B1 => n29142, B2 => 
                           n8919, ZN => n22353);
   U8155 : XOR2_X1 port map( A1 => n30301, A2 => n5762, Z => n24575);
   U8156 : NAND2_X1 port map( A1 => n10231, A2 => n20236, ZN => n13432);
   U8157 : XOR2_X1 port map( A1 => n24643, A2 => n24753, Z => n24419);
   U8159 : NAND2_X2 port map( A1 => n24078, A2 => n24077, ZN => n24643);
   U8162 : NAND2_X2 port map( A1 => n33133, A2 => n31878, ZN => n29898);
   U8163 : NOR3_X2 port map( A1 => n32115, A2 => n32112, A3 => n17849, ZN => 
                           n31571);
   U8164 : NOR3_X2 port map( A1 => n4183, A2 => n25462, A3 => n29116, ZN => 
                           n32112);
   U8165 : AOI21_X2 port map( A1 => n14722, A2 => n14087, B => n33352, ZN => 
                           n5906);
   U8166 : NAND2_X2 port map( A1 => n5820, A2 => n1106, ZN => n23028);
   U8167 : AOI22_X2 port map( A1 => n1232, A2 => n5079, B1 => n5080, B2 => 
                           n29985, ZN => n5284);
   U8170 : NAND2_X2 port map( A1 => n23981, A2 => n421, ZN => n5080);
   U8174 : XOR2_X1 port map( A1 => n6461, A2 => n14613, Z => n32914);
   U8177 : XOR2_X1 port map( A1 => n417, A2 => n32113, Z => n7072);
   U8179 : XOR2_X1 port map( A1 => n33840, A2 => n32114, Z => n32113);
   U8187 : XOR2_X1 port map( A1 => n22225, A2 => n34078, Z => n16897);
   U8190 : XOR2_X1 port map( A1 => n22190, A2 => n22191, Z => n11358);
   U8192 : XOR2_X1 port map( A1 => n7725, A2 => n21892, Z => n22190);
   U8197 : AOI21_X2 port map( A1 => n16001, A2 => n25753, B => n1082, ZN => 
                           n15709);
   U8198 : NAND2_X1 port map( A1 => n25707, A2 => n25705, ZN => n25753);
   U8201 : NAND3_X1 port map( A1 => n11186, A2 => n25905, A3 => n25901, ZN => 
                           n11185);
   U8207 : NAND2_X2 port map( A1 => n21378, A2 => n15751, ZN => n15728);
   U8209 : NAND2_X2 port map( A1 => n21362, A2 => n2230, ZN => n21378);
   U8210 : NOR2_X2 port map( A1 => n33735, A2 => n32116, ZN => n16987);
   U8211 : NOR2_X2 port map( A1 => n1351, A2 => n20447, ZN => n20405);
   U8213 : AOI21_X2 port map( A1 => n32723, A2 => n28982, B => n27373, ZN => 
                           n20447);
   U8214 : XOR2_X1 port map( A1 => n32117, A2 => n24740, Z => n7759);
   U8215 : XOR2_X1 port map( A1 => n33447, A2 => n705, Z => n32117);
   U8217 : XOR2_X1 port map( A1 => n33319, A2 => n32118, Z => n11622);
   U8219 : XOR2_X1 port map( A1 => n11782, A2 => n24803, Z => n32118);
   U8220 : INV_X4 port map( I => n16305, ZN => n32298);
   U8221 : AND2_X1 port map( A1 => n9390, A2 => n13969, Z => n5583);
   U8222 : XOR2_X1 port map( A1 => n21891, A2 => n7289, Z => n9193);
   U8224 : NAND2_X2 port map( A1 => n1678, A2 => n1677, ZN => n33117);
   U8226 : OAI21_X2 port map( A1 => n21465, A2 => n11729, B => n26728, ZN => 
                           n16888);
   U8229 : XOR2_X1 port map( A1 => n2956, A2 => n16520, Z => n210);
   U8234 : NAND3_X2 port map( A1 => n27759, A2 => n33372, A3 => n27760, ZN => 
                           n2956);
   U8238 : XOR2_X1 port map( A1 => n32120, A2 => n25783, Z => Ciphertext(165));
   U8239 : NAND3_X2 port map( A1 => n28989, A2 => n17222, A3 => n26948, ZN => 
                           n32120);
   U8241 : NAND2_X2 port map( A1 => n28073, A2 => n32121, ZN => n19314);
   U8244 : NAND2_X2 port map( A1 => n32150, A2 => n32122, ZN => n23928);
   U8248 : NAND3_X1 port map( A1 => n16186, A2 => n4892, A3 => n23920, ZN => 
                           n32122);
   U8256 : NAND2_X2 port map( A1 => n7146, A2 => n32123, ZN => n9159);
   U8259 : AOI22_X2 port map( A1 => n21320, A2 => n11187, B1 => n21324, B2 => 
                           n28017, ZN => n32123);
   U8260 : XOR2_X1 port map( A1 => n23358, A2 => n23253, Z => n23516);
   U8261 : NAND3_X2 port map( A1 => n22751, A2 => n22750, A3 => n22749, ZN => 
                           n23253);
   U8264 : NAND2_X2 port map( A1 => n32126, A2 => n32125, ZN => n26102);
   U8266 : INV_X2 port map( I => n12594, ZN => n32125);
   U8270 : XOR2_X1 port map( A1 => n13858, A2 => n7880, Z => n32469);
   U8272 : XOR2_X1 port map( A1 => n24545, A2 => n24544, Z => n7880);
   U8275 : BUF_X2 port map( I => n16559, Z => n32127);
   U8281 : NAND2_X2 port map( A1 => n57, A2 => n32128, ZN => n24254);
   U8283 : XOR2_X1 port map( A1 => n19768, A2 => n19703, Z => n19517);
   U8288 : AOI21_X2 port map( A1 => n5654, A2 => n18621, B => n31438, ZN => 
                           n19768);
   U8290 : NAND2_X2 port map( A1 => n10980, A2 => n32129, ZN => n21767);
   U8291 : OR2_X1 port map( A1 => n21051, A2 => n33684, Z => n32129);
   U8294 : OAI21_X2 port map( A1 => n6710, A2 => n6711, B => n6712, ZN => n6799
                           );
   U8295 : NOR2_X2 port map( A1 => n4207, A2 => n6877, ZN => n7078);
   U8296 : AOI21_X2 port map( A1 => n7151, A2 => n14995, B => n972, ZN => n4207
                           );
   U8297 : XOR2_X1 port map( A1 => n348, A2 => n32130, Z => n12805);
   U8299 : NAND2_X1 port map( A1 => n29981, A2 => n11507, ZN => n19984);
   U8300 : NOR2_X2 port map( A1 => n33720, A2 => n25784, ZN => n32874);
   U8301 : NOR3_X2 port map( A1 => n25757, A2 => n3275, A3 => n11899, ZN => 
                           n33720);
   U8302 : OR2_X1 port map( A1 => n8062, A2 => n4897, Z => n4873);
   U8304 : INV_X2 port map( I => n25106, ZN => n7334);
   U8305 : XOR2_X1 port map( A1 => n5601, A2 => n33338, Z => n8964);
   U8309 : XOR2_X1 port map( A1 => n32131, A2 => n32895, Z => n15731);
   U8310 : XOR2_X1 port map( A1 => n32243, A2 => n33265, Z => n32131);
   U8311 : OAI21_X2 port map( A1 => n19051, A2 => n19000, B => n27877, ZN => 
                           n19423);
   U8312 : AOI22_X2 port map( A1 => n18999, A2 => n19217, B1 => n19216, B2 => 
                           n31366, ZN => n27877);
   U8313 : XOR2_X1 port map( A1 => n23312, A2 => n23341, Z => n11039);
   U8314 : NAND2_X1 port map( A1 => n33235, A2 => n24866, ZN => n16850);
   U8315 : XOR2_X1 port map( A1 => n33161, A2 => n14065, Z => n24866);
   U8318 : NOR2_X1 port map( A1 => n25002, A2 => n3232, ZN => n14609);
   U8319 : OAI21_X2 port map( A1 => n15061, A2 => n15062, B => n15059, ZN => 
                           n25002);
   U8320 : XOR2_X1 port map( A1 => n10631, A2 => n3935, Z => n32417);
   U8322 : NOR2_X2 port map( A1 => n14502, A2 => n4959, ZN => n10631);
   U8324 : INV_X4 port map( I => n14001, ZN => n24925);
   U8325 : NAND2_X2 port map( A1 => n8776, A2 => n8777, ZN => n14001);
   U8330 : AOI22_X2 port map( A1 => n23912, A2 => n7005, B1 => n23910, B2 => 
                           n23588, ZN => n33808);
   U8333 : INV_X2 port map( I => n16226, ZN => n21078);
   U8335 : XOR2_X1 port map( A1 => n26954, A2 => n13403, Z => n16226);
   U8336 : NAND2_X2 port map( A1 => n11020, A2 => n32132, ZN => n13960);
   U8346 : XOR2_X1 port map( A1 => n24513, A2 => n30323, Z => n24788);
   U8349 : NAND3_X2 port map( A1 => n4393, A2 => n17493, A3 => n17492, ZN => 
                           n24513);
   U8351 : NOR2_X2 port map( A1 => n12662, A2 => n34127, ZN => n33306);
   U8352 : NAND2_X2 port map( A1 => n7034, A2 => n32133, ZN => n8238);
   U8354 : AOI22_X2 port map( A1 => n7885, A2 => n33589, B1 => n23650, B2 => 
                           n28671, ZN => n32133);
   U8356 : NAND2_X2 port map( A1 => n22399, A2 => n17930, ZN => n23046);
   U8357 : NAND2_X2 port map( A1 => n21980, A2 => n21981, ZN => n22399);
   U8358 : XOR2_X1 port map( A1 => n32134, A2 => n19492, Z => n706);
   U8359 : XOR2_X1 port map( A1 => n27895, A2 => n19577, Z => n32134);
   U8361 : OAI21_X2 port map( A1 => n32135, A2 => n17762, B => n8307, ZN => 
                           n32731);
   U8363 : XOR2_X1 port map( A1 => n32136, A2 => n1431, Z => Ciphertext(163));
   U8366 : NOR3_X1 port map( A1 => n28854, A2 => n14615, A3 => n12395, ZN => 
                           n32136);
   U8369 : XOR2_X1 port map( A1 => n6466, A2 => n32137, Z => n7);
   U8371 : XOR2_X1 port map( A1 => n21893, A2 => n32072, Z => n32137);
   U8372 : NOR2_X2 port map( A1 => n30473, A2 => n24025, ZN => n24936);
   U8374 : OAI22_X2 port map( A1 => n13326, A2 => n14268, B1 => n14042, B2 => 
                           n1221, ZN => n30473);
   U8375 : NAND2_X2 port map( A1 => n32139, A2 => n32138, ZN => n28539);
   U8378 : NOR2_X1 port map( A1 => n31992, A2 => n13160, ZN => n32139);
   U8381 : XOR2_X1 port map( A1 => n32140, A2 => n24407, Z => n17074);
   U8387 : XOR2_X1 port map( A1 => n12422, A2 => n12512, Z => n32140);
   U8388 : BUF_X2 port map( I => n1169, Z => n32141);
   U8389 : NAND2_X2 port map( A1 => n32142, A2 => n9085, ZN => n5973);
   U8394 : NAND3_X2 port map( A1 => n32048, A2 => n22953, A3 => n7544, ZN => 
                           n32142);
   U8395 : XOR2_X1 port map( A1 => n20789, A2 => n20787, Z => n31070);
   U8403 : XOR2_X1 port map( A1 => n10235, A2 => n1507, Z => n28747);
   U8405 : XOR2_X1 port map( A1 => n24842, A2 => n12720, Z => n1507);
   U8406 : NAND2_X1 port map( A1 => n18352, A2 => n9264, ZN => n32769);
   U8409 : AOI22_X2 port map( A1 => n16866, A2 => n22477, B1 => n27207, B2 => 
                           n18098, ZN => n32482);
   U8412 : NAND3_X2 port map( A1 => n3708, A2 => n8799, A3 => n32145, ZN => 
                           n11754);
   U8415 : AOI22_X2 port map( A1 => n4319, A2 => n17694, B1 => n29080, B2 => 
                           n30980, ZN => n32145);
   U8420 : INV_X1 port map( I => n31185, ZN => n20777);
   U8423 : NAND2_X2 port map( A1 => n32288, A2 => n32146, ZN => n1560);
   U8425 : NAND3_X2 port map( A1 => n12429, A2 => n12430, A3 => n32936, ZN => 
                           n32146);
   U8426 : XOR2_X1 port map( A1 => n15517, A2 => n32870, Z => n24746);
   U8435 : NAND2_X2 port map( A1 => n15988, A2 => n13658, ZN => n15517);
   U8437 : NAND2_X1 port map( A1 => n2643, A2 => n14681, ZN => n21469);
   U8438 : NAND2_X2 port map( A1 => n8740, A2 => n21153, ZN => n2643);
   U8439 : NOR2_X1 port map( A1 => n25587, A2 => n25586, ZN => n33500);
   U8441 : OAI21_X1 port map( A1 => n13066, A2 => n9003, B => n9954, ZN => 
                           n30838);
   U8443 : XOR2_X1 port map( A1 => n20861, A2 => n17423, Z => n10169);
   U8445 : NAND2_X2 port map( A1 => n14567, A2 => n14565, ZN => n20861);
   U8448 : NOR2_X1 port map( A1 => n32148, A2 => n861, ZN => n29843);
   U8451 : NOR2_X2 port map( A1 => n32149, A2 => n13212, ZN => n6569);
   U8454 : NAND2_X1 port map( A1 => n32151, A2 => n8760, ZN => n32150);
   U8461 : NOR2_X1 port map( A1 => n23920, A2 => n13361, ZN => n32151);
   U8462 : XOR2_X1 port map( A1 => n32733, A2 => n19679, Z => n8637);
   U8466 : XOR2_X1 port map( A1 => n30547, A2 => n32152, Z => n23916);
   U8473 : XOR2_X1 port map( A1 => n23334, A2 => n14527, Z => n32152);
   U8478 : XOR2_X1 port map( A1 => n20713, A2 => n32153, Z => n21071);
   U8479 : XOR2_X1 port map( A1 => n21020, A2 => n12618, Z => n32153);
   U8481 : NOR2_X2 port map( A1 => n8247, A2 => n8246, ZN => n8245);
   U8483 : AOI22_X2 port map( A1 => n6559, A2 => n20300, B1 => n20358, B2 => 
                           n16011, ZN => n17177);
   U8484 : NOR2_X2 port map( A1 => n20238, A2 => n11453, ZN => n16011);
   U8485 : NOR2_X1 port map( A1 => n33512, A2 => n16304, ZN => n16410);
   U8488 : XOR2_X1 port map( A1 => n32155, A2 => n32156, Z => n33534);
   U8490 : XOR2_X1 port map( A1 => n26462, A2 => n21944, Z => n32156);
   U8493 : XOR2_X1 port map( A1 => n32157, A2 => n25541, Z => Ciphertext(120));
   U8499 : NAND4_X2 port map( A1 => n8805, A2 => n30134, A3 => n8804, A4 => 
                           n25555, ZN => n32157);
   U8500 : NOR2_X1 port map( A1 => n12302, A2 => n27925, ZN => n32566);
   U8501 : AOI22_X2 port map( A1 => n12482, A2 => n17005, B1 => n9294, B2 => 
                           n27990, ZN => n16380);
   U8502 : OAI22_X2 port map( A1 => n9294, A2 => n28591, B1 => n25199, B2 => 
                           n32873, ZN => n12482);
   U8507 : INV_X2 port map( I => n23405, ZN => n33476);
   U8509 : NAND2_X2 port map( A1 => n30982, A2 => n16879, ZN => n23405);
   U8511 : XOR2_X1 port map( A1 => n19390, A2 => n19568, Z => n2951);
   U8512 : XOR2_X1 port map( A1 => n19629, A2 => n19389, Z => n19568);
   U8513 : NAND3_X2 port map( A1 => n20444, A2 => n30496, A3 => n20633, ZN => 
                           n4469);
   U8514 : NAND2_X2 port map( A1 => n30594, A2 => n15162, ZN => n20444);
   U8515 : NOR2_X1 port map( A1 => n31448, A2 => n19936, ZN => n14905);
   U8518 : INV_X2 port map( I => n32158, ZN => n11933);
   U8520 : XNOR2_X1 port map( A1 => n284, A2 => n10051, ZN => n32158);
   U8521 : NAND2_X2 port map( A1 => n12214, A2 => n32159, ZN => n16807);
   U8522 : NAND2_X2 port map( A1 => n18324, A2 => n18567, ZN => n32159);
   U8534 : INV_X2 port map( I => n29261, ZN => n22477);
   U8535 : XOR2_X1 port map( A1 => n32160, A2 => n24689, Z => n24407);
   U8538 : XOR2_X1 port map( A1 => n24785, A2 => n30327, Z => n32160);
   U8541 : NAND2_X2 port map( A1 => n17249, A2 => n32161, ZN => n1266);
   U8544 : NAND3_X2 port map( A1 => n17247, A2 => n17248, A3 => n9620, ZN => 
                           n32161);
   U8547 : XOR2_X1 port map( A1 => n15560, A2 => n22061, Z => n14181);
   U8548 : NAND2_X2 port map( A1 => n26102, A2 => n2777, ZN => n15560);
   U8549 : XOR2_X1 port map( A1 => n27175, A2 => n25783, Z => n102);
   U8551 : NOR3_X2 port map( A1 => n17740, A2 => n12445, A3 => n12444, ZN => 
                           n27175);
   U8552 : NOR2_X2 port map( A1 => n13319, A2 => n13255, ZN => n21381);
   U8560 : AND2_X1 port map( A1 => n17948, A2 => n15212, Z => n29280);
   U8561 : XOR2_X1 port map( A1 => n32162, A2 => n32467, Z => n30492);
   U8564 : NAND2_X2 port map( A1 => n3424, A2 => n30079, ZN => n32467);
   U8565 : INV_X2 port map( I => n11665, ZN => n32162);
   U8567 : XOR2_X1 port map( A1 => n8070, A2 => n8069, Z => n23587);
   U8568 : NOR2_X2 port map( A1 => n23860, A2 => n23556, ZN => n26955);
   U8569 : NAND2_X2 port map( A1 => n28273, A2 => n17661, ZN => n23556);
   U8572 : NAND2_X2 port map( A1 => n18991, A2 => n18992, ZN => n19400);
   U8573 : NOR2_X2 port map( A1 => n13678, A2 => n33583, ZN => n26628);
   U8575 : NAND2_X2 port map( A1 => n206, A2 => n17375, ZN => n30033);
   U8577 : NAND2_X2 port map( A1 => n10939, A2 => n8268, ZN => n20200);
   U8580 : NAND2_X2 port map( A1 => n2495, A2 => n33003, ZN => n10939);
   U8581 : NAND2_X2 port map( A1 => n32163, A2 => n32289, ZN => n31171);
   U8586 : NAND2_X1 port map( A1 => n12208, A2 => n16305, ZN => n32163);
   U8592 : INV_X2 port map( I => n26898, ZN => n23034);
   U8594 : NAND3_X2 port map( A1 => n33901, A2 => n1516, A3 => n30989, ZN => 
                           n26898);
   U8596 : NAND2_X2 port map( A1 => n22474, A2 => n29261, ZN => n13185);
   U8599 : OAI21_X2 port map( A1 => n8230, A2 => n32164, B => n34104, ZN => 
                           n26261);
   U8600 : NAND2_X1 port map( A1 => n6483, A2 => n21580, ZN => n32164);
   U8601 : NAND3_X1 port map( A1 => n4086, A2 => n33097, A3 => n23628, ZN => 
                           n33135);
   U8604 : BUF_X4 port map( I => n28374, Z => n32323);
   U8605 : XOR2_X1 port map( A1 => n4672, A2 => n32165, Z => n5361);
   U8611 : XOR2_X1 port map( A1 => n4671, A2 => n4771, Z => n32165);
   U8628 : XOR2_X1 port map( A1 => Plaintext(20), A2 => Key(20), Z => n18655);
   U8630 : AOI22_X2 port map( A1 => n4774, A2 => n11041, B1 => n12982, B2 => 
                           n24309, ZN => n24199);
   U8636 : OAI22_X2 port map( A1 => n4099, A2 => n6723, B1 => n31982, B2 => 
                           n18204, ZN => n24309);
   U8637 : NOR3_X2 port map( A1 => n33455, A2 => n9335, A3 => n5743, ZN => 
                           n32636);
   U8640 : AOI21_X2 port map( A1 => n32166, A2 => n2993, B => n26545, ZN => 
                           n2158);
   U8642 : XOR2_X1 port map( A1 => n17519, A2 => n22275, Z => n15618);
   U8645 : XOR2_X1 port map( A1 => n14125, A2 => n7808, Z => n17519);
   U8650 : NAND2_X1 port map( A1 => n29614, A2 => n14418, ZN => n32430);
   U8651 : NAND2_X1 port map( A1 => n18133, A2 => n32309, ZN => n23715);
   U8652 : XOR2_X1 port map( A1 => n31237, A2 => n23537, Z => n32309);
   U8655 : XOR2_X1 port map( A1 => n20905, A2 => n27174, Z => n20989);
   U8658 : NAND2_X2 port map( A1 => n5951, A2 => n5949, ZN => n20905);
   U8666 : XOR2_X1 port map( A1 => n32167, A2 => n16775, Z => n28179);
   U8667 : XOR2_X1 port map( A1 => n27729, A2 => n20824, Z => n32167);
   U8668 : XOR2_X1 port map( A1 => n9207, A2 => n27693, Z => n26317);
   U8670 : NOR2_X2 port map( A1 => n29547, A2 => n32168, ZN => n29523);
   U8672 : XOR2_X1 port map( A1 => n26701, A2 => n23186, Z => n23246);
   U8675 : NAND3_X2 port map( A1 => n33777, A2 => n13365, A3 => n14516, ZN => 
                           n26701);
   U8677 : INV_X2 port map( I => n21628, ZN => n21772);
   U8679 : AOI22_X2 port map( A1 => n31524, A2 => n23669, B1 => n23953, B2 => 
                           n33788, ZN => n9995);
   U8680 : NAND2_X2 port map( A1 => n12986, A2 => n32169, ZN => n26585);
   U8682 : OAI21_X2 port map( A1 => n19801, A2 => n19800, B => n19867, ZN => 
                           n32169);
   U8688 : XOR2_X1 port map( A1 => n11218, A2 => n19529, Z => n4578);
   U8696 : XOR2_X1 port map( A1 => n30943, A2 => n19708, Z => n19529);
   U8700 : XOR2_X1 port map( A1 => n21014, A2 => n20718, Z => n32379);
   U8713 : XOR2_X1 port map( A1 => n2789, A2 => n2198, Z => n20718);
   U8714 : OAI21_X1 port map( A1 => n8334, A2 => n22962, B => n22815, ZN => 
                           n33049);
   U8716 : BUF_X2 port map( I => n15917, Z => n32170);
   U8719 : XOR2_X1 port map( A1 => n32171, A2 => n13863, Z => n15205);
   U8723 : XOR2_X1 port map( A1 => n32367, A2 => n27240, Z => n32171);
   U8725 : BUF_X2 port map( I => n32081, Z => n32172);
   U8733 : OAI21_X2 port map( A1 => n30617, A2 => n19761, B => n32173, ZN => 
                           n20312);
   U8734 : AOI22_X2 port map( A1 => n19759, A2 => n20045, B1 => n31715, B2 => 
                           n31823, ZN => n32173);
   U8736 : NAND3_X2 port map( A1 => n29668, A2 => n20414, A3 => n19908, ZN => 
                           n29667);
   U8741 : XOR2_X1 port map( A1 => n19626, A2 => n19624, Z => n17541);
   U8746 : OAI22_X2 port map( A1 => n12271, A2 => n12268, B1 => n7968, B2 => 
                           n18752, ZN => n19626);
   U8749 : NAND2_X2 port map( A1 => n33767, A2 => n32174, ZN => n5211);
   U8750 : AOI22_X2 port map( A1 => n32234, A2 => n32233, B1 => n5821, B2 => 
                           n16976, ZN => n32174);
   U8752 : NAND2_X2 port map( A1 => n31030, A2 => n1333, ZN => n21411);
   U8753 : XOR2_X1 port map( A1 => n14000, A2 => n5539, Z => n24569);
   U8754 : NAND2_X2 port map( A1 => n31039, A2 => n32836, ZN => n5539);
   U8756 : NAND2_X2 port map( A1 => n29502, A2 => n32175, ZN => n11608);
   U8757 : NAND3_X1 port map( A1 => n32917, A2 => n6003, A3 => n23970, ZN => 
                           n32175);
   U8758 : NOR2_X2 port map( A1 => n31979, A2 => n25843, ZN => n25855);
   U8763 : OAI22_X2 port map( A1 => n33196, A2 => n25887, B1 => n7350, B2 => 
                           n25866, ZN => n25843);
   U8770 : OAI22_X2 port map( A1 => n6553, A2 => n896, B1 => n23045, B2 => 
                           n23042, ZN => n13341);
   U8778 : XOR2_X1 port map( A1 => n18365, A2 => Key(49), Z => n32787);
   U8782 : OR2_X1 port map( A1 => n8422, A2 => n9549, Z => n10966);
   U8791 : OAI21_X2 port map( A1 => n31925, A2 => n17039, B => n15444, ZN => 
                           n15443);
   U8795 : NOR2_X1 port map( A1 => n10599, A2 => n10787, ZN => n17039);
   U8798 : XOR2_X1 port map( A1 => n6913, A2 => n19706, Z => n32213);
   U8803 : XOR2_X1 port map( A1 => n2920, A2 => n1944, Z => n19706);
   U8804 : XOR2_X1 port map( A1 => n7674, A2 => n7628, Z => n5321);
   U8807 : XOR2_X1 port map( A1 => n21040, A2 => n33814, Z => n7674);
   U8809 : AOI21_X2 port map( A1 => n11688, A2 => n1377, B => n19309, ZN => 
                           n19311);
   U8811 : XOR2_X1 port map( A1 => n12738, A2 => n27673, Z => n33354);
   U8816 : XOR2_X1 port map( A1 => n20755, A2 => n21016, Z => n20722);
   U8819 : NOR2_X2 port map( A1 => n1929, A2 => n1930, ZN => n21016);
   U8824 : NAND2_X2 port map( A1 => n1472, A2 => n30935, ZN => n32177);
   U8825 : XOR2_X1 port map( A1 => n6373, A2 => n24991, Z => n7211);
   U8829 : NAND2_X2 port map( A1 => n30202, A2 => n33791, ZN => n6373);
   U8835 : NOR2_X2 port map( A1 => n14178, A2 => n19153, ZN => n17528);
   U8837 : XOR2_X1 port map( A1 => n1607, A2 => n28239, Z => n17485);
   U8838 : XOR2_X1 port map( A1 => n19517, A2 => n19518, Z => n1615);
   U8855 : XOR2_X1 port map( A1 => n5775, A2 => n14662, Z => n8556);
   U8858 : XOR2_X1 port map( A1 => n20803, A2 => n32894, Z => n14662);
   U8871 : BUF_X2 port map( I => n26158, Z => n32178);
   U8879 : XOR2_X1 port map( A1 => n32179, A2 => n380, Z => n33903);
   U8882 : XOR2_X1 port map( A1 => n10649, A2 => n12627, Z => n32179);
   U8886 : XOR2_X1 port map( A1 => n20710, A2 => n14522, Z => n26769);
   U8887 : XOR2_X1 port map( A1 => n32180, A2 => n1196, Z => Ciphertext(24));
   U8888 : NOR2_X1 port map( A1 => n32244, A2 => n24989, ZN => n32180);
   U8895 : XOR2_X1 port map( A1 => n15035, A2 => n15036, Z => n15734);
   U8896 : INV_X2 port map( I => n32181, ZN => n499);
   U8897 : XNOR2_X1 port map( A1 => n31411, A2 => n10219, ZN => n32181);
   U8908 : NAND2_X1 port map( A1 => n4525, A2 => n24995, ZN => n315);
   U8916 : NOR2_X1 port map( A1 => n29361, A2 => n21373, ZN => n8856);
   U8917 : XOR2_X1 port map( A1 => n12720, A2 => n17912, Z => n24749);
   U8922 : NAND2_X2 port map( A1 => n16410, A2 => n16409, ZN => n17912);
   U8923 : NOR2_X2 port map( A1 => n32183, A2 => n32182, ZN => n8091);
   U8925 : INV_X2 port map( I => n100, ZN => n32183);
   U8926 : XOR2_X1 port map( A1 => n22063, A2 => n16696, Z => n22064);
   U8929 : NAND2_X2 port map( A1 => n32204, A2 => n9961, ZN => n22063);
   U8932 : XOR2_X1 port map( A1 => n3030, A2 => n27767, Z => n27601);
   U8933 : AND2_X1 port map( A1 => n23082, A2 => n22962, Z => n33294);
   U8936 : XOR2_X1 port map( A1 => n5146, A2 => n139, Z => n2345);
   U8948 : OAI22_X1 port map( A1 => n22697, A2 => n33675, B1 => n22816, B2 => 
                           n27419, ZN => n16463);
   U8955 : XOR2_X1 port map( A1 => n23299, A2 => n12475, Z => n12474);
   U8957 : XOR2_X1 port map( A1 => n27174, A2 => n15877, Z => n20778);
   U8967 : NAND2_X2 port map( A1 => n32385, A2 => n20568, ZN => n27174);
   U8971 : NAND2_X2 port map( A1 => n14184, A2 => n14724, ZN => n24837);
   U8974 : AOI22_X2 port map( A1 => n31228, A2 => n33891, B1 => n3039, B2 => 
                           n3038, ZN => n14184);
   U8975 : AOI21_X2 port map( A1 => n32323, A2 => n33680, B => n30230, ZN => 
                           n26976);
   U8977 : NAND2_X1 port map( A1 => n32976, A2 => n3220, ZN => n1504);
   U8981 : OAI21_X2 port map( A1 => n32185, A2 => n16367, B => n16366, ZN => 
                           n31282);
   U8985 : AOI22_X2 port map( A1 => n239, A2 => n22557, B1 => n22343, B2 => 
                           n7090, ZN => n32185);
   U8986 : AND2_X1 port map( A1 => n33224, A2 => n2957, Z => n12343);
   U8988 : AND2_X1 port map( A1 => n18184, A2 => n32040, Z => n17734);
   U9005 : NAND3_X2 port map( A1 => n17415, A2 => n21345, A3 => n15422, ZN => 
                           n18184);
   U9007 : AOI21_X2 port map( A1 => n820, A2 => n33714, B => n16568, ZN => 
                           n4442);
   U9010 : INV_X1 port map( I => n13913, ZN => n32952);
   U9022 : XNOR2_X1 port map( A1 => n31477, A2 => n20754, ZN => n31185);
   U9023 : XOR2_X1 port map( A1 => n33369, A2 => n26140, Z => n27736);
   U9024 : NAND2_X1 port map( A1 => n23111, A2 => n3103, ZN => n30476);
   U9025 : NAND2_X2 port map( A1 => n29598, A2 => n32518, ZN => n3103);
   U9026 : XOR2_X1 port map( A1 => n13178, A2 => n8160, Z => n13177);
   U9028 : NAND3_X2 port map( A1 => n31998, A2 => n28880, A3 => n19874, ZN => 
                           n27879);
   U9031 : OAI21_X2 port map( A1 => n13950, A2 => n11503, B => n24286, ZN => 
                           n33184);
   U9033 : INV_X2 port map( I => n9624, ZN => n11503);
   U9034 : NAND3_X2 port map( A1 => n32, A2 => n25954, A3 => n6467, ZN => n9624
                           );
   U9036 : XOR2_X1 port map( A1 => n20784, A2 => n20990, Z => n20886);
   U9041 : NOR2_X2 port map( A1 => n12479, A2 => n7033, ZN => n20784);
   U9044 : OAI21_X2 port map( A1 => n28406, A2 => n17985, B => n32187, ZN => 
                           n3313);
   U9045 : NAND2_X2 port map( A1 => n28400, A2 => n17985, ZN => n32187);
   U9053 : OAI21_X2 port map( A1 => n9184, A2 => n32188, B => n23043, ZN => 
                           n23049);
   U9056 : NOR2_X2 port map( A1 => n33007, A2 => n23042, ZN => n32188);
   U9059 : XOR2_X1 port map( A1 => n31769, A2 => n32189, Z => n9626);
   U9060 : XOR2_X1 port map( A1 => n28981, A2 => n10122, Z => n32189);
   U9062 : XOR2_X1 port map( A1 => n30482, A2 => n11326, Z => n5509);
   U9065 : XOR2_X1 port map( A1 => n32190, A2 => n25074, Z => Ciphertext(44));
   U9068 : INV_X2 port map( I => n22689, ZN => n32194);
   U9070 : XOR2_X1 port map( A1 => n9347, A2 => n32195, Z => n29471);
   U9072 : XOR2_X1 port map( A1 => n32715, A2 => n23384, Z => n32195);
   U9074 : XOR2_X1 port map( A1 => n33929, A2 => n32196, Z => n29631);
   U9076 : XOR2_X1 port map( A1 => n12659, A2 => n34112, Z => n32196);
   U9077 : NAND2_X2 port map( A1 => n25980, A2 => n397, ZN => n10286);
   U9078 : NAND2_X2 port map( A1 => n13139, A2 => n32198, ZN => n12374);
   U9080 : AOI22_X2 port map( A1 => n33870, A2 => n975, B1 => n23778, B2 => 
                           n6992, ZN => n32198);
   U9081 : NAND2_X2 port map( A1 => n6503, A2 => n32199, ZN => n11897);
   U9082 : AOI21_X1 port map( A1 => n22901, A2 => n852, B => n26507, ZN => 
                           n32199);
   U9088 : INV_X2 port map( I => n32200, ZN => n27799);
   U9089 : XOR2_X1 port map( A1 => n22518, A2 => n22517, Z => n32200);
   U9095 : XOR2_X1 port map( A1 => n7057, A2 => n11219, Z => n11218);
   U9097 : NAND2_X2 port map( A1 => n11178, A2 => n11177, ZN => n7057);
   U9098 : XOR2_X1 port map( A1 => n30041, A2 => n1417, Z => n27349);
   U9099 : NAND2_X2 port map( A1 => n30182, A2 => n29060, ZN => n30041);
   U9107 : NAND2_X2 port map( A1 => n31983, A2 => n6490, ZN => n14058);
   U9108 : XOR2_X1 port map( A1 => n13843, A2 => n19619, Z => n13842);
   U9109 : NAND2_X2 port map( A1 => n28821, A2 => n21437, ZN => n6544);
   U9110 : NAND2_X2 port map( A1 => n19961, A2 => n27491, ZN => n19962);
   U9111 : XOR2_X1 port map( A1 => n188, A2 => n32703, Z => n11974);
   U9114 : XOR2_X1 port map( A1 => n32124, A2 => n12614, Z => n2900);
   U9120 : INV_X2 port map( I => n32202, ZN => n8422);
   U9121 : XOR2_X1 port map( A1 => Plaintext(61), A2 => Key(61), Z => n32202);
   U9122 : XOR2_X1 port map( A1 => n24469, A2 => n14762, Z => n29809);
   U9123 : XOR2_X1 port map( A1 => n2117, A2 => n24545, Z => n24469);
   U9130 : NAND2_X2 port map( A1 => n13340, A2 => n22758, ZN => n31499);
   U9131 : OAI22_X1 port map( A1 => n9792, A2 => n31231, B1 => n2202, B2 => 
                           n9793, ZN => n32204);
   U9133 : XOR2_X1 port map( A1 => n20906, A2 => n21003, Z => n8026);
   U9135 : XOR2_X1 port map( A1 => n20970, A2 => n21037, Z => n20906);
   U9140 : AOI21_X1 port map( A1 => n22999, A2 => n9280, B => n32635, ZN => 
                           n33640);
   U9141 : INV_X1 port map( I => n18269, ZN => n33613);
   U9146 : NAND2_X2 port map( A1 => n32637, A2 => n32205, ZN => n7831);
   U9147 : XOR2_X1 port map( A1 => n15978, A2 => n32206, Z => n28978);
   U9149 : NOR2_X2 port map( A1 => n27353, A2 => n6188, ZN => n15978);
   U9151 : NAND2_X2 port map( A1 => n11023, A2 => n32207, ZN => n10943);
   U9152 : NOR2_X2 port map( A1 => n448, A2 => n30560, ZN => n32207);
   U9155 : NAND2_X2 port map( A1 => n33551, A2 => n12913, ZN => n32300);
   U9158 : NAND3_X2 port map( A1 => n30587, A2 => n17884, A3 => n17883, ZN => 
                           n32974);
   U9170 : INV_X2 port map( I => n23841, ZN => n32209);
   U9171 : XOR2_X1 port map( A1 => n3736, A2 => n32211, Z => n28605);
   U9173 : XOR2_X1 port map( A1 => n3735, A2 => n12618, Z => n32211);
   U9176 : AOI22_X2 port map( A1 => n32494, A2 => n32212, B1 => n6235, B2 => 
                           n10993, ZN => n24147);
   U9177 : NAND2_X2 port map( A1 => n13031, A2 => n23681, ZN => n32212);
   U9181 : NAND2_X2 port map( A1 => n14752, A2 => n10099, ZN => n24908);
   U9187 : NAND2_X2 port map( A1 => n6471, A2 => n18209, ZN => n14957);
   U9188 : NAND2_X2 port map( A1 => n31995, A2 => n21087, ZN => n18209);
   U9189 : NAND2_X2 port map( A1 => n21688, A2 => n12561, ZN => n21551);
   U9190 : XOR2_X1 port map( A1 => n11332, A2 => n3935, Z => n10235);
   U9194 : NAND3_X2 port map( A1 => n33689, A2 => n29584, A3 => n11331, ZN => 
                           n11332);
   U9196 : NAND3_X2 port map( A1 => n25853, A2 => n15546, A3 => n16673, ZN => 
                           n30071);
   U9211 : NAND2_X2 port map( A1 => n25834, A2 => n14199, ZN => n25853);
   U9212 : XOR2_X1 port map( A1 => n10582, A2 => n32511, Z => n10679);
   U9213 : AOI21_X2 port map( A1 => n22540, A2 => n22539, B => n32448, ZN => 
                           n32447);
   U9214 : NAND2_X2 port map( A1 => n17147, A2 => n22427, ZN => n22539);
   U9218 : NAND2_X2 port map( A1 => n698, A2 => n29127, ZN => n32443);
   U9221 : XOR2_X1 port map( A1 => n6914, A2 => n32213, Z => n15356);
   U9223 : INV_X2 port map( I => n2841, ZN => n14841);
   U9224 : XOR2_X1 port map( A1 => n23335, A2 => n32214, Z => n2841);
   U9225 : INV_X1 port map( I => n6190, ZN => n32820);
   U9228 : NAND2_X2 port map( A1 => n14550, A2 => n14548, ZN => n16554);
   U9229 : NAND2_X2 port map( A1 => n12858, A2 => n27369, ZN => n14550);
   U9233 : NOR2_X2 port map( A1 => n31485, A2 => n32215, ZN => n16280);
   U9237 : NOR2_X2 port map( A1 => n30448, A2 => n33594, ZN => n32216);
   U9240 : OAI21_X1 port map( A1 => n10724, A2 => n22644, B => n1292, ZN => 
                           n32217);
   U9251 : XOR2_X1 port map( A1 => n32220, A2 => n30049, Z => n33487);
   U9253 : XOR2_X1 port map( A1 => n32809, A2 => n32022, Z => n32220);
   U9254 : NAND2_X1 port map( A1 => n22789, A2 => n33388, ZN => n33387);
   U9258 : XOR2_X1 port map( A1 => n23341, A2 => n4564, Z => n4563);
   U9261 : OAI22_X1 port map( A1 => n32221, A2 => n5900, B1 => n5903, B2 => 
                           n17838, ZN => n32235);
   U9268 : NOR2_X1 port map( A1 => n24994, A2 => n7831, ZN => n32221);
   U9269 : XOR2_X1 port map( A1 => n22243, A2 => n22306, Z => n21998);
   U9273 : NAND2_X2 port map( A1 => n16163, A2 => n16164, ZN => n22243);
   U9275 : XOR2_X1 port map( A1 => n5767, A2 => n7605, Z => n12871);
   U9277 : NAND2_X1 port map( A1 => n32819, A2 => n12848, ZN => n23170);
   U9282 : INV_X1 port map( I => n15324, ZN => n32510);
   U9283 : XOR2_X1 port map( A1 => n12659, A2 => n32222, Z => n33662);
   U9284 : XOR2_X1 port map( A1 => n2564, A2 => n14613, Z => n32222);
   U9285 : INV_X2 port map( I => n16554, ZN => n1086);
   U9286 : INV_X2 port map( I => n32550, ZN => n32223);
   U9288 : NOR2_X2 port map( A1 => n32957, A2 => n11513, ZN => n32550);
   U9299 : NAND2_X2 port map( A1 => n12900, A2 => n18026, ZN => n31407);
   U9304 : NAND3_X1 port map( A1 => n25296, A2 => n25344, A3 => n25397, ZN => 
                           n18026);
   U9306 : NOR2_X2 port map( A1 => n24200, A2 => n26027, ZN => n28505);
   U9309 : AOI22_X2 port map( A1 => n738, A2 => n24158, B1 => n7503, B2 => 
                           n24008, ZN => n24200);
   U9313 : OAI21_X1 port map( A1 => n14609, A2 => n25005, B => n42, ZN => 
                           n32227);
   U9316 : NAND3_X1 port map( A1 => n32227, A2 => n14607, A3 => n25004, ZN => 
                           n30063);
   U9317 : NAND3_X2 port map( A1 => n30922, A2 => n30923, A3 => n6999, ZN => 
                           n6997);
   U9318 : NAND2_X2 port map( A1 => n7722, A2 => n32224, ZN => n16954);
   U9320 : AOI22_X2 port map( A1 => n21057, A2 => n11745, B1 => n7721, B2 => 
                           n28406, ZN => n32224);
   U9321 : INV_X2 port map( I => n13970, ZN => n28953);
   U9324 : OAI22_X2 port map( A1 => n7157, A2 => n7154, B1 => n7291, B2 => 
                           n20604, ZN => n13970);
   U9329 : NAND2_X1 port map( A1 => n32225, A2 => n17383, ZN => n16284);
   U9334 : NAND3_X1 port map( A1 => n17089, A2 => n16661, A3 => n16660, ZN => 
                           n32225);
   U9337 : NAND2_X2 port map( A1 => n2529, A2 => n32226, ZN => n8968);
   U9342 : NAND2_X2 port map( A1 => n24289, A2 => n24110, ZN => n32226);
   U9344 : XOR2_X1 port map( A1 => n8761, A2 => n23330, Z => n26279);
   U9345 : XOR2_X1 port map( A1 => n23233, A2 => n23299, Z => n8761);
   U9346 : XOR2_X1 port map( A1 => n23454, A2 => n23474, Z => n23324);
   U9356 : NOR2_X2 port map( A1 => n17585, A2 => n12790, ZN => n23454);
   U9368 : NAND2_X2 port map( A1 => n10784, A2 => n10785, ZN => n32253);
   U9369 : NAND2_X2 port map( A1 => n816, A2 => n17237, ZN => n9986);
   U9370 : NAND3_X2 port map( A1 => n31805, A2 => n8589, A3 => n8592, ZN => 
                           n17237);
   U9372 : CLKBUF_X4 port map( I => n14855, Z => n4728);
   U9379 : AOI22_X2 port map( A1 => n11317, A2 => n8365, B1 => n33563, B2 => 
                           n10296, ZN => n32826);
   U9384 : XOR2_X1 port map( A1 => n4680, A2 => n20835, Z => n20993);
   U9388 : NOR2_X2 port map( A1 => n4534, A2 => n4535, ZN => n4680);
   U9390 : NOR2_X2 port map( A1 => n33972, A2 => n21188, ZN => n4494);
   U9391 : INV_X2 port map( I => n32229, ZN => n32228);
   U9393 : OAI21_X2 port map( A1 => n26120, A2 => n6713, B => n27168, ZN => 
                           n32229);
   U9395 : NOR2_X2 port map( A1 => n4956, A2 => n28403, ZN => n3935);
   U9396 : NAND2_X2 port map( A1 => n18298, A2 => n18299, ZN => n19445);
   U9405 : XOR2_X1 port map( A1 => n12622, A2 => n30038, Z => n625);
   U9406 : NAND2_X2 port map( A1 => n32230, A2 => n16857, ZN => n20733);
   U9410 : AOI21_X2 port map( A1 => n22327, A2 => n722, B => n22328, ZN => 
                           n3512);
   U9411 : XOR2_X1 port map( A1 => n19567, A2 => n32231, Z => n2484);
   U9412 : XOR2_X1 port map( A1 => n19386, A2 => n34119, Z => n19567);
   U9413 : NOR2_X1 port map( A1 => n19061, A2 => n19063, ZN => n28498);
   U9414 : NOR2_X1 port map( A1 => n19108, A2 => n5545, ZN => n19061);
   U9416 : XOR2_X1 port map( A1 => n32232, A2 => n1433, Z => Ciphertext(35));
   U9417 : AOI22_X1 port map( A1 => n25007, A2 => n25008, B1 => n3155, B2 => 
                           n29110, ZN => n32232);
   U9419 : INV_X2 port map( I => n5820, ZN => n32234);
   U9424 : XOR2_X1 port map( A1 => n32235, A2 => n1406, Z => Ciphertext(26));
   U9429 : NAND2_X2 port map( A1 => n29904, A2 => n27840, ZN => n32240);
   U9432 : XOR2_X1 port map( A1 => n12972, A2 => n19529, Z => n19533);
   U9435 : XOR2_X1 port map( A1 => n30539, A2 => n5038, Z => n11850);
   U9437 : XOR2_X1 port map( A1 => n16200, A2 => n33274, Z => n30539);
   U9440 : OAI22_X2 port map( A1 => n14161, A2 => n10978, B1 => n7397, B2 => 
                           n32236, ZN => n10159);
   U9441 : OAI21_X1 port map( A1 => n1353, A2 => n20627, B => n20628, ZN => 
                           n32236);
   U9444 : AOI22_X2 port map( A1 => n9014, A2 => n7552, B1 => n20627, B2 => 
                           n29814, ZN => n10978);
   U9447 : XOR2_X1 port map( A1 => n18929, A2 => n19538, Z => n9636);
   U9455 : NAND2_X2 port map( A1 => n28108, A2 => n9637, ZN => n19538);
   U9461 : NAND2_X2 port map( A1 => n2576, A2 => n16023, ZN => n26386);
   U9465 : OAI21_X2 port map( A1 => n14869, A2 => n14871, B => n21684, ZN => 
                           n22295);
   U9466 : NOR2_X2 port map( A1 => n14292, A2 => n32237, ZN => n2577);
   U9467 : NOR3_X2 port map( A1 => n33641, A2 => n28287, A3 => n11915, ZN => 
                           n32237);
   U9469 : XOR2_X1 port map( A1 => n32238, A2 => n13886, Z => n27503);
   U9470 : XOR2_X1 port map( A1 => n21039, A2 => n20799, Z => n32238);
   U9472 : XOR2_X1 port map( A1 => n2920, A2 => n4362, Z => n9161);
   U9473 : NOR2_X2 port map( A1 => n5872, A2 => n4150, ZN => n2920);
   U9474 : NOR2_X2 port map( A1 => n12522, A2 => n11181, ZN => n11180);
   U9477 : OR2_X2 port map( A1 => n16, A2 => n11913, Z => n4371);
   U9478 : XOR2_X1 port map( A1 => n887, A2 => n5297, Z => n5296);
   U9479 : XNOR2_X1 port map( A1 => n5482, A2 => n34016, ZN => n22164);
   U9480 : NOR2_X2 port map( A1 => n27053, A2 => n21831, ZN => n34016);
   U9482 : AOI22_X2 port map( A1 => n32241, A2 => n21321, B1 => n4382, B2 => 
                           n21324, ZN => n30745);
   U9484 : NOR2_X2 port map( A1 => n15015, A2 => n28017, ZN => n32241);
   U9485 : NAND2_X2 port map( A1 => n21727, A2 => n21728, ZN => n5482);
   U9486 : AOI21_X1 port map( A1 => n5112, A2 => n315, B => n314, ZN => n32244)
                           ;
   U9487 : NAND2_X2 port map( A1 => n5789, A2 => n31948, ZN => n19243);
   U9488 : NAND2_X2 port map( A1 => n5155, A2 => n5154, ZN => n5789);
   U9492 : NAND2_X1 port map( A1 => n23826, A2 => n16467, ZN => n27734);
   U9496 : AOI22_X1 port map( A1 => n17760, A2 => n31907, B1 => n15282, B2 => 
                           n14365, ZN => n14470);
   U9499 : NAND2_X2 port map( A1 => n16804, A2 => n15198, ZN => n31907);
   U9506 : OAI21_X2 port map( A1 => n9652, A2 => n26081, B => n26518, ZN => 
                           n31036);
   U9508 : NOR2_X2 port map( A1 => n33718, A2 => n6290, ZN => n26081);
   U9509 : NAND2_X2 port map( A1 => n27079, A2 => n6189, ZN => n23474);
   U9510 : OAI22_X2 port map( A1 => n23832, A2 => n7005, B1 => n15623, B2 => 
                           n34167, ZN => n13936);
   U9511 : INV_X2 port map( I => n23587, ZN => n7005);
   U9513 : AND2_X1 port map( A1 => n22640, A2 => n11749, Z => n14830);
   U9514 : XOR2_X1 port map( A1 => n23280, A2 => n11326, Z => n47);
   U9517 : XOR2_X1 port map( A1 => n30315, A2 => n23405, Z => n23280);
   U9519 : NAND2_X1 port map( A1 => n22748, A2 => n30231, ZN => n23027);
   U9523 : NOR2_X2 port map( A1 => n22729, A2 => n22731, ZN => n30231);
   U9524 : INV_X1 port map( I => n7052, ZN => n33183);
   U9526 : OAI21_X2 port map( A1 => n11280, A2 => n10828, B => n11278, ZN => 
                           n18669);
   U9527 : XNOR2_X1 port map( A1 => n16641, A2 => n16472, ZN => n32251);
   U9528 : XOR2_X1 port map( A1 => n9877, A2 => n32245, Z => n21330);
   U9531 : XOR2_X1 port map( A1 => n32614, A2 => n30045, Z => n32245);
   U9535 : NOR3_X2 port map( A1 => n32246, A2 => n26465, A3 => n26464, ZN => 
                           n11845);
   U9538 : NOR2_X1 port map( A1 => n3289, A2 => n3288, ZN => n32246);
   U9548 : XOR2_X1 port map( A1 => n30997, A2 => n1396, Z => n6852);
   U9552 : NOR2_X2 port map( A1 => n31032, A2 => n34148, ZN => n30997);
   U9553 : AOI21_X2 port map( A1 => n32247, A2 => n33223, B => n31293, ZN => 
                           n24330);
   U9554 : AOI21_X1 port map( A1 => n33144, A2 => n3860, B => n14335, ZN => 
                           n32247);
   U9555 : NAND2_X2 port map( A1 => n23885, A2 => n15266, ZN => n17777);
   U9556 : NAND2_X1 port map( A1 => n17502, A2 => n32438, ZN => n32338);
   U9557 : XOR2_X1 port map( A1 => n22061, A2 => n22109, Z => n5353);
   U9561 : XOR2_X1 port map( A1 => n1310, A2 => n5476, Z => n22109);
   U9565 : XOR2_X1 port map( A1 => n5186, A2 => n28315, Z => n20716);
   U9566 : XOR2_X1 port map( A1 => n28953, A2 => n2356, Z => n5186);
   U9569 : BUF_X2 port map( I => n17439, Z => n32248);
   U9571 : AOI21_X2 port map( A1 => n20186, A2 => n20187, B => n32249, ZN => 
                           n7889);
   U9574 : XOR2_X1 port map( A1 => n28621, A2 => n32250, Z => n26162);
   U9580 : XOR2_X1 port map( A1 => n20806, A2 => n32251, Z => n32250);
   U9581 : NAND2_X2 port map( A1 => n13989, A2 => n32147, ZN => n29802);
   U9584 : NAND2_X2 port map( A1 => n11300, A2 => n32254, ZN => n32535);
   U9589 : OAI22_X2 port map( A1 => n31604, A2 => n11306, B1 => n12000, B2 => 
                           n32585, ZN => n13483);
   U9590 : INV_X1 port map( I => n27152, ZN => n33943);
   U9594 : OAI21_X2 port map( A1 => n26337, A2 => n11301, B => n29997, ZN => 
                           n32254);
   U9598 : BUF_X4 port map( I => n28278, Z => n33981);
   U9599 : OAI22_X2 port map( A1 => n1125, A2 => n5440, B1 => n22588, B2 => 
                           n22589, ZN => n12899);
   U9600 : XOR2_X1 port map( A1 => n2653, A2 => n32906, Z => n23290);
   U9601 : NAND2_X1 port map( A1 => n8373, A2 => n16154, ZN => n9151);
   U9602 : XOR2_X1 port map( A1 => n28814, A2 => n32256, Z => n4798);
   U9603 : XOR2_X1 port map( A1 => n28354, A2 => n20974, Z => n32256);
   U9607 : OAI22_X2 port map( A1 => n5782, A2 => n27876, B1 => n266, B2 => 
                           n20495, ZN => n5668);
   U9608 : NOR2_X2 port map( A1 => n32257, A2 => n29354, ZN => n28733);
   U9609 : NOR2_X2 port map( A1 => n9364, A2 => n31721, ZN => n32257);
   U9613 : INV_X2 port map( I => n8862, ZN => n33884);
   U9616 : NAND2_X2 port map( A1 => n33022, A2 => n17327, ZN => n32258);
   U9617 : XOR2_X1 port map( A1 => n32259, A2 => n4704, Z => n7896);
   U9619 : OAI21_X2 port map( A1 => n18959, A2 => n4622, B => n4619, ZN => 
                           n32259);
   U9620 : NOR2_X2 port map( A1 => n4390, A2 => n32260, ZN => n21842);
   U9622 : AOI21_X1 port map( A1 => n3916, A2 => n14482, B => n33454, ZN => 
                           n32260);
   U9623 : NAND2_X2 port map( A1 => n1965, A2 => n32261, ZN => n6357);
   U9627 : NOR2_X2 port map( A1 => n1968, A2 => n1967, ZN => n32261);
   U9629 : XOR2_X1 port map( A1 => n32262, A2 => n25993, Z => n19565);
   U9633 : AOI21_X2 port map( A1 => n31349, A2 => n14606, B => n19303, ZN => 
                           n25993);
   U9638 : INV_X2 port map( I => n19483, ZN => n32262);
   U9640 : OAI21_X2 port map( A1 => n13414, A2 => n1519, B => n32754, ZN => 
                           n28839);
   U9643 : OAI21_X2 port map( A1 => n12312, A2 => n32263, B => n6003, ZN => 
                           n31718);
   U9644 : NOR2_X2 port map( A1 => n32264, A2 => n24097, ZN => n32263);
   U9646 : INV_X2 port map( I => n32917, ZN => n32264);
   U9647 : NAND2_X2 port map( A1 => n22765, A2 => n29795, ZN => n29634);
   U9649 : NAND2_X2 port map( A1 => n23631, A2 => n32265, ZN => n24286);
   U9652 : NAND2_X2 port map( A1 => n32426, A2 => n6392, ZN => n32265);
   U9654 : OAI21_X2 port map( A1 => n33470, A2 => n31788, B => n32266, ZN => 
                           n24761);
   U9657 : NAND2_X1 port map( A1 => n1640, A2 => n14447, ZN => n32266);
   U9658 : INV_X2 port map( I => n29540, ZN => n15708);
   U9662 : XOR2_X1 port map( A1 => n32267, A2 => n19368, Z => n29540);
   U9663 : INV_X2 port map( I => n6387, ZN => n32267);
   U9665 : INV_X2 port map( I => n24914, ZN => n24911);
   U9666 : NAND2_X2 port map( A1 => n29877, A2 => n17304, ZN => n24914);
   U9669 : INV_X1 port map( I => n23729, ZN => n30477);
   U9670 : NAND2_X1 port map( A1 => n15722, A2 => n30949, ZN => n23729);
   U9671 : AOI22_X2 port map( A1 => n1219, A2 => n9862, B1 => n837, B2 => n9861
                           , ZN => n33737);
   U9672 : XOR2_X1 port map( A1 => n7250, A2 => n22125, Z => n3395);
   U9673 : NAND2_X2 port map( A1 => n11585, A2 => n6076, ZN => n7250);
   U9676 : XOR2_X1 port map( A1 => n32268, A2 => n23375, Z => n33710);
   U9680 : XOR2_X1 port map( A1 => n23376, A2 => n23475, Z => n32268);
   U9681 : NAND2_X2 port map( A1 => n33239, A2 => n32269, ZN => n24896);
   U9685 : NAND3_X1 port map( A1 => n24477, A2 => n24591, A3 => n25013, ZN => 
                           n32269);
   U9688 : BUF_X2 port map( I => n3964, Z => n32271);
   U9697 : XOR2_X1 port map( A1 => n32272, A2 => n25554, Z => Ciphertext(123));
   U9699 : INV_X1 port map( I => n31389, ZN => n33357);
   U9700 : INV_X2 port map( I => n20581, ZN => n936);
   U9704 : NAND2_X2 port map( A1 => n9449, A2 => n19657, ZN => n20581);
   U9708 : INV_X4 port map( I => n24326, ZN => n24325);
   U9710 : NAND2_X2 port map( A1 => n32274, A2 => n33335, ZN => n33980);
   U9713 : NAND2_X2 port map( A1 => n10353, A2 => n10352, ZN => n32274);
   U9715 : NAND3_X2 port map( A1 => n10261, A2 => n6599, A3 => n28395, ZN => 
                           n33286);
   U9716 : NAND2_X2 port map( A1 => n32275, A2 => n27269, ZN => n17637);
   U9717 : AOI22_X2 port map( A1 => n15979, A2 => n15964, B1 => n24865, B2 => 
                           n26912, ZN => n32275);
   U9720 : NAND2_X2 port map( A1 => n27856, A2 => n27916, ZN => n27419);
   U9721 : INV_X1 port map( I => n20798, ZN => n32392);
   U9723 : NAND2_X1 port map( A1 => n32278, A2 => n32276, ZN => n19457);
   U9727 : INV_X1 port map( I => n8770, ZN => n32277);
   U9728 : NAND2_X1 port map( A1 => n1034, A2 => n8770, ZN => n32278);
   U9732 : NAND2_X2 port map( A1 => n27337, A2 => n21394, ZN => n14095);
   U9735 : OAI21_X1 port map( A1 => n25740, A2 => n27189, B => n32279, ZN => 
                           n6524);
   U9736 : XOR2_X1 port map( A1 => n5024, A2 => n20885, Z => n15875);
   U9738 : NAND2_X2 port map( A1 => n2292, A2 => n2293, ZN => n20549);
   U9739 : AOI21_X2 port map( A1 => n24269, A2 => n24268, B => n11721, ZN => 
                           n11723);
   U9741 : NAND2_X2 port map( A1 => n32280, A2 => n33821, ZN => n26445);
   U9743 : NAND2_X1 port map( A1 => n30562, A2 => n14803, ZN => n32280);
   U9745 : NOR2_X2 port map( A1 => n15326, A2 => n15327, ZN => n33646);
   U9746 : AOI22_X2 port map( A1 => n26633, A2 => n20577, B1 => n20481, B2 => 
                           n20480, ZN => n6228);
   U9754 : INV_X2 port map( I => n12008, ZN => n4674);
   U9757 : NAND2_X1 port map( A1 => n28645, A2 => n20067, ZN => n26741);
   U9763 : NAND2_X2 port map( A1 => n942, A2 => n19947, ZN => n19948);
   U9766 : NAND2_X2 port map( A1 => n7799, A2 => n32281, ZN => n7798);
   U9768 : NAND2_X2 port map( A1 => n20487, A2 => n9808, ZN => n32281);
   U9769 : OR2_X1 port map( A1 => n24153, A2 => n839, Z => n32962);
   U9770 : NOR2_X1 port map( A1 => n6326, A2 => n6325, ZN => n6982);
   U9774 : XOR2_X1 port map( A1 => n32283, A2 => n19412, Z => n1694);
   U9775 : AOI21_X2 port map( A1 => n18938, A2 => n29, B => n18937, ZN => 
                           n19412);
   U9777 : INV_X1 port map( I => n19400, ZN => n32283);
   U9778 : NAND2_X2 port map( A1 => n3983, A2 => n11654, ZN => n31155);
   U9784 : XOR2_X1 port map( A1 => n32284, A2 => n8487, Z => Ciphertext(64));
   U9786 : NAND3_X2 port map( A1 => n8340, A2 => n8928, A3 => n8339, ZN => 
                           n32284);
   U9788 : XOR2_X1 port map( A1 => n32285, A2 => n7665, Z => n7700);
   U9791 : XOR2_X1 port map( A1 => n23424, A2 => n23307, Z => n32285);
   U9793 : AOI22_X2 port map( A1 => n7719, A2 => n16174, B1 => n34052, B2 => 
                           n20515, ZN => n2251);
   U9794 : NAND2_X2 port map( A1 => n3725, A2 => n3724, ZN => n4782);
   U9797 : NOR2_X2 port map( A1 => n9615, A2 => n9609, ZN => n3725);
   U9798 : NAND2_X2 port map( A1 => n31282, A2 => n22464, ZN => n22962);
   U9800 : OAI21_X2 port map( A1 => n16288, A2 => n25999, B => n8233, ZN => 
                           n16068);
   U9802 : XOR2_X1 port map( A1 => n17004, A2 => n9440, Z => n16689);
   U9811 : AND2_X1 port map( A1 => n21357, A2 => n21358, Z => n11655);
   U9814 : NAND2_X2 port map( A1 => n32287, A2 => n3451, ZN => n5915);
   U9815 : OAI21_X2 port map( A1 => n3454, A2 => n3596, B => n31931, ZN => 
                           n32287);
   U9816 : INV_X4 port map( I => n29980, ZN => n28581);
   U9818 : NAND2_X2 port map( A1 => n30972, A2 => n28523, ZN => n29980);
   U9819 : XOR2_X1 port map( A1 => n4883, A2 => n19705, Z => n3416);
   U9820 : XOR2_X1 port map( A1 => n12779, A2 => n16150, Z => n33804);
   U9822 : NAND2_X2 port map( A1 => n8478, A2 => n4114, ZN => n33069);
   U9824 : AOI22_X2 port map( A1 => n31919, A2 => n24292, B1 => n7779, B2 => 
                           n26544, ZN => n32288);
   U9825 : NAND2_X2 port map( A1 => n14711, A2 => n14712, ZN => n20414);
   U9826 : NOR2_X2 port map( A1 => n5820, A2 => n16976, ZN => n22772);
   U9829 : INV_X1 port map( I => n2913, ZN => n32299);
   U9830 : NAND2_X2 port map( A1 => n33458, A2 => n32298, ZN => n32289);
   U9831 : NAND2_X2 port map( A1 => n16787, A2 => n32329, ZN => n26485);
   U9833 : NAND2_X2 port map( A1 => n11035, A2 => n11036, ZN => n16787);
   U9835 : INV_X4 port map( I => n33035, ZN => n15027);
   U9836 : NAND2_X2 port map( A1 => n18170, A2 => n18171, ZN => n20208);
   U9837 : AOI21_X1 port map( A1 => n16444, A2 => n19061, B => n32290, ZN => 
                           n7591);
   U9839 : NOR2_X1 port map( A1 => n29213, A2 => n571, ZN => n29423);
   U9841 : NOR2_X1 port map( A1 => n26406, A2 => n16148, ZN => n32406);
   U9843 : NAND2_X2 port map( A1 => n32291, A2 => n20884, ZN => n21693);
   U9844 : AOI22_X2 port map( A1 => n812, A2 => n20881, B1 => n21163, B2 => 
                           n21367, ZN => n32291);
   U9845 : OAI21_X2 port map( A1 => n33488, A2 => n31239, B => n29964, ZN => 
                           n31497);
   U9846 : OR2_X1 port map( A1 => n19122, A2 => n16361, Z => n32292);
   U9854 : NAND2_X2 port map( A1 => n10043, A2 => n18617, ZN => n18615);
   U9855 : XOR2_X1 port map( A1 => n8392, A2 => n22032, Z => n22154);
   U9856 : NAND2_X2 port map( A1 => n3702, A2 => n33315, ZN => n8392);
   U9858 : XOR2_X1 port map( A1 => n26272, A2 => n6031, Z => n11006);
   U9860 : OAI21_X2 port map( A1 => n14536, A2 => n31115, B => n32294, ZN => 
                           n10055);
   U9863 : XOR2_X1 port map( A1 => n3267, A2 => n32295, Z => n29470);
   U9864 : XOR2_X1 port map( A1 => n17859, A2 => n23400, Z => n32295);
   U9866 : BUF_X2 port map( I => n1164, Z => n32296);
   U9871 : NAND2_X2 port map( A1 => n32297, A2 => n4816, ZN => n15275);
   U9872 : OAI22_X2 port map( A1 => n20479, A2 => n20403, B1 => n20571, B2 => 
                           n31968, ZN => n32297);
   U9873 : XOR2_X1 port map( A1 => n31523, A2 => n16578, Z => n2875);
   U9875 : NAND2_X2 port map( A1 => n4846, A2 => n4847, ZN => n31523);
   U9882 : NOR2_X2 port map( A1 => n26595, A2 => n32300, ZN => n13884);
   U9884 : NOR2_X2 port map( A1 => n32384, A2 => n8029, ZN => n32301);
   U9885 : NOR2_X2 port map( A1 => n10862, A2 => n26410, ZN => n22401);
   U9889 : XOR2_X1 port map( A1 => n28315, A2 => n20873, Z => n32726);
   U9890 : INV_X2 port map( I => n16805, ZN => n18677);
   U9892 : XOR2_X1 port map( A1 => Plaintext(2), A2 => Key(2), Z => n16805);
   U9897 : XOR2_X1 port map( A1 => n9018, A2 => n32302, Z => n33331);
   U9899 : XOR2_X1 port map( A1 => n23355, A2 => n23292, Z => n11249);
   U9900 : XOR2_X1 port map( A1 => n27423, A2 => n18028, Z => n24561);
   U9912 : AOI21_X2 port map( A1 => n342, A2 => n30579, B => n33124, ZN => 
                           n27423);
   U9913 : XOR2_X1 port map( A1 => n32303, A2 => n16497, Z => Ciphertext(108));
   U9918 : NAND3_X1 port map( A1 => n31492, A2 => n25482, A3 => n25458, ZN => 
                           n32303);
   U9920 : NAND2_X2 port map( A1 => n32304, A2 => n31078, ZN => n20996);
   U9921 : NAND2_X2 port map( A1 => n17496, A2 => n32305, ZN => n17497);
   U9932 : AOI22_X2 port map( A1 => n29338, A2 => n34152, B1 => n12075, B2 => 
                           n20052, ZN => n32305);
   U9938 : XOR2_X1 port map( A1 => n24691, A2 => n5762, Z => n30563);
   U9949 : NAND2_X2 port map( A1 => n32725, A2 => n31171, ZN => n24691);
   U9952 : NAND3_X1 port map( A1 => n25285, A2 => n16291, A3 => n25276, ZN => 
                           n11257);
   U9954 : NAND2_X2 port map( A1 => n10743, A2 => n33330, ZN => n16291);
   U9955 : XOR2_X1 port map( A1 => n32306, A2 => n16705, Z => Ciphertext(134));
   U9957 : NAND2_X1 port map( A1 => n13996, A2 => n28775, ZN => n32306);
   U9961 : NAND3_X2 port map( A1 => n29741, A2 => n11109, A3 => n11108, ZN => 
                           n23358);
   U9962 : NAND2_X1 port map( A1 => n15241, A2 => n15242, ZN => n34000);
   U9967 : OAI22_X2 port map( A1 => n19329, A2 => n2040, B1 => n19328, B2 => 
                           n7732, ZN => n18103);
   U9969 : INV_X1 port map( I => n20911, ZN => n32342);
   U9971 : BUF_X4 port map( I => n28839, Z => n33022);
   U9973 : NAND2_X1 port map( A1 => n22885, A2 => n1577, ZN => n32307);
   U9975 : NOR2_X2 port map( A1 => n32308, A2 => n10193, ZN => n6320);
   U9976 : NAND2_X2 port map( A1 => n14412, A2 => n14410, ZN => n11651);
   U9977 : NOR2_X2 port map( A1 => n26079, A2 => n14249, ZN => n14412);
   U9982 : AND2_X1 port map( A1 => n28697, A2 => n22982, Z => n22837);
   U9985 : NAND3_X1 port map( A1 => n12293, A2 => n12295, A3 => n17928, ZN => 
                           n32583);
   U9987 : XOR2_X1 port map( A1 => n22075, A2 => n22141, Z => n22267);
   U9988 : AOI22_X2 port map( A1 => n6968, A2 => n15676, B1 => n12794, B2 => 
                           n6967, ZN => n22141);
   U9989 : NOR2_X2 port map( A1 => n27501, A2 => n24158, ZN => n24067);
   U9990 : XOR2_X1 port map( A1 => n13645, A2 => n19624, Z => n16080);
   U10002 : AOI21_X2 port map( A1 => n8906, A2 => n11955, B => n30209, ZN => 
                           n13645);
   U10003 : NAND2_X2 port map( A1 => n32312, A2 => n32311, ZN => n25816);
   U10006 : INV_X2 port map( I => n32313, ZN => n14661);
   U10009 : XNOR2_X1 port map( A1 => n6721, A2 => n6719, ZN => n32313);
   U10010 : NAND3_X2 port map( A1 => n32314, A2 => n6176, A3 => n16601, ZN => 
                           n18163);
   U10012 : OR2_X2 port map( A1 => n9717, A2 => n32315, Z => n691);
   U10015 : OAI22_X1 port map( A1 => n28283, A2 => n2378, B1 => n12230, B2 => 
                           n10497, ZN => n32315);
   U10017 : AOI22_X2 port map( A1 => n22780, A2 => n11983, B1 => n31824, B2 => 
                           n22848, ZN => n22889);
   U10025 : OR2_X1 port map( A1 => n7581, A2 => n1808, Z => n33894);
   U10033 : NAND2_X2 port map( A1 => n6581, A2 => n32317, ZN => n23981);
   U10035 : XOR2_X1 port map( A1 => n1991, A2 => n32316, Z => n33082);
   U10036 : XOR2_X1 port map( A1 => n1990, A2 => n31928, Z => n32316);
   U10037 : INV_X2 port map( I => n7188, ZN => n32317);
   U10038 : NAND2_X2 port map( A1 => n32453, A2 => n3950, ZN => n6555);
   U10040 : NAND4_X1 port map( A1 => n6730, A2 => n4056, A3 => n25572, A4 => 
                           n25573, ZN => n32702);
   U10050 : NAND2_X2 port map( A1 => n15060, A2 => n11953, ZN => n15059);
   U10052 : NOR2_X2 port map( A1 => n22704, A2 => n32318, ZN => n30532);
   U10053 : XOR2_X1 port map( A1 => n32319, A2 => n3605, Z => n11110);
   U10056 : XOR2_X1 port map( A1 => n22000, A2 => n12882, Z => n32319);
   U10057 : NAND2_X1 port map( A1 => n17240, A2 => n11974, ZN => n24484);
   U10059 : XOR2_X1 port map( A1 => n24638, A2 => n24474, Z => n24773);
   U10061 : AOI22_X2 port map( A1 => n14847, A2 => n29566, B1 => n23781, B2 => 
                           n17280, ZN => n24638);
   U10062 : NAND2_X2 port map( A1 => n32322, A2 => n33171, ZN => n3963);
   U10066 : NAND2_X2 port map( A1 => n32877, A2 => n24060, ZN => n12644);
   U10071 : AND2_X2 port map( A1 => n652, A2 => n23201, Z => n23796);
   U10075 : NAND2_X1 port map( A1 => n15211, A2 => n28078, ZN => n26068);
   U10076 : AOI21_X2 port map( A1 => n29648, A2 => n32089, B => n32324, ZN => 
                           n16635);
   U10079 : XOR2_X1 port map( A1 => n4314, A2 => n19370, Z => n19742);
   U10084 : AOI21_X2 port map( A1 => n7186, A2 => n7187, B => n7185, ZN => 
                           n4314);
   U10088 : XOR2_X1 port map( A1 => n1085, A2 => n5539, Z => n30917);
   U10090 : NOR2_X2 port map( A1 => n17822, A2 => n32325, ZN => n10735);
   U10091 : BUF_X2 port map( I => n32807, Z => n32326);
   U10092 : AOI21_X2 port map( A1 => n13227, A2 => n16485, B => n32327, ZN => 
                           n19583);
   U10096 : AOI21_X2 port map( A1 => n19186, A2 => n13226, B => n13685, ZN => 
                           n32327);
   U10103 : NAND2_X2 port map( A1 => n9995, A2 => n9998, ZN => n24110);
   U10107 : NOR2_X2 port map( A1 => n22483, A2 => n22372, ZN => n33864);
   U10110 : INV_X8 port map( I => n18515, ZN => n829);
   U10112 : AOI22_X2 port map( A1 => n33240, A2 => n11666, B1 => n16492, B2 => 
                           n20227, ZN => n11665);
   U10113 : NOR2_X2 port map( A1 => n32326, A2 => n11364, ZN => n1361);
   U10114 : XOR2_X1 port map( A1 => n27192, A2 => n5322, Z => n32807);
   U10116 : AOI22_X2 port map( A1 => n30507, A2 => n1290, B1 => n22439, B2 => 
                           n12899, ZN => n23018);
   U10125 : NAND2_X2 port map( A1 => n12434, A2 => n27551, ZN => n14619);
   U10127 : NOR2_X1 port map( A1 => n8994, A2 => n20319, ZN => n32440);
   U10128 : AOI21_X2 port map( A1 => n19270, A2 => n19271, B => n19269, ZN => 
                           n19272);
   U10130 : NAND2_X2 port map( A1 => n15961, A2 => n32330, ZN => n21553);
   U10133 : NAND2_X2 port map( A1 => n32670, A2 => n32331, ZN => n9408);
   U10137 : OR2_X1 port map( A1 => n27131, A2 => n19275, Z => n32332);
   U10141 : INV_X4 port map( I => n31579, ZN => n18643);
   U10142 : NOR2_X2 port map( A1 => n1008, A2 => n32333, ZN => n33298);
   U10169 : NAND2_X2 port map( A1 => n10699, A2 => n915, ZN => n32333);
   U10170 : OAI21_X1 port map( A1 => n1581, A2 => n5260, B => n5259, ZN => 
                           n5261);
   U10171 : XOR2_X1 port map( A1 => n11297, A2 => n24520, Z => n24654);
   U10173 : NAND2_X2 port map( A1 => n30732, A2 => n17233, ZN => n11297);
   U10176 : NOR2_X1 port map( A1 => n32335, A2 => n32334, ZN => n8222);
   U10178 : NOR2_X1 port map( A1 => n9456, A2 => n22660, ZN => n32335);
   U10179 : XOR2_X1 port map( A1 => n15606, A2 => n31457, Z => n22182);
   U10185 : NAND2_X2 port map( A1 => n12273, A2 => n9448, ZN => n15606);
   U10192 : NAND3_X2 port map( A1 => n20351, A2 => n28813, A3 => n20350, ZN => 
                           n12364);
   U10194 : OAI22_X2 port map( A1 => n25456, A2 => n32869, B1 => n25454, B2 => 
                           n25455, ZN => n33248);
   U10195 : NOR2_X2 port map( A1 => n408, A2 => n25433, ZN => n25456);
   U10202 : XOR2_X1 port map( A1 => n7889, A2 => n20961, Z => n21025);
   U10247 : NAND3_X1 port map( A1 => n891, A2 => n24221, A3 => n2539, ZN => 
                           n9542);
   U10254 : INV_X1 port map( I => n8168, ZN => n30285);
   U10262 : XOR2_X1 port map( A1 => n6267, A2 => n12083, Z => n17044);
   U10264 : AOI22_X2 port map( A1 => n11566, A2 => n11565, B1 => n11564, B2 => 
                           n22705, ZN => n32705);
   U10265 : NAND2_X2 port map( A1 => n11132, A2 => n25289, ZN => n25290);
   U10270 : NAND2_X2 port map( A1 => n32338, A2 => n22755, ZN => n12821);
   U10271 : OAI22_X2 port map( A1 => n32339, A2 => n8614, B1 => n8613, B2 => 
                           n31271, ZN => n12593);
   U10272 : NOR2_X2 port map( A1 => n1978, A2 => n8615, ZN => n32339);
   U10276 : INV_X1 port map( I => n23369, ZN => n33929);
   U10282 : XOR2_X1 port map( A1 => n24650, A2 => n32340, Z => n28443);
   U10283 : XOR2_X1 port map( A1 => n28579, A2 => n29589, Z => n32340);
   U10284 : XOR2_X1 port map( A1 => n6731, A2 => n19730, Z => n26702);
   U10288 : XOR2_X1 port map( A1 => n19558, A2 => n19474, Z => n19730);
   U10289 : NAND2_X2 port map( A1 => n27832, A2 => n29200, ZN => n33875);
   U10291 : NAND2_X2 port map( A1 => n9610, A2 => n2456, ZN => n3724);
   U10293 : OR2_X2 port map( A1 => n6359, A2 => n2019, Z => n10844);
   U10295 : XOR2_X1 port map( A1 => n1622, A2 => n1621, Z => n11628);
   U10300 : XOR2_X1 port map( A1 => n32342, A2 => n7630, Z => n6159);
   U10303 : NAND2_X2 port map( A1 => n6157, A2 => n4269, ZN => n7630);
   U10305 : AND2_X1 port map( A1 => n20097, A2 => n27832, Z => n8146);
   U10306 : NAND2_X2 port map( A1 => n4708, A2 => n32343, ZN => n5091);
   U10307 : XOR2_X1 port map( A1 => n24021, A2 => n32345, Z => n26126);
   U10308 : XOR2_X1 port map( A1 => n2278, A2 => n32346, Z => n32345);
   U10313 : NAND3_X1 port map( A1 => n5471, A2 => n20375, A3 => n10939, ZN => 
                           n2317);
   U10314 : NAND2_X1 port map( A1 => n9259, A2 => n30838, ZN => n7278);
   U10315 : INV_X2 port map( I => n29215, ZN => n6842);
   U10316 : NAND2_X1 port map( A1 => n32347, A2 => n29215, ZN => n30852);
   U10337 : XOR2_X1 port map( A1 => n6843, A2 => n32464, Z => n29215);
   U10339 : INV_X2 port map( I => n6855, ZN => n32347);
   U10345 : NAND2_X1 port map( A1 => n32617, A2 => n28554, ZN => n22329);
   U10346 : NAND2_X2 port map( A1 => n32348, A2 => n32039, ZN => n21544);
   U10347 : NAND2_X2 port map( A1 => n32506, A2 => n32505, ZN => n26206);
   U10348 : BUF_X2 port map( I => n24207, Z => n32349);
   U10351 : INV_X1 port map( I => n27842, ZN => n32351);
   U10353 : AOI22_X2 port map( A1 => n7262, A2 => n28265, B1 => n707, B2 => 
                           n7263, ZN => n7261);
   U10354 : INV_X2 port map( I => n32352, ZN => n29272);
   U10356 : XNOR2_X1 port map( A1 => n7711, A2 => n33118, ZN => n32352);
   U10357 : XOR2_X1 port map( A1 => n32353, A2 => n3648, Z => n28554);
   U10375 : XOR2_X1 port map( A1 => n33408, A2 => n22070, Z => n32353);
   U10376 : NOR2_X2 port map( A1 => n5570, A2 => n32355, ZN => n17273);
   U10378 : NOR3_X1 port map( A1 => n26015, A2 => n15738, A3 => n25229, ZN => 
                           n32355);
   U10380 : XOR2_X1 port map( A1 => n18929, A2 => n30075, Z => n30074);
   U10384 : XOR2_X1 port map( A1 => n32356, A2 => n23311, Z => n23827);
   U10386 : XOR2_X1 port map( A1 => n33236, A2 => n14841, Z => n32356);
   U10387 : XOR2_X1 port map( A1 => n32722, A2 => n10236, Z => n28514);
   U10388 : OR2_X1 port map( A1 => n32919, A2 => n17439, Z => n2831);
   U10389 : OAI21_X2 port map( A1 => n11976, A2 => n883, B => n32359, ZN => 
                           n29754);
   U10390 : OAI21_X2 port map( A1 => n4318, A2 => n15152, B => n883, ZN => 
                           n32359);
   U10392 : NAND3_X1 port map( A1 => n26206, A2 => n26207, A3 => n1012, ZN => 
                           n32688);
   U10395 : OAI21_X2 port map( A1 => n29758, A2 => n29469, B => n22459, ZN => 
                           n14129);
   U10405 : XOR2_X1 port map( A1 => n8018, A2 => n32360, Z => n31771);
   U10406 : XOR2_X1 port map( A1 => n34047, A2 => n7045, Z => n32360);
   U10409 : INV_X1 port map( I => n21248, ZN => n29142);
   U10411 : NAND2_X1 port map( A1 => n13432, A2 => n13433, ZN => n33133);
   U10412 : OR2_X1 port map( A1 => n28308, A2 => n7368, Z => n3889);
   U10414 : XOR2_X1 port map( A1 => n32361, A2 => n25049, Z => Ciphertext(39));
   U10418 : NAND3_X2 port map( A1 => n25048, A2 => n28220, A3 => n25046, ZN => 
                           n32361);
   U10419 : NOR2_X1 port map( A1 => n23793, A2 => n23794, ZN => n1876);
   U10421 : XOR2_X1 port map( A1 => n32362, A2 => n10951, Z => n589);
   U10424 : XOR2_X1 port map( A1 => n28295, A2 => n25578, Z => n32362);
   U10429 : NAND2_X2 port map( A1 => n27299, A2 => n4241, ZN => n20900);
   U10440 : AOI21_X2 port map( A1 => n23482, A2 => n7220, B => n11956, ZN => 
                           n9212);
   U10443 : AND2_X2 port map( A1 => n15559, A2 => n21193, Z => n21072);
   U10444 : XOR2_X1 port map( A1 => n7880, A2 => n32363, Z => n30173);
   U10448 : XOR2_X1 port map( A1 => n6545, A2 => n2045, Z => n32363);
   U10449 : NAND2_X1 port map( A1 => n29753, A2 => n793, ZN => n32369);
   U10451 : XOR2_X1 port map( A1 => n32364, A2 => n23245, Z => n22935);
   U10452 : XOR2_X1 port map( A1 => n33380, A2 => n22932, Z => n32364);
   U10453 : NOR2_X1 port map( A1 => n4386, A2 => n4387, ZN => n32612);
   U10460 : NOR2_X1 port map( A1 => n22953, A2 => n7544, ZN => n8082);
   U10461 : NAND2_X2 port map( A1 => n16267, A2 => n30584, ZN => n7544);
   U10463 : BUF_X4 port map( I => n3286, Z => n21);
   U10465 : NAND2_X2 port map( A1 => n11710, A2 => n20549, ZN => n20327);
   U10466 : NAND2_X2 port map( A1 => n2285, A2 => n26814, ZN => n11710);
   U10467 : NAND2_X2 port map( A1 => n3760, A2 => n981, ZN => n23815);
   U10468 : AND2_X1 port map( A1 => n11734, A2 => n17522, Z => n2603);
   U10470 : XOR2_X1 port map( A1 => n20803, A2 => n20802, Z => n21012);
   U10474 : NAND2_X2 port map( A1 => n20218, A2 => n20217, ZN => n20803);
   U10476 : XOR2_X1 port map( A1 => n33317, A2 => n26642, Z => n17506);
   U10477 : XOR2_X1 port map( A1 => n32365, A2 => n8464, Z => n14934);
   U10482 : XOR2_X1 port map( A1 => n21033, A2 => n15793, Z => n32365);
   U10483 : XOR2_X1 port map( A1 => n32366, A2 => n4610, Z => n32489);
   U10484 : XOR2_X1 port map( A1 => n27481, A2 => n7046, Z => n32366);
   U10487 : BUF_X2 port map( I => n19749, Z => n32367);
   U10491 : XOR2_X1 port map( A1 => n9440, A2 => n22091, Z => n30070);
   U10493 : XOR2_X1 port map( A1 => n22031, A2 => n22243, Z => n22091);
   U10495 : XOR2_X1 port map( A1 => n24356, A2 => n24403, Z => n17798);
   U10502 : NAND3_X2 port map( A1 => n10176, A2 => n10179, A3 => n10175, ZN => 
                           n24356);
   U10504 : NAND2_X2 port map( A1 => n22737, A2 => n2449, ZN => n22944);
   U10505 : OAI22_X2 port map( A1 => n32369, A2 => n6654, B1 => n24073, B2 => 
                           n737, ZN => n6651);
   U10506 : XOR2_X1 port map( A1 => n23489, A2 => n23435, Z => n30390);
   U10509 : OAI21_X2 port map( A1 => n26526, A2 => n22710, B => n8726, ZN => 
                           n23435);
   U10510 : XOR2_X1 port map( A1 => n18911, A2 => n19466, Z => n10210);
   U10514 : NAND2_X2 port map( A1 => n7420, A2 => n27553, ZN => n18911);
   U10515 : OR2_X1 port map( A1 => n10862, A2 => n17185, Z => n12097);
   U10517 : XOR2_X1 port map( A1 => n25993, A2 => n2388, Z => n5861);
   U10519 : INV_X2 port map( I => n12934, ZN => n23488);
   U10520 : NAND2_X2 port map( A1 => n28401, A2 => n4305, ZN => n12934);
   U10521 : NAND2_X1 port map( A1 => n17134, A2 => n34165, ZN => n15997);
   U10535 : NOR2_X1 port map( A1 => n31033, A2 => n32929, ZN => n30626);
   U10537 : NAND2_X1 port map( A1 => n32373, A2 => n32372, ZN => n9350);
   U10538 : INV_X1 port map( I => n32800, ZN => n32374);
   U10539 : XOR2_X1 port map( A1 => n30411, A2 => n19736, Z => n19574);
   U10540 : OAI21_X2 port map( A1 => n19142, A2 => n19141, B => n16875, ZN => 
                           n19736);
   U10543 : AOI22_X2 port map( A1 => n28585, A2 => n33011, B1 => n23747, B2 => 
                           n16628, ZN => n27168);
   U10546 : NAND2_X2 port map( A1 => n11391, A2 => n11393, ZN => n28585);
   U10550 : OAI21_X2 port map( A1 => n20028, A2 => n1042, B => n20025, ZN => 
                           n8244);
   U10553 : INV_X2 port map( I => n14082, ZN => n1042);
   U10556 : XOR2_X1 port map( A1 => n7297, A2 => n7295, Z => n14082);
   U10558 : NOR2_X2 port map( A1 => n15358, A2 => n32375, ZN => n11208);
   U10562 : OAI22_X2 port map( A1 => n21114, A2 => n33741, B1 => n4989, B2 => 
                           n16072, ZN => n32375);
   U10563 : NAND2_X2 port map( A1 => n7974, A2 => n32376, ZN => n25592);
   U10564 : NAND2_X1 port map( A1 => n33095, A2 => n10248, ZN => n32376);
   U10565 : INV_X2 port map( I => n19920, ZN => n32377);
   U10576 : NAND2_X2 port map( A1 => n32746, A2 => n14761, ZN => n19920);
   U10580 : XOR2_X1 port map( A1 => n32379, A2 => n26401, Z => n13022);
   U10585 : XOR2_X1 port map( A1 => n30058, A2 => n10915, Z => n30057);
   U10588 : AOI22_X1 port map( A1 => n15869, A2 => n19227, B1 => n18974, B2 => 
                           n19226, ZN => n13939);
   U10589 : XOR2_X1 port map( A1 => n20992, A2 => n1339, Z => n20654);
   U10592 : XOR2_X1 port map( A1 => n2953, A2 => n32380, Z => n3392);
   U10593 : XOR2_X1 port map( A1 => n3396, A2 => n3393, Z => n32380);
   U10595 : XOR2_X1 port map( A1 => n32381, A2 => n6175, Z => n5962);
   U10596 : XOR2_X1 port map( A1 => n21912, A2 => n297, Z => n32381);
   U10597 : XOR2_X1 port map( A1 => n28803, A2 => n20999, Z => n17524);
   U10600 : XOR2_X1 port map( A1 => n20839, A2 => n30543, Z => n20999);
   U10602 : XOR2_X1 port map( A1 => n23405, A2 => n1102, Z => n23125);
   U10603 : NOR2_X2 port map( A1 => n33585, A2 => n28338, ZN => n25757);
   U10604 : NAND2_X1 port map( A1 => n33610, A2 => n29597, ZN => n22496);
   U10605 : XOR2_X1 port map( A1 => n6502, A2 => n32382, Z => n9796);
   U10606 : XOR2_X1 port map( A1 => n23458, A2 => n11325, Z => n32382);
   U10611 : AOI21_X2 port map( A1 => n13860, A2 => n18687, B => n32383, ZN => 
                           n2593);
   U10616 : NOR3_X2 port map( A1 => n18687, A2 => n18871, A3 => n29308, ZN => 
                           n32383);
   U10617 : NAND2_X2 port map( A1 => n14387, A2 => n18168, ZN => n6593);
   U10618 : XOR2_X1 port map( A1 => n23451, A2 => n23449, Z => n9782);
   U10621 : XOR2_X1 port map( A1 => n770, A2 => n31727, Z => n23449);
   U10622 : NAND2_X2 port map( A1 => n31759, A2 => n32656, ZN => n33832);
   U10625 : XOR2_X1 port map( A1 => n24788, A2 => n24746, Z => n24024);
   U10626 : AOI22_X2 port map( A1 => n28043, A2 => n28085, B1 => n26399, B2 => 
                           n31863, ZN => n32385);
   U10627 : NAND2_X2 port map( A1 => n8117, A2 => n8118, ZN => n8130);
   U10631 : NAND2_X2 port map( A1 => n5825, A2 => n31991, ZN => n8117);
   U10632 : NAND2_X1 port map( A1 => n23750, A2 => n12848, ZN => n33165);
   U10634 : NOR2_X2 port map( A1 => n29648, A2 => n23070, ZN => n4803);
   U10637 : NOR3_X1 port map( A1 => n31272, A2 => n16743, A3 => n32386, ZN => 
                           n20879);
   U10641 : INV_X1 port map( I => n16938, ZN => n32386);
   U10644 : OAI21_X2 port map( A1 => n27535, A2 => n21778, B => n276, ZN => 
                           n12542);
   U10647 : XOR2_X1 port map( A1 => n4741, A2 => n27000, Z => n4740);
   U10655 : INV_X2 port map( I => n14545, ZN => n1157);
   U10656 : NAND2_X2 port map( A1 => n2674, A2 => n28285, ZN => n14545);
   U10657 : XOR2_X1 port map( A1 => n10320, A2 => n31828, Z => n10708);
   U10660 : NAND2_X2 port map( A1 => n32387, A2 => n23178, ZN => n3147);
   U10665 : NAND2_X2 port map( A1 => n31314, A2 => n30470, ZN => n32387);
   U10667 : XOR2_X1 port map( A1 => n31642, A2 => n30636, Z => n30635);
   U10669 : INV_X2 port map( I => n14756, ZN => n23902);
   U10671 : XOR2_X1 port map( A1 => n15548, A2 => n27106, Z => n4192);
   U10674 : XOR2_X1 port map( A1 => n527, A2 => n9810, Z => n31054);
   U10675 : XOR2_X1 port map( A1 => n22030, A2 => n3550, Z => n527);
   U10676 : XOR2_X1 port map( A1 => n27052, A2 => n3126, Z => n3169);
   U10677 : NOR2_X1 port map( A1 => n1360, A2 => n17456, ZN => n8294);
   U10680 : NAND3_X2 port map( A1 => n32388, A2 => n11761, A3 => n11760, ZN => 
                           n15877);
   U10683 : NAND2_X1 port map( A1 => n30503, A2 => n7035, ZN => n32388);
   U10690 : XOR2_X1 port map( A1 => n1993, A2 => n17837, Z => n20558);
   U10697 : NAND2_X2 port map( A1 => n30450, A2 => n32418, ZN => n1993);
   U10698 : AOI22_X2 port map( A1 => n33522, A2 => n32389, B1 => n4803, B2 => 
                           n29070, ZN => n4801);
   U10701 : NOR2_X2 port map( A1 => n29070, A2 => n29648, ZN => n32389);
   U10702 : NAND2_X2 port map( A1 => n23987, A2 => n32390, ZN => n33124);
   U10711 : NAND3_X2 port map( A1 => n8, A2 => n13268, A3 => n8086, ZN => 
                           n32390);
   U10714 : NAND2_X2 port map( A1 => n25966, A2 => n819, ZN => n10000);
   U10716 : NAND2_X1 port map( A1 => n26806, A2 => n24335, ZN => n29388);
   U10717 : XOR2_X1 port map( A1 => n32391, A2 => n17440, Z => n32919);
   U10720 : XOR2_X1 port map( A1 => n27506, A2 => n32392, Z => n32391);
   U10721 : AOI21_X2 port map( A1 => n21206, A2 => n21289, B => n32393, ZN => 
                           n21207);
   U10722 : AOI22_X2 port map( A1 => n20197, A2 => n20531, B1 => n13499, B2 => 
                           n27755, ZN => n27646);
   U10723 : NOR2_X2 port map( A1 => n1155, A2 => n32903, ZN => n20197);
   U10726 : XOR2_X1 port map( A1 => n31295, A2 => n21015, Z => n2786);
   U10727 : XOR2_X1 port map( A1 => n31704, A2 => n14918, Z => n25110);
   U10730 : XOR2_X1 port map( A1 => n1302, A2 => n17745, Z => n9135);
   U10732 : XOR2_X1 port map( A1 => n26863, A2 => n22013, Z => n1302);
   U10735 : NOR2_X2 port map( A1 => n11710, A2 => n28390, ZN => n20550);
   U10736 : XOR2_X1 port map( A1 => n17798, A2 => n24634, Z => n16989);
   U10739 : XOR2_X1 port map( A1 => n14499, A2 => n9943, Z => n4222);
   U10742 : NAND2_X1 port map( A1 => n32394, A2 => n16094, ZN => n33991);
   U10743 : NAND2_X1 port map( A1 => n28990, A2 => n33020, ZN => n32394);
   U10744 : XOR2_X1 port map( A1 => n32395, A2 => n527, Z => n8154);
   U10745 : XOR2_X1 port map( A1 => n13564, A2 => n33072, Z => n32395);
   U10746 : OAI21_X1 port map( A1 => n26471, A2 => n12872, B => n33149, ZN => 
                           n13000);
   U10747 : NAND2_X1 port map( A1 => n13558, A2 => n7004, ZN => n23105);
   U10748 : NAND3_X2 port map( A1 => n14069, A2 => n22568, A3 => n22569, ZN => 
                           n13558);
   U10756 : XOR2_X1 port map( A1 => n32396, A2 => n24398, Z => n16062);
   U10758 : XOR2_X1 port map( A1 => n24395, A2 => n30607, Z => n32396);
   U10759 : BUF_X2 port map( I => n10720, Z => n32397);
   U10761 : OAI21_X2 port map( A1 => n26198, A2 => n965, B => n24947, ZN => 
                           n32398);
   U10766 : AOI21_X2 port map( A1 => n24161, A2 => n30595, B => n3678, ZN => 
                           n30307);
   U10768 : AND2_X1 port map( A1 => n20584, A2 => n20583, Z => n34045);
   U10769 : AOI22_X2 port map( A1 => n17303, A2 => n17302, B1 => n14671, B2 => 
                           n22411, ZN => n33299);
   U10773 : NOR2_X2 port map( A1 => n26305, A2 => n7023, ZN => n17303);
   U10774 : NAND3_X1 port map( A1 => n16664, A2 => n12100, A3 => n20010, ZN => 
                           n19782);
   U10775 : NOR2_X2 port map( A1 => n1140, A2 => n5018, ZN => n6219);
   U10779 : AOI22_X2 port map( A1 => n27088, A2 => n17739, B1 => n23055, B2 => 
                           n2222, ZN => n26900);
   U10780 : NAND2_X2 port map( A1 => n32400, A2 => n18782, ZN => n15166);
   U10782 : NAND2_X2 port map( A1 => n18187, A2 => n30686, ZN => n32400);
   U10784 : XOR2_X1 port map( A1 => n33291, A2 => n27942, Z => n4330);
   U10786 : XOR2_X1 port map( A1 => n23371, A2 => n11504, Z => n23473);
   U10787 : AOI22_X2 port map( A1 => n3692, A2 => n32964, B1 => n3689, B2 => 
                           n13597, ZN => n23371);
   U10788 : NOR2_X2 port map( A1 => n12759, A2 => n12757, ZN => n16641);
   U10789 : NOR2_X2 port map( A1 => n30873, A2 => n32043, ZN => n12759);
   U10791 : XOR2_X1 port map( A1 => n16030, A2 => n33939, Z => n13180);
   U10793 : XNOR2_X1 port map( A1 => n14507, A2 => n8855, ZN => n32502);
   U10796 : AOI22_X2 port map( A1 => n21372, A2 => n21377, B1 => n33774, B2 => 
                           n32907, ZN => n21573);
   U10797 : NOR2_X2 port map( A1 => n21213, A2 => n12525, ZN => n21372);
   U10802 : INV_X1 port map( I => n24787, ZN => n26795);
   U10803 : NAND2_X2 port map( A1 => n6741, A2 => n33489, ZN => n24787);
   U10805 : NAND2_X2 port map( A1 => n29256, A2 => n21079, ZN => n13712);
   U10807 : NAND2_X2 port map( A1 => n10361, A2 => n23086, ZN => n33791);
   U10809 : XOR2_X1 port map( A1 => n32402, A2 => n19766, Z => n5856);
   U10810 : XOR2_X1 port map( A1 => n32587, A2 => n13480, Z => n32402);
   U10812 : XOR2_X1 port map( A1 => n32403, A2 => n20823, Z => n16770);
   U10815 : XOR2_X1 port map( A1 => n16773, A2 => n17759, Z => n32403);
   U10816 : BUF_X4 port map( I => n9172, Z => n4319);
   U10818 : BUF_X2 port map( I => n33437, Z => n32404);
   U10820 : NAND2_X2 port map( A1 => n33784, A2 => n4206, ZN => n5121);
   U10822 : OAI22_X1 port map( A1 => n576, A2 => n5966, B1 => n29153, B2 => 
                           n4373, ZN => n19924);
   U10824 : NOR2_X2 port map( A1 => n32405, A2 => n30294, ZN => n5317);
   U10825 : NOR3_X1 port map( A1 => n17537, A2 => n16337, A3 => n23351, ZN => 
                           n32405);
   U10826 : NAND2_X2 port map( A1 => n32407, A2 => n12018, ZN => n15863);
   U10834 : NAND3_X2 port map( A1 => n16637, A2 => n27938, A3 => n8292, ZN => 
                           n32528);
   U10839 : OR2_X2 port map( A1 => n9920, A2 => n9490, Z => n23933);
   U10840 : XOR2_X1 port map( A1 => n20788, A2 => n21029, Z => n20983);
   U10841 : NAND2_X2 port map( A1 => n31269, A2 => n20612, ZN => n20788);
   U10845 : NOR2_X1 port map( A1 => n32410, A2 => n18687, ZN => n32409);
   U10846 : INV_X2 port map( I => n18871, ZN => n32411);
   U10854 : NOR2_X2 port map( A1 => n5616, A2 => n5613, ZN => n31893);
   U10857 : XOR2_X1 port map( A1 => n12170, A2 => n12172, Z => n20946);
   U10862 : XOR2_X1 port map( A1 => n23137, A2 => n32975, Z => n23168);
   U10865 : NOR2_X2 port map( A1 => n32741, A2 => n29510, ZN => n30824);
   U10867 : XOR2_X1 port map( A1 => n32412, A2 => n22246, Z => n26484);
   U10871 : XOR2_X1 port map( A1 => n8475, A2 => n13651, Z => n32412);
   U10872 : OAI21_X2 port map( A1 => n7228, A2 => n31522, B => n33820, ZN => 
                           n33819);
   U10873 : AOI21_X1 port map( A1 => n33530, A2 => n33225, B => n33222, ZN => 
                           n33224);
   U10874 : AOI21_X2 port map( A1 => n24294, A2 => n24295, B => n29352, ZN => 
                           n32789);
   U10876 : XOR2_X1 port map( A1 => n32413, A2 => n30514, Z => n11877);
   U10877 : XOR2_X1 port map( A1 => n28584, A2 => n20897, Z => n32413);
   U10883 : BUF_X2 port map( I => n27021, Z => n32414);
   U10885 : XOR2_X1 port map( A1 => n13415, A2 => n23285, Z => n31288);
   U10886 : NAND3_X2 port map( A1 => n9791, A2 => n27544, A3 => n22441, ZN => 
                           n23285);
   U10890 : NAND4_X1 port map( A1 => n19235, A2 => n8119, A3 => n8118, A4 => 
                           n8117, ZN => n19894);
   U10897 : OAI21_X2 port map( A1 => n161, A2 => n27345, B => n3310, ZN => 
                           n19235);
   U10898 : XOR2_X1 port map( A1 => n32415, A2 => n7257, Z => n9126);
   U10899 : XOR2_X1 port map( A1 => n24540, A2 => n17448, Z => n32415);
   U10901 : XOR2_X1 port map( A1 => n14337, A2 => n6974, Z => n12972);
   U10903 : NAND2_X1 port map( A1 => n19835, A2 => n32371, ZN => n32416);
   U10906 : XOR2_X1 port map( A1 => n32417, A2 => n1084, Z => n10632);
   U10914 : NAND2_X1 port map( A1 => n3558, A2 => n20404, ZN => n32418);
   U10918 : OAI21_X2 port map( A1 => n26078, A2 => n6581, B => n32419, ZN => 
                           n4956);
   U10919 : NAND3_X1 port map( A1 => n14770, A2 => n6555, A3 => n7188, ZN => 
                           n32419);
   U10920 : XOR2_X1 port map( A1 => n32420, A2 => n27200, Z => n27453);
   U10922 : XOR2_X1 port map( A1 => n30706, A2 => n27778, Z => n32420);
   U10927 : OR2_X1 port map( A1 => n8965, A2 => n17140, Z => n16412);
   U10933 : XOR2_X1 port map( A1 => n9634, A2 => n9635, Z => n10433);
   U10936 : NAND3_X1 port map( A1 => n25045, A2 => n31640, A3 => n27610, ZN => 
                           n25046);
   U10937 : NAND2_X1 port map( A1 => n32422, A2 => n32421, ZN => n24875);
   U10939 : NAND2_X1 port map( A1 => n25015, A2 => n25012, ZN => n32421);
   U10941 : NAND2_X1 port map( A1 => n17240, A2 => n24975, ZN => n32422);
   U10942 : OR2_X2 port map( A1 => n23742, A2 => n15116, Z => n27459);
   U10950 : AND2_X1 port map( A1 => n21438, A2 => n8398, Z => n30646);
   U10954 : XOR2_X1 port map( A1 => n24691, A2 => n25064, Z => n15792);
   U10959 : NOR2_X2 port map( A1 => n7018, A2 => n14411, ZN => n14410);
   U10960 : XOR2_X1 port map( A1 => n91, A2 => n1416, Z => n9308);
   U10962 : NAND2_X2 port map( A1 => n31643, A2 => n29520, ZN => n91);
   U10966 : AOI21_X2 port map( A1 => n32423, A2 => n31483, B => n29773, ZN => 
                           n10710);
   U10969 : NOR2_X2 port map( A1 => n23809, A2 => n14664, ZN => n32423);
   U10972 : OR2_X1 port map( A1 => n2643, A2 => n26782, Z => n21470);
   U10977 : AOI22_X2 port map( A1 => n32424, A2 => n33591, B1 => n2169, B2 => 
                           n17739, ZN => n4847);
   U10979 : NAND3_X2 port map( A1 => n32425, A2 => n27459, A3 => n23769, ZN => 
                           n8286);
   U10980 : NOR3_X2 port map( A1 => n4714, A2 => n32802, A3 => n1049, ZN => 
                           n29768);
   U10983 : OAI22_X2 port map( A1 => n23901, A2 => n5373, B1 => n1254, B2 => 
                           n667, ZN => n32426);
   U10985 : AOI21_X2 port map( A1 => n24888, A2 => n25149, B => n16293, ZN => 
                           n32427);
   U10986 : XOR2_X1 port map( A1 => n2812, A2 => n32428, Z => n13670);
   U10987 : XOR2_X1 port map( A1 => n16178, A2 => n20974, Z => n32428);
   U10993 : XOR2_X1 port map( A1 => n19686, A2 => n19773, Z => n9327);
   U10995 : NAND2_X2 port map( A1 => n30426, A2 => n5329, ZN => n19686);
   U10996 : NOR3_X1 port map( A1 => n31216, A2 => n28270, A3 => n24857, ZN => 
                           n33084);
   U10999 : INV_X2 port map( I => n32429, ZN => n871);
   U11001 : XOR2_X1 port map( A1 => n10722, A2 => n10723, Z => n32429);
   U11007 : NAND2_X2 port map( A1 => n32430, A2 => n23060, ZN => n17775);
   U11009 : NAND2_X2 port map( A1 => n32431, A2 => n33088, ZN => n2073);
   U11011 : NAND2_X2 port map( A1 => n26758, A2 => n32432, ZN => n7287);
   U11017 : NAND2_X2 port map( A1 => n2383, A2 => n22463, ZN => n32432);
   U11020 : NAND2_X2 port map( A1 => n23919, A2 => n6869, ZN => n5759);
   U11023 : XOR2_X1 port map( A1 => n9474, A2 => n10872, Z => n14845);
   U11025 : NAND2_X2 port map( A1 => n24148, A2 => n24147, ZN => n11346);
   U11028 : NAND2_X2 port map( A1 => n10500, A2 => n23574, ZN => n24148);
   U11032 : XOR2_X1 port map( A1 => n16283, A2 => n32433, Z => n23719);
   U11039 : XOR2_X1 port map( A1 => n23450, A2 => n23062, Z => n32433);
   U11041 : XOR2_X1 port map( A1 => n17504, A2 => n17505, Z => n18075);
   U11042 : AND2_X1 port map( A1 => n5466, A2 => n11571, Z => n14510);
   U11044 : OAI22_X1 port map( A1 => n21412, A2 => n14483, B1 => n13367, B2 => 
                           n11513, ZN => n10135);
   U11045 : XOR2_X1 port map( A1 => n20895, A2 => n14875, Z => n3630);
   U11046 : OR2_X1 port map( A1 => n21085, A2 => n14803, Z => n26988);
   U11048 : NAND2_X2 port map( A1 => n29754, A2 => n34069, ZN => n14359);
   U11052 : NAND2_X2 port map( A1 => n33379, A2 => n10003, ZN => n22798);
   U11056 : OAI21_X2 port map( A1 => n1047, A2 => n18988, B => n5761, ZN => 
                           n10373);
   U11058 : NAND2_X1 port map( A1 => n30643, A2 => n5748, ZN => n20537);
   U11063 : NOR2_X2 port map( A1 => n30031, A2 => n9341, ZN => n30643);
   U11066 : INV_X2 port map( I => n32436, ZN => n24216);
   U11073 : NAND3_X2 port map( A1 => n33431, A2 => n33457, A3 => n14166, ZN => 
                           n32436);
   U11074 : BUF_X2 port map( I => n27921, Z => n32437);
   U11077 : NAND2_X2 port map( A1 => n10046, A2 => n23964, ZN => n24676);
   U11078 : AOI22_X2 port map( A1 => n29293, A2 => n31113, B1 => n10047, B2 => 
                           n10859, ZN => n10046);
   U11079 : AOI22_X2 port map( A1 => n8968, A2 => n24290, B1 => n32985, B2 => 
                           n2444, ZN => n12454);
   U11080 : NAND2_X1 port map( A1 => n12135, A2 => n17501, ZN => n32438);
   U11082 : NAND2_X2 port map( A1 => n25852, A2 => n25851, ZN => n30805);
   U11083 : NOR2_X2 port map( A1 => n10897, A2 => n16673, ZN => n25852);
   U11088 : NAND2_X2 port map( A1 => n32439, A2 => n33396, ZN => n19180);
   U11094 : NAND2_X2 port map( A1 => n11208, A2 => n21797, ZN => n28824);
   U11095 : NOR2_X1 port map( A1 => n33788, A2 => n31916, ZN => n13354);
   U11096 : NOR2_X2 port map( A1 => n14948, A2 => n29721, ZN => n14952);
   U11098 : NOR2_X2 port map( A1 => n32917, A2 => n12356, ZN => n24015);
   U11100 : NAND2_X2 port map( A1 => n21314, A2 => n28565, ZN => n17698);
   U11101 : NOR2_X2 port map( A1 => n32440, A2 => n29560, ZN => n1344);
   U11102 : BUF_X4 port map( I => n14457, Z => n34103);
   U11105 : OAI21_X2 port map( A1 => n32437, A2 => n19111, B => n28996, ZN => 
                           n19629);
   U11106 : NOR3_X2 port map( A1 => n10965, A2 => n18260, A3 => n18370, ZN => 
                           n19360);
   U11107 : NAND2_X2 port map( A1 => n33285, A2 => n1609, ZN => n10087);
   U11110 : NAND2_X2 port map( A1 => n9770, A2 => n32442, ZN => n14123);
   U11113 : XOR2_X1 port map( A1 => n32443, A2 => n31513, Z => Ciphertext(8));
   U11115 : XOR2_X1 port map( A1 => n32445, A2 => n14899, Z => n13716);
   U11125 : XOR2_X1 port map( A1 => n21048, A2 => n5024, Z => n32445);
   U11127 : NOR2_X2 port map( A1 => n32447, A2 => n32446, ZN => n16051);
   U11128 : INV_X2 port map( I => n22429, ZN => n32448);
   U11129 : BUF_X2 port map( I => n22521, Z => n32449);
   U11132 : NAND3_X2 port map( A1 => n30071, A2 => n15544, A3 => n30805, ZN => 
                           n32782);
   U11135 : AOI21_X2 port map( A1 => n32450, A2 => n26173, B => n31001, ZN => 
                           n21929);
   U11136 : BUF_X2 port map( I => n14625, Z => n32451);
   U11138 : OAI21_X2 port map( A1 => n6320, A2 => n6321, B => n28914, ZN => 
                           n32453);
   U11141 : AOI21_X2 port map( A1 => n27625, A2 => n5050, B => n32911, ZN => 
                           n32910);
   U11143 : NAND2_X2 port map( A1 => n18154, A2 => n25019, ZN => n5050);
   U11144 : XOR2_X1 port map( A1 => n19558, A2 => n3131, Z => n17840);
   U11145 : XOR2_X1 port map( A1 => n32458, A2 => n25878, Z => Ciphertext(180))
                           ;
   U11147 : NAND2_X1 port map( A1 => n6047, A2 => n31075, ZN => n32458);
   U11148 : XOR2_X1 port map( A1 => n13471, A2 => n24621, Z => n9467);
   U11150 : XOR2_X1 port map( A1 => n11751, A2 => n3345, Z => n24621);
   U11151 : NAND3_X1 port map( A1 => n1081, A2 => n13428, A3 => n14454, ZN => 
                           n7532);
   U11153 : NAND3_X1 port map( A1 => n10862, A2 => n27390, A3 => n8919, ZN => 
                           n17186);
   U11154 : XOR2_X1 port map( A1 => n22313, A2 => n12980, Z => n21885);
   U11157 : AOI21_X1 port map( A1 => n10653, A2 => n24156, B => n10652, ZN => 
                           n6741);
   U11162 : NOR2_X2 port map( A1 => n12043, A2 => n16240, ZN => n15327);
   U11165 : AOI21_X2 port map( A1 => n5160, A2 => n24093, B => n888, ZN => 
                           n5161);
   U11179 : NOR2_X1 port map( A1 => n16408, A2 => n17601, ZN => n33047);
   U11182 : AOI21_X2 port map( A1 => n9105, A2 => n19814, B => n32460, ZN => 
                           n31533);
   U11184 : NOR2_X1 port map( A1 => n19811, A2 => n19812, ZN => n32460);
   U11190 : XOR2_X1 port map( A1 => n11751, A2 => n16575, Z => n5378);
   U11191 : NAND3_X2 port map( A1 => n27397, A2 => n27396, A3 => n5307, ZN => 
                           n11751);
   U11194 : XNOR2_X1 port map( A1 => n20852, A2 => n20851, ZN => n20930);
   U11196 : AOI22_X2 port map( A1 => n10379, A2 => n20499, B1 => n10992, B2 => 
                           n20497, ZN => n20851);
   U11200 : NOR2_X2 port map( A1 => n11241, A2 => n12991, ZN => n20852);
   U11204 : NAND2_X2 port map( A1 => n29790, A2 => n28035, ZN => n1577);
   U11209 : INV_X4 port map( I => n32461, ZN => n20635);
   U11212 : AND3_X2 port map( A1 => n1812, A2 => n1813, A3 => n1814, Z => 
                           n32461);
   U11214 : NAND4_X2 port map( A1 => n17480, A2 => n17479, A3 => n24353, A4 => 
                           n33343, ZN => n32709);
   U11215 : NAND2_X2 port map( A1 => n32462, A2 => n12237, ZN => n13334);
   U11216 : NAND2_X2 port map( A1 => n32463, A2 => n18142, ZN => n30090);
   U11219 : OAI22_X2 port map( A1 => n1362, A2 => n11911, B1 => n1458, B2 => 
                           n397, ZN => n32463);
   U11223 : XOR2_X1 port map( A1 => n31221, A2 => n22104, Z => n29740);
   U11228 : NAND2_X2 port map( A1 => n17124, A2 => n17122, ZN => n22791);
   U11229 : NOR2_X1 port map( A1 => n26013, A2 => n32778, ZN => n29547);
   U11234 : XOR2_X1 port map( A1 => n13395, A2 => n10628, Z => n32464);
   U11237 : XOR2_X1 port map( A1 => n19578, A2 => n19556, Z => n5768);
   U11239 : BUF_X2 port map( I => n3148, Z => n32465);
   U11241 : NOR2_X1 port map( A1 => n21806, A2 => n21805, ZN => n33985);
   U11243 : NAND2_X2 port map( A1 => n1837, A2 => n1838, ZN => n8636);
   U11246 : NAND2_X2 port map( A1 => n32546, A2 => n337, ZN => n16708);
   U11247 : NAND3_X2 port map( A1 => n32466, A2 => n9232, A3 => n330, ZN => 
                           n33140);
   U11249 : NAND2_X2 port map( A1 => n15394, A2 => n26130, ZN => n32466);
   U11254 : XOR2_X1 port map( A1 => n16448, A2 => n20990, Z => n34038);
   U11256 : NOR2_X2 port map( A1 => n5059, A2 => n5061, ZN => n16448);
   U11258 : NOR2_X2 port map( A1 => n31220, A2 => n29084, ZN => n27535);
   U11259 : NAND2_X2 port map( A1 => n1508, A2 => n32468, ZN => n24810);
   U11261 : AOI22_X2 port map( A1 => n32049, A2 => n24251, B1 => n1511, B2 => 
                           n1513, ZN => n32468);
   U11264 : OAI21_X1 port map( A1 => n787, A2 => n5713, B => n25106, ZN => 
                           n18175);
   U11265 : INV_X2 port map( I => n11360, ZN => n787);
   U11266 : NAND2_X2 port map( A1 => n3223, A2 => n3225, ZN => n11360);
   U11269 : OAI21_X2 port map( A1 => n10645, A2 => n10646, B => n7181, ZN => 
                           n10329);
   U11271 : NAND3_X1 port map( A1 => n8030, A2 => n16925, A3 => n16157, ZN => 
                           n7324);
   U11277 : OR2_X1 port map( A1 => n17637, A2 => n6595, Z => n30523);
   U11278 : INV_X2 port map( I => n1026, ZN => n33631);
   U11286 : NOR2_X2 port map( A1 => n11187, A2 => n1145, ZN => n11091);
   U11287 : INV_X2 port map( I => n10433, ZN => n1145);
   U11289 : AND2_X1 port map( A1 => n21604, A2 => n26439, Z => n34028);
   U11290 : XOR2_X1 port map( A1 => n31493, A2 => n22075, Z => n16150);
   U11291 : XOR2_X1 port map( A1 => n22105, A2 => n27633, Z => n31649);
   U11292 : XOR2_X1 port map( A1 => n17362, A2 => n22012, Z => n22105);
   U11297 : XOR2_X1 port map( A1 => n6771, A2 => n28762, Z => n33203);
   U11304 : OAI21_X2 port map( A1 => n34026, A2 => n21656, B => n32535, ZN => 
                           n28762);
   U11309 : XOR2_X1 port map( A1 => n24618, A2 => n24393, Z => n24504);
   U11314 : NOR2_X2 port map( A1 => n28505, A2 => n12262, ZN => n24618);
   U11315 : OAI22_X2 port map( A1 => n28367, A2 => n10213, B1 => n23873, B2 => 
                           n17133, ZN => n3571);
   U11318 : INV_X1 port map( I => n33996, ZN => n22741);
   U11320 : NAND2_X1 port map( A1 => n22848, A2 => n31854, ZN => n33996);
   U11321 : XOR2_X1 port map( A1 => n30029, A2 => n32469, Z => n24565);
   U11323 : XOR2_X1 port map( A1 => n9011, A2 => n9012, Z => n9010);
   U11324 : NOR2_X2 port map( A1 => n5741, A2 => n29306, ZN => n6769);
   U11325 : INV_X1 port map( I => n18100, ZN => n14593);
   U11326 : XNOR2_X1 port map( A1 => n22137, A2 => n22158, ZN => n18100);
   U11330 : XOR2_X1 port map( A1 => n19565, A2 => n14146, Z => n19429);
   U11331 : OR2_X2 port map( A1 => n499, A2 => n33461, Z => n17579);
   U11332 : NOR2_X2 port map( A1 => n22563, A2 => n14034, ZN => n32654);
   U11333 : NAND2_X2 port map( A1 => n16447, A2 => n15089, ZN => n22563);
   U11334 : XOR2_X1 port map( A1 => n30380, A2 => n23488, Z => n28587);
   U11336 : NOR2_X1 port map( A1 => n15234, A2 => n3080, ZN => n32471);
   U11338 : INV_X2 port map( I => n25444, ZN => n25455);
   U11339 : NAND2_X2 port map( A1 => n33245, A2 => n33258, ZN => n25444);
   U11345 : NOR2_X2 port map( A1 => n32472, A2 => n9725, ZN => n32648);
   U11351 : AOI21_X2 port map( A1 => n19826, A2 => n19827, B => n29972, ZN => 
                           n32472);
   U11353 : INV_X4 port map( I => n32635, ZN => n11956);
   U11354 : INV_X2 port map( I => n18039, ZN => n20097);
   U11355 : XOR2_X1 port map( A1 => n17954, A2 => n17953, Z => n18039);
   U11357 : AOI22_X2 port map( A1 => n5080, A2 => n29985, B1 => n5079, B2 => 
                           n1232, ZN => n30327);
   U11359 : AND3_X1 port map( A1 => n11298, A2 => n14420, A3 => n4184, Z => 
                           n33834);
   U11361 : NAND2_X2 port map( A1 => n11823, A2 => n11824, ZN => n30047);
   U11362 : XOR2_X1 port map( A1 => n20716, A2 => n32473, Z => n7918);
   U11366 : XOR2_X1 port map( A1 => n7594, A2 => n20552, Z => n32473);
   U11369 : XOR2_X1 port map( A1 => n26920, A2 => n28134, Z => n16275);
   U11376 : XOR2_X1 port map( A1 => n61, A2 => n32474, Z => n25963);
   U11383 : XOR2_X1 port map( A1 => n21985, A2 => n15950, Z => n32474);
   U11385 : XOR2_X1 port map( A1 => n4583, A2 => n29458, Z => n4581);
   U11390 : XOR2_X1 port map( A1 => n5090, A2 => n24116, Z => n24793);
   U11393 : NOR2_X2 port map( A1 => n10531, A2 => n12002, ZN => n5090);
   U11403 : XOR2_X1 port map( A1 => n10235, A2 => n24685, Z => n27290);
   U11417 : XOR2_X1 port map( A1 => n24750, A2 => n5090, Z => n24685);
   U11422 : INV_X2 port map( I => n14585, ZN => n16615);
   U11425 : XOR2_X1 port map( A1 => n14580, A2 => n14581, Z => n14585);
   U11431 : NAND4_X2 port map( A1 => n32475, A2 => n22857, A3 => n22859, A4 => 
                           n22860, ZN => n23336);
   U11434 : NAND2_X2 port map( A1 => n7797, A2 => n26667, ZN => n32475);
   U11439 : AND2_X1 port map( A1 => n20097, A2 => n20096, Z => n7997);
   U11441 : AND2_X1 port map( A1 => n25797, A2 => n16112, Z => n14615);
   U11443 : NAND2_X2 port map( A1 => n32476, A2 => n23479, ZN => n29885);
   U11444 : OAI21_X2 port map( A1 => n30825, A2 => n8415, B => n33016, ZN => 
                           n32476);
   U11446 : NOR2_X1 port map( A1 => n28200, A2 => n15323, ZN => n25129);
   U11448 : NAND3_X2 port map( A1 => n14628, A2 => n14631, A3 => n14632, ZN => 
                           n15323);
   U11453 : BUF_X2 port map( I => n13092, Z => n32478);
   U11461 : NOR2_X2 port map( A1 => n30832, A2 => n7811, ZN => n5385);
   U11468 : OAI22_X2 port map( A1 => n21196, A2 => n21195, B1 => n26542, B2 => 
                           n17624, ZN => n30832);
   U11473 : OAI21_X2 port map( A1 => n32479, A2 => n4855, B => n33148, ZN => 
                           n14106);
   U11474 : NAND2_X2 port map( A1 => n2937, A2 => n8308, ZN => n23511);
   U11475 : NAND2_X2 port map( A1 => n33656, A2 => n2912, ZN => n2937);
   U11477 : NAND2_X2 port map( A1 => n11179, A2 => n19008, ZN => n11219);
   U11480 : NAND2_X2 port map( A1 => n32534, A2 => n27368, ZN => n3007);
   U11487 : XOR2_X1 port map( A1 => n32480, A2 => n23295, Z => n81);
   U11491 : NAND2_X2 port map( A1 => n33184, A2 => n2539, ZN => n27396);
   U11493 : NAND3_X2 port map( A1 => n983, A2 => n12259, A3 => n11268, ZN => 
                           n11109);
   U11496 : XOR2_X1 port map( A1 => n22169, A2 => n22168, Z => n2162);
   U11497 : XOR2_X1 port map( A1 => n1309, A2 => n16242, Z => n22169);
   U11498 : INV_X2 port map( I => n4013, ZN => n22132);
   U11499 : NAND2_X2 port map( A1 => n3314, A2 => n3316, ZN => n4013);
   U11500 : NAND2_X1 port map( A1 => n33937, A2 => n28085, ZN => n12808);
   U11505 : XOR2_X1 port map( A1 => n7545, A2 => n22271, Z => n22104);
   U11508 : NOR2_X2 port map( A1 => n17418, A2 => n21347, ZN => n22271);
   U11510 : NAND2_X2 port map( A1 => n26375, A2 => n32482, ZN => n17855);
   U11514 : NAND2_X1 port map( A1 => n23708, A2 => n12680, ZN => n15942);
   U11515 : AOI22_X2 port map( A1 => n28428, A2 => n24134, B1 => n24135, B2 => 
                           n27739, ZN => n27998);
   U11526 : XOR2_X1 port map( A1 => n20918, A2 => n20834, Z => n4949);
   U11527 : XOR2_X1 port map( A1 => n20960, A2 => n1339, Z => n20918);
   U11528 : AOI21_X2 port map( A1 => n27150, A2 => n24925, B => n24920, ZN => 
                           n4867);
   U11529 : INV_X2 port map( I => n24936, ZN => n24920);
   U11531 : NAND2_X2 port map( A1 => n16216, A2 => n16217, ZN => n13573);
   U11532 : INV_X2 port map( I => n6531, ZN => n12263);
   U11533 : AOI22_X2 port map( A1 => n19924, A2 => n26615, B1 => n8934, B2 => 
                           n33187, ZN => n6531);
   U11545 : INV_X2 port map( I => n14737, ZN => n963);
   U11546 : NOR2_X1 port map( A1 => n8535, A2 => n10993, ZN => n32494);
   U11548 : AND2_X1 port map( A1 => n29203, A2 => n23578, Z => n12326);
   U11549 : NOR2_X2 port map( A1 => n13966, A2 => n13965, ZN => n27066);
   U11551 : INV_X2 port map( I => n32484, ZN => n29250);
   U11555 : XNOR2_X1 port map( A1 => n4014, A2 => n4895, ZN => n32484);
   U11558 : NAND3_X1 port map( A1 => n26830, A2 => n13295, A3 => n13390, ZN => 
                           n12114);
   U11559 : NOR2_X2 port map( A1 => n9377, A2 => n23018, ZN => n22473);
   U11567 : NAND2_X1 port map( A1 => n28, A2 => n9793, ZN => n9792);
   U11572 : NAND2_X2 port map( A1 => n32978, A2 => n15925, ZN => n9793);
   U11577 : NAND2_X1 port map( A1 => n1207, A2 => n25277, ZN => n27873);
   U11579 : NAND2_X2 port map( A1 => n22277, A2 => n7, ZN => n11033);
   U11582 : OAI22_X2 port map( A1 => n22411, A2 => n7023, B1 => n645, B2 => 
                           n16225, ZN => n22277);
   U11584 : INV_X2 port map( I => n32486, ZN => n31448);
   U11587 : XNOR2_X1 port map( A1 => n2952, A2 => n2951, ZN => n32486);
   U11588 : NAND2_X2 port map( A1 => n32528, A2 => n20134, ZN => n31157);
   U11590 : INV_X2 port map( I => n32487, ZN => n8028);
   U11591 : XNOR2_X1 port map( A1 => n8026, A2 => n27091, ZN => n32487);
   U11600 : AOI22_X2 port map( A1 => n97, A2 => n98, B1 => n29708, B2 => n32488
                           , ZN => n18146);
   U11604 : NAND2_X2 port map( A1 => n23823, A2 => n23672, ZN => n32488);
   U11606 : XOR2_X1 port map( A1 => n12539, A2 => n14875, Z => n15353);
   U11607 : XOR2_X1 port map( A1 => n32489, A2 => n647, Z => n2200);
   U11608 : NAND2_X2 port map( A1 => n32490, A2 => n29107, ZN => n4542);
   U11610 : OAI22_X2 port map( A1 => n23055, A2 => n17739, B1 => n22878, B2 => 
                           n31437, ZN => n32490);
   U11619 : NAND2_X1 port map( A1 => n29692, A2 => n10623, ZN => n10369);
   U11621 : NOR2_X2 port map( A1 => n32491, A2 => n12768, ZN => n31746);
   U11623 : OAI21_X2 port map( A1 => n12150, A2 => n20412, B => n12149, ZN => 
                           n30219);
   U11624 : XOR2_X1 port map( A1 => n22285, A2 => n32492, Z => n13382);
   U11627 : XOR2_X1 port map( A1 => n2824, A2 => n5099, Z => n32492);
   U11631 : AOI22_X2 port map( A1 => n20308, A2 => n3462, B1 => n2145, B2 => 
                           n33691, ZN => n20309);
   U11633 : BUF_X2 port map( I => n907, Z => n32493);
   U11635 : XOR2_X1 port map( A1 => n33160, A2 => n30495, Z => n10482);
   U11636 : NOR2_X2 port map( A1 => n33409, A2 => n13804, ZN => n30495);
   U11639 : INV_X2 port map( I => n15064, ZN => n19634);
   U11647 : OAI21_X2 port map( A1 => n2411, A2 => n2412, B => n2410, ZN => 
                           n15064);
   U11648 : NAND2_X2 port map( A1 => n19220, A2 => n5610, ZN => n14760);
   U11650 : NAND2_X2 port map( A1 => n18371, A2 => n18372, ZN => n19220);
   U11652 : XOR2_X1 port map( A1 => n4246, A2 => n5732, Z => n9351);
   U11654 : XOR2_X1 port map( A1 => n15161, A2 => n2117, Z => n24674);
   U11655 : AOI21_X2 port map( A1 => n24066, A2 => n14745, B => n3918, ZN => 
                           n15161);
   U11656 : XOR2_X1 port map( A1 => n8328, A2 => n10888, Z => n11620);
   U11658 : INV_X2 port map( I => n8306, ZN => n30528);
   U11659 : NAND2_X2 port map( A1 => n10510, A2 => n10511, ZN => n8306);
   U11660 : AOI22_X2 port map( A1 => n12987, A2 => n20059, B1 => n20058, B2 => 
                           n941, ZN => n12986);
   U11665 : XOR2_X1 port map( A1 => n11358, A2 => n11355, Z => n16885);
   U11666 : NOR3_X2 port map( A1 => n33911, A2 => n33919, A3 => n25295, ZN => 
                           n11258);
   U11667 : NAND2_X2 port map( A1 => n13197, A2 => n7957, ZN => n22921);
   U11669 : NAND2_X2 port map( A1 => n12869, A2 => n17853, ZN => n13197);
   U11670 : NAND3_X2 port map( A1 => n11584, A2 => n32495, A3 => n21667, ZN => 
                           n22125);
   U11671 : OAI21_X2 port map( A1 => n26175, A2 => n4842, B => n28618, ZN => 
                           n32495);
   U11679 : BUF_X2 port map( I => n15172, Z => n13133);
   U11682 : NOR2_X1 port map( A1 => n34012, A2 => n34011, ZN => n3336);
   U11683 : NAND3_X2 port map( A1 => n810, A2 => n21080, A3 => n21365, ZN => 
                           n33551);
   U11685 : OAI22_X2 port map( A1 => n32496, A2 => n30510, B1 => n6482, B2 => 
                           n7090, ZN => n22974);
   U11686 : AOI21_X2 port map( A1 => n32498, A2 => n32497, B => n29595, ZN => 
                           n3634);
   U11688 : NOR2_X2 port map( A1 => n32588, A2 => n32499, ZN => n32498);
   U11691 : XOR2_X1 port map( A1 => n22085, A2 => n22173, Z => n17207);
   U11696 : XOR2_X1 port map( A1 => n32501, A2 => n29420, Z => n4820);
   U11699 : XOR2_X1 port map( A1 => n1865, A2 => n26646, Z => n32501);
   U11701 : NAND2_X2 port map( A1 => n789, A2 => n29331, ZN => n5839);
   U11702 : XOR2_X1 port map( A1 => n16617, A2 => n16618, Z => n8452);
   U11703 : XOR2_X1 port map( A1 => n2969, A2 => n2968, Z => n3012);
   U11705 : NOR2_X2 port map( A1 => n17590, A2 => n17305, ZN => n21162);
   U11706 : XOR2_X1 port map( A1 => n20786, A2 => n20960, Z => n20688);
   U11710 : NOR2_X2 port map( A1 => n14394, A2 => n8264, ZN => n20786);
   U11716 : XOR2_X1 port map( A1 => n32502, A2 => n3793, Z => n33538);
   U11719 : XOR2_X1 port map( A1 => n5356, A2 => n32077, Z => n33934);
   U11726 : NAND2_X1 port map( A1 => n32503, A2 => n14433, ZN => n33873);
   U11729 : NAND2_X1 port map( A1 => n27659, A2 => n14432, ZN => n32503);
   U11734 : INV_X2 port map( I => n32507, ZN => n24603);
   U11736 : XOR2_X1 port map( A1 => n5790, A2 => n24652, Z => n32507);
   U11750 : OAI21_X2 port map( A1 => n2640, A2 => n737, B => n7891, ZN => 
                           n33019);
   U11751 : XOR2_X1 port map( A1 => n32508, A2 => n12754, Z => Ciphertext(155))
                           ;
   U11757 : NAND2_X2 port map( A1 => n28526, A2 => n16934, ZN => n28203);
   U11759 : NAND2_X2 port map( A1 => n3163, A2 => n724, ZN => n28831);
   U11760 : AOI21_X2 port map( A1 => n26688, A2 => n32509, B => n8876, ZN => 
                           n31434);
   U11761 : XOR2_X1 port map( A1 => n20895, A2 => n10581, Z => n32511);
   U11764 : NAND3_X1 port map( A1 => n30945, A2 => n30946, A3 => n23082, ZN => 
                           n33777);
   U11766 : BUF_X2 port map( I => n32605, Z => n32512);
   U11771 : NAND3_X2 port map( A1 => n11814, A2 => n21358, A3 => n21357, ZN => 
                           n33297);
   U11772 : NAND2_X2 port map( A1 => n32514, A2 => n30084, ZN => n2045);
   U11773 : AOI22_X2 port map( A1 => n1634, A2 => n24233, B1 => n5066, B2 => 
                           n974, ZN => n32514);
   U11775 : XOR2_X1 port map( A1 => n32517, A2 => n25358, Z => Ciphertext(98));
   U11776 : NAND2_X1 port map( A1 => n28469, A2 => n28470, ZN => n32517);
   U11779 : OR2_X1 port map( A1 => n13147, A2 => n13180, Z => n11061);
   U11782 : NAND2_X2 port map( A1 => n12452, A2 => n17098, ZN => n21671);
   U11785 : NAND2_X2 port map( A1 => n16851, A2 => n26468, ZN => n12452);
   U11787 : XOR2_X1 port map( A1 => n23371, A2 => n25040, Z => n7411);
   U11789 : XOR2_X1 port map( A1 => n22229, A2 => n8282, Z => n5356);
   U11790 : OR2_X1 port map( A1 => n33934, A2 => n33082, Z => n22430);
   U11793 : NAND2_X2 port map( A1 => n7144, A2 => n8602, ZN => n32519);
   U11794 : NAND2_X1 port map( A1 => n8926, A2 => n25176, ZN => n11468);
   U11798 : NAND2_X2 port map( A1 => n33620, A2 => n11111, ZN => n8926);
   U11803 : XOR2_X1 port map( A1 => n24358, A2 => n16416, Z => n24719);
   U11806 : NAND2_X2 port map( A1 => n14642, A2 => n17053, ZN => n10261);
   U11808 : AND2_X1 port map( A1 => n32926, A2 => n4862, Z => n7429);
   U11809 : XOR2_X1 port map( A1 => n22186, A2 => n9369, Z => n5796);
   U11813 : XOR2_X1 port map( A1 => n14639, A2 => n22080, Z => n22186);
   U11816 : AOI22_X2 port map( A1 => n32088, A2 => n33787, B1 => n7857, B2 => 
                           n28649, ZN => n3170);
   U11823 : NOR2_X2 port map( A1 => n33132, A2 => n25979, ZN => n7857);
   U11829 : NAND2_X2 port map( A1 => n32521, A2 => n17079, ZN => n14640);
   U11830 : NAND2_X2 port map( A1 => n33286, A2 => n9691, ZN => n32881);
   U11832 : NAND3_X2 port map( A1 => n11657, A2 => n14829, A3 => n11656, ZN => 
                           n27130);
   U11834 : NOR2_X2 port map( A1 => n11659, A2 => n11658, ZN => n11657);
   U11838 : AOI21_X2 port map( A1 => n5619, A2 => n5055, B => n5054, ZN => 
                           n12652);
   U11839 : OAI22_X2 port map( A1 => n5618, A2 => n13597, B1 => n22886, B2 => 
                           n12511, ZN => n5054);
   U11842 : XOR2_X1 port map( A1 => n23261, A2 => n23237, Z => n12573);
   U11843 : XOR2_X1 port map( A1 => n7229, A2 => n23120, Z => n23261);
   U11844 : NOR2_X2 port map( A1 => n25446, A2 => n25444, ZN => n25433);
   U11845 : NOR2_X2 port map( A1 => n25058, A2 => n25062, ZN => n17729);
   U11854 : NOR2_X2 port map( A1 => n32523, A2 => n7649, ZN => n6322);
   U11857 : NOR2_X1 port map( A1 => n22596, A2 => n7633, ZN => n32523);
   U11859 : INV_X2 port map( I => n10924, ZN => n887);
   U11861 : NAND2_X2 port map( A1 => n2153, A2 => n2154, ZN => n10924);
   U11864 : XOR2_X1 port map( A1 => n32524, A2 => n25436, Z => Ciphertext(105))
                           ;
   U11873 : NAND2_X1 port map( A1 => n25434, A2 => n33159, ZN => n32524);
   U11877 : NOR2_X2 port map( A1 => n29392, A2 => n32525, ZN => n6400);
   U11879 : XOR2_X1 port map( A1 => n33333, A2 => n22779, Z => n11568);
   U11886 : XOR2_X1 port map( A1 => n4047, A2 => n11668, Z => n22779);
   U11887 : OAI21_X2 port map( A1 => n33963, A2 => n32526, B => n23699, ZN => 
                           n5051);
   U11890 : AOI21_X2 port map( A1 => n2949, A2 => n21771, B => n2948, ZN => 
                           n22173);
   U11892 : OAI22_X2 port map( A1 => n1015, A2 => n38, B1 => n2368, B2 => 
                           n33766, ZN => n21771);
   U11893 : XOR2_X1 port map( A1 => n32527, A2 => n25728, Z => Ciphertext(154))
                           ;
   U11894 : NAND4_X2 port map( A1 => n25727, A2 => n25726, A3 => n34019, A4 => 
                           n25725, ZN => n32527);
   U11896 : NAND2_X2 port map( A1 => n31921, A2 => n13532, ZN => n25593);
   U11897 : XOR2_X1 port map( A1 => n27613, A2 => n1102, Z => n23501);
   U11901 : NAND2_X2 port map( A1 => n7217, A2 => n7724, ZN => n27613);
   U11905 : XOR2_X1 port map( A1 => n14058, A2 => n24819, Z => n16838);
   U11912 : XOR2_X1 port map( A1 => n32529, A2 => n25091, Z => Ciphertext(49));
   U11913 : NOR3_X1 port map( A1 => n16226, A2 => n16933, A3 => n4518, ZN => 
                           n33167);
   U11919 : BUF_X2 port map( I => n18254, Z => n32530);
   U11926 : BUF_X2 port map( I => n22945, Z => n32531);
   U11928 : NOR2_X2 port map( A1 => n11259, A2 => n11258, ZN => n32933);
   U11938 : BUF_X2 port map( I => n34161, Z => n32532);
   U11941 : INV_X1 port map( I => n19167, ZN => n33845);
   U11946 : AOI22_X2 port map( A1 => n22839, A2 => n29329, B1 => n22840, B2 => 
                           n8990, ZN => n33001);
   U11955 : OAI21_X1 port map( A1 => n8923, A2 => n9954, B => n32710, ZN => 
                           n10495);
   U11958 : AOI22_X2 port map( A1 => n17286, A2 => n23786, B1 => n17157, B2 => 
                           n15692, ZN => n841);
   U11960 : NAND2_X2 port map( A1 => n4110, A2 => n22832, ZN => n17503);
   U11971 : NAND2_X2 port map( A1 => n3520, A2 => n29349, ZN => n4110);
   U11974 : XOR2_X1 port map( A1 => n23533, A2 => n23529, Z => n32841);
   U11976 : NAND2_X2 port map( A1 => n4651, A2 => n4650, ZN => n23529);
   U11980 : XOR2_X1 port map( A1 => n32533, A2 => n24399, Z => n34030);
   U11982 : XOR2_X1 port map( A1 => n7574, A2 => n12493, Z => n24399);
   U11983 : INV_X2 port map( I => n15588, ZN => n32533);
   U11985 : NOR2_X2 port map( A1 => n33132, A2 => n30365, ZN => n7797);
   U11987 : NAND3_X2 port map( A1 => n17773, A2 => n27024, A3 => n15655, ZN => 
                           n21276);
   U11989 : NOR3_X2 port map( A1 => n2657, A2 => n2656, A3 => n13143, ZN => 
                           n32534);
   U11992 : NOR2_X1 port map( A1 => n25784, A2 => n33720, ZN => n25779);
   U11994 : NAND2_X1 port map( A1 => n25779, A2 => n25790, ZN => n25780);
   U12002 : NAND4_X2 port map( A1 => n4899, A2 => n3820, A3 => n24365, A4 => 
                           n4898, ZN => n32977);
   U12003 : NAND2_X2 port map( A1 => n32536, A2 => n31531, ZN => n32842);
   U12006 : NAND2_X2 port map( A1 => n29329, A2 => n22978, ZN => n32536);
   U12008 : XNOR2_X1 port map( A1 => n21020, A2 => n20782, ZN => n20168);
   U12012 : XOR2_X1 port map( A1 => n20720, A2 => n10949, Z => n20782);
   U12013 : INV_X2 port map( I => n7, ZN => n630);
   U12014 : NOR2_X2 port map( A1 => n75, A2 => n12929, ZN => n9500);
   U12016 : AOI22_X2 port map( A1 => n32658, A2 => n28314, B1 => n12728, B2 => 
                           n12727, ZN => n30433);
   U12022 : AOI21_X2 port map( A1 => n4375, A2 => n18204, B => n4374, ZN => 
                           n7188);
   U12028 : NAND2_X2 port map( A1 => n25486, A2 => n25462, ZN => n25482);
   U12030 : OR2_X1 port map( A1 => n24335, A2 => n24242, Z => n33669);
   U12031 : AOI21_X2 port map( A1 => n22633, A2 => n11932, B => n32512, ZN => 
                           n7179);
   U12046 : INV_X2 port map( I => n32538, ZN => n22633);
   U12048 : NOR2_X2 port map( A1 => n522, A2 => n17916, ZN => n32538);
   U12049 : NOR2_X1 port map( A1 => n15882, A2 => n31994, ZN => n32717);
   U12054 : NOR2_X2 port map( A1 => n33533, A2 => n29830, ZN => n646);
   U12061 : INV_X2 port map( I => n32539, ZN => n10569);
   U12062 : XOR2_X1 port map( A1 => n2210, A2 => n2211, Z => n32539);
   U12063 : NOR2_X1 port map( A1 => n22785, A2 => n30584, ZN => n29384);
   U12066 : XOR2_X1 port map( A1 => n3368, A2 => n32540, Z => n22199);
   U12068 : XOR2_X1 port map( A1 => n22186, A2 => n28005, Z => n32540);
   U12071 : XOR2_X1 port map( A1 => n23361, A2 => n32633, Z => n29906);
   U12072 : XOR2_X1 port map( A1 => n13216, A2 => n13814, Z => n23361);
   U12073 : NAND2_X2 port map( A1 => n32541, A2 => n2508, ZN => n26969);
   U12074 : NOR2_X2 port map( A1 => n16280, A2 => n7463, ZN => n6190);
   U12076 : NAND2_X1 port map( A1 => n4097, A2 => n28099, ZN => n13828);
   U12078 : NAND2_X2 port map( A1 => n26679, A2 => n34083, ZN => n4097);
   U12079 : NOR2_X2 port map( A1 => n32598, A2 => n32542, ZN => n22249);
   U12080 : AOI21_X2 port map( A1 => n21863, A2 => n21862, B => n1016, ZN => 
                           n32542);
   U12083 : NAND2_X2 port map( A1 => n30649, A2 => n3840, ZN => n11438);
   U12088 : NAND2_X2 port map( A1 => n30448, A2 => n33026, ZN => n9546);
   U12091 : XOR2_X1 port map( A1 => n32543, A2 => n20668, Z => n2881);
   U12102 : XOR2_X1 port map( A1 => n2883, A2 => n31233, Z => n32543);
   U12103 : XOR2_X1 port map( A1 => n12652, A2 => n23200, Z => n23343);
   U12106 : OR2_X1 port map( A1 => n21395, A2 => n6681, Z => n16058);
   U12110 : INV_X2 port map( I => n4862, ZN => n32605);
   U12112 : OAI21_X2 port map( A1 => n21414, A2 => n21413, B => n1332, ZN => 
                           n9905);
   U12116 : NOR2_X2 port map( A1 => n29143, A2 => n28700, ZN => n4287);
   U12119 : AOI22_X2 port map( A1 => n32544, A2 => n21269, B1 => n28642, B2 => 
                           n29460, ZN => n4082);
   U12124 : NOR2_X2 port map( A1 => n28642, A2 => n21267, ZN => n32544);
   U12126 : AND2_X2 port map( A1 => n25198, A2 => n11985, Z => n26015);
   U12127 : NAND2_X2 port map( A1 => n32545, A2 => n7754, ZN => n7753);
   U12131 : NAND2_X1 port map( A1 => n27245, A2 => n27246, ZN => n32545);
   U12133 : BUF_X4 port map( I => n22487, Z => n33046);
   U12134 : NAND2_X2 port map( A1 => n12443, A2 => n14617, ZN => n23295);
   U12137 : NOR2_X1 port map( A1 => n22592, A2 => n17408, ZN => n17212);
   U12139 : AOI21_X2 port map( A1 => n11246, A2 => n28131, B => n26925, ZN => 
                           n22592);
   U12145 : AOI22_X2 port map( A1 => n28128, A2 => n9854, B1 => n20550, B2 => 
                           n125, ZN => n32546);
   U12146 : AND2_X1 port map( A1 => n4281, A2 => n18204, Z => n7263);
   U12148 : AOI21_X2 port map( A1 => n30219, A2 => n20955, B => n2301, ZN => 
                           n21020);
   U12152 : NAND2_X2 port map( A1 => n32957, A2 => n34128, ZN => n21188);
   U12157 : AOI21_X2 port map( A1 => n1257, A2 => n844, B => n23867, ZN => 
                           n32547);
   U12160 : XOR2_X1 port map( A1 => n28747, A2 => n32548, Z => n7624);
   U12161 : XOR2_X1 port map( A1 => n10869, A2 => n7450, Z => n32548);
   U12167 : NOR2_X2 port map( A1 => n21334, A2 => n32549, ZN => n17416);
   U12171 : AOI21_X2 port map( A1 => n21332, A2 => n21331, B => n8378, ZN => 
                           n32549);
   U12173 : XOR2_X1 port map( A1 => n20904, A2 => n20754, Z => n21034);
   U12181 : NAND2_X2 port map( A1 => n162, A2 => n26478, ZN => n20904);
   U12183 : NAND2_X2 port map( A1 => n14805, A2 => n29278, ZN => n12440);
   U12184 : XOR2_X1 port map( A1 => n34160, A2 => n22098, Z => n22229);
   U12188 : INV_X2 port map( I => n24810, ZN => n9209);
   U12200 : XOR2_X1 port map( A1 => n8754, A2 => n32554, Z => n19899);
   U12201 : XOR2_X1 port map( A1 => n7589, A2 => n7590, Z => n32554);
   U12202 : OAI21_X1 port map( A1 => n19322, A2 => n30894, B => n19068, ZN => 
                           n3132);
   U12205 : NAND2_X1 port map( A1 => n21706, A2 => n15414, ZN => n21754);
   U12207 : NAND3_X2 port map( A1 => n15435, A2 => n15436, A3 => n32555, ZN => 
                           n20305);
   U12209 : NAND2_X2 port map( A1 => n29281, A2 => n19998, ZN => n32555);
   U12210 : XOR2_X1 port map( A1 => n22153, A2 => n22190, Z => n5013);
   U12213 : NOR2_X2 port map( A1 => n31940, A2 => n32556, ZN => n33349);
   U12214 : XOR2_X1 port map( A1 => n9914, A2 => n22161, Z => n1938);
   U12229 : XOR2_X1 port map( A1 => n8291, A2 => n3723, Z => n22161);
   U12231 : XOR2_X1 port map( A1 => n24602, A2 => n32557, Z => n30220);
   U12234 : XOR2_X1 port map( A1 => n15264, A2 => n4997, Z => n32557);
   U12236 : OAI22_X2 port map( A1 => n29630, A2 => n29629, B1 => n4886, B2 => 
                           n4885, ZN => n12257);
   U12261 : INV_X2 port map( I => n11173, ZN => n4885);
   U12264 : XOR2_X1 port map( A1 => n10473, A2 => n10475, Z => n11173);
   U12267 : XOR2_X1 port map( A1 => n5253, A2 => n32558, Z => n8939);
   U12290 : XNOR2_X1 port map( A1 => n27114, A2 => n24522, ZN => n5253);
   U12291 : INV_X2 port map( I => n24746, ZN => n32558);
   U12297 : XOR2_X1 port map( A1 => n14058, A2 => n25801, Z => n13520);
   U12298 : OR2_X1 port map( A1 => n10496, A2 => n22945, Z => n32710);
   U12302 : AOI21_X2 port map( A1 => n32560, A2 => n15718, B => n22916, ZN => 
                           n31399);
   U12309 : XOR2_X1 port map( A1 => n5658, A2 => n10989, Z => n5657);
   U12312 : AOI21_X2 port map( A1 => n17860, A2 => n24029, B => n32561, ZN => 
                           n24847);
   U12316 : NOR3_X2 port map( A1 => n28590, A2 => n9066, A3 => n4118, ZN => 
                           n32561);
   U12318 : XOR2_X1 port map( A1 => n32562, A2 => n31098, Z => n26515);
   U12319 : XOR2_X1 port map( A1 => n23459, A2 => n2862, Z => n32562);
   U12325 : AOI21_X2 port map( A1 => n31469, A2 => n31471, B => n111, ZN => 
                           n12991);
   U12327 : XOR2_X1 port map( A1 => n32563, A2 => n17865, Z => n31639);
   U12328 : XOR2_X1 port map( A1 => n34088, A2 => n2278, Z => n32563);
   U12331 : XOR2_X1 port map( A1 => n14058, A2 => n24853, Z => n24854);
   U12333 : NOR2_X2 port map( A1 => n24238, A2 => n24239, ZN => n24853);
   U12335 : INV_X2 port map( I => n23186, ZN => n982);
   U12342 : OAI22_X2 port map( A1 => n17083, A2 => n17639, B1 => n17085, B2 => 
                           n22884, ZN => n23186);
   U12345 : XOR2_X1 port map( A1 => n33606, A2 => n5215, Z => n8251);
   U12347 : NAND2_X2 port map( A1 => n14542, A2 => n32515, ZN => n4458);
   U12351 : OAI22_X2 port map( A1 => n21554, A2 => n32613, B1 => n21555, B2 => 
                           n21556, ZN => n28413);
   U12353 : BUF_X2 port map( I => n22306, Z => n32564);
   U12354 : NAND2_X2 port map( A1 => n974, A2 => n33832, ZN => n24235);
   U12358 : INV_X2 port map( I => n18665, ZN => n2509);
   U12360 : NAND2_X2 port map( A1 => n31972, A2 => n31971, ZN => n18665);
   U12363 : XOR2_X1 port map( A1 => n32566, A2 => n26001, Z => Ciphertext(45));
   U12367 : XOR2_X1 port map( A1 => n12621, A2 => n12624, Z => n30038);
   U12369 : XOR2_X1 port map( A1 => n32567, A2 => n25040, Z => Ciphertext(38));
   U12371 : NAND2_X1 port map( A1 => n6424, A2 => n33145, ZN => n32567);
   U12373 : OAI21_X2 port map( A1 => n32569, A2 => n32568, B => n32483, ZN => 
                           n17001);
   U12374 : NAND2_X2 port map( A1 => n33585, A2 => n32571, ZN => n32570);
   U12375 : INV_X2 port map( I => n28338, ZN => n32571);
   U12377 : XOR2_X1 port map( A1 => n14969, A2 => n32572, Z => n32838);
   U12380 : XOR2_X1 port map( A1 => n22198, A2 => n32573, Z => n32572);
   U12384 : INV_X1 port map( I => n16697, ZN => n32573);
   U12385 : NOR2_X2 port map( A1 => n13696, A2 => n7953, ZN => n20755);
   U12386 : NAND2_X2 port map( A1 => n20459, A2 => n28899, ZN => n162);
   U12387 : OAI22_X2 port map( A1 => n32594, A2 => n27741, B1 => n1158, B2 => 
                           n20614, ZN => n20459);
   U12388 : XOR2_X1 port map( A1 => n4287, A2 => n31311, Z => n6863);
   U12389 : NOR3_X2 port map( A1 => n32574, A2 => n29037, A3 => n9736, ZN => 
                           n33748);
   U12390 : NOR2_X1 port map( A1 => n4423, A2 => n16313, ZN => n4422);
   U12392 : XOR2_X1 port map( A1 => n33267, A2 => n18107, Z => n33391);
   U12396 : XOR2_X1 port map( A1 => n32916, A2 => n32575, Z => n15093);
   U12397 : XOR2_X1 port map( A1 => n24475, A2 => n27115, Z => n24547);
   U12399 : NOR2_X2 port map( A1 => n32576, A2 => n7017, ZN => n22302);
   U12400 : NAND2_X1 port map( A1 => n8174, A2 => n11536, ZN => n32576);
   U12409 : OAI21_X2 port map( A1 => n14245, A2 => n14247, B => n14243, ZN => 
                           n25378);
   U12410 : OAI21_X2 port map( A1 => n31962, A2 => n33915, B => n33914, ZN => 
                           n14245);
   U12411 : NAND2_X2 port map( A1 => n30015, A2 => n12705, ZN => n5003);
   U12414 : XOR2_X1 port map( A1 => n19616, A2 => n19615, Z => n19617);
   U12416 : OAI21_X2 port map( A1 => n17453, A2 => n28120, B => n15253, ZN => 
                           n14288);
   U12419 : XOR2_X1 port map( A1 => n6735, A2 => n32578, Z => n9322);
   U12425 : XOR2_X1 port map( A1 => n6739, A2 => n16178, Z => n32578);
   U12426 : NAND2_X1 port map( A1 => n3772, A2 => n3771, ZN => n32615);
   U12428 : OAI22_X2 port map( A1 => n32579, A2 => n25007, B1 => n3231, B2 => 
                           n3230, ZN => n31182);
   U12429 : AOI21_X2 port map( A1 => n3230, A2 => n25002, B => n31122, ZN => 
                           n32579);
   U12430 : NAND3_X2 port map( A1 => n28776, A2 => n29401, A3 => n32580, ZN => 
                           n23508);
   U12433 : NAND2_X2 port map( A1 => n5091, A2 => n25709, ZN => n4706);
   U12434 : NOR2_X1 port map( A1 => n8086, A2 => n24212, ZN => n26914);
   U12435 : INV_X4 port map( I => n21601, ZN => n5704);
   U12437 : NAND2_X2 port map( A1 => n7651, A2 => n329, ZN => n21601);
   U12444 : XOR2_X1 port map( A1 => n86, A2 => n85, Z => n22656);
   U12445 : NOR2_X2 port map( A1 => n3515, A2 => n6763, ZN => n5032);
   U12449 : XOR2_X1 port map( A1 => n28405, A2 => n32582, Z => n13189);
   U12459 : XOR2_X1 port map( A1 => n14968, A2 => n20640, Z => n32582);
   U12460 : NAND2_X2 port map( A1 => n12577, A2 => n23071, ZN => n6676);
   U12461 : XOR2_X1 port map( A1 => n21001, A2 => n20730, Z => n16175);
   U12464 : OAI21_X2 port map( A1 => n13783, A2 => n13784, B => n13782, ZN => 
                           n21001);
   U12465 : INV_X4 port map( I => n3515, ZN => n2935);
   U12466 : XOR2_X1 port map( A1 => n24807, A2 => n4329, Z => n9571);
   U12474 : NAND2_X2 port map( A1 => n27660, A2 => n27439, ZN => n24807);
   U12476 : NAND2_X2 port map( A1 => n11557, A2 => n12770, ZN => n2958);
   U12477 : AOI22_X2 port map( A1 => n20036, A2 => n2549, B1 => n14210, B2 => 
                           n12337, ZN => n12770);
   U12486 : NAND2_X1 port map( A1 => n13130, A2 => n21506, ZN => n11687);
   U12487 : NAND2_X2 port map( A1 => n33052, A2 => n28485, ZN => n20670);
   U12488 : NAND2_X2 port map( A1 => n8107, A2 => n11872, ZN => n12296);
   U12494 : NAND2_X2 port map( A1 => n20238, A2 => n11453, ZN => n20075);
   U12495 : NOR2_X2 port map( A1 => n11454, A2 => n2387, ZN => n11453);
   U12496 : XOR2_X1 port map( A1 => n7748, A2 => n25274, Z => n4944);
   U12500 : NAND2_X2 port map( A1 => n7108, A2 => n7109, ZN => n7748);
   U12502 : OAI21_X2 port map( A1 => n31507, A2 => n31730, B => n21445, ZN => 
                           n21827);
   U12503 : AOI22_X2 port map( A1 => n21307, A2 => n21305, B1 => n16526, B2 => 
                           n21443, ZN => n21445);
   U12505 : INV_X2 port map( I => n32584, ZN => n29460);
   U12507 : XOR2_X1 port map( A1 => n17281, A2 => n6205, Z => n32584);
   U12514 : OAI21_X2 port map( A1 => n33850, A2 => n9393, B => n9392, ZN => 
                           n32898);
   U12516 : NOR2_X2 port map( A1 => n8380, A2 => n17805, ZN => n24234);
   U12518 : NAND2_X1 port map( A1 => n33383, A2 => n33382, ZN => n7217);
   U12531 : NAND3_X2 port map( A1 => n1873, A2 => n9339, A3 => n9338, ZN => 
                           n30031);
   U12533 : XOR2_X1 port map( A1 => n11490, A2 => n19531, Z => n14316);
   U12536 : NAND2_X2 port map( A1 => n18669, A2 => n18668, ZN => n11490);
   U12539 : NAND2_X2 port map( A1 => n33536, A2 => n31932, ZN => n22455);
   U12540 : XOR2_X1 port map( A1 => n2423, A2 => n32586, Z => n8492);
   U12541 : XOR2_X1 port map( A1 => n17682, A2 => n24752, Z => n32586);
   U12542 : AOI21_X2 port map( A1 => n4071, A2 => n20541, B => n782, ZN => 
                           n10718);
   U12550 : NAND2_X2 port map( A1 => n7123, A2 => n7120, ZN => n30346);
   U12553 : NAND2_X2 port map( A1 => n7118, A2 => n27515, ZN => n7123);
   U12558 : OAI21_X1 port map( A1 => n1628, A2 => n4150, B => n1627, ZN => 
                           n32587);
   U12564 : NOR2_X2 port map( A1 => n30769, A2 => n21697, ZN => n32588);
   U12570 : NAND2_X2 port map( A1 => n19198, A2 => n19200, ZN => n28883);
   U12573 : NAND2_X2 port map( A1 => n5813, A2 => n19199, ZN => n19198);
   U12574 : XOR2_X1 port map( A1 => n14855, A2 => n13470, Z => n4729);
   U12575 : INV_X2 port map( I => n29278, ZN => n32590);
   U12580 : NAND2_X2 port map( A1 => n1214, A2 => n30241, ZN => n32592);
   U12581 : INV_X2 port map( I => n28358, ZN => n25210);
   U12582 : NAND2_X2 port map( A1 => n4533, A2 => n33024, ZN => n28358);
   U12585 : XOR2_X1 port map( A1 => n4354, A2 => n32593, Z => n14911);
   U12587 : XOR2_X1 port map( A1 => n4352, A2 => n4353, Z => n32593);
   U12588 : AND2_X2 port map( A1 => n8838, A2 => n23834, Z => n30060);
   U12589 : BUF_X2 port map( I => n17746, Z => n32594);
   U12593 : NAND3_X1 port map( A1 => n32596, A2 => n849, A3 => n32595, ZN => 
                           n27263);
   U12594 : INV_X2 port map( I => n13807, ZN => n32595);
   U12595 : INV_X1 port map( I => n23066, ZN => n32596);
   U12596 : NAND2_X1 port map( A1 => n18842, A2 => n33232, ZN => n33231);
   U12597 : AOI21_X2 port map( A1 => n3219, A2 => n25974, B => n32597, ZN => 
                           n3234);
   U12601 : AND2_X1 port map( A1 => n3221, A2 => n3222, Z => n32597);
   U12603 : NAND2_X2 port map( A1 => n2727, A2 => n2642, ZN => n25142);
   U12604 : XOR2_X1 port map( A1 => n32111, A2 => n20992, Z => n12330);
   U12611 : INV_X2 port map( I => n31017, ZN => n16623);
   U12612 : XOR2_X1 port map( A1 => n33604, A2 => n4840, Z => n25894);
   U12614 : AOI21_X2 port map( A1 => n30154, A2 => n16241, B => n30152, ZN => 
                           n32598);
   U12615 : XOR2_X1 port map( A1 => n23145, A2 => n6348, Z => n5194);
   U12621 : XOR2_X1 port map( A1 => n23271, A2 => n33971, Z => n6348);
   U12624 : OAI22_X2 port map( A1 => n16623, A2 => n5707, B1 => n20000, B2 => 
                           n10845, ZN => n7281);
   U12631 : INV_X2 port map( I => n10708, ZN => n10845);
   U12633 : NAND2_X2 port map( A1 => n25138, A2 => n32599, ZN => n14189);
   U12635 : NAND2_X2 port map( A1 => n32601, A2 => n32600, ZN => n32599);
   U12636 : NOR2_X2 port map( A1 => n11372, A2 => n9162, ZN => n32600);
   U12637 : INV_X2 port map( I => n17824, ZN => n32601);
   U12638 : XOR2_X1 port map( A1 => n27121, A2 => n14613, Z => n23521);
   U12641 : OAI21_X2 port map( A1 => n32056, A2 => n32603, B => n30817, ZN => 
                           n10297);
   U12642 : NOR2_X1 port map( A1 => n11444, A2 => n6290, ZN => n32603);
   U12643 : BUF_X2 port map( I => n29693, Z => n32604);
   U12644 : INV_X1 port map( I => n10630, ZN => n22631);
   U12646 : NAND2_X2 port map( A1 => n32606, A2 => n32605, ZN => n10630);
   U12647 : INV_X2 port map( I => n7513, ZN => n32606);
   U12650 : NOR2_X2 port map( A1 => n29972, A2 => n20261, ZN => n29528);
   U12652 : NAND2_X2 port map( A1 => n32607, A2 => n27340, ZN => n13412);
   U12653 : NAND2_X1 port map( A1 => n14531, A2 => n7765, ZN => n12458);
   U12657 : XOR2_X1 port map( A1 => n11205, A2 => n15710, Z => n32925);
   U12659 : OAI21_X2 port map( A1 => n7626, A2 => n5895, B => n5893, ZN => 
                           n15710);
   U12662 : NAND3_X2 port map( A1 => n31657, A2 => n14305, A3 => n32608, ZN => 
                           n15825);
   U12663 : NAND3_X2 port map( A1 => n32674, A2 => n8431, A3 => n19547, ZN => 
                           n7102);
   U12665 : INV_X2 port map( I => n12758, ZN => n9404);
   U12666 : NAND2_X2 port map( A1 => n20471, A2 => n32504, ZN => n12758);
   U12667 : NOR2_X1 port map( A1 => n1597, A2 => n25746, ZN => n24431);
   U12671 : NAND2_X2 port map( A1 => n31591, A2 => n27486, ZN => n1597);
   U12672 : AOI22_X2 port map( A1 => n2873, A2 => n15162, B1 => n8998, B2 => 
                           n14568, ZN => n14567);
   U12673 : XOR2_X1 port map( A1 => n1173, A2 => n17091, Z => n19662);
   U12675 : NAND2_X2 port map( A1 => n33407, A2 => n13791, ZN => n17091);
   U12677 : AND2_X1 port map( A1 => n5673, A2 => n4286, Z => n31419);
   U12678 : INV_X2 port map( I => n6479, ZN => n32610);
   U12684 : OAI22_X2 port map( A1 => n32612, A2 => n28806, B1 => n4384, B2 => 
                           n4387, ZN => n10915);
   U12688 : XOR2_X1 port map( A1 => n14206, A2 => n20652, Z => n20710);
   U12690 : NAND2_X2 port map( A1 => n20204, A2 => n20203, ZN => n14206);
   U12691 : INV_X1 port map( I => n22426, ZN => n32988);
   U12692 : INV_X2 port map( I => n7072, ZN => n1805);
   U12699 : AND2_X1 port map( A1 => n7868, A2 => n11401, Z => n6807);
   U12703 : BUF_X2 port map( I => n32800, Z => n32613);
   U12707 : XOR2_X1 port map( A1 => n28897, A2 => n11691, Z => n32614);
   U12708 : NOR2_X2 port map( A1 => n18914, A2 => n27076, ZN => n19483);
   U12710 : XOR2_X1 port map( A1 => n10482, A2 => n1130, Z => n417);
   U12711 : XOR2_X1 port map( A1 => n22127, A2 => n8533, Z => n1130);
   U12715 : XOR2_X1 port map( A1 => n32615, A2 => n16619, Z => Ciphertext(96));
   U12720 : XOR2_X1 port map( A1 => n24650, A2 => n24649, Z => n33663);
   U12722 : XOR2_X1 port map( A1 => n968, A2 => n24799, Z => n24650);
   U12724 : XOR2_X1 port map( A1 => n27516, A2 => n32616, Z => n24511);
   U12731 : XOR2_X1 port map( A1 => n24825, A2 => n24508, Z => n32616);
   U12734 : INV_X2 port map( I => n32617, ZN => n12488);
   U12737 : XNOR2_X1 port map( A1 => n31054, A2 => n3120, ZN => n32617);
   U12739 : NOR2_X1 port map( A1 => n17030, A2 => n17029, ZN => n18412);
   U12740 : NOR3_X2 port map( A1 => n2137, A2 => n2138, A3 => n2135, ZN => 
                           n12375);
   U12743 : OR2_X1 port map( A1 => n27897, A2 => n3536, Z => n22490);
   U12746 : XOR2_X1 port map( A1 => n21907, A2 => n33300, Z => n27897);
   U12747 : AND2_X1 port map( A1 => n15964, A2 => n25586, Z => n24631);
   U12748 : XOR2_X1 port map( A1 => n32255, A2 => n3722, Z => n22037);
   U12751 : BUF_X2 port map( I => n20043, Z => n32618);
   U12752 : BUF_X2 port map( I => n10714, Z => n32619);
   U12756 : XOR2_X1 port map( A1 => n32620, A2 => n31852, Z => n20483);
   U12759 : XOR2_X1 port map( A1 => n20993, A2 => n20482, Z => n32620);
   U12760 : XOR2_X1 port map( A1 => n22251, A2 => n29693, Z => n22150);
   U12763 : OAI22_X2 port map( A1 => n12328, A2 => n6660, B1 => n21776, B2 => 
                           n21775, ZN => n22251);
   U12764 : AND2_X1 port map( A1 => n13667, A2 => n25123, Z => n33413);
   U12768 : OAI21_X2 port map( A1 => n32621, A2 => n4596, B => n19140, ZN => 
                           n4595);
   U12771 : INV_X2 port map( I => n19189, ZN => n32621);
   U12772 : NAND2_X2 port map( A1 => n744, A2 => n13160, ZN => n19189);
   U12777 : INV_X1 port map( I => n31325, ZN => n32837);
   U12778 : NAND3_X2 port map( A1 => n880, A2 => n7732, A3 => n11970, ZN => 
                           n32622);
   U12779 : BUF_X2 port map( I => n21203, Z => n32625);
   U12783 : NAND2_X2 port map( A1 => n17771, A2 => n32626, ZN => n24996);
   U12786 : NAND2_X2 port map( A1 => n34099, A2 => n1559, ZN => n21532);
   U12787 : NOR2_X2 port map( A1 => n22362, A2 => n8471, ZN => n22542);
   U12789 : NAND2_X2 port map( A1 => n10489, A2 => n10486, ZN => n8568);
   U12791 : XOR2_X1 port map( A1 => n32627, A2 => n6903, Z => n7912);
   U12802 : XOR2_X1 port map( A1 => n30482, A2 => n30362, Z => n32627);
   U12803 : AOI22_X2 port map( A1 => n10054, A2 => n19109, B1 => n19110, B2 => 
                           n27921, ZN => n28996);
   U12804 : INV_X2 port map( I => n32628, ZN => n26448);
   U12806 : XNOR2_X1 port map( A1 => n9040, A2 => n9037, ZN => n32628);
   U12812 : XOR2_X1 port map( A1 => n29702, A2 => n19631, Z => n14814);
   U12818 : NAND2_X1 port map( A1 => n22745, A2 => n27166, ZN => n33503);
   U12821 : XOR2_X1 port map( A1 => n31639, A2 => n32629, Z => n24779);
   U12830 : XOR2_X1 port map( A1 => n24619, A2 => n33348, Z => n32629);
   U12840 : AOI21_X1 port map( A1 => n32630, A2 => n16273, B => n12457, ZN => 
                           n12456);
   U12843 : NAND2_X1 port map( A1 => n12458, A2 => n16279, ZN => n32630);
   U12845 : OR2_X1 port map( A1 => n24027, A2 => n32934, Z => n29292);
   U12848 : INV_X2 port map( I => n32631, ZN => n22670);
   U12853 : XOR2_X1 port map( A1 => n24825, A2 => n32632, Z => n27946);
   U12854 : XOR2_X1 port map( A1 => n4240, A2 => n12665, Z => n32632);
   U12855 : XOR2_X1 port map( A1 => n23174, A2 => n23189, Z => n32633);
   U12859 : NAND2_X1 port map( A1 => n4814, A2 => n24976, ZN => n32735);
   U12860 : NAND2_X2 port map( A1 => n12642, A2 => n11214, ZN => n12866);
   U12862 : NOR2_X2 port map( A1 => n29047, A2 => n29093, ZN => n32634);
   U12863 : XOR2_X1 port map( A1 => n19538, A2 => n32184, Z => n14743);
   U12866 : NAND2_X2 port map( A1 => n14749, A2 => n14750, ZN => n32635);
   U12875 : AOI21_X2 port map( A1 => n8499, A2 => n5690, B => n27592, ZN => 
                           n10793);
   U12876 : OAI22_X2 port map( A1 => n9516, A2 => n9334, B1 => n32636, B2 => 
                           n9647, ZN => n22949);
   U12878 : AOI22_X2 port map( A1 => n14993, A2 => n25013, B1 => n24976, B2 => 
                           n14992, ZN => n32637);
   U12882 : OAI22_X2 port map( A1 => n5264, A2 => n1317, B1 => n21821, B2 => 
                           n5546, ZN => n21562);
   U12885 : XOR2_X1 port map( A1 => n29674, A2 => n26371, Z => n30187);
   U12890 : XOR2_X1 port map( A1 => n2809, A2 => n32638, Z => n27894);
   U12895 : XOR2_X1 port map( A1 => n33933, A2 => n32639, Z => n32638);
   U12898 : XOR2_X1 port map( A1 => n9983, A2 => n32640, Z => n33253);
   U12900 : XOR2_X1 port map( A1 => n23331, A2 => n23332, Z => n23437);
   U12901 : NOR2_X2 port map( A1 => n2086, A2 => n32641, ZN => n10523);
   U12902 : AOI21_X2 port map( A1 => n10524, A2 => n20338, B => n20591, ZN => 
                           n32641);
   U12904 : AND2_X1 port map( A1 => n30233, A2 => n32643, Z => n34148);
   U12906 : NOR2_X1 port map( A1 => n33565, A2 => n26615, ZN => n33187);
   U12907 : XOR2_X1 port map( A1 => n19466, A2 => n16584, Z => n19385);
   U12912 : OAI22_X2 port map( A1 => n27420, A2 => n16741, B1 => n7419, B2 => 
                           n18751, ZN => n19466);
   U12916 : BUF_X2 port map( I => n9678, Z => n32644);
   U12917 : NAND2_X2 port map( A1 => n792, A2 => n13601, ZN => n24269);
   U12919 : XOR2_X1 port map( A1 => n11736, A2 => n22227, Z => n22143);
   U12920 : NAND2_X2 port map( A1 => n13029, A2 => n3050, ZN => n11736);
   U12922 : NAND2_X1 port map( A1 => n32712, A2 => n16976, ZN => n26858);
   U12923 : NAND2_X2 port map( A1 => n33044, A2 => n31946, ZN => n7586);
   U12926 : AOI22_X2 port map( A1 => n16673, A2 => n25859, B1 => n14915, B2 => 
                           n25863, ZN => n25836);
   U12932 : XOR2_X1 port map( A1 => n32645, A2 => n23407, Z => n236);
   U12933 : NOR2_X2 port map( A1 => n9277, A2 => n29138, ZN => n10226);
   U12935 : XOR2_X1 port map( A1 => n32646, A2 => n29609, Z => Ciphertext(50));
   U12936 : OAI22_X1 port map( A1 => n29076, A2 => n25097, B1 => n25095, B2 => 
                           n4193, ZN => n32646);
   U12938 : NAND2_X2 port map( A1 => n5897, A2 => n14454, ZN => n15646);
   U12939 : NOR2_X2 port map( A1 => n14281, A2 => n16009, ZN => n7643);
   U12940 : AOI22_X2 port map( A1 => n29180, A2 => n28581, B1 => n10875, B2 => 
                           n9793, ZN => n29577);
   U12941 : OAI21_X1 port map( A1 => n14117, A2 => n18460, B => n15070, ZN => 
                           n15069);
   U12942 : NOR2_X2 port map( A1 => n33688, A2 => n33687, ZN => n14117);
   U12945 : OAI21_X2 port map( A1 => n1278, A2 => n6975, B => n22747, ZN => 
                           n22784);
   U12946 : NAND2_X2 port map( A1 => n15633, A2 => n14540, ZN => n22747);
   U12954 : NOR2_X1 port map( A1 => n31967, A2 => n3084, ZN => n3085);
   U12966 : NAND2_X2 port map( A1 => n33439, A2 => n3061, ZN => n3084);
   U12967 : NOR2_X1 port map( A1 => n18715, A2 => n18716, ZN => n18717);
   U12970 : INV_X1 port map( I => n33153, ZN => n32647);
   U12973 : NAND2_X2 port map( A1 => n7689, A2 => n25891, ZN => n24985);
   U12975 : XOR2_X1 port map( A1 => n24751, A2 => n7135, Z => n2423);
   U12979 : NAND2_X2 port map( A1 => n10848, A2 => n20405, ZN => n5581);
   U12985 : NAND2_X2 port map( A1 => n27965, A2 => n25968, ZN => n8051);
   U12986 : OAI21_X2 port map( A1 => n32649, A2 => n33974, B => n12531, ZN => 
                           n13679);
   U12987 : NOR2_X1 port map( A1 => n12556, A2 => n15911, ZN => n32649);
   U12988 : OR2_X2 port map( A1 => n13427, A2 => n32652, Z => n24888);
   U12994 : XOR2_X1 port map( A1 => n19307, A2 => n14459, Z => n30770);
   U12995 : XOR2_X1 port map( A1 => n29856, A2 => n19403, Z => n29661);
   U13002 : NOR2_X1 port map( A1 => n10433, A2 => n7119, ZN => n21117);
   U13003 : XOR2_X1 port map( A1 => n19598, A2 => n10210, Z => n10079);
   U13004 : XOR2_X1 port map( A1 => n2611, A2 => n19470, Z => n19598);
   U13005 : XOR2_X1 port map( A1 => n32650, A2 => n33778, Z => n11907);
   U13008 : XOR2_X1 port map( A1 => n22166, A2 => n15367, Z => n32650);
   U13011 : XOR2_X1 port map( A1 => n29906, A2 => n13214, Z => n28034);
   U13013 : NOR2_X2 port map( A1 => n20751, A2 => n17341, ZN => n28586);
   U13019 : NAND2_X2 port map( A1 => n32651, A2 => n14019, ZN => n26557);
   U13020 : NAND2_X2 port map( A1 => n30366, A2 => n13077, ZN => n32651);
   U13025 : XOR2_X1 port map( A1 => n19649, A2 => n16349, Z => n19497);
   U13031 : NAND2_X2 port map( A1 => n18421, A2 => n18420, ZN => n19649);
   U13032 : INV_X4 port map( I => n6765, ZN => n11981);
   U13034 : NAND2_X2 port map( A1 => n12506, A2 => n26302, ZN => n6765);
   U13037 : NAND2_X2 port map( A1 => n4800, A2 => n27811, ZN => n7465);
   U13039 : NAND2_X2 port map( A1 => n33165, A2 => n33166, ZN => n4800);
   U13044 : XOR2_X1 port map( A1 => n7808, A2 => n22231, Z => n21993);
   U13046 : NOR2_X2 port map( A1 => n11053, A2 => n30634, ZN => n7808);
   U13053 : OAI21_X2 port map( A1 => n12226, A2 => n12225, B => n10939, ZN => 
                           n12228);
   U13056 : INV_X2 port map( I => n8492, ZN => n32652);
   U13058 : XOR2_X1 port map( A1 => n20917, A2 => n29241, Z => n21017);
   U13060 : OAI21_X2 port map( A1 => n20177, A2 => n20176, B => n20175, ZN => 
                           n29241);
   U13061 : NOR2_X1 port map( A1 => n11876, A2 => n28721, ZN => n32653);
   U13062 : OAI21_X2 port map( A1 => n655, A2 => n34166, B => n23891, ZN => 
                           n1818);
   U13063 : XOR2_X1 port map( A1 => n30421, A2 => n30274, Z => n33651);
   U13065 : XOR2_X1 port map( A1 => n34062, A2 => n30229, Z => n13922);
   U13066 : NOR2_X2 port map( A1 => n24148, A2 => n1775, ZN => n1973);
   U13076 : NOR2_X2 port map( A1 => n14233, A2 => n32485, ZN => n10740);
   U13077 : NOR2_X2 port map( A1 => n32654, A2 => n16232, ZN => n14749);
   U13085 : XNOR2_X1 port map( A1 => n12459, A2 => n16708, ZN => n20746);
   U13086 : OAI21_X2 port map( A1 => n28641, A2 => n7690, B => n15589, ZN => 
                           n32655);
   U13091 : NAND2_X1 port map( A1 => n28329, A2 => n7993, ZN => n23914);
   U13094 : NAND2_X1 port map( A1 => n20565, A2 => n16515, ZN => n11368);
   U13098 : OAI21_X2 port map( A1 => n7710, A2 => n33936, B => n23884, ZN => 
                           n32656);
   U13103 : XOR2_X1 port map( A1 => n20641, A2 => n3350, Z => n3351);
   U13104 : NAND3_X2 port map( A1 => n12846, A2 => n12847, A3 => n14263, ZN => 
                           n20641);
   U13107 : NAND2_X1 port map( A1 => n19991, A2 => n937, ZN => n17036);
   U13109 : INV_X2 port map( I => n22615, ZN => n32658);
   U13111 : NAND2_X2 port map( A1 => n851, A2 => n22810, ZN => n22615);
   U13113 : XOR2_X1 port map( A1 => n29810, A2 => n21000, Z => n15817);
   U13114 : XOR2_X1 port map( A1 => n51, A2 => n26656, Z => n1793);
   U13122 : NOR2_X2 port map( A1 => n3951, A2 => n22652, ZN => n51);
   U13126 : OAI21_X2 port map( A1 => n13230, A2 => n21234, B => n29577, ZN => 
                           n34078);
   U13131 : NAND3_X2 port map( A1 => n1077, A2 => n4407, A3 => n24712, ZN => 
                           n31372);
   U13133 : XOR2_X1 port map( A1 => n9353, A2 => n8949, Z => n24568);
   U13148 : NAND3_X2 port map( A1 => n28703, A2 => n1504, A3 => n27735, ZN => 
                           n9353);
   U13163 : XOR2_X1 port map( A1 => n6904, A2 => n22267, Z => n33214);
   U13165 : XOR2_X1 port map( A1 => n4228, A2 => n7477, Z => n6904);
   U13166 : NAND3_X2 port map( A1 => n19120, A2 => n19181, A3 => n19180, ZN => 
                           n8905);
   U13171 : XOR2_X1 port map( A1 => n1003, A2 => n29121, Z => n7288);
   U13173 : NAND2_X2 port map( A1 => n4880, A2 => n8122, ZN => n29121);
   U13174 : AND2_X2 port map( A1 => n2234, A2 => n29052, Z => n27117);
   U13177 : XOR2_X1 port map( A1 => n32661, A2 => n20902, Z => n5241);
   U13179 : XOR2_X1 port map( A1 => n21046, A2 => n5024, Z => n32661);
   U13180 : OAI21_X2 port map( A1 => n4514, A2 => n23787, B => n30803, ZN => 
                           n7935);
   U13183 : NAND2_X2 port map( A1 => n25210, A2 => n5578, ZN => n7305);
   U13187 : OAI21_X2 port map( A1 => n28688, A2 => n2233, B => n23544, ZN => 
                           n32866);
   U13192 : NAND2_X2 port map( A1 => n32662, A2 => n31967, ZN => n29780);
   U13194 : NAND2_X2 port map( A1 => n26756, A2 => n3084, ZN => n32662);
   U13197 : AOI22_X2 port map( A1 => n1280, A2 => n22981, B1 => n34163, B2 => 
                           n28934, ZN => n29791);
   U13200 : OAI21_X1 port map( A1 => n33500, A2 => n29362, B => n31945, ZN => 
                           n33728);
   U13204 : XOR2_X1 port map( A1 => n15948, A2 => n11995, Z => n25589);
   U13206 : OAI21_X2 port map( A1 => n32663, A2 => n32716, B => n22726, ZN => 
                           n31727);
   U13208 : NAND2_X1 port map( A1 => n22725, A2 => n14555, ZN => n32663);
   U13212 : XOR2_X1 port map( A1 => n22037, A2 => n33217, Z => n12622);
   U13213 : OAI22_X2 port map( A1 => n1998, A2 => n1235, B1 => n1940, B2 => 
                           n24244, ZN => n1997);
   U13215 : NAND2_X2 port map( A1 => n1235, A2 => n28374, ZN => n1940);
   U13216 : BUF_X4 port map( I => n5440, Z => n33320);
   U13219 : XOR2_X1 port map( A1 => n1713, A2 => n32664, Z => n7012);
   U13228 : XOR2_X1 port map( A1 => n34050, A2 => n1712, Z => n32664);
   U13230 : INV_X2 port map( I => n32665, ZN => n17289);
   U13231 : NAND2_X2 port map( A1 => n31539, A2 => n28949, ZN => n32665);
   U13233 : INV_X1 port map( I => n23464, ZN => n33609);
   U13234 : XOR2_X1 port map( A1 => n12796, A2 => n7387, Z => n12795);
   U13238 : NAND2_X2 port map( A1 => n32666, A2 => n31359, ZN => n16060);
   U13239 : NOR2_X2 port map( A1 => n30962, A2 => n30963, ZN => n32666);
   U13242 : NAND2_X2 port map( A1 => n9775, A2 => n9773, ZN => n12478);
   U13244 : XOR2_X1 port map( A1 => n9189, A2 => n30883, Z => n24358);
   U13254 : NOR2_X2 port map( A1 => n32829, A2 => n30000, ZN => n2691);
   U13258 : XOR2_X1 port map( A1 => n15666, A2 => n15669, Z => n15226);
   U13259 : INV_X4 port map( I => n33616, ZN => n26120);
   U13260 : XOR2_X1 port map( A1 => n6758, A2 => n27174, Z => n6757);
   U13262 : NAND2_X2 port map( A1 => n13764, A2 => n25546, ZN => n31360);
   U13267 : NAND3_X2 port map( A1 => n33327, A2 => n25535, A3 => n25534, ZN => 
                           n13764);
   U13269 : NOR3_X2 port map( A1 => n8095, A2 => n30089, A3 => n33867, ZN => 
                           n8094);
   U13275 : NOR2_X1 port map( A1 => n7080, A2 => n4951, ZN => n32667);
   U13277 : NOR2_X2 port map( A1 => n17110, A2 => n32659, ZN => n32668);
   U13283 : NAND2_X2 port map( A1 => n9472, A2 => n21870, ZN => n21632);
   U13284 : NAND2_X2 port map( A1 => n33068, A2 => n33066, ZN => n25387);
   U13285 : NAND2_X2 port map( A1 => n32669, A2 => n4991, ZN => n7384);
   U13287 : NAND2_X2 port map( A1 => n33260, A2 => n33789, ZN => n32669);
   U13289 : NAND2_X2 port map( A1 => n118, A2 => n28058, ZN => n22979);
   U13293 : XOR2_X1 port map( A1 => n1228, A2 => n6168, Z => n24800);
   U13295 : XOR2_X1 port map( A1 => n21019, A2 => n20900, Z => n20984);
   U13299 : NAND2_X2 port map( A1 => n11104, A2 => n33815, ZN => n21019);
   U13300 : NAND2_X2 port map( A1 => n3844, A2 => n30336, ZN => n19275);
   U13301 : XOR2_X1 port map( A1 => n20649, A2 => n26691, Z => n519);
   U13302 : NAND2_X2 port map( A1 => n19232, A2 => n32671, ZN => n32670);
   U13303 : OAI21_X2 port map( A1 => n28856, A2 => n10478, B => n19825, ZN => 
                           n32747);
   U13309 : AOI21_X2 port map( A1 => n1152, A2 => n13920, B => n32672, ZN => 
                           n4534);
   U13310 : OAI21_X2 port map( A1 => n13920, A2 => n13538, B => n13300, ZN => 
                           n32672);
   U13311 : NAND2_X2 port map( A1 => n18206, A2 => n18208, ZN => n6718);
   U13312 : NOR2_X2 port map( A1 => n18207, A2 => n21230, ZN => n18206);
   U13314 : NAND2_X2 port map( A1 => n32673, A2 => n17944, ZN => n6899);
   U13318 : XOR2_X1 port map( A1 => n24394, A2 => n13545, Z => n24619);
   U13319 : BUF_X4 port map( I => n16451, Z => n11703);
   U13327 : NAND2_X2 port map( A1 => n22922, A2 => n22921, ZN => n30868);
   U13328 : NAND2_X2 port map( A1 => n33433, A2 => n252, ZN => n22922);
   U13329 : AOI22_X2 port map( A1 => n5598, A2 => n15394, B1 => n820, B2 => 
                           n26130, ZN => n8406);
   U13332 : INV_X2 port map( I => n27781, ZN => n19691);
   U13333 : NAND2_X2 port map( A1 => n32676, A2 => n32675, ZN => n27781);
   U13335 : NAND2_X1 port map( A1 => n17716, A2 => n32679, ZN => n6145);
   U13337 : OR2_X1 port map( A1 => n2386, A2 => n16077, Z => n32679);
   U13341 : XOR2_X1 port map( A1 => n24805, A2 => n12800, Z => n13471);
   U13342 : NAND2_X2 port map( A1 => n18946, A2 => n18947, ZN => n30443);
   U13343 : AOI22_X2 port map( A1 => n13197, A2 => n22396, B1 => n10757, B2 => 
                           n1124, ZN => n8601);
   U13346 : OAI21_X2 port map( A1 => n7110, A2 => n31152, B => n32681, ZN => 
                           n3057);
   U13355 : NOR2_X2 port map( A1 => n27617, A2 => n27616, ZN => n32681);
   U13363 : NOR2_X2 port map( A1 => n32790, A2 => n13160, ZN => n27420);
   U13364 : NAND2_X2 port map( A1 => n17446, A2 => n6203, ZN => n19260);
   U13365 : AOI21_X2 port map( A1 => n33116, A2 => n20595, B => n817, ZN => 
                           n20176);
   U13366 : XOR2_X1 port map( A1 => n6812, A2 => n22075, Z => n21912);
   U13367 : OAI21_X2 port map( A1 => n32682, A2 => n27987, B => n22959, ZN => 
                           n23286);
   U13373 : NOR2_X1 port map( A1 => n28877, A2 => n28878, ZN => n32682);
   U13374 : NAND2_X2 port map( A1 => n16607, A2 => n2092, ZN => n3842);
   U13377 : XOR2_X1 port map( A1 => n22192, A2 => n32683, Z => n526);
   U13384 : INV_X1 port map( I => n25355, ZN => n32683);
   U13387 : INV_X4 port map( I => n20613, ZN => n1158);
   U13390 : NAND2_X2 port map( A1 => n13954, A2 => n13955, ZN => n20613);
   U13395 : NOR2_X2 port map( A1 => n32684, A2 => n26633, ZN => n26632);
   U13396 : OAI21_X2 port map( A1 => n32671, A2 => n18415, B => n32685, ZN => 
                           n18421);
   U13397 : NAND2_X2 port map( A1 => n33712, A2 => n18419, ZN => n32685);
   U13406 : OAI21_X2 port map( A1 => n32686, A2 => n3163, B => n28970, ZN => 
                           n30753);
   U13407 : INV_X1 port map( I => n32687, ZN => n32686);
   U13416 : NOR2_X1 port map( A1 => n724, A2 => n13694, ZN => n32687);
   U13421 : INV_X2 port map( I => n10948, ZN => n11931);
   U13423 : NAND3_X2 port map( A1 => n15287, A2 => n25580, A3 => n25579, ZN => 
                           n10948);
   U13424 : NOR2_X1 port map( A1 => n30204, A2 => n11366, ZN => n15531);
   U13425 : NAND2_X2 port map( A1 => n32688, A2 => n9884, ZN => n21925);
   U13430 : XOR2_X1 port map( A1 => n32689, A2 => n17914, Z => Ciphertext(85));
   U13431 : AOI22_X1 port map( A1 => n27680, A2 => n25268, B1 => n25286, B2 => 
                           n25280, ZN => n32689);
   U13434 : NAND2_X2 port map( A1 => n33238, A2 => n32690, ZN => n4184);
   U13440 : AND2_X1 port map( A1 => n29620, A2 => n13193, Z => n32690);
   U13443 : INV_X2 port map( I => n24340, ZN => n29567);
   U13444 : NAND2_X2 port map( A1 => n4460, A2 => n20238, ZN => n20302);
   U13451 : NOR2_X2 port map( A1 => n19847, A2 => n31644, ZN => n4460);
   U13453 : NAND2_X2 port map( A1 => n1878, A2 => n32691, ZN => n7232);
   U13454 : NAND2_X2 port map( A1 => n2694, A2 => n15072, ZN => n32691);
   U13455 : NAND2_X1 port map( A1 => n2694, A2 => n19845, ZN => n2693);
   U13458 : NAND2_X1 port map( A1 => n14486, A2 => n14485, ZN => n3788);
   U13459 : NAND2_X2 port map( A1 => n29780, A2 => n16251, ZN => n14486);
   U13462 : AND2_X1 port map( A1 => n24308, A2 => n11041, Z => n28428);
   U13463 : NAND2_X1 port map( A1 => n32693, A2 => n32692, ZN => n7942);
   U13473 : INV_X1 port map( I => n1279, ZN => n32693);
   U13475 : NAND2_X2 port map( A1 => n6512, A2 => n24430, ZN => n25736);
   U13476 : NAND4_X2 port map( A1 => n277, A2 => n25627, A3 => n25584, A4 => 
                           n17863, ZN => n6512);
   U13478 : XOR2_X1 port map( A1 => n32694, A2 => n17564, Z => n8366);
   U13481 : XOR2_X1 port map( A1 => n33509, A2 => n32695, Z => n32694);
   U13482 : OAI21_X2 port map( A1 => n17661, A2 => n11904, B => n1100, ZN => 
                           n155);
   U13483 : XOR2_X1 port map( A1 => n32696, A2 => n22037, Z => n32947);
   U13484 : XOR2_X1 port map( A1 => n4219, A2 => n22283, Z => n9914);
   U13485 : BUF_X2 port map( I => n31568, Z => n32697);
   U13492 : XOR2_X1 port map( A1 => n12785, A2 => n12789, Z => n17745);
   U13493 : NAND2_X2 port map( A1 => n12787, A2 => n12786, ZN => n12789);
   U13494 : NAND2_X2 port map( A1 => n30215, A2 => n27034, ZN => n2449);
   U13498 : XOR2_X1 port map( A1 => n20753, A2 => n20558, Z => n11337);
   U13510 : XOR2_X1 port map( A1 => n23194, A2 => n32698, Z => n23197);
   U13515 : XOR2_X1 port map( A1 => n23210, A2 => n29719, Z => n32698);
   U13516 : AOI21_X2 port map( A1 => n19236, A2 => n3515, B => n31139, ZN => 
                           n2280);
   U13524 : XOR2_X1 port map( A1 => n32699, A2 => n18001, Z => n30131);
   U13525 : XOR2_X1 port map( A1 => n24427, A2 => n8050, Z => n32699);
   U13532 : OAI22_X2 port map( A1 => n30371, A2 => n18515, B1 => n1188, B2 => 
                           n13663, ZN => n6470);
   U13533 : XOR2_X1 port map( A1 => n31892, A2 => n32700, Z => n26930);
   U13534 : XOR2_X1 port map( A1 => n23240, A2 => n23238, Z => n32700);
   U13538 : XOR2_X1 port map( A1 => n23389, A2 => n31523, Z => n23213);
   U13540 : OAI21_X2 port map( A1 => n5681, A2 => n23485, B => n5680, ZN => 
                           n23389);
   U13541 : AOI21_X2 port map( A1 => n22714, A2 => n14188, B => n32701, ZN => 
                           n16160);
   U13542 : OAI22_X2 port map( A1 => n15364, A2 => n14188, B1 => n27389, B2 => 
                           n22836, ZN => n32701);
   U13548 : NAND2_X1 port map( A1 => n16197, A2 => n16198, ZN => n30081);
   U13549 : NAND2_X2 port map( A1 => n32995, A2 => n26501, ZN => n33971);
   U13550 : OAI21_X2 port map( A1 => n28414, A2 => n30869, B => n20429, ZN => 
                           n10992);
   U13552 : XOR2_X1 port map( A1 => n32702, A2 => n16605, Z => Ciphertext(130))
                           ;
   U13553 : XOR2_X1 port map( A1 => n24481, A2 => n24482, Z => n32703);
   U13554 : NAND2_X2 port map( A1 => n29539, A2 => n30277, ZN => n10097);
   U13560 : OAI21_X1 port map( A1 => n14020, A2 => n25014, B => n30461, ZN => 
                           n34043);
   U13561 : NAND2_X2 port map( A1 => n3247, A2 => n31645, ZN => n30314);
   U13562 : AOI22_X2 port map( A1 => n32949, A2 => n8886, B1 => n21585, B2 => 
                           n3248, ZN => n3247);
   U13566 : NOR2_X1 port map( A1 => n33032, A2 => n22873, ZN => n32704);
   U13569 : OAI21_X2 port map( A1 => n22956, A2 => n15601, B => n22955, ZN => 
                           n27988);
   U13574 : INV_X4 port map( I => n28714, ZN => n1020);
   U13577 : OAI21_X2 port map( A1 => n22825, A2 => n22823, B => n32705, ZN => 
                           n23467);
   U13578 : INV_X2 port map( I => n13334, ZN => n719);
   U13580 : NAND2_X2 port map( A1 => n15155, A2 => n2378, ZN => n32950);
   U13582 : XOR2_X1 port map( A1 => n7984, A2 => n28746, Z => n15155);
   U13584 : AOI21_X2 port map( A1 => n5555, A2 => n5556, B => n4306, ZN => 
                           n27104);
   U13587 : NAND2_X1 port map( A1 => n13703, A2 => n34058, ZN => n32706);
   U13594 : NAND2_X2 port map( A1 => n23695, A2 => n14078, ZN => n17578);
   U13596 : NAND3_X2 port map( A1 => n17995, A2 => n29081, A3 => n8344, ZN => 
                           n13530);
   U13597 : XOR2_X1 port map( A1 => n31055, A2 => n23312, Z => n6539);
   U13601 : XOR2_X1 port map( A1 => n22288, A2 => n22266, Z => n11816);
   U13602 : XOR2_X1 port map( A1 => n33437, A2 => n22044, Z => n22266);
   U13605 : XOR2_X1 port map( A1 => n32707, A2 => n27699, Z => n2455);
   U13606 : XOR2_X1 port map( A1 => n22070, A2 => n457, Z => n32707);
   U13608 : OAI21_X2 port map( A1 => n5095, A2 => n5096, B => n29621, ZN => 
                           n30870);
   U13613 : NAND3_X1 port map( A1 => n10010, A2 => n27092, A3 => n10007, ZN => 
                           Ciphertext(126));
   U13618 : XOR2_X1 port map( A1 => n32708, A2 => n23311, Z => n10937);
   U13623 : XOR2_X1 port map( A1 => n28072, A2 => n15055, Z => n32708);
   U13624 : INV_X2 port map( I => n25697, ZN => n1718);
   U13627 : NAND2_X2 port map( A1 => n33628, A2 => n33485, ZN => n3711);
   U13629 : XOR2_X1 port map( A1 => n32709, A2 => n16301, Z => Ciphertext(9));
   U13632 : AOI22_X2 port map( A1 => n8780, A2 => n18219, B1 => n10136, B2 => 
                           n24607, ZN => n29532);
   U13633 : AOI21_X2 port map( A1 => n24161, A2 => n30595, B => n3678, ZN => 
                           n31416);
   U13634 : OAI21_X2 port map( A1 => n16640, A2 => n12066, B => n29739, ZN => 
                           n29997);
   U13639 : INV_X2 port map( I => n26385, ZN => n32711);
   U13640 : NAND2_X2 port map( A1 => n33041, A2 => n3255, ZN => n3253);
   U13641 : XOR2_X1 port map( A1 => n32713, A2 => n16680, Z => Ciphertext(73));
   U13642 : OAI22_X1 port map( A1 => n4613, A2 => n4188, B1 => n25207, B2 => 
                           n4614, ZN => n32713);
   U13645 : XOR2_X1 port map( A1 => n13480, A2 => n19749, Z => n15297);
   U13646 : NAND2_X2 port map( A1 => n7403, A2 => n7402, ZN => n13480);
   U13647 : INV_X2 port map( I => n4735, ZN => n22622);
   U13650 : XOR2_X1 port map( A1 => n3812, A2 => n30901, Z => n4735);
   U13654 : INV_X1 port map( I => n22015, ZN => n11863);
   U13655 : XOR2_X1 port map( A1 => n22015, A2 => n32714, Z => n14796);
   U13656 : NOR2_X2 port map( A1 => n28439, A2 => n9493, ZN => n22015);
   U13662 : NAND2_X2 port map( A1 => n34138, A2 => n32739, ZN => n12376);
   U13664 : NOR2_X2 port map( A1 => n15751, A2 => n4041, ZN => n10973);
   U13668 : NAND2_X2 port map( A1 => n1020, A2 => n17313, ZN => n15751);
   U13671 : NOR2_X2 port map( A1 => n5178, A2 => n11956, ZN => n30167);
   U13678 : NOR2_X2 port map( A1 => n5454, A2 => n24168, ZN => n15253);
   U13679 : NAND2_X2 port map( A1 => n13774, A2 => n8675, ZN => n24168);
   U13680 : XOR2_X1 port map( A1 => n23300, A2 => n23488, Z => n32715);
   U13681 : XOR2_X1 port map( A1 => n30303, A2 => n20924, Z => n7031);
   U13688 : OAI22_X2 port map( A1 => n17228, A2 => n10731, B1 => n15832, B2 => 
                           n20516, ZN => n30303);
   U13691 : AOI21_X2 port map( A1 => n5556, A2 => n5555, B => n4306, ZN => 
                           n32877);
   U13692 : OAI22_X2 port map( A1 => n31266, A2 => n23892, B1 => n707, B2 => 
                           n23715, ZN => n4306);
   U13693 : AOI21_X2 port map( A1 => n23111, A2 => n1264, B => n16254, ZN => 
                           n32716);
   U13699 : OR2_X1 port map( A1 => n13176, A2 => n24216, Z => n10179);
   U13700 : INV_X2 port map( I => n24998, ZN => n31122);
   U13702 : NAND2_X2 port map( A1 => n25003, A2 => n2983, ZN => n24998);
   U13703 : XOR2_X1 port map( A1 => n29740, A2 => n22247, Z => n22340);
   U13704 : NAND2_X2 port map( A1 => n30745, A2 => n29799, ZN => n28181);
   U13707 : AND2_X1 port map( A1 => n15772, A2 => n8140, Z => n4668);
   U13708 : NOR2_X2 port map( A1 => n15883, A2 => n32717, ZN => n25479);
   U13712 : INV_X2 port map( I => n24193, ZN => n13040);
   U13713 : NAND2_X2 port map( A1 => n3484, A2 => n31623, ZN => n24193);
   U13718 : OAI21_X2 port map( A1 => n22842, A2 => n22843, B => n23482, ZN => 
                           n22845);
   U13724 : NAND2_X1 port map( A1 => n33938, A2 => n22626, ZN => n6010);
   U13725 : NOR3_X1 port map( A1 => n33102, A2 => n2480, A3 => n25509, ZN => 
                           n25511);
   U13727 : NOR2_X2 port map( A1 => n32719, A2 => n32718, ZN => n17328);
   U13730 : NAND2_X2 port map( A1 => n13570, A2 => n13571, ZN => n32718);
   U13732 : NAND3_X2 port map( A1 => n32720, A2 => n32849, A3 => n19294, ZN => 
                           n7251);
   U13733 : NOR2_X2 port map( A1 => n3181, A2 => n8125, ZN => n31797);
   U13734 : NAND3_X2 port map( A1 => n3166, A2 => n23835, A3 => n28497, ZN => 
                           n8125);
   U13735 : XOR2_X1 port map( A1 => n20852, A2 => n18102, Z => n6758);
   U13738 : NOR2_X1 port map( A1 => n11985, A2 => n11548, ZN => n15738);
   U13743 : NAND2_X2 port map( A1 => n17816, A2 => n32721, ZN => n6911);
   U13745 : NOR2_X2 port map( A1 => n16862, A2 => n10749, ZN => n32721);
   U13747 : XOR2_X1 port map( A1 => n26045, A2 => n24574, Z => n32722);
   U13750 : NAND2_X1 port map( A1 => n8200, A2 => n8201, ZN => n22620);
   U13753 : NOR2_X2 port map( A1 => n5451, A2 => n5449, ZN => n33329);
   U13757 : XOR2_X1 port map( A1 => n26084, A2 => n19556, Z => n18065);
   U13758 : NAND3_X2 port map( A1 => n2371, A2 => n2664, A3 => n32808, ZN => 
                           n31197);
   U13768 : OR2_X1 port map( A1 => n3860, A2 => n33722, Z => n23566);
   U13774 : OAI22_X1 port map( A1 => n5583, A2 => n33714, B1 => n26130, B2 => 
                           n13969, ZN => n32723);
   U13775 : NAND3_X2 port map( A1 => n25262, A2 => n25263, A3 => n6280, ZN => 
                           n30281);
   U13778 : OAI22_X2 port map( A1 => n1207, A2 => n12431, B1 => n16291, B2 => 
                           n25278, ZN => n25286);
   U13781 : NOR2_X1 port map( A1 => n13720, A2 => n29472, ZN => n7475);
   U13785 : NOR2_X2 port map( A1 => n10202, A2 => n11378, ZN => n3186);
   U13788 : NAND2_X2 port map( A1 => n31813, A2 => n24317, ZN => n32725);
   U13800 : XOR2_X1 port map( A1 => n32726, A2 => n6737, Z => n6735);
   U13801 : XOR2_X1 port map( A1 => n31900, A2 => n14060, Z => n19967);
   U13803 : NAND4_X2 port map( A1 => n30886, A2 => n12883, A3 => n12884, A4 => 
                           n13721, ZN => n16940);
   U13806 : OAI21_X2 port map( A1 => n10247, A2 => n11269, B => n32727, ZN => 
                           n10228);
   U13807 : AOI22_X2 port map( A1 => n17190, A2 => n1439, B1 => n18634, B2 => 
                           n15888, ZN => n32727);
   U13809 : XOR2_X1 port map( A1 => n28640, A2 => n6420, Z => n10954);
   U13810 : INV_X1 port map( I => n33846, ZN => n29437);
   U13812 : OR2_X1 port map( A1 => n33846, A2 => n19267, Z => n15759);
   U13813 : XOR2_X1 port map( A1 => n32728, A2 => n33699, Z => n27790);
   U13816 : XOR2_X1 port map( A1 => n27791, A2 => n12, Z => n32728);
   U13817 : INV_X4 port map( I => n16966, ZN => n32746);
   U13818 : NAND3_X2 port map( A1 => n32729, A2 => n29431, A3 => n3065, ZN => 
                           n12748);
   U13820 : NAND2_X1 port map( A1 => n3069, A2 => n3068, ZN => n32729);
   U13832 : XOR2_X1 port map( A1 => n32730, A2 => n25364, Z => Ciphertext(99));
   U13833 : NAND2_X2 port map( A1 => n34096, A2 => n14308, ZN => n22127);
   U13834 : NAND2_X2 port map( A1 => n21492, A2 => n21566, ZN => n33644);
   U13835 : NAND2_X2 port map( A1 => n987, A2 => n5035, ZN => n16202);
   U13840 : NOR2_X1 port map( A1 => n13295, A2 => n8606, ZN => n15628);
   U13841 : NOR2_X2 port map( A1 => n17515, A2 => n13565, ZN => n13295);
   U13843 : XOR2_X1 port map( A1 => n5884, A2 => n5885, Z => n28545);
   U13844 : AND3_X1 port map( A1 => n14255, A2 => n32170, A3 => n14133, Z => 
                           n27893);
   U13845 : XOR2_X1 port map( A1 => n11862, A2 => n14952, Z => n22252);
   U13850 : NOR2_X2 port map( A1 => n28413, A2 => n30374, ZN => n11862);
   U13851 : XOR2_X1 port map( A1 => n20688, A2 => n11512, Z => n11514);
   U13852 : NAND3_X2 port map( A1 => n24137, A2 => n15011, A3 => n6980, ZN => 
                           n33123);
   U13854 : INV_X4 port map( I => n16286, ZN => n9561);
   U13856 : OAI22_X2 port map( A1 => n3825, A2 => n4308, B1 => n18236, B2 => 
                           n20111, ZN => n20560);
   U13857 : NAND2_X2 port map( A1 => n32731, A2 => n31146, ZN => n3489);
   U13861 : XOR2_X1 port map( A1 => n23145, A2 => n23280, Z => n6388);
   U13862 : XOR2_X1 port map( A1 => n2072, A2 => n32732, Z => n2074);
   U13866 : XOR2_X1 port map( A1 => n32733, A2 => n19470, Z => n32732);
   U13867 : INV_X2 port map( I => n4321, ZN => n32733);
   U13869 : XOR2_X1 port map( A1 => n9848, A2 => n13745, Z => n13743);
   U13870 : XOR2_X1 port map( A1 => n24675, A2 => n3694, Z => n9848);
   U13873 : BUF_X4 port map( I => n11676, Z => n29218);
   U13875 : NAND2_X2 port map( A1 => n28652, A2 => n32734, ZN => n14681);
   U13876 : NAND2_X1 port map( A1 => n15113, A2 => n15112, ZN => n32734);
   U13877 : OAI21_X2 port map( A1 => n32735, A2 => n14021, B => n5624, ZN => 
                           n2983);
   U13878 : AND2_X1 port map( A1 => n16305, A2 => n11845, Z => n24318);
   U13880 : INV_X4 port map( I => n5741, ZN => n1243);
   U13881 : NAND2_X2 port map( A1 => n33789, A2 => n33788, ZN => n34164);
   U13883 : NAND2_X2 port map( A1 => n21559, A2 => n6544, ZN => n21852);
   U13884 : OR2_X1 port map( A1 => n30832, A2 => n7811, Z => n15494);
   U13886 : NOR3_X2 port map( A1 => n33730, A2 => n1347, A3 => n3084, ZN => 
                           n2086);
   U13888 : XOR2_X1 port map( A1 => n13833, A2 => n22224, Z => n13862);
   U13889 : NOR2_X2 port map( A1 => n15458, A2 => n32736, ZN => n28081);
   U13895 : NOR2_X1 port map( A1 => n31490, A2 => n1718, ZN => n32736);
   U13897 : AOI22_X2 port map( A1 => n33779, A2 => n12452, B1 => n26439, B2 => 
                           n21672, ZN => n11991);
   U13900 : NOR2_X1 port map( A1 => n32888, A2 => n12040, ZN => n12085);
   U13901 : XOR2_X1 port map( A1 => n34126, A2 => n14985, Z => n12040);
   U13906 : INV_X4 port map( I => n8057, ZN => n20238);
   U13908 : NAND2_X2 port map( A1 => n31062, A2 => n30790, ZN => n8057);
   U13913 : NOR2_X1 port map( A1 => n33031, A2 => n8733, ZN => n30965);
   U13917 : NAND2_X2 port map( A1 => n18976, A2 => n14892, ZN => n1807);
   U13918 : NOR2_X2 port map( A1 => n17131, A2 => n17130, ZN => n14892);
   U13919 : OAI22_X2 port map( A1 => n33748, A2 => n5040, B1 => n976, B2 => 
                           n4675, ZN => n28945);
   U13921 : OAI22_X2 port map( A1 => n20949, A2 => n5822, B1 => n16633, B2 => 
                           n21239, ZN => n2888);
   U13922 : NAND2_X2 port map( A1 => n2888, A2 => n17699, ZN => n33859);
   U13923 : BUF_X2 port map( I => n24226, Z => n32737);
   U13924 : NAND2_X2 port map( A1 => n25187, A2 => n25234, ZN => n13074);
   U13925 : INV_X2 port map( I => n32738, ZN => n33621);
   U13932 : XNOR2_X1 port map( A1 => n18364, A2 => Key(48), ZN => n32738);
   U13947 : NAND2_X1 port map( A1 => n9876, A2 => n20010, ZN => n19789);
   U13948 : INV_X2 port map( I => n10679, ZN => n12323);
   U13950 : NOR2_X1 port map( A1 => n3760, A2 => n33953, ZN => n16430);
   U13959 : XOR2_X1 port map( A1 => n9230, A2 => n14766, Z => n27571);
   U13960 : XOR2_X1 port map( A1 => n29262, A2 => n5875, Z => n4087);
   U13962 : XOR2_X1 port map( A1 => n22030, A2 => n27837, Z => n29262);
   U13963 : NOR2_X1 port map( A1 => n19907, A2 => n19958, ZN => n29284);
   U13965 : AOI22_X2 port map( A1 => n19996, A2 => n34108, B1 => n6263, B2 => 
                           n1957, ZN => n1956);
   U13966 : INV_X2 port map( I => n17299, ZN => n783);
   U13970 : XNOR2_X1 port map( A1 => n17300, A2 => n19482, ZN => n17299);
   U13972 : NAND2_X2 port map( A1 => n32740, A2 => n19535, ZN => n20401);
   U13981 : AOI21_X1 port map( A1 => n14365, A2 => n3944, B => n20509, ZN => 
                           n19841);
   U13986 : INV_X2 port map( I => n15282, ZN => n20509);
   U13987 : AOI21_X2 port map( A1 => n19832, A2 => n8406, B => n19831, ZN => 
                           n15282);
   U13988 : AOI21_X2 port map( A1 => n27501, A2 => n738, B => n9934, ZN => 
                           n14690);
   U13989 : NAND2_X2 port map( A1 => n3748, A2 => n24120, ZN => n10427);
   U13992 : OR2_X2 port map( A1 => n2978, A2 => n33482, Z => n9852);
   U13994 : XOR2_X1 port map( A1 => n24492, A2 => n24693, Z => n15862);
   U14000 : XOR2_X1 port map( A1 => n15671, A2 => n15508, Z => n24492);
   U14003 : INV_X2 port map( I => n27127, ZN => n1079);
   U14005 : INV_X2 port map( I => n25277, ZN => n25284);
   U14007 : NAND3_X2 port map( A1 => n24588, A2 => n10330, A3 => n24585, ZN => 
                           n25277);
   U14009 : NOR2_X1 port map( A1 => n18874, A2 => n9909, ZN => n14666);
   U14010 : NAND2_X1 port map( A1 => n32938, A2 => n33803, ZN => n23730);
   U14012 : NAND3_X2 port map( A1 => n11629, A2 => n33046, A3 => n2066, ZN => 
                           n22415);
   U14013 : OR2_X1 port map( A1 => n9931, A2 => n7663, Z => n33560);
   U14019 : NOR3_X1 port map( A1 => n31702, A2 => n30783, A3 => n21086, ZN => 
                           n32741);
   U14026 : NOR2_X2 port map( A1 => n27687, A2 => n30271, ZN => n18472);
   U14027 : NOR2_X2 port map( A1 => n4225, A2 => n8285, ZN => n21044);
   U14034 : XOR2_X1 port map( A1 => n32742, A2 => n23213, Z => n284);
   U14036 : XOR2_X1 port map( A1 => n102, A2 => n27763, Z => n32742);
   U14041 : AOI22_X2 port map( A1 => n32743, A2 => n28867, B1 => n5178, B2 => 
                           n5177, ZN => n26767);
   U14042 : NOR2_X2 port map( A1 => n5178, A2 => n28330, ZN => n32743);
   U14046 : NOR2_X2 port map( A1 => n20038, A2 => n20135, ZN => n19964);
   U14048 : NAND2_X2 port map( A1 => n27911, A2 => n20037, ZN => n20038);
   U14049 : XOR2_X1 port map( A1 => n7636, A2 => n7634, Z => n33856);
   U14053 : XOR2_X1 port map( A1 => n19586, A2 => n11817, Z => n7636);
   U14055 : NOR2_X2 port map( A1 => n20453, A2 => n20454, ZN => n16959);
   U14056 : NAND2_X2 port map( A1 => n15176, A2 => n15177, ZN => n20453);
   U14057 : XOR2_X1 port map( A1 => n12376, A2 => n1917, Z => n17128);
   U14064 : XOR2_X1 port map( A1 => n8949, A2 => n24837, Z => n15308);
   U14066 : NOR2_X2 port map( A1 => n10793, A2 => n24172, ZN => n8949);
   U14067 : XOR2_X1 port map( A1 => n20983, A2 => n20686, Z => n15526);
   U14070 : NAND2_X1 port map( A1 => n8927, A2 => n15602, ZN => n11770);
   U14072 : AND2_X1 port map( A1 => n21253, A2 => n21233, Z => n33263);
   U14073 : NAND2_X2 port map( A1 => n12658, A2 => n23901, ZN => n31275);
   U14076 : AOI22_X2 port map( A1 => n26257, A2 => n16959, B1 => n28527, B2 => 
                           n20362, ZN => n28332);
   U14080 : NAND2_X2 port map( A1 => n31960, A2 => n11755, ZN => n10775);
   U14083 : NAND2_X2 port map( A1 => n22358, A2 => n22357, ZN => n22986);
   U14085 : NAND2_X2 port map( A1 => n22510, A2 => n8199, ZN => n22358);
   U14088 : XOR2_X1 port map( A1 => n32744, A2 => n1421, Z => Ciphertext(150));
   U14090 : AOI22_X1 port map( A1 => n1076, A2 => n9552, B1 => n4253, B2 => 
                           n9495, ZN => n32744);
   U14099 : INV_X2 port map( I => n245, ZN => n32745);
   U14100 : NOR2_X1 port map( A1 => n6118, A2 => n18795, ZN => n8315);
   U14101 : XOR2_X1 port map( A1 => n24455, A2 => n24788, Z => n391);
   U14103 : XOR2_X1 port map( A1 => n24790, A2 => n24512, Z => n24455);
   U14106 : XOR2_X1 port map( A1 => n23506, A2 => n23504, Z => n2024);
   U14110 : XOR2_X1 port map( A1 => n4400, A2 => n14293, Z => n19537);
   U14114 : NOR2_X2 port map( A1 => n19250, A2 => n19251, ZN => n4400);
   U14117 : NAND2_X2 port map( A1 => n32748, A2 => n5045, ZN => n23792);
   U14118 : OAI21_X2 port map( A1 => n1973, A2 => n3748, B => n5335, ZN => 
                           n32748);
   U14123 : BUF_X2 port map( I => n27931, Z => n32750);
   U14131 : OAI21_X1 port map( A1 => n21854, A2 => n21559, B => n4356, ZN => 
                           n5264);
   U14132 : NAND2_X2 port map( A1 => n6878, A2 => n6880, ZN => n4356);
   U14134 : NOR2_X2 port map( A1 => n8671, A2 => n32751, ZN => n14331);
   U14136 : NAND3_X2 port map( A1 => n15696, A2 => n18074, A3 => n9512, ZN => 
                           n32751);
   U14142 : NAND2_X2 port map( A1 => n27139, A2 => n17746, ZN => n3487);
   U14144 : AOI22_X2 port map( A1 => n9660, A2 => n937, B1 => n13423, B2 => 
                           n29283, ZN => n17746);
   U14146 : OAI21_X2 port map( A1 => n32752, A2 => n31167, B => n29738, ZN => 
                           n19325);
   U14148 : NOR2_X2 port map( A1 => n9289, A2 => n18671, ZN => n32752);
   U14150 : XOR2_X1 port map( A1 => n14645, A2 => n27167, Z => n3235);
   U14153 : NOR2_X2 port map( A1 => n1997, A2 => n1995, ZN => n27167);
   U14154 : AOI22_X2 port map( A1 => n26301, A2 => n9913, B1 => n13143, B2 => 
                           n11917, ZN => n32754);
   U14156 : BUF_X4 port map( I => n21867, Z => n30152);
   U14158 : XOR2_X1 port map( A1 => n32755, A2 => n24503, Z => n16659);
   U14159 : XOR2_X1 port map( A1 => n10632, A2 => n24241, Z => n32755);
   U14160 : NAND2_X2 port map( A1 => n22613, A2 => n32756, ZN => n16022);
   U14165 : AOI21_X2 port map( A1 => n32045, A2 => n26173, B => n32757, ZN => 
                           n32756);
   U14175 : XOR2_X1 port map( A1 => n13695, A2 => n24479, Z => n14499);
   U14176 : NAND2_X2 port map( A1 => n9398, A2 => n9933, ZN => n13695);
   U14178 : NOR2_X2 port map( A1 => n20312, A2 => n26566, ZN => n20480);
   U14182 : XOR2_X1 port map( A1 => n12972, A2 => n18929, Z => n10861);
   U14185 : XOR2_X1 port map( A1 => n2162, A2 => n2161, Z => n2655);
   U14186 : XOR2_X1 port map( A1 => n22220, A2 => n8617, Z => n13020);
   U14191 : OAI21_X2 port map( A1 => n16371, A2 => n8618, B => n21739, ZN => 
                           n22220);
   U14193 : NAND3_X2 port map( A1 => n16962, A2 => n22415, A3 => n22416, ZN => 
                           n15456);
   U14197 : NAND2_X2 port map( A1 => n6380, A2 => n31428, ZN => n34065);
   U14198 : XOR2_X1 port map( A1 => n20869, A2 => n25457, Z => n2055);
   U14201 : NAND2_X2 port map( A1 => n26632, A2 => n13000, ZN => n20869);
   U14205 : NAND2_X2 port map( A1 => n20312, A2 => n20577, ZN => n20243);
   U14209 : AOI22_X1 port map( A1 => n6807, A2 => n29234, B1 => n32800, B2 => 
                           n27532, ZN => n14308);
   U14210 : NOR2_X2 port map( A1 => n21636, A2 => n21634, ZN => n32800);
   U14211 : INV_X2 port map( I => n28950, ZN => n32760);
   U14215 : NAND2_X2 port map( A1 => n10, A2 => n32762, ZN => n14342);
   U14216 : NAND3_X2 port map( A1 => n14346, A2 => n18637, A3 => n14651, ZN => 
                           n32762);
   U14218 : AOI21_X2 port map( A1 => n28671, A2 => n23760, B => n23756, ZN => 
                           n4026);
   U14221 : NAND2_X2 port map( A1 => n33837, A2 => n32763, ZN => n18974);
   U14223 : XNOR2_X1 port map( A1 => n29042, A2 => n20747, ZN => n20958);
   U14226 : NAND2_X2 port map( A1 => n183, A2 => n7956, ZN => n20747);
   U14227 : AOI21_X2 port map( A1 => n13104, A2 => n13105, B => n22112, ZN => 
                           n22894);
   U14230 : AOI22_X2 port map( A1 => n32764, A2 => n27386, B1 => n13943, B2 => 
                           n20358, ZN => n20963);
   U14234 : OR2_X1 port map( A1 => n7762, A2 => n27600, Z => n32765);
   U14235 : NAND2_X2 port map( A1 => n8968, A2 => n24109, ZN => n28253);
   U14239 : INV_X1 port map( I => n13063, ZN => n32766);
   U14240 : NAND2_X1 port map( A1 => n33023, A2 => n32766, ZN => n5092);
   U14246 : XOR2_X1 port map( A1 => n32767, A2 => n33877, Z => n14439);
   U14248 : XOR2_X1 port map( A1 => n6218, A2 => n6808, Z => n32767);
   U14250 : NAND2_X1 port map( A1 => n33657, A2 => n2911, ZN => n33656);
   U14258 : OAI22_X2 port map( A1 => n21453, A2 => n1143, B1 => n9186, B2 => 
                           n21237, ZN => n33586);
   U14259 : INV_X2 port map( I => n32768, ZN => n29882);
   U14260 : XOR2_X1 port map( A1 => n2054, A2 => n2053, Z => n32768);
   U14261 : AOI21_X2 port map( A1 => n32769, A2 => n33324, B => n15984, ZN => 
                           n19021);
   U14265 : INV_X2 port map( I => n9810, ZN => n9440);
   U14267 : XOR2_X1 port map( A1 => n22306, A2 => n9809, Z => n9810);
   U14268 : NOR2_X1 port map( A1 => n10018, A2 => n3004, ZN => n2560);
   U14269 : NAND2_X2 port map( A1 => n5795, A2 => n21721, ZN => n21806);
   U14270 : NAND3_X2 port map( A1 => n3936, A2 => n10555, A3 => n4179, ZN => 
                           n5795);
   U14275 : NOR2_X2 port map( A1 => n16637, A2 => n1042, ZN => n19903);
   U14277 : OR2_X1 port map( A1 => n10312, A2 => n8057, Z => n19864);
   U14278 : XOR2_X1 port map( A1 => n24812, A2 => n32770, Z => n26365);
   U14281 : XOR2_X1 port map( A1 => n9650, A2 => n24811, Z => n32770);
   U14282 : NAND3_X2 port map( A1 => n21187, A2 => n17640, A3 => n34131, ZN => 
                           n21083);
   U14285 : NAND2_X2 port map( A1 => n5394, A2 => n5395, ZN => n21187);
   U14286 : OAI21_X2 port map( A1 => n33030, A2 => n14276, B => n16728, ZN => 
                           n14274);
   U14290 : OR2_X1 port map( A1 => n31969, A2 => n10312, Z => n31338);
   U14295 : XOR2_X1 port map( A1 => n29624, A2 => n14340, Z => n21232);
   U14297 : AOI21_X2 port map( A1 => n29695, A2 => n20489, B => n20487, ZN => 
                           n17512);
   U14301 : NOR2_X2 port map( A1 => n13015, A2 => n13845, ZN => n12648);
   U14303 : XOR2_X1 port map( A1 => n19642, A2 => n32058, Z => n582);
   U14308 : XOR2_X1 port map( A1 => n32772, A2 => n15679, Z => n32915);
   U14310 : XOR2_X1 port map( A1 => n17220, A2 => n32044, Z => n32772);
   U14311 : XOR2_X1 port map( A1 => n19710, A2 => n19408, Z => n15913);
   U14312 : NOR2_X1 port map( A1 => n12932, A2 => n9146, ZN => n27309);
   U14313 : NOR2_X2 port map( A1 => n17329, A2 => n4647, ZN => n15045);
   U14317 : OAI21_X1 port map( A1 => n22413, A2 => n14160, B => n22486, ZN => 
                           n14010);
   U14320 : XOR2_X1 port map( A1 => n12934, A2 => n23435, Z => n23155);
   U14321 : XOR2_X1 port map( A1 => n24554, A2 => n24556, Z => n1690);
   U14334 : XOR2_X1 port map( A1 => n24846, A2 => n24741, Z => n24554);
   U14335 : INV_X2 port map( I => n25345, ZN => n14246);
   U14339 : NAND2_X2 port map( A1 => n18958, A2 => n18621, ZN => n18962);
   U14343 : XOR2_X1 port map( A1 => n21012, A2 => n21011, Z => n7015);
   U14354 : XOR2_X1 port map( A1 => n15293, A2 => n13930, Z => n30734);
   U14359 : NAND2_X2 port map( A1 => n29464, A2 => n10349, ZN => n15293);
   U14360 : NAND2_X2 port map( A1 => n5428, A2 => n32773, ZN => n8335);
   U14361 : OAI21_X2 port map( A1 => n18750, A2 => n13243, B => n959, ZN => 
                           n32773);
   U14362 : NAND3_X2 port map( A1 => n23002, A2 => n22831, A3 => n13159, ZN => 
                           n12157);
   U14368 : XOR2_X1 port map( A1 => n1994, A2 => n28601, Z => n6913);
   U14369 : XOR2_X1 port map( A1 => n32774, A2 => n590, Z => n21053);
   U14370 : XOR2_X1 port map( A1 => n21026, A2 => n20855, Z => n32774);
   U14375 : AOI22_X2 port map( A1 => n32775, A2 => n8183, B1 => n20060, B2 => 
                           n16789, ZN => n29914);
   U14378 : INV_X1 port map( I => n4327, ZN => n32776);
   U14384 : NAND2_X1 port map( A1 => n27955, A2 => n21396, ZN => n32778);
   U14386 : NAND2_X2 port map( A1 => n9677, A2 => n10228, ZN => n11798);
   U14400 : NAND2_X2 port map( A1 => n30246, A2 => n32779, ZN => n7182);
   U14401 : NAND2_X1 port map( A1 => n3888, A2 => n3889, ZN => n32779);
   U14402 : BUF_X2 port map( I => n20080, Z => n32780);
   U14405 : OAI21_X2 port map( A1 => n31463, A2 => n31464, B => n25872, ZN => 
                           n13053);
   U14408 : INV_X2 port map( I => n32781, ZN => n29444);
   U14413 : NAND2_X2 port map( A1 => n14054, A2 => n8130, ZN => n32781);
   U14416 : XOR2_X1 port map( A1 => n32782, A2 => n25856, Z => Ciphertext(177))
                           ;
   U14422 : XOR2_X1 port map( A1 => n32783, A2 => n465, Z => n6420);
   U14424 : XOR2_X1 port map( A1 => n30524, A2 => n16373, Z => n32783);
   U14427 : INV_X2 port map( I => n28278, ZN => n1322);
   U14428 : INV_X2 port map( I => n32784, ZN => n18920);
   U14430 : NAND3_X2 port map( A1 => n18833, A2 => n32786, A3 => n32785, ZN => 
                           n32784);
   U14434 : NOR3_X1 port map( A1 => n27262, A2 => n1202, A3 => n32856, ZN => 
                           n27528);
   U14436 : OR2_X1 port map( A1 => n16606, A2 => n20566, Z => n33937);
   U14437 : OR3_X1 port map( A1 => n28430, A2 => n20008, A3 => n29882, Z => 
                           n1873);
   U14443 : XOR2_X1 port map( A1 => n9507, A2 => n20976, Z => n2812);
   U14450 : INV_X2 port map( I => n15516, ZN => n9507);
   U14453 : XOR2_X1 port map( A1 => n21009, A2 => n20873, Z => n15516);
   U14455 : NAND2_X2 port map( A1 => n32789, A2 => n3780, ZN => n18028);
   U14461 : BUF_X2 port map( I => n33373, Z => n32791);
   U14463 : NAND2_X2 port map( A1 => n32792, A2 => n16978, ZN => n20565);
   U14472 : NAND2_X2 port map( A1 => n32793, A2 => n18270, ZN => n21028);
   U14474 : OAI22_X2 port map( A1 => n27901, A2 => n27902, B1 => n8819, B2 => 
                           n12999, ZN => n32793);
   U14476 : NAND2_X2 port map( A1 => n32794, A2 => n13106, ZN => n3055);
   U14477 : NAND2_X2 port map( A1 => n3057, A2 => n5139, ZN => n13106);
   U14482 : OR2_X1 port map( A1 => n3060, A2 => n3059, Z => n32794);
   U14486 : XOR2_X1 port map( A1 => n33427, A2 => n1540, Z => n11720);
   U14495 : XOR2_X1 port map( A1 => n20889, A2 => n32795, Z => n27000);
   U14496 : XOR2_X1 port map( A1 => n10159, A2 => n32796, Z => n32795);
   U14499 : XOR2_X1 port map( A1 => n28587, A2 => n15424, Z => n27234);
   U14501 : NAND2_X2 port map( A1 => n7881, A2 => n23065, ZN => n22827);
   U14503 : NOR3_X2 port map( A1 => n29455, A2 => n31073, A3 => n16722, ZN => 
                           n21913);
   U14505 : NOR2_X1 port map( A1 => n7993, A2 => n28329, ZN => n5678);
   U14506 : NOR2_X1 port map( A1 => n1773, A2 => n22551, ZN => n22314);
   U14509 : NAND3_X2 port map( A1 => n24233, A2 => n1634, A3 => n24236, ZN => 
                           n23699);
   U14512 : XOR2_X1 port map( A1 => n29137, A2 => n9412, Z => n17395);
   U14518 : AOI22_X2 port map( A1 => n1771, A2 => n1770, B1 => n1769, B2 => 
                           n2551, ZN => n9412);
   U14523 : XOR2_X1 port map( A1 => n20743, A2 => n1545, Z => n7431);
   U14524 : XOR2_X1 port map( A1 => n3009, A2 => n21047, Z => n20743);
   U14525 : OAI22_X2 port map( A1 => n20288, A2 => n10351, B1 => n20324, B2 => 
                           n20519, ZN => n7255);
   U14529 : XOR2_X1 port map( A1 => n9701, A2 => n33678, Z => n22597);
   U14532 : BUF_X4 port map( I => n18655, Z => n17843);
   U14538 : AND2_X1 port map( A1 => n10847, A2 => n8870, Z => n30004);
   U14548 : XOR2_X1 port map( A1 => n18100, A2 => n22191, Z => n6515);
   U14551 : NAND2_X2 port map( A1 => n11359, A2 => n11728, ZN => n22191);
   U14556 : BUF_X2 port map( I => n32069, Z => n32799);
   U14557 : NAND2_X2 port map( A1 => n22497, A2 => n16306, ZN => n33010);
   U14560 : OAI22_X2 port map( A1 => n22762, A2 => n22715, B1 => n22694, B2 => 
                           n851, ZN => n33008);
   U14565 : XOR2_X1 port map( A1 => n17369, A2 => n16429, Z => n18929);
   U14566 : OR2_X1 port map( A1 => n18098, A2 => n22476, Z => n30384);
   U14568 : XOR2_X1 port map( A1 => n14215, A2 => n19475, Z => n11092);
   U14570 : XOR2_X1 port map( A1 => n14214, A2 => n19367, Z => n14215);
   U14573 : OAI22_X2 port map( A1 => n12509, A2 => n32801, B1 => n23448, B2 => 
                           n28210, ZN => n16215);
   U14575 : BUF_X2 port map( I => n19325, Z => n32802);
   U14581 : INV_X2 port map( I => n32803, ZN => n4145);
   U14588 : XOR2_X1 port map( A1 => n33916, A2 => n1704, Z => n32803);
   U14589 : XOR2_X1 port map( A1 => n32804, A2 => n19575, Z => n13305);
   U14593 : XOR2_X1 port map( A1 => n26617, A2 => n8633, Z => n32804);
   U14602 : XOR2_X1 port map( A1 => n17351, A2 => n17350, Z => n33152);
   U14603 : XOR2_X1 port map( A1 => n4728, A2 => n31843, Z => n5523);
   U14604 : NAND2_X2 port map( A1 => n11266, A2 => n11265, ZN => n21559);
   U14605 : NAND2_X2 port map( A1 => n2355, A2 => n33664, ZN => n22283);
   U14606 : OAI21_X2 port map( A1 => n375, A2 => n29040, B => n20092, ZN => 
                           n31280);
   U14608 : NAND2_X2 port map( A1 => n33286, A2 => n9691, ZN => n14639);
   U14610 : XOR2_X1 port map( A1 => n26255, A2 => n11636, Z => n31575);
   U14611 : XOR2_X1 port map( A1 => n33111, A2 => n23219, Z => n15487);
   U14612 : XOR2_X1 port map( A1 => n20912, A2 => n7458, Z => n26954);
   U14615 : XOR2_X1 port map( A1 => n8997, A2 => n20781, Z => n7458);
   U14616 : NOR3_X2 port map( A1 => n33985, A2 => n4117, A3 => n7349, ZN => 
                           n7348);
   U14622 : XOR2_X1 port map( A1 => n29936, A2 => n30676, Z => n13427);
   U14627 : XOR2_X1 port map( A1 => n21027, A2 => n21026, Z => n12272);
   U14632 : NAND2_X2 port map( A1 => n7007, A2 => n28190, ZN => n10149);
   U14638 : AND2_X1 port map( A1 => n25891, A2 => n25890, Z => n33473);
   U14640 : NAND2_X2 port map( A1 => n32806, A2 => n15631, ZN => n7868);
   U14642 : OAI21_X2 port map( A1 => n30694, A2 => n10483, B => n926, ZN => 
                           n32806);
   U14644 : NOR2_X2 port map( A1 => n32108, A2 => n33621, ZN => n18800);
   U14646 : OR2_X1 port map( A1 => n17131, A2 => n17130, Z => n28361);
   U14648 : OAI22_X2 port map( A1 => n11049, A2 => n23608, B1 => n24285, B2 => 
                           n17068, ZN => n27793);
   U14649 : XOR2_X1 port map( A1 => n14762, A2 => n24826, Z => n24808);
   U14650 : NAND2_X2 port map( A1 => n29924, A2 => n2401, ZN => n14762);
   U14656 : NAND2_X2 port map( A1 => n2036, A2 => n32843, ZN => n27931);
   U14664 : OAI22_X2 port map( A1 => n33567, A2 => n33568, B1 => n9945, B2 => 
                           n10416, ZN => n12720);
   U14666 : NAND2_X1 port map( A1 => n11379, A2 => n14898, ZN => n3436);
   U14668 : NAND2_X1 port map( A1 => n26330, A2 => n22634, ZN => n22612);
   U14669 : NOR2_X1 port map( A1 => n33283, A2 => n858, ZN => n33282);
   U14675 : NAND2_X1 port map( A1 => n33282, A2 => n33280, ZN => n33901);
   U14681 : NAND2_X2 port map( A1 => n12358, A2 => n25890, ZN => n30019);
   U14684 : XOR2_X1 port map( A1 => n3576, A2 => n3574, Z => n18182);
   U14685 : XOR2_X1 port map( A1 => n32810, A2 => n24553, Z => n9189);
   U14688 : OAI21_X2 port map( A1 => n18127, A2 => n18128, B => n24227, ZN => 
                           n24553);
   U14690 : INV_X2 port map( I => n24847, ZN => n32810);
   U14692 : BUF_X4 port map( I => n15296, Z => n29180);
   U14702 : OAI22_X2 port map( A1 => n32601, A2 => n25205, B1 => n13273, B2 => 
                           n25239, ZN => n33494);
   U14706 : NAND2_X1 port map( A1 => n10287, A2 => n33566, ZN => n4341);
   U14710 : XOR2_X1 port map( A1 => n12272, A2 => n21032, Z => n33566);
   U14711 : NAND2_X2 port map( A1 => n21674, A2 => n16345, ZN => n28111);
   U14713 : NAND2_X2 port map( A1 => n33810, A2 => n21604, ZN => n21674);
   U14719 : XOR2_X1 port map( A1 => n31486, A2 => n32811, Z => n28107);
   U14720 : XOR2_X1 port map( A1 => n30628, A2 => n21996, Z => n32811);
   U14724 : XOR2_X1 port map( A1 => n7107, A2 => n32812, Z => n31737);
   U14725 : XOR2_X1 port map( A1 => n34100, A2 => n32813, Z => n32812);
   U14728 : INV_X1 port map( I => n25541, ZN => n32813);
   U14733 : NOR2_X2 port map( A1 => n25165, A2 => n25175, ZN => n25173);
   U14735 : CLKBUF_X8 port map( I => n13473, Z => n33007);
   U14739 : NAND2_X2 port map( A1 => n29043, A2 => n8125, ZN => n421);
   U14740 : XOR2_X1 port map( A1 => n8067, A2 => n8065, Z => n9490);
   U14743 : NAND3_X2 port map( A1 => n31933, A2 => n1117, A3 => n7561, ZN => 
                           n27856);
   U14751 : NAND3_X2 port map( A1 => n17532, A2 => n20489, A3 => n4254, ZN => 
                           n7799);
   U14753 : OR2_X1 port map( A1 => n19101, A2 => n18923, Z => n17444);
   U14754 : NOR2_X1 port map( A1 => n10103, A2 => n10104, ZN => n33601);
   U14763 : BUF_X2 port map( I => n13286, Z => n32816);
   U14768 : NAND2_X2 port map( A1 => n14959, A2 => n25013, ZN => n14846);
   U14774 : NAND2_X2 port map( A1 => n15277, A2 => n14799, ZN => n33288);
   U14776 : XOR2_X1 port map( A1 => n32817, A2 => n1198, Z => Ciphertext(138));
   U14778 : AOI22_X1 port map( A1 => n28631, A2 => n11212, B1 => n9365, B2 => 
                           n734, ZN => n32817);
   U14782 : NAND2_X2 port map( A1 => n33304, A2 => n28194, ZN => n16286);
   U14792 : XOR2_X1 port map( A1 => n15691, A2 => n32818, Z => n26630);
   U14793 : XOR2_X1 port map( A1 => n23504, A2 => n15690, Z => n32818);
   U14795 : NAND2_X2 port map( A1 => n3379, A2 => n777, ZN => n34084);
   U14796 : OAI22_X2 port map( A1 => n21438, A2 => n21224, B1 => n21223, B2 => 
                           n8398, ZN => n11232);
   U14802 : NAND3_X1 port map( A1 => n16091, A2 => n8045, A3 => n30059, ZN => 
                           n32819);
   U14804 : NOR2_X2 port map( A1 => n8970, A2 => n279, ZN => n32983);
   U14807 : NAND2_X2 port map( A1 => n4289, A2 => n20401, ZN => n31079);
   U14808 : XOR2_X1 port map( A1 => n10758, A2 => n23164, Z => n4446);
   U14811 : XOR2_X1 port map( A1 => n23441, A2 => n23211, Z => n23164);
   U14812 : INV_X2 port map( I => n28374, ZN => n26806);
   U14813 : NAND2_X2 port map( A1 => n32821, A2 => n23802, ZN => n28374);
   U14818 : AND2_X1 port map( A1 => n23803, A2 => n23801, Z => n32821);
   U14819 : XOR2_X1 port map( A1 => n19772, A2 => n19399, Z => n19733);
   U14821 : NAND2_X2 port map( A1 => n8576, A2 => n8857, ZN => n9106);
   U14831 : OR2_X1 port map( A1 => n26448, A2 => n21258, Z => n33683);
   U14832 : NOR2_X2 port map( A1 => n9195, A2 => n25701, ZN => n25766);
   U14833 : NAND2_X1 port map( A1 => n16170, A2 => n25, ZN => n2258);
   U14841 : OR2_X1 port map( A1 => n29342, A2 => n22398, Z => n33190);
   U14844 : BUF_X2 port map( I => n2483, Z => n32822);
   U14846 : XOR2_X1 port map( A1 => n24528, A2 => n549, Z => n28746);
   U14847 : XOR2_X1 port map( A1 => n4662, A2 => n4661, Z => n16536);
   U14854 : XOR2_X1 port map( A1 => n32824, A2 => n23239, Z => Ciphertext(75));
   U14857 : NAND3_X2 port map( A1 => n10942, A2 => n32990, A3 => n10940, ZN => 
                           n32824);
   U14858 : XOR2_X1 port map( A1 => n15877, A2 => n10159, Z => n30985);
   U14860 : XOR2_X1 port map( A1 => n31899, A2 => n10729, Z => n5229);
   U14862 : INV_X4 port map( I => n25235, ZN => n34115);
   U14867 : XOR2_X1 port map( A1 => n23137, A2 => n23532, Z => n23219);
   U14870 : OAI21_X2 port map( A1 => n11064, A2 => n10687, B => n28467, ZN => 
                           n10811);
   U14872 : OAI22_X2 port map( A1 => n32826, A2 => n2773, B1 => n2775, B2 => 
                           n11317, ZN => n3519);
   U14877 : NAND2_X2 port map( A1 => n4967, A2 => n14055, ZN => n32828);
   U14879 : NAND2_X2 port map( A1 => n29334, A2 => n15318, ZN => n4967);
   U14881 : OAI21_X1 port map( A1 => n5492, A2 => n24996, B => n7940, ZN => 
                           n9478);
   U14882 : NAND2_X2 port map( A1 => n28647, A2 => n19530, ZN => n28108);
   U14884 : NAND2_X2 port map( A1 => n3266, A2 => n11967, ZN => n28523);
   U14885 : NOR2_X2 port map( A1 => n1940, A2 => n1233, ZN => n32829);
   U14886 : NAND2_X2 port map( A1 => n15253, A2 => n13472, ZN => n6354);
   U14888 : XOR2_X1 port map( A1 => n31727, A2 => n16705, Z => n12924);
   U14890 : INV_X2 port map( I => n11845, ZN => n24316);
   U14891 : OAI22_X1 port map( A1 => n23946, A2 => n30359, B1 => n11676, B2 => 
                           n10187, ZN => n8675);
   U14892 : OAI22_X2 port map( A1 => n15225, A2 => n20381, B1 => n15162, B2 => 
                           n20633, ZN => n11241);
   U14898 : NAND2_X2 port map( A1 => n20445, A2 => n20384, ZN => n20633);
   U14901 : BUF_X2 port map( I => n19901, Z => n8421);
   U14906 : XOR2_X1 port map( A1 => n20930, A2 => n20929, Z => n33673);
   U14908 : NAND3_X2 port map( A1 => n16235, A2 => n30152, A3 => n32832, ZN => 
                           n21588);
   U14909 : INV_X2 port map( I => n21866, ZN => n32833);
   U14910 : XOR2_X1 port map( A1 => n32516, A2 => n25098, Z => n23398);
   U14916 : OAI21_X2 port map( A1 => n21254, A2 => n32644, B => n32834, ZN => 
                           n29854);
   U14923 : AOI22_X2 port map( A1 => n15932, A2 => n9699, B1 => n15931, B2 => 
                           n27462, ZN => n32834);
   U14926 : BUF_X2 port map( I => n22979, Z => n27814);
   U14927 : BUF_X4 port map( I => n16568, Z => n330);
   U14934 : XOR2_X1 port map( A1 => n19637, A2 => n8633, Z => n19433);
   U14936 : NAND2_X2 port map( A1 => n14697, A2 => n19246, ZN => n19637);
   U14937 : BUF_X4 port map( I => n23904, Z => n6414);
   U14938 : XOR2_X1 port map( A1 => n22171, A2 => n3781, Z => n175);
   U14939 : XOR2_X1 port map( A1 => n30999, A2 => n22211, Z => n3781);
   U14944 : NAND2_X2 port map( A1 => n16421, A2 => n8434, ZN => n20780);
   U14945 : NAND3_X1 port map( A1 => n31103, A2 => n29250, A3 => n19808, ZN => 
                           n19809);
   U14950 : OAI22_X2 port map( A1 => n14725, A2 => n27104, B1 => n31228, B2 => 
                           n2798, ZN => n24383);
   U14953 : NAND2_X2 port map( A1 => n31218, A2 => n7893, ZN => n7892);
   U14954 : OAI21_X2 port map( A1 => n3224, A2 => n1213, B => n33493, ZN => 
                           n3223);
   U14967 : XOR2_X1 port map( A1 => n13455, A2 => n13456, Z => n27257);
   U14970 : NAND2_X1 port map( A1 => n28657, A2 => n28655, ZN => n10823);
   U14976 : NAND2_X1 port map( A1 => n4733, A2 => n14056, ZN => n18625);
   U14978 : NAND2_X2 port map( A1 => n26962, A2 => n16564, ZN => n4733);
   U14984 : AND2_X1 port map( A1 => n21426, A2 => n13286, Z => n33418);
   U14986 : XOR2_X1 port map( A1 => n7597, A2 => n7599, Z => n22598);
   U14987 : XOR2_X1 port map( A1 => n14277, A2 => n31552, Z => n675);
   U14988 : XOR2_X1 port map( A1 => n17798, A2 => n24494, Z => n10685);
   U14994 : XOR2_X1 port map( A1 => n24811, A2 => n24553, Z => n24494);
   U15001 : NAND3_X2 port map( A1 => n23711, A2 => n23709, A3 => n23710, ZN => 
                           n12981);
   U15017 : BUF_X2 port map( I => n17338, Z => n31850);
   U15020 : XOR2_X1 port map( A1 => n32835, A2 => n13899, Z => n21198);
   U15022 : XOR2_X1 port map( A1 => n32892, A2 => n13898, Z => n32835);
   U15026 : AOI22_X2 port map( A1 => n17139, A2 => n28429, B1 => n30506, B2 => 
                           n28450, ZN => n21488);
   U15030 : OAI21_X2 port map( A1 => n5377, A2 => n5376, B => n26516, ZN => 
                           n32836);
   U15031 : NAND2_X2 port map( A1 => n17561, A2 => n4349, ZN => n24095);
   U15033 : AND2_X1 port map( A1 => n25563, A2 => n28093, Z => n25520);
   U15034 : INV_X1 port map( I => n30252, ZN => n33813);
   U15039 : AND2_X1 port map( A1 => n30252, A2 => n23833, Z => n33812);
   U15044 : INV_X1 port map( I => n17280, ZN => n31801);
   U15057 : NOR2_X2 port map( A1 => n2209, A2 => n25686, ZN => n14732);
   U15059 : NAND2_X2 port map( A1 => n715, A2 => n28651, ZN => n14795);
   U15060 : NOR2_X1 port map( A1 => n32837, A2 => n27007, ZN => n11566);
   U15061 : NAND2_X2 port map( A1 => n13535, A2 => n30631, ZN => n27007);
   U15065 : AOI21_X2 port map( A1 => n23601, A2 => n5357, B => n27049, ZN => 
                           n14548);
   U15077 : XOR2_X1 port map( A1 => n6329, A2 => n32838, Z => n32924);
   U15089 : INV_X2 port map( I => n522, ZN => n32926);
   U15091 : XOR2_X1 port map( A1 => n19558, A2 => n19755, Z => n19611);
   U15094 : NAND3_X2 port map( A1 => n18526, A2 => n18527, A3 => n18528, ZN => 
                           n19755);
   U15095 : NOR2_X2 port map( A1 => n5704, A2 => n7592, ZN => n21711);
   U15098 : XOR2_X1 port map( A1 => n602, A2 => n2756, Z => n4327);
   U15099 : XOR2_X1 port map( A1 => n29832, A2 => n20684, Z => n602);
   U15101 : XOR2_X1 port map( A1 => n20956, A2 => n32839, Z => n29303);
   U15103 : XOR2_X1 port map( A1 => n27054, A2 => n20896, Z => n32839);
   U15110 : NAND2_X2 port map( A1 => n15344, A2 => n32840, ZN => n34004);
   U15111 : NAND2_X2 port map( A1 => n25592, A2 => n9862, ZN => n388);
   U15113 : INV_X4 port map( I => n9219, ZN => n24292);
   U15118 : OAI21_X2 port map( A1 => n2325, A2 => n32323, B => n24127, ZN => 
                           n34093);
   U15120 : XOR2_X1 port map( A1 => n32841, A2 => n23264, Z => n27667);
   U15122 : NOR2_X2 port map( A1 => n16922, A2 => n22743, ZN => n23395);
   U15129 : BUF_X4 port map( I => n29321, Z => n33992);
   U15131 : XOR2_X1 port map( A1 => n19686, A2 => n32844, Z => n19586);
   U15132 : INV_X2 port map( I => n19341, ZN => n32844);
   U15135 : NAND2_X1 port map( A1 => n33853, A2 => n29568, ZN => n14838);
   U15138 : INV_X2 port map( I => n13073, ZN => n21414);
   U15139 : NOR2_X1 port map( A1 => n29322, A2 => n6176, ZN => n2219);
   U15141 : INV_X2 port map( I => n6275, ZN => n16848);
   U15142 : NAND2_X1 port map( A1 => n12564, A2 => n33218, ZN => n124);
   U15143 : NOR2_X1 port map( A1 => n32852, A2 => n9480, ZN => n27968);
   U15154 : NOR2_X1 port map( A1 => n9052, A2 => n33643, ZN => n27099);
   U15172 : OAI21_X1 port map( A1 => n25053, A2 => n27610, B => n32845, ZN => 
                           n25055);
   U15174 : AOI22_X1 port map( A1 => n17728, A2 => n25062, B1 => n17729, B2 => 
                           n27610, ZN => n32845);
   U15177 : NAND2_X2 port map( A1 => n27624, A2 => n1164, ZN => n10272);
   U15178 : OAI21_X2 port map( A1 => n31822, A2 => n25890, B => n30811, ZN => 
                           n31378);
   U15182 : NAND2_X2 port map( A1 => n22655, A2 => n22951, ZN => n22952);
   U15185 : NAND2_X2 port map( A1 => n22258, A2 => n6540, ZN => n22655);
   U15187 : OAI21_X2 port map( A1 => n10221, A2 => n6981, B => n1223, ZN => 
                           n33197);
   U15188 : XOR2_X1 port map( A1 => n32846, A2 => n30156, Z => n31650);
   U15190 : XOR2_X1 port map( A1 => n23123, A2 => n23124, Z => n32846);
   U15192 : XOR2_X1 port map( A1 => n21995, A2 => n22282, Z => n15727);
   U15193 : XOR2_X1 port map( A1 => n33150, A2 => n22255, Z => n21995);
   U15200 : INV_X2 port map( I => n11805, ZN => n33739);
   U15205 : AOI21_X2 port map( A1 => n6802, A2 => n6675, B => n6674, ZN => 
                           n32860);
   U15206 : XOR2_X1 port map( A1 => n32847, A2 => n25259, Z => Ciphertext(83));
   U15210 : AOI22_X1 port map( A1 => n26497, A2 => n27429, B1 => n8035, B2 => 
                           n8036, ZN => n32847);
   U15215 : NAND2_X2 port map( A1 => n32848, A2 => n5888, ZN => n17236);
   U15221 : NAND2_X1 port map( A1 => n14988, A2 => n28912, ZN => n32848);
   U15223 : NAND2_X1 port map( A1 => n5789, A2 => n28885, ZN => n19205);
   U15224 : OAI22_X2 port map( A1 => n9645, A2 => n843, B1 => n5764, B2 => n548
                           , ZN => n9616);
   U15226 : AOI22_X2 port map( A1 => n10145, A2 => n843, B1 => n9172, B2 => 
                           n11968, ZN => n5764);
   U15227 : NAND3_X2 port map( A1 => n29521, A2 => n15670, A3 => n10066, ZN => 
                           n10469);
   U15231 : NAND2_X2 port map( A1 => n11571, A2 => n15054, ZN => n7871);
   U15234 : OR2_X1 port map( A1 => n33189, A2 => n29230, Z => n34121);
   U15235 : NAND2_X2 port map( A1 => n26903, A2 => n28664, ZN => n33146);
   U15239 : NOR2_X2 port map( A1 => n11695, A2 => n11698, ZN => n25670);
   U15242 : NAND3_X1 port map( A1 => n19292, A2 => n18682, A3 => n746, ZN => 
                           n32849);
   U15247 : XOR2_X1 port map( A1 => n32850, A2 => n29550, Z => n16401);
   U15250 : XOR2_X1 port map( A1 => n572, A2 => n33742, Z => n32850);
   U15252 : OR2_X1 port map( A1 => n14780, A2 => n26447, Z => n25684);
   U15255 : INV_X4 port map( I => n11956, ZN => n28867);
   U15257 : INV_X2 port map( I => n32851, ZN => n34167);
   U15258 : XOR2_X1 port map( A1 => n6848, A2 => n28062, Z => n32851);
   U15260 : XOR2_X1 port map( A1 => n23506, A2 => n23126, Z => n8071);
   U15263 : XOR2_X1 port map( A1 => n29885, A2 => n23293, Z => n23506);
   U15264 : NOR2_X1 port map( A1 => n9479, A2 => n9478, ZN => n32852);
   U15272 : NAND2_X1 port map( A1 => n32853, A2 => n30740, ZN => n7336);
   U15274 : NAND2_X1 port map( A1 => n7341, A2 => n26744, ZN => n32853);
   U15275 : AND3_X1 port map( A1 => n15807, A2 => n21297, A3 => n4989, Z => 
                           n26025);
   U15280 : XOR2_X1 port map( A1 => n5149, A2 => n32854, Z => n19527);
   U15281 : XOR2_X1 port map( A1 => n8561, A2 => n26794, Z => n32854);
   U15284 : BUF_X4 port map( I => n13670, Z => n11187);
   U15285 : OR2_X1 port map( A1 => n26374, A2 => n24340, Z => n24343);
   U15288 : OAI21_X2 port map( A1 => n11757, A2 => n11949, B => n783, ZN => 
                           n33323);
   U15290 : INV_X2 port map( I => n9958, ZN => n14137);
   U15291 : BUF_X4 port map( I => n31721, Z => n33301);
   U15292 : NAND2_X2 port map( A1 => n24933, A2 => n24351, ZN => n17479);
   U15296 : BUF_X4 port map( I => n25051, Z => n31640);
   U15301 : NAND3_X1 port map( A1 => n8766, A2 => n32897, A3 => n33399, ZN => 
                           n4325);
   U15302 : INV_X1 port map( I => n888, ZN => n24101);
   U15305 : NAND3_X1 port map( A1 => n5160, A2 => n24104, A3 => n888, ZN => 
                           n28524);
   U15306 : OAI21_X1 port map( A1 => n24102, A2 => n12098, B => n888, ZN => 
                           n4928);
   U15318 : NAND2_X1 port map( A1 => n24667, A2 => n25536, ZN => n9915);
   U15319 : OAI21_X1 port map( A1 => n24667, A2 => n25536, B => n736, ZN => 
                           n26921);
   U15322 : NOR2_X1 port map( A1 => n8062, A2 => n11200, ZN => n11201);
   U15325 : NAND2_X1 port map( A1 => n3925, A2 => n20142, ZN => n33003);
   U15328 : NAND3_X1 port map( A1 => n10266, A2 => n10265, A3 => n10268, ZN => 
                           n33513);
   U15329 : NOR2_X1 port map( A1 => n26566, A2 => n20577, ZN => n33149);
   U15334 : INV_X1 port map( I => n26566, ZN => n8528);
   U15336 : NOR2_X1 port map( A1 => n6230, A2 => n26566, ZN => n27806);
   U15338 : OAI21_X1 port map( A1 => n29271, A2 => n26415, B => n30125, ZN => 
                           n26221);
   U15344 : OAI21_X1 port map( A1 => n33400, A2 => n33399, B => n1204, ZN => 
                           n33957);
   U15345 : NOR2_X2 port map( A1 => n24888, A2 => n2092, ZN => n28706);
   U15350 : NAND2_X1 port map( A1 => n4243, A2 => n33480, ZN => n24724);
   U15358 : INV_X2 port map( I => n10622, ZN => n998);
   U15359 : NAND2_X1 port map( A1 => n797, A2 => n24150, ZN => n12208);
   U15367 : OAI21_X1 port map( A1 => n797, A2 => n2744, B => n26545, ZN => 
                           n2746);
   U15368 : NOR2_X1 port map( A1 => n10042, A2 => n12423, ZN => n30569);
   U15369 : NAND2_X1 port map( A1 => n1209, A2 => n16798, ZN => n1472);
   U15381 : OR2_X1 port map( A1 => n14490, A2 => n15065, Z => n14491);
   U15382 : AOI22_X1 port map( A1 => n8263, A2 => n14490, B1 => n15818, B2 => 
                           n15996, ZN => n3845);
   U15383 : OAI22_X1 port map( A1 => n24176, A2 => n15790, B1 => n14052, B2 => 
                           n14490, ZN => n3256);
   U15385 : NAND2_X1 port map( A1 => n1007, A2 => n2386, ZN => n33367);
   U15387 : CLKBUF_X2 port map( I => n18818, Z => n16393);
   U15388 : INV_X1 port map( I => n18818, ZN => n18639);
   U15392 : NAND2_X1 port map( A1 => n22883, A2 => n22882, ZN => n33383);
   U15393 : NAND2_X1 port map( A1 => n22883, A2 => n13274, ZN => n3778);
   U15400 : AOI21_X1 port map( A1 => n10045, A2 => n23795, B => n5777, ZN => 
                           n5776);
   U15406 : INV_X2 port map( I => n23795, ZN => n845);
   U15409 : NAND2_X1 port map( A1 => n13698, A2 => n25297, ZN => n33956);
   U15412 : NOR2_X1 port map( A1 => n6869, A2 => n23917, ZN => n4197);
   U15413 : BUF_X1 port map( I => n25546, Z => n8320);
   U15414 : NOR2_X1 port map( A1 => n13334, A2 => n27168, ZN => n6654);
   U15415 : INV_X1 port map( I => n5790, ZN => n11868);
   U15416 : NAND2_X1 port map( A1 => n7501, A2 => n6483, ZN => n33955);
   U15417 : INV_X2 port map( I => n14650, ZN => n25066);
   U15421 : INV_X1 port map( I => n30323, ZN => n29670);
   U15422 : NAND2_X1 port map( A1 => n25568, A2 => n3638, ZN => n10959);
   U15423 : AOI21_X1 port map( A1 => n9022, A2 => n33237, B => n9910, ZN => 
                           n7904);
   U15429 : NOR2_X1 port map( A1 => n20575, A2 => n27785, ZN => n27902);
   U15430 : NAND2_X1 port map( A1 => n1463, A2 => n886, ZN => n1462);
   U15434 : INV_X1 port map( I => n678, ZN => n886);
   U15444 : CLKBUF_X4 port map( I => n18494, Z => n16564);
   U15445 : NOR2_X2 port map( A1 => n23539, A2 => n23538, ZN => n12547);
   U15446 : BUF_X2 port map( I => n4287, Z => n28579);
   U15447 : OAI21_X1 port map( A1 => n23950, A2 => n30359, B => n23620, ZN => 
                           n13774);
   U15455 : AND2_X1 port map( A1 => n13308, A2 => n23949, Z => n23620);
   U15456 : NOR2_X1 port map( A1 => n13698, A2 => n8105, ZN => n15785);
   U15459 : NOR2_X1 port map( A1 => n33460, A2 => n8105, ZN => n15481);
   U15463 : OAI21_X1 port map( A1 => n25537, A2 => n16826, B => n8105, ZN => 
                           n34033);
   U15464 : NOR2_X1 port map( A1 => n33480, A2 => n18242, ZN => n17815);
   U15468 : AOI21_X1 port map( A1 => n17815, A2 => n25902, B => n10792, ZN => 
                           n12420);
   U15469 : INV_X1 port map( I => n17815, ZN => n11186);
   U15471 : AOI22_X1 port map( A1 => n10303, A2 => n22547, B1 => n22551, B2 => 
                           n27402, ZN => n27416);
   U15472 : NAND2_X1 port map( A1 => n25800, A2 => n25799, ZN => n25802);
   U15475 : OR2_X2 port map( A1 => n28557, A2 => n7806, Z => n32855);
   U15477 : OR2_X2 port map( A1 => n28557, A2 => n7806, Z => n32856);
   U15480 : NAND2_X1 port map( A1 => n22784, A2 => n3898, ZN => n17900);
   U15482 : AND2_X1 port map( A1 => n3515, A2 => n3340, Z => n6780);
   U15483 : INV_X2 port map( I => n7555, ZN => n788);
   U15489 : OAI21_X1 port map( A1 => n8178, A2 => n1239, B => n29056, ZN => 
                           n29863);
   U15495 : NAND3_X1 port map( A1 => n30280, A2 => n29056, A3 => n7809, ZN => 
                           n7727);
   U15496 : CLKBUF_X8 port map( I => n8238, Z => n32917);
   U15497 : OR2_X1 port map( A1 => n7993, A2 => n2022, Z => n23858);
   U15499 : INV_X2 port map( I => n7889, ZN => n13457);
   U15500 : NOR2_X1 port map( A1 => n34109, A2 => n5466, ZN => n25237);
   U15502 : NAND2_X1 port map( A1 => n6074, A2 => n21466, ZN => n21283);
   U15503 : CLKBUF_X2 port map( I => n6074, Z => n26728);
   U15504 : OAI21_X1 port map( A1 => n27104, A2 => n24060, B => n13601, ZN => 
                           n3039);
   U15506 : INV_X1 port map( I => n16422, ZN => n16112);
   U15513 : INV_X1 port map( I => n16529, ZN => n1113);
   U15516 : OAI21_X1 port map( A1 => n22567, A2 => n28692, B => n22683, ZN => 
                           n22568);
   U15519 : NOR2_X1 port map( A1 => n9939, A2 => n23936, ZN => n15098);
   U15521 : INV_X2 port map( I => n9939, ZN => n13242);
   U15529 : AOI21_X1 port map( A1 => n17166, A2 => n33205, B => n16287, ZN => 
                           n4505);
   U15535 : NOR2_X1 port map( A1 => n16287, A2 => n31417, ZN => n18864);
   U15540 : NAND2_X1 port map( A1 => n14194, A2 => n11203, ZN => n18842);
   U15541 : INV_X1 port map( I => n14194, ZN => n19216);
   U15543 : NAND2_X1 port map( A1 => n7557, A2 => n14194, ZN => n16336);
   U15552 : OR2_X1 port map( A1 => n13413, A2 => n16384, Z => n23590);
   U15565 : INV_X1 port map( I => n25258, ZN => n25250);
   U15566 : AND2_X1 port map( A1 => n13532, A2 => n32875, Z => n9861);
   U15568 : OAI22_X1 port map( A1 => n28952, A2 => n16793, B1 => n25514, B2 => 
                           n2480, ZN => n33401);
   U15570 : INV_X1 port map( I => n24643, ZN => n242);
   U15577 : OAI21_X1 port map( A1 => n13078, A2 => n9065, B => n22595, ZN => 
                           n22596);
   U15584 : NAND3_X1 port map( A1 => n30708, A2 => n25102, A3 => n3824, ZN => 
                           n32984);
   U15588 : NOR2_X1 port map( A1 => n27233, A2 => n25951, ZN => n27232);
   U15589 : NAND2_X1 port map( A1 => n24232, A2 => n972, ZN => n27381);
   U15598 : AOI22_X1 port map( A1 => n6772, A2 => n29120, B1 => n24232, B2 => 
                           n14399, ZN => n3633);
   U15599 : AOI22_X1 port map( A1 => n2558, A2 => n24232, B1 => n6476, B2 => 
                           n14399, ZN => n29836);
   U15605 : NAND2_X1 port map( A1 => n25586, A2 => n34169, ZN => n25530);
   U15606 : NOR2_X1 port map( A1 => n25590, A2 => n25586, ZN => n13560);
   U15607 : INV_X1 port map( I => n12042, ZN => n967);
   U15617 : NAND2_X1 port map( A1 => n1786, A2 => n12476, ZN => n25113);
   U15629 : CLKBUF_X1 port map( I => n16380, Z => n31207);
   U15630 : NAND2_X1 port map( A1 => n25066, A2 => n31207, ZN => n16836);
   U15632 : INV_X1 port map( I => n22832, ZN => n806);
   U15635 : OR2_X2 port map( A1 => n22832, A2 => n4110, Z => n4731);
   U15637 : CLKBUF_X4 port map( I => n9301, Z => n9195);
   U15638 : INV_X1 port map( I => n9870, ZN => n22580);
   U15642 : INV_X1 port map( I => n25128, ZN => n25130);
   U15653 : NAND2_X1 port map( A1 => n25128, A2 => n1075, ZN => n31617);
   U15654 : CLKBUF_X4 port map( I => n15012, Z => n14454);
   U15655 : NAND2_X1 port map( A1 => n4655, A2 => n14147, ZN => n24092);
   U15657 : INV_X2 port map( I => n14147, ZN => n28694);
   U15659 : OR3_X1 port map( A1 => n7081, A2 => n25337, A3 => n11132, Z => 
                           n25342);
   U15660 : INV_X1 port map( I => n30991, ZN => n23955);
   U15661 : OAI21_X1 port map( A1 => n15974, A2 => n29056, B => n24263, ZN => 
                           n13616);
   U15666 : NOR2_X2 port map( A1 => n27854, A2 => n26949, ZN => n13615);
   U15667 : NAND2_X1 port map( A1 => n18143, A2 => n22499, ZN => n32858);
   U15669 : NAND2_X2 port map( A1 => n22500, A2 => n22691, ZN => n18143);
   U15670 : OR2_X1 port map( A1 => n25621, A2 => n25620, Z => n16001);
   U15673 : NAND2_X1 port map( A1 => n23026, A2 => n26169, ZN => n11495);
   U15677 : CLKBUF_X4 port map( I => n23706, Z => n14080);
   U15679 : INV_X1 port map( I => n25624, ZN => n1219);
   U15682 : OAI21_X1 port map( A1 => n24327, A2 => n24328, B => n24326, ZN => 
                           n28030);
   U15684 : INV_X1 port map( I => n12746, ZN => n33926);
   U15688 : INV_X2 port map( I => n11912, ZN => n12746);
   U15689 : BUF_X2 port map( I => n23834, Z => n16424);
   U15690 : INV_X1 port map( I => n16424, ZN => n33166);
   U15691 : NAND3_X1 port map( A1 => n2640, A2 => n27038, A3 => n31615, ZN => 
                           n668);
   U15699 : NOR3_X1 port map( A1 => n793, A2 => n26120, A3 => n27038, ZN => 
                           n17747);
   U15700 : NOR2_X1 port map( A1 => n26120, A2 => n6713, ZN => n8142);
   U15702 : NAND2_X1 port map( A1 => n7753, A2 => n15414, ZN => n21613);
   U15710 : OAI21_X1 port map( A1 => n1316, A2 => n21752, B => n15414, ZN => 
                           n13662);
   U15714 : CLKBUF_X4 port map( I => n25654, Z => n7083);
   U15715 : NAND2_X1 port map( A1 => n8924, A2 => n31835, ZN => n21151);
   U15716 : INV_X2 port map( I => n21395, ZN => n12325);
   U15718 : INV_X4 port map( I => n23767, ZN => n23770);
   U15719 : NOR2_X1 port map( A1 => n9399, A2 => n22483, ZN => n33021);
   U15720 : NAND3_X1 port map( A1 => n9399, A2 => n22483, A3 => n8287, ZN => 
                           n28463);
   U15723 : AOI21_X1 port map( A1 => n12586, A2 => n22982, B => n28234, ZN => 
                           n8037);
   U15728 : NAND2_X1 port map( A1 => n25760, A2 => n4407, ZN => n30221);
   U15733 : OAI21_X1 port map( A1 => n11898, A2 => n33278, B => n24611, ZN => 
                           n8648);
   U15736 : OAI21_X1 port map( A1 => n1300, A2 => n22497, B => n31933, ZN => 
                           n22020);
   U15740 : NAND2_X1 port map( A1 => n22628, A2 => n31933, ZN => n33938);
   U15741 : AND3_X2 port map( A1 => n32998, A2 => n3004, A3 => n23942, Z => 
                           n10019);
   U15742 : CLKBUF_X2 port map( I => n2635, Z => n33596);
   U15744 : NOR2_X1 port map( A1 => n13995, A2 => n2635, ZN => n30488);
   U15750 : NAND2_X1 port map( A1 => n20429, A2 => n2928, ZN => n31111);
   U15753 : NAND2_X1 port map( A1 => n28414, A2 => n20429, ZN => n17808);
   U15754 : INV_X1 port map( I => n20429, ZN => n20498);
   U15761 : NOR2_X1 port map( A1 => n20429, A2 => n2928, ZN => n20259);
   U15764 : AND2_X2 port map( A1 => n19901, A2 => n27655, Z => n31593);
   U15768 : NOR2_X1 port map( A1 => n6605, A2 => n30976, ZN => n11925);
   U15787 : NAND2_X1 port map( A1 => n25326, A2 => n16528, ZN => n33921);
   U15792 : INV_X1 port map( I => n25796, ZN => n25781);
   U15798 : OAI21_X1 port map( A1 => n12395, A2 => n25797, B => n25796, ZN => 
                           n25800);
   U15801 : NOR2_X1 port map( A1 => n19451, A2 => n16317, ZN => n3591);
   U15808 : NAND2_X1 port map( A1 => n7335, A2 => n32909, ZN => n30708);
   U15810 : NAND2_X1 port map( A1 => n1127, A2 => n2547, ZN => n22669);
   U15812 : NOR2_X1 port map( A1 => n2141, A2 => n24242, ZN => n3947);
   U15813 : NAND2_X1 port map( A1 => n5141, A2 => n21426, ZN => n28342);
   U15819 : NAND2_X1 port map( A1 => n21426, A2 => n17624, ZN => n30091);
   U15821 : OAI22_X1 port map( A1 => n30091, A2 => n28211, B1 => n21426, B2 => 
                           n28594, ZN => n21195);
   U15823 : OAI21_X1 port map( A1 => n17624, A2 => n21426, B => n28342, ZN => 
                           n21196);
   U15824 : INV_X1 port map( I => n15806, ZN => n23069);
   U15825 : NAND2_X1 port map( A1 => n23070, A2 => n15806, ZN => n4806);
   U15830 : NAND2_X1 port map( A1 => n22905, A2 => n15806, ZN => n22907);
   U15831 : INV_X1 port map( I => n15296, ZN => n18079);
   U15835 : AOI22_X1 port map( A1 => n11058, A2 => n11059, B1 => n4067, B2 => 
                           n7181, ZN => n11057);
   U15837 : OAI21_X1 port map( A1 => n903, A2 => n4100, B => n3810, ZN => n9158
                           );
   U15838 : NAND2_X2 port map( A1 => n5741, A2 => n24193, ZN => n5690);
   U15844 : NAND3_X1 port map( A1 => n18220, A2 => n25697, A3 => n25695, ZN => 
                           n33119);
   U15856 : AND3_X1 port map( A1 => n25082, A2 => n25107, A3 => n787, Z => 
                           n24857);
   U15858 : NAND2_X1 port map( A1 => n33616, A2 => n27168, ZN => n29753);
   U15860 : AOI22_X1 port map( A1 => n8049, A2 => n719, B1 => n26120, B2 => 
                           n7891, ZN => n11388);
   U15863 : OAI22_X1 port map( A1 => n26120, A2 => n737, B1 => n793, B2 => 
                           n27168, ZN => n8049);
   U15866 : NAND2_X1 port map( A1 => n34009, A2 => n4069, ZN => n17880);
   U15873 : AOI22_X1 port map( A1 => n25013, A2 => n25014, B1 => n25015, B2 => 
                           n17240, ZN => n6283);
   U15879 : INV_X2 port map( I => n11401, ZN => n21642);
   U15882 : CLKBUF_X1 port map( I => n19938, Z => n28644);
   U15886 : OR2_X1 port map( A1 => n11548, A2 => n18075, Z => n25260);
   U15887 : NAND3_X1 port map( A1 => n16393, A2 => n18815, A3 => n18515, ZN => 
                           n4645);
   U15889 : NOR2_X1 port map( A1 => n15296, A2 => n9793, ZN => n3248);
   U15893 : INV_X1 port map( I => n5708, ZN => n33567);
   U15895 : NAND3_X2 port map( A1 => n1243, A2 => n24272, A3 => n8412, ZN => 
                           n24495);
   U15896 : NAND2_X2 port map( A1 => n6400, A2 => n30123, ZN => n32861);
   U15913 : XNOR2_X1 port map( A1 => n24695, A2 => n24740, ZN => n29545);
   U15915 : NAND2_X1 port map( A1 => n6400, A2 => n30123, ZN => n17052);
   U15922 : OAI21_X1 port map( A1 => n25755, A2 => n717, B => n11899, ZN => 
                           n30877);
   U15927 : NAND2_X1 port map( A1 => n13472, A2 => n2654, ZN => n24279);
   U15931 : INV_X2 port map( I => n665, ZN => n34008);
   U15932 : AOI22_X1 port map( A1 => n20269, A2 => n5781, B1 => n17693, B2 => 
                           n20494, ZN => n20650);
   U15935 : NAND2_X1 port map( A1 => n15250, A2 => n15249, ZN => n33958);
   U15936 : INV_X2 port map( I => n10281, ZN => n32862);
   U15939 : NOR3_X1 port map( A1 => n10606, A2 => n10605, A3 => n30018, ZN => 
                           n27060);
   U15940 : INV_X1 port map( I => n4886, ZN => n5755);
   U15948 : BUF_X2 port map( I => n28119, Z => n32878);
   U15953 : INV_X1 port map( I => n23067, ZN => n18159);
   U15961 : NOR2_X1 port map( A1 => n23067, A2 => n23070, ZN => n30967);
   U15962 : OAI22_X1 port map( A1 => n12043, A2 => n31914, B1 => n29626, B2 => 
                           n22639, ZN => n33610);
   U15963 : INV_X1 port map( I => n24829, ZN => n11842);
   U15968 : NOR2_X1 port map( A1 => n24250, A2 => n24248, ZN => n31664);
   U15972 : NAND2_X1 port map( A1 => n6512, A2 => n24430, ZN => n32863);
   U15973 : AOI22_X1 port map( A1 => n1219, A2 => n31921, B1 => n16397, B2 => 
                           n32896, ZN => n33773);
   U15981 : NOR2_X1 port map( A1 => n3487, A2 => n16959, ZN => n27020);
   U15985 : INV_X2 port map( I => n16959, ZN => n28899);
   U15987 : INV_X1 port map( I => n25014, ZN => n24976);
   U15990 : AOI21_X1 port map( A1 => n901, A2 => n8314, B => n1728, ZN => 
                           n26803);
   U15998 : NOR2_X1 port map( A1 => n8766, A2 => n1209, ZN => n33102);
   U16001 : INV_X1 port map( I => n25302, ZN => n32864);
   U16004 : OAI21_X1 port map( A1 => n11255, A2 => n24325, B => n30186, ZN => 
                           n9826);
   U16005 : NAND2_X1 port map( A1 => n3729, A2 => n1083, ZN => n3728);
   U16008 : CLKBUF_X1 port map( I => n19284, Z => n30501);
   U16009 : CLKBUF_X12 port map( I => n20137, Z => n27911);
   U16010 : AOI22_X1 port map( A1 => n23957, A2 => n13720, B1 => n14232, B2 => 
                           n23825, ZN => n29811);
   U16019 : NAND2_X1 port map( A1 => n14133, A2 => n13720, ZN => n13981);
   U16022 : AOI22_X1 port map( A1 => n29541, A2 => n998, B1 => n905, B2 => 
                           n22467, ZN => n29790);
   U16023 : NAND3_X1 port map( A1 => n32868, A2 => n27622, A3 => n5915, ZN => 
                           n12071);
   U16026 : OR2_X1 port map( A1 => n17936, A2 => n11920, Z => n18094);
   U16027 : NOR2_X1 port map( A1 => n18098, A2 => n11920, ZN => n16866);
   U16030 : INV_X2 port map( I => n7492, ZN => n11000);
   U16032 : INV_X2 port map( I => n17273, ZN => n11571);
   U16034 : CLKBUF_X1 port map( I => n28196, Z => n33851);
   U16036 : INV_X2 port map( I => n11559, ZN => n11904);
   U16037 : NOR3_X1 port map( A1 => n23806, A2 => n11904, A3 => n1247, ZN => 
                           n29705);
   U16040 : NAND2_X1 port map( A1 => n1247, A2 => n11904, ZN => n12248);
   U16050 : OAI21_X1 port map( A1 => n1247, A2 => n11904, B => n23806, ZN => 
                           n15683);
   U16051 : AOI21_X1 port map( A1 => n1100, A2 => n11904, B => n28273, ZN => 
                           n18167);
   U16053 : NAND2_X1 port map( A1 => n1850, A2 => n12476, ZN => n12295);
   U16057 : INV_X2 port map( I => n11987, ZN => n25199);
   U16061 : CLKBUF_X4 port map( I => n25014, Z => n14959);
   U16072 : INV_X1 port map( I => n386, ZN => n17396);
   U16074 : NOR2_X1 port map( A1 => n9778, A2 => n5035, ZN => n28877);
   U16076 : INV_X1 port map( I => n3093, ZN => n32932);
   U16084 : NAND2_X1 port map( A1 => n3093, A2 => n5455, ZN => n19313);
   U16093 : NAND2_X1 port map( A1 => n10999, A2 => n3093, ZN => n33261);
   U16094 : CLKBUF_X4 port map( I => n5612, Z => n25991);
   U16095 : NAND2_X1 port map( A1 => n25308, A2 => n32096, ZN => n33169);
   U16096 : OAI21_X1 port map( A1 => n25391, A2 => n17717, B => n25962, ZN => 
                           n9548);
   U16098 : NAND2_X1 port map( A1 => n17717, A2 => n25962, ZN => n18099);
   U16099 : NOR2_X1 port map( A1 => n25487, A2 => n25462, ZN => n17199);
   U16100 : NOR2_X1 port map( A1 => n32750, A2 => n3748, ZN => n33568);
   U16101 : INV_X1 port map( I => n13648, ZN => n23068);
   U16105 : INV_X2 port map( I => n4580, ZN => n23070);
   U16107 : NAND2_X1 port map( A1 => n11754, A2 => n30505, ZN => n14530);
   U16108 : CLKBUF_X4 port map( I => n8374, Z => n2879);
   U16109 : NOR2_X1 port map( A1 => n25296, A2 => n16650, ZN => n28186);
   U16110 : AND2_X2 port map( A1 => n2570, A2 => n30403, Z => n32865);
   U16114 : NOR2_X1 port map( A1 => n987, A2 => n22957, ZN => n22901);
   U16115 : BUF_X2 port map( I => n17947, Z => n29695);
   U16116 : AND2_X2 port map( A1 => n25409, A2 => n15496, Z => n25329);
   U16117 : NOR2_X1 port map( A1 => n25995, A2 => n14737, ZN => n7272);
   U16120 : NAND2_X1 port map( A1 => n22886, A2 => n23093, ZN => n13618);
   U16123 : NAND3_X1 port map( A1 => n10376, A2 => n789, A3 => n13684, ZN => 
                           n25727);
   U16130 : OAI21_X1 port map( A1 => n25731, A2 => n16494, B => n10376, ZN => 
                           n1896);
   U16140 : CLKBUF_X4 port map( I => n25145, Z => n29976);
   U16141 : NAND2_X1 port map( A1 => n14972, A2 => n25973, ZN => n28703);
   U16144 : NAND2_X1 port map( A1 => n2456, A2 => n25234, ZN => n8841);
   U16145 : NAND2_X1 port map( A1 => n8784, A2 => n21579, ZN => n3472);
   U16146 : OAI22_X1 port map( A1 => n19010, A2 => n17445, B1 => n944, B2 => 
                           n17444, ZN => n27460);
   U16164 : OR2_X2 port map( A1 => n944, A2 => n18913, Z => n5139);
   U16166 : OR2_X1 port map( A1 => n8412, A2 => n29306, Z => n15537);
   U16167 : AND3_X2 port map( A1 => n30930, A2 => n30555, A3 => n28217, Z => 
                           n32867);
   U16173 : NAND3_X1 port map( A1 => n753, A2 => n17717, A3 => n28136, ZN => 
                           n30555);
   U16175 : NAND3_X1 port map( A1 => n29388, A2 => n33680, A3 => n33540, ZN => 
                           n1475);
   U16185 : NAND2_X1 port map( A1 => n25058, A2 => n25044, ZN => n25059);
   U16187 : INV_X1 port map( I => n22856, ZN => n986);
   U16188 : NAND2_X1 port map( A1 => n13859, A2 => n6275, ZN => n3940);
   U16189 : CLKBUF_X2 port map( I => n9133, Z => n33147);
   U16192 : NOR2_X1 port map( A1 => n19058, A2 => n945, ZN => n5709);
   U16193 : AOI21_X1 port map( A1 => n9982, A2 => n25615, B => n10174, ZN => 
                           n9981);
   U16199 : OAI21_X1 port map( A1 => n21642, A2 => n21651, B => n31511, ZN => 
                           n21555);
   U16202 : INV_X1 port map( I => n24289, ZN => n15977);
   U16204 : NOR2_X1 port map( A1 => n21358, A2 => n5018, ZN => n28882);
   U16205 : INV_X2 port map( I => n21358, ZN => n1140);
   U16216 : AND3_X1 port map( A1 => n16254, A2 => n23109, A3 => n23111, Z => 
                           n78);
   U16227 : NOR2_X2 port map( A1 => n31795, A2 => n28853, ZN => n13006);
   U16229 : NAND2_X1 port map( A1 => n23052, A2 => n23051, ZN => n4006);
   U16237 : AOI21_X1 port map( A1 => n1108, A2 => n23052, B => n25994, ZN => 
                           n4487);
   U16239 : NAND2_X1 port map( A1 => n23052, A2 => n23053, ZN => n1745);
   U16244 : OAI21_X1 port map( A1 => n16054, A2 => n23052, B => n31129, ZN => 
                           n9949);
   U16245 : INV_X2 port map( I => n15038, ZN => n9736);
   U16256 : INV_X2 port map( I => n16589, ZN => n25187);
   U16257 : OAI21_X1 port map( A1 => n25235, A2 => n8219, B => n16589, ZN => 
                           n3729);
   U16258 : INV_X2 port map( I => n25563, ZN => n765);
   U16261 : INV_X1 port map( I => n25563, ZN => n33394);
   U16271 : NAND2_X1 port map( A1 => n25592, A2 => n25624, ZN => n8854);
   U16277 : NOR2_X2 port map( A1 => n25429, A2 => n11640, ZN => n408);
   U16278 : NAND2_X1 port map( A1 => n6662, A2 => n15600, ZN => n7034);
   U16279 : NAND3_X1 port map( A1 => n33078, A2 => n19180, A3 => n19178, ZN => 
                           n13011);
   U16281 : AOI22_X1 port map( A1 => n19177, A2 => n19180, B1 => n18114, B2 => 
                           n784, ZN => n2126);
   U16283 : CLKBUF_X4 port map( I => n25903, Z => n28455);
   U16288 : OAI21_X1 port map( A1 => n25180, A2 => n25179, B => n33428, ZN => 
                           n25181);
   U16289 : OAI22_X1 port map( A1 => n21159, A2 => n26133, B1 => n21158, B2 => 
                           n1020, ZN => n28038);
   U16294 : OAI21_X1 port map( A1 => n33507, A2 => n715, B => n15462, ZN => 
                           n7303);
   U16302 : NOR3_X1 port map( A1 => n5926, A2 => n25571, A3 => n27113, ZN => 
                           n30200);
   U16303 : NAND3_X1 port map( A1 => n13660, A2 => n11937, A3 => n24198, ZN => 
                           n17494);
   U16305 : CLKBUF_X12 port map( I => n22602, Z => n16665);
   U16310 : NAND2_X1 port map( A1 => n33107, A2 => n20419, ZN => n10322);
   U16315 : NAND2_X1 port map( A1 => n24056, A2 => n24002, ZN => n24162);
   U16318 : INV_X2 port map( I => n24056, ZN => n29566);
   U16320 : NAND2_X2 port map( A1 => n21909, A2 => n32021, ZN => n22730);
   U16323 : OR2_X2 port map( A1 => n21688, A2 => n12561, Z => n27073);
   U16329 : NAND2_X1 port map( A1 => n28839, A2 => n13063, ZN => n5374);
   U16333 : NAND2_X1 port map( A1 => n12904, A2 => n18146, ZN => n24144);
   U16334 : XNOR2_X1 port map( A1 => n5023, A2 => n5022, ZN => n32873);
   U16338 : OAI21_X1 port map( A1 => n7334, A2 => n5713, B => n25107, ZN => 
                           n32909);
   U16340 : NAND2_X1 port map( A1 => n8926, A2 => n25174, ZN => n8925);
   U16341 : NAND3_X2 port map( A1 => n1213, A2 => n9162, A3 => n6034, ZN => 
                           n25138);
   U16348 : CLKBUF_X4 port map( I => n10943, Z => n34005);
   U16356 : INV_X1 port map( I => n13349, ZN => n33598);
   U16360 : OAI21_X1 port map( A1 => n21162, A2 => n21161, B => n21139, ZN => 
                           n21140);
   U16363 : NAND2_X1 port map( A1 => n21466, A2 => n31085, ZN => n9666);
   U16365 : XNOR2_X1 port map( A1 => n30749, A2 => n10332, ZN => n20967);
   U16366 : INV_X1 port map( I => n10332, ZN => n1345);
   U16370 : INV_X2 port map( I => n1294, ZN => n13703);
   U16371 : AOI21_X1 port map( A1 => n24718, A2 => n12266, B => n11735, ZN => 
                           n17304);
   U16378 : NAND2_X1 port map( A1 => n20427, A2 => n12421, ZN => n14620);
   U16379 : NAND2_X1 port map( A1 => n28376, A2 => n12421, ZN => n19827);
   U16382 : AOI21_X1 port map( A1 => n12482, A2 => n12247, B => n15274, ZN => 
                           n11759);
   U16390 : XOR2_X1 port map( A1 => n16989, A2 => n27896, Z => n32875);
   U16394 : INV_X1 port map( I => n221, ZN => n32876);
   U16399 : NOR2_X1 port map( A1 => n24339, A2 => n24056, ZN => n29018);
   U16401 : INV_X2 port map( I => n25176, ZN => n16273);
   U16402 : NOR2_X1 port map( A1 => n33353, A2 => n25257, ZN => n32954);
   U16404 : XNOR2_X1 port map( A1 => n24826, A2 => n24532, ZN => n24673);
   U16416 : AND2_X2 port map( A1 => n29681, A2 => n30802, Z => n32879);
   U16417 : NAND2_X2 port map( A1 => n33443, A2 => n33442, ZN => n30802);
   U16418 : NAND2_X1 port map( A1 => n33126, A2 => n11382, ZN => n32880);
   U16425 : XOR2_X1 port map( A1 => n13504, A2 => n12749, Z => n32883);
   U16426 : INV_X1 port map( I => n5118, ZN => n19011);
   U16429 : AOI21_X1 port map( A1 => n22899, A2 => n22592, B => n22705, ZN => 
                           n10896);
   U16430 : INV_X1 port map( I => n12238, ZN => n10126);
   U16431 : AOI21_X1 port map( A1 => n32869, A2 => n25444, B => n31263, ZN => 
                           n15498);
   U16435 : NAND2_X2 port map( A1 => n33243, A2 => n33644, ZN => n32885);
   U16436 : XNOR2_X1 port map( A1 => n32885, A2 => n10075, ZN => n30671);
   U16438 : NAND2_X1 port map( A1 => n33243, A2 => n33644, ZN => n22059);
   U16441 : INV_X2 port map( I => n25175, ZN => n14531);
   U16450 : INV_X1 port map( I => n19899, ZN => n20033);
   U16463 : INV_X1 port map( I => n20577, ZN => n32989);
   U16464 : NOR2_X1 port map( A1 => n20312, A2 => n20577, ZN => n17647);
   U16470 : NAND2_X1 port map( A1 => n4396, A2 => n33281, ZN => n33280);
   U16474 : OAI21_X1 port map( A1 => n22558, A2 => n4396, B => n9630, ZN => 
                           n32955);
   U16476 : INV_X1 port map( I => n4396, ZN => n22671);
   U16484 : OAI21_X1 port map( A1 => n1140, A2 => n30267, B => n11967, ZN => 
                           n21273);
   U16489 : NOR2_X1 port map( A1 => n12037, A2 => n11967, ZN => n12492);
   U16490 : INV_X2 port map( I => n11967, ZN => n1331);
   U16491 : INV_X1 port map( I => n7699, ZN => n10142);
   U16493 : NAND2_X1 port map( A1 => n20494, A2 => n17497, ZN => n5779);
   U16501 : INV_X2 port map( I => n17497, ZN => n20268);
   U16502 : NOR3_X1 port map( A1 => n27752, A2 => n30293, A3 => n28680, ZN => 
                           n13431);
   U16506 : OAI22_X1 port map( A1 => n6074, A2 => n14012, B1 => n16127, B2 => 
                           n32073, ZN => n21600);
   U16510 : OAI21_X1 port map( A1 => n30318, A2 => n3489, B => n747, ZN => 
                           n7341);
   U16511 : AND2_X1 port map( A1 => n26551, A2 => n3816, Z => n19944);
   U16514 : INV_X1 port map( I => n22138, ZN => n16210);
   U16517 : INV_X1 port map( I => n23813, ZN => n23852);
   U16521 : CLKBUF_X12 port map( I => n11845, Z => n26545);
   U16524 : NAND2_X1 port map( A1 => n230, A2 => n21512, ZN => n5787);
   U16527 : INV_X1 port map( I => n10219, ZN => n33200);
   U16528 : NAND2_X1 port map( A1 => n31566, A2 => n3007, ZN => n23058);
   U16530 : NAND3_X1 port map( A1 => n21392, A2 => n17522, A3 => n21163, ZN => 
                           n4784);
   U16535 : AOI21_X1 port map( A1 => n21163, A2 => n21392, B => n17522, ZN => 
                           n2604);
   U16538 : XNOR2_X1 port map( A1 => Plaintext(31), A2 => Key(31), ZN => n18139
                           );
   U16539 : OAI21_X1 port map( A1 => n20533, A2 => n20463, B => n28028, ZN => 
                           n4077);
   U16540 : XOR2_X1 port map( A1 => n17498, A2 => n6397, Z => n32886);
   U16542 : AOI21_X2 port map( A1 => n5810, A2 => n8186, B => n32992, ZN => 
                           n32887);
   U16544 : INV_X1 port map( I => n24276, ZN => n34137);
   U16551 : AOI21_X1 port map( A1 => n3984, A2 => n24276, B => n7068, ZN => 
                           n24169);
   U16552 : AND2_X1 port map( A1 => n31939, A2 => n9486, Z => n7065);
   U16557 : AOI21_X1 port map( A1 => n6662, A2 => n26115, B => n5191, ZN => 
                           n13906);
   U16561 : NAND2_X1 port map( A1 => n24002, A2 => n2826, ZN => n7171);
   U16565 : NOR2_X1 port map( A1 => n25806, A2 => n25820, ZN => n25817);
   U16566 : INV_X2 port map( I => n9126, ZN => n16113);
   U16572 : NOR2_X1 port map( A1 => n10967, A2 => n23862, ZN => n30736);
   U16575 : INV_X1 port map( I => n23862, ZN => n13031);
   U16576 : INV_X2 port map( I => n9252, ZN => n580);
   U16577 : AND2_X1 port map( A1 => n14600, A2 => n15299, Z => n10405);
   U16579 : INV_X2 port map( I => n32096, ZN => n25391);
   U16581 : AOI21_X1 port map( A1 => n794, A2 => n4604, B => n11049, ZN => 
                           n13552);
   U16593 : NAND2_X1 port map( A1 => n33857, A2 => n17888, ZN => n27707);
   U16594 : NAND3_X1 port map( A1 => n25043, A2 => n25062, A3 => n25042, ZN => 
                           n28220);
   U16595 : NAND3_X1 port map( A1 => n25731, A2 => n25724, A3 => n13640, ZN => 
                           n25725);
   U16596 : INV_X2 port map( I => n23888, ZN => n23887);
   U16602 : CLKBUF_X4 port map( I => n23888, Z => n29240);
   U16612 : NOR2_X1 port map( A1 => n9405, A2 => n21452, ZN => n9324);
   U16618 : NOR2_X1 port map( A1 => n7291, A2 => n7852, ZN => n20397);
   U16619 : XOR2_X1 port map( A1 => n27976, A2 => n30016, Z => n32888);
   U16620 : AND3_X2 port map( A1 => n7279, A2 => n14161, A3 => n20627, Z => 
                           n31291);
   U16624 : AOI21_X1 port map( A1 => n28736, A2 => n14810, B => n788, ZN => 
                           n8723);
   U16629 : INV_X2 port map( I => n16981, ZN => n14232);
   U16631 : NAND2_X1 port map( A1 => n16981, A2 => n11096, ZN => n15616);
   U16632 : NOR2_X1 port map( A1 => n30584, A2 => n3909, ZN => n8083);
   U16633 : INV_X1 port map( I => n32452, ZN => n7044);
   U16637 : OAI21_X1 port map( A1 => n27685, A2 => n30832, B => n9472, ZN => 
                           n5495);
   U16650 : OAI21_X1 port map( A1 => n5863, A2 => n7811, B => n21872, ZN => 
                           n12390);
   U16655 : NAND2_X1 port map( A1 => n5863, A2 => n9472, ZN => n12354);
   U16660 : NOR2_X1 port map( A1 => n17720, A2 => n32858, ZN => n12107);
   U16661 : INV_X2 port map( I => n17720, ZN => n15601);
   U16662 : CLKBUF_X4 port map( I => n16798, Z => n8766);
   U16663 : INV_X2 port map( I => n16798, ZN => n749);
   U16664 : INV_X1 port map( I => n10858, ZN => n25193);
   U16665 : NAND2_X1 port map( A1 => n19320, A2 => n19274, ZN => n33389);
   U16666 : NAND2_X1 port map( A1 => n29317, A2 => n4908, ZN => n8954);
   U16667 : NAND2_X1 port map( A1 => n29317, A2 => n13694, ZN => n23072);
   U16669 : AOI21_X1 port map( A1 => n916, A2 => n196, B => n11755, ZN => n9898
                           );
   U16673 : AOI21_X1 port map( A1 => n5850, A2 => n27954, B => n11755, ZN => 
                           n5849);
   U16676 : INV_X1 port map( I => n17305, ZN => n32907);
   U16677 : NAND2_X1 port map( A1 => n21161, A2 => n17305, ZN => n7050);
   U16678 : INV_X1 port map( I => n3286, ZN => n17644);
   U16679 : INV_X2 port map( I => n12657, ZN => n5371);
   U16687 : NAND2_X1 port map( A1 => n13574, A2 => n29173, ZN => n1561);
   U16692 : CLKBUF_X12 port map( I => n2655, Z => n123);
   U16694 : AOI21_X1 port map( A1 => n13059, A2 => n14811, B => n12548, ZN => 
                           n6188);
   U16695 : BUF_X2 port map( I => n18076, Z => n11097);
   U16700 : INV_X1 port map( I => n18076, ZN => n31669);
   U16705 : INV_X1 port map( I => n18861, ZN => n18863);
   U16706 : XOR2_X1 port map( A1 => n30767, A2 => n7071, Z => n32890);
   U16707 : NAND3_X1 port map( A1 => n14752, A2 => n10755, A3 => n27248, ZN => 
                           n24365);
   U16710 : INV_X2 port map( I => n22979, ZN => n31531);
   U16712 : NAND2_X1 port map( A1 => n22978, A2 => n22979, ZN => n28348);
   U16721 : OR2_X2 port map( A1 => n29908, A2 => n11364, Z => n3005);
   U16722 : NAND2_X1 port map( A1 => n3169, A2 => n17150, ZN => n12848);
   U16727 : OR2_X1 port map( A1 => n28811, A2 => n16776, Z => n23728);
   U16729 : OAI21_X1 port map( A1 => n25987, A2 => n16776, B => n23728, ZN => 
                           n17134);
   U16733 : INV_X1 port map( I => n30045, ZN => n32892);
   U16734 : OR2_X2 port map( A1 => n32891, A2 => n8327, Z => n6109);
   U16735 : OR2_X1 port map( A1 => n31922, A2 => n32891, Z => n9033);
   U16736 : NAND2_X1 port map( A1 => n535, A2 => n23197, ZN => n23804);
   U16740 : AOI21_X2 port map( A1 => n23006, A2 => n3999, B => n23004, ZN => 
                           n32893);
   U16741 : AOI21_X2 port map( A1 => n16883, A2 => n20220, B => n30530, ZN => 
                           n32894);
   U16745 : XOR2_X1 port map( A1 => n22970, A2 => n23375, Z => n32895);
   U16749 : NOR3_X1 port map( A1 => n15139, A2 => n18006, A3 => n18007, ZN => 
                           n18005);
   U16757 : INV_X1 port map( I => n14132, ZN => n9568);
   U16759 : CLKBUF_X12 port map( I => n16309, Z => n26766);
   U16761 : OAI21_X1 port map( A1 => n14627, A2 => n17987, B => n15641, ZN => 
                           n15331);
   U16764 : NOR2_X1 port map( A1 => n4897, A2 => n15227, ZN => n27963);
   U16766 : AOI21_X1 port map( A1 => n9687, A2 => n14490, B => n4897, ZN => 
                           n33390);
   U16767 : INV_X2 port map( I => n10612, ZN => n31345);
   U16772 : INV_X1 port map( I => n837, ZN => n32896);
   U16774 : NAND2_X2 port map( A1 => n6656, A2 => n26614, ZN => n32897);
   U16776 : NAND2_X1 port map( A1 => n6656, A2 => n26614, ZN => n25515);
   U16778 : NAND2_X2 port map( A1 => n24864, A2 => n16397, ZN => n6656);
   U16780 : NOR2_X2 port map( A1 => n8149, A2 => n8150, ZN => n32899);
   U16782 : OAI21_X1 port map( A1 => n33850, A2 => n9393, B => n9392, ZN => 
                           n8323);
   U16785 : INV_X2 port map( I => n1877, ZN => n31522);
   U16786 : BUF_X2 port map( I => n8088, Z => n28737);
   U16787 : NOR2_X1 port map( A1 => n723, A2 => n31325, ZN => n11564);
   U16789 : NAND2_X1 port map( A1 => n27719, A2 => n31325, ZN => n10884);
   U16799 : NAND2_X1 port map( A1 => n723, A2 => n31325, ZN => n3830);
   U16801 : INV_X1 port map( I => n24803, ZN => n33100);
   U16803 : NOR2_X1 port map( A1 => n1269, A2 => n7287, ZN => n2579);
   U16809 : AND2_X2 port map( A1 => n27880, A2 => n1284, Z => n27889);
   U16815 : CLKBUF_X12 port map( I => n7881, Z => n28689);
   U16816 : NOR2_X1 port map( A1 => n32595, A2 => n7881, ZN => n16560);
   U16830 : NAND2_X1 port map( A1 => n14133, A2 => n29472, ZN => n23958);
   U16831 : INV_X1 port map( I => n25790, ZN => n16422);
   U16836 : INV_X2 port map( I => n25790, ZN => n25788);
   U16838 : NAND2_X1 port map( A1 => n24062, A2 => n30651, ZN => n6287);
   U16841 : NOR3_X1 port map( A1 => n796, A2 => n30651, A3 => n24207, ZN => 
                           n10652);
   U16845 : INV_X1 port map( I => n30651, ZN => n970);
   U16849 : NAND2_X1 port map( A1 => n7778, A2 => n9220, ZN => n5673);
   U16850 : NAND2_X1 port map( A1 => n25515, A2 => n6595, ZN => n25510);
   U16852 : NOR2_X1 port map( A1 => n22951, A2 => n13762, ZN => n3202);
   U16854 : NOR2_X1 port map( A1 => n2654, A2 => n5454, ZN => n9581);
   U16861 : CLKBUF_X4 port map( I => n5454, Z => n31461);
   U16863 : OR2_X2 port map( A1 => n22565, A2 => n14676, Z => n22680);
   U16867 : NAND3_X1 port map( A1 => n25804, A2 => n25818, A3 => n11003, ZN => 
                           n18246);
   U16871 : AOI22_X1 port map( A1 => n25807, A2 => n25816, B1 => n25804, B2 => 
                           n25817, ZN => n14009);
   U16873 : NAND2_X1 port map( A1 => n15340, A2 => n28358, ZN => n33507);
   U16875 : NOR2_X1 port map( A1 => n28358, A2 => n15340, ZN => n25207);
   U16876 : NAND2_X1 port map( A1 => n3581, A2 => n30333, ZN => n33227);
   U16880 : INV_X1 port map( I => n30333, ZN => n34039);
   U16892 : NOR2_X1 port map( A1 => n31263, A2 => n17948, ZN => n25432);
   U16894 : NAND2_X1 port map( A1 => n17948, A2 => n25437, ZN => n25445);
   U16902 : INV_X1 port map( I => n17948, ZN => n25425);
   U16910 : OAI21_X2 port map( A1 => n6204, A2 => n28706, B => n24889, ZN => 
                           n32900);
   U16914 : INV_X1 port map( I => n9301, ZN => n33681);
   U16916 : XOR2_X1 port map( A1 => Plaintext(110), A2 => Key(110), Z => n32901
                           );
   U16917 : XOR2_X1 port map( A1 => n10707, A2 => n27766, Z => n32902);
   U16918 : OR2_X1 port map( A1 => n23018, A2 => n9575, Z => n13274);
   U16927 : NAND2_X1 port map( A1 => n21811, A2 => n8140, ZN => n15774);
   U16928 : OAI22_X2 port map( A1 => n3866, A2 => n3867, B1 => n6568, B2 => 
                           n10096, ZN => n32904);
   U16930 : OR2_X2 port map( A1 => n32904, A2 => n21601, Z => n6238);
   U16931 : CLKBUF_X12 port map( I => n31497, Z => n31113);
   U16932 : AOI21_X1 port map( A1 => n2444, A2 => n24216, B => n31497, ZN => 
                           n10047);
   U16934 : NOR2_X1 port map( A1 => n889, A2 => n31497, ZN => n6225);
   U16936 : AND3_X2 port map( A1 => n25975, A2 => n21715, A3 => n5704, Z => 
                           n9591);
   U16937 : NOR2_X1 port map( A1 => n8270, A2 => n843, ZN => n23788);
   U16938 : XOR2_X1 port map( A1 => n17400, A2 => n32050, Z => n32905);
   U16941 : AOI22_X2 port map( A1 => n32010, A2 => n4110, B1 => n31942, B2 => 
                           n22383, ZN => n8418);
   U16942 : XOR2_X1 port map( A1 => n23475, A2 => n23417, Z => n32906);
   U16943 : XOR2_X1 port map( A1 => n22231, A2 => n22303, Z => n30402);
   U16949 : NAND2_X2 port map( A1 => n15847, A2 => n15846, ZN => n22231);
   U16951 : XOR2_X1 port map( A1 => n22240, A2 => n22197, Z => n22167);
   U16953 : NOR2_X2 port map( A1 => n21600, A2 => n21599, ZN => n22240);
   U16954 : INV_X4 port map( I => n7892, ZN => n20607);
   U16959 : XNOR2_X1 port map( A1 => n33952, A2 => n31116, ZN => n8434);
   U16961 : AOI22_X1 port map( A1 => n25367, A2 => n30302, B1 => n3300, B2 => 
                           n25376, ZN => n25380);
   U16964 : XOR2_X1 port map( A1 => n19497, A2 => n17931, Z => n12653);
   U16967 : NAND2_X2 port map( A1 => n7647, A2 => n6494, ZN => n5713);
   U16969 : NAND2_X2 port map( A1 => n31309, A2 => n5228, ZN => n21933);
   U16971 : NAND2_X1 port map( A1 => n21213, A2 => n32907, ZN => n17375);
   U16974 : NOR2_X2 port map( A1 => n21160, A2 => n32902, ZN => n21213);
   U16975 : INV_X2 port map( I => n20472, ZN => n20317);
   U16978 : NAND2_X2 port map( A1 => n19382, A2 => n27196, ZN => n20472);
   U16982 : NOR2_X1 port map( A1 => n1018, A2 => n21358, ZN => n27828);
   U16987 : XOR2_X1 port map( A1 => n29833, A2 => n33311, Z => n1018);
   U16999 : XOR2_X1 port map( A1 => n23367, A2 => n15941, Z => n10758);
   U17001 : NOR2_X2 port map( A1 => n31823, A2 => n16298, ZN => n19759);
   U17004 : INV_X2 port map( I => n32910, ZN => n28602);
   U17006 : INV_X2 port map( I => n560, ZN => n32911);
   U17007 : XOR2_X1 port map( A1 => n32912, A2 => n10064, Z => n8277);
   U17009 : XOR2_X1 port map( A1 => n27667, A2 => n10459, Z => n32912);
   U17011 : NAND3_X2 port map( A1 => n17108, A2 => n32913, A3 => n30151, ZN => 
                           n25665);
   U17014 : NAND2_X2 port map( A1 => n3774, A2 => n755, ZN => n32913);
   U17017 : XOR2_X1 port map( A1 => n32914, A2 => n14527, Z => n15433);
   U17023 : NAND2_X1 port map( A1 => n32086, A2 => n2226, ZN => n2225);
   U17025 : INV_X1 port map( I => n13472, ZN => n969);
   U17028 : NAND2_X2 port map( A1 => n7613, A2 => n29788, ZN => n13472);
   U17029 : XOR2_X1 port map( A1 => n13794, A2 => n13792, Z => n17037);
   U17040 : NAND2_X2 port map( A1 => n17639, A2 => n22814, ZN => n17085);
   U17045 : INV_X2 port map( I => n19908, ZN => n870);
   U17047 : NAND2_X1 port map( A1 => n6549, A2 => n3967, ZN => n19908);
   U17051 : XOR2_X1 port map( A1 => n33348, A2 => n33588, Z => n32916);
   U17061 : INV_X2 port map( I => n32919, ZN => n8469);
   U17063 : XOR2_X1 port map( A1 => n32921, A2 => n2651, Z => n28611);
   U17065 : XOR2_X1 port map( A1 => n2653, A2 => n32922, Z => n32921);
   U17069 : AOI21_X1 port map( A1 => n28715, A2 => n24340, B => n16552, ZN => 
                           n14847);
   U17071 : INV_X1 port map( I => n2653, ZN => n1865);
   U17078 : XOR2_X1 port map( A1 => n31499, A2 => n29927, Z => n2653);
   U17082 : NAND3_X2 port map( A1 => n23772, A2 => n33668, A3 => n15402, ZN => 
                           n7093);
   U17084 : XOR2_X1 port map( A1 => n32923, A2 => n21014, Z => n12557);
   U17085 : XOR2_X1 port map( A1 => n13681, A2 => n12559, Z => n32923);
   U17086 : NOR2_X1 port map( A1 => n16868, A2 => n24254, ZN => n17802);
   U17093 : XOR2_X1 port map( A1 => n31133, A2 => n22250, Z => n27693);
   U17094 : XOR2_X1 port map( A1 => n31081, A2 => n23490, Z => n28847);
   U17095 : INV_X2 port map( I => n32924, ZN => n7513);
   U17096 : XOR2_X1 port map( A1 => n32925, A2 => n10052, Z => n31844);
   U17104 : NOR2_X2 port map( A1 => n32045, A2 => n1291, ZN => n7398);
   U17105 : XOR2_X1 port map( A1 => n5703, A2 => n4173, Z => n4718);
   U17109 : NAND2_X2 port map( A1 => n24496, A2 => n24495, ZN => n24498);
   U17110 : NAND2_X2 port map( A1 => n12753, A2 => n32927, ZN => n12785);
   U17111 : NAND3_X2 port map( A1 => n15494, A2 => n12788, A3 => n7813, ZN => 
                           n32927);
   U17121 : XOR2_X1 port map( A1 => n12637, A2 => n32928, Z => n17117);
   U17124 : XOR2_X1 port map( A1 => n12636, A2 => n13309, Z => n32928);
   U17128 : NOR2_X1 port map( A1 => n1379, A2 => n19132, ZN => n7418);
   U17129 : NAND2_X1 port map( A1 => n4405, A2 => n19249, ZN => n19132);
   U17133 : XOR2_X1 port map( A1 => n10902, A2 => n32930, Z => n33770);
   U17135 : XOR2_X1 port map( A1 => n27098, A2 => n19654, Z => n10902);
   U17138 : XOR2_X1 port map( A1 => n10006, A2 => n22274, Z => n22084);
   U17140 : INV_X2 port map( I => n21925, ZN => n10006);
   U17150 : OAI21_X1 port map( A1 => n28388, A2 => n10835, B => n692, ZN => 
                           n27342);
   U17151 : NAND2_X2 port map( A1 => n33560, A2 => n27676, ZN => n24008);
   U17158 : NAND2_X1 port map( A1 => n32931, A2 => n17087, ZN => n23927);
   U17159 : AOI22_X2 port map( A1 => n11971, A2 => n20154, B1 => n20153, B2 => 
                           n8259, ZN => n4420);
   U17160 : NOR2_X2 port map( A1 => n19914, A2 => n31951, ZN => n11971);
   U17161 : NOR2_X1 port map( A1 => n31915, A2 => n26641, ZN => n29037);
   U17166 : OAI21_X2 port map( A1 => n31962, A2 => n24557, B => n32933, ZN => 
                           n25285);
   U17168 : AOI22_X1 port map( A1 => n20076, A2 => n12408, B1 => n6444, B2 => 
                           n2499, ZN => n3624);
   U17169 : NAND2_X1 port map( A1 => n2654, A2 => n5454, ZN => n8664);
   U17171 : OAI21_X1 port map( A1 => n16474, A2 => n28344, B => n18805, ZN => 
                           n26909);
   U17174 : AOI22_X2 port map( A1 => n32062, A2 => n32934, B1 => n24308, B2 => 
                           n24135, ZN => n11830);
   U17177 : INV_X2 port map( I => n23714, ZN => n32934);
   U17181 : XOR2_X1 port map( A1 => n14781, A2 => n14783, Z => n16603);
   U17182 : AND3_X1 port map( A1 => n28641, A2 => n5595, A3 => n21223, Z => 
                           n33352);
   U17185 : NAND2_X2 port map( A1 => n1700, A2 => n32920, ZN => n15768);
   U17186 : INV_X2 port map( I => n22108, ZN => n7725);
   U17187 : NAND2_X2 port map( A1 => n8078, A2 => n8077, ZN => n22108);
   U17188 : XOR2_X1 port map( A1 => n32937, A2 => n33017, Z => n28615);
   U17189 : XOR2_X1 port map( A1 => n23330, A2 => n23277, Z => n32937);
   U17198 : INV_X2 port map( I => n32938, ZN => n15722);
   U17202 : XNOR2_X1 port map( A1 => n15507, A2 => n23377, ZN => n32938);
   U17205 : INV_X2 port map( I => n20531, ZN => n32940);
   U17206 : INV_X1 port map( I => n28064, ZN => n32941);
   U17208 : OAI21_X2 port map( A1 => n28786, A2 => n1170, B => n33241, ZN => 
                           n28064);
   U17211 : OAI21_X2 port map( A1 => n10621, A2 => n10620, B => n32942, ZN => 
                           n10281);
   U17212 : AND2_X1 port map( A1 => n5274, A2 => n8365, Z => n26195);
   U17215 : NAND2_X2 port map( A1 => n17008, A2 => n17006, ZN => n5274);
   U17217 : NAND2_X2 port map( A1 => n10760, A2 => n10759, ZN => n15941);
   U17218 : NAND2_X2 port map( A1 => n19310, A2 => n10828, ZN => n18667);
   U17221 : AOI21_X2 port map( A1 => n7662, A2 => n6366, B => n32943, ZN => 
                           n7660);
   U17222 : INV_X2 port map( I => n32945, ZN => n3193);
   U17224 : XOR2_X1 port map( A1 => n3298, A2 => n509, Z => n32945);
   U17225 : XOR2_X1 port map( A1 => n15360, A2 => n11193, Z => n16998);
   U17230 : NOR2_X2 port map( A1 => n22556, A2 => n15362, ZN => n15360);
   U17231 : XOR2_X1 port map( A1 => n10516, A2 => n2074, Z => n10514);
   U17235 : NAND2_X1 port map( A1 => n14633, A2 => n33701, ZN => Ciphertext(57)
                           );
   U17242 : NAND2_X2 port map( A1 => n30870, A2 => n5092, ZN => n13415);
   U17248 : XOR2_X1 port map( A1 => n30284, A2 => n22123, Z => n1971);
   U17252 : NAND2_X2 port map( A1 => n12997, A2 => n14907, ZN => n12982);
   U17255 : NAND2_X2 port map( A1 => n29368, A2 => n30409, ZN => n12997);
   U17256 : XOR2_X1 port map( A1 => n15373, A2 => n17051, Z => n33303);
   U17257 : NAND2_X2 port map( A1 => n33987, A2 => n32946, ZN => n25106);
   U17260 : NAND2_X1 port map( A1 => n15331, A2 => n15332, ZN => n32946);
   U17261 : XOR2_X1 port map( A1 => n24674, A2 => n24673, Z => n24679);
   U17265 : NAND2_X2 port map( A1 => n1749, A2 => n29982, ZN => n23052);
   U17266 : XOR2_X1 port map( A1 => n32947, A2 => n22040, Z => n22535);
   U17267 : INV_X2 port map( I => n13623, ZN => n7361);
   U17270 : NAND4_X2 port map( A1 => n3744, A2 => n7075, A3 => n7074, A4 => 
                           n7076, ZN => n13623);
   U17272 : XOR2_X1 port map( A1 => n23324, A2 => n32948, Z => n11225);
   U17274 : XOR2_X1 port map( A1 => n11227, A2 => n29082, Z => n32948);
   U17276 : INV_X2 port map( I => n3250, ZN => n32949);
   U17280 : NAND2_X2 port map( A1 => n28581, A2 => n15302, ZN => n3250);
   U17281 : OAI21_X2 port map( A1 => n28096, A2 => n18151, B => n32950, ZN => 
                           n12856);
   U17283 : XOR2_X1 port map( A1 => n5932, A2 => n6547, Z => n15674);
   U17290 : NAND2_X2 port map( A1 => n5933, A2 => n5935, ZN => n5932);
   U17291 : XOR2_X1 port map( A1 => n12310, A2 => n23388, Z => n23220);
   U17292 : NAND3_X2 port map( A1 => n12180, A2 => n5136, A3 => n9918, ZN => 
                           n12310);
   U17296 : NAND2_X2 port map( A1 => n4571, A2 => n9835, ZN => n29781);
   U17305 : NOR2_X1 port map( A1 => n16041, A2 => n25322, ZN => n6234);
   U17308 : NAND3_X2 port map( A1 => n30930, A2 => n30555, A3 => n28217, ZN => 
                           n25322);
   U17310 : NAND2_X2 port map( A1 => n23101, A2 => n11956, ZN => n22783);
   U17311 : NAND2_X1 port map( A1 => n32954, A2 => n11569, ZN => n107);
   U17319 : OAI22_X2 port map( A1 => n24149, A2 => n32750, B1 => n9946, B2 => 
                           n24063, ZN => n24064);
   U17320 : INV_X4 port map( I => n1775, ZN => n9946);
   U17325 : NAND2_X2 port map( A1 => n27064, A2 => n1776, ZN => n1775);
   U17329 : NAND2_X2 port map( A1 => n32956, A2 => n11505, ZN => n7552);
   U17333 : BUF_X2 port map( I => n33153, Z => n32957);
   U17335 : OR2_X1 port map( A1 => n33942, A2 => n30200, Z => n31489);
   U17336 : XOR2_X1 port map( A1 => n23296, A2 => n17766, Z => n26371);
   U17338 : XOR2_X1 port map( A1 => n19741, A2 => n19625, Z => n19571);
   U17339 : NOR2_X2 port map( A1 => n30670, A2 => n30768, ZN => n19741);
   U17340 : XOR2_X1 port map( A1 => n32958, A2 => n24918, Z => Ciphertext(5));
   U17343 : AOI22_X1 port map( A1 => n8278, A2 => n10099, B1 => n24915, B2 => 
                           n24916, ZN => n32958);
   U17345 : XOR2_X1 port map( A1 => n24356, A2 => n24370, Z => n24390);
   U17346 : INV_X2 port map( I => n28415, ZN => n32960);
   U17349 : XOR2_X1 port map( A1 => n2435, A2 => n32961, Z => n22350);
   U17357 : XOR2_X1 port map( A1 => n21984, A2 => n29418, Z => n32961);
   U17359 : NOR2_X2 port map( A1 => n745, A2 => n17817, ZN => n19195);
   U17363 : NAND2_X2 port map( A1 => n33122, A2 => n12826, ZN => n17817);
   U17377 : NAND3_X2 port map( A1 => n32963, A2 => n32962, A3 => n363, ZN => 
                           n16045);
   U17379 : NAND3_X2 port map( A1 => n5367, A2 => n5366, A3 => n28833, ZN => 
                           n32963);
   U17381 : NAND2_X2 port map( A1 => n5124, A2 => n32965, ZN => n16960);
   U17383 : AOI22_X2 port map( A1 => n18578, A2 => n18855, B1 => n6873, B2 => 
                           n18854, ZN => n32965);
   U17388 : XOR2_X1 port map( A1 => n29209, A2 => n11416, Z => n16384);
   U17401 : XOR2_X1 port map( A1 => n32966, A2 => n15338, Z => n15153);
   U17402 : XOR2_X1 port map( A1 => n15337, A2 => n20818, Z => n32966);
   U17405 : NAND3_X2 port map( A1 => n24079, A2 => n24080, A3 => n24081, ZN => 
                           n24083);
   U17407 : NAND2_X2 port map( A1 => n18754, A2 => n15193, ZN => n19386);
   U17408 : AND2_X1 port map( A1 => n18830, A2 => n6256, Z => n17054);
   U17414 : XOR2_X1 port map( A1 => n31092, A2 => n30126, Z => n27435);
   U17422 : NOR2_X2 port map( A1 => n22894, A2 => n6605, ZN => n33023);
   U17429 : NAND2_X2 port map( A1 => n29608, A2 => n33982, ZN => n6605);
   U17432 : OAI22_X2 port map( A1 => n18901, A2 => n9787, B1 => n30995, B2 => 
                           n1378, ZN => n5872);
   U17435 : NAND2_X2 port map( A1 => n1378, A2 => n29146, ZN => n18901);
   U17436 : NAND2_X1 port map( A1 => n16372, A2 => n12863, ZN => n12875);
   U17442 : XOR2_X1 port map( A1 => n32968, A2 => n17918, Z => n16618);
   U17443 : XOR2_X1 port map( A1 => n13651, A2 => n22048, Z => n32968);
   U17445 : XOR2_X1 port map( A1 => n24793, A2 => n11217, Z => n30393);
   U17446 : AOI21_X2 port map( A1 => n32969, A2 => n11381, B => n32013, ZN => 
                           n22085);
   U17451 : OR2_X1 port map( A1 => n31859, A2 => n31484, Z => n32969);
   U17457 : OAI21_X2 port map( A1 => n8991, A2 => n10138, B => n10137, ZN => 
                           n22978);
   U17458 : XOR2_X1 port map( A1 => n31901, A2 => n17904, Z => n3503);
   U17462 : XOR2_X1 port map( A1 => n22252, A2 => n14796, Z => n8993);
   U17464 : XOR2_X1 port map( A1 => n21769, A2 => n32970, Z => n29287);
   U17471 : XOR2_X1 port map( A1 => n21921, A2 => n22242, Z => n32970);
   U17476 : NAND2_X2 port map( A1 => n33516, A2 => n32971, ZN => n25806);
   U17477 : NAND3_X1 port map( A1 => n13819, A2 => n1211, A3 => n24710, ZN => 
                           n32971);
   U17478 : OAI21_X2 port map( A1 => n32973, A2 => n23778, B => n32972, ZN => 
                           n23354);
   U17480 : NOR2_X2 port map( A1 => n9181, A2 => n17642, ZN => n25812);
   U17483 : AOI22_X2 port map( A1 => n24102, A2 => n24101, B1 => n14375, B2 => 
                           n24103, ZN => n33505);
   U17486 : AOI22_X2 port map( A1 => n11003, A2 => n9181, B1 => n25818, B2 => 
                           n25823, ZN => n25825);
   U17487 : NAND2_X1 port map( A1 => n28256, A2 => n28255, ZN => n33450);
   U17488 : XOR2_X1 port map( A1 => n32974, A2 => n16622, Z => Ciphertext(3));
   U17492 : NAND2_X2 port map( A1 => n14828, A2 => n16782, ZN => n18830);
   U17494 : AND2_X1 port map( A1 => n29139, A2 => n33175, Z => n32986);
   U17495 : XOR2_X1 port map( A1 => n32977, A2 => n24748, Z => Ciphertext(4));
   U17496 : XOR2_X1 port map( A1 => n10210, A2 => n19504, Z => n5862);
   U17499 : NOR2_X1 port map( A1 => n33155, A2 => n25889, ZN => n11735);
   U17500 : NOR2_X2 port map( A1 => n32980, A2 => n32979, ZN => n32978);
   U17502 : OR2_X1 port map( A1 => n8412, A2 => n24271, Z => n8499);
   U17503 : XOR2_X1 port map( A1 => n12494, A2 => n32981, Z => n516);
   U17504 : NAND2_X2 port map( A1 => n8940, A2 => n29835, ZN => n12494);
   U17506 : XOR2_X1 port map( A1 => n23140, A2 => n33073, Z => n23144);
   U17507 : NAND2_X2 port map( A1 => n32983, A2 => n33667, ZN => n22197);
   U17511 : XOR2_X1 port map( A1 => n32984, A2 => n25104, Z => Ciphertext(51));
   U17522 : OAI21_X2 port map( A1 => n1244, A2 => n889, B => n24289, ZN => 
                           n32985);
   U17523 : NAND3_X1 port map( A1 => n8614, A2 => n3860, A3 => n33722, ZN => 
                           n29964);
   U17528 : NOR2_X2 port map( A1 => n15718, A2 => n22873, ZN => n9460);
   U17532 : INV_X4 port map( I => n865, ZN => n33888);
   U17533 : OAI22_X1 port map( A1 => n22952, A2 => n13762, B1 => n6801, B2 => 
                           n22951, ZN => n6674);
   U17536 : NAND2_X2 port map( A1 => n23915, A2 => n13521, ZN => n7991);
   U17544 : BUF_X4 port map( I => n11676, Z => n33659);
   U17546 : NAND2_X2 port map( A1 => n32987, A2 => n11746, ZN => n22729);
   U17548 : AOI21_X2 port map( A1 => n30658, A2 => n1726, B => n32988, ZN => 
                           n29610);
   U17555 : CLKBUF_X4 port map( I => n14290, Z => n33641);
   U17557 : NAND2_X2 port map( A1 => n30119, A2 => n19735, ZN => n26566);
   U17558 : NAND2_X2 port map( A1 => n7204, A2 => n7207, ZN => n21579);
   U17559 : XOR2_X1 port map( A1 => n9369, A2 => n22150, Z => n4589);
   U17560 : AOI22_X2 port map( A1 => n5912, A2 => n17261, B1 => n10188, B2 => 
                           n5913, ZN => n33041);
   U17561 : NOR2_X2 port map( A1 => n24004, A2 => n841, ZN => n10188);
   U17562 : NAND3_X1 port map( A1 => n5043, A2 => n28358, A3 => n15340, ZN => 
                           n32990);
   U17564 : NAND2_X1 port map( A1 => n23092, A2 => n13597, ZN => n33931);
   U17565 : NAND2_X2 port map( A1 => n12147, A2 => n12148, ZN => n20955);
   U17566 : NOR2_X1 port map( A1 => n23942, A2 => n11933, ZN => n15451);
   U17567 : XOR2_X1 port map( A1 => n283, A2 => n24801, Z => n24649);
   U17574 : NAND2_X2 port map( A1 => n6165, A2 => n30509, ZN => n24801);
   U17577 : XOR2_X1 port map( A1 => n27145, A2 => n24478, Z => n24551);
   U17580 : NAND2_X1 port map( A1 => n14184, A2 => n14724, ZN => n27145);
   U17581 : XOR2_X1 port map( A1 => n32991, A2 => n2739, Z => n2859);
   U17582 : XOR2_X1 port map( A1 => n20777, A2 => n10412, Z => n32991);
   U17585 : NAND3_X2 port map( A1 => n11952, A2 => n20042, A3 => n410, ZN => 
                           n16248);
   U17586 : NAND2_X1 port map( A1 => n27110, A2 => n1169, ZN => n20039);
   U17588 : XOR2_X1 port map( A1 => n1615, A2 => n1616, Z => n27110);
   U17589 : OAI22_X2 port map( A1 => n14547, A2 => n25708, B1 => n17092, B2 => 
                           n25752, ZN => n32992);
   U17591 : AOI22_X2 port map( A1 => n8587, A2 => n29207, B1 => n34059, B2 => 
                           n32993, ZN => n2790);
   U17594 : NAND2_X1 port map( A1 => n17522, A2 => n28607, ZN => n32993);
   U17597 : NAND3_X2 port map( A1 => n7276, A2 => n28995, A3 => n32994, ZN => 
                           n22274);
   U17599 : AOI22_X2 port map( A1 => n31935, A2 => n29242, B1 => n11330, B2 => 
                           n29314, ZN => n32995);
   U17600 : XOR2_X1 port map( A1 => n6348, A2 => n33465, Z => n5703);
   U17602 : XNOR2_X1 port map( A1 => n20859, A2 => n10081, ZN => n5518);
   U17604 : XOR2_X1 port map( A1 => n33234, A2 => n9141, Z => n10081);
   U17607 : AOI21_X2 port map( A1 => n20327, A2 => n20328, B => n1149, ZN => 
                           n32996);
   U17611 : INV_X2 port map( I => n28975, ZN => n32998);
   U17619 : NOR2_X2 port map( A1 => n24925, A2 => n24936, ZN => n24921);
   U17620 : AOI22_X2 port map( A1 => n13258, A2 => n25712, B1 => n13924, B2 => 
                           n12314, ZN => n33537);
   U17623 : XOR2_X1 port map( A1 => n30104, A2 => n32997, Z => n4682);
   U17624 : XOR2_X1 port map( A1 => n15508, A2 => n7511, Z => n32997);
   U17627 : OAI21_X1 port map( A1 => n5867, A2 => n10822, B => n25072, ZN => 
                           n5866);
   U17628 : NOR2_X2 port map( A1 => n13551, A2 => n13552, ZN => n24394);
   U17639 : AOI22_X2 port map( A1 => n5678, A2 => n1920, B1 => n2021, B2 => 
                           n845, ZN => n33244);
   U17642 : NAND2_X2 port map( A1 => n32999, A2 => n32998, ZN => n23672);
   U17644 : INV_X2 port map( I => n23942, ZN => n32999);
   U17645 : AOI22_X2 port map( A1 => n30725, A2 => n26882, B1 => n23871, B2 => 
                           n3571, ZN => n12841);
   U17646 : XOR2_X1 port map( A1 => n11349, A2 => n16708, Z => n5337);
   U17647 : OAI21_X2 port map( A1 => n2251, A2 => n2250, B => n12115, ZN => 
                           n11349);
   U17649 : NAND2_X2 port map( A1 => n33001, A2 => n34007, ZN => n27252);
   U17652 : NAND2_X2 port map( A1 => n8821, A2 => n8822, ZN => n18017);
   U17658 : OAI21_X2 port map( A1 => n8307, A2 => n5292, B => n33002, ZN => 
                           n25784);
   U17659 : XOR2_X1 port map( A1 => n33004, A2 => n572, Z => n10663);
   U17661 : XOR2_X1 port map( A1 => n358, A2 => n14908, Z => n33004);
   U17662 : INV_X1 port map( I => n33006, ZN => n11077);
   U17665 : NAND2_X2 port map( A1 => n32093, A2 => n33006, ZN => n33005);
   U17666 : NAND2_X2 port map( A1 => n33670, A2 => n16333, ZN => n33006);
   U17668 : XOR2_X1 port map( A1 => n20851, A2 => n20928, Z => n33332);
   U17670 : AOI21_X2 port map( A1 => n12782, A2 => n851, B => n33008, ZN => 
                           n23318);
   U17671 : OAI21_X2 port map( A1 => n22908, A2 => n29329, B => n22981, ZN => 
                           n22910);
   U17673 : INV_X2 port map( I => n33009, ZN => n17124);
   U17674 : AOI21_X2 port map( A1 => n1300, A2 => n22626, B => n33010, ZN => 
                           n33009);
   U17677 : XOR2_X1 port map( A1 => n13651, A2 => n16242, Z => n22000);
   U17678 : NAND2_X2 port map( A1 => n15698, A2 => n21873, ZN => n16242);
   U17682 : AOI21_X1 port map( A1 => n14524, A2 => n14525, B => n17139, ZN => 
                           n14151);
   U17685 : NAND2_X2 port map( A1 => n6178, A2 => n6177, ZN => n21626);
   U17694 : XOR2_X1 port map( A1 => n15517, A2 => n24616, Z => n24539);
   U17695 : NAND2_X2 port map( A1 => n33012, A2 => n24208, ZN => n24830);
   U17698 : OAI21_X2 port map( A1 => n2463, A2 => n24206, B => n33549, ZN => 
                           n33012);
   U17699 : XOR2_X1 port map( A1 => n27567, A2 => n33013, Z => n9789);
   U17705 : XOR2_X1 port map( A1 => n10519, A2 => n623, Z => n33013);
   U17709 : OAI21_X1 port map( A1 => n29335, A2 => n11895, B => n22553, ZN => 
                           n14776);
   U17712 : XOR2_X1 port map( A1 => n33014, A2 => n24754, Z => n7794);
   U17713 : XOR2_X1 port map( A1 => n9281, A2 => n27852, Z => n33014);
   U17715 : XNOR2_X1 port map( A1 => n24516, A2 => n25598, ZN => n33128);
   U17718 : NAND3_X2 port map( A1 => n27495, A2 => n2548, A3 => n33015, ZN => 
                           n2813);
   U17720 : XOR2_X1 port map( A1 => n20835, A2 => n16641, Z => n5630);
   U17726 : BUF_X2 port map( I => n31894, Z => n33016);
   U17732 : XOR2_X1 port map( A1 => n31860, A2 => n20765, Z => n17804);
   U17733 : XOR2_X1 port map( A1 => n28100, A2 => n532, Z => n33017);
   U17739 : NOR2_X2 port map( A1 => n8094, A2 => n33018, ZN => n33616);
   U17743 : OR2_X2 port map( A1 => n10327, A2 => n14238, Z => n25905);
   U17745 : XOR2_X1 port map( A1 => n33351, A2 => n28819, Z => n10327);
   U17749 : XOR2_X1 port map( A1 => n22148, A2 => n22318, Z => n10598);
   U17752 : NAND2_X2 port map( A1 => n21484, A2 => n21485, ZN => n22148);
   U17754 : NAND2_X1 port map( A1 => n28992, A2 => n25650, ZN => n33020);
   U17757 : AOI22_X2 port map( A1 => n29281, A2 => n7609, B1 => n10804, B2 => 
                           n10805, ZN => n29615);
   U17764 : XOR2_X1 port map( A1 => n24813, A2 => n7837, Z => n7838);
   U17766 : NAND2_X2 port map( A1 => n11388, A2 => n11387, ZN => n24813);
   U17768 : XOR2_X1 port map( A1 => n15384, A2 => n22036, Z => n17918);
   U17769 : AOI21_X2 port map( A1 => n21275, A2 => n21732, B => n15385, ZN => 
                           n15384);
   U17775 : XNOR2_X1 port map( A1 => n25224, A2 => n28898, ZN => n33579);
   U17779 : NOR3_X2 port map( A1 => n30758, A2 => n33021, A3 => n3934, ZN => 
                           n28077);
   U17780 : NAND3_X2 port map( A1 => n4823, A2 => n4822, A3 => n4824, ZN => 
                           n24257);
   U17784 : AOI22_X2 port map( A1 => n23954, A2 => n4991, B1 => n7140, B2 => 
                           n13998, ZN => n4822);
   U17787 : INV_X1 port map( I => n33023, ZN => n9446);
   U17791 : NAND3_X2 port map( A1 => n2348, A2 => n33945, A3 => n22344, ZN => 
                           n23009);
   U17794 : NOR2_X2 port map( A1 => n14594, A2 => n14595, ZN => n21964);
   U17797 : NAND2_X1 port map( A1 => n24162, A2 => n24340, ZN => n23781);
   U17803 : AOI22_X1 port map( A1 => n11069, A2 => n25292, B1 => n25196, B2 => 
                           n7081, ZN => n33024);
   U17804 : NAND2_X2 port map( A1 => n21680, A2 => n21681, ZN => n17362);
   U17805 : NAND3_X1 port map( A1 => n2342, A2 => n14540, A3 => n11626, ZN => 
                           n33686);
   U17808 : XOR2_X1 port map( A1 => n13041, A2 => n7653, Z => n21033);
   U17812 : NAND2_X2 port map( A1 => n13851, A2 => n30892, ZN => n7653);
   U17816 : NOR2_X2 port map( A1 => n33075, A2 => n29499, ZN => n9890);
   U17817 : NAND2_X2 port map( A1 => n9452, A2 => n9451, ZN => n4834);
   U17818 : XOR2_X1 port map( A1 => n33025, A2 => n10773, Z => n23188);
   U17821 : XOR2_X1 port map( A1 => n23368, A2 => n23247, Z => n33025);
   U17824 : OAI21_X1 port map( A1 => n14627, A2 => n1218, B => n17987, ZN => 
                           n33030);
   U17827 : XOR2_X1 port map( A1 => n24536, A2 => n33027, Z => n27490);
   U17828 : XOR2_X1 port map( A1 => n8413, A2 => n33028, Z => n33027);
   U17835 : NAND2_X2 port map( A1 => n33029, A2 => n21104, ZN => n15414);
   U17843 : OAI21_X2 port map( A1 => n26735, A2 => n26736, B => n21251, ZN => 
                           n33029);
   U17845 : NOR2_X1 port map( A1 => n22743, A2 => n16922, ZN => n30315);
   U17851 : XOR2_X1 port map( A1 => n29858, A2 => n17203, Z => n17204);
   U17856 : AOI21_X2 port map( A1 => n30050, A2 => n28502, B => n31999, ZN => 
                           n17079);
   U17857 : NAND2_X2 port map( A1 => n15584, A2 => n33043, ZN => n11041);
   U17860 : NOR2_X2 port map( A1 => n23037, A2 => n28415, ZN => n12444);
   U17867 : NAND2_X2 port map( A1 => n13412, A2 => n9964, ZN => n24044);
   U17869 : NAND2_X2 port map( A1 => n9589, A2 => n21480, ZN => n16269);
   U17873 : BUF_X2 port map( I => n16051, Z => n33032);
   U17874 : NOR2_X2 port map( A1 => n29246, A2 => n10955, ZN => n28855);
   U17881 : INV_X2 port map( I => n18235, ZN => n21692);
   U17882 : NAND2_X2 port map( A1 => n5628, A2 => n3286, ZN => n18235);
   U17886 : OAI21_X2 port map( A1 => n33034, A2 => n33033, B => n15149, ZN => 
                           n29975);
   U17900 : NOR2_X2 port map( A1 => n7238, A2 => n349, ZN => n33033);
   U17904 : INV_X2 port map( I => n21219, ZN => n33034);
   U17905 : NOR2_X2 port map( A1 => n29305, A2 => n654, ZN => n23705);
   U17912 : INV_X2 port map( I => n376, ZN => n654);
   U17913 : XOR2_X1 port map( A1 => n12579, A2 => n28031, Z => n376);
   U17916 : AOI21_X2 port map( A1 => n6704, A2 => n29905, B => n31048, ZN => 
                           n33035);
   U17917 : XOR2_X1 port map( A1 => n27875, A2 => n33036, Z => n11223);
   U17919 : XOR2_X1 port map( A1 => n33823, A2 => n23391, Z => n33036);
   U17928 : XOR2_X1 port map( A1 => n10460, A2 => n20692, Z => n20863);
   U17930 : NOR2_X2 port map( A1 => n30612, A2 => n33037, ZN => n16364);
   U17932 : NOR2_X1 port map( A1 => n20206, A2 => n20464, ZN => n20207);
   U17933 : INV_X2 port map( I => n33038, ZN => n15438);
   U17937 : XOR2_X1 port map( A1 => n3253, A2 => n12945, Z => n33038);
   U17941 : NAND2_X1 port map( A1 => n31522, A2 => n20257, ZN => n33820);
   U17944 : BUF_X2 port map( I => n881, Z => n33039);
   U17951 : XOR2_X1 port map( A1 => n1307, A2 => n3704, Z => n12627);
   U17960 : NOR2_X2 port map( A1 => n9088, A2 => n33483, ZN => n16237);
   U17961 : NAND2_X2 port map( A1 => n6926, A2 => n29008, ZN => n28028);
   U17967 : NAND2_X1 port map( A1 => n19986, A2 => n16, ZN => n19459);
   U17968 : XOR2_X1 port map( A1 => n11580, A2 => n14621, Z => n16);
   U17969 : XOR2_X1 port map( A1 => n22143, A2 => n22144, Z => n4627);
   U17978 : XNOR2_X1 port map( A1 => n4529, A2 => n4530, ZN => n33376);
   U17979 : OAI21_X2 port map( A1 => n16372, A2 => n18554, B => n9555, ZN => 
                           n19249);
   U17981 : XOR2_X1 port map( A1 => n22267, A2 => n22191, Z => n30250);
   U17982 : NAND3_X2 port map( A1 => n33228, A2 => n33229, A3 => n18956, ZN => 
                           n19558);
   U17983 : AOI21_X1 port map( A1 => n21228, A2 => n21305, B => n21132, ZN => 
                           n31728);
   U17986 : NAND2_X1 port map( A1 => n4834, A2 => n23086, ZN => n17669);
   U17987 : XOR2_X1 port map( A1 => n29501, A2 => n22102, Z => n22180);
   U17989 : NAND2_X2 port map( A1 => n5289, A2 => n18218, ZN => n13028);
   U17996 : NAND2_X2 port map( A1 => n31989, A2 => n5836, ZN => n5289);
   U17998 : XOR2_X1 port map( A1 => n26889, A2 => n33042, Z => n29075);
   U18002 : XOR2_X1 port map( A1 => n11996, A2 => n23236, Z => n33042);
   U18006 : NAND2_X2 port map( A1 => n10149, A2 => n21379, ZN => n10148);
   U18007 : OAI22_X2 port map( A1 => n20458, A2 => n20459, B1 => n20457, B2 => 
                           n3487, ZN => n21040);
   U18009 : NAND2_X2 port map( A1 => n9976, A2 => n9977, ZN => n24161);
   U18011 : NAND3_X2 port map( A1 => n33045, A2 => n24295, A3 => n15520, ZN => 
                           n6165);
   U18015 : NAND2_X2 port map( A1 => n7779, A2 => n5631, ZN => n33045);
   U18016 : NAND2_X2 port map( A1 => n30185, A2 => n11418, ZN => n2826);
   U18019 : OAI21_X2 port map( A1 => n24009, A2 => n17602, B => n33047, ZN => 
                           n9708);
   U18020 : AOI22_X2 port map( A1 => n22906, A2 => n33522, B1 => n989, B2 => 
                           n22907, ZN => n5343);
   U18025 : NOR2_X2 port map( A1 => n23069, A2 => n22865, ZN => n22906);
   U18033 : XOR2_X1 port map( A1 => n33048, A2 => n12717, Z => n27042);
   U18037 : XOR2_X1 port map( A1 => n23272, A2 => n15114, Z => n33048);
   U18039 : NAND3_X2 port map( A1 => n33049, A2 => n22701, A3 => n12646, ZN => 
                           n23417);
   U18041 : INV_X1 port map( I => n22960, ZN => n33050);
   U18043 : OR2_X1 port map( A1 => n29952, A2 => n33050, Z => n22701);
   U18045 : XOR2_X1 port map( A1 => n22084, A2 => n27943, Z => n27942);
   U18051 : AOI21_X1 port map( A1 => n22332, A2 => n8420, B => n28692, ZN => 
                           n29823);
   U18054 : XOR2_X1 port map( A1 => n33051, A2 => n23194, Z => n27441);
   U18058 : XOR2_X1 port map( A1 => n31567, A2 => n29012, Z => n33051);
   U18059 : NAND2_X2 port map( A1 => n10806, A2 => n33136, ZN => n28840);
   U18065 : NOR2_X2 port map( A1 => n16847, A2 => n19053, ZN => n2584);
   U18067 : XOR2_X1 port map( A1 => n27413, A2 => n27412, Z => n28702);
   U18074 : BUF_X2 port map( I => n24610, Z => n33053);
   U18077 : AND3_X1 port map( A1 => n24243, A2 => n28374, A3 => n24242, Z => 
                           n30000);
   U18078 : XOR2_X1 port map( A1 => n33054, A2 => n25373, Z => Ciphertext(100))
                           ;
   U18081 : NAND3_X2 port map( A1 => n25372, A2 => n25371, A3 => n25370, ZN => 
                           n33054);
   U18083 : OAI22_X2 port map( A1 => n33055, A2 => n1528, B1 => n11708, B2 => 
                           n29294, ZN => n31707);
   U18086 : INV_X4 port map( I => n6357, ZN => n21832);
   U18091 : XOR2_X1 port map( A1 => n23439, A2 => n10535, Z => n23277);
   U18093 : NAND2_X2 port map( A1 => n33728, A2 => n13559, ZN => n15212);
   U18094 : OAI21_X2 port map( A1 => n32493, A2 => n28669, B => n629, ZN => 
                           n33056);
   U18095 : XOR2_X1 port map( A1 => n20664, A2 => n5647, Z => n6701);
   U18097 : XOR2_X1 port map( A1 => n20849, A2 => n20658, Z => n20664);
   U18098 : XOR2_X1 port map( A1 => n23790, A2 => n33057, Z => n30398);
   U18099 : XOR2_X1 port map( A1 => n9907, A2 => n33058, Z => n33057);
   U18100 : XOR2_X1 port map( A1 => n33059, A2 => n25355, Z => Ciphertext(97));
   U18101 : OAI22_X1 port map( A1 => n25353, A2 => n25354, B1 => n25380, B2 => 
                           n25360, ZN => n33059);
   U18103 : OAI22_X1 port map( A1 => n24904, A2 => n24905, B1 => n24903, B2 => 
                           n10099, ZN => n33717);
   U18105 : NAND2_X2 port map( A1 => n33060, A2 => n23644, ZN => n24226);
   U18107 : NAND2_X1 port map( A1 => n3757, A2 => n34075, ZN => n33060);
   U18109 : INV_X2 port map( I => n24219, ZN => n1096);
   U18110 : OAI21_X2 port map( A1 => n14037, A2 => n23604, B => n32008, ZN => 
                           n24219);
   U18111 : NOR2_X2 port map( A1 => n23033, A2 => n6605, ZN => n23035);
   U18118 : INV_X2 port map( I => n11933, ZN => n33583);
   U18124 : XOR2_X1 port map( A1 => n1988, A2 => n33062, Z => n21455);
   U18132 : XOR2_X1 port map( A1 => n21034, A2 => n1986, Z => n33062);
   U18137 : XOR2_X1 port map( A1 => n33063, A2 => n25428, Z => Ciphertext(104))
                           ;
   U18139 : NAND2_X1 port map( A1 => n33546, A2 => n25427, ZN => n33063);
   U18143 : NAND2_X1 port map( A1 => n25425, A2 => n25455, ZN => n15500);
   U18146 : NAND2_X2 port map( A1 => n15783, A2 => n33064, ZN => n17948);
   U18148 : XOR2_X1 port map( A1 => n12714, A2 => n23408, Z => n3280);
   U18151 : NAND2_X2 port map( A1 => n3282, A2 => n3281, ZN => n12714);
   U18152 : OAI21_X2 port map( A1 => n8279, A2 => n24118, B => n33065, ZN => 
                           n8502);
   U18154 : NAND2_X2 port map( A1 => n24224, A2 => n24222, ZN => n33065);
   U18156 : XOR2_X1 port map( A1 => n8050, A2 => n24816, Z => n24593);
   U18162 : NAND2_X2 port map( A1 => n23610, A2 => n23609, ZN => n8050);
   U18164 : NAND2_X1 port map( A1 => n25383, A2 => n25561, ZN => n33068);
   U18167 : NOR3_X2 port map( A1 => n7776, A2 => n7775, A3 => n7232, ZN => 
                           n1877);
   U18174 : AOI22_X2 port map( A1 => n25925, A2 => n7701, B1 => n5411, B2 => 
                           n25923, ZN => n25927);
   U18177 : NAND2_X2 port map( A1 => n33071, A2 => n33070, ZN => n2558);
   U18189 : OAI21_X2 port map( A1 => n2563, A2 => n13402, B => n26965, ZN => 
                           n33070);
   U18193 : AND2_X1 port map( A1 => n16625, A2 => n33430, Z => n19801);
   U18194 : OAI21_X2 port map( A1 => n15905, A2 => n1337, B => n33209, ZN => 
                           n12221);
   U18195 : XOR2_X1 port map( A1 => n11324, A2 => n23165, Z => n33073);
   U18202 : AND2_X1 port map( A1 => n17770, A2 => n17787, Z => n33074);
   U18203 : XOR2_X1 port map( A1 => n19728, A2 => n32184, Z => n17954);
   U18209 : XOR2_X1 port map( A1 => n30943, A2 => n26751, Z => n19728);
   U18212 : XOR2_X1 port map( A1 => n20912, A2 => n20833, Z => n30107);
   U18213 : XOR2_X1 port map( A1 => n21040, A2 => n21018, Z => n20912);
   U18216 : OAI22_X2 port map( A1 => n17374, A2 => n2752, B1 => n1100, B2 => 
                           n23555, ZN => n33075);
   U18217 : XOR2_X1 port map( A1 => n23274, A2 => n1260, Z => n23459);
   U18220 : NOR2_X2 port map( A1 => n7921, A2 => n33076, ZN => n7762);
   U18228 : OAI22_X2 port map( A1 => n19862, A2 => n7920, B1 => n7922, B2 => 
                           n16694, ZN => n33076);
   U18233 : NAND2_X2 port map( A1 => n6123, A2 => n31148, ZN => n14953);
   U18234 : NOR2_X2 port map( A1 => n21719, A2 => n6718, ZN => n17716);
   U18236 : NAND2_X2 port map( A1 => n19249, A2 => n4436, ZN => n19248);
   U18239 : XOR2_X1 port map( A1 => n8921, A2 => n19585, Z => n4169);
   U18240 : XOR2_X1 port map( A1 => n1372, A2 => n19679, Z => n19585);
   U18243 : XOR2_X1 port map( A1 => n33077, A2 => n1402, Z => Ciphertext(153));
   U18244 : NOR2_X1 port map( A1 => n31833, A2 => n5784, ZN => n33077);
   U18250 : NOR2_X2 port map( A1 => n18006, A2 => n13846, ZN => n18470);
   U18253 : XOR2_X1 port map( A1 => n12674, A2 => n32889, Z => n10628);
   U18254 : NOR2_X2 port map( A1 => n31290, A2 => n31291, ZN => n20792);
   U18263 : NAND2_X2 port map( A1 => n9966, A2 => n9965, ZN => n27114);
   U18266 : XOR2_X1 port map( A1 => Plaintext(110), A2 => Key(110), Z => n33094
                           );
   U18268 : NAND2_X1 port map( A1 => n33069, A2 => n19120, ZN => n18956);
   U18273 : INV_X2 port map( I => n19118, ZN => n33078);
   U18274 : XOR2_X1 port map( A1 => n33079, A2 => n19686, Z => n17835);
   U18276 : XOR2_X1 port map( A1 => n31731, A2 => n25578, Z => n33079);
   U18279 : NAND2_X2 port map( A1 => n33080, A2 => n33732, ZN => n30130);
   U18280 : OAI22_X2 port map( A1 => n20035, A2 => n20034, B1 => n16243, B2 => 
                           n2795, ZN => n33080);
   U18287 : XOR2_X1 port map( A1 => n33081, A2 => n16672, Z => Ciphertext(15));
   U18288 : INV_X2 port map( I => n33082, ZN => n10438);
   U18290 : NAND2_X1 port map( A1 => n17977, A2 => n17978, ZN => n33431);
   U18293 : XOR2_X1 port map( A1 => n705, A2 => n24813, Z => n24797);
   U18296 : NOR2_X2 port map( A1 => n13217, A2 => n8204, ZN => n705);
   U18299 : AND2_X1 port map( A1 => n12221, A2 => n33083, Z => n17226);
   U18300 : XOR2_X1 port map( A1 => n22183, A2 => n27190, Z => n5976);
   U18301 : XOR2_X1 port map( A1 => n33084, A2 => n28462, Z => Ciphertext(52));
   U18302 : INV_X2 port map( I => n34128, ZN => n13073);
   U18304 : XOR2_X1 port map( A1 => n33358, A2 => n33085, Z => n34128);
   U18305 : XOR2_X1 port map( A1 => n26530, A2 => n20860, Z => n20668);
   U18312 : NOR2_X2 port map( A1 => n8959, A2 => n8960, ZN => n26530);
   U18313 : OAI21_X2 port map( A1 => n22671, A2 => n27357, B => n2311, ZN => 
                           n30297);
   U18315 : NOR2_X2 port map( A1 => n26663, A2 => n26784, ZN => n4254);
   U18316 : NAND2_X2 port map( A1 => n12496, A2 => n22503, ZN => n22530);
   U18319 : NOR3_X1 port map( A1 => n8902, A2 => n16798, A3 => n1204, ZN => 
                           n16793);
   U18322 : OR2_X1 port map( A1 => n3339, A2 => n25111, Z => n33314);
   U18323 : XOR2_X1 port map( A1 => n19409, A2 => n19398, Z => n6731);
   U18325 : NAND2_X2 port map( A1 => n10741, A2 => n10739, ZN => n19409);
   U18327 : XOR2_X1 port map( A1 => n15556, A2 => n29443, Z => n30094);
   U18342 : XOR2_X1 port map( A1 => n33086, A2 => n19496, Z => n3283);
   U18345 : XOR2_X1 port map( A1 => n29890, A2 => n1045, Z => n33086);
   U18349 : XOR2_X1 port map( A1 => n23459, A2 => n8974, Z => n8973);
   U18356 : NAND2_X2 port map( A1 => n25330, A2 => n6411, ZN => n25375);
   U18357 : NAND2_X2 port map( A1 => n33087, A2 => n25017, ZN => n25058);
   U18361 : OAI21_X2 port map( A1 => n11977, A2 => n14959, B => n14846, ZN => 
                           n33087);
   U18364 : NAND2_X2 port map( A1 => n9826, A2 => n9825, ZN => n24545);
   U18365 : XOR2_X1 port map( A1 => n17095, A2 => n17096, Z => n17094);
   U18366 : NAND3_X1 port map( A1 => n14232, A2 => n27577, A3 => n13720, ZN => 
                           n12883);
   U18373 : AOI21_X1 port map( A1 => n33310, A2 => n18085, B => n1182, ZN => 
                           n15928);
   U18374 : OR2_X1 port map( A1 => n1279, A2 => n4135, Z => n7946);
   U18375 : NAND3_X2 port map( A1 => n33089, A2 => n33750, A3 => n16225, ZN => 
                           n21974);
   U18376 : NAND2_X2 port map( A1 => n31551, A2 => n630, ZN => n33089);
   U18377 : NAND2_X2 port map( A1 => n263, A2 => n262, ZN => n7293);
   U18392 : NOR2_X2 port map( A1 => n1557, A2 => n26328, ZN => n34099);
   U18393 : OAI21_X2 port map( A1 => n33441, A2 => n13978, B => n17136, ZN => 
                           n33527);
   U18395 : XOR2_X1 port map( A1 => n23375, A2 => n22970, Z => n23517);
   U18401 : NOR2_X2 port map( A1 => n27566, A2 => n7945, ZN => n23375);
   U18402 : NAND2_X2 port map( A1 => n21163, A2 => n11734, ZN => n13593);
   U18403 : XOR2_X1 port map( A1 => n33090, A2 => n24445, Z => n27526);
   U18412 : XOR2_X1 port map( A1 => n24691, A2 => n8050, Z => n24525);
   U18415 : NAND3_X2 port map( A1 => n11964, A2 => n13630, A3 => n13628, ZN => 
                           n25988);
   U18417 : INV_X2 port map( I => n33092, ZN => n9064);
   U18419 : XNOR2_X1 port map( A1 => n33636, A2 => n7640, ZN => n33092);
   U18422 : NOR2_X2 port map( A1 => n29769, A2 => n19118, ZN => n19119);
   U18423 : NAND2_X2 port map( A1 => n926, A2 => n6520, ZN => n10730);
   U18428 : XOR2_X1 port map( A1 => n12454, A2 => n24836, Z => n30493);
   U18432 : INV_X2 port map( I => n12748, ZN => n26778);
   U18439 : NAND2_X2 port map( A1 => n14501, A2 => n24059, ZN => n13470);
   U18444 : NAND3_X2 port map( A1 => n6354, A2 => n7069, A3 => n13306, ZN => 
                           n14501);
   U18446 : XOR2_X1 port map( A1 => n4312, A2 => n287, Z => n9375);
   U18448 : OR2_X1 port map( A1 => n12551, A2 => n3222, Z => n24071);
   U18459 : XOR2_X1 port map( A1 => n30131, A2 => n4682, Z => n25696);
   U18466 : AOI22_X2 port map( A1 => n28585, A2 => n33011, B1 => n23747, B2 => 
                           n16628, ZN => n23748);
   U18468 : INV_X1 port map( I => n686, ZN => n33095);
   U18469 : OR2_X1 port map( A1 => n22999, A2 => n16297, Z => n7219);
   U18472 : NOR2_X2 port map( A1 => n17922, A2 => n33096, ZN => n26883);
   U18474 : OR2_X1 port map( A1 => n33766, A2 => n31958, Z => n14209);
   U18479 : BUF_X2 port map( I => n16569, Z => n33098);
   U18480 : XOR2_X1 port map( A1 => n15297, A2 => n28710, Z => n34118);
   U18481 : NOR2_X2 port map( A1 => n20589, A2 => n31967, ZN => n15638);
   U18482 : XOR2_X1 port map( A1 => n33099, A2 => n6620, Z => n33617);
   U18483 : XOR2_X1 port map( A1 => n33100, A2 => n30917, Z => n33099);
   U18486 : XOR2_X1 port map( A1 => n3964, A2 => n19341, Z => n31414);
   U18489 : NOR2_X2 port map( A1 => n19162, A2 => n19161, ZN => n19341);
   U18490 : NAND3_X2 port map( A1 => n17692, A2 => n21747, A3 => n21746, ZN => 
                           n4034);
   U18493 : AOI21_X2 port map( A1 => n29632, A2 => n8176, B => n21968, ZN => 
                           n33115);
   U18507 : XOR2_X1 port map( A1 => n20720, A2 => n31966, Z => n20757);
   U18511 : NOR2_X2 port map( A1 => n13597, A2 => n22964, ZN => n12662);
   U18512 : XOR2_X1 port map( A1 => n20558, A2 => n20718, Z => n10391);
   U18513 : OAI22_X2 port map( A1 => n7426, A2 => n33105, B1 => n7427, B2 => 
                           n15740, ZN => n16315);
   U18514 : BUF_X2 port map( I => n4568, Z => n33106);
   U18516 : INV_X4 port map( I => n8130, ZN => n1350);
   U18518 : NAND2_X1 port map( A1 => n14545, A2 => n8130, ZN => n33107);
   U18520 : NOR2_X1 port map( A1 => n15340, A2 => n5578, ZN => n5173);
   U18527 : OAI21_X1 port map( A1 => n33432, A2 => n19275, B => n33108, ZN => 
                           n18971);
   U18536 : XOR2_X1 port map( A1 => n33109, A2 => n10332, Z => n29828);
   U18540 : XOR2_X1 port map( A1 => n20802, A2 => n25311, Z => n33109);
   U18541 : XOR2_X1 port map( A1 => n4321, A2 => n2388, Z => n29028);
   U18549 : NOR3_X2 port map( A1 => n6024, A2 => n11581, A3 => n6023, ZN => 
                           n4321);
   U18557 : NAND2_X1 port map( A1 => n21530, A2 => n29980, ZN => n6231);
   U18562 : NOR2_X2 port map( A1 => n28299, A2 => n28298, ZN => n21530);
   U18567 : XOR2_X1 port map( A1 => n2349, A2 => n1129, Z => n22187);
   U18578 : OAI21_X2 port map( A1 => n33113, A2 => n33112, B => n2574, ZN => 
                           n8391);
   U18584 : NOR2_X1 port map( A1 => n1632, A2 => n17439, ZN => n33112);
   U18587 : INV_X2 port map( I => n33114, ZN => n23706);
   U18591 : XNOR2_X1 port map( A1 => n17826, A2 => n33490, ZN => n33114);
   U18594 : AND2_X1 port map( A1 => n29980, A2 => n21530, Z => n16952);
   U18603 : NAND2_X2 port map( A1 => n14717, A2 => n12221, ZN => n27595);
   U18606 : XOR2_X1 port map( A1 => n24852, A2 => n8480, Z => n24427);
   U18608 : NAND3_X2 port map( A1 => n11962, A2 => n3021, A3 => n24071, ZN => 
                           n24852);
   U18610 : NOR2_X1 port map( A1 => n31664, A2 => n24069, ZN => n31663);
   U18612 : XOR2_X1 port map( A1 => n15588, A2 => n24600, Z => n1441);
   U18614 : NAND2_X1 port map( A1 => n28414, A2 => n27697, ZN => n26800);
   U18615 : NAND2_X2 port map( A1 => n2934, A2 => n19807, ZN => n27697);
   U18617 : XOR2_X1 port map( A1 => n23402, A2 => n27552, Z => n33606);
   U18621 : NOR2_X2 port map( A1 => n23052, A2 => n22798, ZN => n6099);
   U18623 : XOR2_X1 port map( A1 => n23415, A2 => n23414, Z => n33118);
   U18625 : XOR2_X1 port map( A1 => n24569, A2 => n15438, Z => n10196);
   U18627 : OAI21_X2 port map( A1 => n13642, A2 => n13641, B => n33119, ZN => 
                           n13637);
   U18628 : NOR2_X2 port map( A1 => n33786, A2 => n4350, ZN => n4349);
   U18630 : XOR2_X1 port map( A1 => n5904, A2 => n23292, Z => n33465);
   U18637 : OR2_X1 port map( A1 => n17503, A2 => n31943, Z => n13231);
   U18639 : XOR2_X1 port map( A1 => n12252, A2 => n23196, Z => n23451);
   U18650 : NAND2_X2 port map( A1 => n22767, A2 => n22768, ZN => n12252);
   U18653 : XOR2_X1 port map( A1 => n33121, A2 => n11822, Z => n27570);
   U18660 : XOR2_X1 port map( A1 => n31611, A2 => n23296, Z => n33121);
   U18661 : OAI21_X2 port map( A1 => n8315, A2 => n14091, B => n6119, ZN => 
                           n33122);
   U18663 : NAND2_X2 port map( A1 => n33708, A2 => n8463, ZN => n22232);
   U18664 : XOR2_X1 port map( A1 => n19625, A2 => n16429, Z => n17540);
   U18665 : NOR2_X2 port map( A1 => n27718, A2 => n19077, ZN => n19625);
   U18666 : NAND2_X2 port map( A1 => n21083, A2 => n7620, ZN => n12827);
   U18669 : XOR2_X1 port map( A1 => n5185, A2 => n31887, Z => n33153);
   U18670 : NAND2_X2 port map( A1 => n16297, A2 => n22999, ZN => n5682);
   U18672 : XOR2_X1 port map( A1 => n10005, A2 => n13873, Z => n10004);
   U18680 : NAND2_X2 port map( A1 => n33125, A2 => n33859, ZN => n11755);
   U18687 : AOI21_X2 port map( A1 => n21312, A2 => n13194, B => n34159, ZN => 
                           n33125);
   U18688 : NAND2_X1 port map( A1 => n9917, A2 => n17044, ZN => n9916);
   U18690 : NAND2_X2 port map( A1 => n21390, A2 => n6179, ZN => n6177);
   U18691 : NAND2_X1 port map( A1 => n16716, A2 => n22889, ZN => n33126);
   U18693 : XOR2_X1 port map( A1 => n28448, A2 => n33127, Z => n30526);
   U18696 : XOR2_X1 port map( A1 => n24418, A2 => n33128, Z => n33127);
   U18701 : AOI21_X2 port map( A1 => n9689, A2 => n33515, B => n33129, ZN => 
                           n12902);
   U18705 : NOR3_X2 port map( A1 => n33515, A2 => n13300, A3 => n1154, ZN => 
                           n33129);
   U18712 : XOR2_X1 port map( A1 => n15823, A2 => n33130, Z => n10800);
   U18714 : XOR2_X1 port map( A1 => n31584, A2 => n31884, Z => n33130);
   U18717 : OAI21_X1 port map( A1 => n33144, A2 => n14335, B => n33722, ZN => 
                           n3289);
   U18720 : INV_X2 port map( I => n8166, ZN => n14335);
   U18721 : XOR2_X1 port map( A1 => n33866, A2 => n1436, Z => n8166);
   U18722 : NAND2_X2 port map( A1 => n33131, A2 => n15624, ZN => n31793);
   U18723 : NAND2_X2 port map( A1 => n30561, A2 => n31149, ZN => n33131);
   U18724 : NAND2_X2 port map( A1 => n28253, A2 => n30826, ZN => n13545);
   U18726 : AOI22_X2 port map( A1 => n33180, A2 => n22483, B1 => n9022, B2 => 
                           n22297, ZN => n4221);
   U18728 : OAI21_X1 port map( A1 => n21705, A2 => n26782, B => n2643, ZN => 
                           n26479);
   U18731 : INV_X2 port map( I => n33134, ZN => n10325);
   U18732 : XNOR2_X1 port map( A1 => Plaintext(4), A2 => Key(4), ZN => n33134);
   U18734 : NAND3_X1 port map( A1 => n31977, A2 => n33277, A3 => n24611, ZN => 
                           n24613);
   U18739 : OAI22_X2 port map( A1 => n23811, A2 => n23559, B1 => n23558, B2 => 
                           n23947, ZN => n23560);
   U18743 : NAND2_X2 port map( A1 => n33135, A2 => n18117, ZN => n5306);
   U18745 : NOR2_X2 port map( A1 => n23007, A2 => n23013, ZN => n10528);
   U18754 : OAI22_X2 port map( A1 => n22348, A2 => n996, B1 => n7965, B2 => 
                           n22450, ZN => n23013);
   U18758 : OAI21_X1 port map( A1 => n8757, A2 => n21054, B => n33137, ZN => 
                           n33142);
   U18759 : NAND2_X1 port map( A1 => n15323, A2 => n6402, ZN => n33138);
   U18761 : XOR2_X1 port map( A1 => n20690, A2 => n21047, Z => n5775);
   U18763 : INV_X2 port map( I => n30191, ZN => n24268);
   U18768 : NAND3_X2 port map( A1 => n31691, A2 => n31690, A3 => n11670, ZN => 
                           n30191);
   U18769 : NAND3_X2 port map( A1 => n2167, A2 => n10152, A3 => n31173, ZN => 
                           n26363);
   U18771 : NAND2_X2 port map( A1 => n33797, A2 => n33694, ZN => n10312);
   U18775 : XOR2_X1 port map( A1 => n2820, A2 => n2819, Z => n31101);
   U18776 : NOR2_X1 port map( A1 => n23694, A2 => n28367, ZN => n33226);
   U18779 : OAI21_X2 port map( A1 => n9233, A2 => n18172, B => n33140, ZN => 
                           n29763);
   U18781 : AOI22_X2 port map( A1 => n33141, A2 => n17238, B1 => n12249, B2 => 
                           n12497, ZN => n19463);
   U18782 : OAI21_X2 port map( A1 => n12249, A2 => n12500, B => n18135, ZN => 
                           n33141);
   U18788 : NAND2_X2 port map( A1 => n33142, A2 => n31848, ZN => n21719);
   U18789 : AOI22_X2 port map( A1 => n21771, A2 => n26904, B1 => n2718, B2 => 
                           n38, ZN => n4219);
   U18790 : BUF_X4 port map( I => n23499, Z => n33293);
   U18802 : BUF_X2 port map( I => n18919, Z => n33143);
   U18805 : BUF_X2 port map( I => n23813, Z => n33144);
   U18809 : NAND2_X1 port map( A1 => n11983, A2 => n31854, ZN => n13575);
   U18815 : NAND2_X2 port map( A1 => n22011, A2 => n26394, ZN => n31854);
   U18817 : INV_X2 port map( I => n7515, ZN => n715);
   U18818 : NAND2_X2 port map( A1 => n26380, A2 => n1859, ZN => n7515);
   U18820 : XOR2_X1 port map( A1 => n4732, A2 => n32860, Z => n23312);
   U18822 : OAI22_X2 port map( A1 => n29789, A2 => n29922, B1 => n33690, B2 => 
                           n28263, ZN => n14540);
   U18829 : XOR2_X1 port map( A1 => n28323, A2 => n30041, Z => n29643);
   U18839 : OAI21_X1 port map( A1 => n31661, A2 => n31662, B => n28070, ZN => 
                           n33145);
   U18848 : NOR2_X1 port map( A1 => n31932, A2 => n10197, ZN => n12213);
   U18852 : NAND3_X1 port map( A1 => n8206, A2 => n32240, A3 => n20534, ZN => 
                           n20354);
   U18856 : XOR2_X1 port map( A1 => n5472, A2 => n20813, Z => n33508);
   U18861 : NAND2_X2 port map( A1 => n2316, A2 => n2318, ZN => n5472);
   U18865 : XNOR2_X1 port map( A1 => n5742, A2 => n25054, ZN => n33960);
   U18871 : NOR2_X2 port map( A1 => n9201, A2 => n20067, ZN => n11052);
   U18874 : NOR2_X1 port map( A1 => n31263, A2 => n25452, ZN => n25420);
   U18875 : XOR2_X1 port map( A1 => n6863, A2 => n6862, Z => n2557);
   U18876 : NOR2_X1 port map( A1 => n28343, A2 => n31357, ZN => n23773);
   U18879 : NAND2_X2 port map( A1 => n30990, A2 => n26579, ZN => n5454);
   U18880 : NOR2_X1 port map( A1 => n8912, A2 => n16745, ZN => n22335);
   U18881 : XOR2_X1 port map( A1 => n13347, A2 => n23274, Z => n17565);
   U18883 : NAND2_X2 port map( A1 => n28355, A2 => n29114, ZN => n23274);
   U18884 : NAND4_X2 port map( A1 => n7091, A2 => n7094, A3 => n23988, A4 => 
                           n7095, ZN => n10331);
   U18886 : OAI21_X1 port map( A1 => n2066, A2 => n31964, B => n1288, ZN => 
                           n7819);
   U18888 : BUF_X2 port map( I => n30997, Z => n33150);
   U18889 : XOR2_X1 port map( A1 => n22173, A2 => n33151, Z => n28000);
   U18891 : XOR2_X1 port map( A1 => n33152, A2 => n23447, Z => n17352);
   U18894 : OR2_X1 port map( A1 => n18919, A2 => n18626, Z => n33965);
   U18896 : BUF_X2 port map( I => n27741, Z => n33154);
   U18899 : NAND2_X2 port map( A1 => n33156, A2 => n28340, ZN => n21569);
   U18903 : NOR2_X2 port map( A1 => n4284, A2 => n4283, ZN => n33156);
   U18908 : NAND2_X2 port map( A1 => n14485, A2 => n14486, ZN => n20992);
   U18909 : XOR2_X1 port map( A1 => n12609, A2 => n33157, Z => n7566);
   U18914 : XOR2_X1 port map( A1 => n8284, A2 => n32889, Z => n33157);
   U18924 : NOR2_X1 port map( A1 => n25060, A2 => n25062, ZN => n3122);
   U18925 : OAI21_X2 port map( A1 => n20055, A2 => n8616, B => n33158, ZN => 
                           n17715);
   U18927 : NAND2_X2 port map( A1 => n3005, A2 => n8616, ZN => n33158);
   U18930 : XOR2_X1 port map( A1 => n33756, A2 => n9464, Z => n4727);
   U18932 : XOR2_X1 port map( A1 => n29481, A2 => n31043, Z => n9464);
   U18937 : OAI21_X1 port map( A1 => n31142, A2 => n25444, B => n31141, ZN => 
                           n33159);
   U18942 : AND2_X1 port map( A1 => n15623, A2 => n34167, Z => n16540);
   U18943 : NAND3_X2 port map( A1 => n7282, A2 => n7176, A3 => n19245, ZN => 
                           n7109);
   U18945 : NAND2_X2 port map( A1 => n3183, A2 => n22848, ZN => n22937);
   U18949 : NAND2_X2 port map( A1 => n3187, A2 => n2252, ZN => n3183);
   U18959 : XOR2_X1 port map( A1 => n15823, A2 => n29482, Z => n27413);
   U18964 : XOR2_X1 port map( A1 => n30749, A2 => n20670, Z => n15823);
   U18966 : OAI22_X2 port map( A1 => n4505, A2 => n4506, B1 => n18865, B2 => 
                           n18864, ZN => n30865);
   U18969 : XOR2_X1 port map( A1 => n14819, A2 => n23253, Z => n23184);
   U18971 : NAND3_X2 port map( A1 => n22943, A2 => n60, A3 => n22942, ZN => 
                           n14819);
   U18978 : XOR2_X1 port map( A1 => n14584, A2 => n23119, Z => n6848);
   U18991 : XOR2_X1 port map( A1 => n24651, A2 => n24653, Z => n33161);
   U18996 : NOR3_X1 port map( A1 => n25996, A2 => n652, A3 => n14193, ZN => 
                           n27233);
   U19005 : NOR2_X2 port map( A1 => n33162, A2 => n3947, ZN => n1995);
   U19007 : NAND2_X1 port map( A1 => n11563, A2 => n24244, ZN => n33162);
   U19013 : XOR2_X1 port map( A1 => n18125, A2 => n19783, Z => n30757);
   U19016 : INV_X2 port map( I => n19708, ZN => n18125);
   U19024 : NOR2_X2 port map( A1 => n16907, A2 => n16909, ZN => n19708);
   U19027 : INV_X1 port map( I => n33163, ZN => n12201);
   U19030 : NOR2_X1 port map( A1 => n24970, A2 => n3843, ZN => n33163);
   U19031 : NAND2_X2 port map( A1 => n33666, A2 => n30928, ZN => n3843);
   U19032 : NOR2_X1 port map( A1 => n4750, A2 => n8365, ZN => n22879);
   U19039 : XOR2_X1 port map( A1 => n23331, A2 => n23256, Z => n30156);
   U19040 : XOR2_X1 port map( A1 => n23438, A2 => n23534, Z => n23256);
   U19048 : NAND2_X2 port map( A1 => n28489, A2 => n33164, ZN => n31129);
   U19053 : NAND2_X2 port map( A1 => n5770, A2 => n5771, ZN => n33164);
   U19055 : OAI21_X2 port map( A1 => n19036, A2 => n26603, B => n33168, ZN => 
                           n5418);
   U19056 : NOR2_X2 port map( A1 => n29962, A2 => n29963, ZN => n33168);
   U19057 : OAI21_X2 port map( A1 => n28136, A2 => n16451, B => n33169, ZN => 
                           n11705);
   U19058 : NAND2_X1 port map( A1 => n28530, A2 => n26570, ZN => n29934);
   U19063 : XOR2_X1 port map( A1 => n33170, A2 => n5722, Z => n6894);
   U19067 : XOR2_X1 port map( A1 => n5724, A2 => n21045, Z => n33170);
   U19070 : NAND2_X1 port map( A1 => n24286, A2 => n17361, ZN => n29576);
   U19074 : XOR2_X1 port map( A1 => n16200, A2 => n23312, Z => n11143);
   U19087 : AOI21_X2 port map( A1 => n31978, A2 => n29552, B => n33172, ZN => 
                           n2215);
   U19090 : NOR3_X2 port map( A1 => n2217, A2 => n21628, A3 => n33992, ZN => 
                           n33172);
   U19093 : NAND2_X2 port map( A1 => n16413, A2 => n6939, ZN => n14547);
   U19095 : NAND2_X2 port map( A1 => n33173, A2 => n28506, ZN => n24084);
   U19098 : AOI21_X2 port map( A1 => n14155, A2 => n28676, B => n33174, ZN => 
                           n33173);
   U19119 : INV_X1 port map( I => n23724, ZN => n33174);
   U19122 : NAND2_X1 port map( A1 => n14598, A2 => n21341, ZN => n33417);
   U19129 : XOR2_X1 port map( A1 => n23429, A2 => n16053, Z => n4792);
   U19130 : NAND2_X2 port map( A1 => n31365, A2 => n30433, ZN => n16053);
   U19131 : INV_X2 port map( I => n33175, ZN => n28329);
   U19138 : XNOR2_X1 port map( A1 => n2024, A2 => n30190, ZN => n33175);
   U19139 : XOR2_X1 port map( A1 => n28999, A2 => n24388, Z => n34073);
   U19140 : XOR2_X1 port map( A1 => n24478, A2 => n24622, Z => n24388);
   U19143 : NAND4_X1 port map( A1 => n14637, A2 => n14763, A3 => n16578, A4 => 
                           n14635, ZN => n33701);
   U19144 : AOI21_X2 port map( A1 => n28330, A2 => n5178, B => n7047, ZN => 
                           n11466);
   U19147 : XOR2_X1 port map( A1 => n10960, A2 => n30098, Z => n21970);
   U19152 : INV_X1 port map( I => n15559, ZN => n33215);
   U19154 : NOR2_X2 port map( A1 => n22732, A2 => n22730, ZN => n3668);
   U19155 : AOI21_X2 port map( A1 => n21902, A2 => n22488, B => n31551, ZN => 
                           n22732);
   U19156 : NOR2_X2 port map( A1 => n23326, A2 => n33177, ZN => n31772);
   U19163 : OAI21_X2 port map( A1 => n32006, A2 => n27219, B => n33178, ZN => 
                           n33177);
   U19165 : NAND2_X2 port map( A1 => n23322, A2 => n27219, ZN => n33178);
   U19167 : NOR2_X2 port map( A1 => n33179, A2 => n4453, ZN => n23143);
   U19170 : AOI22_X1 port map( A1 => n25008, A2 => n24998, B1 => n15016, B2 => 
                           n15078, ZN => n25000);
   U19171 : NAND2_X2 port map( A1 => n10612, A2 => n9737, ZN => n22372);
   U19173 : XOR2_X1 port map( A1 => n2192, A2 => n1482, Z => n1481);
   U19178 : XOR2_X1 port map( A1 => n2198, A2 => n16331, Z => n2192);
   U19179 : AOI21_X2 port map( A1 => n16295, A2 => n2778, B => n6295, ZN => 
                           n15808);
   U19180 : NAND2_X2 port map( A1 => n18711, A2 => n328, ZN => n2778);
   U19182 : XOR2_X1 port map( A1 => n11781, A2 => n33181, Z => n11780);
   U19183 : XOR2_X1 port map( A1 => n6454, A2 => n2896, Z => n33181);
   U19188 : NOR2_X2 port map( A1 => n15054, A2 => n25247, ZN => n33353);
   U19189 : INV_X2 port map( I => n5544, ZN => n25247);
   U19193 : NAND3_X2 port map( A1 => n28117, A2 => n2214, A3 => n17925, ZN => 
                           n5544);
   U19195 : OR2_X1 port map( A1 => n15790, A2 => n33182, Z => n23999);
   U19197 : OR2_X1 port map( A1 => n33183, A2 => n22443, Z => n6837);
   U19203 : XOR2_X1 port map( A1 => n22282, A2 => n3395, Z => n33202);
   U19204 : XOR2_X1 port map( A1 => n22274, A2 => n22028, Z => n22282);
   U19207 : NOR2_X2 port map( A1 => n31640, A2 => n25062, ZN => n25041);
   U19210 : XOR2_X1 port map( A1 => n17552, A2 => n19536, Z => n11251);
   U19212 : NAND2_X1 port map( A1 => n25644, A2 => n34094, ZN => n25646);
   U19215 : OAI22_X2 port map( A1 => n33185, A2 => n1962, B1 => n20551, B2 => 
                           n26343, ZN => n21009);
   U19219 : NOR3_X2 port map( A1 => n20550, A2 => n31232, A3 => n125, ZN => 
                           n33185);
   U19221 : OAI21_X2 port map( A1 => n14437, A2 => n13796, B => n33186, ZN => 
                           n19241);
   U19225 : OAI21_X2 port map( A1 => n1054, A2 => n26603, B => n13796, ZN => 
                           n33186);
   U19227 : AOI22_X1 port map( A1 => n25432, A2 => n11640, B1 => n25453, B2 => 
                           n25433, ZN => n25434);
   U19229 : XNOR2_X1 port map( A1 => n231, A2 => n7619, ZN => n33264);
   U19230 : NAND2_X2 port map( A1 => n33980, A2 => n29801, ZN => n5462);
   U19231 : NOR2_X2 port map( A1 => n27973, A2 => n33188, ZN => n27504);
   U19241 : OAI22_X2 port map( A1 => n17438, A2 => n21060, B1 => n21222, B2 => 
                           n21061, ZN => n33188);
   U19244 : INV_X2 port map( I => n33189, ZN => n11063);
   U19248 : XNOR2_X1 port map( A1 => n26769, A2 => n4263, ZN => n33189);
   U19254 : NAND3_X2 port map( A1 => n33191, A2 => n22299, A3 => n33190, ZN => 
                           n13622);
   U19257 : NAND2_X1 port map( A1 => n8136, A2 => n10757, ZN => n33191);
   U19258 : NOR2_X2 port map( A1 => n21566, A2 => n17274, ZN => n33611);
   U19260 : NAND2_X2 port map( A1 => n33192, A2 => n1788, ZN => n1787);
   U19265 : AOI21_X2 port map( A1 => n1774, A2 => n20200, B => n1789, ZN => 
                           n33193);
   U19267 : XOR2_X1 port map( A1 => n8581, A2 => n11691, Z => n20762);
   U19275 : NOR2_X2 port map( A1 => n13573, A2 => n13572, ZN => n8581);
   U19280 : AOI21_X1 port map( A1 => n18737, A2 => n12166, B => n16287, ZN => 
                           n13026);
   U19286 : NAND2_X2 port map( A1 => n33195, A2 => n33194, ZN => n14027);
   U19289 : NOR2_X1 port map( A1 => n17240, A2 => n24975, ZN => n26020);
   U19291 : NOR2_X1 port map( A1 => n14812, A2 => n14811, ZN => n6637);
   U19294 : NAND2_X2 port map( A1 => n17253, A2 => n17254, ZN => n14812);
   U19301 : AND2_X2 port map( A1 => n14001, A2 => n10371, Z => n24351);
   U19304 : NOR2_X2 port map( A1 => n23877, A2 => n23878, ZN => n15245);
   U19306 : NOR2_X1 port map( A1 => n3565, A2 => n25763, ZN => n24448);
   U19308 : XOR2_X1 port map( A1 => n24619, A2 => n5253, Z => n8656);
   U19309 : NAND2_X2 port map( A1 => n6982, A2 => n33197, ZN => n7198);
   U19310 : INV_X2 port map( I => n31942, ZN => n17501);
   U19312 : NAND2_X2 port map( A1 => n33863, A2 => n92, ZN => n23005);
   U19319 : XOR2_X1 port map( A1 => n23454, A2 => n7520, Z => n28493);
   U19324 : NAND2_X1 port map( A1 => n33198, A2 => n14164, ZN => n15207);
   U19325 : NAND2_X1 port map( A1 => n23578, A2 => n16981, ZN => n33198);
   U19330 : NAND2_X1 port map( A1 => n11898, A2 => n24610, ZN => n33199);
   U19332 : XOR2_X1 port map( A1 => n1003, A2 => n22028, Z => n22275);
   U19336 : XOR2_X1 port map( A1 => n33201, A2 => n33200, Z => n30042);
   U19337 : XOR2_X1 port map( A1 => n14733, A2 => n6833, Z => n33201);
   U19343 : AND2_X1 port map( A1 => n29158, A2 => n28924, Z => n33865);
   U19349 : NAND3_X1 port map( A1 => n10295, A2 => n4750, A3 => n5274, ZN => 
                           n27544);
   U19353 : XOR2_X1 port map( A1 => n33203, A2 => n16060, Z => n22285);
   U19354 : NAND2_X2 port map( A1 => n1874, A2 => n11595, ZN => n7066);
   U19355 : NAND2_X2 port map( A1 => n5593, A2 => n7103, ZN => n13347);
   U19357 : XOR2_X1 port map( A1 => n26872, A2 => n34146, Z => n9690);
   U19361 : XOR2_X1 port map( A1 => n4285, A2 => n22138, Z => n12980);
   U19368 : NOR2_X2 port map( A1 => n3578, A2 => n3579, ZN => n4285);
   U19370 : AOI22_X1 port map( A1 => n6830, A2 => n6829, B1 => n6828, B2 => 
                           n1075, ZN => n6827);
   U19373 : XOR2_X1 port map( A1 => n8885, A2 => n32083, Z => n21248);
   U19374 : XOR2_X1 port map( A1 => n20837, A2 => n33204, Z => n30778);
   U19381 : INV_X2 port map( I => n21007, ZN => n33204);
   U19390 : NAND2_X2 port map( A1 => n17431, A2 => n9076, ZN => n11619);
   U19404 : NAND2_X2 port map( A1 => n33262, A2 => n30105, ZN => n15806);
   U19405 : OAI21_X1 port map( A1 => n18738, A2 => n33208, B => n33207, ZN => 
                           n18736);
   U19407 : OAI21_X1 port map( A1 => n26369, A2 => n11792, B => n21233, ZN => 
                           n33209);
   U19410 : XOR2_X1 port map( A1 => n33210, A2 => n24798, Z => n18155);
   U19412 : XOR2_X1 port map( A1 => n24797, A2 => n31440, Z => n33210);
   U19415 : NAND2_X2 port map( A1 => n33212, A2 => n33211, ZN => n15787);
   U19419 : AOI22_X1 port map( A1 => n18907, A2 => n1056, B1 => n12128, B2 => 
                           n10227, ZN => n33211);
   U19430 : NAND2_X1 port map( A1 => n2517, A2 => n764, ZN => n33212);
   U19431 : XOR2_X1 port map( A1 => n33213, A2 => n32930, Z => n31296);
   U19439 : XOR2_X1 port map( A1 => n19487, A2 => n19737, Z => n33213);
   U19440 : XOR2_X1 port map( A1 => n33214, A2 => n30951, Z => n29064);
   U19451 : INV_X4 port map( I => n9575, ZN => n33382);
   U19453 : XOR2_X1 port map( A1 => n15, A2 => n2989, Z => n1986);
   U19455 : NAND2_X2 port map( A1 => n21240, A2 => n11601, ZN => n13152);
   U19456 : OAI22_X2 port map( A1 => n21431, A2 => n21070, B1 => n21241, B2 => 
                           n606, ZN => n21240);
   U19457 : NAND2_X2 port map( A1 => n31418, A2 => n27411, ZN => n4580);
   U19461 : INV_X1 port map( I => n28177, ZN => n23424);
   U19462 : INV_X2 port map( I => n3260, ZN => n10294);
   U19466 : OAI22_X2 port map( A1 => n9711, A2 => n9677, B1 => n9710, B2 => 
                           n9709, ZN => n3260);
   U19471 : NAND2_X2 port map( A1 => n26404, A2 => n15019, ZN => n23087);
   U19475 : NAND2_X2 port map( A1 => n15831, A2 => n32002, ZN => n17334);
   U19481 : NAND2_X2 port map( A1 => n31264, A2 => n11954, ZN => n12548);
   U19484 : NAND2_X2 port map( A1 => n23998, A2 => n23997, ZN => n14490);
   U19486 : NAND3_X2 port map( A1 => n14047, A2 => n23914, A3 => n26221, ZN => 
                           n23998);
   U19488 : XOR2_X1 port map( A1 => n16060, A2 => n3682, Z => n33217);
   U19489 : NAND3_X1 port map( A1 => n11710, A2 => n13693, A3 => n28390, ZN => 
                           n33218);
   U19493 : BUF_X2 port map( I => n16331, Z => n33219);
   U19494 : XOR2_X1 port map( A1 => n11124, A2 => n33220, Z => n11175);
   U19498 : XOR2_X1 port map( A1 => n30671, A2 => n11126, Z => n33220);
   U19505 : XOR2_X1 port map( A1 => n23324, A2 => n3322, Z => n23041);
   U19506 : NAND2_X1 port map( A1 => n25430, A2 => n25444, ZN => n31141);
   U19507 : NOR2_X1 port map( A1 => n8219, A2 => n3339, ZN => n3732);
   U19511 : XOR2_X1 port map( A1 => n24689, A2 => n27153, Z => n24758);
   U19516 : NAND2_X2 port map( A1 => n2691, A2 => n31553, ZN => n24689);
   U19519 : INV_X4 port map( I => n10899, ZN => n13349);
   U19524 : XOR2_X1 port map( A1 => n12557, A2 => n33673, Z => n14798);
   U19532 : INV_X1 port map( I => n1892, ZN => n33223);
   U19534 : XOR2_X1 port map( A1 => n22104, A2 => n28612, Z => n6466);
   U19537 : NOR2_X2 port map( A1 => n33226, A2 => n31396, ZN => n33284);
   U19541 : NAND2_X1 port map( A1 => n22500, A2 => n33227, ZN => n26762);
   U19544 : XOR2_X1 port map( A1 => n27792, A2 => n5126, Z => n30333);
   U19552 : OAI21_X1 port map( A1 => n16430, A2 => n3759, B => n11888, ZN => 
                           n34075);
   U19554 : XOR2_X1 port map( A1 => n33233, A2 => n33975, Z => n22367);
   U19556 : XOR2_X1 port map( A1 => n12370, A2 => n22301, Z => n33233);
   U19563 : NAND3_X1 port map( A1 => n33962, A2 => n736, A3 => n33961, ZN => 
                           n25336);
   U19567 : NAND2_X1 port map( A1 => n4983, A2 => n2486, ZN => n33379);
   U19569 : NAND2_X2 port map( A1 => n8178, A2 => n1931, ZN => n24263);
   U19571 : NAND2_X1 port map( A1 => n24254, A2 => n2558, ZN => n24255);
   U19573 : NAND2_X2 port map( A1 => n16957, A2 => n25334, ZN => n13698);
   U19582 : NAND2_X1 port map( A1 => n17028, A2 => n66, ZN => n28531);
   U19583 : NAND2_X2 port map( A1 => n16041, A2 => n72, ZN => n25316);
   U19585 : XOR2_X1 port map( A1 => n2345, A2 => n17048, Z => n33235);
   U19586 : XOR2_X1 port map( A1 => n23310, A2 => n13888, Z => n33236);
   U19590 : OR2_X1 port map( A1 => n29494, A2 => n26098, Z => n33238);
   U19593 : NAND2_X1 port map( A1 => n31052, A2 => n7003, ZN => n2636);
   U19601 : NOR2_X2 port map( A1 => n6364, A2 => n6365, ZN => n33239);
   U19602 : AOI22_X2 port map( A1 => n19944, A2 => n2694, B1 => n17882, B2 => 
                           n16681, ZN => n33241);
   U19603 : NAND3_X2 port map( A1 => n22920, A2 => n12887, A3 => n22924, ZN => 
                           n9963);
   U19605 : NAND2_X2 port map( A1 => n29507, A2 => n12888, ZN => n22920);
   U19606 : AOI22_X2 port map( A1 => n22880, A2 => n33344, B1 => n32092, B2 => 
                           n8365, ZN => n9791);
   U19608 : AND2_X1 port map( A1 => n14335, A2 => n13147, Z => n3288);
   U19618 : NOR2_X2 port map( A1 => n33611, A2 => n29875, ZN => n33243);
   U19621 : OAI21_X2 port map( A1 => n5679, A2 => n5954, B => n33244, ZN => 
                           n4151);
   U19622 : XOR2_X1 port map( A1 => n33892, A2 => n600, Z => n6627);
   U19629 : NOR3_X1 port map( A1 => n23841, A2 => n23840, A3 => n17234, ZN => 
                           n31083);
   U19630 : INV_X2 port map( I => n33246, ZN => n34156);
   U19634 : XOR2_X1 port map( A1 => n5321, A2 => n30427, Z => n33246);
   U19635 : INV_X2 port map( I => n33247, ZN => n23767);
   U19636 : XOR2_X1 port map( A1 => n10347, A2 => n12331, Z => n33247);
   U19637 : XOR2_X1 port map( A1 => n13496, A2 => n15438, Z => n10200);
   U19638 : NAND3_X2 port map( A1 => n17036, A2 => n19931, A3 => n17035, ZN => 
                           n16515);
   U19643 : XOR2_X1 port map( A1 => n7078, A2 => n27922, Z => n26812);
   U19644 : XOR2_X1 port map( A1 => n23291, A2 => n5512, Z => n5511);
   U19645 : OAI22_X2 port map( A1 => n27835, A2 => n27834, B1 => n22614, B2 => 
                           n22813, ZN => n23291);
   U19648 : OAI21_X2 port map( A1 => n2722, A2 => n5289, B => n2721, ZN => 
                           n33766);
   U19649 : XOR2_X1 port map( A1 => n33248, A2 => n25457, Z => Ciphertext(107))
                           ;
   U19650 : NAND2_X2 port map( A1 => n29920, A2 => n33249, ZN => n26881);
   U19651 : XOR2_X1 port map( A1 => n22100, A2 => n22121, Z => n17586);
   U19653 : NAND2_X2 port map( A1 => n21725, A2 => n21724, ZN => n22100);
   U19654 : XOR2_X1 port map( A1 => n17797, A2 => n33250, Z => n23944);
   U19659 : XOR2_X1 port map( A1 => n33895, A2 => n23316, Z => n33250);
   U19669 : NAND2_X2 port map( A1 => n33251, A2 => n6311, ZN => n17423);
   U19683 : AOI22_X2 port map( A1 => n8242, A2 => n9014, B1 => n20629, B2 => 
                           n9255, ZN => n33251);
   U19693 : NAND2_X2 port map( A1 => n13196, A2 => n23953, ZN => n4823);
   U19695 : XOR2_X1 port map( A1 => n33253, A2 => n33252, Z => n33269);
   U19698 : NAND2_X2 port map( A1 => n25490, A2 => n25473, ZN => n25464);
   U19700 : NOR2_X2 port map( A1 => n84, A2 => n24672, ZN => n25490);
   U19703 : AOI21_X1 port map( A1 => n29748, A2 => n24052, B => n24182, ZN => 
                           n18179);
   U19712 : OAI21_X2 port map( A1 => n33255, A2 => n33254, B => n18889, ZN => 
                           n11302);
   U19713 : NOR2_X2 port map( A1 => n18886, A2 => n18887, ZN => n33254);
   U19714 : NOR2_X2 port map( A1 => n13349, A2 => n4993, ZN => n15555);
   U19722 : INV_X2 port map( I => n33256, ZN => n9630);
   U19723 : XOR2_X1 port map( A1 => n4395, A2 => n22292, Z => n33256);
   U19731 : OAI21_X1 port map( A1 => n33257, A2 => n28246, B => n16957, ZN => 
                           n30025);
   U19732 : INV_X1 port map( I => n16850, ZN => n33257);
   U19739 : OAI21_X2 port map( A1 => n26038, A2 => n419, B => n28279, ZN => 
                           n33258);
   U19741 : XOR2_X1 port map( A1 => n23361, A2 => n23362, Z => n23366);
   U19742 : XOR2_X1 port map( A1 => n23328, A2 => n7070, Z => n23362);
   U19744 : NOR2_X2 port map( A1 => n29328, A2 => n31531, ZN => n2130);
   U19748 : OAI22_X2 port map( A1 => n26422, A2 => n3999, B1 => n23002, B2 => 
                           n13159, ZN => n23004);
   U19764 : XOR2_X1 port map( A1 => n33259, A2 => n29108, Z => n2108);
   U19769 : XOR2_X1 port map( A1 => n33860, A2 => n24593, Z => n33259);
   U19770 : OAI21_X2 port map( A1 => n32011, A2 => n33261, B => n17606, ZN => 
                           n28674);
   U19771 : OAI22_X2 port map( A1 => n1595, A2 => n21692, B1 => n21691, B2 => 
                           n2708, ZN => n22113);
   U19777 : INV_X2 port map( I => n24031, ZN => n1241);
   U19778 : OAI21_X2 port map( A1 => n7384, A2 => n7383, B => n6308, ZN => 
                           n24031);
   U19780 : OAI22_X2 port map( A1 => n34080, A2 => n17975, B1 => n19841, B2 => 
                           n10057, ZN => n2198);
   U19782 : NOR2_X1 port map( A1 => n28037, A2 => n33263, ZN => n5858);
   U19786 : NAND2_X1 port map( A1 => n32111, A2 => n26974, ZN => n1734);
   U19787 : XOR2_X1 port map( A1 => n24620, A2 => n12800, Z => n24489);
   U19796 : NAND2_X2 port map( A1 => n10777, A2 => n15570, ZN => n24620);
   U19797 : XOR2_X1 port map( A1 => n23291, A2 => n5212, Z => n23403);
   U19798 : NAND2_X2 port map( A1 => n9243, A2 => n9244, ZN => n5212);
   U19802 : NOR2_X2 port map( A1 => n31930, A2 => n18079, ZN => n11659);
   U19804 : BUF_X2 port map( I => n15710, Z => n33265);
   U19806 : OAI21_X2 port map( A1 => n18970, A2 => n18600, B => n33266, ZN => 
                           n28806);
   U19812 : AOI22_X2 port map( A1 => n6639, A2 => n19156, B1 => n6637, B2 => 
                           n6638, ZN => n33266);
   U19814 : NAND2_X2 port map( A1 => n5343, A2 => n17873, ZN => n15114);
   U19822 : XOR2_X1 port map( A1 => n22779, A2 => n23400, Z => n33267);
   U19829 : XOR2_X1 port map( A1 => n11514, A2 => n33268, Z => n30570);
   U19836 : XOR2_X1 port map( A1 => n30792, A2 => n1741, Z => n33268);
   U19839 : INV_X2 port map( I => n33269, ZN => n17157);
   U19840 : XOR2_X1 port map( A1 => n3395, A2 => n27601, Z => n2953);
   U19842 : NAND2_X2 port map( A1 => n11904, A2 => n17661, ZN => n17374);
   U19843 : XOR2_X1 port map( A1 => n1923, A2 => n29167, Z => n20870);
   U19844 : XOR2_X1 port map( A1 => n5148, A2 => n101, Z => n17380);
   U19846 : XOR2_X1 port map( A1 => n5150, A2 => n29130, Z => n5148);
   U19847 : INV_X2 port map( I => n33270, ZN => n34157);
   U19850 : XOR2_X1 port map( A1 => n14887, A2 => n17643, Z => n33270);
   U19851 : XOR2_X1 port map( A1 => n10780, A2 => n19486, Z => n12145);
   U19854 : XOR2_X1 port map( A1 => n26778, A2 => n11691, Z => n20772);
   U19861 : AOI22_X2 port map( A1 => n26466, A2 => n7041, B1 => n7064, B2 => 
                           n25704, ZN => n9496);
   U19863 : NAND2_X2 port map( A1 => n29503, A2 => n10733, ZN => n28429);
   U19864 : NOR2_X2 port map( A1 => n33272, A2 => n33271, ZN => n26814);
   U19871 : NOR2_X2 port map( A1 => n5825, A2 => n2288, ZN => n33272);
   U19873 : NOR2_X2 port map( A1 => n15150, A2 => n33273, ZN => n24909);
   U19876 : AOI21_X2 port map( A1 => n24362, A2 => n11945, B => n33053, ZN => 
                           n33273);
   U19877 : OR2_X1 port map( A1 => n12290, A2 => n14926, Z => n28383);
   U19879 : INV_X1 port map( I => n4790, ZN => n33274);
   U19881 : XOR2_X1 port map( A1 => n23388, A2 => n23499, Z => n4790);
   U19893 : XOR2_X1 port map( A1 => n17235, A2 => n33275, Z => n23886);
   U19896 : XOR2_X1 port map( A1 => n23460, A2 => n643, Z => n33275);
   U19897 : XOR2_X1 port map( A1 => n23469, A2 => n33276, Z => n28031);
   U19898 : XOR2_X1 port map( A1 => n31354, A2 => n23388, Z => n33276);
   U19904 : NAND2_X1 port map( A1 => n24974, A2 => n33278, ZN => n33277);
   U19911 : INV_X2 port map( I => n24610, ZN => n33278);
   U19915 : XOR2_X1 port map( A1 => n24692, A2 => n29639, Z => n29638);
   U19919 : XOR2_X1 port map( A1 => n24533, A2 => n16141, Z => n24692);
   U19922 : INV_X2 port map( I => n33279, ZN => n7993);
   U19925 : XNOR2_X1 port map( A1 => n5158, A2 => n5159, ZN => n33279);
   U19927 : NAND2_X2 port map( A1 => n33284, A2 => n5258, ZN => n1808);
   U19934 : NAND2_X2 port map( A1 => n21996, A2 => n8269, ZN => n33285);
   U19935 : NAND3_X2 port map( A1 => n22512, A2 => n22513, A3 => n22600, ZN => 
                           n14044);
   U19937 : NAND2_X2 port map( A1 => n6837, A2 => n33287, ZN => n31894);
   U19941 : NAND4_X2 port map( A1 => n22569, A2 => n7053, A3 => n22443, A4 => 
                           n22442, ZN => n33287);
   U19944 : NOR2_X1 port map( A1 => n9059, A2 => n7753, ZN => n9058);
   U19950 : OAI22_X2 port map( A1 => n21445, A2 => n6277, B1 => n21101, B2 => 
                           n16526, ZN => n26622);
   U19954 : XOR2_X1 port map( A1 => n23478, A2 => n12714, Z => n27866);
   U19956 : XOR2_X1 port map( A1 => n22157, A2 => n30275, Z => n7911);
   U19958 : NAND2_X2 port map( A1 => n115, A2 => n34084, ZN => n30275);
   U19966 : NAND2_X1 port map( A1 => n12006, A2 => n32901, ZN => n18695);
   U19970 : XOR2_X1 port map( A1 => n7045, A2 => n15183, Z => n23145);
   U19971 : INV_X2 port map( I => n33289, ZN => n26712);
   U19981 : XNOR2_X1 port map( A1 => n13294, A2 => n13293, ZN => n33289);
   U19990 : XOR2_X1 port map( A1 => n6090, A2 => n33290, Z => n31411);
   U19991 : XOR2_X1 port map( A1 => n31499, A2 => n33823, Z => n33290);
   U19996 : NAND2_X2 port map( A1 => n7817, A2 => n135, ZN => n22832);
   U20001 : AOI22_X2 port map( A1 => n7169, A2 => n10498, B1 => n17580, B2 => 
                           n23885, ZN => n24248);
   U20007 : XOR2_X1 port map( A1 => n21891, A2 => n22256, Z => n33291);
   U20010 : XOR2_X1 port map( A1 => n5925, A2 => n19727, Z => n29486);
   U20011 : XOR2_X1 port map( A1 => n19386, A2 => n19403, Z => n19727);
   U20019 : INV_X2 port map( I => n33292, ZN => n4378);
   U20023 : XOR2_X1 port map( A1 => n4379, A2 => n4380, Z => n33292);
   U20024 : XOR2_X1 port map( A1 => n12785, A2 => n16662, Z => n14237);
   U20025 : NOR2_X2 port map( A1 => n20636, A2 => n26907, ZN => n20652);
   U20026 : AOI22_X2 port map( A1 => n33294, A2 => n6985, B1 => n13411, B2 => 
                           n13592, ZN => n3786);
   U20030 : XOR2_X1 port map( A1 => n2894, A2 => n30331, Z => n13198);
   U20037 : NAND2_X2 port map( A1 => n26261, A2 => n3469, ZN => n30331);
   U20040 : XOR2_X1 port map( A1 => n10650, A2 => n33437, Z => n22118);
   U20045 : NAND2_X2 port map( A1 => n33676, A2 => n16014, ZN => n33437);
   U20046 : BUF_X2 port map( I => n24138, Z => n33295);
   U20047 : NAND3_X2 port map( A1 => n31025, A2 => n8046, A3 => n14618, ZN => 
                           n21738);
   U20050 : INV_X2 port map( I => n33296, ZN => n26084);
   U20055 : XOR2_X1 port map( A1 => n19395, A2 => n19230, Z => n33296);
   U20061 : NAND2_X2 port map( A1 => n31583, A2 => n33297, ZN => n31473);
   U20067 : AOI21_X2 port map( A1 => n8712, A2 => n8711, B => n25633, ZN => 
                           n31830);
   U20073 : NAND2_X2 port map( A1 => n6835, A2 => n6836, ZN => n29317);
   U20076 : OAI21_X2 port map( A1 => n2986, A2 => n2987, B => n29821, ZN => 
                           n13320);
   U20089 : OR2_X1 port map( A1 => n31034, A2 => n26170, Z => n6309);
   U20100 : NAND2_X2 port map( A1 => n10832, A2 => n33299, ZN => n31325);
   U20102 : XOR2_X1 port map( A1 => n21903, A2 => n31606, Z => n33300);
   U20106 : NAND2_X2 port map( A1 => n1567, A2 => n25152, ZN => n30615);
   U20107 : NAND2_X2 port map( A1 => n13028, A2 => n21498, ZN => n13113);
   U20108 : BUF_X2 port map( I => n23807, Z => n33302);
   U20109 : AND2_X1 port map( A1 => n30282, A2 => n31915, Z => n6042);
   U20111 : XOR2_X1 port map( A1 => n33303, A2 => n3739, Z => n15372);
   U20114 : NAND2_X1 port map( A1 => n25177, A2 => n8929, ZN => n33428);
   U20115 : OAI22_X2 port map( A1 => n9404, A2 => n20165, B1 => n20164, B2 => 
                           n20476, ZN => n33373);
   U20116 : NOR2_X2 port map( A1 => n23966, A2 => n23967, ZN => n29767);
   U20122 : NOR2_X2 port map( A1 => n29834, A2 => n23771, ZN => n23966);
   U20128 : AOI22_X2 port map( A1 => n33221, A2 => n28306, B1 => n23722, B2 => 
                           n847, ZN => n33304);
   U20131 : XOR2_X1 port map( A1 => n16837, A2 => n536, Z => n6175);
   U20143 : NAND2_X2 port map( A1 => n33305, A2 => n5926, ZN => n10385);
   U20144 : NAND2_X1 port map( A1 => n9885, A2 => n15411, ZN => n13252);
   U20145 : OAI22_X2 port map( A1 => n1449, A2 => n34141, B1 => n26378, B2 => 
                           n1446, ZN => n15411);
   U20151 : NAND2_X2 port map( A1 => n33306, A2 => n22699, ZN => n23282);
   U20152 : NOR2_X2 port map( A1 => n33314, A2 => n34115, ZN => n31895);
   U20159 : INV_X2 port map( I => n14612, ZN => n12715);
   U20160 : NAND3_X2 port map( A1 => n12418, A2 => n12781, A3 => n12417, ZN => 
                           n14612);
   U20166 : NAND2_X1 port map( A1 => n33308, A2 => n7023, ZN => n11031);
   U20170 : OAI21_X1 port map( A1 => n22491, A2 => n16225, B => n27897, ZN => 
                           n33308);
   U20171 : NOR2_X1 port map( A1 => n29098, A2 => n29099, ZN => n33569);
   U20172 : XOR2_X1 port map( A1 => n28822, A2 => n29042, Z => n20443);
   U20175 : INV_X2 port map( I => n11097, ZN => n33310);
   U20176 : INV_X1 port map( I => n1018, ZN => n30267);
   U20194 : INV_X4 port map( I => n21780, ZN => n31220);
   U20196 : NAND2_X2 port map( A1 => n15443, A2 => n33695, ZN => n21780);
   U20202 : XOR2_X1 port map( A1 => n3847, A2 => n12765, Z => n12764);
   U20209 : BUF_X2 port map( I => n22537, Z => n33312);
   U20212 : NAND2_X2 port map( A1 => n33313, A2 => n23727, ZN => n3880);
   U20214 : NAND3_X1 port map( A1 => n7269, A2 => n7425, A3 => n7268, ZN => 
                           n33318);
   U20219 : OAI21_X1 port map( A1 => n996, A2 => n22667, B => n22580, ZN => 
                           n4994);
   U20221 : OAI21_X2 port map( A1 => n31926, A2 => n32588, B => n32499, ZN => 
                           n33315);
   U20223 : INV_X2 port map( I => n11754, ZN => n24118);
   U20224 : XOR2_X1 port map( A1 => n12980, A2 => n33316, Z => n8885);
   U20226 : XOR2_X1 port map( A1 => n1308, A2 => n21892, Z => n33316);
   U20237 : XOR2_X1 port map( A1 => n9131, A2 => n23470, Z => n33317);
   U20238 : INV_X4 port map( I => n654, ZN => n34009);
   U20242 : OAI22_X2 port map( A1 => n29342, A2 => n1124, B1 => n22542, B2 => 
                           n22397, ZN => n8991);
   U20247 : NAND2_X2 port map( A1 => n6257, A2 => n33739, ZN => n29342);
   U20248 : NAND3_X1 port map( A1 => n33318, A2 => n7265, A3 => n7266, ZN => 
                           Ciphertext(181));
   U20251 : XOR2_X1 port map( A1 => n14532, A2 => n24806, Z => n33319);
   U20252 : AOI21_X2 port map( A1 => n27947, A2 => n25630, B => n31974, ZN => 
                           n31604);
   U20253 : NAND2_X2 port map( A1 => n26585, A2 => n17497, ZN => n20495);
   U20257 : AOI22_X2 port map( A1 => n12161, A2 => n34046, B1 => n396, B2 => 
                           n29454, ZN => n33321);
   U20258 : INV_X1 port map( I => n2618, ZN => n1348);
   U20259 : NAND2_X2 port map( A1 => n9403, A2 => n33288, ZN => n2618);
   U20267 : NAND2_X2 port map( A1 => n33323, A2 => n30857, ZN => n14720);
   U20268 : NAND2_X1 port map( A1 => n29339, A2 => n29250, ZN => n29872);
   U20271 : XOR2_X1 port map( A1 => n8728, A2 => n13606, Z => n20977);
   U20281 : NAND3_X2 port map( A1 => n5734, A2 => n20408, A3 => n10290, ZN => 
                           n13606);
   U20283 : AND2_X1 port map( A1 => n33325, A2 => n15296, Z => n21531);
   U20286 : NAND2_X2 port map( A1 => n17715, A2 => n10925, ZN => n29337);
   U20287 : XOR2_X1 port map( A1 => Plaintext(10), A2 => Key(10), Z => n8213);
   U20290 : XOR2_X1 port map( A1 => n33326, A2 => n20916, Z => n52);
   U20293 : XOR2_X1 port map( A1 => n20792, A2 => n30163, Z => n33326);
   U20295 : NAND2_X2 port map( A1 => n7780, A2 => n29606, ZN => n7778);
   U20297 : OR2_X1 port map( A1 => n11820, A2 => n25531, Z => n33327);
   U20299 : OR2_X1 port map( A1 => n25724, A2 => n13640, Z => n2962);
   U20301 : NOR2_X2 port map( A1 => n11511, A2 => n14352, ZN => n25724);
   U20304 : XOR2_X1 port map( A1 => n33328, A2 => n19648, Z => n31900);
   U20305 : XOR2_X1 port map( A1 => n17129, A2 => n25993, Z => n33328);
   U20306 : NAND3_X2 port map( A1 => n33302, A2 => n23850, A3 => n3241, ZN => 
                           n33457);
   U20310 : INV_X2 port map( I => n33329, ZN => n758);
   U20317 : NAND2_X2 port map( A1 => n22810, A2 => n12729, ZN => n22694);
   U20324 : NAND2_X2 port map( A1 => n13972, A2 => n22424, ZN => n22810);
   U20326 : OAI21_X2 port map( A1 => n10747, A2 => n25233, B => n11132, ZN => 
                           n33330);
   U20327 : XOR2_X1 port map( A1 => n1707, A2 => n33331, Z => n15865);
   U20328 : AND2_X1 port map( A1 => n6118, A2 => n9766, Z => n7726);
   U20329 : NAND2_X2 port map( A1 => n16920, A2 => n16918, ZN => n23355);
   U20333 : AOI22_X2 port map( A1 => n30243, A2 => n29286, B1 => n15747, B2 => 
                           n21514, ZN => n10233);
   U20336 : AOI21_X2 port map( A1 => n23006, A2 => n3999, B => n23004, ZN => 
                           n7070);
   U20338 : XOR2_X1 port map( A1 => n20987, A2 => n33332, Z => n3298);
   U20342 : OAI22_X2 port map( A1 => n14996, A2 => n14997, B1 => n14999, B2 => 
                           n14998, ZN => n21761);
   U20348 : XOR2_X1 port map( A1 => n32516, A2 => n29155, Z => n33333);
   U20349 : XOR2_X1 port map( A1 => n9464, A2 => n33334, Z => n30214);
   U20350 : XOR2_X1 port map( A1 => n26715, A2 => n28295, Z => n33334);
   U20352 : BUF_X2 port map( I => n30781, Z => n33335);
   U20355 : NAND2_X2 port map( A1 => n1816, A2 => n1819, ZN => n24220);
   U20371 : NAND2_X2 port map( A1 => n30354, A2 => n14463, ZN => n1816);
   U20374 : NAND2_X2 port map( A1 => n33336, A2 => n27270, ZN => n3266);
   U20377 : XOR2_X1 port map( A1 => n5600, A2 => n22027, Z => n33338);
   U20381 : XOR2_X1 port map( A1 => n9904, A2 => n11102, Z => n33339);
   U20383 : NAND2_X2 port map( A1 => n11492, A2 => n11491, ZN => n30651);
   U20384 : XOR2_X1 port map( A1 => n15889, A2 => n15891, Z => n14029);
   U20387 : XOR2_X1 port map( A1 => n20848, A2 => n20729, Z => n5724);
   U20388 : NAND2_X2 port map( A1 => n26212, A2 => n29672, ZN => n20848);
   U20389 : XOR2_X1 port map( A1 => n5979, A2 => n3957, Z => n9203);
   U20401 : NAND2_X2 port map( A1 => n3440, A2 => n3439, ZN => n13357);
   U20403 : NOR3_X2 port map( A1 => n28276, A2 => n26969, A3 => n1180, ZN => 
                           n31246);
   U20408 : OR2_X1 port map( A1 => n3468, A2 => n8784, Z => n26265);
   U20414 : NAND2_X2 port map( A1 => n4878, A2 => n18897, ZN => n29030);
   U20419 : NAND3_X2 port map( A1 => n4611, A2 => n33686, A3 => n17774, ZN => 
                           n15183);
   U20420 : NAND2_X1 port map( A1 => n7751, A2 => n33069, ZN => n8193);
   U20421 : NAND2_X2 port map( A1 => n33342, A2 => n28888, ZN => n3994);
   U20424 : NOR2_X2 port map( A1 => n9016, A2 => n9017, ZN => n33342);
   U20426 : NAND3_X1 port map( A1 => n24924, A2 => n30328, A3 => n24925, ZN => 
                           n33343);
   U20428 : XOR2_X1 port map( A1 => n10196, A2 => n10194, Z => n18220);
   U20429 : XOR2_X1 port map( A1 => n22015, A2 => n4342, Z => n12614);
   U20430 : NAND3_X1 port map( A1 => n25449, A2 => n33658, A3 => n25447, ZN => 
                           n33469);
   U20436 : NAND2_X2 port map( A1 => n23864, A2 => n10993, ZN => n23930);
   U20438 : XOR2_X1 port map( A1 => n2917, A2 => n2918, Z => n29288);
   U20439 : NOR2_X1 port map( A1 => n25818, A2 => n25804, ZN => n25811);
   U20448 : NAND2_X2 port map( A1 => n11185, A2 => n12420, ZN => n25804);
   U20450 : NAND3_X2 port map( A1 => n22620, A2 => n33347, A3 => n33346, ZN => 
                           n16073);
   U20462 : NAND2_X2 port map( A1 => n33349, A2 => n31403, ZN => n25863);
   U20463 : AOI21_X1 port map( A1 => n21503, A2 => n13028, B => n30346, ZN => 
                           n21504);
   U20465 : NAND2_X2 port map( A1 => n2570, A2 => n30403, ZN => n34046);
   U20469 : XOR2_X1 port map( A1 => n24801, A2 => n7603, Z => n24567);
   U20471 : AOI21_X2 port map( A1 => n4786, A2 => n11732, B => n33350, ZN => 
                           n4785);
   U20486 : XOR2_X1 port map( A1 => n19728, A2 => n12223, Z => n17193);
   U20487 : XOR2_X1 port map( A1 => n19625, A2 => n19530, Z => n12223);
   U20499 : XOR2_X1 port map( A1 => n24388, A2 => n29140, Z => n4418);
   U20500 : NAND3_X2 port map( A1 => n12605, A2 => n12604, A3 => n5384, ZN => 
                           n9536);
   U20502 : NOR2_X1 port map( A1 => n34009, A2 => n32308, ZN => n8849);
   U20504 : NAND2_X2 port map( A1 => n8848, A2 => n8851, ZN => n24159);
   U20506 : XOR2_X1 port map( A1 => n17153, A2 => n8109, Z => n33351);
   U20514 : XNOR2_X1 port map( A1 => n16897, A2 => n21888, ZN => n33975);
   U20516 : NAND2_X2 port map( A1 => n1579, A2 => n1580, ZN => n22960);
   U20517 : NAND2_X1 port map( A1 => n28722, A2 => n7083, ZN => n28990);
   U20518 : NAND2_X1 port map( A1 => n25657, A2 => n25665, ZN => n28722);
   U20519 : INV_X2 port map( I => n29042, ZN => n30163);
   U20522 : NAND2_X2 port map( A1 => n2620, A2 => n11412, ZN => n29042);
   U20525 : INV_X2 port map( I => n24779, ZN => n14627);
   U20530 : NAND2_X1 port map( A1 => n13650, A2 => n13649, ZN => n2293);
   U20531 : INV_X2 port map( I => n23385, ZN => n26426);
   U20537 : NAND2_X2 port map( A1 => n14466, A2 => n14465, ZN => n23385);
   U20540 : INV_X2 port map( I => n33354, ZN => n10193);
   U20541 : XOR2_X1 port map( A1 => n7191, A2 => n33355, Z => n15057);
   U20545 : XOR2_X1 port map( A1 => n7193, A2 => n15157, Z => n33355);
   U20546 : OAI22_X2 port map( A1 => n33357, A2 => n33356, B1 => n13325, B2 => 
                           n26343, ZN => n13696);
   U20547 : INV_X1 port map( I => n6475, ZN => n33356);
   U20554 : XOR2_X1 port map( A1 => n21027, A2 => n13338, Z => n33358);
   U20559 : XOR2_X1 port map( A1 => n24505, A2 => n6897, Z => n33359);
   U20564 : AOI22_X2 port map( A1 => n11705, A2 => n11704, B1 => n9548, B2 => 
                           n11703, ZN => n16509);
   U20567 : NAND2_X2 port map( A1 => n21087, A2 => n21209, ZN => n21382);
   U20571 : OR2_X1 port map( A1 => n18064, A2 => n12895, Z => n9661);
   U20573 : NAND2_X2 port map( A1 => n19910, A2 => n17633, ZN => n20960);
   U20577 : NAND2_X1 port map( A1 => n4066, A2 => n19158, ZN => n13059);
   U20578 : NAND3_X1 port map( A1 => n7968, A2 => n25999, A3 => n8233, ZN => 
                           n19130);
   U20579 : NAND2_X1 port map( A1 => n33360, A2 => n15456, ZN => n26705);
   U20582 : NAND2_X2 port map( A1 => n16134, A2 => n16133, ZN => n14485);
   U20584 : XOR2_X1 port map( A1 => n33361, A2 => n25929, Z => Ciphertext(191))
                           ;
   U20586 : OAI22_X1 port map( A1 => n25927, A2 => n25926, B1 => n25924, B2 => 
                           n25925, ZN => n33361);
   U20590 : NAND2_X2 port map( A1 => n20433, A2 => n20431, ZN => n14365);
   U20591 : XOR2_X1 port map( A1 => n33362, A2 => n14584, Z => n5692);
   U20593 : XOR2_X1 port map( A1 => n34120, A2 => n23533, Z => n33362);
   U20598 : XOR2_X1 port map( A1 => n5522, A2 => n5523, Z => n29936);
   U20605 : INV_X2 port map( I => n33363, ZN => n11784);
   U20607 : XOR2_X1 port map( A1 => n22063, A2 => n9960, Z => n33363);
   U20621 : NAND2_X2 port map( A1 => n33365, A2 => n33364, ZN => n21742);
   U20625 : NAND2_X2 port map( A1 => n33367, A2 => n33366, ZN => n33365);
   U20628 : INV_X2 port map( I => n423, ZN => n33366);
   U20633 : NAND2_X2 port map( A1 => n3854, A2 => n33368, ZN => n33869);
   U20634 : XOR2_X1 port map( A1 => n17765, A2 => n15821, Z => n17879);
   U20636 : XOR2_X1 port map( A1 => n23438, A2 => n23439, Z => n3514);
   U20637 : NAND2_X2 port map( A1 => n17460, A2 => n17458, ZN => n23438);
   U20644 : INV_X2 port map( I => n2940, ZN => n8924);
   U20648 : XOR2_X1 port map( A1 => n2926, A2 => n2924, Z => n2940);
   U20649 : XOR2_X1 port map( A1 => n22229, A2 => n22230, Z => n11282);
   U20654 : XOR2_X1 port map( A1 => n22305, A2 => n22308, Z => n22230);
   U20656 : XOR2_X1 port map( A1 => n7057, A2 => n1984, Z => n19578);
   U20658 : AOI21_X2 port map( A1 => n33555, A2 => n19003, B => n7749, ZN => 
                           n1984);
   U20663 : XOR2_X1 port map( A1 => n32478, A2 => n21028, Z => n20787);
   U20666 : INV_X2 port map( I => n29296, ZN => n30504);
   U20669 : OAI21_X2 port map( A1 => n6631, A2 => n20144, B => n6630, ZN => 
                           n29296);
   U20671 : XNOR2_X1 port map( A1 => n16303, A2 => n4028, ZN => n33427);
   U20672 : NAND2_X2 port map( A1 => n23556, A2 => n5685, ZN => n29499);
   U20674 : XOR2_X1 port map( A1 => n6348, A2 => n1708, Z => n1707);
   U20685 : XOR2_X1 port map( A1 => n20778, A2 => n31185, Z => n33369);
   U20694 : NAND2_X2 port map( A1 => n30222, A2 => n26576, ZN => n31477);
   U20696 : NAND2_X2 port map( A1 => n12315, A2 => n3614, ZN => n22762);
   U20700 : NAND2_X2 port map( A1 => n22418, A2 => n33582, ZN => n12315);
   U20701 : OAI21_X2 port map( A1 => n11714, A2 => n11715, B => n19009, ZN => 
                           n11177);
   U20706 : INV_X2 port map( I => n31511, ZN => n31007);
   U20708 : NAND2_X2 port map( A1 => n13292, A2 => n34158, ZN => n31511);
   U20717 : NOR3_X1 port map( A1 => n22634, A2 => n28979, A3 => n7513, ZN => 
                           n18012);
   U20718 : NAND2_X2 port map( A1 => n33370, A2 => n17387, ZN => n24250);
   U20725 : OR2_X2 port map( A1 => n8444, A2 => n9968, Z => n24361);
   U20728 : NAND2_X2 port map( A1 => n16639, A2 => n26712, ZN => n21326);
   U20729 : XOR2_X1 port map( A1 => n10758, A2 => n33371, Z => n17014);
   U20731 : XOR2_X1 port map( A1 => n23441, A2 => n23442, Z => n33371);
   U20734 : NAND2_X1 port map( A1 => n27594, A2 => n3016, ZN => n33372);
   U20748 : NAND3_X1 port map( A1 => n18752, A2 => n18753, A3 => n18983, ZN => 
                           n18754);
   U20753 : NAND2_X2 port map( A1 => n31850, A2 => n16288, ZN => n18752);
   U20754 : XOR2_X1 port map( A1 => n15093, A2 => n15934, Z => n27182);
   U20758 : OAI21_X2 port map( A1 => n15650, A2 => n4850, B => n30106, ZN => 
                           n30105);
   U20760 : XOR2_X1 port map( A1 => n23363, A2 => n23385, Z => n23463);
   U20762 : NAND2_X2 port map( A1 => n29266, A2 => n16635, ZN => n23363);
   U20765 : XOR2_X1 port map( A1 => n33374, A2 => n19371, Z => n19439);
   U20766 : INV_X2 port map( I => n19599, ZN => n33374);
   U20769 : NAND2_X2 port map( A1 => n7440, A2 => n7439, ZN => n19371);
   U20770 : XOR2_X1 port map( A1 => n33375, A2 => n24787, Z => n8152);
   U20771 : NAND2_X2 port map( A1 => n14309, A2 => n5115, ZN => n24995);
   U20776 : XOR2_X1 port map( A1 => n33377, A2 => n33376, Z => n26284);
   U20780 : XOR2_X1 port map( A1 => n9346, A2 => n31252, Z => n33377);
   U20784 : NAND2_X2 port map( A1 => n33832, A2 => n7581, ZN => n24091);
   U20795 : XOR2_X1 port map( A1 => n33378, A2 => n29447, Z => n11248);
   U20801 : XOR2_X1 port map( A1 => n19493, A2 => n34071, Z => n33378);
   U20803 : INV_X1 port map( I => n25891, ZN => n33474);
   U20807 : OAI21_X2 port map( A1 => n10556, A2 => n16795, B => n20043, ZN => 
                           n17241);
   U20808 : XOR2_X1 port map( A1 => n4020, A2 => n23537, Z => n28407);
   U20809 : INV_X2 port map( I => n16310, ZN => n33687);
   U20811 : XOR2_X1 port map( A1 => n33381, A2 => n7572, Z => n1942);
   U20812 : XOR2_X1 port map( A1 => n5127, A2 => n31410, Z => n33381);
   U20813 : OAI21_X2 port map( A1 => n28543, A2 => n28544, B => n33206, ZN => 
                           n3900);
   U20819 : NOR2_X1 port map( A1 => n4180, A2 => n29908, ZN => n17714);
   U20820 : XOR2_X1 port map( A1 => n22044, A2 => n9536, Z => n8630);
   U20822 : NAND2_X2 port map( A1 => n33384, A2 => n24613, ZN => n8622);
   U20829 : OAI21_X2 port map( A1 => n15231, A2 => n28815, B => n15232, ZN => 
                           n33384);
   U20837 : NAND2_X2 port map( A1 => n33738, A2 => n33385, ZN => n14002);
   U20841 : BUF_X2 port map( I => n13684, Z => n33386);
   U20842 : AND2_X1 port map( A1 => n25711, A2 => n4449, Z => n13924);
   U20845 : NAND2_X2 port map( A1 => n30044, A2 => n14856, ZN => n14201);
   U20846 : AOI21_X1 port map( A1 => n3717, A2 => n15522, B => n12323, ZN => 
                           n21058);
   U20848 : AOI22_X2 port map( A1 => n13026, A2 => n17599, B1 => n13025, B2 => 
                           n13024, ZN => n19274);
   U20849 : NAND2_X2 port map( A1 => n28484, A2 => n28829, ZN => n20990);
   U20856 : XNOR2_X1 port map( A1 => n19389, A2 => n31882, ZN => n26300);
   U20857 : OAI21_X1 port map( A1 => n29432, A2 => n17964, B => n742, ZN => 
                           n15168);
   U20859 : NOR2_X2 port map( A1 => n33390, A2 => n26874, ZN => n16321);
   U20862 : INV_X2 port map( I => n33391, ZN => n26641);
   U20864 : NAND2_X2 port map( A1 => n25332, A2 => n16783, ZN => n15624);
   U20866 : NAND2_X2 port map( A1 => n33394, A2 => n33393, ZN => n25332);
   U20873 : INV_X2 port map( I => n28093, ZN => n33393);
   U20876 : NAND2_X2 port map( A1 => n31886, A2 => n31572, ZN => n34116);
   U20891 : OR2_X1 port map( A1 => n26345, A2 => n4755, Z => n12441);
   U20893 : OAI21_X2 port map( A1 => n327, A2 => n17473, B => n22443, ZN => 
                           n13127);
   U20894 : NAND2_X2 port map( A1 => n327, A2 => n27959, ZN => n22443);
   U20896 : NOR2_X2 port map( A1 => n11235, A2 => n22748, ZN => n17707);
   U20905 : AOI22_X2 port map( A1 => n33398, A2 => n33397, B1 => n7290, B2 => 
                           n15217, ZN => n13547);
   U20910 : XOR2_X1 port map( A1 => n33401, A2 => n16674, Z => Ciphertext(118))
                           ;
   U20911 : XOR2_X1 port map( A1 => n2854, A2 => n7832, Z => n2857);
   U20912 : NAND2_X2 port map( A1 => n6945, A2 => n33402, ZN => n22945);
   U20914 : NAND2_X1 port map( A1 => n9991, A2 => n10754, ZN => n9990);
   U20916 : XOR2_X1 port map( A1 => n14588, A2 => n1464, Z => n9006);
   U20921 : NAND2_X2 port map( A1 => n29581, A2 => n29580, ZN => n1464);
   U20923 : AND3_X1 port map( A1 => n20109, A2 => n33848, A3 => n8421, Z => 
                           n2906);
   U20933 : BUF_X2 port map( I => n21755, Z => n33403);
   U20935 : XOR2_X1 port map( A1 => n31495, A2 => n33404, Z => n31453);
   U20949 : XOR2_X1 port map( A1 => n19541, A2 => n19471, Z => n33404);
   U20954 : NOR2_X2 port map( A1 => n33405, A2 => n13610, ZN => n20545);
   U20955 : OAI21_X2 port map( A1 => n11414, A2 => n33419, B => n5470, ZN => 
                           n13610);
   U20956 : INV_X1 port map( I => n33406, ZN => n33405);
   U20957 : NAND2_X1 port map( A1 => n13611, A2 => n12078, ZN => n33406);
   U20959 : NOR2_X2 port map( A1 => n14649, A2 => n26890, ZN => n33407);
   U20961 : XOR2_X1 port map( A1 => n23337, A2 => n23146, Z => n2842);
   U20962 : XOR2_X1 port map( A1 => n17775, A2 => n14077, Z => n23337);
   U20965 : XOR2_X1 port map( A1 => n1607, A2 => n30407, Z => n33408);
   U20968 : XOR2_X1 port map( A1 => n4728, A2 => n24839, Z => n31340);
   U20980 : NAND2_X2 port map( A1 => n3234, A2 => n28522, ZN => n24839);
   U20982 : OAI22_X2 port map( A1 => n21666, A2 => n1134, B1 => n31089, B2 => 
                           n1136, ZN => n33409);
   U20983 : OAI21_X2 port map( A1 => n33411, A2 => n33410, B => n983, ZN => 
                           n22768);
   U20984 : NOR2_X1 port map( A1 => n33818, A2 => n641, ZN => n33410);
   U20985 : INV_X1 port map( I => n6227, ZN => n33411);
   U20988 : NOR2_X2 port map( A1 => n24001, A2 => n24000, ZN => n3220);
   U20990 : NAND3_X2 port map( A1 => n15957, A2 => n18632, A3 => n33412, ZN => 
                           n30781);
   U20991 : NAND2_X2 port map( A1 => n33413, A2 => n33650, ZN => n28736);
   U20992 : OR2_X1 port map( A1 => n22491, A2 => n630, Z => n21902);
   U20994 : INV_X2 port map( I => n33415, ZN => n18496);
   U20998 : NOR2_X2 port map( A1 => n17223, A2 => n17255, ZN => n33415);
   U21000 : NOR3_X2 port map( A1 => n5549, A2 => n5550, A3 => n33416, ZN => 
                           n5548);
   U21003 : NOR3_X2 port map( A1 => n30554, A2 => n19926, A3 => n4587, ZN => 
                           n33416);
   U21007 : XOR2_X1 port map( A1 => n14662, A2 => n8343, Z => n28027);
   U21011 : AND2_X1 port map( A1 => n386, A2 => n23745, Z => n30895);
   U21012 : XOR2_X1 port map( A1 => n2335, A2 => n28039, Z => n13510);
   U21016 : OAI22_X2 port map( A1 => n11538, A2 => n11539, B1 => n30875, B2 => 
                           n11540, ZN => n23456);
   U21020 : XOR2_X1 port map( A1 => n10758, A2 => n9671, Z => n9670);
   U21023 : XOR2_X1 port map( A1 => n23229, A2 => n26108, Z => n28286);
   U21024 : XOR2_X1 port map( A1 => n23419, A2 => n646, Z => n23229);
   U21028 : NAND2_X2 port map( A1 => n27272, A2 => n11752, ZN => n18084);
   U21035 : INV_X4 port map( I => n33420, ZN => n3944);
   U21036 : NOR2_X2 port map( A1 => n3946, A2 => n3945, ZN => n33420);
   U21043 : AND2_X1 port map( A1 => n20375, A2 => n20374, Z => n12225);
   U21053 : NAND2_X2 port map( A1 => n30996, A2 => n2492, ZN => n20375);
   U21055 : NAND2_X2 port map( A1 => n33423, A2 => n27711, ZN => n10732);
   U21059 : XOR2_X1 port map( A1 => n20862, A2 => n16831, Z => n21049);
   U21060 : NOR2_X2 port map( A1 => n29993, A2 => n4061, ZN => n20862);
   U21062 : XOR2_X1 port map( A1 => n31200, A2 => n33424, Z => n8694);
   U21064 : XOR2_X1 port map( A1 => n16382, A2 => n23342, Z => n33424);
   U21071 : INV_X1 port map( I => n33446, ZN => n23851);
   U21072 : AND2_X1 port map( A1 => n33446, A2 => n663, Z => n5817);
   U21078 : NAND2_X2 port map( A1 => n11385, A2 => n4760, ZN => n2611);
   U21080 : XOR2_X1 port map( A1 => n30535, A2 => n33426, Z => n33803);
   U21082 : XOR2_X1 port map( A1 => n23359, A2 => n32015, Z => n33426);
   U21086 : XOR2_X1 port map( A1 => n17307, A2 => n17308, Z => n6434);
   U21087 : XOR2_X1 port map( A1 => n12454, A2 => n12414, Z => n24838);
   U21094 : XNOR2_X1 port map( A1 => n7016, A2 => n21010, ZN => n33521);
   U21105 : INV_X2 port map( I => n33429, ZN => n34153);
   U21107 : XOR2_X1 port map( A1 => n3070, A2 => n3074, Z => n33429);
   U21111 : XOR2_X1 port map( A1 => n8637, A2 => n2072, Z => n31395);
   U21113 : INV_X2 port map( I => n33430, ZN => n29252);
   U21121 : XOR2_X1 port map( A1 => n19407, A2 => n8383, Z => n33430);
   U21124 : NAND2_X2 port map( A1 => n31970, A2 => n7197, ZN => n11072);
   U21126 : NAND2_X1 port map( A1 => n3979, A2 => n7502, ZN => n33954);
   U21127 : OAI21_X2 port map( A1 => n10757, A2 => n1124, B => n10288, ZN => 
                           n33433);
   U21132 : NOR2_X2 port map( A1 => n26474, A2 => n17431, ZN => n17428);
   U21133 : NAND2_X2 port map( A1 => n27016, A2 => n33435, ZN => n16278);
   U21137 : AOI22_X2 port map( A1 => n7115, A2 => n21427, B1 => n21072, B2 => 
                           n21341, ZN => n33435);
   U21140 : AOI21_X2 port map( A1 => n20598, A2 => n5993, B => n31401, ZN => 
                           n20913);
   U21142 : XOR2_X1 port map( A1 => n10026, A2 => n19627, Z => n19723);
   U21144 : NAND2_X1 port map( A1 => n33436, A2 => n8171, ZN => n27585);
   U21145 : NOR2_X1 port map( A1 => n27806, A2 => n20578, ZN => n33436);
   U21149 : NOR2_X2 port map( A1 => n10227, A2 => n764, ZN => n18907);
   U21150 : NAND2_X1 port map( A1 => n33586, A2 => n8957, ZN => n8955);
   U21156 : OAI21_X2 port map( A1 => n23112, A2 => n17099, B => n33438, ZN => 
                           n9041);
   U21166 : NAND3_X1 port map( A1 => n6453, A2 => n23109, A3 => n16022, ZN => 
                           n33438);
   U21168 : INV_X2 port map( I => n28702, ZN => n4274);
   U21173 : XOR2_X1 port map( A1 => n5138, A2 => n5137, Z => n5188);
   U21176 : XOR2_X1 port map( A1 => n2808, A2 => n33715, Z => n17245);
   U21180 : XNOR2_X1 port map( A1 => n23272, A2 => n23441, ZN => n13190);
   U21185 : NAND2_X2 port map( A1 => n4174, A2 => n5233, ZN => n23272);
   U21186 : NAND2_X1 port map( A1 => n7973, A2 => n33440, ZN => n387);
   U21192 : AOI21_X1 port map( A1 => n16397, A2 => n837, B => n13763, ZN => 
                           n33440);
   U21197 : INV_X2 port map( I => n19102, ZN => n27617);
   U21199 : NAND2_X2 port map( A1 => n18923, A2 => n19101, ZN => n19102);
   U21207 : NAND2_X2 port map( A1 => n28139, A2 => n5250, ZN => n17888);
   U21208 : AND2_X1 port map( A1 => n2697, A2 => n1119, Z => n33854);
   U21210 : OR2_X1 port map( A1 => n29944, A2 => n19991, Z => n33441);
   U21213 : NOR2_X2 port map( A1 => n30833, A2 => n12213, ZN => n23007);
   U21225 : NAND2_X2 port map( A1 => n18473, A2 => n15148, ZN => n19057);
   U21226 : XOR2_X1 port map( A1 => n3599, A2 => n19513, Z => n19731);
   U21247 : NAND2_X2 port map( A1 => n18928, A2 => n18927, ZN => n19513);
   U21249 : NAND2_X1 port map( A1 => n25621, A2 => n17499, ZN => n33442);
   U21251 : INV_X1 port map( I => n31569, ZN => n33443);
   U21256 : AOI22_X2 port map( A1 => n18226, A2 => n18731, B1 => n18733, B2 => 
                           n18730, ZN => n18225);
   U21259 : NOR2_X2 port map( A1 => n957, A2 => n26155, ZN => n18226);
   U21268 : INV_X2 port map( I => n33849, ZN => n34089);
   U21270 : XOR2_X1 port map( A1 => n13122, A2 => n32067, Z => n33849);
   U21272 : NOR2_X2 port map( A1 => n33444, A2 => n24012, ZN => n31919);
   U21273 : NAND3_X2 port map( A1 => n33445, A2 => n8591, A3 => n2391, ZN => 
                           n31805);
   U21303 : NAND2_X2 port map( A1 => n940, A2 => n4233, ZN => n33445);
   U21306 : NOR2_X2 port map( A1 => n13147, A2 => n17799, ZN => n33446);
   U21307 : INV_X2 port map( I => n27894, ZN => n10899);
   U21310 : XOR2_X1 port map( A1 => n23476, A2 => n25881, Z => n30955);
   U21311 : NAND2_X2 port map( A1 => n2636, A2 => n2637, ZN => n23476);
   U21316 : XOR2_X1 port map( A1 => n19163, A2 => n19446, Z => n4052);
   U21323 : XOR2_X1 port map( A1 => n33448, A2 => n15117, Z => n19163);
   U21325 : INV_X2 port map( I => n31731, ZN => n33448);
   U21327 : XOR2_X1 port map( A1 => n27362, A2 => n11483, Z => n11548);
   U21332 : XOR2_X1 port map( A1 => n19469, A2 => n33449, Z => n10696);
   U21334 : XOR2_X1 port map( A1 => n16792, A2 => n9503, Z => n33449);
   U21345 : NAND2_X2 port map( A1 => n4635, A2 => n4638, ZN => n28011);
   U21346 : AOI22_X2 port map( A1 => n7773, A2 => n8041, B1 => n5858, B2 => 
                           n5857, ZN => n21512);
   U21347 : XOR2_X1 port map( A1 => n26865, A2 => n7380, Z => n2915);
   U21349 : XOR2_X1 port map( A1 => n24450, A2 => n24409, Z => n8691);
   U21352 : NAND2_X2 port map( A1 => n1960, A2 => n1963, ZN => n20873);
   U21353 : NOR2_X2 port map( A1 => n1926, A2 => n1805, ZN => n22280);
   U21358 : OAI22_X2 port map( A1 => n33450, A2 => n20249, B1 => n16308, B2 => 
                           n28257, ZN => n21743);
   U21364 : NOR2_X1 port map( A1 => n15172, A2 => n21581, ZN => n30652);
   U21366 : NAND2_X2 port map( A1 => n14704, A2 => n15997, ZN => n15720);
   U21367 : OAI21_X2 port map( A1 => n4435, A2 => n4434, B => n33451, ZN => 
                           n22036);
   U21377 : AOI22_X2 port map( A1 => n4432, A2 => n33242, B1 => n21697, B2 => 
                           n4433, ZN => n33451);
   U21383 : XOR2_X1 port map( A1 => n19598, A2 => n19647, Z => n15776);
   U21384 : XOR2_X1 port map( A1 => n4437, A2 => n33452, Z => n16272);
   U21389 : XOR2_X1 port map( A1 => n28441, A2 => n31754, Z => n33452);
   U21392 : BUF_X2 port map( I => n24635, Z => n33453);
   U21393 : AOI22_X2 port map( A1 => n31080, A2 => n1681, B1 => n4301, B2 => 
                           n14927, ZN => n1680);
   U21401 : OAI22_X2 port map( A1 => n33456, A2 => n33455, B1 => n9647, B2 => 
                           n16529, ZN => n4084);
   U21416 : OAI21_X1 port map( A1 => n28240, A2 => n24031, B => n24304, ZN => 
                           n24033);
   U21421 : XOR2_X1 port map( A1 => n30273, A2 => n29169, Z => n31251);
   U21423 : XOR2_X1 port map( A1 => n22005, A2 => n22067, Z => n22288);
   U21427 : NAND2_X2 port map( A1 => n2913, A2 => n24316, ZN => n33458);
   U21433 : XOR2_X1 port map( A1 => n23419, A2 => n4732, Z => n4564);
   U21435 : NAND2_X2 port map( A1 => n31434, A2 => n14769, ZN => n23419);
   U21442 : NAND2_X2 port map( A1 => n33462, A2 => n11340, ZN => n30795);
   U21444 : NOR2_X2 port map( A1 => n28391, A2 => n32094, ZN => n33462);
   U21466 : AOI22_X2 port map( A1 => n33463, A2 => n6649, B1 => n13369, B2 => 
                           n29823, ZN => n29952);
   U21467 : NOR2_X1 port map( A1 => n16290, A2 => n26061, ZN => n33464);
   U21469 : XOR2_X1 port map( A1 => n33465, A2 => n23501, Z => n33550);
   U21470 : NAND2_X2 port map( A1 => n26883, A2 => n17923, ZN => n24207);
   U21484 : XOR2_X1 port map( A1 => n24504, A2 => n24681, Z => n6898);
   U21489 : XOR2_X1 port map( A1 => n24830, A2 => n27114, Z => n24681);
   U21492 : INV_X2 port map( I => n21326, ZN => n1142);
   U21493 : XOR2_X1 port map( A1 => n9218, A2 => n20964, Z => n9217);
   U21496 : NAND2_X1 port map( A1 => n5672, A2 => n5632, ZN => n5671);
   U21498 : XOR2_X1 port map( A1 => n17745, A2 => n22046, Z => n3303);
   U21499 : OAI21_X1 port map( A1 => n2858, A2 => n5961, B => n33466, ZN => 
                           n33485);
   U21508 : INV_X2 port map( I => n22606, ZN => n33466);
   U21517 : NAND2_X2 port map( A1 => n11402, A2 => n33467, ZN => n12421);
   U21518 : OAI21_X2 port map( A1 => n12397, A2 => n19819, B => n12396, ZN => 
                           n33467);
   U21520 : AOI22_X2 port map( A1 => n22566, A2 => n13409, B1 => n22564, B2 => 
                           n16490, ZN => n22971);
   U21521 : NAND2_X2 port map( A1 => n11874, A2 => n12530, ZN => n13409);
   U21524 : NOR2_X2 port map( A1 => n28379, A2 => n19137, ZN => n28543);
   U21525 : XOR2_X1 port map( A1 => n23470, A2 => n33960, Z => n33959);
   U21538 : NAND2_X2 port map( A1 => n27701, A2 => n2803, ZN => n23470);
   U21539 : AOI22_X2 port map( A1 => n3494, A2 => n31345, B1 => n3911, B2 => 
                           n3495, ZN => n28083);
   U21547 : NOR2_X2 port map( A1 => n28378, A2 => n10612, ZN => n3911);
   U21548 : NOR2_X1 port map( A1 => n3348, A2 => n33503, ZN => n28002);
   U21550 : XOR2_X1 port map( A1 => n13802, A2 => n21898, Z => n7114);
   U21557 : OAI22_X2 port map( A1 => n12151, A2 => n28773, B1 => n12153, B2 => 
                           n33687, ZN => n27021);
   U21569 : XOR2_X1 port map( A1 => n33469, A2 => n25450, Z => Ciphertext(106))
                           ;
   U21573 : NAND2_X2 port map( A1 => n33471, A2 => n6514, ZN => n22158);
   U21574 : INV_X2 port map( I => n4029, ZN => n8784);
   U21576 : NAND2_X2 port map( A1 => n29106, A2 => n7543, ZN => n4029);
   U21577 : OAI21_X2 port map( A1 => n33473, A2 => n31822, B => n716, ZN => 
                           n17022);
   U21585 : XOR2_X1 port map( A1 => n31165, A2 => n22197, Z => n14969);
   U21586 : NAND2_X2 port map( A1 => n31037, A2 => n33475, ZN => n24965);
   U21591 : NAND3_X1 port map( A1 => n2886, A2 => n1221, A3 => n716, ZN => 
                           n33475);
   U21595 : XOR2_X1 port map( A1 => n33476, A2 => n34056, Z => n33638);
   U21597 : OAI21_X2 port map( A1 => n29570, A2 => n34168, B => n32004, ZN => 
                           n30394);
   U21599 : XOR2_X1 port map( A1 => n33477, A2 => n20870, Z => n14887);
   U21601 : XOR2_X1 port map( A1 => n2055, A2 => n20955, Z => n33477);
   U21610 : XOR2_X1 port map( A1 => n3987, A2 => n33478, Z => n29762);
   U21612 : XOR2_X1 port map( A1 => n33574, A2 => n4997, Z => n33478);
   U21618 : XOR2_X1 port map( A1 => n33479, A2 => n12284, Z => n31272);
   U21623 : XOR2_X1 port map( A1 => n30492, A2 => n3617, Z => n33479);
   U21624 : XOR2_X1 port map( A1 => n14612, A2 => n23191, Z => n23192);
   U21626 : INV_X2 port map( I => n6552, ZN => n33480);
   U21629 : INV_X2 port map( I => n33482, ZN => n10086);
   U21635 : XNOR2_X1 port map( A1 => n2366, A2 => n2364, ZN => n33482);
   U21636 : NOR2_X1 port map( A1 => n15680, A2 => n21546, ZN => n33483);
   U21640 : INV_X2 port map( I => n23150, ZN => n1261);
   U21641 : NAND3_X2 port map( A1 => n393, A2 => n18239, A3 => n28178, ZN => 
                           n23150);
   U21642 : XOR2_X1 port map( A1 => n10946, A2 => n11862, Z => n12915);
   U21647 : XOR2_X1 port map( A1 => n33484, A2 => n12896, Z => n34122);
   U21649 : XOR2_X1 port map( A1 => n19557, A2 => n27884, Z => n33484);
   U21670 : XOR2_X1 port map( A1 => n11781, A2 => n33486, Z => n11641);
   U21678 : XOR2_X1 port map( A1 => n10946, A2 => n22141, Z => n33486);
   U21692 : XOR2_X1 port map( A1 => n24810, A2 => n7879, Z => n13858);
   U21697 : NAND2_X2 port map( A1 => n6110, A2 => n5960, ZN => n33760);
   U21701 : INV_X2 port map( I => n33487, ZN => n29153);
   U21705 : NAND2_X2 port map( A1 => n9171, A2 => n11785, ZN => n33909);
   U21712 : AOI21_X2 port map( A1 => n23812, A2 => n3860, B => n11061, ZN => 
                           n33488);
   U21717 : NOR2_X1 port map( A1 => n33867, A2 => n23595, ZN => n23584);
   U21718 : NAND2_X1 port map( A1 => n9283, A2 => n9282, ZN => n33489);
   U21722 : XOR2_X1 port map( A1 => n23422, A2 => n23421, Z => n33490);
   U21736 : NOR2_X2 port map( A1 => n10973, A2 => n33491, ZN => n10721);
   U21744 : NOR3_X1 port map( A1 => n7007, A2 => n21379, A3 => n17313, ZN => 
                           n33491);
   U21745 : XOR2_X1 port map( A1 => n24562, A2 => n24563, Z => n24564);
   U21746 : XOR2_X1 port map( A1 => n26795, A2 => n24819, Z => n24562);
   U21748 : NOR2_X2 port map( A1 => n14189, A2 => n33494, ZN => n25175);
   U21749 : XOR2_X1 port map( A1 => n32648, A2 => n31950, Z => n2785);
   U21753 : NAND2_X2 port map( A1 => n349, A2 => n21218, ZN => n33495);
   U21754 : OAI22_X2 port map( A1 => n10871, A2 => n28825, B1 => n22606, B2 => 
                           n5961, ZN => n6110);
   U21755 : XOR2_X1 port map( A1 => n5186, A2 => n21011, Z => n5185);
   U21767 : NOR2_X2 port map( A1 => n33497, A2 => n31811, ZN => n7154);
   U21768 : NOR2_X2 port map( A1 => n20607, A2 => n7577, ZN => n33497);
   U21771 : INV_X1 port map( I => n33501, ZN => n17322);
   U21782 : AND2_X1 port map( A1 => n1465, A2 => n33501, Z => n34080);
   U21783 : INV_X2 port map( I => n13644, ZN => n13681);
   U21794 : NAND2_X2 port map( A1 => n7800, A2 => n31496, ZN => n13644);
   U21796 : OR2_X1 port map( A1 => n21392, A2 => n20882, Z => n20883);
   U21800 : NOR2_X2 port map( A1 => n20511, A2 => n16774, ZN => n20730);
   U21803 : XOR2_X1 port map( A1 => n33448, A2 => n19508, Z => n19588);
   U21807 : NAND2_X2 port map( A1 => n17507, A2 => n17509, ZN => n19508);
   U21812 : NAND2_X2 port map( A1 => n1684, A2 => n7392, ZN => n20970);
   U21820 : OR2_X1 port map( A1 => n18677, A2 => n18888, Z => n10367);
   U21825 : NAND2_X2 port map( A1 => n29089, A2 => n7316, ZN => n5150);
   U21831 : OAI22_X2 port map( A1 => n4994, A2 => n33502, B1 => n4996, B2 => 
                           n26878, ZN => n15501);
   U21832 : XOR2_X1 port map( A1 => n31597, A2 => n18189, Z => n27633);
   U21842 : NAND2_X2 port map( A1 => n10705, A2 => n14868, ZN => n18189);
   U21845 : XOR2_X1 port map( A1 => n8659, A2 => n23455, Z => n7178);
   U21848 : NAND2_X2 port map( A1 => n14371, A2 => n33505, ZN => n17301);
   U21851 : NAND2_X2 port map( A1 => n24189, A2 => n24186, ZN => n8412);
   U21856 : XOR2_X1 port map( A1 => n12653, A2 => n31638, Z => n31468);
   U21862 : XOR2_X1 port map( A1 => n33506, A2 => n16666, Z => Ciphertext(81));
   U21863 : NAND2_X1 port map( A1 => n4226, A2 => n31281, ZN => n33506);
   U21865 : INV_X2 port map( I => n33508, ZN => n11869);
   U21870 : NOR2_X2 port map( A1 => n5000, A2 => n5002, ZN => n9300);
   U21871 : INV_X2 port map( I => n33510, ZN => n29462);
   U21900 : XOR2_X1 port map( A1 => n30747, A2 => n5482, Z => n10519);
   U21902 : XOR2_X1 port map( A1 => n33511, A2 => n4555, Z => n17857);
   U21903 : XOR2_X1 port map( A1 => n4554, A2 => n4559, Z => n33511);
   U21906 : NOR2_X2 port map( A1 => n5668, A2 => n5669, ZN => n20690);
   U21908 : NAND2_X1 port map( A1 => n33499, A2 => n17181, ZN => n26570);
   U21909 : AND2_X1 port map( A1 => n16809, A2 => n16380, Z => n1949);
   U21910 : NAND2_X2 port map( A1 => n24894, A2 => n14274, ZN => n16809);
   U21911 : XOR2_X1 port map( A1 => n33513, A2 => n16322, Z => Ciphertext(136))
                           ;
   U21912 : XOR2_X1 port map( A1 => n22141, A2 => n22055, Z => n22206);
   U21914 : INV_X2 port map( I => n33514, ZN => n12058);
   U21923 : NAND2_X2 port map( A1 => n29976, A2 => n15641, ZN => n33514);
   U21926 : NAND2_X1 port map( A1 => n21427, A2 => n21338, ZN => n21339);
   U21935 : NOR2_X2 port map( A1 => n9994, A2 => n21826, ZN => n28278);
   U21938 : NAND2_X2 port map( A1 => n34015, A2 => n5687, ZN => n21826);
   U21944 : BUF_X2 port map( I => n7102, Z => n33515);
   U21946 : INV_X2 port map( I => n10001, ZN => n819);
   U21947 : OAI22_X2 port map( A1 => n1976, A2 => n16491, B1 => n1974, B2 => 
                           n10742, ZN => n10001);
   U21948 : AND2_X1 port map( A1 => n31437, A2 => n17462, Z => n28777);
   U21954 : XOR2_X1 port map( A1 => n2388, A2 => n19403, Z => n19543);
   U21955 : OAI21_X2 port map( A1 => n1871, A2 => n2390, B => n16788, ZN => 
                           n2388);
   U21956 : XOR2_X1 port map( A1 => n33517, A2 => n24766, Z => n15106);
   U21960 : XOR2_X1 port map( A1 => n30358, A2 => n24764, Z => n33517);
   U21966 : XOR2_X1 port map( A1 => n30532, A2 => n23282, Z => n23173);
   U21971 : XOR2_X1 port map( A1 => n2072, A2 => n33518, Z => n26854);
   U21973 : XOR2_X1 port map( A1 => n8741, A2 => n29876, Z => n33518);
   U21974 : NAND2_X2 port map( A1 => n28463, A2 => n31006, ZN => n3614);
   U21975 : XOR2_X1 port map( A1 => Plaintext(168), A2 => Key(168), Z => n17030
                           );
   U21978 : XOR2_X1 port map( A1 => n7015, A2 => n33521, Z => n3879);
   U21979 : XOR2_X1 port map( A1 => n10075, A2 => n10935, Z => n12621);
   U21981 : NAND2_X2 port map( A1 => n29729, A2 => n33524, ZN => n6865);
   U21993 : NAND2_X2 port map( A1 => n33526, A2 => n33525, ZN => n33524);
   U22001 : NAND2_X2 port map( A1 => n33527, A2 => n3087, ZN => n3086);
   U22003 : NOR2_X2 port map( A1 => n29659, A2 => n33558, ZN => n33528);
   U22004 : NAND2_X2 port map( A1 => n33529, A2 => n33730, ZN => n3036);
   U22005 : INV_X2 port map( I => n10524, ZN => n33529);
   U22007 : NAND2_X2 port map( A1 => n31967, A2 => n3084, ZN => n10524);
   U22020 : XOR2_X1 port map( A1 => n1787, A2 => n14428, Z => n11532);
   U22028 : AND2_X1 port map( A1 => n24324, A2 => n30579, Z => n2360);
   U22031 : NAND2_X2 port map( A1 => n8, A2 => n8086, ZN => n30579);
   U22032 : BUF_X2 port map( I => n29763, Z => n33530);
   U22037 : XOR2_X1 port map( A1 => n23529, A2 => n23287, Z => n14584);
   U22038 : XOR2_X1 port map( A1 => n4627, A2 => n15686, Z => n17151);
   U22044 : INV_X2 port map( I => n33531, ZN => n29688);
   U22045 : XOR2_X1 port map( A1 => n5607, A2 => n5609, Z => n33531);
   U22053 : XOR2_X1 port map( A1 => n24760, A2 => n10084, Z => n24743);
   U22056 : NAND3_X2 port map( A1 => n8000, A2 => n8001, A3 => n24228, ZN => 
                           n24760);
   U22070 : NAND3_X1 port map( A1 => n4916, A2 => n34058, A3 => n14251, ZN => 
                           n22351);
   U22074 : NOR2_X2 port map( A1 => n16559, A2 => n12074, ZN => n18641);
   U22077 : OR2_X1 port map( A1 => n13431, A2 => n13430, Z => n33533);
   U22084 : INV_X2 port map( I => n33534, ZN => n4916);
   U22091 : NAND2_X2 port map( A1 => n275, A2 => n9299, ZN => n22318);
   U22092 : AOI21_X2 port map( A1 => n11309, A2 => n23697, B => n33535, ZN => 
                           n11287);
   U22099 : XOR2_X1 port map( A1 => n24422, A2 => n24423, Z => n10172);
   U22102 : CLKBUF_X12 port map( I => n9870, Z => n33536);
   U22105 : XOR2_X1 port map( A1 => n21029, A2 => n12342, Z => n20764);
   U22110 : NOR2_X2 port map( A1 => n12343, A2 => n12344, ZN => n12342);
   U22113 : NAND2_X2 port map( A1 => n2961, A2 => n33537, ZN => n13684);
   U22114 : INV_X2 port map( I => n33538, ZN => n21160);
   U22117 : OAI22_X2 port map( A1 => n18277, A2 => n18641, B1 => n18276, B2 => 
                           n4626, ZN => n18279);
   U22132 : XOR2_X1 port map( A1 => n14908, A2 => n16502, Z => n15990);
   U22140 : NAND2_X2 port map( A1 => n11070, A2 => n30743, ZN => n14908);
   U22152 : AND2_X1 port map( A1 => n17590, A2 => n21160, Z => n12521);
   U22155 : XOR2_X1 port map( A1 => n33539, A2 => n24798, Z => n10209);
   U22166 : XOR2_X1 port map( A1 => n24597, A2 => n27283, Z => n33539);
   U22183 : NAND2_X1 port map( A1 => n27514, A2 => n30673, ZN => n33650);
   U22185 : OAI22_X2 port map( A1 => n17767, A2 => n21078, B1 => n21079, B2 => 
                           n16933, ZN => n15622);
   U22189 : NAND2_X2 port map( A1 => n33541, A2 => n10928, ZN => n23065);
   U22190 : NAND2_X1 port map( A1 => n8427, A2 => n10654, ZN => n33541);
   U22218 : AOI21_X2 port map( A1 => n33542, A2 => n33830, B => n23584, ZN => 
                           n16643);
   U22225 : NOR2_X2 port map( A1 => n6082, A2 => n21401, ZN => n28426);
   U22230 : NAND2_X2 port map( A1 => n21403, A2 => n596, ZN => n21401);
   U22231 : NOR2_X2 port map( A1 => n20070, A2 => n18036, ZN => n27600);
   U22236 : XOR2_X1 port map( A1 => n2520, A2 => n25879, Z => n30421);
   U22242 : OAI22_X2 port map( A1 => n2404, A2 => n2405, B1 => n17202, B2 => 
                           n22895, ZN => n2520);
   U22245 : XOR2_X1 port map( A1 => n2626, A2 => n33545, Z => n18090);
   U22247 : XOR2_X1 port map( A1 => n2628, A2 => n15188, Z => n33545);
   U22248 : NAND2_X2 port map( A1 => n18677, A2 => n10325, ZN => n10364);
   U22249 : XOR2_X1 port map( A1 => n23258, A2 => n23376, Z => n23181);
   U22254 : OAI21_X2 port map( A1 => n12529, A2 => n22906, B => n14914, ZN => 
                           n23258);
   U22260 : XOR2_X1 port map( A1 => n32697, A2 => n19461, Z => n5921);
   U22261 : NAND3_X2 port map( A1 => n28372, A2 => n28371, A3 => n6193, ZN => 
                           n31568);
   U22264 : INV_X1 port map( I => n1652, ZN => n21461);
   U22265 : OAI22_X2 port map( A1 => n28396, A2 => n21058, B1 => n21263, B2 => 
                           n11745, ZN => n1652);
   U22266 : NAND2_X1 port map( A1 => n15500, A2 => n15498, ZN => n33546);
   U22269 : XOR2_X1 port map( A1 => n18058, A2 => n22255, Z => n17486);
   U22270 : XOR2_X1 port map( A1 => n33547, A2 => n25567, Z => Ciphertext(128))
                           ;
   U22280 : NAND4_X2 port map( A1 => n10035, A2 => n37, A3 => n10039, A4 => n36
                           , ZN => n33547);
   U22281 : NOR2_X2 port map( A1 => n12525, A2 => n20780, ZN => n28420);
   U22282 : NAND2_X1 port map( A1 => n10511, A2 => n10510, ZN => n27282);
   U22285 : NAND3_X2 port map( A1 => n10446, A2 => n10448, A3 => n10450, ZN => 
                           n5762);
   U22288 : NAND3_X1 port map( A1 => n22463, A2 => n22462, A3 => n22557, ZN => 
                           n22464);
   U22294 : NAND2_X2 port map( A1 => n22462, A2 => n22460, ZN => n22463);
   U22297 : XOR2_X1 port map( A1 => n31884, A2 => n16958, Z => n2925);
   U22302 : NAND2_X2 port map( A1 => n6775, A2 => n14366, ZN => n16958);
   U22303 : NAND2_X2 port map( A1 => n25025, A2 => n16293, ZN => n25123);
   U22305 : OAI22_X2 port map( A1 => n21571, A2 => n29806, B1 => n1012, B2 => 
                           n32039, ZN => n3578);
   U22310 : XOR2_X1 port map( A1 => n33550, A2 => n9550, Z => n665);
   U22313 : XOR2_X1 port map( A1 => n33552, A2 => n7596, Z => n28236);
   U22315 : XOR2_X1 port map( A1 => n30778, A2 => n3559, Z => n33552);
   U22316 : XOR2_X1 port map( A1 => n17301, A2 => n24442, Z => n24825);
   U22318 : XOR2_X1 port map( A1 => n7603, A2 => n24532, Z => n7135);
   U22326 : NOR2_X2 port map( A1 => n6334, A2 => n17067, ZN => n24532);
   U22327 : AND2_X1 port map( A1 => n18405, A2 => n5139, Z => n3052);
   U22335 : OAI21_X2 port map( A1 => n33553, A2 => n33909, B => n5717, ZN => 
                           n8087);
   U22336 : XOR2_X1 port map( A1 => n24749, A2 => n33554, Z => n7695);
   U22337 : XOR2_X1 port map( A1 => n11651, A2 => n10070, Z => n33554);
   U22339 : XOR2_X1 port map( A1 => n16175, A2 => n20798, Z => n9674);
   U22345 : XNOR2_X1 port map( A1 => n31279, A2 => n25856, ZN => n33838);
   U22348 : NAND3_X2 port map( A1 => n5485, A2 => n2935, A3 => n19039, ZN => 
                           n33555);
   U22349 : NAND2_X2 port map( A1 => n33556, A2 => n26767, ZN => n7045);
   U22352 : BUF_X2 port map( I => n24224, Z => n33557);
   U22354 : NAND3_X1 port map( A1 => n801, A2 => n28367, A3 => n23695, ZN => 
                           n10160);
   U22355 : INV_X4 port map( I => n17930, ZN => n896);
   U22356 : NAND2_X2 port map( A1 => n3711, A2 => n34053, ZN => n17930);
   U22360 : NOR2_X2 port map( A1 => n33645, A2 => n7602, ZN => n7604);
   U22365 : XOR2_X1 port map( A1 => n20999, A2 => n21000, Z => n21005);
   U22366 : INV_X2 port map( I => n28010, ZN => n33558);
   U22378 : BUF_X2 port map( I => n578, Z => n33561);
   U22379 : NOR2_X2 port map( A1 => n33595, A2 => n29705, ZN => n2005);
   U22381 : XOR2_X1 port map( A1 => n1536, A2 => n1538, Z => n7699);
   U22385 : XOR2_X1 port map( A1 => n14181, A2 => n15561, Z => n28312);
   U22390 : NAND2_X2 port map( A1 => n11317, A2 => n4750, ZN => n33562);
   U22392 : INV_X2 port map( I => n1112, ZN => n33563);
   U22394 : XOR2_X1 port map( A1 => n6746, A2 => n33575, Z => n14398);
   U22398 : NAND2_X2 port map( A1 => n7541, A2 => n33564, ZN => n7802);
   U22402 : AOI22_X2 port map( A1 => n13665, A2 => n13664, B1 => n26878, B2 => 
                           n908, ZN => n33564);
   U22422 : NOR2_X2 port map( A1 => n12168, A2 => n33264, ZN => n33565);
   U22431 : NOR2_X2 port map( A1 => n13541, A2 => n10398, ZN => n19530);
   U22438 : XOR2_X1 port map( A1 => n19672, A2 => n26683, Z => n6156);
   U22441 : NAND2_X2 port map( A1 => n28237, A2 => n14735, ZN => n19672);
   U22443 : INV_X2 port map( I => n14321, ZN => n24994);
   U22445 : NAND2_X2 port map( A1 => n12679, A2 => n12678, ZN => n14321);
   U22454 : AOI21_X2 port map( A1 => n16873, A2 => n4210, B => n16870, ZN => 
                           n30411);
   U22456 : OR3_X1 port map( A1 => n29695, A2 => n28812, A3 => n20489, Z => 
                           n20254);
   U22459 : INV_X2 port map( I => n33570, ZN => n27343);
   U22464 : BUF_X2 port map( I => n21820, Z => n33571);
   U22466 : BUF_X2 port map( I => n22317, Z => n33572);
   U22468 : NAND2_X2 port map( A1 => n33573, A2 => n11008, ZN => n13694);
   U22472 : NAND2_X1 port map( A1 => n11010, A2 => n8252, ZN => n33573);
   U22473 : NAND2_X1 port map( A1 => n1619, A2 => n6003, ZN => n33727);
   U22478 : XOR2_X1 port map( A1 => n6745, A2 => n15424, Z => n33575);
   U22485 : NAND2_X2 port map( A1 => n33576, A2 => n9794, ZN => n16147);
   U22488 : NOR2_X2 port map( A1 => n2724, A2 => n2725, ZN => n33576);
   U22491 : NAND2_X2 port map( A1 => n384, A2 => n11103, ZN => n16134);
   U22492 : NAND2_X2 port map( A1 => n33577, A2 => n6663, ZN => n7852);
   U22503 : AOI22_X2 port map( A1 => n29284, A2 => n16298, B1 => n20116, B2 => 
                           n20118, ZN => n33577);
   U22505 : XOR2_X1 port map( A1 => n33578, A2 => n32074, Z => n30445);
   U22509 : XOR2_X1 port map( A1 => n6218, A2 => n20979, Z => n33578);
   U22513 : XOR2_X1 port map( A1 => n24419, A2 => n33579, Z => n28819);
   U22516 : OAI21_X1 port map( A1 => n9251, A2 => n786, B => n33580, ZN => 
                           n10587);
   U22517 : AOI22_X1 port map( A1 => n3988, A2 => n4953, B1 => n4952, B2 => 
                           n27149, ZN => n33580);
   U22520 : BUF_X2 port map( I => n946, Z => n33581);
   U22521 : NAND2_X1 port map( A1 => n30384, A2 => n30383, ZN => n33582);
   U22525 : XOR2_X1 port map( A1 => n12721, A2 => n20775, Z => n20756);
   U22527 : NAND2_X2 port map( A1 => n34045, A2 => n20585, ZN => n12721);
   U22528 : XOR2_X1 port map( A1 => n11897, A2 => n23519, Z => n26338);
   U22532 : XOR2_X1 port map( A1 => n12478, A2 => n20784, Z => n20925);
   U22533 : XOR2_X1 port map( A1 => n28968, A2 => n17869, Z => n17867);
   U22534 : XOR2_X1 port map( A1 => n27344, A2 => n33584, Z => n28496);
   U22535 : XOR2_X1 port map( A1 => n24800, A2 => n1227, Z => n33584);
   U22536 : NOR3_X1 port map( A1 => n15134, A2 => n13764, A3 => n31236, ZN => 
                           n15133);
   U22537 : OAI22_X1 port map( A1 => n8722, A2 => n25130, B1 => n8723, B2 => 
                           n712, ZN => n27664);
   U22540 : XOR2_X1 port map( A1 => n18042, A2 => n24647, Z => n9868);
   U22548 : XOR2_X1 port map( A1 => n6547, A2 => n24573, Z => n24647);
   U22549 : AOI21_X2 port map( A1 => n33615, A2 => n27443, B => n32020, ZN => 
                           n25317);
   U22561 : XOR2_X1 port map( A1 => n11862, A2 => n33587, Z => n21918);
   U22564 : INV_X1 port map( I => n24861, ZN => n33587);
   U22565 : NAND3_X2 port map( A1 => n9473, A2 => n12156, A3 => n12157, ZN => 
                           n23271);
   U22567 : BUF_X2 port map( I => n12493, Z => n33588);
   U22570 : NOR2_X2 port map( A1 => n6661, A2 => n14092, ZN => n33589);
   U22582 : XOR2_X1 port map( A1 => n23518, A2 => n33590, Z => n31751);
   U22587 : XOR2_X1 port map( A1 => n8068, A2 => n16373, Z => n23518);
   U22598 : XOR2_X1 port map( A1 => n30528, A2 => n16693, Z => n29772);
   U22605 : NOR2_X2 port map( A1 => n28782, A2 => n28783, ZN => n17460);
   U22606 : NAND3_X1 port map( A1 => n22642, A2 => n6297, A3 => n22645, ZN => 
                           n22337);
   U22612 : XOR2_X1 port map( A1 => n32404, A2 => n33593, Z => n31380);
   U22626 : NAND2_X2 port map( A1 => n29605, A2 => n5671, ZN => n12800);
   U22635 : AND2_X1 port map( A1 => n10673, A2 => n23706, Z => n23634);
   U22636 : BUF_X2 port map( I => n5226, Z => n33597);
   U22643 : NAND2_X1 port map( A1 => n26390, A2 => n9127, ZN => n33599);
   U22648 : NAND2_X2 port map( A1 => n10926, A2 => n27879, ZN => n20471);
   U22649 : NAND2_X2 port map( A1 => n695, A2 => n33600, ZN => n2236);
   U22653 : NOR2_X2 port map( A1 => n10251, A2 => n32023, ZN => n33600);
   U22657 : NOR2_X2 port map( A1 => n33602, A2 => n33601, ZN => n5790);
   U22661 : NAND2_X2 port map( A1 => n28351, A2 => n33603, ZN => n33602);
   U22663 : NAND3_X2 port map( A1 => n26667, A2 => n33132, A3 => n18261, ZN => 
                           n1564);
   U22669 : NOR2_X1 port map( A1 => n7868, A2 => n11401, ZN => n21556);
   U22672 : NAND2_X2 port map( A1 => n13152, A2 => n13150, ZN => n11401);
   U22676 : NOR2_X1 port map( A1 => n17956, A2 => n21220, ZN => n10837);
   U22677 : XOR2_X1 port map( A1 => n17400, A2 => n32050, Z => n17766);
   U22679 : XOR2_X1 port map( A1 => n31340, A2 => n24624, Z => n33604);
   U22681 : XOR2_X1 port map( A1 => n4790, A2 => n2142, Z => n7665);
   U22683 : XOR2_X1 port map( A1 => n20789, A2 => n20890, Z => n28405);
   U22685 : NAND2_X2 port map( A1 => n21545, A2 => n21544, ZN => n22157);
   U22686 : NOR2_X2 port map( A1 => n18672, A2 => n18881, ZN => n18517);
   U22687 : INV_X2 port map( I => n18879, ZN => n18672);
   U22689 : XOR2_X1 port map( A1 => n18354, A2 => Key(8), Z => n18879);
   U22690 : NAND2_X2 port map( A1 => n3137, A2 => n33605, ZN => n3629);
   U22692 : NOR2_X2 port map( A1 => n28269, A2 => n28268, ZN => n33605);
   U22694 : XOR2_X1 port map( A1 => n7705, A2 => n21028, Z => n21031);
   U22715 : XOR2_X1 port map( A1 => n33607, A2 => n10249, Z => n10303);
   U22716 : XOR2_X1 port map( A1 => n7288, A2 => n33747, Z => n33607);
   U22724 : BUF_X2 port map( I => n29757, Z => n33608);
   U22726 : AOI22_X1 port map( A1 => n1830, A2 => n1832, B1 => n1833, B2 => 
                           n7555, ZN => n33612);
   U22731 : NAND2_X2 port map( A1 => n5075, A2 => n5077, ZN => n8617);
   U22736 : XOR2_X1 port map( A1 => n33609, A2 => n23315, Z => n17797);
   U22740 : XOR2_X1 port map( A1 => n29299, A2 => n23332, Z => n23315);
   U22743 : XOR2_X1 port map( A1 => n33612, A2 => n1390, Z => Ciphertext(58));
   U22745 : XOR2_X1 port map( A1 => n33613, A2 => n33614, Z => n29916);
   U22747 : XOR2_X1 port map( A1 => n11062, A2 => n29955, Z => n33614);
   U22752 : OAI21_X2 port map( A1 => n33761, A2 => n13985, B => n31060, ZN => 
                           n33615);
   U22757 : INV_X2 port map( I => n33617, ZN => n18156);
   U22761 : XOR2_X1 port map( A1 => n33618, A2 => n20918, Z => n28998);
   U22763 : XOR2_X1 port map( A1 => n29918, A2 => n20652, Z => n33618);
   U22772 : XOR2_X1 port map( A1 => n8973, A2 => n8975, Z => n27960);
   U22784 : NAND2_X1 port map( A1 => n30888, A2 => n3901, ZN => n33767);
   U22791 : NAND2_X2 port map( A1 => n31629, A2 => n33619, ZN => n2860);
   U22793 : AOI22_X2 port map( A1 => n19188, A2 => n33672, B1 => n12316, B2 => 
                           n9538, ZN => n31682);
   U22794 : NOR2_X2 port map( A1 => n1883, A2 => n14597, ZN => n19188);
   U22796 : OAI21_X2 port map( A1 => n11112, A2 => n11409, B => n25306, ZN => 
                           n33620);
   U22800 : XOR2_X1 port map( A1 => n24173, A2 => n33622, Z => n24181);
   U22801 : XOR2_X1 port map( A1 => n15368, A2 => n6050, Z => n33622);
   U22802 : INV_X2 port map( I => n28181, ZN => n15772);
   U22803 : OR2_X1 port map( A1 => n28181, A2 => n17416, Z => n21348);
   U22805 : INV_X1 port map( I => n22271, ZN => n22218);
   U22806 : XOR2_X1 port map( A1 => n22271, A2 => n24759, Z => n29350);
   U22810 : XOR2_X1 port map( A1 => n16073, A2 => n23336, Z => n23496);
   U22812 : NAND2_X2 port map( A1 => n20594, A2 => n20599, ZN => n10379);
   U22815 : INV_X4 port map( I => n25806, ZN => n9181);
   U22819 : NAND2_X2 port map( A1 => n8759, A2 => n33623, ZN => n20577);
   U22821 : AOI22_X2 port map( A1 => n11587, A2 => n17696, B1 => n16243, B2 => 
                           n19971, ZN => n33623);
   U22828 : XOR2_X1 port map( A1 => n33905, A2 => n31725, Z => n28142);
   U22831 : OAI21_X2 port map( A1 => n31082, A2 => n30060, B => n6932, ZN => 
                           n29785);
   U22836 : NAND2_X2 port map( A1 => n33626, A2 => n33625, ZN => n33752);
   U22837 : BUF_X2 port map( I => n34151, Z => n33627);
   U22838 : XOR2_X1 port map( A1 => n24646, A2 => n15508, Z => n24563);
   U22841 : NAND2_X2 port map( A1 => n7884, A2 => n7883, ZN => n24646);
   U22846 : AOI21_X2 port map( A1 => n29849, A2 => n3236, B => n7377, ZN => 
                           n7620);
   U22851 : NOR2_X2 port map( A1 => n5395, A2 => n505, ZN => n7377);
   U22861 : BUF_X2 port map( I => n10871, Z => n33628);
   U22862 : AOI22_X2 port map( A1 => n24467, A2 => n27128, B1 => n31378, B2 => 
                           n1221, ZN => n24947);
   U22863 : NOR2_X1 port map( A1 => n29666, A2 => n19885, ZN => n20058);
   U22868 : XOR2_X1 port map( A1 => n392, A2 => n32085, Z => n21356);
   U22873 : XOR2_X1 port map( A1 => n33995, A2 => n28082, Z => n13817);
   U22874 : NOR2_X2 port map( A1 => n6590, A2 => n33629, ZN => n2971);
   U22876 : OAI22_X2 port map( A1 => n34066, A2 => n6587, B1 => n829, B2 => 
                           n785, ZN => n33629);
   U22878 : AOI21_X2 port map( A1 => n21558, A2 => n38, B => n33630, ZN => 
                           n22317);
   U22881 : OAI22_X2 port map( A1 => n32079, A2 => n21817, B1 => n21820, B2 => 
                           n1015, ZN => n33630);
   U22883 : XOR2_X1 port map( A1 => n8761, A2 => n27548, Z => n8765);
   U22887 : XOR2_X1 port map( A1 => n20733, A2 => n20843, Z => n21003);
   U22889 : NOR2_X2 port map( A1 => n16858, A2 => n20496, ZN => n20843);
   U22892 : OAI22_X2 port map( A1 => n33631, A2 => n1028, B1 => n7228, B2 => 
                           n12917, ZN => n7253);
   U22899 : NAND2_X2 port map( A1 => n25845, A2 => n13944, ZN => n25851);
   U22908 : NAND2_X2 port map( A1 => n34044, A2 => n3447, ZN => n3718);
   U22919 : BUF_X2 port map( I => n1944, Z => n33633);
   U22932 : AOI21_X2 port map( A1 => n6063, A2 => n6064, B => n33634, ZN => 
                           n22361);
   U22938 : INV_X4 port map( I => n28553, ZN => n24249);
   U22940 : NAND2_X2 port map( A1 => n7357, A2 => n7356, ZN => n17400);
   U22941 : XOR2_X1 port map( A1 => n6545, A2 => n24770, Z => n2667);
   U22942 : NOR2_X2 port map( A1 => n17747, A2 => n6651, ZN => n6545);
   U22949 : XOR2_X1 port map( A1 => n16917, A2 => n13299, Z => n4291);
   U22951 : OAI21_X2 port map( A1 => n3305, A2 => n2045, B => n30248, ZN => 
                           n16917);
   U22952 : XOR2_X1 port map( A1 => n23391, A2 => n9153, Z => n10289);
   U22953 : AND2_X1 port map( A1 => n9578, A2 => n12952, Z => n15920);
   U22964 : XOR2_X1 port map( A1 => n27211, A2 => n24693, Z => n27851);
   U22971 : XOR2_X1 port map( A1 => n24753, A2 => n24853, Z => n24693);
   U22972 : OR2_X1 port map( A1 => n26120, A2 => n23748, Z => n24074);
   U22974 : XOR2_X1 port map( A1 => n7638, A2 => n7639, Z => n33636);
   U22983 : XOR2_X1 port map( A1 => n33637, A2 => n16738, Z => n31655);
   U22990 : XOR2_X1 port map( A1 => n27458, A2 => n7466, Z => n33637);
   U22994 : XOR2_X1 port map( A1 => n33638, A2 => n23314, Z => n7616);
   U23000 : OAI21_X2 port map( A1 => n31768, A2 => n111, B => n8998, ZN => 
                           n33639);
   U23001 : NOR2_X2 port map( A1 => n21858, A2 => n29523, ZN => n21856);
   U23006 : AOI21_X2 port map( A1 => n30067, A2 => n29911, B => n24099, ZN => 
                           n24927);
   U23008 : XOR2_X1 port map( A1 => n33642, A2 => n20711, Z => n15047);
   U23009 : XOR2_X1 port map( A1 => n2356, A2 => n1343, Z => n33642);
   U23011 : AND2_X2 port map( A1 => n4224, A2 => n33856, Z => n13859);
   U23024 : OR2_X1 port map( A1 => n22831, A2 => n4110, Z => n9473);
   U23025 : NOR2_X1 port map( A1 => n34064, A2 => n11215, ZN => n1557);
   U23037 : XOR2_X1 port map( A1 => n11665, A2 => n7705, Z => n8189);
   U23039 : NOR2_X1 port map( A1 => n15039, A2 => n32119, ZN => n23092);
   U23040 : NAND3_X2 port map( A1 => n23964, A2 => n10046, A3 => n18120, ZN => 
                           n33645);
   U23042 : NOR2_X2 port map( A1 => n33646, A2 => n15328, ZN => n15324);
   U23047 : XOR2_X1 port map( A1 => n20767, A2 => n20768, Z => n10707);
   U23054 : XOR2_X1 port map( A1 => n21009, A2 => n20715, Z => n20768);
   U23059 : XOR2_X1 port map( A1 => n19599, A2 => n2483, Z => n19542);
   U23062 : NAND2_X1 port map( A1 => n33647, A2 => n21175, ZN => n13316);
   U23064 : NAND2_X1 port map( A1 => n31894, A2 => n985, ZN => n7221);
   U23066 : OR2_X1 port map( A1 => n4327, A2 => n11677, Z => n25943);
   U23070 : NOR2_X1 port map( A1 => n1480, A2 => n1235, ZN => n33648);
   U23077 : OAI21_X2 port map( A1 => n25886, A2 => n4318, B => n2182, ZN => 
                           n34069);
   U23080 : XOR2_X1 port map( A1 => n2592, A2 => n8138, Z => n26511);
   U23087 : XOR2_X1 port map( A1 => n9222, A2 => n23237, Z => n26889);
   U23093 : XOR2_X1 port map( A1 => n8695, A2 => n23430, Z => n23237);
   U23095 : XOR2_X1 port map( A1 => n27850, A2 => n22132, Z => n22183);
   U23096 : XOR2_X1 port map( A1 => n33651, A2 => n23505, Z => n30964);
   U23108 : XOR2_X1 port map( A1 => n31251, A2 => n33652, Z => n9744);
   U23120 : XOR2_X1 port map( A1 => n20711, A2 => n20642, Z => n33652);
   U23121 : OR2_X2 port map( A1 => n2655, A2 => n33536, Z => n22450);
   U23127 : NAND2_X2 port map( A1 => n33654, A2 => n33653, ZN => n23679);
   U23130 : NAND2_X2 port map( A1 => n24198, A2 => n33655, ZN => n33654);
   U23132 : NAND2_X2 port map( A1 => n1241, A2 => n24304, ZN => n24198);
   U23133 : OR2_X1 port map( A1 => n7287, A2 => n14402, Z => n33657);
   U23134 : XOR2_X1 port map( A1 => n19536, A2 => n400, Z => n30016);
   U23135 : XOR2_X1 port map( A1 => n19676, A2 => n19779, Z => n19536);
   U23144 : XOR2_X1 port map( A1 => n19409, A2 => n25598, Z => n8055);
   U23146 : NAND2_X1 port map( A1 => n27531, A2 => n25445, ZN => n33658);
   U23149 : XOR2_X1 port map( A1 => n27055, A2 => n11422, Z => n8133);
   U23152 : NAND2_X2 port map( A1 => n23354, A2 => n31058, ZN => n24106);
   U23157 : NAND2_X2 port map( A1 => n33660, A2 => n29575, ZN => n17361);
   U23165 : NOR2_X2 port map( A1 => n15245, A2 => n30717, ZN => n33660);
   U23168 : NAND2_X2 port map( A1 => n20309, A2 => n33661, ZN => n30749);
   U23176 : AOI22_X2 port map( A1 => n29432, A2 => n31961, B1 => n28626, B2 => 
                           n2134, ZN => n33661);
   U23184 : XOR2_X1 port map( A1 => n33662, A2 => n23188, Z => n23025);
   U23185 : XOR2_X1 port map( A1 => n9369, A2 => n30550, Z => n9235);
   U23194 : XOR2_X1 port map( A1 => n11481, A2 => n5476, Z => n9369);
   U23196 : XOR2_X1 port map( A1 => n15630, A2 => n17830, Z => n8464);
   U23198 : XOR2_X1 port map( A1 => n30013, A2 => n31477, Z => n17830);
   U23202 : XOR2_X1 port map( A1 => n33663, A2 => n15484, Z => n17047);
   U23205 : NAND2_X2 port map( A1 => n18379, A2 => n12534, ZN => n29146);
   U23206 : OR2_X1 port map( A1 => n25116, A2 => n18156, Z => n25117);
   U23209 : XOR2_X1 port map( A1 => n31568, A2 => n6488, Z => n33665);
   U23212 : NAND2_X2 port map( A1 => n11442, A2 => n31124, ZN => n30234);
   U23213 : XOR2_X1 port map( A1 => n9300, A2 => n13508, Z => n24624);
   U23215 : NAND3_X2 port map( A1 => n34079, A2 => n17943, A3 => n24266, ZN => 
                           n13508);
   U23217 : XOR2_X1 port map( A1 => n29652, A2 => n10332, Z => n20711);
   U23227 : OAI22_X2 port map( A1 => n10324, A2 => n11839, B1 => n11840, B2 => 
                           n4077, ZN => n29652);
   U23229 : AOI22_X2 port map( A1 => n1573, A2 => n24873, B1 => n5662, B2 => 
                           n8758, ZN => n33666);
   U23230 : AOI21_X2 port map( A1 => n1446, A2 => n8395, B => n18800, ZN => 
                           n1449);
   U23231 : NOR2_X1 port map( A1 => n3790, A2 => n10465, ZN => n19381);
   U23234 : OAI21_X2 port map( A1 => n12322, A2 => n8611, B => n5347, ZN => 
                           n14179);
   U23258 : OAI21_X2 port map( A1 => n15405, A2 => n15404, B => n8095, ZN => 
                           n33668);
   U23262 : NAND3_X2 port map( A1 => n2004, A2 => n2003, A3 => n2005, ZN => 
                           n2396);
   U23282 : NAND2_X1 port map( A1 => n2141, A2 => n33669, ZN => n2398);
   U23283 : XOR2_X1 port map( A1 => n23535, A2 => n27708, Z => n23234);
   U23291 : NAND2_X2 port map( A1 => n3513, A2 => n3512, ZN => n23535);
   U23295 : AOI22_X2 port map( A1 => n33671, A2 => n18621, B1 => n18626, B2 => 
                           n26550, ZN => n4619);
   U23304 : OAI21_X1 port map( A1 => n15660, A2 => n14939, B => n10470, ZN => 
                           n23973);
   U23306 : NOR2_X2 port map( A1 => n30282, A2 => n976, ZN => n15660);
   U23308 : BUF_X2 port map( I => n9885, Z => n33672);
   U23309 : XOR2_X1 port map( A1 => n19632, A2 => n31415, Z => n17552);
   U23323 : NAND2_X2 port map( A1 => n33775, A2 => n33674, ZN => n3181);
   U23329 : AOI22_X2 port map( A1 => n7407, A2 => n23901, B1 => n7406, B2 => 
                           n1254, ZN => n33674);
   U23336 : XOR2_X1 port map( A1 => n19503, A2 => n9161, Z => n9160);
   U23349 : XOR2_X1 port map( A1 => n26623, A2 => n31057, Z => n19503);
   U23358 : AOI22_X2 port map( A1 => n18376, A2 => n4626, B1 => n32127, B2 => 
                           n18375, ZN => n12534);
   U23362 : XOR2_X1 port map( A1 => n33677, A2 => n1392, Z => Ciphertext(54));
   U23364 : NOR3_X2 port map( A1 => n29227, A2 => n6814, A3 => n27518, ZN => 
                           n33677);
   U23366 : XOR2_X1 port map( A1 => n526, A2 => n6571, Z => n33678);
   U23375 : OR3_X1 port map( A1 => n12952, A2 => n22597, A3 => n4378, Z => 
                           n22512);
   U23376 : AOI21_X1 port map( A1 => n11113, A2 => n29815, B => n15291, ZN => 
                           n33719);
   U23377 : NOR2_X2 port map( A1 => n7233, A2 => n12051, ZN => n29815);
   U23378 : INV_X2 port map( I => n2396, ZN => n33680);
   U23379 : NAND2_X2 port map( A1 => n31707, A2 => n1525, ZN => n24243);
   U23380 : NAND2_X2 port map( A1 => n347, A2 => n2577, ZN => n2576);
   U23383 : NAND3_X2 port map( A1 => n4922, A2 => n4920, A3 => n14860, ZN => 
                           n347);
   U23384 : NAND2_X2 port map( A1 => n29681, A2 => n30802, ZN => n2209);
   U23388 : NAND2_X2 port map( A1 => n3592, A2 => n3590, ZN => n30763);
   U23389 : INV_X1 port map( I => n25703, ZN => n7041);
   U23394 : NAND2_X1 port map( A1 => n25703, A2 => n33681, ZN => n11595);
   U23396 : XOR2_X1 port map( A1 => n17653, A2 => n24392, Z => n25703);
   U23403 : XNOR2_X1 port map( A1 => n3028, A2 => n3026, ZN => n33950);
   U23413 : XOR2_X1 port map( A1 => n21007, A2 => n25218, Z => n15802);
   U23416 : NAND2_X2 port map( A1 => n27611, A2 => n4965, ZN => n21007);
   U23417 : XOR2_X1 port map( A1 => n4701, A2 => n34118, Z => n11364);
   U23422 : NAND2_X1 port map( A1 => n4049, A2 => n28281, ZN => n33689);
   U23446 : XOR2_X1 port map( A1 => n33685, A2 => n23289, Z => n27882);
   U23465 : XOR2_X1 port map( A1 => n7011, A2 => n29082, Z => n33685);
   U23484 : XNOR2_X1 port map( A1 => n15801, A2 => n16803, ZN => n28254);
   U23486 : NAND2_X1 port map( A1 => n31561, A2 => n31467, ZN => n29360);
   U23502 : NAND2_X2 port map( A1 => n19290, A2 => n19021, ZN => n2799);
   U23506 : AOI22_X2 port map( A1 => n17394, A2 => n10206, B1 => n1286, B2 => 
                           n856, ZN => n33690);
   U23507 : NOR2_X2 port map( A1 => n7283, A2 => n26164, ZN => n7108);
   U23511 : BUF_X2 port map( I => n28471, Z => n33691);
   U23514 : NAND2_X2 port map( A1 => n33692, A2 => n8391, ZN => n21707);
   U23515 : NAND2_X1 port map( A1 => n8468, A2 => n8466, ZN => n33692);
   U23517 : XOR2_X1 port map( A1 => n33698, A2 => n33693, Z => n479);
   U23520 : NAND3_X2 port map( A1 => n15109, A2 => n15111, A3 => n30355, ZN => 
                           n33694);
   U23522 : NAND2_X1 port map( A1 => n15441, A2 => n9518, ZN => n33695);
   U23529 : OAI21_X1 port map( A1 => n18537, A2 => n1184, B => n18539, ZN => 
                           n9420);
   U23532 : NOR2_X2 port map( A1 => n14624, A2 => n14198, ZN => n19359);
   U23548 : NAND2_X2 port map( A1 => n33696, A2 => n13172, ZN => n31290);
   U23551 : OAI21_X2 port map( A1 => n29774, A2 => n30022, B => n32481, ZN => 
                           n33696);
   U23554 : OAI22_X2 port map( A1 => n9176, A2 => n18969, B1 => n17593, B2 => 
                           n10472, ZN => n33749);
   U23567 : XOR2_X1 port map( A1 => n33697, A2 => n14701, Z => n29642);
   U23568 : XOR2_X1 port map( A1 => n30338, A2 => n32065, Z => n33697);
   U23570 : XOR2_X1 port map( A1 => n5051, A2 => n14665, Z => n24473);
   U23573 : NAND2_X2 port map( A1 => n23703, A2 => n23702, ZN => n14665);
   U23576 : NAND3_X2 port map( A1 => n34001, A2 => n21576, A3 => n34000, ZN => 
                           n7545);
   U23577 : NAND2_X2 port map( A1 => n33981, A2 => n5170, ZN => n8753);
   U23580 : BUF_X2 port map( I => n3345, Z => n33700);
   U23587 : NOR2_X2 port map( A1 => n24218, A2 => n16554, ZN => n14386);
   U23594 : NOR2_X2 port map( A1 => n1355, A2 => n3944, ZN => n30603);
   U23595 : NAND2_X2 port map( A1 => n14974, A2 => n23786, ZN => n23877);
   U23596 : NAND2_X1 port map( A1 => n33703, A2 => n14443, ZN => n23703);
   U23598 : NAND2_X1 port map( A1 => n5437, A2 => n26674, ZN => n33703);
   U23599 : NOR2_X2 port map( A1 => n517, A2 => n21743, ZN => n21778);
   U23600 : XOR2_X1 port map( A1 => n33704, A2 => n1801, Z => n26345);
   U23601 : XOR2_X1 port map( A1 => n33984, A2 => n20887, Z => n33704);
   U23602 : INV_X2 port map( I => n19950, ZN => n6580);
   U23606 : XOR2_X1 port map( A1 => n22324, A2 => n33706, Z => n9168);
   U23609 : XOR2_X1 port map( A1 => n22322, A2 => n33707, Z => n33706);
   U23622 : XNOR2_X1 port map( A1 => n27860, A2 => n721, ZN => n33895);
   U23629 : AOI22_X2 port map( A1 => n27595, A2 => n31954, B1 => n2386, B2 => 
                           n14794, ZN => n33708);
   U23636 : NOR2_X1 port map( A1 => n33709, A2 => n11902, ZN => n15277);
   U23639 : NOR2_X1 port map( A1 => n29872, A2 => n579, ZN => n33709);
   U23641 : OAI21_X2 port map( A1 => n30477, A2 => n27329, B => n31959, ZN => 
                           n15521);
   U23646 : XOR2_X1 port map( A1 => n33710, A2 => n33711, Z => n15507);
   U23647 : XOR2_X1 port map( A1 => n2838, A2 => n29879, Z => n27506);
   U23653 : AND2_X1 port map( A1 => n9939, A2 => n15722, Z => n23688);
   U23658 : NOR3_X1 port map( A1 => n4286, A2 => n12593, A3 => n9220, ZN => 
                           n29370);
   U23663 : INV_X2 port map( I => n21553, ZN => n31042);
   U23664 : XOR2_X1 port map( A1 => n31523, A2 => n24968, Z => n33711);
   U23666 : AOI21_X2 port map( A1 => n31861, A2 => n33713, B => n12824, ZN => 
                           n12823);
   U23668 : OAI22_X2 port map( A1 => n22873, A2 => n18241, B1 => n27090, B2 => 
                           n4113, ZN => n33713);
   U23674 : XOR2_X1 port map( A1 => n33796, A2 => n19748, Z => n29986);
   U23675 : XOR2_X1 port map( A1 => n19436, A2 => n19583, Z => n19748);
   U23684 : NAND2_X2 port map( A1 => n29071, A2 => n11519, ZN => n19040);
   U23687 : XOR2_X1 port map( A1 => n15788, A2 => n19497, Z => n11580);
   U23688 : NAND2_X2 port map( A1 => n8645, A2 => n27628, ZN => n30894);
   U23690 : XOR2_X1 port map( A1 => n23173, A2 => n23247, Z => n23369);
   U23693 : NAND2_X2 port map( A1 => n33760, A2 => n13983, ZN => n22816);
   U23694 : XOR2_X1 port map( A1 => n23314, A2 => n26123, Z => n33715);
   U23696 : NAND3_X2 port map( A1 => n14708, A2 => n12114, A3 => n14709, ZN => 
                           n8633);
   U23697 : XOR2_X1 port map( A1 => n12750, A2 => n33716, Z => n29908);
   U23698 : XOR2_X1 port map( A1 => n30765, A2 => n32026, Z => n33716);
   U23705 : NAND2_X2 port map( A1 => n17756, A2 => n931, ZN => n20247);
   U23706 : NAND2_X2 port map( A1 => n32504, A2 => n5003, ZN => n17756);
   U23711 : NAND2_X2 port map( A1 => n3114, A2 => n3116, ZN => n3964);
   U23712 : AND2_X1 port map( A1 => n17245, A2 => n23944, Z => n23322);
   U23726 : OAI21_X1 port map( A1 => n10214, A2 => n24906, B => n33717, ZN => 
                           n9969);
   U23729 : NAND2_X1 port map( A1 => n792, A2 => n30289, ZN => n15175);
   U23731 : INV_X2 port map( I => n31650, ZN => n23912);
   U23740 : NAND2_X1 port map( A1 => n29965, A2 => n31650, ZN => n31667);
   U23743 : XOR2_X1 port map( A1 => n17889, A2 => n22223, Z => n17891);
   U23746 : NAND2_X2 port map( A1 => n4106, A2 => n29517, ZN => n24262);
   U23747 : XOR2_X1 port map( A1 => n23264, A2 => n6169, Z => n9644);
   U23749 : AOI21_X2 port map( A1 => n5261, A2 => n8127, B => n8126, ZN => 
                           n23264);
   U23754 : AOI21_X1 port map( A1 => n19851, A2 => n19987, B => n20000, ZN => 
                           n34101);
   U23763 : XOR2_X1 port map( A1 => n33959, A2 => n5445, Z => n34134);
   U23764 : INV_X2 port map( I => n13180, ZN => n33722);
   U23771 : NOR2_X2 port map( A1 => n28002, A2 => n30633, ZN => n23224);
   U23775 : XOR2_X1 port map( A1 => n23266, A2 => n23267, Z => n12538);
   U23779 : AOI22_X2 port map( A1 => n22853, A2 => n22888, B1 => n22852, B2 => 
                           n22851, ZN => n23266);
   U23780 : NAND3_X2 port map( A1 => n15312, A2 => n15313, A3 => n32014, ZN => 
                           n20371);
   U23793 : NAND3_X2 port map( A1 => n9186, A2 => n21237, A3 => n780, ZN => 
                           n34015);
   U23794 : XOR2_X1 port map( A1 => n13545, A2 => n25567, Z => n15986);
   U23795 : NAND2_X2 port map( A1 => n14957, A2 => n29369, ZN => n21688);
   U23808 : OAI21_X2 port map( A1 => n2793, A2 => n16137, B => n33723, ZN => 
                           n2502);
   U23809 : NAND2_X2 port map( A1 => n16137, A2 => n7090, ZN => n33723);
   U23813 : NOR2_X2 port map( A1 => n25234, A2 => n25235, ZN => n5611);
   U23815 : XOR2_X1 port map( A1 => n23534, A2 => n27860, Z => n23411);
   U23817 : NOR2_X2 port map( A1 => n33793, A2 => n34010, ZN => n10398);
   U23827 : XOR2_X1 port map( A1 => n2192, A2 => n20856, Z => n12736);
   U23855 : XOR2_X1 port map( A1 => n1993, A2 => n2989, Z => n20856);
   U23856 : INV_X2 port map( I => n25517, ZN => n1209);
   U23862 : NAND2_X2 port map( A1 => n33956, A2 => n26277, ZN => n25517);
   U23874 : OAI21_X2 port map( A1 => n12992, A2 => n9879, B => n4119, ZN => 
                           n26524);
   U23878 : XOR2_X1 port map( A1 => n30069, A2 => n30290, Z => n29720);
   U23879 : XOR2_X1 port map( A1 => n29241, A2 => n20775, Z => n20723);
   U23883 : XOR2_X1 port map( A1 => n33725, A2 => n25507, Z => Ciphertext(116))
                           ;
   U23884 : NOR3_X2 port map( A1 => n25504, A2 => n30165, A3 => n33772, ZN => 
                           n33725);
   U23889 : XOR2_X1 port map( A1 => n27790, A2 => n33726, Z => n25228);
   U23893 : XOR2_X1 port map( A1 => n24575, A2 => n28807, Z => n33726);
   U23898 : XOR2_X1 port map( A1 => n29912, A2 => n4302, Z => n25111);
   U23901 : AND2_X1 port map( A1 => n21218, A2 => n21220, Z => n29900);
   U23911 : OAI21_X2 port map( A1 => n3643, A2 => n32060, B => n13796, ZN => 
                           n30174);
   U23912 : NAND3_X2 port map( A1 => n31868, A2 => n26488, A3 => n33912, ZN => 
                           n3694);
   U23914 : NAND2_X2 port map( A1 => n8905, A2 => n13647, ZN => n30209);
   U23917 : NAND2_X1 port map( A1 => n29690, A2 => n7182, ZN => n10442);
   U23922 : NAND2_X2 port map( A1 => n31960, A2 => n6442, ZN => n21518);
   U23929 : NAND2_X1 port map( A1 => n33729, A2 => n18631, ZN => n3251);
   U23930 : XOR2_X1 port map( A1 => n17622, A2 => Key(124), Z => n18631);
   U23931 : INV_X1 port map( I => n17143, ZN => n33729);
   U23941 : OR2_X1 port map( A1 => n33731, A2 => n5795, Z => n3979);
   U23945 : NAND2_X2 port map( A1 => n8442, A2 => n25521, ZN => n31236);
   U23950 : XOR2_X1 port map( A1 => Plaintext(185), A2 => Key(185), Z => n18869
                           );
   U23967 : OR2_X1 port map( A1 => n22340, A2 => n16306, Z => n22024);
   U23969 : OAI22_X2 port map( A1 => n14690, A2 => n1246, B1 => n24200, B2 => 
                           n24311, ZN => n3345);
   U23970 : NAND2_X2 port map( A1 => n31619, A2 => n20780, ZN => n33774);
   U23974 : NOR2_X1 port map( A1 => n31504, A2 => n29763, ZN => n8650);
   U23975 : AOI22_X2 port map( A1 => n21652, A2 => n29234, B1 => n31511, B2 => 
                           n17354, ZN => n34096);
   U23980 : NAND2_X2 port map( A1 => n261, A2 => n28567, ZN => n22951);
   U23983 : XOR2_X1 port map( A1 => n33733, A2 => n25190, Z => Ciphertext(67));
   U23987 : NAND3_X2 port map( A1 => n9705, A2 => n9704, A3 => n25189, ZN => 
                           n33733);
   U23991 : XOR2_X1 port map( A1 => n7348, A2 => n25252, Z => n22208);
   U23998 : XOR2_X1 port map( A1 => n24761, A2 => n24796, Z => n24695);
   U24002 : INV_X2 port map( I => n33734, ZN => n29365);
   U24003 : NAND2_X2 port map( A1 => n9856, A2 => n33737, ZN => n25557);
   U24005 : NOR2_X1 port map( A1 => n7236, A2 => n7237, ZN => n33738);
   U24008 : NAND2_X2 port map( A1 => n25387, A2 => n33876, ZN => n25452);
   U24021 : OR2_X2 port map( A1 => n17405, A2 => n31248, Z => n1699);
   U24022 : XNOR2_X1 port map( A1 => n3781, A2 => n22166, ZN => n2309);
   U24024 : NAND2_X2 port map( A1 => n33906, A2 => n4498, ZN => n9252);
   U24028 : INV_X2 port map( I => n30731, ZN => n33740);
   U24038 : INV_X2 port map( I => n22978, ZN => n6433);
   U24039 : NAND2_X2 port map( A1 => n17432, A2 => n31777, ZN => n17431);
   U24041 : XNOR2_X1 port map( A1 => n10935, A2 => n5848, ZN => n22061);
   U24042 : AOI22_X2 port map( A1 => n3226, A2 => n33691, B1 => n3227, B2 => 
                           n26567, ZN => n3439);
   U24048 : INV_X2 port map( I => n12478, ZN => n21048);
   U24059 : INV_X1 port map( I => n6611, ZN => n30404);
   U24060 : NAND2_X2 port map( A1 => n28087, A2 => n34153, ZN => n6611);
   U24062 : NAND2_X2 port map( A1 => n27285, A2 => n31965, ZN => n10546);
   U24066 : NAND2_X2 port map( A1 => n19235, A2 => n8119, ZN => n14054);
   U24068 : NAND2_X2 port map( A1 => n3403, A2 => n3402, ZN => n21045);
   U24070 : XOR2_X1 port map( A1 => n19627, A2 => n28601, Z => n33742);
   U24077 : XOR2_X1 port map( A1 => n19642, A2 => n29988, Z => n9103);
   U24079 : BUF_X2 port map( I => n14083, Z => n33743);
   U24081 : XOR2_X1 port map( A1 => n22149, A2 => n22192, Z => n10703);
   U24085 : NAND3_X2 port map( A1 => n6426, A2 => n21935, A3 => n21936, ZN => 
                           n22192);
   U24096 : XOR2_X1 port map( A1 => n28632, A2 => n25878, Z => n26765);
   U24098 : NAND2_X2 port map( A1 => n31889, A2 => n29878, ZN => n28632);
   U24099 : NOR2_X2 port map( A1 => n33744, A2 => n3798, ZN => n10705);
   U24100 : NAND2_X2 port map( A1 => n14153, A2 => n21574, ZN => n33744);
   U24101 : INV_X2 port map( I => n22810, ZN => n22715);
   U24104 : NOR2_X2 port map( A1 => n9071, A2 => n29717, ZN => n31309);
   U24108 : NAND2_X2 port map( A1 => n18322, A2 => n18321, ZN => n34082);
   U24110 : XOR2_X1 port map( A1 => n17798, A2 => n24849, Z => n5023);
   U24114 : NAND2_X2 port map( A1 => n27589, A2 => n22882, ZN => n27588);
   U24123 : AOI21_X2 port map( A1 => n33746, A2 => n4358, B => n8007, ZN => 
                           n1544);
   U24131 : NAND2_X2 port map( A1 => n936, A2 => n6255, ZN => n15053);
   U24136 : XOR2_X1 port map( A1 => n6852, A2 => n14125, Z => n33747);
   U24138 : XOR2_X1 port map( A1 => n9222, A2 => n7832, Z => n2969);
   U24144 : XOR2_X1 port map( A1 => n12821, A2 => n23253, Z => n7832);
   U24154 : XOR2_X1 port map( A1 => n33751, A2 => n20696, Z => n21184);
   U24157 : XOR2_X1 port map( A1 => n21042, A2 => n20796, Z => n33751);
   U24162 : NOR2_X2 port map( A1 => n31028, A2 => n33752, ZN => n26157);
   U24164 : OAI21_X1 port map( A1 => n33854, A2 => n22388, B => n33753, ZN => 
                           n22382);
   U24165 : NAND2_X2 port map( A1 => n30467, A2 => n33754, ZN => n12585);
   U24179 : AOI22_X1 port map( A1 => n33799, A2 => n18767, B1 => n18768, B2 => 
                           n28238, ZN => n33754);
   U24184 : NAND3_X2 port map( A1 => n317, A2 => n31149, A3 => n25331, ZN => 
                           n33874);
   U24185 : XOR2_X1 port map( A1 => n22029, A2 => n22216, Z => n22144);
   U24188 : AOI21_X2 port map( A1 => n33954, A2 => n33955, B => n21722, ZN => 
                           n22029);
   U24194 : NAND2_X1 port map( A1 => n31114, A2 => n16668, ZN => n33755);
   U24217 : XOR2_X1 port map( A1 => n20832, A2 => n31966, Z => n33756);
   U24219 : AND2_X1 port map( A1 => n8901, A2 => n11820, Z => n10454);
   U24221 : NOR2_X2 port map( A1 => n28227, A2 => n31549, ZN => n5252);
   U24229 : AOI21_X2 port map( A1 => n34043, A2 => n14964, B => n33757, ZN => 
                           n14960);
   U24234 : NOR2_X2 port map( A1 => n29339, A2 => n16491, ZN => n19932);
   U24239 : NAND2_X2 port map( A1 => n33758, A2 => n14896, ZN => n8790);
   U24247 : OAI21_X2 port map( A1 => n34081, A2 => n21439, B => n29933, ZN => 
                           n33758);
   U24248 : XOR2_X1 port map( A1 => n22107, A2 => n31649, Z => n28014);
   U24260 : NAND2_X2 port map( A1 => n23974, A2 => n23973, ZN => n26750);
   U24269 : NAND2_X2 port map( A1 => n33759, A2 => n23131, ZN => n3077);
   U24270 : NAND2_X2 port map( A1 => n9397, A2 => n9396, ZN => n28099);
   U24271 : NAND2_X2 port map( A1 => n33762, A2 => n11871, ZN => n6610);
   U24272 : OAI21_X2 port map( A1 => n17573, A2 => n17574, B => n11958, ZN => 
                           n33762);
   U24273 : BUF_X2 port map( I => n9919, Z => n33763);
   U24286 : OR2_X1 port map( A1 => n5032, A2 => n5034, Z => n1768);
   U24297 : XOR2_X1 port map( A1 => n23143, A2 => n6461, Z => n22385);
   U24309 : XOR2_X1 port map( A1 => n33764, A2 => n5145, Z => n17476);
   U24315 : XOR2_X1 port map( A1 => n29772, A2 => n24743, Z => n33764);
   U24318 : XOR2_X1 port map( A1 => n33765, A2 => n11784, Z => n31346);
   U24319 : XOR2_X1 port map( A1 => n28574, A2 => n28162, Z => n33765);
   U24328 : XNOR2_X1 port map( A1 => n23429, A2 => n1261, ZN => n28177);
   U24334 : OAI21_X2 port map( A1 => n9384, A2 => n5571, B => n4231, ZN => 
                           n23429);
   U24352 : NAND2_X1 port map( A1 => n1106, A2 => n16280, ZN => n14016);
   U24353 : XOR2_X1 port map( A1 => n20690, A2 => n1394, Z => n9274);
   U24361 : NAND2_X2 port map( A1 => n21974, A2 => n21975, ZN => n22795);
   U24368 : NAND2_X2 port map( A1 => n26961, A2 => n33768, ZN => n20492);
   U24370 : XOR2_X1 port map( A1 => n33770, A2 => n30899, Z => n30593);
   U24377 : INV_X4 port map( I => n6290, ZN => n19165);
   U24382 : NAND2_X2 port map( A1 => n7285, A2 => n7286, ZN => n6290);
   U24383 : OAI21_X2 port map( A1 => n29240, A2 => n739, B => n33771, ZN => 
                           n15585);
   U24391 : NAND2_X1 port map( A1 => n23888, A2 => n23713, ZN => n33771);
   U24395 : NOR2_X1 port map( A1 => n25510, A2 => n8766, ZN => n33772);
   U24397 : NAND2_X2 port map( A1 => n11180, A2 => n33773, ZN => n25657);
   U24399 : NOR3_X2 port map( A1 => n330, A2 => n783, A3 => n26130, ZN => 
                           n30546);
   U24443 : OAI21_X2 port map( A1 => n9137, A2 => n27474, B => n4340, ZN => 
                           n33775);
   U24447 : AOI21_X2 port map( A1 => n20296, A2 => n16218, B => n33776, ZN => 
                           n20299);
   U24452 : NAND2_X2 port map( A1 => n24212, A2 => n3718, ZN => n13458);
   U24453 : NAND2_X2 port map( A1 => n9986, A2 => n27904, ZN => n20479);
   U24454 : XOR2_X1 port map( A1 => n13321, A2 => n23511, Z => n13930);
   U24458 : NAND3_X1 port map( A1 => n28167, A2 => n32066, A3 => n5460, ZN => 
                           n26212);
   U24490 : NOR2_X1 port map( A1 => n29539, A2 => n686, ZN => n30998);
   U24502 : NAND2_X2 port map( A1 => n4488, A2 => n28487, ZN => n5512);
   U24503 : NAND2_X2 port map( A1 => n3748, A2 => n1775, ZN => n24149);
   U24507 : XOR2_X1 port map( A1 => n31660, A2 => n4831, Z => n33778);
   U24513 : AOI22_X2 port map( A1 => n29407, A2 => n32499, B1 => n21696, B2 => 
                           n21697, ZN => n21698);
   U24518 : NAND2_X1 port map( A1 => n13654, A2 => n10845, ZN => n34143);
   U24525 : INV_X2 port map( I => n17098, ZN => n33779);
   U24533 : NOR2_X2 port map( A1 => n26413, A2 => n5396, ZN => n17098);
   U24541 : XOR2_X1 port map( A1 => n3519, A2 => n23297, Z => n17859);
   U24542 : NAND2_X2 port map( A1 => n22618, A2 => n18056, ZN => n23297);
   U24547 : NAND3_X1 port map( A1 => n5239, A2 => n5395, A3 => n26677, ZN => 
                           n5238);
   U24551 : XOR2_X1 port map( A1 => n19557, A2 => n18072, Z => n1698);
   U24553 : XOR2_X1 port map( A1 => n33995, A2 => n8785, Z => n19557);
   U24565 : NAND3_X1 port map( A1 => n24340, A2 => n16552, A3 => n14840, ZN => 
                           n24341);
   U24567 : OAI21_X2 port map( A1 => n14314, A2 => n16395, B => n33780, ZN => 
                           n15144);
   U24568 : OAI21_X2 port map( A1 => n15789, A2 => n17623, B => n13554, ZN => 
                           n33780);
   U24571 : OAI21_X2 port map( A1 => n33781, A2 => n29282, B => n27491, ZN => 
                           n31218);
   U24572 : NOR2_X2 port map( A1 => n431, A2 => n28767, ZN => n33781);
   U24579 : XOR2_X1 port map( A1 => n33782, A2 => n11834, Z => n23899);
   U24581 : XOR2_X1 port map( A1 => n23390, A2 => n26888, Z => n33782);
   U24586 : XOR2_X1 port map( A1 => n2415, A2 => n2414, Z => n8398);
   U24588 : AOI21_X2 port map( A1 => n18431, A2 => n13554, B => n30001, ZN => 
                           n34107);
   U24590 : NOR2_X1 port map( A1 => n34101, A2 => n12300, ZN => n31062);
   U24592 : NAND2_X2 port map( A1 => n829, A2 => n33785, ZN => n33784);
   U24595 : NOR2_X2 port map( A1 => n13663, A2 => n11918, ZN => n33785);
   U24613 : BUF_X2 port map( I => n25979, Z => n33787);
   U24614 : OAI21_X2 port map( A1 => n23828, A2 => n1250, B => n34164, ZN => 
                           n3482);
   U24615 : INV_X2 port map( I => n29268, ZN => n33788);
   U24616 : INV_X2 port map( I => n33790, ZN => n10181);
   U24622 : XOR2_X1 port map( A1 => Plaintext(175), A2 => Key(175), Z => n33790
                           );
   U24639 : XOR2_X1 port map( A1 => n11218, A2 => n11222, Z => n11221);
   U24642 : OAI21_X2 port map( A1 => n32003, A2 => n33792, B => n33093, ZN => 
                           n8550);
   U24647 : NAND2_X1 port map( A1 => n33795, A2 => n33794, ZN => n33793);
   U24654 : INV_X1 port map( I => n29815, ZN => n33794);
   U24662 : XOR2_X1 port map( A1 => n33633, A2 => n30435, Z => n33796);
   U24671 : XOR2_X1 port map( A1 => n24674, A2 => n17811, Z => n5529);
   U24674 : INV_X2 port map( I => n9757, ZN => n34125);
   U24683 : NAND2_X1 port map( A1 => n28020, A2 => n28022, ZN => n33797);
   U24684 : AOI21_X2 port map( A1 => n33798, A2 => n1088, B => n24126, ZN => 
                           n10539);
   U24689 : NAND2_X2 port map( A1 => n24123, A2 => n17100, ZN => n33798);
   U24693 : OAI21_X2 port map( A1 => n29553, A2 => n27600, B => n20301, ZN => 
                           n13943);
   U24699 : NAND3_X2 port map( A1 => n32862, A2 => n974, A3 => n24234, ZN => 
                           n24030);
   U24700 : XOR2_X1 port map( A1 => n3416, A2 => n26456, Z => n19455);
   U24705 : INV_X2 port map( I => n33800, ZN => n29369);
   U24722 : NOR2_X2 port map( A1 => n21087, A2 => n28886, ZN => n33800);
   U24723 : XOR2_X1 port map( A1 => n7931, A2 => n33801, Z => n28608);
   U24726 : XOR2_X1 port map( A1 => n7178, A2 => n23452, Z => n33801);
   U24727 : AND2_X1 port map( A1 => n13318, A2 => n15467, Z => n29789);
   U24728 : INV_X2 port map( I => n33803, ZN => n9939);
   U24730 : XOR2_X1 port map( A1 => n9432, A2 => n26388, Z => n17899);
   U24733 : XOR2_X1 port map( A1 => n11667, A2 => n17775, Z => n33806);
   U24745 : NAND2_X2 port map( A1 => n2631, A2 => n2632, ZN => n11667);
   U24752 : XOR2_X1 port map( A1 => n33804, A2 => n11780, Z => n11083);
   U24756 : OAI21_X2 port map( A1 => n29355, A2 => n29626, B => n33805, ZN => 
                           n21981);
   U24767 : OAI21_X2 port map( A1 => n29597, A2 => n16240, B => n29626, ZN => 
                           n33805);
   U24781 : AND2_X1 port map( A1 => n5433, A2 => n33561, Z => n6953);
   U24786 : XOR2_X1 port map( A1 => n33806, A2 => n450, Z => n1454);
   U24788 : XOR2_X1 port map( A1 => n10585, A2 => n19518, Z => n5436);
   U24798 : XOR2_X1 port map( A1 => n10294, A2 => n19743, Z => n10585);
   U24799 : NAND2_X2 port map( A1 => n10383, A2 => n10382, ZN => n24053);
   U24809 : XOR2_X1 port map( A1 => n33807, A2 => n24968, Z => Ciphertext(21));
   U24811 : NAND3_X1 port map( A1 => n17330, A2 => n699, A3 => n3846, ZN => 
                           n33807);
   U24816 : NAND2_X2 port map( A1 => n16121, A2 => n1489, ZN => n23766);
   U24836 : INV_X2 port map( I => n33809, ZN => n29282);
   U24843 : NAND2_X2 port map( A1 => n16154, A2 => n8576, ZN => n33809);
   U24844 : AOI22_X1 port map( A1 => n22832, A2 => n17501, B1 => n22753, B2 => 
                           n15421, ZN => n30207);
   U24847 : XOR2_X1 port map( A1 => n23206, A2 => n33811, Z => n16829);
   U24853 : XOR2_X1 port map( A1 => n23262, A2 => n9153, Z => n23206);
   U24855 : NAND2_X2 port map( A1 => n24117, A2 => n24226, ZN => n24224);
   U24858 : NAND2_X2 port map( A1 => n18044, A2 => n15206, ZN => n24117);
   U24863 : NAND2_X2 port map( A1 => n7789, A2 => n30924, ZN => n22075);
   U24865 : XOR2_X1 port map( A1 => n20699, A2 => n1828, Z => n20593);
   U24868 : XOR2_X1 port map( A1 => Plaintext(76), A2 => Key(76), Z => n31099);
   U24871 : OAI22_X2 port map( A1 => n23903, A2 => n17157, B1 => n14975, B2 => 
                           n23786, ZN => n23448);
   U24873 : XNOR2_X1 port map( A1 => n22313, A2 => n7664, ZN => n33816);
   U24876 : AOI21_X2 port map( A1 => n20592, A2 => n1347, B => n30882, ZN => 
                           n33815);
   U24878 : NAND2_X1 port map( A1 => n10248, A2 => n686, ZN => n25624);
   U24879 : XOR2_X1 port map( A1 => n21726, A2 => n22145, Z => n21906);
   U24881 : NOR2_X2 port map( A1 => n26690, A2 => n6253, ZN => n22145);
   U24894 : XOR2_X1 port map( A1 => n2104, A2 => n33816, Z => n30994);
   U24898 : NAND2_X1 port map( A1 => n33818, A2 => n33817, ZN => n26109);
   U24901 : INV_X1 port map( I => n14600, ZN => n33818);
   U24906 : NAND2_X2 port map( A1 => n33819, A2 => n7698, ZN => n7717);
   U24908 : XOR2_X1 port map( A1 => n24473, A2 => n1507, Z => n10277);
   U24916 : AOI22_X2 port map( A1 => n2172, A2 => n30988, B1 => n2088, B2 => 
                           n2173, ZN => n33821);
   U24923 : BUF_X2 port map( I => n23417, Z => n33823);
   U24934 : NOR3_X2 port map( A1 => n19992, A2 => n28293, A3 => n17882, ZN => 
                           n7775);
   U24935 : XOR2_X1 port map( A1 => n30449, A2 => n27669, Z => n28109);
   U24954 : NAND3_X2 port map( A1 => n19850, A2 => n4663, A3 => n27345, ZN => 
                           n8016);
   U24958 : NAND2_X2 port map( A1 => n21134, A2 => n33826, ZN => n21715);
   U24965 : NAND2_X2 port map( A1 => n33829, A2 => n28265, ZN => n33828);
   U24966 : XOR2_X1 port map( A1 => n9670, A2 => n9672, Z => n11413);
   U24967 : NOR2_X1 port map( A1 => n12336, A2 => n14523, ZN => n33830);
   U24968 : OR2_X1 port map( A1 => n30172, A2 => n23770, Z => n33831);
   U24971 : NAND2_X2 port map( A1 => n13934, A2 => n27134, ZN => n3006);
   U24972 : AOI21_X2 port map( A1 => n1120, A2 => n34035, B => n28170, ZN => 
                           n2253);
   U24973 : INV_X2 port map( I => n29687, ZN => n21039);
   U24974 : XNOR2_X1 port map( A1 => n20766, A2 => n32467, ZN => n29687);
   U24986 : BUF_X2 port map( I => n8965, Z => n34035);
   U24987 : AOI21_X2 port map( A1 => n6138, A2 => n13788, B => n15406, ZN => 
                           n13202);
   U24988 : OAI21_X2 port map( A1 => n8937, A2 => n30730, B => n33888, ZN => 
                           n6784);
   U25003 : XOR2_X1 port map( A1 => n20993, A2 => n33836, Z => n13504);
   U25004 : XOR2_X1 port map( A1 => n8581, A2 => n29870, Z => n33836);
   U25008 : AOI22_X2 port map( A1 => n13448, A2 => n27941, B1 => n13450, B2 => 
                           n13449, ZN => n34119);
   U25018 : NAND2_X2 port map( A1 => n18443, A2 => n18881, ZN => n33837);
   U25029 : XOR2_X1 port map( A1 => n24372, A2 => n24829, Z => n8791);
   U25030 : XOR2_X1 port map( A1 => n24830, A2 => n24747, Z => n24372);
   U25032 : NAND2_X1 port map( A1 => n18537, A2 => n16042, ZN => n18538);
   U25033 : XOR2_X1 port map( A1 => n19579, A2 => n33838, Z => n231);
   U25040 : XOR2_X1 port map( A1 => n19658, A2 => n19698, Z => n19579);
   U25041 : XOR2_X1 port map( A1 => n23443, A2 => n32905, Z => n3635);
   U25043 : XOR2_X1 port map( A1 => n33839, A2 => n16355, Z => Ciphertext(70));
   U25044 : OAI22_X1 port map( A1 => n9675, A2 => n9676, B1 => n11365, B2 => 
                           n12060, ZN => n33839);
   U25045 : XOR2_X1 port map( A1 => n32604, A2 => n22208, Z => n33840);
   U25057 : XOR2_X1 port map( A1 => n2989, A2 => n20801, Z => n20987);
   U25058 : NAND2_X2 port map( A1 => n3035, A2 => n3036, ZN => n20801);
   U25061 : NAND2_X2 port map( A1 => n9905, A2 => n9906, ZN => n29937);
   U25062 : OAI21_X2 port map( A1 => n2368, A2 => n33842, B => n33841, ZN => 
                           n21558);
   U25063 : AOI21_X2 port map( A1 => n22910, A2 => n6433, B => n5345, ZN => 
                           n17871);
   U25065 : INV_X2 port map( I => n25571, ZN => n25577);
   U25066 : OAI22_X2 port map( A1 => n6640, A2 => n5929, B1 => n5930, B2 => 
                           n6641, ZN => n25571);
   U25069 : XOR2_X1 port map( A1 => n23271, A2 => n5904, Z => n23458);
   U25070 : XOR2_X1 port map( A1 => n17859, A2 => n23495, Z => n3518);
   U25072 : OR2_X1 port map( A1 => n25565, A2 => n25582, Z => n1473);
   U25073 : NOR2_X2 port map( A1 => n33844, A2 => n18907, ZN => n29801);
   U25080 : NOR2_X2 port map( A1 => n11798, A2 => n33845, ZN => n33844);
   U25087 : NOR2_X2 port map( A1 => n19268, A2 => n18974, ZN => n33846);
   U25091 : XOR2_X1 port map( A1 => n33847, A2 => n28896, Z => n11089);
   U25093 : XOR2_X1 port map( A1 => n24561, A2 => n24451, Z => n33847);
   U25096 : XOR2_X1 port map( A1 => n24756, A2 => n13496, Z => n13163);
   U25097 : XOR2_X1 port map( A1 => n3295, A2 => n13060, Z => n24756);
   U25098 : XOR2_X1 port map( A1 => n13724, A2 => n34111, Z => n13723);
   U25104 : AOI21_X2 port map( A1 => n8957, A2 => n34054, B => n9395, ZN => 
                           n33850);
   U25108 : NAND2_X2 port map( A1 => n20010, A2 => n20008, ZN => n13585);
   U25112 : XOR2_X1 port map( A1 => n34024, A2 => n10985, Z => n5675);
   U25113 : XOR2_X1 port map( A1 => n3260, A2 => n19403, Z => n19504);
   U25115 : OAI21_X2 port map( A1 => n18789, A2 => n18790, B => n18788, ZN => 
                           n19403);
   U25129 : NOR2_X2 port map( A1 => n6530, A2 => n20325, ZN => n20324);
   U25135 : NAND2_X2 port map( A1 => n5225, A2 => n32051, ZN => n33999);
   U25140 : NAND2_X2 port map( A1 => n33852, A2 => n30012, ZN => n19520);
   U25141 : NAND2_X2 port map( A1 => n23766, A2 => n28676, ZN => n28745);
   U25142 : XOR2_X1 port map( A1 => n24683, A2 => n24579, Z => n17505);
   U25151 : XOR2_X1 port map( A1 => n2278, A2 => n32871, Z => n24579);
   U25154 : INV_X2 port map( I => n11576, ZN => n865);
   U25155 : XOR2_X1 port map( A1 => n5500, A2 => n11577, Z => n11576);
   U25160 : NAND2_X2 port map( A1 => n3501, A2 => n33855, ZN => n13191);
   U25163 : INV_X2 port map( I => n21876, ZN => n33857);
   U25170 : OR2_X1 port map( A1 => n17888, A2 => n33857, Z => n21590);
   U25176 : NAND2_X2 port map( A1 => n30798, A2 => n14262, ZN => n20892);
   U25192 : OAI22_X2 port map( A1 => n29422, A2 => n33858, B1 => n4443, B2 => 
                           n4442, ZN => n15715);
   U25196 : NOR2_X2 port map( A1 => n330, A2 => n4441, ZN => n33858);
   U25198 : XNOR2_X1 port map( A1 => n10169, A2 => n26030, ZN => n6604);
   U25206 : INV_X2 port map( I => n29322, ZN => n21629);
   U25208 : XOR2_X1 port map( A1 => n13520, A2 => n27950, Z => n33860);
   U25214 : OAI21_X2 port map( A1 => n33862, A2 => n33861, B => n29325, ZN => 
                           n3852);
   U25219 : AOI21_X2 port map( A1 => n33865, A2 => n22483, B => n33864, ZN => 
                           n33863);
   U25220 : OR2_X1 port map( A1 => n28723, A2 => n11089, Z => n8711);
   U25224 : XOR2_X1 port map( A1 => n16992, A2 => n23229, Z => n33866);
   U25232 : BUF_X2 port map( I => n29767, Z => n33868);
   U25235 : NAND3_X2 port map( A1 => n23636, A2 => n5227, A3 => n23635, ZN => 
                           n5226);
   U25244 : NOR2_X2 port map( A1 => n33869, A2 => n22366, ZN => n9377);
   U25245 : XOR2_X1 port map( A1 => n23496, A2 => n23494, Z => n3517);
   U25246 : NOR2_X2 port map( A1 => n5913, A2 => n31096, ZN => n33871);
   U25255 : XOR2_X1 port map( A1 => n3504, A2 => n7679, Z => n11217);
   U25257 : NAND3_X2 port map( A1 => n7668, A2 => n3216, A3 => n3217, ZN => 
                           n7679);
   U25263 : XOR2_X1 port map( A1 => n33873, A2 => n25911, Z => Ciphertext(189))
                           ;
   U25268 : NAND2_X2 port map( A1 => n13979, A2 => n33874, ZN => n30144);
   U25270 : XOR2_X1 port map( A1 => n19400, A2 => n19399, Z => n19546);
   U25286 : INV_X2 port map( I => n33875, ZN => n20065);
   U25292 : NAND3_X2 port map( A1 => n32029, A2 => n14139, A3 => n6551, ZN => 
                           n33876);
   U25296 : XOR2_X1 port map( A1 => n20588, A2 => n29850, Z => n33877);
   U25299 : NOR2_X2 port map( A1 => n30144, A2 => n33878, ZN => n25488);
   U25303 : NOR3_X2 port map( A1 => n28866, A2 => n25520, A3 => n25561, ZN => 
                           n33878);
   U25304 : NAND3_X1 port map( A1 => n14149, A2 => n25485, A3 => n33879, ZN => 
                           Ciphertext(112));
   U25306 : NAND3_X1 port map( A1 => n25481, A2 => n30117, A3 => n30118, ZN => 
                           n33879);
   U25313 : INV_X2 port map( I => n15212, ZN => n25446);
   U25314 : NAND3_X2 port map( A1 => n6818, A2 => n6817, A3 => n6990, ZN => 
                           n12868);
   U25316 : NAND2_X2 port map( A1 => n15529, A2 => n33880, ZN => n25276);
   U25321 : XOR2_X1 port map( A1 => n33881, A2 => n14526, Z => Ciphertext(89));
   U25327 : AOI22_X1 port map( A1 => n16291, A2 => n11294, B1 => n25286, B2 => 
                           n28532, ZN => n33881);
   U25330 : XOR2_X1 port map( A1 => n11304, A2 => n20977, Z => n6615);
   U25335 : XOR2_X1 port map( A1 => n13844, A2 => n23368, Z => n14527);
   U25349 : OAI21_X2 port map( A1 => n26732, A2 => n26731, B => n26710, ZN => 
                           n8078);
   U25355 : NAND2_X2 port map( A1 => n33883, A2 => n12527, ZN => n12617);
   U25359 : NAND2_X2 port map( A1 => n30720, A2 => n17580, ZN => n33883);
   U25362 : AOI22_X2 port map( A1 => n2039, A2 => n2040, B1 => n33885, B2 => 
                           n33884, ZN => n2037);
   U25368 : NOR2_X2 port map( A1 => n879, A2 => n880, ZN => n33885);
   U25369 : XOR2_X1 port map( A1 => n31234, A2 => n7137, Z => n27012);
   U25371 : OR2_X1 port map( A1 => n16987, A2 => n30346, Z => n21843);
   U25372 : NOR2_X1 port map( A1 => n8632, A2 => n31040, ZN => n30730);
   U25373 : OAI21_X2 port map( A1 => n33887, A2 => n10113, B => n33886, ZN => 
                           n8740);
   U25376 : INV_X2 port map( I => n21149, ZN => n33889);
   U25378 : INV_X2 port map( I => n33890, ZN => n17255);
   U25385 : XNOR2_X1 port map( A1 => Plaintext(78), A2 => Key(78), ZN => n33890
                           );
   U25386 : XOR2_X1 port map( A1 => n24675, A2 => n24487, Z => n24488);
   U25393 : NAND3_X2 port map( A1 => n12319, A2 => n10827, A3 => n12318, ZN => 
                           n24675);
   U25394 : NOR2_X1 port map( A1 => n11390, A2 => n18676, ZN => n2105);
   U25397 : INV_X1 port map( I => n12282, ZN => n18676);
   U25400 : XOR2_X1 port map( A1 => Key(14), A2 => Plaintext(14), Z => n12282);
   U25410 : NOR3_X1 port map( A1 => n30935, A2 => n749, A3 => n1204, ZN => 
                           n30165);
   U25419 : INV_X2 port map( I => n4782, ZN => n4953);
   U25422 : XOR2_X1 port map( A1 => n9218, A2 => n33893, Z => n26236);
   U25424 : XOR2_X1 port map( A1 => n21035, A2 => n5009, Z => n33893);
   U25428 : NAND2_X1 port map( A1 => n12900, A2 => n18026, ZN => n72);
   U25429 : AOI21_X1 port map( A1 => n27931, A2 => n26158, B => n24120, ZN => 
                           n10449);
   U25434 : OAI21_X2 port map( A1 => n5952, A2 => n5953, B => n15213, ZN => 
                           n5951);
   U25440 : NAND2_X2 port map( A1 => n33896, A2 => n6931, ZN => n20534);
   U25445 : XOR2_X1 port map( A1 => n16608, A2 => n32053, Z => n34135);
   U25450 : XOR2_X1 port map( A1 => n4321, A2 => n2611, Z => n16608);
   U25457 : XOR2_X1 port map( A1 => n33897, A2 => n15712, Z => n15711);
   U25463 : XOR2_X1 port map( A1 => n15293, A2 => n30565, Z => n33897);
   U25471 : NAND2_X1 port map( A1 => n33898, A2 => n19118, ZN => n13647);
   U25473 : OAI21_X2 port map( A1 => n3856, A2 => n18513, B => n18512, ZN => 
                           n19118);
   U25474 : NOR2_X1 port map( A1 => n19120, A2 => n13646, ZN => n33898);
   U25480 : NOR2_X1 port map( A1 => n27060, A2 => n10603, ZN => n33913);
   U25481 : NAND2_X2 port map( A1 => n1982, A2 => n13151, ZN => n21636);
   U25483 : NAND2_X2 port map( A1 => n34054, A2 => n5575, ZN => n13151);
   U25484 : INV_X1 port map( I => n16374, ZN => n20298);
   U25486 : NAND2_X1 port map( A1 => n33902, A2 => n16374, ZN => n29201);
   U25487 : NAND2_X2 port map( A1 => n34032, A2 => n17346, ZN => n16374);
   U25490 : INV_X2 port map( I => n28166, ZN => n33902);
   U25493 : INV_X2 port map( I => n33903, ZN => n28263);
   U25496 : XOR2_X1 port map( A1 => n16641, A2 => n13357, Z => n3209);
   U25498 : NAND2_X2 port map( A1 => n8502, A2 => n12629, ZN => n24836);
   U25508 : NAND2_X1 port map( A1 => n9058, A2 => n21509, ZN => n9057);
   U25513 : XOR2_X1 port map( A1 => n23246, A2 => n23244, Z => n30912);
   U25517 : XOR2_X1 port map( A1 => n15360, A2 => n13638, Z => n23244);
   U25519 : AOI21_X1 port map( A1 => n6475, A2 => n12563, B => n13693, ZN => 
                           n1962);
   U25520 : XOR2_X1 port map( A1 => n1825, A2 => n23230, Z => n23370);
   U25543 : NOR2_X2 port map( A1 => n26607, A2 => n6150, ZN => n1825);
   U25555 : XOR2_X1 port map( A1 => n17811, A2 => n24439, Z => n33905);
   U25556 : AOI22_X2 port map( A1 => n6016, A2 => n34154, B1 => n4855, B2 => 
                           n6961, ZN => n33906);
   U25559 : OAI21_X2 port map( A1 => n8235, A2 => n12090, B => n12602, ZN => 
                           n24171);
   U25563 : XOR2_X1 port map( A1 => n17973, A2 => n33910, Z => n26846);
   U25568 : XOR2_X1 port map( A1 => n17722, A2 => n32070, Z => n33910);
   U25575 : BUF_X2 port map( I => n27182, Z => n33911);
   U25578 : OAI22_X1 port map( A1 => n33913, A2 => n10600, B1 => n10604, B2 => 
                           n16653, ZN => Ciphertext(88));
   U25581 : NAND2_X2 port map( A1 => n33915, A2 => n33911, ZN => n33914);
   U25583 : INV_X4 port map( I => n16650, ZN => n33915);
   U25589 : AOI22_X2 port map( A1 => n3596, A2 => n22691, B1 => n1122, B2 => 
                           n30436, ZN => n28489);
   U25594 : XOR2_X1 port map( A1 => n5501, A2 => n31576, Z => n5504);
   U25605 : XOR2_X1 port map( A1 => n3117, A2 => n3118, Z => n33916);
   U25618 : NAND2_X2 port map( A1 => n3247, A2 => n31645, ZN => n27767);
   U25623 : XOR2_X1 port map( A1 => n11651, A2 => n3544, Z => n29538);
   U25629 : XOR2_X1 port map( A1 => n16971, A2 => n33917, Z => n27567);
   U25630 : XOR2_X1 port map( A1 => n22243, A2 => n33918, Z => n33917);
   U25631 : INV_X1 port map( I => n25364, ZN => n33918);
   U25632 : NAND3_X2 port map( A1 => n3310, A2 => n3309, A3 => n1036, ZN => 
                           n1678);
   U25633 : NAND2_X1 port map( A1 => n23771, A2 => n15116, ZN => n23772);
   U25635 : NAND2_X2 port map( A1 => n27459, A2 => n1610, ZN => n23771);
   U25638 : XOR2_X1 port map( A1 => n13727, A2 => n33920, Z => n34111);
   U25641 : XOR2_X1 port map( A1 => n31526, A2 => n1993, Z => n33920);
   U25642 : XOR2_X1 port map( A1 => n19378, A2 => n18102, Z => n4986);
   U25646 : NOR2_X2 port map( A1 => n26503, A2 => n18103, ZN => n19378);
   U25648 : NAND2_X2 port map( A1 => n26370, A2 => n7703, ZN => n22076);
   U25649 : INV_X2 port map( I => n33922, ZN => n14248);
   U25650 : XOR2_X1 port map( A1 => Plaintext(122), A2 => Key(122), Z => n33922
                           );
   U25652 : NAND2_X2 port map( A1 => n15303, A2 => n24007, ZN => n24442);
   U25653 : AND2_X1 port map( A1 => n10561, A2 => n18615, Z => n26442);
   U25655 : NAND3_X2 port map( A1 => n24867, A2 => n24667, A3 => n25536, ZN => 
                           n26277);
   U25657 : NAND2_X2 port map( A1 => n13693, A2 => n20329, ZN => n20410);
   U25661 : NAND2_X2 port map( A1 => n9413, A2 => n9097, ZN => n13693);
   U25663 : NAND2_X2 port map( A1 => n26012, A2 => n6131, ZN => n7809);
   U25665 : INV_X2 port map( I => n33928, ZN => n34163);
   U25666 : NAND3_X2 port map( A1 => n17001, A2 => n22555, A3 => n413, ZN => 
                           n33928);
   U25673 : XOR2_X1 port map( A1 => n33930, A2 => n2015, Z => n2013);
   U25676 : XOR2_X1 port map( A1 => n24493, A2 => n705, Z => n33930);
   U25678 : NAND4_X2 port map( A1 => n13598, A2 => n33932, A3 => n23094, A4 => 
                           n33931, ZN => n17278);
   U25679 : XOR2_X1 port map( A1 => n15161, A2 => n24770, Z => n33933);
   U25680 : INV_X2 port map( I => n33934, ZN => n25);
   U25690 : OR2_X1 port map( A1 => n31911, A2 => n21655, Z => n29947);
   U25694 : XOR2_X1 port map( A1 => n12923, A2 => n12921, Z => n33939);
   U25700 : XOR2_X1 port map( A1 => n22061, A2 => n33940, Z => n21990);
   U25703 : XOR2_X1 port map( A1 => n6771, A2 => n26942, Z => n33940);
   U25704 : NAND2_X2 port map( A1 => n27586, A2 => n25404, ZN => n1700);
   U25717 : OAI21_X2 port map( A1 => n16306, A2 => n22497, B => n25, ZN => 
                           n9108);
   U25725 : NAND2_X2 port map( A1 => n3801, A2 => n6455, ZN => n7881);
   U25726 : AND2_X1 port map( A1 => n17143, A2 => n14248, Z => n18821);
   U25728 : NAND3_X2 port map( A1 => n6597, A2 => n1853, A3 => n18511, ZN => 
                           n19042);
   U25734 : AOI21_X2 port map( A1 => n11949, A2 => n20147, B => n20148, ZN => 
                           n28911);
   U25741 : NOR3_X1 port map( A1 => n221, A2 => n25575, A3 => n5942, ZN => 
                           n33942);
   U25759 : XOR2_X1 port map( A1 => n33943, A2 => n24543, Z => n6008);
   U25762 : XOR2_X1 port map( A1 => n12313, A2 => n14762, Z => n24543);
   U25778 : XOR2_X1 port map( A1 => n28082, A2 => n19754, Z => n19476);
   U25781 : NAND2_X2 port map( A1 => n11801, A2 => n11800, ZN => n28082);
   U25783 : NOR2_X1 port map( A1 => n2613, A2 => n28344, ZN => n11880);
   U25788 : NAND2_X2 port map( A1 => n3124, A2 => n9801, ZN => n4908);
   U25789 : NAND2_X2 port map( A1 => n12891, A2 => n12894, ZN => n14214);
   U25793 : OR2_X1 port map( A1 => n32888, A2 => n14457, Z => n19851);
   U25801 : XOR2_X1 port map( A1 => n30258, A2 => n31857, Z => n30257);
   U25802 : NAND3_X2 port map( A1 => n15910, A2 => n29093, A3 => n19096, ZN => 
                           n13889);
   U25804 : NAND2_X1 port map( A1 => n15964, A2 => n25566, ZN => n13421);
   U25805 : INV_X2 port map( I => n33945, ZN => n6482);
   U25809 : XOR2_X1 port map( A1 => n28709, A2 => n22078, Z => n22079);
   U25810 : NAND2_X2 port map( A1 => n31263, A2 => n25444, ZN => n25418);
   U25811 : XOR2_X1 port map( A1 => n23521, A2 => n23522, Z => n23526);
   U25812 : AOI21_X2 port map( A1 => n31981, A2 => n14973, B => n23880, ZN => 
                           n17387);
   U25814 : NAND3_X2 port map( A1 => n33948, A2 => n14066, A3 => n33947, ZN => 
                           n16486);
   U25819 : NAND2_X2 port map( A1 => n29222, A2 => n30065, ZN => n33947);
   U25825 : BUF_X2 port map( I => n16440, Z => n33949);
   U25829 : INV_X2 port map( I => n8335, ZN => n19154);
   U25830 : XNOR2_X1 port map( A1 => n23404, A2 => n13638, ZN => n23502);
   U25832 : NAND2_X2 port map( A1 => n30853, A2 => n27695, ZN => n23404);
   U25833 : NOR2_X2 port map( A1 => n27814, A2 => n22981, ZN => n22839);
   U25836 : XOR2_X1 port map( A1 => n2143, A2 => n33950, Z => n30125);
   U25837 : NAND3_X2 port map( A1 => n24044, A2 => n24043, A3 => n33951, ZN => 
                           n24522);
   U25839 : NAND3_X2 port map( A1 => n4510, A2 => n34003, A3 => n13881, ZN => 
                           n13807);
   U25840 : NAND2_X2 port map( A1 => n25844, A2 => n25846, ZN => n16673);
   U25841 : NAND2_X2 port map( A1 => n25839, A2 => n25901, ZN => n25844);
   U25846 : XOR2_X1 port map( A1 => n12559, A2 => n20857, Z => n31295);
   U25848 : XOR2_X1 port map( A1 => n34067, A2 => n24751, Z => n27523);
   U25849 : XOR2_X1 port map( A1 => n24531, A2 => n2424, Z => n24751);
   U25851 : AOI22_X2 port map( A1 => n20093, A2 => n15192, B1 => n6027, B2 => 
                           n10768, ZN => n4075);
   U25852 : NAND2_X1 port map( A1 => n13242, A2 => n25987, ZN => n27265);
   U25853 : XOR2_X1 port map( A1 => n1848, A2 => n30664, Z => n33952);
   U25854 : XOR2_X1 port map( A1 => n30393, A2 => n29033, Z => n25118);
   U25856 : INV_X2 port map( I => n33953, ZN => n981);
   U25859 : XOR2_X1 port map( A1 => n15731, A2 => n6485, Z => n33953);
   U25862 : NOR2_X1 port map( A1 => n23816, A2 => n6759, ZN => n23817);
   U25863 : NAND2_X2 port map( A1 => n15732, A2 => n16431, ZN => n23816);
   U25864 : XOR2_X1 port map( A1 => n24843, A2 => n14645, Z => n10869);
   U25865 : NOR2_X2 port map( A1 => n7358, A2 => n28029, ZN => n14645);
   U25867 : XOR2_X1 port map( A1 => n8993, A2 => n4251, Z => n6407);
   U25869 : NAND2_X1 port map( A1 => n23938, A2 => n9939, ZN => n34165);
   U25875 : NOR2_X1 port map( A1 => n386, A2 => n11567, ZN => n10409);
   U25879 : INV_X2 port map( I => n2855, ZN => n386);
   U25880 : XOR2_X1 port map( A1 => n2857, A2 => n28286, Z => n2855);
   U25884 : MUX2_X1 port map( I0 => n24960, I1 => n24955, S => n24947, Z => 
                           n11428);
   U25888 : NAND2_X1 port map( A1 => n33957, A2 => n30523, ZN => n28952);
   U25889 : XOR2_X1 port map( A1 => n33958, A2 => n24953, Z => Ciphertext(14));
   U25896 : NAND2_X1 port map( A1 => n24667, A2 => n25390, ZN => n33961);
   U25897 : NAND2_X1 port map( A1 => n14763, A2 => n14635, ZN => n14634);
   U25899 : NAND2_X1 port map( A1 => n9227, A2 => n788, ZN => n14635);
   U25904 : NOR2_X1 port map( A1 => n14810, A2 => n28736, ZN => n6831);
   U25905 : NOR2_X2 port map( A1 => n27575, A2 => n34090, ZN => n7554);
   U25906 : AOI22_X2 port map( A1 => n18962, A2 => n16592, B1 => n31819, B2 => 
                           n33965, ZN => n19711);
   U25907 : XOR2_X1 port map( A1 => n24695, A2 => n24576, Z => n27362);
   U25908 : XOR2_X1 port map( A1 => n22075, A2 => n1433, Z => n7685);
   U25910 : NAND4_X2 port map( A1 => n26720, A2 => n20354, A3 => n26722, A4 => 
                           n20353, ZN => n20766);
   U25913 : XOR2_X1 port map( A1 => n26236, A2 => n33970, Z => n5392);
   U25916 : XOR2_X1 port map( A1 => n20785, A2 => n449, Z => n33970);
   U25919 : NAND3_X2 port map( A1 => n6865, A2 => n6866, A3 => n9015, ZN => 
                           n9287);
   U25926 : NAND3_X2 port map( A1 => n16514, A2 => n11204, A3 => n7625, ZN => 
                           n11205);
   U25928 : XOR2_X1 port map( A1 => n23344, A2 => n33973, Z => n3576);
   U25929 : XOR2_X1 port map( A1 => n1263, A2 => n23457, Z => n33973);
   U25930 : OAI21_X1 port map( A1 => n13032, A2 => n10497, B => n28097, ZN => 
                           n10393);
   U25931 : INV_X2 port map( I => n10392, ZN => n10497);
   U25932 : XOR2_X1 port map( A1 => n27526, A2 => n17159, Z => n10392);
   U25933 : AOI21_X2 port map( A1 => n16752, A2 => n25142, B => n1547, ZN => 
                           n25051);
   U25937 : INV_X2 port map( I => n14126, ZN => n31867);
   U25945 : NAND3_X2 port map( A1 => n29551, A2 => n22351, A3 => n10611, ZN => 
                           n14126);
   U25947 : NAND2_X2 port map( A1 => n8455, A2 => n26796, ZN => n23499);
   U25950 : XOR2_X1 port map( A1 => n22017, A2 => n31616, Z => n27669);
   U25959 : NAND3_X2 port map( A1 => n6145, A2 => n6146, A3 => n27529, ZN => 
                           n22225);
   U25960 : XOR2_X1 port map( A1 => n13067, A2 => n16584, Z => n31590);
   U25962 : OAI21_X2 port map( A1 => n29737, A2 => n16195, B => n21564, ZN => 
                           n13067);
   U25963 : NAND3_X2 port map( A1 => n4715, A2 => n4716, A3 => n9646, ZN => 
                           n4760);
   U25965 : INV_X2 port map( I => n33977, ZN => n30282);
   U25967 : XOR2_X1 port map( A1 => n30539, A2 => n5038, Z => n33977);
   U25968 : XOR2_X1 port map( A1 => n1762, A2 => n33978, Z => n16124);
   U25969 : XOR2_X1 port map( A1 => n26996, A2 => n22004, Z => n33978);
   U25970 : XOR2_X1 port map( A1 => n2117, A2 => n30795, Z => n7562);
   U25971 : NAND3_X1 port map( A1 => n785, A2 => n18515, A3 => n18639, ZN => 
                           n29492);
   U25978 : NAND2_X2 port map( A1 => n3919, A2 => n26391, ZN => n4655);
   U25979 : XOR2_X1 port map( A1 => n23343, A2 => n11249, Z => n13375);
   U25980 : XOR2_X1 port map( A1 => n34030, A2 => n30398, Z => n25883);
   U25981 : XOR2_X1 port map( A1 => n31288, A2 => n1980, Z => n16992);
   U25988 : AND3_X1 port map( A1 => n9328, A2 => n32890, A3 => n30820, Z => 
                           n29773);
   U25989 : XOR2_X1 port map( A1 => n7695, A2 => n29543, Z => n10420);
   U25990 : AOI21_X2 port map( A1 => n9177, A2 => n19146, B => n33983, ZN => 
                           n9904);
   U25994 : NAND2_X2 port map( A1 => n13548, A2 => n15146, ZN => n18546);
   U25995 : OAI22_X1 port map( A1 => n29323, A2 => n11922, B1 => n23755, B2 => 
                           n15399, ZN => n16224);
   U25996 : XOR2_X1 port map( A1 => n26929, A2 => n20885, Z => n33984);
   U26000 : NOR2_X2 port map( A1 => n8736, A2 => n8734, ZN => n33986);
   U26004 : NOR2_X1 port map( A1 => n21463, A2 => n33810, ZN => n26051);
   U26007 : XOR2_X1 port map( A1 => n2667, A2 => n2666, Z => n2665);
   U26008 : OR3_X1 port map( A1 => n1358, A2 => n16489, A3 => n17495, Z => 
                           n29844);
   U26009 : AOI21_X2 port map( A1 => n18691, A2 => n33988, B => n31987, ZN => 
                           n18694);
   U26011 : NAND2_X2 port map( A1 => n33989, A2 => n31971, ZN => n33988);
   U26014 : XOR2_X1 port map( A1 => n33991, A2 => n16604, Z => Ciphertext(142))
                           ;
   U26015 : NOR2_X2 port map( A1 => n29678, A2 => n15321, ZN => n15302);
   U26019 : NOR2_X2 port map( A1 => n33993, A2 => n27534, ZN => n12983);
   U26020 : NOR2_X1 port map( A1 => n14677, A2 => n9561, ZN => n33993);
   U26022 : XOR2_X1 port map( A1 => n24639, A2 => n33994, Z => n11843);
   U26026 : XOR2_X1 port map( A1 => n9145, A2 => n24638, Z => n33994);
   U26028 : OAI22_X2 port map( A1 => n7568, A2 => n7008, B1 => n19185, B2 => 
                           n29440, ZN => n8785);
   U26029 : NOR2_X2 port map( A1 => n8636, A2 => n9068, ZN => n8480);
   U26031 : NOR2_X1 port map( A1 => n34106, A2 => n27343, ZN => n34105);
   U26032 : NAND2_X2 port map( A1 => n2704, A2 => n9304, ZN => n29757);
   U26035 : NOR2_X2 port map( A1 => n9215, A2 => n33998, ZN => n33997);
   U26038 : OAI21_X2 port map( A1 => n7170, A2 => n32019, B => n7167, ZN => 
                           n28553);
   U26039 : XOR2_X1 port map( A1 => n14422, A2 => n8358, Z => n26934);
   U26040 : NOR2_X1 port map( A1 => n3782, A2 => n15255, ZN => n29362);
   U26041 : AOI21_X2 port map( A1 => n7400, A2 => n1291, B => n34002, ZN => 
                           n3801);
   U26042 : NAND3_X1 port map( A1 => n22637, A2 => n29626, A3 => n22636, ZN => 
                           n34003);
   U26045 : NOR2_X2 port map( A1 => n34004, A2 => n31022, ZN => n20819);
   U26049 : XOR2_X1 port map( A1 => n22067, A2 => n17555, Z => n21946);
   U26053 : NAND2_X2 port map( A1 => n2299, A2 => n2297, ZN => n17555);
   U26055 : XOR2_X1 port map( A1 => n10841, A2 => n6293, Z => n28950);
   U26058 : XOR2_X1 port map( A1 => n11102, A2 => n25500, Z => n3131);
   U26061 : NAND2_X2 port map( A1 => n3133, A2 => n3132, ZN => n11102);
   U26063 : XOR2_X1 port map( A1 => n16930, A2 => n14842, Z => n29919);
   U26064 : AND2_X1 port map( A1 => n20450, A2 => n20375, Z => n20201);
   U26065 : XOR2_X1 port map( A1 => n322, A2 => n24917, Z => n16717);
   U26077 : NAND2_X2 port map( A1 => n13834, A2 => n17411, ZN => n23376);
   U26081 : XOR2_X1 port map( A1 => n7469, A2 => n7472, Z => n25185);
   U26086 : NAND3_X2 port map( A1 => n16898, A2 => n27814, A3 => n29427, ZN => 
                           n34007);
   U26089 : XOR2_X1 port map( A1 => n4169, A2 => n8922, Z => n8933);
   U26093 : XOR2_X1 port map( A1 => n20888, A2 => n15268, Z => n4741);
   U26100 : XOR2_X1 port map( A1 => n20717, A2 => n30430, Z => n15268);
   U26104 : NOR2_X1 port map( A1 => n24347, A2 => n24346, ZN => n34011);
   U26105 : XOR2_X1 port map( A1 => n12494, A2 => n20825, Z => n21026);
   U26106 : INV_X1 port map( I => n22164, ZN => n1303);
   U26108 : XOR2_X1 port map( A1 => n22164, A2 => n34014, Z => n5884);
   U26109 : NOR2_X2 port map( A1 => n4124, A2 => n22978, ZN => n34017);
   U26111 : BUF_X2 port map( I => n19002, Z => n34018);
   U26123 : NAND3_X1 port map( A1 => n25729, A2 => n9495, A3 => n29331, ZN => 
                           n34019);
   U26127 : AOI21_X2 port map( A1 => n21367, A2 => n21369, B => n21163, ZN => 
                           n34059);
   U26135 : XOR2_X1 port map( A1 => n34020, A2 => n22307, Z => n2095);
   U26140 : XOR2_X1 port map( A1 => n32564, A2 => n4057, Z => n34020);
   U26141 : XOR2_X1 port map( A1 => n29644, A2 => n19627, Z => n19628);
   U26144 : NAND2_X2 port map( A1 => n26987, A2 => n26986, ZN => n20742);
   U26145 : INV_X2 port map( I => n11206, ZN => n859);
   U26150 : XOR2_X1 port map( A1 => n11206, A2 => n34021, Z => n22177);
   U26156 : INV_X1 port map( I => n16672, ZN => n34021);
   U26158 : NAND2_X2 port map( A1 => n28431, A2 => n10874, ZN => n11206);
   U26164 : NAND2_X1 port map( A1 => n10470, A2 => n26641, ZN => n2728);
   U26165 : XOR2_X1 port map( A1 => n34022, A2 => n20866, Z => n21210);
   U26169 : XOR2_X1 port map( A1 => n29734, A2 => n6465, Z => n34022);
   U26173 : NOR2_X2 port map( A1 => n11990, A2 => n28186, ZN => n12900);
   U26178 : NAND2_X2 port map( A1 => n18551, A2 => n30192, ZN => n4436);
   U26179 : XOR2_X1 port map( A1 => n27152, A2 => n34023, Z => n27360);
   U26180 : XOR2_X1 port map( A1 => n9585, A2 => n24532, Z => n34023);
   U26181 : XOR2_X1 port map( A1 => n8637, A2 => n8504, Z => n34024);
   U26184 : AOI21_X1 port map( A1 => n32414, A2 => n25999, B => n18983, ZN => 
                           n5477);
   U26188 : XOR2_X1 port map( A1 => n9006, A2 => n479, Z => n9005);
   U26189 : XOR2_X1 port map( A1 => n29709, A2 => n23119, Z => n22969);
   U26197 : OAI21_X2 port map( A1 => n32037, A2 => n32858, B => n2002, ZN => 
                           n22822);
   U26203 : NAND2_X2 port map( A1 => n34025, A2 => n26682, ZN => n13063);
   U26204 : NAND2_X1 port map( A1 => n12439, A2 => n6657, ZN => n34025);
   U26206 : AOI22_X2 port map( A1 => n30769, A2 => n1013, B1 => n32252, B2 => 
                           n27635, ZN => n34026);
   U26209 : AOI22_X2 port map( A1 => n20278, A2 => n20562, B1 => n20280, B2 => 
                           n15213, ZN => n17633);
   U26210 : XOR2_X1 port map( A1 => n5253, A2 => n12011, Z => n5256);
   U26212 : NAND2_X2 port map( A1 => n10812, A2 => n9374, ZN => n11064);
   U26216 : OAI21_X2 port map( A1 => n34028, A2 => n34027, B => n28923, ZN => 
                           n17680);
   U26217 : NOR2_X1 port map( A1 => n21604, A2 => n33810, ZN => n34027);
   U26218 : XOR2_X1 port map( A1 => n34029, A2 => n29007, Z => n5187);
   U26219 : XOR2_X1 port map( A1 => n19611, A2 => n5190, Z => n34029);
   U26223 : NAND2_X2 port map( A1 => n27440, A2 => n13621, ZN => n29321);
   U26224 : INV_X2 port map( I => n34031, ZN => n29398);
   U26232 : AOI21_X2 port map( A1 => n24285, A2 => n794, B => n24041, ZN => 
                           n13551);
   U26233 : NAND2_X2 port map( A1 => n26389, A2 => n1475, ZN => n7574);
   U26234 : XOR2_X1 port map( A1 => n20781, A2 => n20985, Z => n7452);
   U26237 : NAND2_X2 port map( A1 => n20287, A2 => n27478, ZN => n20985);
   U26239 : NOR2_X1 port map( A1 => n6831, A2 => n25129, ZN => n6830);
   U26242 : NOR2_X2 port map( A1 => n10699, A2 => n11499, ZN => n17822);
   U26245 : NAND2_X2 port map( A1 => n34033, A2 => n16827, ZN => n25542);
   U26246 : XOR2_X1 port map( A1 => n7828, A2 => n34034, Z => n29000);
   U26257 : INV_X1 port map( I => n24843, ZN => n34034);
   U26260 : NAND3_X2 port map( A1 => n13205, A2 => n13204, A3 => n32016, ZN => 
                           n24843);
   U26263 : XNOR2_X1 port map( A1 => n7045, A2 => n7046, ZN => n23344);
   U26264 : NOR2_X2 port map( A1 => n3200, A2 => n4609, ZN => n7046);
   U26266 : NAND3_X1 port map( A1 => n767, A2 => n24340, A3 => n24163, ZN => 
                           n11331);
   U26270 : OAI21_X2 port map( A1 => n20283, A2 => n20282, B => n20281, ZN => 
                           n20781);
   U26271 : XOR2_X1 port map( A1 => n34038, A2 => n21048, Z => n14340);
   U26273 : INV_X2 port map( I => n9852, ZN => n19996);
   U26280 : OAI22_X2 port map( A1 => n13816, A2 => n21840, B1 => n16386, B2 => 
                           n30346, ZN => n21748);
   U26282 : NAND2_X2 port map( A1 => n21497, A2 => n21499, ZN => n21840);
   U26286 : XOR2_X1 port map( A1 => n15791, A2 => n14110, Z => n34085);
   U26290 : NOR3_X1 port map( A1 => n7935, A2 => n10513, A3 => n30651, ZN => 
                           n16408);
   U26296 : NAND2_X2 port map( A1 => n11033, A2 => n11031, ZN => n30584);
   U26298 : XOR2_X1 port map( A1 => n10585, A2 => n32047, Z => n27717);
   U26299 : NAND2_X2 port map( A1 => n13199, A2 => n15677, ZN => n22055);
   U26301 : INV_X2 port map( I => n3581, ZN => n6882);
   U26307 : NAND2_X1 port map( A1 => n34039, A2 => n3581, ZN => n31127);
   U26308 : XOR2_X1 port map( A1 => n29260, A2 => n3584, Z => n3581);
   U26309 : NAND3_X2 port map( A1 => n21882, A2 => n21883, A3 => n12019, ZN => 
                           n22737);
   U26310 : NAND2_X2 port map( A1 => n9646, A2 => n19325, ZN => n13913);
   U26311 : XOR2_X1 port map( A1 => n34041, A2 => n30881, Z => Ciphertext(20));
   U26315 : AOI22_X1 port map( A1 => n12203, A2 => n1208, B1 => n12201, B2 => 
                           n12202, ZN => n34041);
   U26316 : XOR2_X1 port map( A1 => n6020, A2 => n34042, Z => n11986);
   U26317 : XOR2_X1 port map( A1 => n6018, A2 => n31253, Z => n34042);
   U26322 : XOR2_X1 port map( A1 => n5067, A2 => n5068, Z => n5070);
   U26323 : NAND2_X2 port map( A1 => n1773, A2 => n15260, ZN => n9411);
   U26325 : NOR2_X2 port map( A1 => n3446, A2 => n3445, ZN => n34044);
   U26327 : AOI21_X1 port map( A1 => n3650, A2 => n33345, B => n33216, ZN => 
                           n3667);
   U26331 : XOR2_X1 port map( A1 => n14742, A2 => n19722, Z => n10024);
   U26332 : XOR2_X1 port map( A1 => n5127, A2 => n1368, Z => n14742);
   U26333 : NAND2_X1 port map( A1 => n4908, A2 => n5696, ZN => n22913);
   U26336 : XOR2_X1 port map( A1 => Plaintext(157), A2 => Key(157), Z => n16614
                           );
   U26342 : INV_X2 port map( I => n10354, ZN => n34048);
   U26348 : NAND2_X2 port map( A1 => n639, A2 => n34048, ZN => n29395);
   U26353 : NAND3_X2 port map( A1 => n34049, A2 => n26176, A3 => n18341, ZN => 
                           n10423);
   U26360 : NAND2_X2 port map( A1 => n18185, A2 => n16426, ZN => n34049);
   U26361 : XOR2_X1 port map( A1 => n29589, A2 => n6545, Z => n30807);
   U26363 : XOR2_X1 port map( A1 => n31491, A2 => n12310, Z => n30733);
   U26364 : NAND2_X2 port map( A1 => n6110, A2 => n4100, ZN => n34053);
   U26367 : XOR2_X1 port map( A1 => n20727, A2 => n32162, Z => n10164);
   U26369 : XOR2_X1 port map( A1 => n6388, A2 => n6572, Z => n13361);
   U26370 : NAND2_X2 port map( A1 => n30846, A2 => n6619, ZN => n6771);
   U26371 : NAND2_X2 port map( A1 => n34055, A2 => n14561, ZN => n16222);
   U26372 : NAND3_X2 port map( A1 => n7205, A2 => n14560, A3 => n7830, ZN => 
                           n34055);
   U26376 : BUF_X2 port map( I => n11193, Z => n34056);
   U26379 : BUF_X2 port map( I => n16293, Z => n34057);
   U26383 : NOR2_X2 port map( A1 => n26387, A2 => n4151, ZN => n11049);
   U26386 : NOR2_X2 port map( A1 => n847, A2 => n23721, ZN => n28306);
   U26387 : INV_X2 port map( I => n13361, ZN => n847);
   U26393 : NOR2_X2 port map( A1 => n23929, A2 => n23928, ZN => n4897);
   U26396 : NOR3_X2 port map( A1 => n4197, A2 => n11812, A3 => n847, ZN => 
                           n23929);
   U26397 : NAND2_X2 port map( A1 => n1601, A2 => n1600, ZN => n27189);
   U26398 : NOR2_X2 port map( A1 => n31245, A2 => n4531, ZN => n1601);
   U26402 : XOR2_X1 port map( A1 => n30273, A2 => n30487, Z => n30486);
   U26407 : XOR2_X1 port map( A1 => n16829, A2 => n34060, Z => n23925);
   U26408 : XOR2_X1 port map( A1 => n14733, A2 => n29194, Z => n34060);
   U26409 : XOR2_X1 port map( A1 => n22240, A2 => n22210, Z => n21985);
   U26410 : XOR2_X1 port map( A1 => n23261, A2 => n551, Z => n5737);
   U26422 : XOR2_X1 port map( A1 => n24579, A2 => n34061, Z => n31132);
   U26427 : XOR2_X1 port map( A1 => n11370, A2 => n7574, Z => n34061);
   U26429 : NOR2_X1 port map( A1 => n3646, A2 => n5466, ZN => n25251);
   U26432 : XOR2_X1 port map( A1 => n19552, A2 => n31908, Z => n34062);
   U26433 : NAND2_X2 port map( A1 => n5995, A2 => n5996, ZN => n5994);
   U26436 : XOR2_X1 port map( A1 => n34063, A2 => n22141, Z => n30449);
   U26437 : NAND2_X1 port map( A1 => n16034, A2 => n1017, ZN => n34064);
   U26439 : NAND2_X2 port map( A1 => n34065, A2 => n10829, ZN => n16801);
   U26445 : NOR2_X2 port map( A1 => n16393, A2 => n18515, ZN => n34066);
   U26448 : XOR2_X1 port map( A1 => n23143, A2 => n23273, Z => n4554);
   U26453 : XOR2_X1 port map( A1 => n20674, A2 => n20841, Z => n17738);
   U26455 : XOR2_X1 port map( A1 => n21037, A2 => n20892, Z => n20841);
   U26463 : XOR2_X1 port map( A1 => n4567, A2 => n4566, Z => n34067);
   U26465 : NAND2_X2 port map( A1 => n22382, A2 => n17357, ZN => n15421);
   U26474 : INV_X4 port map( I => n8087, ZN => n13920);
   U26476 : NAND2_X2 port map( A1 => n34068, A2 => n26336, ZN => n23536);
   U26477 : NAND2_X1 port map( A1 => n2031, A2 => n2032, ZN => n34068);
   U26478 : OAI21_X2 port map( A1 => n18821, A2 => n12976, B => n16352, ZN => 
                           n12975);
   U26481 : XOR2_X1 port map( A1 => n34070, A2 => n16530, Z => Ciphertext(166))
                           ;
   U26482 : XOR2_X1 port map( A1 => n11726, A2 => n19754, Z => n34071);
   U26485 : OR2_X1 port map( A1 => n16855, A2 => n6634, Z => n6659);
   U26487 : NOR2_X1 port map( A1 => n31783, A2 => n11985, ZN => n7655);
   U26488 : INV_X2 port map( I => n11548, ZN => n31783);
   U26489 : XOR2_X1 port map( A1 => n24754, A2 => n34072, Z => n24536);
   U26501 : XOR2_X1 port map( A1 => n242, A2 => n27750, Z => n34072);
   U26507 : XOR2_X1 port map( A1 => n34073, A2 => n24369, Z => n9125);
   U26510 : INV_X2 port map( I => n981, ZN => n15732);
   U26511 : XOR2_X1 port map( A1 => n19391, A2 => n34076, Z => n29653);
   U26518 : XOR2_X1 port map( A1 => n207, A2 => n34077, Z => n34076);
   U26519 : INV_X2 port map( I => n19769, ZN => n34077);
   U26520 : XOR2_X1 port map( A1 => n26351, A2 => n22145, Z => n22202);
   U26523 : NAND3_X2 port map( A1 => n17941, A2 => n17940, A3 => n5913, ZN => 
                           n34079);
   U26524 : XOR2_X1 port map( A1 => n18028, A2 => n12797, Z => n4332);
   U26525 : AOI21_X2 port map( A1 => n18268, A2 => n19147, B => n18267, ZN => 
                           n19368);
   U26527 : XOR2_X1 port map( A1 => n5737, A2 => n29807, Z => n26170);
   U26528 : NAND2_X2 port map( A1 => n26326, A2 => n2239, ZN => n21497);
   U26531 : XOR2_X1 port map( A1 => n9327, A2 => n29540, Z => n5563);
   U26532 : XOR2_X1 port map( A1 => n34085, A2 => n27851, Z => n15235);
   U26533 : OR2_X1 port map( A1 => n21862, A2 => n13652, Z => n13653);
   U26536 : NAND2_X2 port map( A1 => n21738, A2 => n21866, ZN => n21862);
   U26537 : AOI21_X2 port map( A1 => n21361, A2 => n15728, B => n4906, ZN => 
                           n29302);
   U26538 : XOR2_X1 port map( A1 => n34086, A2 => n24435, Z => Ciphertext(159))
                           ;
   U26539 : NOR2_X1 port map( A1 => n24433, A2 => n24434, ZN => n34086);
   U26540 : INV_X2 port map( I => n2132, ZN => n13966);
   U26541 : NAND2_X1 port map( A1 => n34162, A2 => n13862, ZN => n2132);
   U26542 : XOR2_X1 port map( A1 => n17040, A2 => n23121, Z => n3081);
   U26549 : XOR2_X1 port map( A1 => n23306, A2 => n23420, Z => n23121);
   U26551 : OAI21_X2 port map( A1 => n14767, A2 => n14768, B => n8325, ZN => 
                           n20961);
   U26555 : INV_X2 port map( I => n17426, ZN => n24212);
   U26556 : OAI22_X2 port map( A1 => n14746, A2 => n23651, B1 => n8330, B2 => 
                           n23650, ZN => n17426);
   U26557 : BUF_X2 port map( I => n14236, Z => n34087);
   U26560 : XOR2_X1 port map( A1 => n11867, A2 => n27144, Z => n19684);
   U26563 : XOR2_X1 port map( A1 => n335, A2 => n14685, Z => n22638);
   U26565 : XOR2_X1 port map( A1 => n6607, A2 => n6608, Z => n10675);
   U26566 : NOR2_X2 port map( A1 => n29359, A2 => n5825, ZN => n7776);
   U26569 : XOR2_X1 port map( A1 => n11297, A2 => n25001, Z => n34088);
   U26570 : NAND2_X2 port map( A1 => n8418, A2 => n13231, ZN => n23367);
   U26574 : NOR2_X2 port map( A1 => n25968, A2 => n8787, ZN => n13806);
   U26577 : NOR2_X2 port map( A1 => n26432, A2 => n12247, ZN => n34090);
   U26578 : XOR2_X1 port map( A1 => n24854, A2 => n27423, Z => n26435);
   U26581 : XOR2_X1 port map( A1 => n24377, A2 => n34091, Z => n10901);
   U26582 : XOR2_X1 port map( A1 => n24559, A2 => n27750, Z => n34091);
   U26584 : NAND2_X2 port map( A1 => n28699, A2 => n34092, ZN => n7811);
   U26585 : AOI22_X2 port map( A1 => n1889, A2 => n17341, B1 => n5039, B2 => 
                           n18218, ZN => n34092);
   U26589 : OR2_X1 port map( A1 => n16042, A2 => n14156, Z => n3344);
   U26593 : AOI21_X2 port map( A1 => n2324, A2 => n26976, B => n34093, ZN => 
                           n16693);
   U26595 : BUF_X2 port map( I => n25665, Z => n34094);
   U26596 : XOR2_X1 port map( A1 => n23465, A2 => n34095, Z => n4312);
   U26597 : XOR2_X1 port map( A1 => n23488, A2 => n16548, Z => n34095);
   U26598 : NAND2_X2 port map( A1 => n3489, A2 => n2536, ZN => n5410);
   U26600 : AND2_X1 port map( A1 => n13525, A2 => n4916, Z => n29736);
   U26601 : OR2_X1 port map( A1 => n6286, A2 => n8178, Z => n2245);
   U26602 : AOI22_X2 port map( A1 => n5387, A2 => n25893, B1 => n16113, B2 => 
                           n28910, ZN => n29521);
   U26604 : NAND2_X2 port map( A1 => n19866, A2 => n17177, ZN => n20692);
   U26605 : OAI21_X2 port map( A1 => n3656, A2 => n32499, B => n34102, ZN => 
                           n10824);
   U26606 : NOR2_X2 port map( A1 => n26913, A2 => n27836, ZN => n34102);
   U26609 : NOR2_X2 port map( A1 => n18510, A2 => n34110, ZN => n15789);
   U26610 : INV_X2 port map( I => n18820, ZN => n34110);
   U26611 : XOR2_X1 port map( A1 => n18393, A2 => Key(120), Z => n18820);
   U26614 : XOR2_X1 port map( A1 => n19764, A2 => n18453, Z => n19620);
   U26615 : NAND2_X2 port map( A1 => n17997, A2 => n17996, ZN => n18453);
   U26618 : XNOR2_X1 port map( A1 => n15419, A2 => n6867, ZN => n12008);
   U26629 : XOR2_X1 port map( A1 => n27349, A2 => n23274, Z => n34112);
   U26630 : NAND3_X1 port map( A1 => n27336, A2 => n26445, A3 => n31458, ZN => 
                           n21564);
   U26633 : NAND2_X2 port map( A1 => n1687, A2 => n1688, ZN => n27336);
   U26634 : NAND2_X2 port map( A1 => n34114, A2 => n15069, ZN => n16209);
   U26635 : OR2_X1 port map( A1 => n15071, A2 => n34139, Z => n34114);
   U26641 : XOR2_X1 port map( A1 => n8741, A2 => n19484, Z => n19518);
   U26643 : OAI21_X2 port map( A1 => n18459, A2 => n6597, B => n956, ZN => 
                           n11519);
   U26650 : OR3_X1 port map( A1 => n25236, A2 => n8219, A3 => n34115, Z => 
                           n16398);
   U26651 : XOR2_X1 port map( A1 => n24489, A2 => n10474, Z => n10473);
   U26652 : AOI21_X2 port map( A1 => n2743, A2 => n12448, B => n34116, ZN => 
                           n21992);
   U26656 : XOR2_X1 port map( A1 => n34117, A2 => n25815, Z => Ciphertext(171))
                           ;
   U26663 : NAND2_X1 port map( A1 => n25813, A2 => n25814, ZN => n34117);
   U26668 : XOR2_X1 port map( A1 => n11349, A2 => n7717, Z => n2592);
   U26670 : XOR2_X1 port map( A1 => n24407, A2 => n30986, Z => n24408);
   U26671 : BUF_X2 port map( I => n16073, Z => n34120);
   U26672 : INV_X2 port map( I => n34122, ZN => n12895);
   U26674 : XOR2_X1 port map( A1 => n9914, A2 => n3683, Z => n6948);
   U26675 : OR2_X1 port map( A1 => n7345, A2 => n19057, Z => n16832);
   U26676 : INV_X2 port map( I => n34123, ZN => n34169);
   U26678 : XOR2_X1 port map( A1 => n8896, A2 => n8894, Z => n34123);
   U26679 : XOR2_X1 port map( A1 => n34124, A2 => n23411, Z => n7711);
   U26685 : XOR2_X1 port map( A1 => n23412, A2 => n32893, Z => n34124);
   U26687 : NAND2_X1 port map( A1 => n34125, A2 => n31692, ZN => n9271);
   U26693 : XOR2_X1 port map( A1 => n10184, A2 => n31100, Z => n31692);
   U26696 : XOR2_X1 port map( A1 => n17323, A2 => n15044, Z => n34126);
   U26697 : OAI21_X2 port map( A1 => n27520, A2 => n5089, B => n24655, ZN => 
                           n30323);
   U26698 : NOR2_X2 port map( A1 => n12511, A2 => n15852, ZN => n34127);
   U26699 : XOR2_X1 port map( A1 => n236, A2 => n34129, Z => n2312);
   U26700 : XOR2_X1 port map( A1 => n23408, A2 => n32027, Z => n34129);
   U26701 : OR2_X1 port map( A1 => n29139, A2 => n27485, Z => n23793);
   U26702 : NAND2_X2 port map( A1 => n2687, A2 => n34130, ZN => n11266);
   U26703 : XOR2_X1 port map( A1 => n34133, A2 => n17793, Z => n7987);
   U26704 : XOR2_X1 port map( A1 => n32111, A2 => n16708, Z => n34133);
   U26705 : XOR2_X1 port map( A1 => n26214, A2 => n6395, Z => n27933);
   U26706 : NOR2_X1 port map( A1 => n8678, A2 => n32874, ZN => n25789);
   U26707 : NOR2_X2 port map( A1 => n15709, A2 => n15276, ZN => n8678);
   U26708 : INV_X2 port map( I => n34134, ZN => n13147);
   U26709 : INV_X2 port map( I => n6549, ZN => n16811);
   U26710 : XOR2_X1 port map( A1 => n34135, A2 => n8532, Z => n6549);
   U26711 : OAI21_X2 port map( A1 => n31461, A2 => n24195, B => n34136, ZN => 
                           n1857);
   U26712 : AOI22_X2 port map( A1 => n1315, A2 => n11981, B1 => n4331, B2 => 
                           n21700, ZN => n34138);
   U26713 : INV_X1 port map( I => n18295, ZN => n30934);
   U26714 : XOR2_X1 port map( A1 => Plaintext(84), A2 => Key(84), Z => n18295);
   U26715 : INV_X2 port map( I => n15194, ZN => n34139);
   U26716 : XOR2_X1 port map( A1 => n20928, A2 => n15877, Z => n20753);
   U26717 : AOI21_X2 port map( A1 => n20557, A2 => n20556, B => n15749, ZN => 
                           n20928);
   U26718 : AOI22_X2 port map( A1 => n21624, A2 => n17748, B1 => n21623, B2 => 
                           n28387, ZN => n7477);
   U26719 : BUF_X2 port map( I => n12074, Z => n34140);
   U26720 : BUF_X2 port map( I => n18801, Z => n34141);
   U26721 : AOI22_X2 port map( A1 => n34142, A2 => n28056, B1 => n18739, B2 => 
                           n16287, ZN => n8203);
   U26722 : NOR2_X1 port map( A1 => n18587, A2 => n18737, ZN => n34142);
   U26723 : XOR2_X1 port map( A1 => n23419, A2 => n27186, Z => n23422);
   U26724 : NAND2_X2 port map( A1 => n4776, A2 => n4778, ZN => n27186);
   U26725 : XOR2_X1 port map( A1 => n19556, A2 => n4992, Z => n5607);
   U26726 : OAI21_X2 port map( A1 => n13656, A2 => n13655, B => n34143, ZN => 
                           n10806);
   U26727 : NAND2_X2 port map( A1 => n9508, A2 => n9512, ZN => n4405);
   U26728 : XOR2_X1 port map( A1 => n15028, A2 => n9434, Z => n9586);
   U26729 : NAND2_X2 port map( A1 => n8829, A2 => n8828, ZN => n9434);
   U26730 : XOR2_X1 port map( A1 => n10111, A2 => n12414, Z => n29140);
   U26731 : NAND2_X2 port map( A1 => n4520, A2 => n4519, ZN => n10111);
   U26732 : INV_X2 port map( I => n34144, ZN => n9663);
   U26733 : XOR2_X1 port map( A1 => n10437, A2 => n10436, Z => n34144);
   U26734 : XOR2_X1 port map( A1 => n34145, A2 => n24619, Z => n8845);
   U26735 : XOR2_X1 port map( A1 => n24747, A2 => n31866, Z => n34145);
   U26736 : NAND2_X1 port map( A1 => n28414, A2 => n31533, ZN => n31112);
   U26737 : AND2_X1 port map( A1 => n651, A2 => n16333, Z => n10619);
   U26738 : NAND3_X2 port map( A1 => n8003, A2 => n8005, A3 => n24030, ZN => 
                           n10084);
   U26739 : XOR2_X1 port map( A1 => n1884, A2 => n31626, Z => n8059);
   U26740 : OAI22_X2 port map( A1 => n8653, A2 => n31260, B1 => n8651, B2 => 
                           n16157, ZN => n29693);
   U26741 : XOR2_X1 port map( A1 => n19543, A2 => n19542, Z => n34146);
   U26742 : XOR2_X1 port map( A1 => n21903, A2 => n21911, Z => n14506);
   U26743 : XOR2_X1 port map( A1 => n1305, A2 => n22291, Z => n21911);
   U26744 : XOR2_X1 port map( A1 => n9907, A2 => n24636, Z => n24521);
   U26745 : OAI21_X2 port map( A1 => n18179, A2 => n34147, B => n11461, ZN => 
                           n24826);
   U26746 : OAI22_X2 port map( A1 => n24183, A2 => n28691, B1 => n10381, B2 => 
                           n24052, ZN => n34147);
   U26747 : OR2_X1 port map( A1 => n14080, A2 => n10217, Z => n28507);
   U26748 : BUF_X2 port map( I => n25889, Z => n34149);
   U26749 : XOR2_X1 port map( A1 => n22222, A2 => n8324, Z => n17889);
   U26750 : XOR2_X1 port map( A1 => n26931, A2 => n22147, Z => n22222);
   U26751 : XNOR2_X1 port map( A1 => n3511, A2 => n27599, ZN => n34151);
   U26752 : INV_X2 port map( I => n14456, ZN => n31017);
   U26753 : NOR2_X1 port map( A1 => n29213, A2 => n5837, ZN => n34152);
   U26754 : INV_X2 port map( I => n27110, ZN => n20037);
   U26755 : INV_X2 port map( I => n12670, ZN => n17767);
   U26756 : INV_X4 port map( I => n8530, ZN => n21865);
   U26757 : NAND2_X2 port map( A1 => n8490, A2 => n31965, ZN => n21506);
   U26758 : INV_X2 port map( I => n4274, ZN => n8539);
   U26759 : AND2_X2 port map( A1 => n30984, A2 => n31026, Z => n34160);
   U26760 : INV_X2 port map( I => n11805, ZN => n22397);
   U26761 : XOR2_X1 port map( A1 => n14753, A2 => n11327, Z => n34161);
   U26762 : XNOR2_X1 port map( A1 => n6055, A2 => n28872, ZN => n34162);
   U26763 : BUF_X2 port map( I => n22598, Z => n16432);
   U26764 : INV_X2 port map( I => n8365, ZN => n10295);
   U26765 : INV_X2 port map( I => n6093, ZN => n28825);
   U26766 : NOR2_X2 port map( A1 => n9041, A2 => n9042, ZN => n30321);
   U26767 : INV_X2 port map( I => n17932, ZN => n23786);
   U26768 : AND2_X1 port map( A1 => n32309, A2 => n23894, Z => n34166);
   U26769 : AND3_X1 port map( A1 => n8694, A2 => n14078, A3 => n6474, Z => 
                           n34168);
   U26770 : INV_X4 port map( I => n2967, ZN => n11899);
   U26771 : AND2_X1 port map( A1 => n24958, A2 => n24939, Z => n34170);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_SPEEDY_Top.all;

entity SPEEDY_Top is

   port( clk : in std_logic;  Plaintext, Key : in std_logic_vector (191 downto 
         0);  Ciphertext : out std_logic_vector (191 downto 0));

end SPEEDY_Top;

architecture SYN_Behavioral of SPEEDY_Top is

   component DFFRNQ_X1
      port( D, CLK, RN : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFSNQ_X1
      port( D, CLK, SN : in std_logic;  Q : out std_logic);
   end component;
   
   component SPEEDY_Rounds6_0
      port( Plaintext, Key : in std_logic_vector (191 downto 0);  Ciphertext : 
            out std_logic_vector (191 downto 0));
   end component;
   
   signal reg_in_191_port, reg_in_190_port, reg_in_189_port, reg_in_188_port, 
      reg_in_187_port, reg_in_186_port, reg_in_185_port, reg_in_184_port, 
      reg_in_183_port, reg_in_182_port, reg_in_181_port, reg_in_180_port, 
      reg_in_179_port, reg_in_178_port, reg_in_177_port, reg_in_176_port, 
      reg_in_175_port, reg_in_174_port, reg_in_173_port, reg_in_172_port, 
      reg_in_171_port, reg_in_170_port, reg_in_169_port, reg_in_168_port, 
      reg_in_167_port, reg_in_166_port, reg_in_165_port, reg_in_164_port, 
      reg_in_163_port, reg_in_162_port, reg_in_161_port, reg_in_160_port, 
      reg_in_159_port, reg_in_158_port, reg_in_157_port, reg_in_156_port, 
      reg_in_155_port, reg_in_154_port, reg_in_153_port, reg_in_152_port, 
      reg_in_151_port, reg_in_150_port, reg_in_149_port, reg_in_148_port, 
      reg_in_147_port, reg_in_146_port, reg_in_145_port, reg_in_144_port, 
      reg_in_143_port, reg_in_142_port, reg_in_141_port, reg_in_140_port, 
      reg_in_139_port, reg_in_138_port, reg_in_137_port, reg_in_136_port, 
      reg_in_135_port, reg_in_134_port, reg_in_133_port, reg_in_132_port, 
      reg_in_131_port, reg_in_130_port, reg_in_129_port, reg_in_128_port, 
      reg_in_127_port, reg_in_126_port, reg_in_125_port, reg_in_124_port, 
      reg_in_123_port, reg_in_122_port, reg_in_121_port, reg_in_120_port, 
      reg_in_119_port, reg_in_118_port, reg_in_117_port, reg_in_116_port, 
      reg_in_115_port, reg_in_114_port, reg_in_113_port, reg_in_112_port, 
      reg_in_111_port, reg_in_110_port, reg_in_109_port, reg_in_108_port, 
      reg_in_107_port, reg_in_106_port, reg_in_105_port, reg_in_104_port, 
      reg_in_103_port, reg_in_102_port, reg_in_101_port, reg_in_100_port, 
      reg_in_99_port, reg_in_98_port, reg_in_97_port, reg_in_96_port, 
      reg_in_95_port, reg_in_94_port, reg_in_93_port, reg_in_92_port, 
      reg_in_91_port, reg_in_90_port, reg_in_89_port, reg_in_88_port, 
      reg_in_87_port, reg_in_86_port, reg_in_85_port, reg_in_84_port, 
      reg_in_83_port, reg_in_82_port, reg_in_81_port, reg_in_80_port, 
      reg_in_79_port, reg_in_78_port, reg_in_77_port, reg_in_76_port, 
      reg_in_75_port, reg_in_74_port, reg_in_73_port, reg_in_72_port, 
      reg_in_71_port, reg_in_70_port, reg_in_69_port, reg_in_68_port, 
      reg_in_67_port, reg_in_66_port, reg_in_65_port, reg_in_64_port, 
      reg_in_63_port, reg_in_62_port, reg_in_61_port, reg_in_60_port, 
      reg_in_59_port, reg_in_58_port, reg_in_57_port, reg_in_56_port, 
      reg_in_55_port, reg_in_54_port, reg_in_53_port, reg_in_52_port, 
      reg_in_51_port, reg_in_50_port, reg_in_49_port, reg_in_48_port, 
      reg_in_47_port, reg_in_46_port, reg_in_45_port, reg_in_44_port, 
      reg_in_43_port, reg_in_42_port, reg_in_41_port, reg_in_40_port, 
      reg_in_39_port, reg_in_38_port, reg_in_37_port, reg_in_36_port, 
      reg_in_35_port, reg_in_34_port, reg_in_33_port, reg_in_32_port, 
      reg_in_31_port, reg_in_30_port, reg_in_29_port, reg_in_28_port, 
      reg_in_27_port, reg_in_26_port, reg_in_25_port, reg_in_24_port, 
      reg_in_23_port, reg_in_22_port, reg_in_21_port, reg_in_20_port, 
      reg_in_19_port, reg_in_18_port, reg_in_17_port, reg_in_16_port, 
      reg_in_15_port, reg_in_14_port, reg_in_13_port, reg_in_12_port, 
      reg_in_11_port, reg_in_10_port, reg_in_9_port, reg_in_8_port, 
      reg_in_7_port, reg_in_6_port, reg_in_5_port, reg_in_4_port, reg_in_3_port
      , reg_in_2_port, reg_in_1_port, reg_in_0_port, reg_key_191_port, 
      reg_key_190_port, reg_key_189_port, reg_key_188_port, reg_key_187_port, 
      reg_key_186_port, reg_key_185_port, reg_key_184_port, reg_key_183_port, 
      reg_key_182_port, reg_key_181_port, reg_key_180_port, reg_key_179_port, 
      reg_key_178_port, reg_key_177_port, reg_key_176_port, reg_key_175_port, 
      reg_key_174_port, reg_key_173_port, reg_key_172_port, reg_key_171_port, 
      reg_key_170_port, reg_key_169_port, reg_key_168_port, reg_key_167_port, 
      reg_key_166_port, reg_key_165_port, reg_key_164_port, reg_key_163_port, 
      reg_key_162_port, reg_key_161_port, reg_key_160_port, reg_key_159_port, 
      reg_key_158_port, reg_key_157_port, reg_key_156_port, reg_key_155_port, 
      reg_key_154_port, reg_key_153_port, reg_key_152_port, reg_key_151_port, 
      reg_key_150_port, reg_key_149_port, reg_key_148_port, reg_key_147_port, 
      reg_key_146_port, reg_key_145_port, reg_key_144_port, reg_key_143_port, 
      reg_key_142_port, reg_key_141_port, reg_key_140_port, reg_key_139_port, 
      reg_key_138_port, reg_key_137_port, reg_key_136_port, reg_key_135_port, 
      reg_key_134_port, reg_key_133_port, reg_key_132_port, reg_key_131_port, 
      reg_key_130_port, reg_key_129_port, reg_key_128_port, reg_key_127_port, 
      reg_key_126_port, reg_key_125_port, reg_key_124_port, reg_key_123_port, 
      reg_key_122_port, reg_key_121_port, reg_key_120_port, reg_key_119_port, 
      reg_key_118_port, reg_key_117_port, reg_key_116_port, reg_key_115_port, 
      reg_key_114_port, reg_key_113_port, reg_key_112_port, reg_key_111_port, 
      reg_key_110_port, reg_key_109_port, reg_key_108_port, reg_key_107_port, 
      reg_key_106_port, reg_key_105_port, reg_key_104_port, reg_key_103_port, 
      reg_key_102_port, reg_key_101_port, reg_key_100_port, reg_key_99_port, 
      reg_key_98_port, reg_key_97_port, reg_key_96_port, reg_key_95_port, 
      reg_key_94_port, reg_key_93_port, reg_key_92_port, reg_key_91_port, 
      reg_key_90_port, reg_key_89_port, reg_key_88_port, reg_key_87_port, 
      reg_key_86_port, reg_key_85_port, reg_key_84_port, reg_key_83_port, 
      reg_key_82_port, reg_key_81_port, reg_key_80_port, reg_key_79_port, 
      reg_key_78_port, reg_key_77_port, reg_key_76_port, reg_key_75_port, 
      reg_key_74_port, reg_key_73_port, reg_key_72_port, reg_key_71_port, 
      reg_key_70_port, reg_key_69_port, reg_key_68_port, reg_key_67_port, 
      reg_key_66_port, reg_key_65_port, reg_key_64_port, reg_key_63_port, 
      reg_key_62_port, reg_key_61_port, reg_key_60_port, reg_key_59_port, 
      reg_key_58_port, reg_key_57_port, reg_key_56_port, reg_key_55_port, 
      reg_key_54_port, reg_key_53_port, reg_key_52_port, reg_key_51_port, 
      reg_key_50_port, reg_key_49_port, reg_key_48_port, reg_key_47_port, 
      reg_key_46_port, reg_key_45_port, reg_key_44_port, reg_key_43_port, 
      reg_key_42_port, reg_key_41_port, reg_key_40_port, reg_key_39_port, 
      reg_key_38_port, reg_key_37_port, reg_key_36_port, reg_key_35_port, 
      reg_key_34_port, reg_key_33_port, reg_key_32_port, reg_key_31_port, 
      reg_key_30_port, reg_key_29_port, reg_key_28_port, reg_key_27_port, 
      reg_key_26_port, reg_key_25_port, reg_key_24_port, reg_key_23_port, 
      reg_key_22_port, reg_key_21_port, reg_key_20_port, reg_key_19_port, 
      reg_key_18_port, reg_key_17_port, reg_key_16_port, reg_key_15_port, 
      reg_key_14_port, reg_key_13_port, reg_key_12_port, reg_key_11_port, 
      reg_key_10_port, reg_key_9_port, reg_key_8_port, reg_key_7_port, 
      reg_key_6_port, reg_key_5_port, reg_key_4_port, reg_key_3_port, 
      reg_key_2_port, reg_key_1_port, reg_key_0_port, reg_out_191_port, 
      reg_out_190_port, reg_out_189_port, reg_out_188_port, reg_out_187_port, 
      reg_out_186_port, reg_out_185_port, reg_out_184_port, reg_out_183_port, 
      reg_out_182_port, reg_out_181_port, reg_out_180_port, reg_out_179_port, 
      reg_out_178_port, reg_out_177_port, reg_out_176_port, reg_out_175_port, 
      reg_out_174_port, reg_out_173_port, reg_out_172_port, reg_out_171_port, 
      reg_out_170_port, reg_out_169_port, reg_out_168_port, reg_out_167_port, 
      reg_out_166_port, reg_out_165_port, reg_out_164_port, reg_out_163_port, 
      reg_out_162_port, reg_out_161_port, reg_out_160_port, reg_out_159_port, 
      reg_out_158_port, reg_out_157_port, reg_out_156_port, reg_out_155_port, 
      reg_out_154_port, reg_out_153_port, reg_out_152_port, reg_out_151_port, 
      reg_out_150_port, reg_out_149_port, reg_out_148_port, reg_out_147_port, 
      reg_out_146_port, reg_out_145_port, reg_out_144_port, reg_out_143_port, 
      reg_out_142_port, reg_out_141_port, reg_out_140_port, reg_out_139_port, 
      reg_out_138_port, reg_out_137_port, reg_out_136_port, reg_out_135_port, 
      reg_out_134_port, reg_out_133_port, reg_out_132_port, reg_out_131_port, 
      reg_out_130_port, reg_out_129_port, reg_out_128_port, reg_out_127_port, 
      reg_out_126_port, reg_out_125_port, reg_out_124_port, reg_out_123_port, 
      reg_out_122_port, reg_out_121_port, reg_out_120_port, reg_out_119_port, 
      reg_out_118_port, reg_out_117_port, reg_out_116_port, reg_out_115_port, 
      reg_out_114_port, reg_out_113_port, reg_out_112_port, reg_out_111_port, 
      reg_out_110_port, reg_out_109_port, reg_out_108_port, reg_out_107_port, 
      reg_out_106_port, reg_out_105_port, reg_out_104_port, reg_out_103_port, 
      reg_out_102_port, reg_out_101_port, reg_out_100_port, reg_out_99_port, 
      reg_out_98_port, reg_out_97_port, reg_out_96_port, reg_out_95_port, 
      reg_out_94_port, reg_out_93_port, reg_out_92_port, reg_out_91_port, 
      reg_out_90_port, reg_out_89_port, reg_out_88_port, reg_out_87_port, 
      reg_out_86_port, reg_out_85_port, reg_out_84_port, reg_out_83_port, 
      reg_out_82_port, reg_out_81_port, reg_out_80_port, reg_out_79_port, 
      reg_out_78_port, reg_out_77_port, reg_out_76_port, reg_out_75_port, 
      reg_out_74_port, reg_out_73_port, reg_out_72_port, reg_out_71_port, 
      reg_out_70_port, reg_out_69_port, reg_out_68_port, reg_out_67_port, 
      reg_out_66_port, reg_out_65_port, reg_out_64_port, reg_out_63_port, 
      reg_out_62_port, reg_out_61_port, reg_out_60_port, reg_out_59_port, 
      reg_out_58_port, reg_out_57_port, reg_out_56_port, reg_out_55_port, 
      reg_out_54_port, reg_out_53_port, reg_out_52_port, reg_out_51_port, 
      reg_out_50_port, reg_out_49_port, reg_out_48_port, reg_out_47_port, 
      reg_out_46_port, reg_out_45_port, reg_out_44_port, reg_out_43_port, 
      reg_out_42_port, reg_out_41_port, reg_out_40_port, reg_out_39_port, 
      reg_out_38_port, reg_out_37_port, reg_out_36_port, reg_out_35_port, 
      reg_out_34_port, reg_out_33_port, reg_out_32_port, reg_out_31_port, 
      reg_out_30_port, reg_out_29_port, reg_out_28_port, reg_out_27_port, 
      reg_out_26_port, reg_out_25_port, reg_out_24_port, reg_out_23_port, 
      reg_out_22_port, reg_out_21_port, reg_out_20_port, reg_out_19_port, 
      reg_out_18_port, reg_out_17_port, reg_out_16_port, reg_out_15_port, 
      reg_out_14_port, reg_out_13_port, reg_out_12_port, reg_out_11_port, 
      reg_out_10_port, reg_out_9_port, reg_out_8_port, reg_out_7_port, 
      reg_out_6_port, reg_out_5_port, reg_out_4_port, reg_out_3_port, 
      reg_out_2_port, reg_out_1_port, reg_out_0_port, n5, n9, n10, n11, n12, 
      n16, n19, n20, n21, n24, n27, n29, n33, n34, n46, n48, n51, n53, n54, n55
      , n59, n63, n64, n65, n66, n69, n70, n71, n73, n76, n77, n80, n82, n83, 
      n86, n88, n90, n92, n93, n94, n95, n96, n100, n104, n108, n109, n119, 
      n120, n137, n139, n141, n142, n145, n149, n151, n154, n155, n156, n157, 
      n161, n164, n165, n166, n167, n170, n171, n173, n184, n185, n189, n191, 
      n193, n194, n195, n196, n197, n198, n199, n200, n202, n203, n204, n205, 
      n206, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n466, n467, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n497, n498, n499, n500, 
      n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, 
      n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, 
      n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, 
      n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n571, n572, n573, 
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
      n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
      n635, n636, n637, n638, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, 
      n673, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
      n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711 : std_logic;

begin
   
   reg_in_regx191x : DFFSNQ_X1 port map( D => Plaintext(191), CLK => clk, SN =>
                           n576, Q => reg_in_191_port);
   reg_in_regx190x : DFFSNQ_X1 port map( D => Plaintext(190), CLK => clk, SN =>
                           n575, Q => reg_in_190_port);
   reg_in_regx189x : DFFSNQ_X1 port map( D => Plaintext(189), CLK => clk, SN =>
                           n574, Q => reg_in_189_port);
   reg_in_regx188x : DFFSNQ_X1 port map( D => Plaintext(188), CLK => clk, SN =>
                           n573, Q => reg_in_188_port);
   reg_in_regx187x : DFFSNQ_X1 port map( D => Plaintext(187), CLK => clk, SN =>
                           n572, Q => reg_in_187_port);
   reg_in_regx186x : DFFSNQ_X1 port map( D => Plaintext(186), CLK => clk, SN =>
                           n571, Q => reg_in_186_port);
   reg_in_regx184x : DFFSNQ_X1 port map( D => Plaintext(184), CLK => clk, SN =>
                           n569, Q => reg_in_184_port);
   reg_in_regx183x : DFFSNQ_X1 port map( D => Plaintext(183), CLK => clk, SN =>
                           n568, Q => reg_in_183_port);
   reg_in_regx182x : DFFSNQ_X1 port map( D => Plaintext(182), CLK => clk, SN =>
                           n567, Q => reg_in_182_port);
   reg_in_regx181x : DFFSNQ_X1 port map( D => Plaintext(181), CLK => clk, SN =>
                           n566, Q => reg_in_181_port);
   reg_in_regx180x : DFFSNQ_X1 port map( D => Plaintext(180), CLK => clk, SN =>
                           n565, Q => reg_in_180_port);
   reg_in_regx179x : DFFSNQ_X1 port map( D => Plaintext(179), CLK => clk, SN =>
                           n564, Q => reg_in_179_port);
   reg_in_regx178x : DFFSNQ_X1 port map( D => Plaintext(178), CLK => clk, SN =>
                           n563, Q => reg_in_178_port);
   reg_in_regx177x : DFFSNQ_X1 port map( D => Plaintext(177), CLK => clk, SN =>
                           n562, Q => reg_in_177_port);
   reg_in_regx176x : DFFSNQ_X1 port map( D => Plaintext(176), CLK => clk, SN =>
                           n561, Q => reg_in_176_port);
   reg_in_regx175x : DFFSNQ_X1 port map( D => Plaintext(175), CLK => clk, SN =>
                           n560, Q => reg_in_175_port);
   reg_in_regx174x : DFFSNQ_X1 port map( D => Plaintext(174), CLK => clk, SN =>
                           n559, Q => reg_in_174_port);
   reg_in_regx173x : DFFSNQ_X1 port map( D => Plaintext(173), CLK => clk, SN =>
                           n558, Q => reg_in_173_port);
   reg_in_regx172x : DFFSNQ_X1 port map( D => Plaintext(172), CLK => clk, SN =>
                           n557, Q => reg_in_172_port);
   reg_in_regx171x : DFFSNQ_X1 port map( D => Plaintext(171), CLK => clk, SN =>
                           n556, Q => reg_in_171_port);
   reg_in_regx170x : DFFSNQ_X1 port map( D => Plaintext(170), CLK => clk, SN =>
                           n555, Q => reg_in_170_port);
   reg_in_regx169x : DFFSNQ_X1 port map( D => Plaintext(169), CLK => clk, SN =>
                           n554, Q => reg_in_169_port);
   reg_in_regx168x : DFFSNQ_X1 port map( D => Plaintext(168), CLK => clk, SN =>
                           n553, Q => reg_in_168_port);
   reg_in_regx167x : DFFSNQ_X1 port map( D => Plaintext(167), CLK => clk, SN =>
                           n552, Q => reg_in_167_port);
   reg_in_regx166x : DFFSNQ_X1 port map( D => Plaintext(166), CLK => clk, SN =>
                           n551, Q => reg_in_166_port);
   reg_in_regx165x : DFFSNQ_X1 port map( D => Plaintext(165), CLK => clk, SN =>
                           n550, Q => reg_in_165_port);
   reg_in_regx164x : DFFSNQ_X1 port map( D => Plaintext(164), CLK => clk, SN =>
                           n549, Q => reg_in_164_port);
   reg_in_regx163x : DFFSNQ_X1 port map( D => Plaintext(163), CLK => clk, SN =>
                           n548, Q => reg_in_163_port);
   reg_in_regx162x : DFFSNQ_X1 port map( D => Plaintext(162), CLK => clk, SN =>
                           n547, Q => reg_in_162_port);
   reg_in_regx161x : DFFSNQ_X1 port map( D => Plaintext(161), CLK => clk, SN =>
                           n546, Q => reg_in_161_port);
   reg_in_regx160x : DFFSNQ_X1 port map( D => Plaintext(160), CLK => clk, SN =>
                           n545, Q => reg_in_160_port);
   reg_in_regx159x : DFFSNQ_X1 port map( D => Plaintext(159), CLK => clk, SN =>
                           n544, Q => reg_in_159_port);
   reg_in_regx158x : DFFSNQ_X1 port map( D => Plaintext(158), CLK => clk, SN =>
                           n543, Q => reg_in_158_port);
   reg_in_regx157x : DFFSNQ_X1 port map( D => Plaintext(157), CLK => clk, SN =>
                           n542, Q => reg_in_157_port);
   reg_in_regx156x : DFFSNQ_X1 port map( D => Plaintext(156), CLK => clk, SN =>
                           n541, Q => reg_in_156_port);
   reg_in_regx155x : DFFSNQ_X1 port map( D => Plaintext(155), CLK => clk, SN =>
                           n540, Q => reg_in_155_port);
   reg_in_regx154x : DFFSNQ_X1 port map( D => Plaintext(154), CLK => clk, SN =>
                           n539, Q => reg_in_154_port);
   reg_in_regx153x : DFFSNQ_X1 port map( D => Plaintext(153), CLK => clk, SN =>
                           n538, Q => reg_in_153_port);
   reg_in_regx152x : DFFSNQ_X1 port map( D => Plaintext(152), CLK => clk, SN =>
                           n537, Q => reg_in_152_port);
   reg_in_regx151x : DFFSNQ_X1 port map( D => Plaintext(151), CLK => clk, SN =>
                           n536, Q => reg_in_151_port);
   reg_in_regx150x : DFFSNQ_X1 port map( D => Plaintext(150), CLK => clk, SN =>
                           n535, Q => reg_in_150_port);
   reg_in_regx149x : DFFSNQ_X1 port map( D => Plaintext(149), CLK => clk, SN =>
                           n534, Q => reg_in_149_port);
   reg_in_regx148x : DFFSNQ_X1 port map( D => Plaintext(148), CLK => clk, SN =>
                           n533, Q => reg_in_148_port);
   reg_in_regx147x : DFFSNQ_X1 port map( D => Plaintext(147), CLK => clk, SN =>
                           n532, Q => reg_in_147_port);
   reg_in_regx146x : DFFSNQ_X1 port map( D => Plaintext(146), CLK => clk, SN =>
                           n531, Q => reg_in_146_port);
   reg_in_regx145x : DFFSNQ_X1 port map( D => Plaintext(145), CLK => clk, SN =>
                           n530, Q => reg_in_145_port);
   reg_in_regx144x : DFFSNQ_X1 port map( D => Plaintext(144), CLK => clk, SN =>
                           n529, Q => reg_in_144_port);
   reg_in_regx143x : DFFSNQ_X1 port map( D => Plaintext(143), CLK => clk, SN =>
                           n528, Q => reg_in_143_port);
   reg_in_regx142x : DFFSNQ_X1 port map( D => Plaintext(142), CLK => clk, SN =>
                           n527, Q => reg_in_142_port);
   reg_in_regx141x : DFFSNQ_X1 port map( D => Plaintext(141), CLK => clk, SN =>
                           n526, Q => reg_in_141_port);
   reg_in_regx140x : DFFSNQ_X1 port map( D => Plaintext(140), CLK => clk, SN =>
                           n525, Q => reg_in_140_port);
   reg_in_regx139x : DFFSNQ_X1 port map( D => Plaintext(139), CLK => clk, SN =>
                           n524, Q => reg_in_139_port);
   reg_in_regx138x : DFFSNQ_X1 port map( D => Plaintext(138), CLK => clk, SN =>
                           n523, Q => reg_in_138_port);
   reg_in_regx137x : DFFSNQ_X1 port map( D => Plaintext(137), CLK => clk, SN =>
                           n522, Q => reg_in_137_port);
   reg_in_regx136x : DFFSNQ_X1 port map( D => Plaintext(136), CLK => clk, SN =>
                           n521, Q => reg_in_136_port);
   reg_in_regx135x : DFFSNQ_X1 port map( D => Plaintext(135), CLK => clk, SN =>
                           n520, Q => reg_in_135_port);
   reg_in_regx134x : DFFSNQ_X1 port map( D => Plaintext(134), CLK => clk, SN =>
                           n519, Q => reg_in_134_port);
   reg_in_regx133x : DFFSNQ_X1 port map( D => Plaintext(133), CLK => clk, SN =>
                           n518, Q => reg_in_133_port);
   reg_in_regx132x : DFFSNQ_X1 port map( D => Plaintext(132), CLK => clk, SN =>
                           n517, Q => reg_in_132_port);
   reg_in_regx131x : DFFSNQ_X1 port map( D => Plaintext(131), CLK => clk, SN =>
                           n516, Q => reg_in_131_port);
   reg_in_regx130x : DFFSNQ_X1 port map( D => Plaintext(130), CLK => clk, SN =>
                           n515, Q => reg_in_130_port);
   reg_in_regx129x : DFFSNQ_X1 port map( D => Plaintext(129), CLK => clk, SN =>
                           n514, Q => reg_in_129_port);
   reg_in_regx128x : DFFSNQ_X1 port map( D => Plaintext(128), CLK => clk, SN =>
                           n513, Q => reg_in_128_port);
   reg_in_regx127x : DFFSNQ_X1 port map( D => Plaintext(127), CLK => clk, SN =>
                           n512, Q => reg_in_127_port);
   reg_in_regx126x : DFFSNQ_X1 port map( D => Plaintext(126), CLK => clk, SN =>
                           n511, Q => reg_in_126_port);
   reg_in_regx125x : DFFSNQ_X1 port map( D => Plaintext(125), CLK => clk, SN =>
                           n510, Q => reg_in_125_port);
   reg_in_regx124x : DFFSNQ_X1 port map( D => Plaintext(124), CLK => clk, SN =>
                           n509, Q => reg_in_124_port);
   reg_in_regx123x : DFFSNQ_X1 port map( D => Plaintext(123), CLK => clk, SN =>
                           n508, Q => reg_in_123_port);
   reg_in_regx122x : DFFSNQ_X1 port map( D => Plaintext(122), CLK => clk, SN =>
                           n507, Q => reg_in_122_port);
   reg_in_regx121x : DFFSNQ_X1 port map( D => Plaintext(121), CLK => clk, SN =>
                           n506, Q => reg_in_121_port);
   reg_in_regx120x : DFFSNQ_X1 port map( D => Plaintext(120), CLK => clk, SN =>
                           n505, Q => reg_in_120_port);
   reg_in_regx119x : DFFSNQ_X1 port map( D => Plaintext(119), CLK => clk, SN =>
                           n504, Q => reg_in_119_port);
   reg_in_regx118x : DFFSNQ_X1 port map( D => Plaintext(118), CLK => clk, SN =>
                           n503, Q => reg_in_118_port);
   reg_in_regx117x : DFFSNQ_X1 port map( D => Plaintext(117), CLK => clk, SN =>
                           n502, Q => reg_in_117_port);
   reg_in_regx116x : DFFSNQ_X1 port map( D => Plaintext(116), CLK => clk, SN =>
                           n501, Q => reg_in_116_port);
   reg_in_regx115x : DFFSNQ_X1 port map( D => Plaintext(115), CLK => clk, SN =>
                           n500, Q => reg_in_115_port);
   reg_in_regx114x : DFFSNQ_X1 port map( D => Plaintext(114), CLK => clk, SN =>
                           n499, Q => reg_in_114_port);
   reg_in_regx113x : DFFSNQ_X1 port map( D => Plaintext(113), CLK => clk, SN =>
                           n498, Q => reg_in_113_port);
   reg_in_regx112x : DFFSNQ_X1 port map( D => Plaintext(112), CLK => clk, SN =>
                           n497, Q => reg_in_112_port);
   reg_in_regx110x : DFFSNQ_X1 port map( D => Plaintext(110), CLK => clk, SN =>
                           n495, Q => reg_in_110_port);
   reg_in_regx109x : DFFSNQ_X1 port map( D => Plaintext(109), CLK => clk, SN =>
                           n494, Q => reg_in_109_port);
   reg_in_regx108x : DFFSNQ_X1 port map( D => Plaintext(108), CLK => clk, SN =>
                           n493, Q => reg_in_108_port);
   reg_in_regx107x : DFFSNQ_X1 port map( D => Plaintext(107), CLK => clk, SN =>
                           n492, Q => reg_in_107_port);
   reg_in_regx106x : DFFSNQ_X1 port map( D => Plaintext(106), CLK => clk, SN =>
                           n491, Q => reg_in_106_port);
   reg_in_regx105x : DFFSNQ_X1 port map( D => Plaintext(105), CLK => clk, SN =>
                           n490, Q => reg_in_105_port);
   reg_in_regx104x : DFFSNQ_X1 port map( D => Plaintext(104), CLK => clk, SN =>
                           n489, Q => reg_in_104_port);
   reg_in_regx103x : DFFSNQ_X1 port map( D => Plaintext(103), CLK => clk, SN =>
                           n488, Q => reg_in_103_port);
   reg_in_regx102x : DFFSNQ_X1 port map( D => Plaintext(102), CLK => clk, SN =>
                           n487, Q => reg_in_102_port);
   reg_in_regx100x : DFFSNQ_X1 port map( D => Plaintext(100), CLK => clk, SN =>
                           n485, Q => reg_in_100_port);
   reg_in_regx99x : DFFSNQ_X1 port map( D => Plaintext(99), CLK => clk, SN => 
                           n484, Q => reg_in_99_port);
   reg_in_regx98x : DFFSNQ_X1 port map( D => Plaintext(98), CLK => clk, SN => 
                           n483, Q => reg_in_98_port);
   reg_in_regx97x : DFFSNQ_X1 port map( D => Plaintext(97), CLK => clk, SN => 
                           n482, Q => reg_in_97_port);
   reg_in_regx96x : DFFSNQ_X1 port map( D => Plaintext(96), CLK => clk, SN => 
                           n481, Q => reg_in_96_port);
   reg_in_regx95x : DFFSNQ_X1 port map( D => Plaintext(95), CLK => clk, SN => 
                           n480, Q => reg_in_95_port);
   reg_in_regx94x : DFFSNQ_X1 port map( D => Plaintext(94), CLK => clk, SN => 
                           n479, Q => reg_in_94_port);
   reg_in_regx93x : DFFSNQ_X1 port map( D => Plaintext(93), CLK => clk, SN => 
                           n478, Q => reg_in_93_port);
   reg_in_regx92x : DFFSNQ_X1 port map( D => Plaintext(92), CLK => clk, SN => 
                           n477, Q => reg_in_92_port);
   reg_in_regx91x : DFFSNQ_X1 port map( D => Plaintext(91), CLK => clk, SN => 
                           n476, Q => reg_in_91_port);
   reg_in_regx90x : DFFSNQ_X1 port map( D => Plaintext(90), CLK => clk, SN => 
                           n475, Q => reg_in_90_port);
   reg_in_regx89x : DFFSNQ_X1 port map( D => Plaintext(89), CLK => clk, SN => 
                           n474, Q => reg_in_89_port);
   reg_in_regx88x : DFFSNQ_X1 port map( D => Plaintext(88), CLK => clk, SN => 
                           n473, Q => reg_in_88_port);
   reg_in_regx87x : DFFSNQ_X1 port map( D => Plaintext(87), CLK => clk, SN => 
                           n472, Q => reg_in_87_port);
   reg_in_regx86x : DFFSNQ_X1 port map( D => Plaintext(86), CLK => clk, SN => 
                           n471, Q => reg_in_86_port);
   reg_in_regx85x : DFFSNQ_X1 port map( D => Plaintext(85), CLK => clk, SN => 
                           n470, Q => reg_in_85_port);
   reg_in_regx84x : DFFSNQ_X1 port map( D => Plaintext(84), CLK => clk, SN => 
                           n469, Q => reg_in_84_port);
   reg_in_regx82x : DFFSNQ_X1 port map( D => Plaintext(82), CLK => clk, SN => 
                           n467, Q => reg_in_82_port);
   reg_in_regx81x : DFFSNQ_X1 port map( D => Plaintext(81), CLK => clk, SN => 
                           n466, Q => reg_in_81_port);
   reg_in_regx79x : DFFSNQ_X1 port map( D => Plaintext(79), CLK => clk, SN => 
                           n464, Q => reg_in_79_port);
   reg_in_regx78x : DFFSNQ_X1 port map( D => Plaintext(78), CLK => clk, SN => 
                           n463, Q => reg_in_78_port);
   reg_in_regx77x : DFFSNQ_X1 port map( D => Plaintext(77), CLK => clk, SN => 
                           n462, Q => reg_in_77_port);
   reg_in_regx76x : DFFSNQ_X1 port map( D => Plaintext(76), CLK => clk, SN => 
                           n461, Q => reg_in_76_port);
   reg_in_regx75x : DFFSNQ_X1 port map( D => Plaintext(75), CLK => clk, SN => 
                           n460, Q => reg_in_75_port);
   reg_in_regx74x : DFFSNQ_X1 port map( D => Plaintext(74), CLK => clk, SN => 
                           n459, Q => reg_in_74_port);
   reg_in_regx73x : DFFSNQ_X1 port map( D => Plaintext(73), CLK => clk, SN => 
                           n458, Q => reg_in_73_port);
   reg_in_regx72x : DFFSNQ_X1 port map( D => Plaintext(72), CLK => clk, SN => 
                           n457, Q => reg_in_72_port);
   reg_in_regx71x : DFFSNQ_X1 port map( D => Plaintext(71), CLK => clk, SN => 
                           n456, Q => reg_in_71_port);
   reg_in_regx70x : DFFSNQ_X1 port map( D => Plaintext(70), CLK => clk, SN => 
                           n455, Q => reg_in_70_port);
   reg_in_regx69x : DFFSNQ_X1 port map( D => Plaintext(69), CLK => clk, SN => 
                           n454, Q => reg_in_69_port);
   reg_in_regx68x : DFFSNQ_X1 port map( D => Plaintext(68), CLK => clk, SN => 
                           n453, Q => reg_in_68_port);
   reg_in_regx67x : DFFSNQ_X1 port map( D => Plaintext(67), CLK => clk, SN => 
                           n452, Q => reg_in_67_port);
   reg_in_regx66x : DFFSNQ_X1 port map( D => Plaintext(66), CLK => clk, SN => 
                           n451, Q => reg_in_66_port);
   reg_in_regx65x : DFFSNQ_X1 port map( D => Plaintext(65), CLK => clk, SN => 
                           n450, Q => reg_in_65_port);
   reg_in_regx64x : DFFSNQ_X1 port map( D => Plaintext(64), CLK => clk, SN => 
                           n449, Q => reg_in_64_port);
   reg_in_regx63x : DFFSNQ_X1 port map( D => Plaintext(63), CLK => clk, SN => 
                           n448, Q => reg_in_63_port);
   reg_in_regx62x : DFFSNQ_X1 port map( D => Plaintext(62), CLK => clk, SN => 
                           n447, Q => reg_in_62_port);
   reg_in_regx61x : DFFSNQ_X1 port map( D => Plaintext(61), CLK => clk, SN => 
                           n446, Q => reg_in_61_port);
   reg_in_regx60x : DFFSNQ_X1 port map( D => Plaintext(60), CLK => clk, SN => 
                           n445, Q => reg_in_60_port);
   reg_in_regx58x : DFFSNQ_X1 port map( D => Plaintext(58), CLK => clk, SN => 
                           n443, Q => reg_in_58_port);
   reg_in_regx57x : DFFSNQ_X1 port map( D => Plaintext(57), CLK => clk, SN => 
                           n442, Q => reg_in_57_port);
   reg_in_regx56x : DFFSNQ_X1 port map( D => Plaintext(56), CLK => clk, SN => 
                           n441, Q => reg_in_56_port);
   reg_in_regx55x : DFFSNQ_X1 port map( D => Plaintext(55), CLK => clk, SN => 
                           n440, Q => reg_in_55_port);
   reg_in_regx54x : DFFSNQ_X1 port map( D => Plaintext(54), CLK => clk, SN => 
                           n439, Q => reg_in_54_port);
   reg_in_regx53x : DFFSNQ_X1 port map( D => Plaintext(53), CLK => clk, SN => 
                           n438, Q => reg_in_53_port);
   reg_in_regx52x : DFFSNQ_X1 port map( D => Plaintext(52), CLK => clk, SN => 
                           n437, Q => reg_in_52_port);
   reg_in_regx51x : DFFSNQ_X1 port map( D => Plaintext(51), CLK => clk, SN => 
                           n436, Q => reg_in_51_port);
   reg_in_regx50x : DFFSNQ_X1 port map( D => Plaintext(50), CLK => clk, SN => 
                           n435, Q => reg_in_50_port);
   reg_in_regx49x : DFFSNQ_X1 port map( D => Plaintext(49), CLK => clk, SN => 
                           n434, Q => reg_in_49_port);
   reg_in_regx48x : DFFSNQ_X1 port map( D => Plaintext(48), CLK => clk, SN => 
                           n433, Q => reg_in_48_port);
   reg_in_regx47x : DFFSNQ_X1 port map( D => Plaintext(47), CLK => clk, SN => 
                           n432, Q => reg_in_47_port);
   reg_in_regx46x : DFFSNQ_X1 port map( D => Plaintext(46), CLK => clk, SN => 
                           n431, Q => reg_in_46_port);
   reg_in_regx45x : DFFSNQ_X1 port map( D => Plaintext(45), CLK => clk, SN => 
                           n430, Q => reg_in_45_port);
   reg_in_regx44x : DFFSNQ_X1 port map( D => Plaintext(44), CLK => clk, SN => 
                           n429, Q => reg_in_44_port);
   reg_in_regx43x : DFFSNQ_X1 port map( D => Plaintext(43), CLK => clk, SN => 
                           n428, Q => reg_in_43_port);
   reg_in_regx42x : DFFSNQ_X1 port map( D => Plaintext(42), CLK => clk, SN => 
                           n427, Q => reg_in_42_port);
   reg_in_regx41x : DFFSNQ_X1 port map( D => Plaintext(41), CLK => clk, SN => 
                           n426, Q => reg_in_41_port);
   reg_in_regx40x : DFFSNQ_X1 port map( D => Plaintext(40), CLK => clk, SN => 
                           n425, Q => reg_in_40_port);
   reg_in_regx39x : DFFSNQ_X1 port map( D => Plaintext(39), CLK => clk, SN => 
                           n424, Q => reg_in_39_port);
   reg_in_regx38x : DFFSNQ_X1 port map( D => Plaintext(38), CLK => clk, SN => 
                           n423, Q => reg_in_38_port);
   reg_in_regx37x : DFFSNQ_X1 port map( D => Plaintext(37), CLK => clk, SN => 
                           n422, Q => reg_in_37_port);
   reg_in_regx36x : DFFSNQ_X1 port map( D => Plaintext(36), CLK => clk, SN => 
                           n421, Q => reg_in_36_port);
   reg_in_regx35x : DFFSNQ_X1 port map( D => Plaintext(35), CLK => clk, SN => 
                           n420, Q => reg_in_35_port);
   reg_in_regx34x : DFFSNQ_X1 port map( D => Plaintext(34), CLK => clk, SN => 
                           n419, Q => reg_in_34_port);
   reg_in_regx33x : DFFSNQ_X1 port map( D => Plaintext(33), CLK => clk, SN => 
                           n418, Q => reg_in_33_port);
   reg_in_regx32x : DFFSNQ_X1 port map( D => Plaintext(32), CLK => clk, SN => 
                           n417, Q => reg_in_32_port);
   reg_in_regx31x : DFFSNQ_X1 port map( D => Plaintext(31), CLK => clk, SN => 
                           n416, Q => reg_in_31_port);
   reg_in_regx30x : DFFSNQ_X1 port map( D => Plaintext(30), CLK => clk, SN => 
                           n415, Q => reg_in_30_port);
   reg_in_regx29x : DFFSNQ_X1 port map( D => Plaintext(29), CLK => clk, SN => 
                           n414, Q => reg_in_29_port);
   reg_in_regx28x : DFFSNQ_X1 port map( D => Plaintext(28), CLK => clk, SN => 
                           n413, Q => reg_in_28_port);
   reg_in_regx27x : DFFSNQ_X1 port map( D => Plaintext(27), CLK => clk, SN => 
                           n412, Q => reg_in_27_port);
   reg_in_regx26x : DFFSNQ_X1 port map( D => Plaintext(26), CLK => clk, SN => 
                           n411, Q => reg_in_26_port);
   reg_in_regx25x : DFFSNQ_X1 port map( D => Plaintext(25), CLK => clk, SN => 
                           n410, Q => reg_in_25_port);
   reg_in_regx24x : DFFSNQ_X1 port map( D => Plaintext(24), CLK => clk, SN => 
                           n409, Q => reg_in_24_port);
   reg_in_regx23x : DFFSNQ_X1 port map( D => Plaintext(23), CLK => clk, SN => 
                           n408, Q => reg_in_23_port);
   reg_in_regx22x : DFFSNQ_X1 port map( D => Plaintext(22), CLK => clk, SN => 
                           n407, Q => reg_in_22_port);
   reg_in_regx21x : DFFSNQ_X1 port map( D => Plaintext(21), CLK => clk, SN => 
                           n406, Q => reg_in_21_port);
   reg_in_regx20x : DFFSNQ_X1 port map( D => Plaintext(20), CLK => clk, SN => 
                           n405, Q => reg_in_20_port);
   reg_in_regx19x : DFFSNQ_X1 port map( D => Plaintext(19), CLK => clk, SN => 
                           n404, Q => reg_in_19_port);
   reg_in_regx18x : DFFSNQ_X1 port map( D => Plaintext(18), CLK => clk, SN => 
                           n403, Q => reg_in_18_port);
   reg_in_regx17x : DFFSNQ_X1 port map( D => Plaintext(17), CLK => clk, SN => 
                           n402, Q => reg_in_17_port);
   reg_in_regx16x : DFFSNQ_X1 port map( D => Plaintext(16), CLK => clk, SN => 
                           n401, Q => reg_in_16_port);
   reg_in_regx15x : DFFSNQ_X1 port map( D => Plaintext(15), CLK => clk, SN => 
                           n400, Q => reg_in_15_port);
   reg_in_regx14x : DFFSNQ_X1 port map( D => Plaintext(14), CLK => clk, SN => 
                           n399, Q => reg_in_14_port);
   reg_in_regx13x : DFFSNQ_X1 port map( D => Plaintext(13), CLK => clk, SN => 
                           n398, Q => reg_in_13_port);
   reg_in_regx12x : DFFSNQ_X1 port map( D => Plaintext(12), CLK => clk, SN => 
                           n397, Q => reg_in_12_port);
   reg_in_regx11x : DFFSNQ_X1 port map( D => Plaintext(11), CLK => clk, SN => 
                           n396, Q => reg_in_11_port);
   reg_in_regx10x : DFFSNQ_X1 port map( D => Plaintext(10), CLK => clk, SN => 
                           n395, Q => reg_in_10_port);
   reg_in_regx9x : DFFSNQ_X1 port map( D => Plaintext(9), CLK => clk, SN => 
                           n394, Q => reg_in_9_port);
   reg_in_regx8x : DFFSNQ_X1 port map( D => Plaintext(8), CLK => clk, SN => 
                           n393, Q => reg_in_8_port);
   reg_in_regx7x : DFFSNQ_X1 port map( D => Plaintext(7), CLK => clk, SN => 
                           n392, Q => reg_in_7_port);
   reg_in_regx6x : DFFSNQ_X1 port map( D => Plaintext(6), CLK => clk, SN => 
                           n391, Q => reg_in_6_port);
   reg_in_regx5x : DFFSNQ_X1 port map( D => Plaintext(5), CLK => clk, SN => 
                           n390, Q => reg_in_5_port);
   reg_in_regx4x : DFFSNQ_X1 port map( D => Plaintext(4), CLK => clk, SN => 
                           n389, Q => reg_in_4_port);
   reg_in_regx3x : DFFSNQ_X1 port map( D => Plaintext(3), CLK => clk, SN => 
                           n388, Q => reg_in_3_port);
   reg_in_regx2x : DFFSNQ_X1 port map( D => Plaintext(2), CLK => clk, SN => 
                           n387, Q => reg_in_2_port);
   reg_in_regx1x : DFFSNQ_X1 port map( D => Plaintext(1), CLK => clk, SN => 
                           n386, Q => reg_in_1_port);
   reg_in_regx0x : DFFSNQ_X1 port map( D => Plaintext(0), CLK => clk, SN => 
                           n385, Q => reg_in_0_port);
   reg_key_regx191x : DFFSNQ_X1 port map( D => Key(191), CLK => clk, SN => n384
                           , Q => reg_key_191_port);
   reg_key_regx190x : DFFSNQ_X1 port map( D => Key(190), CLK => clk, SN => n383
                           , Q => reg_key_190_port);
   reg_key_regx189x : DFFSNQ_X1 port map( D => Key(189), CLK => clk, SN => n382
                           , Q => reg_key_189_port);
   reg_key_regx188x : DFFSNQ_X1 port map( D => Key(188), CLK => clk, SN => n381
                           , Q => reg_key_188_port);
   reg_key_regx187x : DFFSNQ_X1 port map( D => Key(187), CLK => clk, SN => n380
                           , Q => reg_key_187_port);
   reg_key_regx186x : DFFSNQ_X1 port map( D => Key(186), CLK => clk, SN => n379
                           , Q => reg_key_186_port);
   reg_key_regx185x : DFFSNQ_X1 port map( D => Key(185), CLK => clk, SN => n378
                           , Q => reg_key_185_port);
   reg_key_regx184x : DFFSNQ_X1 port map( D => Key(184), CLK => clk, SN => n377
                           , Q => reg_key_184_port);
   reg_key_regx183x : DFFSNQ_X1 port map( D => Key(183), CLK => clk, SN => n376
                           , Q => reg_key_183_port);
   reg_key_regx182x : DFFSNQ_X1 port map( D => Key(182), CLK => clk, SN => n375
                           , Q => reg_key_182_port);
   reg_key_regx181x : DFFSNQ_X1 port map( D => Key(181), CLK => clk, SN => n374
                           , Q => reg_key_181_port);
   reg_key_regx180x : DFFSNQ_X1 port map( D => Key(180), CLK => clk, SN => n373
                           , Q => reg_key_180_port);
   reg_key_regx179x : DFFSNQ_X1 port map( D => Key(179), CLK => clk, SN => n372
                           , Q => reg_key_179_port);
   reg_key_regx178x : DFFSNQ_X1 port map( D => Key(178), CLK => clk, SN => n371
                           , Q => reg_key_178_port);
   reg_key_regx177x : DFFSNQ_X1 port map( D => Key(177), CLK => clk, SN => n370
                           , Q => reg_key_177_port);
   reg_key_regx176x : DFFSNQ_X1 port map( D => Key(176), CLK => clk, SN => n369
                           , Q => reg_key_176_port);
   reg_key_regx175x : DFFSNQ_X1 port map( D => Key(175), CLK => clk, SN => n368
                           , Q => reg_key_175_port);
   reg_key_regx174x : DFFSNQ_X1 port map( D => Key(174), CLK => clk, SN => n367
                           , Q => reg_key_174_port);
   reg_key_regx173x : DFFSNQ_X1 port map( D => Key(173), CLK => clk, SN => n366
                           , Q => reg_key_173_port);
   reg_key_regx172x : DFFSNQ_X1 port map( D => Key(172), CLK => clk, SN => n365
                           , Q => reg_key_172_port);
   reg_key_regx171x : DFFSNQ_X1 port map( D => Key(171), CLK => clk, SN => n364
                           , Q => reg_key_171_port);
   reg_key_regx170x : DFFSNQ_X1 port map( D => Key(170), CLK => clk, SN => n363
                           , Q => reg_key_170_port);
   reg_key_regx169x : DFFSNQ_X1 port map( D => Key(169), CLK => clk, SN => n362
                           , Q => reg_key_169_port);
   reg_key_regx168x : DFFSNQ_X1 port map( D => Key(168), CLK => clk, SN => n361
                           , Q => reg_key_168_port);
   reg_key_regx167x : DFFSNQ_X1 port map( D => Key(167), CLK => clk, SN => n360
                           , Q => reg_key_167_port);
   reg_key_regx166x : DFFSNQ_X1 port map( D => Key(166), CLK => clk, SN => n359
                           , Q => reg_key_166_port);
   reg_key_regx165x : DFFSNQ_X1 port map( D => Key(165), CLK => clk, SN => n358
                           , Q => reg_key_165_port);
   reg_key_regx164x : DFFSNQ_X1 port map( D => Key(164), CLK => clk, SN => n357
                           , Q => reg_key_164_port);
   reg_key_regx163x : DFFSNQ_X1 port map( D => Key(163), CLK => clk, SN => n356
                           , Q => reg_key_163_port);
   reg_key_regx162x : DFFSNQ_X1 port map( D => Key(162), CLK => clk, SN => n355
                           , Q => reg_key_162_port);
   reg_key_regx161x : DFFSNQ_X1 port map( D => Key(161), CLK => clk, SN => n354
                           , Q => reg_key_161_port);
   reg_key_regx160x : DFFSNQ_X1 port map( D => Key(160), CLK => clk, SN => n353
                           , Q => reg_key_160_port);
   reg_key_regx159x : DFFSNQ_X1 port map( D => Key(159), CLK => clk, SN => n352
                           , Q => reg_key_159_port);
   reg_key_regx158x : DFFSNQ_X1 port map( D => Key(158), CLK => clk, SN => n351
                           , Q => reg_key_158_port);
   reg_key_regx157x : DFFSNQ_X1 port map( D => Key(157), CLK => clk, SN => n350
                           , Q => reg_key_157_port);
   reg_key_regx156x : DFFSNQ_X1 port map( D => Key(156), CLK => clk, SN => n349
                           , Q => reg_key_156_port);
   reg_key_regx155x : DFFSNQ_X1 port map( D => Key(155), CLK => clk, SN => n348
                           , Q => reg_key_155_port);
   reg_key_regx154x : DFFSNQ_X1 port map( D => Key(154), CLK => clk, SN => n347
                           , Q => reg_key_154_port);
   reg_key_regx153x : DFFSNQ_X1 port map( D => Key(153), CLK => clk, SN => n346
                           , Q => reg_key_153_port);
   reg_key_regx152x : DFFSNQ_X1 port map( D => Key(152), CLK => clk, SN => n345
                           , Q => reg_key_152_port);
   reg_key_regx151x : DFFSNQ_X1 port map( D => Key(151), CLK => clk, SN => n344
                           , Q => reg_key_151_port);
   reg_key_regx150x : DFFSNQ_X1 port map( D => Key(150), CLK => clk, SN => n343
                           , Q => reg_key_150_port);
   reg_key_regx149x : DFFSNQ_X1 port map( D => Key(149), CLK => clk, SN => n342
                           , Q => reg_key_149_port);
   reg_key_regx148x : DFFSNQ_X1 port map( D => Key(148), CLK => clk, SN => n341
                           , Q => reg_key_148_port);
   reg_key_regx147x : DFFSNQ_X1 port map( D => Key(147), CLK => clk, SN => n340
                           , Q => reg_key_147_port);
   reg_key_regx146x : DFFSNQ_X1 port map( D => Key(146), CLK => clk, SN => n339
                           , Q => reg_key_146_port);
   reg_key_regx145x : DFFSNQ_X1 port map( D => Key(145), CLK => clk, SN => n338
                           , Q => reg_key_145_port);
   reg_key_regx144x : DFFSNQ_X1 port map( D => Key(144), CLK => clk, SN => n337
                           , Q => reg_key_144_port);
   reg_key_regx143x : DFFSNQ_X1 port map( D => Key(143), CLK => clk, SN => n336
                           , Q => reg_key_143_port);
   reg_key_regx142x : DFFSNQ_X1 port map( D => Key(142), CLK => clk, SN => n335
                           , Q => reg_key_142_port);
   reg_key_regx141x : DFFSNQ_X1 port map( D => Key(141), CLK => clk, SN => n334
                           , Q => reg_key_141_port);
   reg_key_regx140x : DFFSNQ_X1 port map( D => Key(140), CLK => clk, SN => n333
                           , Q => reg_key_140_port);
   reg_key_regx139x : DFFSNQ_X1 port map( D => Key(139), CLK => clk, SN => n332
                           , Q => reg_key_139_port);
   reg_key_regx138x : DFFSNQ_X1 port map( D => Key(138), CLK => clk, SN => n331
                           , Q => reg_key_138_port);
   reg_key_regx137x : DFFSNQ_X1 port map( D => Key(137), CLK => clk, SN => n330
                           , Q => reg_key_137_port);
   reg_key_regx136x : DFFSNQ_X1 port map( D => Key(136), CLK => clk, SN => n329
                           , Q => reg_key_136_port);
   reg_key_regx135x : DFFSNQ_X1 port map( D => Key(135), CLK => clk, SN => n328
                           , Q => reg_key_135_port);
   reg_key_regx134x : DFFSNQ_X1 port map( D => Key(134), CLK => clk, SN => n327
                           , Q => reg_key_134_port);
   reg_key_regx133x : DFFSNQ_X1 port map( D => Key(133), CLK => clk, SN => n326
                           , Q => reg_key_133_port);
   reg_key_regx132x : DFFSNQ_X1 port map( D => Key(132), CLK => clk, SN => n325
                           , Q => reg_key_132_port);
   reg_key_regx131x : DFFSNQ_X1 port map( D => Key(131), CLK => clk, SN => n324
                           , Q => reg_key_131_port);
   reg_key_regx130x : DFFSNQ_X1 port map( D => Key(130), CLK => clk, SN => n323
                           , Q => reg_key_130_port);
   reg_key_regx129x : DFFSNQ_X1 port map( D => Key(129), CLK => clk, SN => n322
                           , Q => reg_key_129_port);
   reg_key_regx128x : DFFSNQ_X1 port map( D => Key(128), CLK => clk, SN => n321
                           , Q => reg_key_128_port);
   reg_key_regx127x : DFFSNQ_X1 port map( D => Key(127), CLK => clk, SN => n320
                           , Q => reg_key_127_port);
   reg_key_regx126x : DFFSNQ_X1 port map( D => Key(126), CLK => clk, SN => n319
                           , Q => reg_key_126_port);
   reg_key_regx125x : DFFSNQ_X1 port map( D => Key(125), CLK => clk, SN => n318
                           , Q => reg_key_125_port);
   reg_key_regx124x : DFFSNQ_X1 port map( D => Key(124), CLK => clk, SN => n317
                           , Q => reg_key_124_port);
   reg_key_regx123x : DFFSNQ_X1 port map( D => Key(123), CLK => clk, SN => n316
                           , Q => reg_key_123_port);
   reg_key_regx122x : DFFSNQ_X1 port map( D => Key(122), CLK => clk, SN => n315
                           , Q => reg_key_122_port);
   reg_key_regx121x : DFFSNQ_X1 port map( D => Key(121), CLK => clk, SN => n314
                           , Q => reg_key_121_port);
   reg_key_regx120x : DFFSNQ_X1 port map( D => Key(120), CLK => clk, SN => n313
                           , Q => reg_key_120_port);
   reg_key_regx119x : DFFSNQ_X1 port map( D => Key(119), CLK => clk, SN => n312
                           , Q => reg_key_119_port);
   reg_key_regx118x : DFFSNQ_X1 port map( D => Key(118), CLK => clk, SN => n311
                           , Q => reg_key_118_port);
   reg_key_regx117x : DFFSNQ_X1 port map( D => Key(117), CLK => clk, SN => n310
                           , Q => reg_key_117_port);
   reg_key_regx116x : DFFSNQ_X1 port map( D => Key(116), CLK => clk, SN => n309
                           , Q => reg_key_116_port);
   reg_key_regx115x : DFFSNQ_X1 port map( D => Key(115), CLK => clk, SN => n308
                           , Q => reg_key_115_port);
   reg_key_regx114x : DFFSNQ_X1 port map( D => Key(114), CLK => clk, SN => n307
                           , Q => reg_key_114_port);
   reg_key_regx113x : DFFSNQ_X1 port map( D => Key(113), CLK => clk, SN => n306
                           , Q => reg_key_113_port);
   reg_key_regx112x : DFFSNQ_X1 port map( D => Key(112), CLK => clk, SN => n305
                           , Q => reg_key_112_port);
   reg_key_regx111x : DFFSNQ_X1 port map( D => Key(111), CLK => clk, SN => n304
                           , Q => reg_key_111_port);
   reg_key_regx110x : DFFSNQ_X1 port map( D => Key(110), CLK => clk, SN => n303
                           , Q => reg_key_110_port);
   reg_key_regx109x : DFFSNQ_X1 port map( D => Key(109), CLK => clk, SN => n302
                           , Q => reg_key_109_port);
   reg_key_regx108x : DFFSNQ_X1 port map( D => Key(108), CLK => clk, SN => n301
                           , Q => reg_key_108_port);
   reg_key_regx107x : DFFSNQ_X1 port map( D => Key(107), CLK => clk, SN => n300
                           , Q => reg_key_107_port);
   reg_key_regx106x : DFFSNQ_X1 port map( D => Key(106), CLK => clk, SN => n299
                           , Q => reg_key_106_port);
   reg_key_regx105x : DFFSNQ_X1 port map( D => Key(105), CLK => clk, SN => n298
                           , Q => reg_key_105_port);
   reg_key_regx104x : DFFSNQ_X1 port map( D => Key(104), CLK => clk, SN => n297
                           , Q => reg_key_104_port);
   reg_key_regx103x : DFFSNQ_X1 port map( D => Key(103), CLK => clk, SN => n296
                           , Q => reg_key_103_port);
   reg_key_regx102x : DFFSNQ_X1 port map( D => Key(102), CLK => clk, SN => n295
                           , Q => reg_key_102_port);
   reg_key_regx101x : DFFSNQ_X1 port map( D => Key(101), CLK => clk, SN => n294
                           , Q => reg_key_101_port);
   reg_key_regx100x : DFFSNQ_X1 port map( D => Key(100), CLK => clk, SN => n293
                           , Q => reg_key_100_port);
   reg_key_regx99x : DFFSNQ_X1 port map( D => Key(99), CLK => clk, SN => n292, 
                           Q => reg_key_99_port);
   reg_key_regx98x : DFFSNQ_X1 port map( D => Key(98), CLK => clk, SN => n291, 
                           Q => reg_key_98_port);
   reg_key_regx97x : DFFSNQ_X1 port map( D => Key(97), CLK => clk, SN => n290, 
                           Q => reg_key_97_port);
   reg_key_regx96x : DFFSNQ_X1 port map( D => Key(96), CLK => clk, SN => n289, 
                           Q => reg_key_96_port);
   reg_key_regx95x : DFFSNQ_X1 port map( D => Key(95), CLK => clk, SN => n288, 
                           Q => reg_key_95_port);
   reg_key_regx94x : DFFSNQ_X1 port map( D => Key(94), CLK => clk, SN => n287, 
                           Q => reg_key_94_port);
   reg_key_regx93x : DFFSNQ_X1 port map( D => Key(93), CLK => clk, SN => n286, 
                           Q => reg_key_93_port);
   reg_key_regx92x : DFFSNQ_X1 port map( D => Key(92), CLK => clk, SN => n285, 
                           Q => reg_key_92_port);
   reg_key_regx91x : DFFSNQ_X1 port map( D => Key(91), CLK => clk, SN => n284, 
                           Q => reg_key_91_port);
   reg_key_regx90x : DFFSNQ_X1 port map( D => Key(90), CLK => clk, SN => n283, 
                           Q => reg_key_90_port);
   reg_key_regx89x : DFFSNQ_X1 port map( D => Key(89), CLK => clk, SN => n282, 
                           Q => reg_key_89_port);
   reg_key_regx88x : DFFSNQ_X1 port map( D => Key(88), CLK => clk, SN => n281, 
                           Q => reg_key_88_port);
   reg_key_regx87x : DFFSNQ_X1 port map( D => Key(87), CLK => clk, SN => n280, 
                           Q => reg_key_87_port);
   reg_key_regx86x : DFFSNQ_X1 port map( D => Key(86), CLK => clk, SN => n279, 
                           Q => reg_key_86_port);
   reg_key_regx85x : DFFSNQ_X1 port map( D => Key(85), CLK => clk, SN => n278, 
                           Q => reg_key_85_port);
   reg_key_regx84x : DFFSNQ_X1 port map( D => Key(84), CLK => clk, SN => n277, 
                           Q => reg_key_84_port);
   reg_key_regx83x : DFFSNQ_X1 port map( D => Key(83), CLK => clk, SN => n276, 
                           Q => reg_key_83_port);
   reg_key_regx82x : DFFSNQ_X1 port map( D => Key(82), CLK => clk, SN => n275, 
                           Q => reg_key_82_port);
   reg_key_regx81x : DFFSNQ_X1 port map( D => Key(81), CLK => clk, SN => n274, 
                           Q => reg_key_81_port);
   reg_key_regx80x : DFFSNQ_X1 port map( D => Key(80), CLK => clk, SN => n273, 
                           Q => reg_key_80_port);
   reg_key_regx79x : DFFSNQ_X1 port map( D => Key(79), CLK => clk, SN => n272, 
                           Q => reg_key_79_port);
   reg_key_regx78x : DFFSNQ_X1 port map( D => Key(78), CLK => clk, SN => n271, 
                           Q => reg_key_78_port);
   reg_key_regx77x : DFFSNQ_X1 port map( D => Key(77), CLK => clk, SN => n270, 
                           Q => reg_key_77_port);
   reg_key_regx76x : DFFSNQ_X1 port map( D => Key(76), CLK => clk, SN => n269, 
                           Q => reg_key_76_port);
   reg_key_regx75x : DFFSNQ_X1 port map( D => Key(75), CLK => clk, SN => n268, 
                           Q => reg_key_75_port);
   reg_key_regx74x : DFFSNQ_X1 port map( D => Key(74), CLK => clk, SN => n267, 
                           Q => reg_key_74_port);
   reg_key_regx73x : DFFSNQ_X1 port map( D => Key(73), CLK => clk, SN => n266, 
                           Q => reg_key_73_port);
   reg_key_regx72x : DFFSNQ_X1 port map( D => Key(72), CLK => clk, SN => n265, 
                           Q => reg_key_72_port);
   reg_key_regx71x : DFFSNQ_X1 port map( D => Key(71), CLK => clk, SN => n264, 
                           Q => reg_key_71_port);
   reg_key_regx70x : DFFSNQ_X1 port map( D => Key(70), CLK => clk, SN => n263, 
                           Q => reg_key_70_port);
   reg_key_regx69x : DFFSNQ_X1 port map( D => Key(69), CLK => clk, SN => n262, 
                           Q => reg_key_69_port);
   reg_key_regx68x : DFFSNQ_X1 port map( D => Key(68), CLK => clk, SN => n261, 
                           Q => reg_key_68_port);
   reg_key_regx67x : DFFSNQ_X1 port map( D => Key(67), CLK => clk, SN => n260, 
                           Q => reg_key_67_port);
   reg_key_regx66x : DFFSNQ_X1 port map( D => Key(66), CLK => clk, SN => n259, 
                           Q => reg_key_66_port);
   reg_key_regx65x : DFFSNQ_X1 port map( D => Key(65), CLK => clk, SN => n258, 
                           Q => reg_key_65_port);
   reg_key_regx64x : DFFSNQ_X1 port map( D => Key(64), CLK => clk, SN => n257, 
                           Q => reg_key_64_port);
   reg_key_regx63x : DFFSNQ_X1 port map( D => Key(63), CLK => clk, SN => n256, 
                           Q => reg_key_63_port);
   reg_key_regx62x : DFFSNQ_X1 port map( D => Key(62), CLK => clk, SN => n255, 
                           Q => reg_key_62_port);
   reg_key_regx61x : DFFSNQ_X1 port map( D => Key(61), CLK => clk, SN => n254, 
                           Q => reg_key_61_port);
   reg_key_regx60x : DFFSNQ_X1 port map( D => Key(60), CLK => clk, SN => n253, 
                           Q => reg_key_60_port);
   reg_key_regx59x : DFFSNQ_X1 port map( D => Key(59), CLK => clk, SN => n252, 
                           Q => reg_key_59_port);
   reg_key_regx58x : DFFSNQ_X1 port map( D => Key(58), CLK => clk, SN => n251, 
                           Q => reg_key_58_port);
   reg_key_regx57x : DFFSNQ_X1 port map( D => Key(57), CLK => clk, SN => n250, 
                           Q => reg_key_57_port);
   reg_key_regx56x : DFFSNQ_X1 port map( D => Key(56), CLK => clk, SN => n249, 
                           Q => reg_key_56_port);
   reg_key_regx55x : DFFSNQ_X1 port map( D => Key(55), CLK => clk, SN => n248, 
                           Q => reg_key_55_port);
   reg_key_regx54x : DFFSNQ_X1 port map( D => Key(54), CLK => clk, SN => n247, 
                           Q => reg_key_54_port);
   reg_key_regx53x : DFFSNQ_X1 port map( D => Key(53), CLK => clk, SN => n246, 
                           Q => reg_key_53_port);
   reg_key_regx52x : DFFSNQ_X1 port map( D => Key(52), CLK => clk, SN => n245, 
                           Q => reg_key_52_port);
   reg_key_regx51x : DFFSNQ_X1 port map( D => Key(51), CLK => clk, SN => n244, 
                           Q => reg_key_51_port);
   reg_key_regx50x : DFFSNQ_X1 port map( D => Key(50), CLK => clk, SN => n243, 
                           Q => reg_key_50_port);
   reg_key_regx49x : DFFSNQ_X1 port map( D => Key(49), CLK => clk, SN => n242, 
                           Q => reg_key_49_port);
   reg_key_regx48x : DFFSNQ_X1 port map( D => Key(48), CLK => clk, SN => n241, 
                           Q => reg_key_48_port);
   reg_key_regx46x : DFFSNQ_X1 port map( D => Key(46), CLK => clk, SN => n239, 
                           Q => reg_key_46_port);
   reg_key_regx45x : DFFSNQ_X1 port map( D => Key(45), CLK => clk, SN => n238, 
                           Q => reg_key_45_port);
   reg_key_regx44x : DFFSNQ_X1 port map( D => Key(44), CLK => clk, SN => n237, 
                           Q => reg_key_44_port);
   reg_key_regx43x : DFFSNQ_X1 port map( D => Key(43), CLK => clk, SN => n236, 
                           Q => reg_key_43_port);
   reg_key_regx42x : DFFSNQ_X1 port map( D => Key(42), CLK => clk, SN => n235, 
                           Q => reg_key_42_port);
   reg_key_regx41x : DFFSNQ_X1 port map( D => Key(41), CLK => clk, SN => n234, 
                           Q => reg_key_41_port);
   reg_key_regx40x : DFFSNQ_X1 port map( D => Key(40), CLK => clk, SN => n233, 
                           Q => reg_key_40_port);
   reg_key_regx39x : DFFSNQ_X1 port map( D => Key(39), CLK => clk, SN => n232, 
                           Q => reg_key_39_port);
   reg_key_regx38x : DFFSNQ_X1 port map( D => Key(38), CLK => clk, SN => n231, 
                           Q => reg_key_38_port);
   reg_key_regx37x : DFFSNQ_X1 port map( D => Key(37), CLK => clk, SN => n230, 
                           Q => reg_key_37_port);
   reg_key_regx36x : DFFSNQ_X1 port map( D => Key(36), CLK => clk, SN => n229, 
                           Q => reg_key_36_port);
   reg_key_regx35x : DFFSNQ_X1 port map( D => Key(35), CLK => clk, SN => n228, 
                           Q => reg_key_35_port);
   reg_key_regx34x : DFFSNQ_X1 port map( D => Key(34), CLK => clk, SN => n227, 
                           Q => reg_key_34_port);
   reg_key_regx33x : DFFSNQ_X1 port map( D => Key(33), CLK => clk, SN => n226, 
                           Q => reg_key_33_port);
   reg_key_regx32x : DFFSNQ_X1 port map( D => Key(32), CLK => clk, SN => n225, 
                           Q => reg_key_32_port);
   reg_key_regx31x : DFFSNQ_X1 port map( D => Key(31), CLK => clk, SN => n224, 
                           Q => reg_key_31_port);
   reg_key_regx30x : DFFSNQ_X1 port map( D => Key(30), CLK => clk, SN => n223, 
                           Q => reg_key_30_port);
   reg_key_regx29x : DFFSNQ_X1 port map( D => Key(29), CLK => clk, SN => n222, 
                           Q => reg_key_29_port);
   reg_key_regx28x : DFFSNQ_X1 port map( D => Key(28), CLK => clk, SN => n221, 
                           Q => reg_key_28_port);
   reg_key_regx27x : DFFSNQ_X1 port map( D => Key(27), CLK => clk, SN => n220, 
                           Q => reg_key_27_port);
   reg_key_regx26x : DFFSNQ_X1 port map( D => Key(26), CLK => clk, SN => n219, 
                           Q => reg_key_26_port);
   reg_key_regx25x : DFFSNQ_X1 port map( D => Key(25), CLK => clk, SN => n218, 
                           Q => reg_key_25_port);
   reg_key_regx24x : DFFSNQ_X1 port map( D => Key(24), CLK => clk, SN => n217, 
                           Q => reg_key_24_port);
   reg_key_regx23x : DFFSNQ_X1 port map( D => Key(23), CLK => clk, SN => n216, 
                           Q => reg_key_23_port);
   reg_key_regx22x : DFFSNQ_X1 port map( D => Key(22), CLK => clk, SN => n215, 
                           Q => reg_key_22_port);
   reg_key_regx21x : DFFSNQ_X1 port map( D => Key(21), CLK => clk, SN => n214, 
                           Q => reg_key_21_port);
   reg_key_regx20x : DFFSNQ_X1 port map( D => Key(20), CLK => clk, SN => n213, 
                           Q => reg_key_20_port);
   reg_key_regx19x : DFFSNQ_X1 port map( D => Key(19), CLK => clk, SN => n212, 
                           Q => reg_key_19_port);
   reg_key_regx18x : DFFSNQ_X1 port map( D => Key(18), CLK => clk, SN => n211, 
                           Q => reg_key_18_port);
   reg_key_regx17x : DFFSNQ_X1 port map( D => Key(17), CLK => clk, SN => n210, 
                           Q => reg_key_17_port);
   reg_key_regx16x : DFFSNQ_X1 port map( D => Key(16), CLK => clk, SN => n209, 
                           Q => reg_key_16_port);
   reg_key_regx15x : DFFSNQ_X1 port map( D => Key(15), CLK => clk, SN => n208, 
                           Q => reg_key_15_port);
   reg_key_regx13x : DFFSNQ_X1 port map( D => Key(13), CLK => clk, SN => n206, 
                           Q => reg_key_13_port);
   reg_key_regx12x : DFFSNQ_X1 port map( D => Key(12), CLK => clk, SN => n205, 
                           Q => reg_key_12_port);
   reg_key_regx11x : DFFSNQ_X1 port map( D => Key(11), CLK => clk, SN => n204, 
                           Q => reg_key_11_port);
   reg_key_regx10x : DFFSNQ_X1 port map( D => Key(10), CLK => clk, SN => n203, 
                           Q => reg_key_10_port);
   reg_key_regx9x : DFFSNQ_X1 port map( D => Key(9), CLK => clk, SN => n202, Q 
                           => reg_key_9_port);
   reg_key_regx7x : DFFSNQ_X1 port map( D => Key(7), CLK => clk, SN => n200, Q 
                           => reg_key_7_port);
   reg_key_regx6x : DFFSNQ_X1 port map( D => Key(6), CLK => clk, SN => n199, Q 
                           => reg_key_6_port);
   reg_key_regx5x : DFFSNQ_X1 port map( D => Key(5), CLK => clk, SN => n198, Q 
                           => reg_key_5_port);
   reg_key_regx4x : DFFSNQ_X1 port map( D => Key(4), CLK => clk, SN => n197, Q 
                           => reg_key_4_port);
   reg_key_regx3x : DFFSNQ_X1 port map( D => Key(3), CLK => clk, SN => n196, Q 
                           => reg_key_3_port);
   reg_key_regx2x : DFFSNQ_X1 port map( D => Key(2), CLK => clk, SN => n195, Q 
                           => reg_key_2_port);
   reg_key_regx1x : DFFSNQ_X1 port map( D => Key(1), CLK => clk, SN => n194, Q 
                           => reg_key_1_port);
   reg_key_regx0x : DFFSNQ_X1 port map( D => Key(0), CLK => clk, SN => n193, Q 
                           => reg_key_0_port);
   Ciphertext_regx190x : DFFSNQ_X1 port map( D => reg_out_190_port, CLK => clk,
                           SN => n191, Q => Ciphertext(190));
   Ciphertext_regx188x : DFFSNQ_X1 port map( D => reg_out_188_port, CLK => clk,
                           SN => n189, Q => Ciphertext(188));
   Ciphertext_regx184x : DFFSNQ_X1 port map( D => reg_out_184_port, CLK => clk,
                           SN => n185, Q => Ciphertext(184));
   Ciphertext_regx183x : DFFSNQ_X1 port map( D => reg_out_183_port, CLK => clk,
                           SN => n184, Q => Ciphertext(183));
   Ciphertext_regx172x : DFFSNQ_X1 port map( D => reg_out_172_port, CLK => clk,
                           SN => n173, Q => Ciphertext(172));
   Ciphertext_regx170x : DFFSNQ_X1 port map( D => reg_out_170_port, CLK => clk,
                           SN => n171, Q => Ciphertext(170));
   Ciphertext_regx169x : DFFSNQ_X1 port map( D => reg_out_169_port, CLK => clk,
                           SN => n170, Q => Ciphertext(169));
   Ciphertext_regx166x : DFFSNQ_X1 port map( D => reg_out_166_port, CLK => clk,
                           SN => n167, Q => Ciphertext(166));
   Ciphertext_regx165x : DFFSNQ_X1 port map( D => reg_out_165_port, CLK => clk,
                           SN => n166, Q => Ciphertext(165));
   Ciphertext_regx164x : DFFSNQ_X1 port map( D => reg_out_164_port, CLK => clk,
                           SN => n165, Q => Ciphertext(164));
   Ciphertext_regx163x : DFFSNQ_X1 port map( D => reg_out_163_port, CLK => clk,
                           SN => n164, Q => Ciphertext(163));
   Ciphertext_regx160x : DFFSNQ_X1 port map( D => reg_out_160_port, CLK => clk,
                           SN => n161, Q => Ciphertext(160));
   Ciphertext_regx156x : DFFSNQ_X1 port map( D => reg_out_156_port, CLK => clk,
                           SN => n157, Q => Ciphertext(156));
   Ciphertext_regx155x : DFFSNQ_X1 port map( D => reg_out_155_port, CLK => clk,
                           SN => n156, Q => Ciphertext(155));
   Ciphertext_regx154x : DFFSNQ_X1 port map( D => reg_out_154_port, CLK => clk,
                           SN => n155, Q => Ciphertext(154));
   Ciphertext_regx153x : DFFSNQ_X1 port map( D => reg_out_153_port, CLK => clk,
                           SN => n154, Q => Ciphertext(153));
   Ciphertext_regx150x : DFFSNQ_X1 port map( D => reg_out_150_port, CLK => clk,
                           SN => n151, Q => Ciphertext(150));
   Ciphertext_regx148x : DFFSNQ_X1 port map( D => reg_out_148_port, CLK => clk,
                           SN => n149, Q => Ciphertext(148));
   Ciphertext_regx144x : DFFSNQ_X1 port map( D => reg_out_144_port, CLK => clk,
                           SN => n145, Q => Ciphertext(144));
   Ciphertext_regx141x : DFFSNQ_X1 port map( D => reg_out_141_port, CLK => clk,
                           SN => n142, Q => Ciphertext(141));
   Ciphertext_regx140x : DFFSNQ_X1 port map( D => reg_out_140_port, CLK => clk,
                           SN => n141, Q => Ciphertext(140));
   Ciphertext_regx138x : DFFSNQ_X1 port map( D => reg_out_138_port, CLK => clk,
                           SN => n139, Q => Ciphertext(138));
   Ciphertext_regx136x : DFFSNQ_X1 port map( D => reg_out_136_port, CLK => clk,
                           SN => n137, Q => Ciphertext(136));
   Ciphertext_regx119x : DFFSNQ_X1 port map( D => reg_out_119_port, CLK => clk,
                           SN => n120, Q => Ciphertext(119));
   Ciphertext_regx118x : DFFSNQ_X1 port map( D => reg_out_118_port, CLK => clk,
                           SN => n119, Q => Ciphertext(118));
   Ciphertext_regx108x : DFFSNQ_X1 port map( D => reg_out_108_port, CLK => clk,
                           SN => n109, Q => Ciphertext(108));
   Ciphertext_regx107x : DFFSNQ_X1 port map( D => reg_out_107_port, CLK => clk,
                           SN => n108, Q => Ciphertext(107));
   Ciphertext_regx103x : DFFSNQ_X1 port map( D => reg_out_103_port, CLK => clk,
                           SN => n104, Q => Ciphertext(103));
   Ciphertext_regx99x : DFFSNQ_X1 port map( D => reg_out_99_port, CLK => clk, 
                           SN => n100, Q => Ciphertext(99));
   Ciphertext_regx95x : DFFSNQ_X1 port map( D => reg_out_95_port, CLK => clk, 
                           SN => n96, Q => Ciphertext(95));
   Ciphertext_regx94x : DFFSNQ_X1 port map( D => reg_out_94_port, CLK => clk, 
                           SN => n95, Q => Ciphertext(94));
   Ciphertext_regx93x : DFFSNQ_X1 port map( D => reg_out_93_port, CLK => clk, 
                           SN => n94, Q => Ciphertext(93));
   Ciphertext_regx92x : DFFSNQ_X1 port map( D => reg_out_92_port, CLK => clk, 
                           SN => n93, Q => Ciphertext(92));
   Ciphertext_regx91x : DFFSNQ_X1 port map( D => reg_out_91_port, CLK => clk, 
                           SN => n92, Q => Ciphertext(91));
   Ciphertext_regx89x : DFFSNQ_X1 port map( D => reg_out_89_port, CLK => clk, 
                           SN => n90, Q => Ciphertext(89));
   Ciphertext_regx87x : DFFSNQ_X1 port map( D => reg_out_87_port, CLK => clk, 
                           SN => n88, Q => Ciphertext(87));
   Ciphertext_regx85x : DFFSNQ_X1 port map( D => reg_out_85_port, CLK => clk, 
                           SN => n86, Q => Ciphertext(85));
   Ciphertext_regx82x : DFFSNQ_X1 port map( D => reg_out_82_port, CLK => clk, 
                           SN => n83, Q => Ciphertext(82));
   Ciphertext_regx81x : DFFSNQ_X1 port map( D => reg_out_81_port, CLK => clk, 
                           SN => n82, Q => Ciphertext(81));
   Ciphertext_regx79x : DFFSNQ_X1 port map( D => reg_out_79_port, CLK => clk, 
                           SN => n80, Q => Ciphertext(79));
   Ciphertext_regx76x : DFFSNQ_X1 port map( D => reg_out_76_port, CLK => clk, 
                           SN => n77, Q => Ciphertext(76));
   Ciphertext_regx75x : DFFSNQ_X1 port map( D => reg_out_75_port, CLK => clk, 
                           SN => n76, Q => Ciphertext(75));
   Ciphertext_regx72x : DFFSNQ_X1 port map( D => reg_out_72_port, CLK => clk, 
                           SN => n73, Q => Ciphertext(72));
   Ciphertext_regx70x : DFFSNQ_X1 port map( D => reg_out_70_port, CLK => clk, 
                           SN => n71, Q => Ciphertext(70));
   Ciphertext_regx69x : DFFSNQ_X1 port map( D => reg_out_69_port, CLK => clk, 
                           SN => n70, Q => Ciphertext(69));
   Ciphertext_regx68x : DFFSNQ_X1 port map( D => reg_out_68_port, CLK => clk, 
                           SN => n69, Q => Ciphertext(68));
   Ciphertext_regx65x : DFFSNQ_X1 port map( D => reg_out_65_port, CLK => clk, 
                           SN => n66, Q => Ciphertext(65));
   Ciphertext_regx64x : DFFSNQ_X1 port map( D => reg_out_64_port, CLK => clk, 
                           SN => n65, Q => Ciphertext(64));
   Ciphertext_regx63x : DFFSNQ_X1 port map( D => reg_out_63_port, CLK => clk, 
                           SN => n64, Q => Ciphertext(63));
   Ciphertext_regx62x : DFFSNQ_X1 port map( D => reg_out_62_port, CLK => clk, 
                           SN => n63, Q => Ciphertext(62));
   Ciphertext_regx58x : DFFSNQ_X1 port map( D => reg_out_58_port, CLK => clk, 
                           SN => n59, Q => Ciphertext(58));
   Ciphertext_regx54x : DFFSNQ_X1 port map( D => reg_out_54_port, CLK => clk, 
                           SN => n55, Q => Ciphertext(54));
   Ciphertext_regx53x : DFFSNQ_X1 port map( D => reg_out_53_port, CLK => clk, 
                           SN => n54, Q => Ciphertext(53));
   Ciphertext_regx52x : DFFSNQ_X1 port map( D => reg_out_52_port, CLK => clk, 
                           SN => n53, Q => Ciphertext(52));
   Ciphertext_regx50x : DFFSNQ_X1 port map( D => reg_out_50_port, CLK => clk, 
                           SN => n51, Q => Ciphertext(50));
   Ciphertext_regx47x : DFFSNQ_X1 port map( D => reg_out_47_port, CLK => clk, 
                           SN => n48, Q => Ciphertext(47));
   Ciphertext_regx45x : DFFSNQ_X1 port map( D => reg_out_45_port, CLK => clk, 
                           SN => n46, Q => Ciphertext(45));
   Ciphertext_regx33x : DFFSNQ_X1 port map( D => reg_out_33_port, CLK => clk, 
                           SN => n34, Q => Ciphertext(33));
   Ciphertext_regx32x : DFFSNQ_X1 port map( D => reg_out_32_port, CLK => clk, 
                           SN => n33, Q => Ciphertext(32));
   Ciphertext_regx28x : DFFSNQ_X1 port map( D => reg_out_28_port, CLK => clk, 
                           SN => n29, Q => Ciphertext(28));
   Ciphertext_regx26x : DFFSNQ_X1 port map( D => reg_out_26_port, CLK => clk, 
                           SN => n27, Q => Ciphertext(26));
   Ciphertext_regx23x : DFFSNQ_X1 port map( D => reg_out_23_port, CLK => clk, 
                           SN => n24, Q => Ciphertext(23));
   Ciphertext_regx20x : DFFSNQ_X1 port map( D => reg_out_20_port, CLK => clk, 
                           SN => n21, Q => Ciphertext(20));
   Ciphertext_regx19x : DFFSNQ_X1 port map( D => reg_out_19_port, CLK => clk, 
                           SN => n20, Q => Ciphertext(19));
   Ciphertext_regx18x : DFFSNQ_X1 port map( D => reg_out_18_port, CLK => clk, 
                           SN => n19, Q => Ciphertext(18));
   Ciphertext_regx15x : DFFSNQ_X1 port map( D => reg_out_15_port, CLK => clk, 
                           SN => n16, Q => Ciphertext(15));
   Ciphertext_regx11x : DFFSNQ_X1 port map( D => reg_out_11_port, CLK => clk, 
                           SN => n12, Q => Ciphertext(11));
   Ciphertext_regx10x : DFFSNQ_X1 port map( D => reg_out_10_port, CLK => clk, 
                           SN => n11, Q => Ciphertext(10));
   Ciphertext_regx9x : DFFSNQ_X1 port map( D => reg_out_9_port, CLK => clk, SN 
                           => n10, Q => Ciphertext(9));
   Ciphertext_regx8x : DFFSNQ_X1 port map( D => reg_out_8_port, CLK => clk, SN 
                           => n9, Q => Ciphertext(8));
   Ciphertext_regx4x : DFFSNQ_X1 port map( D => reg_out_4_port, CLK => clk, SN 
                           => n5, Q => Ciphertext(4));
   n5 <= '1';
   n9 <= '1';
   n10 <= '1';
   n11 <= '1';
   n12 <= '1';
   n16 <= '1';
   n19 <= '1';
   n20 <= '1';
   n21 <= '1';
   n24 <= '1';
   n27 <= '1';
   n29 <= '1';
   n33 <= '1';
   n34 <= '1';
   n46 <= '1';
   n48 <= '1';
   n51 <= '1';
   n53 <= '1';
   n54 <= '1';
   n55 <= '1';
   n59 <= '1';
   n63 <= '1';
   n64 <= '1';
   n65 <= '1';
   n66 <= '1';
   n69 <= '1';
   n70 <= '1';
   n71 <= '1';
   n73 <= '1';
   n76 <= '1';
   n77 <= '1';
   n80 <= '1';
   n82 <= '1';
   n83 <= '1';
   n86 <= '1';
   n88 <= '1';
   n90 <= '1';
   n92 <= '1';
   n93 <= '1';
   n94 <= '1';
   n95 <= '1';
   n96 <= '1';
   n100 <= '1';
   n104 <= '1';
   n108 <= '1';
   n109 <= '1';
   n119 <= '1';
   n120 <= '1';
   n137 <= '1';
   n139 <= '1';
   n141 <= '1';
   n142 <= '1';
   n145 <= '1';
   n149 <= '1';
   n151 <= '1';
   n154 <= '1';
   n155 <= '1';
   n156 <= '1';
   n157 <= '1';
   n161 <= '1';
   n164 <= '1';
   n165 <= '1';
   n166 <= '1';
   n167 <= '1';
   n170 <= '1';
   n171 <= '1';
   n173 <= '1';
   n184 <= '1';
   n185 <= '1';
   n189 <= '1';
   n191 <= '1';
   n193 <= '1';
   n194 <= '1';
   n195 <= '1';
   n196 <= '1';
   n197 <= '1';
   n198 <= '1';
   n199 <= '1';
   n200 <= '1';
   n202 <= '1';
   n203 <= '1';
   n204 <= '1';
   n205 <= '1';
   n206 <= '1';
   n208 <= '1';
   n209 <= '1';
   n210 <= '1';
   n211 <= '1';
   n212 <= '1';
   n213 <= '1';
   n214 <= '1';
   n215 <= '1';
   n216 <= '1';
   n217 <= '1';
   n218 <= '1';
   n219 <= '1';
   n220 <= '1';
   n221 <= '1';
   n222 <= '1';
   n223 <= '1';
   n224 <= '1';
   n225 <= '1';
   n226 <= '1';
   n227 <= '1';
   n228 <= '1';
   n229 <= '1';
   n230 <= '1';
   n231 <= '1';
   n232 <= '1';
   n233 <= '1';
   n234 <= '1';
   n235 <= '1';
   n236 <= '1';
   n237 <= '1';
   n238 <= '1';
   n239 <= '1';
   n241 <= '1';
   n242 <= '1';
   n243 <= '1';
   n244 <= '1';
   n245 <= '1';
   n246 <= '1';
   n247 <= '1';
   n248 <= '1';
   n249 <= '1';
   n250 <= '1';
   n251 <= '1';
   n252 <= '1';
   n253 <= '1';
   n254 <= '1';
   n255 <= '1';
   n256 <= '1';
   n257 <= '1';
   n258 <= '1';
   n259 <= '1';
   n260 <= '1';
   n261 <= '1';
   n262 <= '1';
   n263 <= '1';
   n264 <= '1';
   n265 <= '1';
   n266 <= '1';
   n267 <= '1';
   n268 <= '1';
   n269 <= '1';
   n270 <= '1';
   n271 <= '1';
   n272 <= '1';
   n273 <= '1';
   n274 <= '1';
   n275 <= '1';
   n276 <= '1';
   n277 <= '1';
   n278 <= '1';
   n279 <= '1';
   n280 <= '1';
   n281 <= '1';
   n282 <= '1';
   n283 <= '1';
   n284 <= '1';
   n285 <= '1';
   n286 <= '1';
   n287 <= '1';
   n288 <= '1';
   n289 <= '1';
   n290 <= '1';
   n291 <= '1';
   n292 <= '1';
   n293 <= '1';
   n294 <= '1';
   n295 <= '1';
   n296 <= '1';
   n297 <= '1';
   n298 <= '1';
   n299 <= '1';
   n300 <= '1';
   n301 <= '1';
   n302 <= '1';
   n303 <= '1';
   n304 <= '1';
   n305 <= '1';
   n306 <= '1';
   n307 <= '1';
   n308 <= '1';
   n309 <= '1';
   n310 <= '1';
   n311 <= '1';
   n312 <= '1';
   n313 <= '1';
   n314 <= '1';
   n315 <= '1';
   n316 <= '1';
   n317 <= '1';
   n318 <= '1';
   n319 <= '1';
   n320 <= '1';
   n321 <= '1';
   n322 <= '1';
   n323 <= '1';
   n324 <= '1';
   n325 <= '1';
   n326 <= '1';
   n327 <= '1';
   n328 <= '1';
   n329 <= '1';
   n330 <= '1';
   n331 <= '1';
   n332 <= '1';
   n333 <= '1';
   n334 <= '1';
   n335 <= '1';
   n336 <= '1';
   n337 <= '1';
   n338 <= '1';
   n339 <= '1';
   n340 <= '1';
   n341 <= '1';
   n342 <= '1';
   n343 <= '1';
   n344 <= '1';
   n345 <= '1';
   n346 <= '1';
   n347 <= '1';
   n348 <= '1';
   n349 <= '1';
   n350 <= '1';
   n351 <= '1';
   n352 <= '1';
   n353 <= '1';
   n354 <= '1';
   n355 <= '1';
   n356 <= '1';
   n357 <= '1';
   n358 <= '1';
   n359 <= '1';
   n360 <= '1';
   n361 <= '1';
   n362 <= '1';
   n363 <= '1';
   n364 <= '1';
   n365 <= '1';
   n366 <= '1';
   n367 <= '1';
   n368 <= '1';
   n369 <= '1';
   n370 <= '1';
   n371 <= '1';
   n372 <= '1';
   n373 <= '1';
   n374 <= '1';
   n375 <= '1';
   n376 <= '1';
   n377 <= '1';
   n378 <= '1';
   n379 <= '1';
   n380 <= '1';
   n381 <= '1';
   n382 <= '1';
   n383 <= '1';
   n384 <= '1';
   n385 <= '1';
   n386 <= '1';
   n387 <= '1';
   n388 <= '1';
   n389 <= '1';
   n390 <= '1';
   n391 <= '1';
   n392 <= '1';
   n393 <= '1';
   n394 <= '1';
   n395 <= '1';
   n396 <= '1';
   n397 <= '1';
   n398 <= '1';
   n399 <= '1';
   n400 <= '1';
   n401 <= '1';
   n402 <= '1';
   n403 <= '1';
   n404 <= '1';
   n405 <= '1';
   n406 <= '1';
   n407 <= '1';
   n408 <= '1';
   n409 <= '1';
   n410 <= '1';
   n411 <= '1';
   n412 <= '1';
   n413 <= '1';
   n414 <= '1';
   n415 <= '1';
   n416 <= '1';
   n417 <= '1';
   n418 <= '1';
   n419 <= '1';
   n420 <= '1';
   n421 <= '1';
   n422 <= '1';
   n423 <= '1';
   n424 <= '1';
   n425 <= '1';
   n426 <= '1';
   n427 <= '1';
   n428 <= '1';
   n429 <= '1';
   n430 <= '1';
   n431 <= '1';
   n432 <= '1';
   n433 <= '1';
   n434 <= '1';
   n435 <= '1';
   n436 <= '1';
   n437 <= '1';
   n438 <= '1';
   n439 <= '1';
   n440 <= '1';
   n441 <= '1';
   n442 <= '1';
   n443 <= '1';
   n445 <= '1';
   n446 <= '1';
   n447 <= '1';
   n448 <= '1';
   n449 <= '1';
   n450 <= '1';
   n451 <= '1';
   n452 <= '1';
   n453 <= '1';
   n454 <= '1';
   n455 <= '1';
   n456 <= '1';
   n457 <= '1';
   n458 <= '1';
   n459 <= '1';
   n460 <= '1';
   n461 <= '1';
   n462 <= '1';
   n463 <= '1';
   n464 <= '1';
   n466 <= '1';
   n467 <= '1';
   n469 <= '1';
   n470 <= '1';
   n471 <= '1';
   n472 <= '1';
   n473 <= '1';
   n474 <= '1';
   n475 <= '1';
   n476 <= '1';
   n477 <= '1';
   n478 <= '1';
   n479 <= '1';
   n480 <= '1';
   n481 <= '1';
   n482 <= '1';
   n483 <= '1';
   n484 <= '1';
   n485 <= '1';
   n487 <= '1';
   n488 <= '1';
   n489 <= '1';
   n490 <= '1';
   n491 <= '1';
   n492 <= '1';
   n493 <= '1';
   n494 <= '1';
   n495 <= '1';
   n497 <= '1';
   n498 <= '1';
   n499 <= '1';
   n500 <= '1';
   n501 <= '1';
   n502 <= '1';
   n503 <= '1';
   n504 <= '1';
   n505 <= '1';
   n506 <= '1';
   n507 <= '1';
   n508 <= '1';
   n509 <= '1';
   n510 <= '1';
   n511 <= '1';
   n512 <= '1';
   n513 <= '1';
   n514 <= '1';
   n515 <= '1';
   n516 <= '1';
   n517 <= '1';
   n518 <= '1';
   n519 <= '1';
   n520 <= '1';
   n521 <= '1';
   n522 <= '1';
   n523 <= '1';
   n524 <= '1';
   n525 <= '1';
   n526 <= '1';
   n527 <= '1';
   n528 <= '1';
   n529 <= '1';
   n530 <= '1';
   n531 <= '1';
   n532 <= '1';
   n533 <= '1';
   n534 <= '1';
   n535 <= '1';
   n536 <= '1';
   n537 <= '1';
   n538 <= '1';
   n539 <= '1';
   n540 <= '1';
   n541 <= '1';
   n542 <= '1';
   n543 <= '1';
   n544 <= '1';
   n545 <= '1';
   n546 <= '1';
   n547 <= '1';
   n548 <= '1';
   n549 <= '1';
   n550 <= '1';
   n551 <= '1';
   n552 <= '1';
   n553 <= '1';
   n554 <= '1';
   n555 <= '1';
   n556 <= '1';
   n557 <= '1';
   n558 <= '1';
   n559 <= '1';
   n560 <= '1';
   n561 <= '1';
   n562 <= '1';
   n563 <= '1';
   n564 <= '1';
   n565 <= '1';
   n566 <= '1';
   n567 <= '1';
   n568 <= '1';
   n569 <= '1';
   n571 <= '1';
   n572 <= '1';
   n573 <= '1';
   n574 <= '1';
   n575 <= '1';
   n576 <= '1';
   Ciphertext_regx17x : DFFRNQ_X1 port map( D => reg_out_17_port, CLK => clk, 
                           RN => n680, Q => Ciphertext(17));
   Ciphertext_regx112x : DFFRNQ_X1 port map( D => reg_out_112_port, CLK => clk,
                           RN => n679, Q => Ciphertext(112));
   Ciphertext_regx174x : DFFRNQ_X1 port map( D => reg_out_174_port, CLK => clk,
                           RN => n678, Q => Ciphertext(174));
   Ciphertext_regx105x : DFFRNQ_X1 port map( D => reg_out_105_port, CLK => clk,
                           RN => n677, Q => Ciphertext(105));
   Ciphertext_regx181x : DFFRNQ_X1 port map( D => reg_out_181_port, CLK => clk,
                           RN => n676, Q => Ciphertext(181));
   Ciphertext_regx36x : DFFRNQ_X1 port map( D => reg_out_36_port, CLK => clk, 
                           RN => n675, Q => Ciphertext(36));
   Ciphertext_regx34x : DFFRNQ_X1 port map( D => reg_out_34_port, CLK => clk, 
                           RN => n673, Q => Ciphertext(34));
   Ciphertext_regx106x : DFFRNQ_X1 port map( D => reg_out_106_port, CLK => clk,
                           RN => n672, Q => Ciphertext(106));
   Ciphertext_regx41x : DFFRNQ_X1 port map( D => reg_out_41_port, CLK => clk, 
                           RN => n671, Q => Ciphertext(41));
   Ciphertext_regx157x : DFFRNQ_X1 port map( D => reg_out_157_port, CLK => clk,
                           RN => n670, Q => Ciphertext(157));
   Ciphertext_regx145x : DFFRNQ_X1 port map( D => reg_out_145_port, CLK => clk,
                           RN => n669, Q => Ciphertext(145));
   Ciphertext_regx114x : DFFRNQ_X1 port map( D => reg_out_114_port, CLK => clk,
                           RN => n668, Q => Ciphertext(114));
   Ciphertext_regx14x : DFFRNQ_X1 port map( D => reg_out_14_port, CLK => clk, 
                           RN => n667, Q => Ciphertext(14));
   Ciphertext_regx122x : DFFRNQ_X1 port map( D => reg_out_122_port, CLK => clk,
                           RN => n666, Q => Ciphertext(122));
   Ciphertext_regx124x : DFFRNQ_X1 port map( D => reg_out_124_port, CLK => clk,
                           RN => n665, Q => Ciphertext(124));
   Ciphertext_regx88x : DFFRNQ_X1 port map( D => reg_out_88_port, CLK => clk, 
                           RN => n664, Q => Ciphertext(88));
   Ciphertext_regx29x : DFFRNQ_X1 port map( D => reg_out_29_port, CLK => clk, 
                           RN => n663, Q => Ciphertext(29));
   Ciphertext_regx42x : DFFRNQ_X1 port map( D => reg_out_42_port, CLK => clk, 
                           RN => n661, Q => Ciphertext(42));
   Ciphertext_regx176x : DFFRNQ_X1 port map( D => reg_out_176_port, CLK => clk,
                           RN => n660, Q => Ciphertext(176));
   Ciphertext_regx98x : DFFRNQ_X1 port map( D => reg_out_98_port, CLK => clk, 
                           RN => n659, Q => Ciphertext(98));
   Ciphertext_regx111x : DFFRNQ_X1 port map( D => reg_out_111_port, CLK => clk,
                           RN => n658, Q => Ciphertext(111));
   Ciphertext_regx37x : DFFRNQ_X1 port map( D => reg_out_37_port, CLK => clk, 
                           RN => n657, Q => Ciphertext(37));
   Ciphertext_regx143x : DFFRNQ_X1 port map( D => reg_out_143_port, CLK => clk,
                           RN => n656, Q => Ciphertext(143));
   Ciphertext_regx130x : DFFRNQ_X1 port map( D => reg_out_130_port, CLK => clk,
                           RN => n655, Q => Ciphertext(130));
   Ciphertext_regx59x : DFFRNQ_X1 port map( D => reg_out_59_port, CLK => clk, 
                           RN => n654, Q => Ciphertext(59));
   Ciphertext_regx129x : DFFRNQ_X1 port map( D => reg_out_129_port, CLK => clk,
                           RN => n653, Q => Ciphertext(129));
   Ciphertext_regx13x : DFFRNQ_X1 port map( D => reg_out_13_port, CLK => clk, 
                           RN => n652, Q => Ciphertext(13));
   Ciphertext_regx115x : DFFRNQ_X1 port map( D => reg_out_115_port, CLK => clk,
                           RN => n651, Q => Ciphertext(115));
   Ciphertext_regx177x : DFFRNQ_X1 port map( D => reg_out_177_port, CLK => clk,
                           RN => n650, Q => Ciphertext(177));
   Ciphertext_regx44x : DFFRNQ_X1 port map( D => reg_out_44_port, CLK => clk, 
                           RN => n649, Q => Ciphertext(44));
   Ciphertext_regx55x : DFFRNQ_X1 port map( D => reg_out_55_port, CLK => clk, 
                           RN => n648, Q => Ciphertext(55));
   Ciphertext_regx116x : DFFRNQ_X1 port map( D => reg_out_116_port, CLK => clk,
                           RN => n647, Q => Ciphertext(116));
   Ciphertext_regx40x : DFFRNQ_X1 port map( D => reg_out_40_port, CLK => clk, 
                           RN => n646, Q => Ciphertext(40));
   Ciphertext_regx25x : DFFRNQ_X1 port map( D => reg_out_25_port, CLK => clk, 
                           RN => n645, Q => Ciphertext(25));
   Ciphertext_regx187x : DFFRNQ_X1 port map( D => reg_out_187_port, CLK => clk,
                           RN => n644, Q => Ciphertext(187));
   Ciphertext_regx38x : DFFRNQ_X1 port map( D => reg_out_38_port, CLK => clk, 
                           RN => n643, Q => Ciphertext(38));
   Ciphertext_regx83x : DFFRNQ_X1 port map( D => reg_out_83_port, CLK => clk, 
                           RN => n642, Q => Ciphertext(83));
   Ciphertext_regx30x : DFFRNQ_X1 port map( D => reg_out_30_port, CLK => clk, 
                           RN => n641, Q => Ciphertext(30));
   Ciphertext_regx185x : DFFRNQ_X1 port map( D => reg_out_185_port, CLK => clk,
                           RN => n640, Q => Ciphertext(185));
   Ciphertext_regx178x : DFFRNQ_X1 port map( D => reg_out_178_port, CLK => clk,
                           RN => n638, Q => Ciphertext(178));
   Ciphertext_regx120x : DFFRNQ_X1 port map( D => reg_out_120_port, CLK => clk,
                           RN => n637, Q => Ciphertext(120));
   Ciphertext_regx133x : DFFRNQ_X1 port map( D => reg_out_133_port, CLK => clk,
                           RN => n636, Q => Ciphertext(133));
   Ciphertext_regx24x : DFFRNQ_X1 port map( D => reg_out_24_port, CLK => clk, 
                           RN => n635, Q => Ciphertext(24));
   Ciphertext_regx123x : DFFRNQ_X1 port map( D => reg_out_123_port, CLK => clk,
                           RN => n634, Q => Ciphertext(123));
   Ciphertext_regx101x : DFFRNQ_X1 port map( D => reg_out_101_port, CLK => clk,
                           RN => n633, Q => Ciphertext(101));
   Ciphertext_regx167x : DFFRNQ_X1 port map( D => reg_out_167_port, CLK => clk,
                           RN => n632, Q => Ciphertext(167));
   Ciphertext_regx2x : DFFRNQ_X1 port map( D => reg_out_2_port, CLK => clk, RN 
                           => n631, Q => Ciphertext(2));
   Ciphertext_regx158x : DFFRNQ_X1 port map( D => reg_out_158_port, CLK => clk,
                           RN => n630, Q => Ciphertext(158));
   Ciphertext_regx125x : DFFRNQ_X1 port map( D => reg_out_125_port, CLK => clk,
                           RN => n629, Q => Ciphertext(125));
   Ciphertext_regx121x : DFFRNQ_X1 port map( D => reg_out_121_port, CLK => clk,
                           RN => n628, Q => Ciphertext(121));
   Ciphertext_regx102x : DFFRNQ_X1 port map( D => reg_out_102_port, CLK => clk,
                           RN => n627, Q => Ciphertext(102));
   Ciphertext_regx131x : DFFRNQ_X1 port map( D => reg_out_131_port, CLK => clk,
                           RN => n626, Q => Ciphertext(131));
   Ciphertext_regx66x : DFFRNQ_X1 port map( D => reg_out_66_port, CLK => clk, 
                           RN => n625, Q => Ciphertext(66));
   Ciphertext_regx22x : DFFRNQ_X1 port map( D => reg_out_22_port, CLK => clk, 
                           RN => n624, Q => Ciphertext(22));
   Ciphertext_regx182x : DFFRNQ_X1 port map( D => reg_out_182_port, CLK => clk,
                           RN => n623, Q => Ciphertext(182));
   Ciphertext_regx97x : DFFRNQ_X1 port map( D => reg_out_97_port, CLK => clk, 
                           RN => n622, Q => Ciphertext(97));
   Ciphertext_regx180x : DFFRNQ_X1 port map( D => reg_out_180_port, CLK => clk,
                           RN => n621, Q => Ciphertext(180));
   Ciphertext_regx73x : DFFRNQ_X1 port map( D => reg_out_73_port, CLK => clk, 
                           RN => n620, Q => Ciphertext(73));
   Ciphertext_regx117x : DFFRNQ_X1 port map( D => reg_out_117_port, CLK => clk,
                           RN => n619, Q => Ciphertext(117));
   Ciphertext_regx78x : DFFRNQ_X1 port map( D => reg_out_78_port, CLK => clk, 
                           RN => n618, Q => Ciphertext(78));
   Ciphertext_regx152x : DFFRNQ_X1 port map( D => reg_out_152_port, CLK => clk,
                           RN => n617, Q => Ciphertext(152));
   Ciphertext_regx39x : DFFRNQ_X1 port map( D => reg_out_39_port, CLK => clk, 
                           RN => n616, Q => Ciphertext(39));
   Ciphertext_regx74x : DFFRNQ_X1 port map( D => reg_out_74_port, CLK => clk, 
                           RN => n615, Q => Ciphertext(74));
   Ciphertext_regx179x : DFFRNQ_X1 port map( D => reg_out_179_port, CLK => clk,
                           RN => n614, Q => Ciphertext(179));
   Ciphertext_regx132x : DFFRNQ_X1 port map( D => reg_out_132_port, CLK => clk,
                           RN => n613, Q => Ciphertext(132));
   Ciphertext_regx109x : DFFRNQ_X1 port map( D => reg_out_109_port, CLK => clk,
                           RN => n612, Q => Ciphertext(109));
   Ciphertext_regx61x : DFFRNQ_X1 port map( D => reg_out_61_port, CLK => clk, 
                           RN => n611, Q => Ciphertext(61));
   Ciphertext_regx16x : DFFRNQ_X1 port map( D => reg_out_16_port, CLK => clk, 
                           RN => n610, Q => Ciphertext(16));
   Ciphertext_regx134x : DFFRNQ_X1 port map( D => reg_out_134_port, CLK => clk,
                           RN => n609, Q => Ciphertext(134));
   Ciphertext_regx80x : DFFRNQ_X1 port map( D => reg_out_80_port, CLK => clk, 
                           RN => n608, Q => Ciphertext(80));
   Ciphertext_regx46x : DFFRNQ_X1 port map( D => reg_out_46_port, CLK => clk, 
                           RN => n607, Q => Ciphertext(46));
   Ciphertext_regx43x : DFFRNQ_X1 port map( D => reg_out_43_port, CLK => clk, 
                           RN => n606, Q => Ciphertext(43));
   Ciphertext_regx7x : DFFRNQ_X1 port map( D => reg_out_7_port, CLK => clk, RN 
                           => n605, Q => Ciphertext(7));
   Ciphertext_regx110x : DFFRNQ_X1 port map( D => reg_out_110_port, CLK => clk,
                           RN => n604, Q => Ciphertext(110));
   Ciphertext_regx149x : DFFRNQ_X1 port map( D => reg_out_149_port, CLK => clk,
                           RN => n603, Q => Ciphertext(149));
   Ciphertext_regx175x : DFFRNQ_X1 port map( D => reg_out_175_port, CLK => clk,
                           RN => n602, Q => Ciphertext(175));
   Ciphertext_regx128x : DFFRNQ_X1 port map( D => reg_out_128_port, CLK => clk,
                           RN => n601, Q => Ciphertext(128));
   Ciphertext_regx127x : DFFRNQ_X1 port map( D => reg_out_127_port, CLK => clk,
                           RN => n600, Q => Ciphertext(127));
   Ciphertext_regx31x : DFFRNQ_X1 port map( D => reg_out_31_port, CLK => clk, 
                           RN => n599, Q => Ciphertext(31));
   Ciphertext_regx96x : DFFRNQ_X1 port map( D => reg_out_96_port, CLK => clk, 
                           RN => n598, Q => Ciphertext(96));
   Ciphertext_regx113x : DFFRNQ_X1 port map( D => reg_out_113_port, CLK => clk,
                           RN => n597, Q => Ciphertext(113));
   Ciphertext_regx6x : DFFRNQ_X1 port map( D => reg_out_6_port, CLK => clk, RN 
                           => n596, Q => Ciphertext(6));
   Ciphertext_regx191x : DFFRNQ_X1 port map( D => reg_out_191_port, CLK => clk,
                           RN => n595, Q => Ciphertext(191));
   Ciphertext_regx77x : DFFRNQ_X1 port map( D => reg_out_77_port, CLK => clk, 
                           RN => n594, Q => Ciphertext(77));
   Ciphertext_regx104x : DFFRNQ_X1 port map( D => reg_out_104_port, CLK => clk,
                           RN => n593, Q => Ciphertext(104));
   Ciphertext_regx71x : DFFRNQ_X1 port map( D => reg_out_71_port, CLK => clk, 
                           RN => n592, Q => Ciphertext(71));
   Ciphertext_regx1x : DFFRNQ_X1 port map( D => reg_out_1_port, CLK => clk, RN 
                           => n591, Q => Ciphertext(1));
   Ciphertext_regx60x : DFFRNQ_X1 port map( D => reg_out_60_port, CLK => clk, 
                           RN => n590, Q => Ciphertext(60));
   Ciphertext_regx86x : DFFRNQ_X1 port map( D => reg_out_86_port, CLK => clk, 
                           RN => n589, Q => Ciphertext(86));
   Ciphertext_regx139x : DFFRNQ_X1 port map( D => reg_out_139_port, CLK => clk,
                           RN => n588, Q => Ciphertext(139));
   Ciphertext_regx49x : DFFRNQ_X1 port map( D => reg_out_49_port, CLK => clk, 
                           RN => n587, Q => Ciphertext(49));
   Ciphertext_regx173x : DFFRNQ_X1 port map( D => reg_out_173_port, CLK => clk,
                           RN => n586, Q => Ciphertext(173));
   Ciphertext_regx84x : DFFRNQ_X1 port map( D => reg_out_84_port, CLK => clk, 
                           RN => n584, Q => Ciphertext(84));
   Ciphertext_regx35x : DFFRNQ_X1 port map( D => reg_out_35_port, CLK => clk, 
                           RN => n583, Q => Ciphertext(35));
   Ciphertext_regx12x : DFFRNQ_X1 port map( D => reg_out_12_port, CLK => clk, 
                           RN => n582, Q => Ciphertext(12));
   Ciphertext_regx146x : DFFRNQ_X1 port map( D => reg_out_146_port, CLK => clk,
                           RN => n581, Q => Ciphertext(146));
   Ciphertext_regx189x : DFFRNQ_X1 port map( D => reg_out_189_port, CLK => clk,
                           RN => n580, Q => Ciphertext(189));
   Ciphertext_regx137x : DFFRNQ_X1 port map( D => reg_out_137_port, CLK => clk,
                           RN => n579, Q => Ciphertext(137));
   Ciphertext_regx3x : DFFRNQ_X1 port map( D => reg_out_3_port, CLK => clk, RN 
                           => n578, Q => Ciphertext(3));
   Ciphertext_regx142x : DFFRNQ_X1 port map( D => reg_out_142_port, CLK => clk,
                           RN => n577, Q => Ciphertext(142));
   n577 <= '1';
   n578 <= '1';
   n579 <= '1';
   n580 <= '1';
   n581 <= '1';
   n582 <= '1';
   n583 <= '1';
   n584 <= '1';
   n586 <= '1';
   n587 <= '1';
   n588 <= '1';
   n589 <= '1';
   n590 <= '1';
   n591 <= '1';
   n592 <= '1';
   n593 <= '1';
   n594 <= '1';
   n595 <= '1';
   n596 <= '1';
   n597 <= '1';
   n598 <= '1';
   n599 <= '1';
   n600 <= '1';
   n601 <= '1';
   n602 <= '1';
   n603 <= '1';
   n604 <= '1';
   n605 <= '1';
   n606 <= '1';
   n607 <= '1';
   n608 <= '1';
   n609 <= '1';
   n610 <= '1';
   n611 <= '1';
   n612 <= '1';
   n613 <= '1';
   n614 <= '1';
   n615 <= '1';
   n616 <= '1';
   n617 <= '1';
   n618 <= '1';
   n619 <= '1';
   n620 <= '1';
   n621 <= '1';
   n622 <= '1';
   n623 <= '1';
   n624 <= '1';
   n625 <= '1';
   n626 <= '1';
   n627 <= '1';
   n628 <= '1';
   n629 <= '1';
   n630 <= '1';
   n631 <= '1';
   n632 <= '1';
   n633 <= '1';
   n634 <= '1';
   n635 <= '1';
   n636 <= '1';
   n637 <= '1';
   n638 <= '1';
   n640 <= '1';
   n641 <= '1';
   n642 <= '1';
   n643 <= '1';
   n644 <= '1';
   n645 <= '1';
   n646 <= '1';
   n647 <= '1';
   n648 <= '1';
   n649 <= '1';
   n650 <= '1';
   n651 <= '1';
   n652 <= '1';
   n653 <= '1';
   n654 <= '1';
   n655 <= '1';
   n656 <= '1';
   n657 <= '1';
   n658 <= '1';
   n659 <= '1';
   n660 <= '1';
   n661 <= '1';
   n663 <= '1';
   n664 <= '1';
   n665 <= '1';
   n666 <= '1';
   n667 <= '1';
   n668 <= '1';
   n669 <= '1';
   n670 <= '1';
   n671 <= '1';
   n672 <= '1';
   n673 <= '1';
   n675 <= '1';
   n676 <= '1';
   n677 <= '1';
   n678 <= '1';
   n679 <= '1';
   n680 <= '1';
   Ciphertext_regx126x : DFFRNQ_X1 port map( D => reg_out_126_port, CLK => clk,
                           RN => n693, Q => Ciphertext(126));
   Ciphertext_regx162x : DFFRNQ_X1 port map( D => reg_out_162_port, CLK => clk,
                           RN => n692, Q => Ciphertext(162));
   Ciphertext_regx56x : DFFRNQ_X1 port map( D => reg_out_56_port, CLK => clk, 
                           RN => n691, Q => Ciphertext(56));
   Ciphertext_regx5x : DFFRNQ_X1 port map( D => reg_out_5_port, CLK => clk, RN 
                           => n690, Q => Ciphertext(5));
   Ciphertext_regx135x : DFFRNQ_X1 port map( D => reg_out_135_port, CLK => clk,
                           RN => n689, Q => Ciphertext(135));
   Ciphertext_regx57x : DFFRNQ_X1 port map( D => reg_out_57_port, CLK => clk, 
                           RN => n688, Q => Ciphertext(57));
   Ciphertext_regx27x : DFFRNQ_X1 port map( D => reg_out_27_port, CLK => clk, 
                           RN => n687, Q => Ciphertext(27));
   Ciphertext_regx90x : DFFRNQ_X1 port map( D => reg_out_90_port, CLK => clk, 
                           RN => n686, Q => Ciphertext(90));
   reg_key_regx47x : DFFRNQ_X1 port map( D => Key(47), CLK => clk, RN => n685, 
                           Q => reg_key_47_port);
   Ciphertext_regx0x : DFFRNQ_X1 port map( D => reg_out_0_port, CLK => clk, RN 
                           => n684, Q => Ciphertext(0));
   Ciphertext_regx151x : DFFRNQ_X1 port map( D => reg_out_151_port, CLK => clk,
                           RN => n683, Q => Ciphertext(151));
   reg_in_regx101x : DFFRNQ_X1 port map( D => Plaintext(101), CLK => clk, RN =>
                           n682, Q => reg_in_101_port);
   reg_in_regx59x : DFFRNQ_X1 port map( D => Plaintext(59), CLK => clk, RN => 
                           n681, Q => reg_in_59_port);
   n681 <= '1';
   n682 <= '1';
   n683 <= '1';
   n684 <= '1';
   n685 <= '1';
   n686 <= '1';
   n687 <= '1';
   n688 <= '1';
   n689 <= '1';
   n690 <= '1';
   n691 <= '1';
   n692 <= '1';
   n693 <= '1';
   Ciphertext_regx161x : DFFSNQ_X1 port map( D => reg_out_161_port, CLK => clk,
                           SN => n701, Q => Ciphertext(161));
   Ciphertext_regx67x : DFFSNQ_X1 port map( D => reg_out_67_port, CLK => clk, 
                           SN => n700, Q => Ciphertext(67));
   Ciphertext_regx48x : DFFSNQ_X1 port map( D => reg_out_48_port, CLK => clk, 
                           SN => n699, Q => Ciphertext(48));
   reg_in_regx80x : DFFRNQ_X1 port map( D => Plaintext(80), CLK => clk, RN => 
                           n697, Q => reg_in_80_port);
   reg_key_regx14x : DFFRNQ_X1 port map( D => Key(14), CLK => clk, RN => n696, 
                           Q => reg_key_14_port);
   reg_in_regx185x : DFFRNQ_X1 port map( D => Plaintext(185), CLK => clk, RN =>
                           n695, Q => reg_in_185_port);
   Ciphertext_regx168x : DFFRNQ_X1 port map( D => reg_out_168_port, CLK => clk,
                           RN => n694, Q => Ciphertext(168));
   n694 <= '1';
   n695 <= '1';
   n696 <= '1';
   n697 <= '1';
   n699 <= '1';
   n700 <= '1';
   n701 <= '1';
   SPEEDY_instance : SPEEDY_Rounds6_0 port map( Plaintext(191) => 
                           reg_in_191_port, Plaintext(190) => reg_in_190_port, 
                           Plaintext(189) => reg_in_189_port, Plaintext(188) =>
                           reg_in_188_port, Plaintext(187) => reg_in_187_port, 
                           Plaintext(186) => reg_in_186_port, Plaintext(185) =>
                           reg_in_185_port, Plaintext(184) => reg_in_184_port, 
                           Plaintext(183) => reg_in_183_port, Plaintext(182) =>
                           reg_in_182_port, Plaintext(181) => reg_in_181_port, 
                           Plaintext(180) => reg_in_180_port, Plaintext(179) =>
                           reg_in_179_port, Plaintext(178) => reg_in_178_port, 
                           Plaintext(177) => reg_in_177_port, Plaintext(176) =>
                           reg_in_176_port, Plaintext(175) => reg_in_175_port, 
                           Plaintext(174) => reg_in_174_port, Plaintext(173) =>
                           reg_in_173_port, Plaintext(172) => reg_in_172_port, 
                           Plaintext(171) => reg_in_171_port, Plaintext(170) =>
                           reg_in_170_port, Plaintext(169) => reg_in_169_port, 
                           Plaintext(168) => reg_in_168_port, Plaintext(167) =>
                           reg_in_167_port, Plaintext(166) => reg_in_166_port, 
                           Plaintext(165) => reg_in_165_port, Plaintext(164) =>
                           reg_in_164_port, Plaintext(163) => reg_in_163_port, 
                           Plaintext(162) => reg_in_162_port, Plaintext(161) =>
                           reg_in_161_port, Plaintext(160) => reg_in_160_port, 
                           Plaintext(159) => reg_in_159_port, Plaintext(158) =>
                           reg_in_158_port, Plaintext(157) => reg_in_157_port, 
                           Plaintext(156) => reg_in_156_port, Plaintext(155) =>
                           reg_in_155_port, Plaintext(154) => reg_in_154_port, 
                           Plaintext(153) => reg_in_153_port, Plaintext(152) =>
                           reg_in_152_port, Plaintext(151) => reg_in_151_port, 
                           Plaintext(150) => reg_in_150_port, Plaintext(149) =>
                           reg_in_149_port, Plaintext(148) => reg_in_148_port, 
                           Plaintext(147) => reg_in_147_port, Plaintext(146) =>
                           reg_in_146_port, Plaintext(145) => reg_in_145_port, 
                           Plaintext(144) => reg_in_144_port, Plaintext(143) =>
                           reg_in_143_port, Plaintext(142) => reg_in_142_port, 
                           Plaintext(141) => reg_in_141_port, Plaintext(140) =>
                           reg_in_140_port, Plaintext(139) => reg_in_139_port, 
                           Plaintext(138) => reg_in_138_port, Plaintext(137) =>
                           reg_in_137_port, Plaintext(136) => reg_in_136_port, 
                           Plaintext(135) => reg_in_135_port, Plaintext(134) =>
                           reg_in_134_port, Plaintext(133) => reg_in_133_port, 
                           Plaintext(132) => reg_in_132_port, Plaintext(131) =>
                           reg_in_131_port, Plaintext(130) => reg_in_130_port, 
                           Plaintext(129) => reg_in_129_port, Plaintext(128) =>
                           reg_in_128_port, Plaintext(127) => reg_in_127_port, 
                           Plaintext(126) => reg_in_126_port, Plaintext(125) =>
                           reg_in_125_port, Plaintext(124) => reg_in_124_port, 
                           Plaintext(123) => reg_in_123_port, Plaintext(122) =>
                           reg_in_122_port, Plaintext(121) => reg_in_121_port, 
                           Plaintext(120) => reg_in_120_port, Plaintext(119) =>
                           reg_in_119_port, Plaintext(118) => reg_in_118_port, 
                           Plaintext(117) => reg_in_117_port, Plaintext(116) =>
                           reg_in_116_port, Plaintext(115) => reg_in_115_port, 
                           Plaintext(114) => reg_in_114_port, Plaintext(113) =>
                           reg_in_113_port, Plaintext(112) => reg_in_112_port, 
                           Plaintext(111) => reg_in_111_port, Plaintext(110) =>
                           reg_in_110_port, Plaintext(109) => reg_in_109_port, 
                           Plaintext(108) => reg_in_108_port, Plaintext(107) =>
                           reg_in_107_port, Plaintext(106) => reg_in_106_port, 
                           Plaintext(105) => reg_in_105_port, Plaintext(104) =>
                           reg_in_104_port, Plaintext(103) => reg_in_103_port, 
                           Plaintext(102) => reg_in_102_port, Plaintext(101) =>
                           reg_in_101_port, Plaintext(100) => reg_in_100_port, 
                           Plaintext(99) => reg_in_99_port, Plaintext(98) => 
                           reg_in_98_port, Plaintext(97) => reg_in_97_port, 
                           Plaintext(96) => reg_in_96_port, Plaintext(95) => 
                           reg_in_95_port, Plaintext(94) => reg_in_94_port, 
                           Plaintext(93) => reg_in_93_port, Plaintext(92) => 
                           reg_in_92_port, Plaintext(91) => reg_in_91_port, 
                           Plaintext(90) => reg_in_90_port, Plaintext(89) => 
                           reg_in_89_port, Plaintext(88) => reg_in_88_port, 
                           Plaintext(87) => reg_in_87_port, Plaintext(86) => 
                           reg_in_86_port, Plaintext(85) => reg_in_85_port, 
                           Plaintext(84) => reg_in_84_port, Plaintext(83) => 
                           reg_in_83_port, Plaintext(82) => reg_in_82_port, 
                           Plaintext(81) => reg_in_81_port, Plaintext(80) => 
                           reg_in_80_port, Plaintext(79) => reg_in_79_port, 
                           Plaintext(78) => reg_in_78_port, Plaintext(77) => 
                           reg_in_77_port, Plaintext(76) => reg_in_76_port, 
                           Plaintext(75) => reg_in_75_port, Plaintext(74) => 
                           reg_in_74_port, Plaintext(73) => reg_in_73_port, 
                           Plaintext(72) => reg_in_72_port, Plaintext(71) => 
                           reg_in_71_port, Plaintext(70) => reg_in_70_port, 
                           Plaintext(69) => reg_in_69_port, Plaintext(68) => 
                           reg_in_68_port, Plaintext(67) => reg_in_67_port, 
                           Plaintext(66) => reg_in_66_port, Plaintext(65) => 
                           reg_in_65_port, Plaintext(64) => reg_in_64_port, 
                           Plaintext(63) => reg_in_63_port, Plaintext(62) => 
                           reg_in_62_port, Plaintext(61) => reg_in_61_port, 
                           Plaintext(60) => reg_in_60_port, Plaintext(59) => 
                           reg_in_59_port, Plaintext(58) => reg_in_58_port, 
                           Plaintext(57) => reg_in_57_port, Plaintext(56) => 
                           reg_in_56_port, Plaintext(55) => reg_in_55_port, 
                           Plaintext(54) => reg_in_54_port, Plaintext(53) => 
                           reg_in_53_port, Plaintext(52) => reg_in_52_port, 
                           Plaintext(51) => reg_in_51_port, Plaintext(50) => 
                           reg_in_50_port, Plaintext(49) => reg_in_49_port, 
                           Plaintext(48) => reg_in_48_port, Plaintext(47) => 
                           reg_in_47_port, Plaintext(46) => reg_in_46_port, 
                           Plaintext(45) => reg_in_45_port, Plaintext(44) => 
                           reg_in_44_port, Plaintext(43) => reg_in_43_port, 
                           Plaintext(42) => reg_in_42_port, Plaintext(41) => 
                           reg_in_41_port, Plaintext(40) => reg_in_40_port, 
                           Plaintext(39) => reg_in_39_port, Plaintext(38) => 
                           reg_in_38_port, Plaintext(37) => reg_in_37_port, 
                           Plaintext(36) => reg_in_36_port, Plaintext(35) => 
                           reg_in_35_port, Plaintext(34) => reg_in_34_port, 
                           Plaintext(33) => reg_in_33_port, Plaintext(32) => 
                           reg_in_32_port, Plaintext(31) => reg_in_31_port, 
                           Plaintext(30) => reg_in_30_port, Plaintext(29) => 
                           reg_in_29_port, Plaintext(28) => reg_in_28_port, 
                           Plaintext(27) => reg_in_27_port, Plaintext(26) => 
                           reg_in_26_port, Plaintext(25) => reg_in_25_port, 
                           Plaintext(24) => reg_in_24_port, Plaintext(23) => 
                           reg_in_23_port, Plaintext(22) => reg_in_22_port, 
                           Plaintext(21) => reg_in_21_port, Plaintext(20) => 
                           reg_in_20_port, Plaintext(19) => reg_in_19_port, 
                           Plaintext(18) => reg_in_18_port, Plaintext(17) => 
                           reg_in_17_port, Plaintext(16) => reg_in_16_port, 
                           Plaintext(15) => reg_in_15_port, Plaintext(14) => 
                           reg_in_14_port, Plaintext(13) => reg_in_13_port, 
                           Plaintext(12) => reg_in_12_port, Plaintext(11) => 
                           reg_in_11_port, Plaintext(10) => reg_in_10_port, 
                           Plaintext(9) => reg_in_9_port, Plaintext(8) => 
                           reg_in_8_port, Plaintext(7) => reg_in_7_port, 
                           Plaintext(6) => reg_in_6_port, Plaintext(5) => 
                           reg_in_5_port, Plaintext(4) => reg_in_4_port, 
                           Plaintext(3) => reg_in_3_port, Plaintext(2) => 
                           reg_in_2_port, Plaintext(1) => reg_in_1_port, 
                           Plaintext(0) => reg_in_0_port, Key(191) => 
                           reg_key_191_port, Key(190) => reg_key_190_port, 
                           Key(189) => reg_key_189_port, Key(188) => 
                           reg_key_188_port, Key(187) => reg_key_187_port, 
                           Key(186) => reg_key_186_port, Key(185) => 
                           reg_key_185_port, Key(184) => reg_key_184_port, 
                           Key(183) => reg_key_183_port, Key(182) => 
                           reg_key_182_port, Key(181) => reg_key_181_port, 
                           Key(180) => reg_key_180_port, Key(179) => 
                           reg_key_179_port, Key(178) => reg_key_178_port, 
                           Key(177) => reg_key_177_port, Key(176) => 
                           reg_key_176_port, Key(175) => reg_key_175_port, 
                           Key(174) => reg_key_174_port, Key(173) => 
                           reg_key_173_port, Key(172) => reg_key_172_port, 
                           Key(171) => reg_key_171_port, Key(170) => 
                           reg_key_170_port, Key(169) => reg_key_169_port, 
                           Key(168) => reg_key_168_port, Key(167) => 
                           reg_key_167_port, Key(166) => reg_key_166_port, 
                           Key(165) => reg_key_165_port, Key(164) => 
                           reg_key_164_port, Key(163) => reg_key_163_port, 
                           Key(162) => reg_key_162_port, Key(161) => 
                           reg_key_161_port, Key(160) => reg_key_160_port, 
                           Key(159) => reg_key_159_port, Key(158) => 
                           reg_key_158_port, Key(157) => reg_key_157_port, 
                           Key(156) => reg_key_156_port, Key(155) => 
                           reg_key_155_port, Key(154) => reg_key_154_port, 
                           Key(153) => reg_key_153_port, Key(152) => 
                           reg_key_152_port, Key(151) => reg_key_151_port, 
                           Key(150) => reg_key_150_port, Key(149) => 
                           reg_key_149_port, Key(148) => reg_key_148_port, 
                           Key(147) => reg_key_147_port, Key(146) => 
                           reg_key_146_port, Key(145) => reg_key_145_port, 
                           Key(144) => reg_key_144_port, Key(143) => 
                           reg_key_143_port, Key(142) => reg_key_142_port, 
                           Key(141) => reg_key_141_port, Key(140) => 
                           reg_key_140_port, Key(139) => reg_key_139_port, 
                           Key(138) => reg_key_138_port, Key(137) => 
                           reg_key_137_port, Key(136) => reg_key_136_port, 
                           Key(135) => reg_key_135_port, Key(134) => 
                           reg_key_134_port, Key(133) => reg_key_133_port, 
                           Key(132) => reg_key_132_port, Key(131) => 
                           reg_key_131_port, Key(130) => reg_key_130_port, 
                           Key(129) => reg_key_129_port, Key(128) => 
                           reg_key_128_port, Key(127) => reg_key_127_port, 
                           Key(126) => reg_key_126_port, Key(125) => 
                           reg_key_125_port, Key(124) => reg_key_124_port, 
                           Key(123) => reg_key_123_port, Key(122) => 
                           reg_key_122_port, Key(121) => reg_key_121_port, 
                           Key(120) => reg_key_120_port, Key(119) => 
                           reg_key_119_port, Key(118) => reg_key_118_port, 
                           Key(117) => reg_key_117_port, Key(116) => 
                           reg_key_116_port, Key(115) => reg_key_115_port, 
                           Key(114) => reg_key_114_port, Key(113) => 
                           reg_key_113_port, Key(112) => reg_key_112_port, 
                           Key(111) => reg_key_111_port, Key(110) => 
                           reg_key_110_port, Key(109) => reg_key_109_port, 
                           Key(108) => reg_key_108_port, Key(107) => 
                           reg_key_107_port, Key(106) => reg_key_106_port, 
                           Key(105) => reg_key_105_port, Key(104) => 
                           reg_key_104_port, Key(103) => reg_key_103_port, 
                           Key(102) => reg_key_102_port, Key(101) => 
                           reg_key_101_port, Key(100) => reg_key_100_port, 
                           Key(99) => reg_key_99_port, Key(98) => 
                           reg_key_98_port, Key(97) => reg_key_97_port, Key(96)
                           => reg_key_96_port, Key(95) => reg_key_95_port, 
                           Key(94) => reg_key_94_port, Key(93) => 
                           reg_key_93_port, Key(92) => reg_key_92_port, Key(91)
                           => reg_key_91_port, Key(90) => reg_key_90_port, 
                           Key(89) => reg_key_89_port, Key(88) => 
                           reg_key_88_port, Key(87) => reg_key_87_port, Key(86)
                           => reg_key_86_port, Key(85) => reg_key_85_port, 
                           Key(84) => reg_key_84_port, Key(83) => 
                           reg_key_83_port, Key(82) => reg_key_82_port, Key(81)
                           => reg_key_81_port, Key(80) => reg_key_80_port, 
                           Key(79) => reg_key_79_port, Key(78) => 
                           reg_key_78_port, Key(77) => reg_key_77_port, Key(76)
                           => reg_key_76_port, Key(75) => reg_key_75_port, 
                           Key(74) => reg_key_74_port, Key(73) => 
                           reg_key_73_port, Key(72) => reg_key_72_port, Key(71)
                           => reg_key_71_port, Key(70) => reg_key_70_port, 
                           Key(69) => reg_key_69_port, Key(68) => 
                           reg_key_68_port, Key(67) => reg_key_67_port, Key(66)
                           => reg_key_66_port, Key(65) => reg_key_65_port, 
                           Key(64) => reg_key_64_port, Key(63) => 
                           reg_key_63_port, Key(62) => reg_key_62_port, Key(61)
                           => reg_key_61_port, Key(60) => reg_key_60_port, 
                           Key(59) => reg_key_59_port, Key(58) => 
                           reg_key_58_port, Key(57) => reg_key_57_port, Key(56)
                           => reg_key_56_port, Key(55) => reg_key_55_port, 
                           Key(54) => reg_key_54_port, Key(53) => 
                           reg_key_53_port, Key(52) => reg_key_52_port, Key(51)
                           => reg_key_51_port, Key(50) => reg_key_50_port, 
                           Key(49) => reg_key_49_port, Key(48) => 
                           reg_key_48_port, Key(47) => reg_key_47_port, Key(46)
                           => reg_key_46_port, Key(45) => reg_key_45_port, 
                           Key(44) => reg_key_44_port, Key(43) => 
                           reg_key_43_port, Key(42) => reg_key_42_port, Key(41)
                           => reg_key_41_port, Key(40) => reg_key_40_port, 
                           Key(39) => reg_key_39_port, Key(38) => 
                           reg_key_38_port, Key(37) => reg_key_37_port, Key(36)
                           => reg_key_36_port, Key(35) => reg_key_35_port, 
                           Key(34) => reg_key_34_port, Key(33) => 
                           reg_key_33_port, Key(32) => reg_key_32_port, Key(31)
                           => reg_key_31_port, Key(30) => reg_key_30_port, 
                           Key(29) => reg_key_29_port, Key(28) => 
                           reg_key_28_port, Key(27) => reg_key_27_port, Key(26)
                           => reg_key_26_port, Key(25) => reg_key_25_port, 
                           Key(24) => reg_key_24_port, Key(23) => 
                           reg_key_23_port, Key(22) => reg_key_22_port, Key(21)
                           => reg_key_21_port, Key(20) => reg_key_20_port, 
                           Key(19) => reg_key_19_port, Key(18) => 
                           reg_key_18_port, Key(17) => reg_key_17_port, Key(16)
                           => reg_key_16_port, Key(15) => reg_key_15_port, 
                           Key(14) => reg_key_14_port, Key(13) => 
                           reg_key_13_port, Key(12) => reg_key_12_port, Key(11)
                           => reg_key_11_port, Key(10) => reg_key_10_port, 
                           Key(9) => reg_key_9_port, Key(8) => reg_key_8_port, 
                           Key(7) => reg_key_7_port, Key(6) => reg_key_6_port, 
                           Key(5) => reg_key_5_port, Key(4) => reg_key_4_port, 
                           Key(3) => reg_key_3_port, Key(2) => reg_key_2_port, 
                           Key(1) => reg_key_1_port, Key(0) => reg_key_0_port, 
                           Ciphertext(191) => reg_out_191_port, Ciphertext(190)
                           => reg_out_190_port, Ciphertext(189) => 
                           reg_out_189_port, Ciphertext(188) => 
                           reg_out_188_port, Ciphertext(187) => 
                           reg_out_187_port, Ciphertext(186) => 
                           reg_out_186_port, Ciphertext(185) => 
                           reg_out_185_port, Ciphertext(184) => 
                           reg_out_184_port, Ciphertext(183) => 
                           reg_out_183_port, Ciphertext(182) => 
                           reg_out_182_port, Ciphertext(181) => 
                           reg_out_181_port, Ciphertext(180) => 
                           reg_out_180_port, Ciphertext(179) => 
                           reg_out_179_port, Ciphertext(178) => 
                           reg_out_178_port, Ciphertext(177) => 
                           reg_out_177_port, Ciphertext(176) => 
                           reg_out_176_port, Ciphertext(175) => 
                           reg_out_175_port, Ciphertext(174) => 
                           reg_out_174_port, Ciphertext(173) => 
                           reg_out_173_port, Ciphertext(172) => 
                           reg_out_172_port, Ciphertext(171) => 
                           reg_out_171_port, Ciphertext(170) => 
                           reg_out_170_port, Ciphertext(169) => 
                           reg_out_169_port, Ciphertext(168) => 
                           reg_out_168_port, Ciphertext(167) => 
                           reg_out_167_port, Ciphertext(166) => 
                           reg_out_166_port, Ciphertext(165) => 
                           reg_out_165_port, Ciphertext(164) => 
                           reg_out_164_port, Ciphertext(163) => 
                           reg_out_163_port, Ciphertext(162) => 
                           reg_out_162_port, Ciphertext(161) => 
                           reg_out_161_port, Ciphertext(160) => 
                           reg_out_160_port, Ciphertext(159) => 
                           reg_out_159_port, Ciphertext(158) => 
                           reg_out_158_port, Ciphertext(157) => 
                           reg_out_157_port, Ciphertext(156) => 
                           reg_out_156_port, Ciphertext(155) => 
                           reg_out_155_port, Ciphertext(154) => 
                           reg_out_154_port, Ciphertext(153) => 
                           reg_out_153_port, Ciphertext(152) => 
                           reg_out_152_port, Ciphertext(151) => 
                           reg_out_151_port, Ciphertext(150) => 
                           reg_out_150_port, Ciphertext(149) => 
                           reg_out_149_port, Ciphertext(148) => 
                           reg_out_148_port, Ciphertext(147) => 
                           reg_out_147_port, Ciphertext(146) => 
                           reg_out_146_port, Ciphertext(145) => 
                           reg_out_145_port, Ciphertext(144) => 
                           reg_out_144_port, Ciphertext(143) => 
                           reg_out_143_port, Ciphertext(142) => 
                           reg_out_142_port, Ciphertext(141) => 
                           reg_out_141_port, Ciphertext(140) => 
                           reg_out_140_port, Ciphertext(139) => 
                           reg_out_139_port, Ciphertext(138) => 
                           reg_out_138_port, Ciphertext(137) => 
                           reg_out_137_port, Ciphertext(136) => 
                           reg_out_136_port, Ciphertext(135) => 
                           reg_out_135_port, Ciphertext(134) => 
                           reg_out_134_port, Ciphertext(133) => 
                           reg_out_133_port, Ciphertext(132) => 
                           reg_out_132_port, Ciphertext(131) => 
                           reg_out_131_port, Ciphertext(130) => 
                           reg_out_130_port, Ciphertext(129) => 
                           reg_out_129_port, Ciphertext(128) => 
                           reg_out_128_port, Ciphertext(127) => 
                           reg_out_127_port, Ciphertext(126) => 
                           reg_out_126_port, Ciphertext(125) => 
                           reg_out_125_port, Ciphertext(124) => 
                           reg_out_124_port, Ciphertext(123) => 
                           reg_out_123_port, Ciphertext(122) => 
                           reg_out_122_port, Ciphertext(121) => 
                           reg_out_121_port, Ciphertext(120) => 
                           reg_out_120_port, Ciphertext(119) => 
                           reg_out_119_port, Ciphertext(118) => 
                           reg_out_118_port, Ciphertext(117) => 
                           reg_out_117_port, Ciphertext(116) => 
                           reg_out_116_port, Ciphertext(115) => 
                           reg_out_115_port, Ciphertext(114) => 
                           reg_out_114_port, Ciphertext(113) => 
                           reg_out_113_port, Ciphertext(112) => 
                           reg_out_112_port, Ciphertext(111) => 
                           reg_out_111_port, Ciphertext(110) => 
                           reg_out_110_port, Ciphertext(109) => 
                           reg_out_109_port, Ciphertext(108) => 
                           reg_out_108_port, Ciphertext(107) => 
                           reg_out_107_port, Ciphertext(106) => 
                           reg_out_106_port, Ciphertext(105) => 
                           reg_out_105_port, Ciphertext(104) => 
                           reg_out_104_port, Ciphertext(103) => 
                           reg_out_103_port, Ciphertext(102) => 
                           reg_out_102_port, Ciphertext(101) => 
                           reg_out_101_port, Ciphertext(100) => 
                           reg_out_100_port, Ciphertext(99) => reg_out_99_port,
                           Ciphertext(98) => reg_out_98_port, Ciphertext(97) =>
                           reg_out_97_port, Ciphertext(96) => reg_out_96_port, 
                           Ciphertext(95) => reg_out_95_port, Ciphertext(94) =>
                           reg_out_94_port, Ciphertext(93) => reg_out_93_port, 
                           Ciphertext(92) => reg_out_92_port, Ciphertext(91) =>
                           reg_out_91_port, Ciphertext(90) => reg_out_90_port, 
                           Ciphertext(89) => reg_out_89_port, Ciphertext(88) =>
                           reg_out_88_port, Ciphertext(87) => reg_out_87_port, 
                           Ciphertext(86) => reg_out_86_port, Ciphertext(85) =>
                           reg_out_85_port, Ciphertext(84) => reg_out_84_port, 
                           Ciphertext(83) => reg_out_83_port, Ciphertext(82) =>
                           reg_out_82_port, Ciphertext(81) => reg_out_81_port, 
                           Ciphertext(80) => reg_out_80_port, Ciphertext(79) =>
                           reg_out_79_port, Ciphertext(78) => reg_out_78_port, 
                           Ciphertext(77) => reg_out_77_port, Ciphertext(76) =>
                           reg_out_76_port, Ciphertext(75) => reg_out_75_port, 
                           Ciphertext(74) => reg_out_74_port, Ciphertext(73) =>
                           reg_out_73_port, Ciphertext(72) => reg_out_72_port, 
                           Ciphertext(71) => reg_out_71_port, Ciphertext(70) =>
                           reg_out_70_port, Ciphertext(69) => reg_out_69_port, 
                           Ciphertext(68) => reg_out_68_port, Ciphertext(67) =>
                           reg_out_67_port, Ciphertext(66) => reg_out_66_port, 
                           Ciphertext(65) => reg_out_65_port, Ciphertext(64) =>
                           reg_out_64_port, Ciphertext(63) => reg_out_63_port, 
                           Ciphertext(62) => reg_out_62_port, Ciphertext(61) =>
                           reg_out_61_port, Ciphertext(60) => reg_out_60_port, 
                           Ciphertext(59) => reg_out_59_port, Ciphertext(58) =>
                           reg_out_58_port, Ciphertext(57) => reg_out_57_port, 
                           Ciphertext(56) => reg_out_56_port, Ciphertext(55) =>
                           reg_out_55_port, Ciphertext(54) => reg_out_54_port, 
                           Ciphertext(53) => reg_out_53_port, Ciphertext(52) =>
                           reg_out_52_port, Ciphertext(51) => reg_out_51_port, 
                           Ciphertext(50) => reg_out_50_port, Ciphertext(49) =>
                           reg_out_49_port, Ciphertext(48) => reg_out_48_port, 
                           Ciphertext(47) => reg_out_47_port, Ciphertext(46) =>
                           reg_out_46_port, Ciphertext(45) => reg_out_45_port, 
                           Ciphertext(44) => reg_out_44_port, Ciphertext(43) =>
                           reg_out_43_port, Ciphertext(42) => reg_out_42_port, 
                           Ciphertext(41) => reg_out_41_port, Ciphertext(40) =>
                           reg_out_40_port, Ciphertext(39) => reg_out_39_port, 
                           Ciphertext(38) => reg_out_38_port, Ciphertext(37) =>
                           reg_out_37_port, Ciphertext(36) => reg_out_36_port, 
                           Ciphertext(35) => reg_out_35_port, Ciphertext(34) =>
                           reg_out_34_port, Ciphertext(33) => reg_out_33_port, 
                           Ciphertext(32) => reg_out_32_port, Ciphertext(31) =>
                           reg_out_31_port, Ciphertext(30) => reg_out_30_port, 
                           Ciphertext(29) => reg_out_29_port, Ciphertext(28) =>
                           reg_out_28_port, Ciphertext(27) => reg_out_27_port, 
                           Ciphertext(26) => reg_out_26_port, Ciphertext(25) =>
                           reg_out_25_port, Ciphertext(24) => reg_out_24_port, 
                           Ciphertext(23) => reg_out_23_port, Ciphertext(22) =>
                           reg_out_22_port, Ciphertext(21) => reg_out_21_port, 
                           Ciphertext(20) => reg_out_20_port, Ciphertext(19) =>
                           reg_out_19_port, Ciphertext(18) => reg_out_18_port, 
                           Ciphertext(17) => reg_out_17_port, Ciphertext(16) =>
                           reg_out_16_port, Ciphertext(15) => reg_out_15_port, 
                           Ciphertext(14) => reg_out_14_port, Ciphertext(13) =>
                           reg_out_13_port, Ciphertext(12) => reg_out_12_port, 
                           Ciphertext(11) => reg_out_11_port, Ciphertext(10) =>
                           reg_out_10_port, Ciphertext(9) => reg_out_9_port, 
                           Ciphertext(8) => reg_out_8_port, Ciphertext(7) => 
                           reg_out_7_port, Ciphertext(6) => reg_out_6_port, 
                           Ciphertext(5) => reg_out_5_port, Ciphertext(4) => 
                           reg_out_4_port, Ciphertext(3) => reg_out_3_port, 
                           Ciphertext(2) => reg_out_2_port, Ciphertext(1) => 
                           reg_out_1_port, Ciphertext(0) => reg_out_0_port);
   Ciphertext_regx186x : DFFRNQ_X1 port map( D => reg_out_186_port, CLK => clk,
                           RN => n711, Q => Ciphertext(186));
   Ciphertext_regx147x : DFFRNQ_X1 port map( D => reg_out_147_port, CLK => clk,
                           RN => n710, Q => Ciphertext(147));
   Ciphertext_regx21x : DFFRNQ_X1 port map( D => reg_out_21_port, CLK => clk, 
                           RN => n709, Q => Ciphertext(21));
   reg_key_regx8x : DFFSNQ_X1 port map( D => Key(8), CLK => clk, SN => n708, Q 
                           => reg_key_8_port);
   reg_in_regx111x : DFFRNQ_X1 port map( D => Plaintext(111), CLK => clk, RN =>
                           n707, Q => reg_in_111_port);
   Ciphertext_regx100x : DFFSNQ_X1 port map( D => reg_out_100_port, CLK => clk,
                           SN => n706, Q => Ciphertext(100));
   Ciphertext_regx51x : DFFRNQ_X1 port map( D => reg_out_51_port, CLK => clk, 
                           RN => n705, Q => Ciphertext(51));
   Ciphertext_regx159x : DFFSNQ_X1 port map( D => reg_out_159_port, CLK => clk,
                           SN => n704, Q => Ciphertext(159));
   Ciphertext_regx171x : DFFRNQ_X1 port map( D => reg_out_171_port, CLK => clk,
                           RN => n703, Q => Ciphertext(171));
   reg_in_regx83x : DFFRNQ_X1 port map( D => Plaintext(83), CLK => clk, RN => 
                           n702, Q => reg_in_83_port);
   n702 <= '1';
   n703 <= '1';
   n704 <= '1';
   n705 <= '1';
   n706 <= '1';
   n707 <= '1';
   n708 <= '1';
   n709 <= '1';
   n710 <= '1';
   n711 <= '1';

end SYN_Behavioral;
